

module b17_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P1_MEMORYFETCH_REG_SCAN_IN, 
        DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, 
        DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, 
        DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, 
        DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, 
        DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, 
        DATAI_0_, HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_,
         DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_,
         DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_,
         DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_,
         DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_,
         DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_,
         HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN,
         P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN,
         P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN,
         P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN,
         P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN,
         P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN,
         P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN,
         P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN,
         P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN,
         P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN,
         P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN,
         P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN,
         P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN,
         P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN,
         P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN,
         P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN,
         P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN,
         P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN,
         P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN,
         P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN,
         P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN,
         P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN,
         P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN,
         P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN,
         P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN,
         P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN,
         P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN,
         P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN,
         P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN,
         P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN,
         P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN,
         P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN,
         P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN,
         P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN,
         P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN,
         P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN,
         P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN,
         P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN,
         P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN,
         P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN,
         P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN,
         P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN,
         P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN,
         P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN,
         P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN,
         P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN,
         P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN,
         P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN,
         P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN,
         P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN,
         P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11012, n11013, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
         n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
         n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
         n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
         n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
         n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
         n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
         n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
         n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
         n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479,
         n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
         n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495,
         n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503,
         n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
         n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
         n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
         n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543,
         n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551,
         n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
         n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567,
         n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575,
         n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
         n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
         n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
         n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607,
         n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
         n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623,
         n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
         n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
         n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
         n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
         n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
         n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
         n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
         n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
         n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
         n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
         n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719,
         n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
         n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735,
         n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743,
         n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751,
         n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
         n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
         n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
         n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783,
         n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791,
         n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807,
         n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815,
         n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823,
         n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831,
         n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839,
         n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
         n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855,
         n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863,
         n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871,
         n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879,
         n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887,
         n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895,
         n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903,
         n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911,
         n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919,
         n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927,
         n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935,
         n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943,
         n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951,
         n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959,
         n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967,
         n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975,
         n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983,
         n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991,
         n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999,
         n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007,
         n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015,
         n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023,
         n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031,
         n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039,
         n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047,
         n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055,
         n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063,
         n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071,
         n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079,
         n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087,
         n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095,
         n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103,
         n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
         n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119,
         n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127,
         n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135,
         n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143,
         n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151,
         n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159,
         n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167,
         n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175,
         n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
         n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191,
         n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199,
         n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
         n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215,
         n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223,
         n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231,
         n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239,
         n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247,
         n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255,
         n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263,
         n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271,
         n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
         n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287,
         n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295,
         n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303,
         n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311,
         n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319,
         n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327,
         n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335,
         n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343,
         n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
         n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359,
         n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367,
         n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375,
         n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383,
         n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391,
         n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399,
         n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
         n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415,
         n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
         n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431,
         n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439,
         n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447,
         n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455,
         n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463,
         n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471,
         n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479,
         n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487,
         n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
         n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503,
         n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511,
         n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519,
         n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527,
         n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535,
         n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543,
         n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551,
         n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559,
         n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567,
         n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575,
         n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583,
         n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591,
         n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599,
         n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607,
         n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615,
         n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623,
         n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631,
         n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639,
         n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647,
         n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655,
         n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663,
         n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671,
         n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679,
         n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687,
         n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695,
         n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703,
         n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
         n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719,
         n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727,
         n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735,
         n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743,
         n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751,
         n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759,
         n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767,
         n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775,
         n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
         n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791,
         n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799,
         n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807,
         n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
         n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823,
         n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831,
         n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839,
         n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847,
         n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855,
         n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863,
         n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871,
         n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879,
         n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887,
         n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895,
         n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903,
         n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911,
         n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919,
         n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927,
         n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935,
         n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943,
         n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951,
         n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959,
         n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967,
         n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975,
         n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983,
         n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991,
         n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999,
         n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007,
         n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015,
         n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023,
         n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031,
         n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039,
         n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047,
         n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,
         n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,
         n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,
         n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
         n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088,
         n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096,
         n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104,
         n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,
         n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
         n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
         n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,
         n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
         n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160,
         n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168,
         n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176,
         n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,
         n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,
         n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,
         n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
         n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,
         n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
         n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232,
         n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240,
         n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,
         n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,
         n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,
         n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272,
         n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
         n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,
         n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,
         n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304,
         n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312,
         n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,
         n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
         n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
         n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,
         n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
         n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,
         n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,
         n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,
         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,
         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,
         n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
         n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,
         n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,
         n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,
         n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528,
         n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,
         n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,
         n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,
         n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560,
         n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
         n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576,
         n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584,
         n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592,
         n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600,
         n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,
         n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,
         n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
         n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632,
         n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,
         n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648,
         n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,
         n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,
         n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672,
         n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680,
         n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
         n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696,
         n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704,
         n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,
         n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720,
         n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,
         n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736,
         n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,
         n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752,
         n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,
         n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,
         n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776,
         n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,
         n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,
         n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,
         n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,
         n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816,
         n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,
         n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,
         n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840,
         n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848,
         n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,
         n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,
         n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,
         n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,
         n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888,
         n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896,
         n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,
         n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,
         n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920,
         n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,
         n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,
         n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944,
         n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952,
         n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960,
         n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968,
         n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
         n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984,
         n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992,
         n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,
         n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008,
         n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,
         n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024,
         n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032,
         n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040,
         n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048,
         n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056,
         n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064,
         n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,
         n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080,
         n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
         n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096,
         n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104,
         n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112,
         n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,
         n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128,
         n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136,
         n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,
         n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152,
         n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160,
         n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168,
         n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176,
         n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184,
         n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192,
         n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200,
         n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208,
         n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216,
         n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224,
         n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232,
         n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240,
         n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248,
         n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256,
         n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264,
         n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272,
         n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280,
         n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288,
         n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296,
         n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304,
         n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312,
         n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320,
         n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328,
         n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336,
         n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344,
         n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352,
         n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360,
         n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368,
         n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376,
         n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384,
         n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392,
         n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400,
         n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408,
         n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416,
         n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424,
         n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432,
         n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440,
         n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448,
         n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456,
         n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464,
         n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472,
         n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480,
         n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488,
         n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496,
         n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504,
         n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512,
         n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520,
         n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528,
         n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536,
         n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544,
         n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552,
         n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560,
         n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568,
         n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,
         n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584,
         n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592,
         n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600,
         n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608,
         n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616,
         n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624,
         n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632,
         n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640,
         n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648,
         n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656,
         n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664,
         n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672,
         n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680,
         n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,
         n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,
         n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704,
         n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712,
         n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720,
         n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728,
         n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
         n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744,
         n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752,
         n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760,
         n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
         n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776,
         n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784,
         n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792,
         n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
         n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
         n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816,
         n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824,
         n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832,
         n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,
         n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848,
         n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856,
         n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864,
         n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872,
         n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880,
         n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888,
         n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896,
         n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,
         n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912,
         n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920,
         n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928,
         n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936,
         n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944,
         n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952,
         n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960,
         n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968,
         n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976,
         n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984,
         n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992,
         n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000,
         n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008,
         n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016,
         n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024,
         n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032,
         n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040,
         n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048,
         n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056,
         n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064,
         n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072,
         n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080,
         n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088,
         n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096,
         n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104,
         n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112,
         n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120,
         n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128,
         n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136,
         n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144,
         n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152,
         n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160,
         n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168,
         n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176,
         n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184,
         n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192,
         n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,
         n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208,
         n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216,
         n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224,
         n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232,
         n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240,
         n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248,
         n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256,
         n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264,
         n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
         n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280,
         n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288,
         n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296,
         n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304,
         n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312,
         n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320,
         n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328,
         n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336,
         n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344,
         n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352,
         n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360,
         n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368,
         n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376,
         n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384,
         n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392,
         n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400,
         n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408,
         n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416,
         n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424,
         n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432,
         n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440,
         n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448,
         n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456,
         n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464,
         n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472,
         n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480,
         n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488,
         n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496,
         n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504,
         n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512,
         n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520,
         n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528,
         n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536,
         n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544,
         n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552,
         n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560,
         n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568,
         n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576,
         n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,
         n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592,
         n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600,
         n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608,
         n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616,
         n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624,
         n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632,
         n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640,
         n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648,
         n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656,
         n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664,
         n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672,
         n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680,
         n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688,
         n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696,
         n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704,
         n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712,
         n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720,
         n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728,
         n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736,
         n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744,
         n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752,
         n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760,
         n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768,
         n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
         n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784,
         n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792,
         n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800,
         n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808,
         n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816,
         n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824,
         n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832,
         n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840,
         n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848,
         n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856,
         n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864,
         n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872,
         n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880,
         n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888,
         n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896,
         n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904,
         n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912,
         n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920,
         n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928,
         n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936,
         n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944,
         n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952,
         n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960,
         n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968,
         n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976,
         n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984,
         n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992,
         n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000,
         n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008,
         n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016,
         n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024,
         n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032,
         n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040,
         n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048,
         n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056,
         n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064,
         n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072,
         n21073, n21074, n21075, n21076, n21077, n21078, n21079, n21080,
         n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088,
         n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096,
         n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104,
         n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112,
         n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120,
         n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128,
         n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136,
         n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144,
         n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152,
         n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160,
         n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21168,
         n21169, n21170, n21171, n21172, n21173, n21174, n21175, n21176,
         n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184,
         n21185, n21186, n21187, n21188, n21189, n21190, n21191, n21192,
         n21193, n21194, n21195, n21196, n21197, n21198, n21199, n21200,
         n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208,
         n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216,
         n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224,
         n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232,
         n21233, n21234, n21235, n21236, n21237, n21238, n21239, n21240,
         n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248,
         n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256,
         n21257, n21258, n21259, n21260, n21261, n21262, n21263, n21264,
         n21265, n21266, n21267, n21268, n21269, n21270, n21271, n21272,
         n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280,
         n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288,
         n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296,
         n21297, n21298, n21299, n21300, n21301, n21302, n21303, n21304,
         n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312,
         n21313, n21314, n21315, n21316, n21317, n21318, n21319, n21320,
         n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328,
         n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336,
         n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344,
         n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352,
         n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360,
         n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368,
         n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376,
         n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384,
         n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392,
         n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400,
         n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408,
         n21409, n21410, n21411, n21412, n21413, n21414, n21415, n21416,
         n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424,
         n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432,
         n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440,
         n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448,
         n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456,
         n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464,
         n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472,
         n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480,
         n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488,
         n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496,
         n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504,
         n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512,
         n21513, n21514, n21515, n21516, n21517, n21518, n21519, n21520,
         n21521, n21522, n21523, n21524, n21525, n21526, n21527, n21528,
         n21529, n21530, n21531, n21532, n21533, n21534, n21535, n21536,
         n21537, n21538, n21539, n21540, n21541, n21542, n21543, n21544,
         n21545, n21546, n21547, n21548, n21549, n21550, n21551, n21552,
         n21553, n21554, n21555, n21556, n21557, n21558, n21559, n21560,
         n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568,
         n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576,
         n21577, n21578, n21579, n21580, n21581, n21582, n21583, n21584,
         n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592,
         n21593, n21594, n21595, n21596, n21597, n21598, n21599, n21600,
         n21601, n21602, n21603, n21604, n21605, n21606, n21607, n21608,
         n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616,
         n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624,
         n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632,
         n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640,
         n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648,
         n21649, n21650, n21651, n21652, n21653, n21654, n21655, n21656,
         n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664,
         n21665, n21666, n21667, n21668, n21669, n21670, n21671, n21672,
         n21673, n21674, n21675, n21676, n21677, n21678, n21679, n21680,
         n21681, n21682, n21683, n21684, n21685, n21686, n21687, n21688,
         n21689, n21690, n21691, n21692, n21693, n21694, n21695, n21696,
         n21697, n21698, n21699, n21700, n21701, n21702, n21703, n21704,
         n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712,
         n21713, n21714, n21715, n21716, n21717, n21718, n21719, n21720,
         n21721, n21722, n21723, n21724, n21725, n21726, n21727, n21728,
         n21729, n21730, n21731, n21732, n21733, n21734, n21735, n21736,
         n21737, n21738, n21739, n21740, n21741, n21742, n21743, n21744,
         n21745, n21746, n21747, n21748, n21749, n21750, n21751, n21752,
         n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760,
         n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768,
         n21769, n21770, n21771, n21772, n21773, n21774, n21775, n21776,
         n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784,
         n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792,
         n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21800,
         n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808,
         n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816,
         n21817, n21818, n21819, n21820, n21821, n21822, n21823, n21824,
         n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832,
         n21833, n21834, n21835, n21836, n21837, n21838, n21839, n21840,
         n21841, n21842, n21843, n21844, n21845, n21846, n21847, n21848,
         n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856,
         n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864,
         n21865, n21866, n21867, n21868, n21869, n21870, n21871, n21872,
         n21873, n21874, n21875, n21876, n21877, n21878, n21879, n21880,
         n21881, n21882, n21883, n21884, n21885, n21886, n21887, n21888,
         n21889, n21890, n21891, n21892, n21893, n21894, n21895, n21896,
         n21897, n21898, n21899, n21900, n21901, n21902, n21903, n21904,
         n21905, n21906, n21907, n21908, n21909, n21910, n21911, n21912,
         n21913, n21914, n21915, n21916, n21917, n21918, n21919, n21920,
         n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928,
         n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936,
         n21937, n21938, n21939, n21940, n21941, n21942, n21943, n21944,
         n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952,
         n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960,
         n21961, n21962, n21963, n21964, n21965, n21966, n21967, n21968,
         n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21976,
         n21977, n21978, n21979, n21980, n21981, n21982, n21983, n21984,
         n21985, n21986, n21987, n21988, n21989, n21990, n21991, n21992,
         n21993, n21994, n21995, n21996, n21997, n21998, n21999, n22000,
         n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008,
         n22009, n22010, n22011, n22012, n22013, n22014, n22015, n22016,
         n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024,
         n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032,
         n22033, n22034, n22035, n22036, n22037, n22038, n22039, n22040,
         n22041, n22042, n22043, n22044, n22045, n22046, n22047, n22048,
         n22049, n22050, n22051, n22052, n22053, n22054, n22055, n22056,
         n22057, n22058, n22059, n22060, n22061, n22062, n22063, n22064,
         n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072,
         n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080,
         n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088,
         n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096,
         n22097, n22098, n22099, n22100, n22101, n22102, n22103, n22104,
         n22105, n22106, n22107, n22108, n22109, n22110, n22111, n22112,
         n22113, n22114, n22115, n22116, n22117, n22118, n22119, n22120,
         n22121, n22122, n22123, n22124, n22125, n22126, n22127, n22128,
         n22129, n22130, n22131, n22132, n22133, n22134, n22135, n22136,
         n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144,
         n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152,
         n22153, n22154, n22155, n22156, n22157, n22158, n22159, n22160,
         n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168,
         n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176,
         n22177, n22178, n22179, n22180, n22181, n22182, n22183, n22184,
         n22185, n22186, n22187, n22188, n22189, n22190, n22191, n22192,
         n22193, n22194, n22195, n22196, n22197, n22198, n22199, n22200,
         n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22208,
         n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216,
         n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224,
         n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232,
         n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240,
         n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248,
         n22249, n22250, n22251, n22252, n22253, n22254, n22255, n22256,
         n22257, n22258, n22259, n22260, n22261, n22262, n22263, n22264,
         n22265, n22266, n22267, n22268, n22269, n22270, n22271, n22272,
         n22273, n22274, n22275, n22276, n22277, n22278, n22279, n22280,
         n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288,
         n22289, n22290, n22291, n22292, n22293, n22294, n22295, n22296,
         n22297, n22298, n22299, n22300, n22301, n22302, n22303, n22304,
         n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312,
         n22313, n22314, n22315, n22316, n22317, n22318, n22319, n22320,
         n22321, n22322, n22323, n22324, n22325, n22326, n22327, n22328,
         n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336,
         n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344,
         n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352,
         n22353, n22354, n22355, n22356, n22357, n22358, n22359, n22360,
         n22361, n22362, n22363, n22364, n22365, n22366, n22367, n22368,
         n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376,
         n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384,
         n22385, n22386, n22387, n22388, n22389, n22390, n22391, n22392,
         n22393, n22394, n22395, n22396, n22397, n22398, n22399, n22400,
         n22401;

  INV_X1 U11062 ( .A(n18297), .ZN(n18304) );
  OAI22_X1 U11063 ( .A1(n16660), .A2(n11177), .B1(n11180), .B2(n14440), .ZN(
        n16639) );
  AND2_X1 U11064 ( .A1(n14553), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n15942)
         );
  NOR2_X1 U11065 ( .A1(n18219), .A2(n21247), .ZN(n18218) );
  NAND2_X1 U11066 ( .A1(n14511), .A2(n14512), .ZN(n14510) );
  INV_X1 U11067 ( .A(n16382), .ZN(n20182) );
  OR2_X2 U11068 ( .A1(n16233), .A2(n16173), .ZN(n16175) );
  NAND2_X1 U11069 ( .A1(n15514), .A2(n15513), .ZN(n15512) );
  NAND2_X1 U11070 ( .A1(n12203), .A2(n11589), .ZN(n15520) );
  NAND2_X1 U11071 ( .A1(n18253), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n18296) );
  CLKBUF_X1 U11072 ( .A(n19793), .Z(n10959) );
  CLKBUF_X1 U11073 ( .A(n12979), .Z(n13070) );
  NOR3_X1 U11074 ( .A1(n11480), .A2(n11479), .A3(n11478), .ZN(n11506) );
  AND3_X1 U11075 ( .A1(n11482), .A2(n11487), .A3(n16033), .ZN(n19439) );
  OR2_X1 U11076 ( .A1(n11496), .A2(n11492), .ZN(n19447) );
  NAND2_X1 U11077 ( .A1(n18093), .A2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n18186) );
  OR2_X1 U11078 ( .A1(n12714), .A2(n12640), .ZN(n12667) );
  NAND2_X1 U11079 ( .A1(n11130), .A2(n11128), .ZN(n20502) );
  INV_X2 U11080 ( .A(n15053), .ZN(n17890) );
  NAND2_X1 U11081 ( .A1(n12666), .A2(n12838), .ZN(n13129) );
  CLKBUF_X2 U11082 ( .A(n13835), .Z(n18013) );
  CLKBUF_X3 U11083 ( .A(n13789), .Z(n18047) );
  BUF_X1 U11084 ( .A(n11427), .Z(n11832) );
  CLKBUF_X1 U11085 ( .A(n11916), .Z(n12181) );
  NOR2_X4 U11086 ( .A1(n21012), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13835) );
  CLKBUF_X1 U11087 ( .A(n13789), .Z(n10960) );
  CLKBUF_X1 U11088 ( .A(n13839), .Z(n17908) );
  CLKBUF_X2 U11089 ( .A(n13790), .Z(n18025) );
  CLKBUF_X1 U11090 ( .A(n13778), .Z(n18032) );
  AND2_X1 U11091 ( .A1(n15340), .A2(n11414), .ZN(n11461) );
  AND2_X1 U11092 ( .A1(n14453), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14253) );
  AND2_X2 U11093 ( .A1(n10962), .A2(n11374), .ZN(n14271) );
  INV_X2 U11094 ( .A(n15313), .ZN(n11394) );
  AND2_X1 U11095 ( .A1(n14303), .A2(n15283), .ZN(n14273) );
  INV_X1 U11096 ( .A(n11379), .ZN(n14099) );
  BUF_X1 U11097 ( .A(n12967), .Z(n15401) );
  AND2_X2 U11098 ( .A1(n12971), .A2(n12601), .ZN(n13074) );
  NOR2_X1 U11099 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11268) );
  NAND3_X1 U11100 ( .A1(n11208), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14477) );
  AND2_X1 U11101 ( .A1(n12454), .A2(n12455), .ZN(n12687) );
  AND4_X1 U11102 ( .A1(n11209), .A2(n12447), .A3(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A4(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12527) );
  AND2_X1 U11103 ( .A1(n11091), .A2(n15211), .ZN(n12686) );
  AND2_X1 U11104 ( .A1(n11091), .A2(n15213), .ZN(n12507) );
  INV_X1 U11105 ( .A(n12460), .ZN(n11021) );
  INV_X2 U11106 ( .A(n12460), .ZN(n12612) );
  AND2_X1 U11107 ( .A1(n11394), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11414) );
  CLKBUF_X2 U11109 ( .A(n12527), .Z(n13579) );
  NOR2_X1 U11110 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12455) );
  CLKBUF_X2 U11111 ( .A(n11366), .Z(n14481) );
  NOR2_X2 U11112 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11261) );
  INV_X1 U11113 ( .A(n14477), .ZN(n11341) );
  AND2_X1 U11114 ( .A1(n15211), .A2(n12455), .ZN(n12629) );
  AND4_X1 U11115 ( .A1(n12451), .A2(n12450), .A3(n12449), .A4(n12448), .ZN(
        n11257) );
  INV_X1 U11116 ( .A(n12460), .ZN(n11022) );
  AND2_X1 U11117 ( .A1(n14303), .A2(n11267), .ZN(n14288) );
  AND2_X1 U11118 ( .A1(n14303), .A2(n11261), .ZN(n14272) );
  INV_X1 U11119 ( .A(n14477), .ZN(n10961) );
  INV_X1 U11120 ( .A(n14477), .ZN(n10962) );
  BUF_X1 U11121 ( .A(n11365), .Z(n14480) );
  NAND2_X1 U11122 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21021) );
  NAND2_X1 U11123 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21006), .ZN(
        n13760) );
  NAND2_X2 U11124 ( .A1(n12972), .A2(n11020), .ZN(n13052) );
  NAND2_X1 U11125 ( .A1(n12840), .A2(n12839), .ZN(n12850) );
  AND2_X1 U11126 ( .A1(n11925), .A2(n11399), .ZN(n11934) );
  INV_X1 U11127 ( .A(n12202), .ZN(n13735) );
  INV_X1 U11128 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11374) );
  AOI21_X1 U11129 ( .B1(n14008), .B2(n13870), .A(n18371), .ZN(n18339) );
  NAND2_X1 U11131 ( .A1(n16145), .A2(n16215), .ZN(n16127) );
  NAND2_X1 U11132 ( .A1(n12682), .A2(n14890), .ZN(n22063) );
  OR2_X1 U11133 ( .A1(n18771), .A2(n18784), .ZN(n16613) );
  NAND2_X1 U11134 ( .A1(n12339), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12354) );
  AOI211_X1 U11136 ( .C1(n18876), .C2(n16044), .A(n16775), .B(n16043), .ZN(
        n16048) );
  INV_X2 U11137 ( .A(n12181), .ZN(n19633) );
  AND2_X1 U11138 ( .A1(n11126), .A2(n20592), .ZN(n11037) );
  INV_X1 U11139 ( .A(n20351), .ZN(n19216) );
  INV_X1 U11140 ( .A(n13074), .ZN(n14535) );
  NOR2_X2 U11141 ( .A1(n15925), .A2(n13021), .ZN(n16514) );
  BUF_X1 U11142 ( .A(n16103), .Z(n16114) );
  BUF_X1 U11143 ( .A(n16127), .Z(n16214) );
  INV_X1 U11144 ( .A(n12966), .ZN(n15178) );
  NAND2_X1 U11147 ( .A1(n15640), .A2(n15641), .ZN(n15642) );
  XNOR2_X1 U11148 ( .A(n13663), .B(n13662), .ZN(n16044) );
  OAI21_X1 U11149 ( .B1(n16787), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n16045), .ZN(n15992) );
  NAND2_X1 U11150 ( .A1(n15175), .A2(n13635), .ZN(n14744) );
  AOI22_X1 U11151 ( .A1(n21577), .A2(n21596), .B1(n21595), .B2(n21576), .ZN(
        n21584) );
  OR2_X1 U11152 ( .A1(n18917), .A2(n10959), .ZN(n17670) );
  INV_X1 U11153 ( .A(n18613), .ZN(n11489) );
  INV_X1 U11154 ( .A(n17850), .ZN(n10957) );
  INV_X1 U11155 ( .A(n13840), .ZN(n17850) );
  OR2_X1 U11156 ( .A1(n16517), .A2(n13033), .ZN(n10955) );
  BUF_X1 U11157 ( .A(n13908), .Z(n18049) );
  NAND2_X2 U11158 ( .A1(n15887), .A2(n11043), .ZN(n11103) );
  NOR2_X4 U11159 ( .A1(n20502), .A2(n20519), .ZN(n18100) );
  AOI211_X2 U11160 ( .C1(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n21748), .A(
        n13655), .B(n13654), .ZN(n13656) );
  OR2_X2 U11161 ( .A1(n12267), .A2(n12265), .ZN(n12262) );
  AND3_X4 U11162 ( .A1(n12483), .A2(n12482), .A3(n12481), .ZN(n12558) );
  AND2_X2 U11163 ( .A1(n12559), .A2(n12971), .ZN(n12952) );
  OR2_X2 U11164 ( .A1(n12471), .A2(n12470), .ZN(n12971) );
  AND2_X2 U11165 ( .A1(n12562), .A2(n12558), .ZN(n14810) );
  NOR2_X4 U11166 ( .A1(n18368), .A2(n21374), .ZN(n18312) );
  AND2_X2 U11167 ( .A1(n15735), .A2(n15749), .ZN(n15640) );
  NAND2_X2 U11169 ( .A1(n11704), .A2(n11664), .ZN(n11711) );
  NOR2_X2 U11170 ( .A1(n20343), .A2(n13758), .ZN(n13839) );
  NAND3_X2 U11172 ( .A1(n11036), .A2(n11275), .A3(n11096), .ZN(n12002) );
  BUF_X8 U11174 ( .A(n18049), .Z(n10956) );
  AND4_X2 U11175 ( .A1(n12497), .A2(n12496), .A3(n12495), .A4(n12494), .ZN(
        n11034) );
  NAND3_X2 U11176 ( .A1(n11459), .A2(n11458), .A3(n11457), .ZN(n11826) );
  NAND2_X2 U11177 ( .A1(n11117), .A2(n12727), .ZN(n12750) );
  NOR2_X1 U11178 ( .A1(n13759), .A2(n21021), .ZN(n13840) );
  NAND2_X2 U11181 ( .A1(n11257), .A2(n11255), .ZN(n14860) );
  OAI211_X1 U11182 ( .C1(n11832), .C2(n17662), .A(n11039), .B(n11417), .ZN(
        n11440) );
  AOI211_X2 U11183 ( .C1(n20192), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n20162), .B(n20161), .ZN(n20163) );
  NAND2_X2 U11184 ( .A1(n21001), .A2(n21020), .ZN(n20343) );
  AOI21_X2 U11185 ( .B1(n15512), .B2(n12230), .A(n11237), .ZN(n15766) );
  NOR2_X1 U11186 ( .A1(n13761), .A2(n13758), .ZN(n13789) );
  AND2_X4 U11187 ( .A1(n12883), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12454) );
  XNOR2_X2 U11189 ( .A(n11614), .B(n11615), .ZN(n15692) );
  NAND2_X2 U11190 ( .A1(n15520), .A2(n11591), .ZN(n11614) );
  INV_X1 U11191 ( .A(n10962), .ZN(n10963) );
  INV_X1 U11192 ( .A(n14477), .ZN(n14452) );
  NAND2_X2 U11193 ( .A1(n11203), .A2(n11202), .ZN(n11450) );
  NOR2_X2 U11194 ( .A1(n18452), .A2(n13852), .ZN(n21078) );
  NOR2_X1 U11195 ( .A1(n16889), .A2(n16877), .ZN(n16876) );
  CLKBUF_X1 U11196 ( .A(n16639), .Z(n16646) );
  OR2_X1 U11197 ( .A1(n20935), .A2(n20936), .ZN(n20937) );
  OR2_X1 U11198 ( .A1(n18224), .A2(n18258), .ZN(n18220) );
  NOR2_X1 U11199 ( .A1(n16614), .A2(n16613), .ZN(n16612) );
  OR2_X1 U11200 ( .A1(n16175), .A2(n16162), .ZN(n10973) );
  BUF_X1 U11201 ( .A(n18463), .Z(n11018) );
  NAND2_X1 U11202 ( .A1(n21475), .A2(n21446), .ZN(n21505) );
  INV_X2 U11203 ( .A(n21343), .ZN(n21437) );
  NAND2_X1 U11204 ( .A1(n14000), .A2(n21025), .ZN(n21003) );
  NOR2_X1 U11205 ( .A1(n12246), .A2(n12245), .ZN(n12247) );
  INV_X1 U11206 ( .A(n12361), .ZN(n10983) );
  INV_X2 U11207 ( .A(n16651), .ZN(n16689) );
  NOR2_X1 U11208 ( .A1(n14899), .A2(n14900), .ZN(n14898) );
  CLKBUF_X2 U11209 ( .A(n12390), .Z(n13678) );
  INV_X1 U11210 ( .A(n12354), .ZN(n10985) );
  CLKBUF_X1 U11211 ( .A(n11420), .Z(n15280) );
  INV_X1 U11212 ( .A(n11973), .ZN(n11007) );
  BUF_X1 U11213 ( .A(n11404), .Z(n15340) );
  NAND2_X2 U11214 ( .A1(n11785), .A2(n15313), .ZN(n11921) );
  INV_X2 U11215 ( .A(n20801), .ZN(n20971) );
  INV_X1 U11216 ( .A(n15869), .ZN(n13121) );
  NOR2_X2 U11217 ( .A1(n12913), .A2(n15411), .ZN(n12935) );
  NOR2_X1 U11218 ( .A1(n11398), .A2(n15313), .ZN(n11399) );
  NAND2_X4 U11219 ( .A1(n14636), .A2(n11383), .ZN(n15313) );
  BUF_X1 U11220 ( .A(n11381), .Z(n19592) );
  INV_X4 U11221 ( .A(n13961), .ZN(n18031) );
  INV_X4 U11222 ( .A(n15306), .ZN(n14287) );
  CLKBUF_X2 U11223 ( .A(n11369), .Z(n14482) );
  BUF_X2 U11224 ( .A(n12507), .Z(n13418) );
  CLKBUF_X2 U11225 ( .A(n12686), .Z(n13564) );
  BUF_X2 U11226 ( .A(n12687), .Z(n13585) );
  BUF_X2 U11227 ( .A(n13908), .Z(n18026) );
  BUF_X2 U11228 ( .A(n12518), .Z(n13584) );
  CLKBUF_X2 U11229 ( .A(n20031), .Z(n21515) );
  INV_X2 U11230 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n21461) );
  INV_X2 U11231 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12883) );
  AND2_X1 U11232 ( .A1(n13622), .A2(n13621), .ZN(n16325) );
  NAND2_X1 U11233 ( .A1(n11038), .A2(n13688), .ZN(n16258) );
  AOI21_X1 U11234 ( .B1(n15979), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15978), .ZN(n15982) );
  XNOR2_X1 U11235 ( .A(n16559), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n20160) );
  XNOR2_X1 U11236 ( .A(n15977), .B(n13720), .ZN(n15979) );
  AOI21_X1 U11237 ( .B1(n16779), .B2(n17668), .A(n16778), .ZN(n16780) );
  AND2_X1 U11238 ( .A1(n10988), .A2(n10989), .ZN(n12865) );
  NAND2_X1 U11239 ( .A1(n11198), .A2(n11195), .ZN(n11194) );
  NOR2_X1 U11240 ( .A1(n11033), .A2(n16381), .ZN(n16510) );
  NAND2_X1 U11241 ( .A1(n16895), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16889) );
  CLKBUF_X1 U11242 ( .A(n15612), .Z(n16557) );
  NOR2_X1 U11243 ( .A1(n16930), .A2(n17069), .ZN(n16895) );
  XNOR2_X1 U11244 ( .A(n13675), .B(n13676), .ZN(n15993) );
  OR2_X1 U11245 ( .A1(n16903), .A2(n16900), .ZN(n16860) );
  NAND2_X1 U11246 ( .A1(n11745), .A2(n14506), .ZN(n13749) );
  NAND2_X1 U11247 ( .A1(n13663), .A2(n12433), .ZN(n16074) );
  NAND2_X1 U11248 ( .A1(n11181), .A2(n11176), .ZN(n16647) );
  OR2_X1 U11249 ( .A1(n16703), .A2(n16702), .ZN(n18856) );
  AND2_X1 U11250 ( .A1(n15980), .A2(n13723), .ZN(n10977) );
  NAND2_X1 U11251 ( .A1(n16663), .A2(n11024), .ZN(n14396) );
  AOI21_X1 U11252 ( .B1(n13632), .B2(n13631), .A(n13630), .ZN(n13633) );
  OR2_X1 U11253 ( .A1(n16395), .A2(n16398), .ZN(n16390) );
  NAND2_X1 U11254 ( .A1(n16665), .A2(n16664), .ZN(n16663) );
  NAND2_X1 U11255 ( .A1(n18833), .A2(n18832), .ZN(n16602) );
  OR2_X1 U11256 ( .A1(n14536), .A2(n13629), .ZN(n16415) );
  AND2_X1 U11257 ( .A1(n12850), .A2(n12852), .ZN(n16392) );
  OR2_X2 U11258 ( .A1(n16116), .A2(n16100), .ZN(n16102) );
  INV_X2 U11259 ( .A(n12850), .ZN(n16382) );
  NAND2_X1 U11260 ( .A1(n16129), .A2(n16117), .ZN(n16116) );
  XNOR2_X1 U11261 ( .A(n12840), .B(n12827), .ZN(n13186) );
  NOR2_X1 U11262 ( .A1(n15797), .A2(n15880), .ZN(n15878) );
  AND2_X1 U11263 ( .A1(n12290), .A2(n12295), .ZN(n10978) );
  XNOR2_X1 U11264 ( .A(n13711), .B(n13710), .ZN(n18828) );
  NAND2_X1 U11265 ( .A1(n12816), .A2(n12815), .ZN(n12840) );
  OR2_X1 U11266 ( .A1(n15578), .A2(n15634), .ZN(n15706) );
  NAND2_X1 U11267 ( .A1(n12789), .A2(n12790), .ZN(n12818) );
  NAND2_X1 U11268 ( .A1(n11190), .A2(n11189), .ZN(n15946) );
  OR2_X1 U11269 ( .A1(n20667), .A2(n20668), .ZN(n11122) );
  NAND2_X1 U11270 ( .A1(n12766), .A2(n12765), .ZN(n12792) );
  NAND2_X1 U11271 ( .A1(n18311), .A2(n18315), .ZN(n18310) );
  NAND2_X1 U11272 ( .A1(n20967), .A2(P3_EAX_REG_15__SCAN_IN), .ZN(n20965) );
  NOR2_X1 U11273 ( .A1(n18321), .A2(n13871), .ZN(n21208) );
  NOR3_X2 U11274 ( .A1(n20859), .A2(n20858), .A3(n20857), .ZN(n20967) );
  NAND2_X1 U11275 ( .A1(n11157), .A2(n11156), .ZN(n14797) );
  NAND2_X1 U11276 ( .A1(n20970), .A2(P3_EAX_REG_7__SCAN_IN), .ZN(n20859) );
  NAND2_X1 U11277 ( .A1(n13133), .A2(n13132), .ZN(n14909) );
  AOI21_X1 U11278 ( .B1(n13874), .B2(n13873), .A(n18258), .ZN(n13877) );
  NOR2_X1 U11279 ( .A1(n18327), .A2(n21166), .ZN(n21170) );
  AND2_X1 U11280 ( .A1(n11124), .A2(n11123), .ZN(n20654) );
  NAND2_X1 U11281 ( .A1(n11125), .A2(n20592), .ZN(n11124) );
  CLKBUF_X1 U11282 ( .A(n15870), .Z(n16296) );
  NAND2_X1 U11283 ( .A1(n20828), .A2(P3_EAX_REG_1__SCAN_IN), .ZN(n20981) );
  AOI22_X1 U11284 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19439), .B1(
        n11508), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11515) );
  NAND2_X1 U11285 ( .A1(n13648), .A2(n13647), .ZN(n21622) );
  OAI21_X1 U11286 ( .B1(n22063), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n12700), 
        .ZN(n12701) );
  INV_X1 U11287 ( .A(n20985), .ZN(n20828) );
  AOI211_X1 U11288 ( .C1(n17356), .C2(n15174), .A(n14867), .B(n14866), .ZN(
        n21796) );
  OR2_X1 U11289 ( .A1(n20628), .A2(n20629), .ZN(n11125) );
  CLKBUF_X1 U11290 ( .A(n11638), .Z(n19417) );
  XNOR2_X1 U11291 ( .A(n14890), .B(n15081), .ZN(n22015) );
  INV_X1 U11292 ( .A(n19447), .ZN(n19450) );
  NAND2_X1 U11293 ( .A1(n16514), .A2(n13029), .ZN(n16517) );
  OR2_X1 U11294 ( .A1(n11628), .A2(n14329), .ZN(n11518) );
  AOI21_X1 U11295 ( .B1(n17318), .B2(n20284), .A(n17300), .ZN(n20797) );
  OR2_X2 U11296 ( .A1(n11496), .A2(n11497), .ZN(n11624) );
  OR2_X1 U11297 ( .A1(n12681), .A2(n12680), .ZN(n12682) );
  NAND2_X1 U11298 ( .A1(n12681), .A2(n12680), .ZN(n14890) );
  NOR2_X2 U11299 ( .A1(n12368), .A2(n14525), .ZN(n12370) );
  NAND2_X1 U11300 ( .A1(n16136), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15163) );
  OR2_X2 U11301 ( .A1(n12366), .A2(n12365), .ZN(n12368) );
  CLKBUF_X3 U11302 ( .A(n20615), .Z(n20765) );
  NAND2_X1 U11303 ( .A1(n14113), .A2(n14125), .ZN(n14916) );
  INV_X1 U11304 ( .A(n21003), .ZN(n13998) );
  OR2_X1 U11305 ( .A1(n12363), .A2(n16811), .ZN(n12366) );
  NOR2_X2 U11306 ( .A1(n20132), .A2(n20131), .ZN(n20134) );
  NOR2_X1 U11307 ( .A1(n15648), .A2(n19376), .ZN(n19583) );
  NAND2_X1 U11308 ( .A1(n12990), .A2(n12989), .ZN(n20132) );
  NAND2_X1 U11309 ( .A1(n17302), .A2(n20284), .ZN(n21440) );
  AND2_X1 U11310 ( .A1(n11454), .A2(n11444), .ZN(n18600) );
  NAND2_X1 U11311 ( .A1(n12337), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12361) );
  NOR2_X2 U11312 ( .A1(n19751), .A2(n19837), .ZN(n19752) );
  INV_X2 U11313 ( .A(n20285), .ZN(n20335) );
  NOR2_X2 U11314 ( .A1(n19378), .A2(n19837), .ZN(n19379) );
  NOR2_X2 U11315 ( .A1(n19631), .A2(n19837), .ZN(n19632) );
  NOR2_X2 U11316 ( .A1(n12360), .A2(n12331), .ZN(n12337) );
  NOR2_X2 U11317 ( .A1(n19672), .A2(n19837), .ZN(n19673) );
  INV_X1 U11318 ( .A(n11454), .ZN(n11470) );
  NOR2_X2 U11319 ( .A1(n19712), .A2(n19837), .ZN(n19713) );
  OAI21_X1 U11320 ( .B1(n13989), .B2(n21469), .A(n21476), .ZN(n17317) );
  INV_X2 U11321 ( .A(n18070), .ZN(n18043) );
  NAND2_X1 U11322 ( .A1(n12338), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12360) );
  NAND2_X1 U11323 ( .A1(n11120), .A2(n11434), .ZN(n11453) );
  NAND2_X1 U11324 ( .A1(n14722), .A2(n14721), .ZN(n14720) );
  NAND2_X1 U11325 ( .A1(n12607), .A2(n11106), .ZN(n12642) );
  NAND2_X1 U11326 ( .A1(n11460), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11204) );
  XNOR2_X1 U11327 ( .A(n14734), .B(n11986), .ZN(n14722) );
  NAND2_X1 U11328 ( .A1(n18197), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n18227) );
  AND2_X1 U11329 ( .A1(n14062), .A2(n13985), .ZN(n21469) );
  NAND2_X1 U11330 ( .A1(n14736), .A2(n14735), .ZN(n14734) );
  NOR2_X2 U11331 ( .A1(n12355), .A2(n12330), .ZN(n12358) );
  AND2_X1 U11332 ( .A1(n11201), .A2(n11056), .ZN(n11202) );
  NAND2_X1 U11333 ( .A1(n11390), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11427) );
  NOR2_X1 U11334 ( .A1(n12211), .A2(n12178), .ZN(n12221) );
  NAND2_X1 U11335 ( .A1(n10986), .A2(n10985), .ZN(n12355) );
  AND2_X1 U11336 ( .A1(n12982), .A2(n12981), .ZN(n14900) );
  NAND2_X1 U11337 ( .A1(n12976), .A2(n12975), .ZN(n12978) );
  NAND2_X1 U11338 ( .A1(n11152), .A2(n11151), .ZN(n14736) );
  AND4_X1 U11339 ( .A1(n13098), .A2(n12606), .A3(n12605), .A4(n12604), .ZN(
        n12607) );
  AOI21_X1 U11340 ( .B1(n14695), .B2(n12557), .A(n12968), .ZN(n12572) );
  CLKBUF_X1 U11341 ( .A(n12595), .Z(n12956) );
  BUF_X2 U11342 ( .A(n11464), .Z(n11833) );
  INV_X1 U11343 ( .A(n11991), .ZN(n11986) );
  NAND2_X1 U11344 ( .A1(n14886), .A2(n13074), .ZN(n13071) );
  NAND2_X1 U11345 ( .A1(n11981), .A2(n11031), .ZN(n14735) );
  AND2_X1 U11346 ( .A1(n11406), .A2(n11405), .ZN(n11944) );
  AND2_X1 U11347 ( .A1(n11985), .A2(n11984), .ZN(n11991) );
  AND2_X1 U11348 ( .A1(n20584), .A2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18093) );
  AND2_X1 U11349 ( .A1(n11378), .A2(n11923), .ZN(n11926) );
  INV_X2 U11350 ( .A(n12973), .ZN(n14886) );
  NOR2_X1 U11351 ( .A1(n19055), .A2(n20856), .ZN(n20804) );
  OAI21_X1 U11352 ( .B1(n12914), .B2(n12913), .A(n12915), .ZN(n12919) );
  INV_X1 U11353 ( .A(n20855), .ZN(n19055) );
  AND2_X1 U11354 ( .A1(n11922), .A2(n11397), .ZN(n11412) );
  INV_X1 U11355 ( .A(n15156), .ZN(n14806) );
  BUF_X4 U11356 ( .A(n12973), .Z(n11020) );
  NAND2_X1 U11357 ( .A1(n18100), .A2(n20562), .ZN(n18303) );
  NAND2_X1 U11358 ( .A1(n11403), .A2(n11348), .ZN(n13741) );
  NAND2_X1 U11359 ( .A1(n13623), .A2(n14811), .ZN(n15869) );
  NAND3_X1 U11360 ( .A1(n13970), .A2(n13969), .A3(n13968), .ZN(n20801) );
  INV_X1 U11361 ( .A(n12599), .ZN(n21510) );
  INV_X1 U11362 ( .A(n15215), .ZN(n15228) );
  INV_X1 U11363 ( .A(n14057), .ZN(n20856) );
  INV_X2 U11364 ( .A(n11982), .ZN(n13660) );
  AND3_X1 U11365 ( .A1(n12952), .A2(n12513), .A3(n14700), .ZN(n12947) );
  NAND2_X1 U11366 ( .A1(n15411), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12684) );
  INV_X1 U11367 ( .A(n11800), .ZN(n11348) );
  AND2_X1 U11368 ( .A1(n11384), .A2(n11408), .ZN(n11385) );
  NAND2_X1 U11369 ( .A1(n14099), .A2(n11916), .ZN(n11800) );
  INV_X1 U11370 ( .A(n12601), .ZN(n12967) );
  AND2_X1 U11371 ( .A1(n11193), .A2(n11798), .ZN(n11192) );
  NAND2_X1 U11372 ( .A1(n11577), .A2(n11576), .ZN(n12170) );
  AND2_X1 U11373 ( .A1(n12342), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12340) );
  NAND2_X1 U11374 ( .A1(n11975), .A2(n11392), .ZN(n11408) );
  NAND2_X1 U11375 ( .A1(n11391), .A2(n11381), .ZN(n11801) );
  BUF_X2 U11376 ( .A(n12611), .Z(n15411) );
  NOR2_X1 U11377 ( .A1(n13980), .A2(n13979), .ZN(n19133) );
  AND2_X1 U11378 ( .A1(n14099), .A2(n19674), .ZN(n11191) );
  NOR2_X2 U11379 ( .A1(n13929), .A2(n13928), .ZN(n19174) );
  BUF_X1 U11380 ( .A(n11379), .Z(n11381) );
  INV_X1 U11381 ( .A(n11916), .ZN(n11391) );
  NOR2_X2 U11382 ( .A1(n13939), .A2(n13938), .ZN(n17389) );
  NAND2_X1 U11383 ( .A1(n11379), .A2(n11916), .ZN(n11975) );
  INV_X1 U11384 ( .A(n12971), .ZN(n15096) );
  INV_X2 U11385 ( .A(n14860), .ZN(n12559) );
  AND2_X2 U11386 ( .A1(n11377), .A2(n19753), .ZN(n11923) );
  INV_X1 U11387 ( .A(n14715), .ZN(n19380) );
  NAND2_X1 U11388 ( .A1(n12512), .A2(n11256), .ZN(n12561) );
  AND2_X1 U11389 ( .A1(n12545), .A2(n12544), .ZN(n12556) );
  INV_X2 U11390 ( .A(U212), .ZN(n10964) );
  NAND2_X2 U11391 ( .A1(U214), .A2(n20207), .ZN(n20271) );
  AND4_X1 U11392 ( .A1(n12476), .A2(n12477), .A3(n12475), .A4(n12474), .ZN(
        n12483) );
  OR2_X2 U11393 ( .A1(n12493), .A2(n12492), .ZN(n14811) );
  AND2_X2 U11394 ( .A1(n11299), .A2(n11298), .ZN(n19674) );
  INV_X2 U11395 ( .A(n14230), .ZN(n14278) );
  NAND2_X1 U11396 ( .A1(n12343), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12349) );
  OAI21_X1 U11397 ( .B1(n11292), .B2(n11291), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11299) );
  NOR2_X2 U11398 ( .A1(n18399), .A2(n18397), .ZN(n20414) );
  INV_X2 U11399 ( .A(n19054), .ZN(n19215) );
  AND4_X1 U11400 ( .A1(n12526), .A2(n12525), .A3(n12524), .A4(n12523), .ZN(
        n12533) );
  AND4_X1 U11401 ( .A1(n12517), .A2(n12516), .A3(n12515), .A4(n12514), .ZN(
        n12535) );
  OR2_X2 U11402 ( .A1(n21835), .A2(n22401), .ZN(n17343) );
  INV_X2 U11403 ( .A(n20068), .ZN(n10965) );
  INV_X2 U11404 ( .A(n17850), .ZN(n17909) );
  AND2_X2 U11405 ( .A1(n14482), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14151) );
  NAND2_X1 U11406 ( .A1(n12348), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12347) );
  AND2_X2 U11407 ( .A1(n14483), .A2(n11374), .ZN(n14270) );
  AND4_X1 U11408 ( .A1(n12553), .A2(n12552), .A3(n12551), .A4(n12550), .ZN(
        n12554) );
  INV_X1 U11409 ( .A(n11009), .ZN(n11010) );
  AND4_X1 U11410 ( .A1(n12522), .A2(n12521), .A3(n12520), .A4(n12519), .ZN(
        n12534) );
  INV_X2 U11411 ( .A(n11013), .ZN(n10966) );
  NAND2_X1 U11412 ( .A1(n11093), .A2(n11092), .ZN(n11291) );
  INV_X2 U11413 ( .A(n11012), .ZN(n10967) );
  AND3_X1 U11414 ( .A1(n11325), .A2(n11324), .A3(n11323), .ZN(n11329) );
  AND2_X1 U11415 ( .A1(n11327), .A2(n11326), .ZN(n11328) );
  AND4_X1 U11417 ( .A1(n12501), .A2(n12500), .A3(n12499), .A4(n12498), .ZN(
        n12502) );
  AND4_X1 U11418 ( .A1(n12539), .A2(n12538), .A3(n12537), .A4(n12536), .ZN(
        n12545) );
  AND3_X1 U11419 ( .A1(n12480), .A2(n12479), .A3(n12478), .ZN(n12481) );
  NAND2_X1 U11420 ( .A1(n18413), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18399) );
  AND4_X1 U11421 ( .A1(n12531), .A2(n12530), .A3(n12529), .A4(n12528), .ZN(
        n12532) );
  INV_X1 U11422 ( .A(n12465), .ZN(n13286) );
  NOR2_X1 U11423 ( .A1(n20997), .A2(n18464), .ZN(n21489) );
  INV_X1 U11424 ( .A(n12465), .ZN(n13187) );
  NAND2_X2 U11425 ( .A1(n14480), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14285) );
  NOR2_X2 U11426 ( .A1(n12345), .A2(n17622), .ZN(n12348) );
  INV_X1 U11427 ( .A(n18412), .ZN(n18413) );
  CLKBUF_X3 U11428 ( .A(n13778), .Z(n18056) );
  AND2_X1 U11429 ( .A1(n18358), .A2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n20480) );
  INV_X2 U11430 ( .A(n18571), .ZN(n18553) );
  NAND2_X2 U11431 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n21855), .ZN(n17762) );
  CLKBUF_X2 U11432 ( .A(n13837), .Z(n18034) );
  INV_X2 U11433 ( .A(n19257), .ZN(U215) );
  AND2_X2 U11434 ( .A1(n12452), .A2(n15213), .ZN(n12685) );
  AND2_X1 U11435 ( .A1(n12453), .A2(n12455), .ZN(n12518) );
  BUF_X4 U11436 ( .A(n13848), .Z(n10969) );
  NAND2_X1 U11437 ( .A1(n12453), .A2(n11091), .ZN(n12465) );
  INV_X2 U11438 ( .A(n22398), .ZN(n22401) );
  NAND2_X1 U11439 ( .A1(n12346), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12345) );
  NOR2_X2 U11440 ( .A1(n21461), .A2(n21012), .ZN(n13908) );
  NOR2_X1 U11441 ( .A1(n13761), .A2(n13760), .ZN(n13778) );
  CLKBUF_X1 U11442 ( .A(n13813), .Z(n10970) );
  BUF_X8 U11443 ( .A(n13842), .Z(n10971) );
  NOR2_X2 U11444 ( .A1(n12344), .A2(n15681), .ZN(n12346) );
  CLKBUF_X1 U11445 ( .A(n22117), .Z(n22059) );
  AND2_X2 U11446 ( .A1(n15212), .A2(n15213), .ZN(n12808) );
  NOR2_X2 U11447 ( .A1(n12445), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12452) );
  NAND2_X1 U11448 ( .A1(n21461), .A2(n21006), .ZN(n21022) );
  NAND2_X1 U11449 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21001), .ZN(
        n13761) );
  NAND2_X1 U11450 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n21020), .ZN(
        n13759) );
  NAND2_X1 U11451 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n21461), .ZN(
        n13758) );
  INV_X2 U11452 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n21020) );
  AND2_X2 U11453 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11271) );
  NAND2_X1 U11454 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12344) );
  AND2_X2 U11455 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15213) );
  INV_X1 U11456 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11208) );
  INV_X1 U11457 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11418) );
  NAND2_X1 U11459 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21028) );
  INV_X1 U11460 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n15681) );
  AND2_X1 U11461 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15229) );
  INV_X2 U11462 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12447) );
  AND2_X1 U11463 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18373) );
  NOR2_X1 U11464 ( .A1(n16175), .A2(n16162), .ZN(n10972) );
  INV_X1 U11465 ( .A(n13007), .ZN(n10974) );
  NAND2_X1 U11466 ( .A1(n10975), .A2(n15624), .ZN(n15925) );
  NOR2_X1 U11467 ( .A1(n13015), .A2(n10974), .ZN(n10975) );
  NOR2_X2 U11468 ( .A1(n16175), .A2(n16162), .ZN(n16161) );
  NOR2_X2 U11469 ( .A1(n16219), .A2(n16130), .ZN(n16129) );
  AND2_X1 U11470 ( .A1(n20134), .A2(n12999), .ZN(n15624) );
  OR2_X1 U11471 ( .A1(n12966), .A2(n12601), .ZN(n12599) );
  AND2_X1 U11472 ( .A1(n12967), .A2(n12966), .ZN(n15156) );
  CLKBUF_X1 U11473 ( .A(n16988), .Z(n10976) );
  NOR2_X1 U11474 ( .A1(n16006), .A2(n16005), .ZN(n16007) );
  NAND2_X1 U11475 ( .A1(n11121), .A2(n10977), .ZN(n13730) );
  NAND2_X1 U11476 ( .A1(n16917), .A2(n10978), .ZN(n11206) );
  NAND2_X1 U11478 ( .A1(n12836), .A2(n12835), .ZN(n10980) );
  CLKBUF_X1 U11479 ( .A(n14924), .Z(n10981) );
  NAND2_X1 U11480 ( .A1(n12836), .A2(n12835), .ZN(n15583) );
  NAND2_X1 U11481 ( .A1(n12863), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10982) );
  XNOR2_X1 U11483 ( .A(n12750), .B(n12728), .ZN(n14924) );
  AND2_X1 U11484 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10984) );
  AND2_X1 U11485 ( .A1(n10983), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12335) );
  AND2_X1 U11486 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10986) );
  AND2_X1 U11487 ( .A1(n10985), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12356) );
  NAND2_X1 U11488 ( .A1(n12358), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12357) );
  OR3_X1 U11489 ( .A1(n18224), .A2(n18151), .A3(n11140), .ZN(n11139) );
  NAND2_X2 U11490 ( .A1(n18152), .A2(n18090), .ZN(n18084) );
  NOR2_X1 U11491 ( .A1(n18389), .A2(n13869), .ZN(n14008) );
  AND2_X1 U11492 ( .A1(n11211), .A2(n12667), .ZN(n12702) );
  CLKBUF_X1 U11493 ( .A(n15556), .Z(n10987) );
  NAND2_X1 U11494 ( .A1(n16366), .A2(n10991), .ZN(n10988) );
  OR2_X1 U11495 ( .A1(n10990), .A2(n20182), .ZN(n10989) );
  INV_X1 U11496 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10990) );
  AND2_X1 U11497 ( .A1(n12860), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10991) );
  AND2_X1 U11498 ( .A1(n10982), .A2(n16334), .ZN(n10992) );
  NAND2_X1 U11499 ( .A1(n12824), .A2(n12823), .ZN(n15556) );
  INV_X2 U11500 ( .A(n13749), .ZN(n16807) );
  OAI21_X2 U11501 ( .B1(n17247), .B2(n11148), .A(n11146), .ZN(n16988) );
  NAND4_X1 U11502 ( .A1(n11205), .A2(n11204), .A3(n11202), .A4(n11203), .ZN(
        n11446) );
  INV_X1 U11503 ( .A(n10995), .ZN(n10993) );
  XNOR2_X1 U11504 ( .A(n12591), .B(n12590), .ZN(n15125) );
  NAND2_X2 U11505 ( .A1(n11149), .A2(n11711), .ZN(n11710) );
  INV_X1 U11506 ( .A(n11427), .ZN(n10994) );
  INV_X1 U11507 ( .A(n11427), .ZN(n11460) );
  AND2_X2 U11508 ( .A1(n15363), .A2(n11047), .ZN(n15469) );
  NAND2_X1 U11511 ( .A1(n12864), .A2(n16334), .ZN(n16304) );
  NOR2_X2 U11512 ( .A1(n13883), .A2(n21306), .ZN(n18248) );
  INV_X1 U11513 ( .A(n15125), .ZN(n10995) );
  INV_X2 U11514 ( .A(n12558), .ZN(n13623) );
  NAND2_X1 U11515 ( .A1(n12571), .A2(n12570), .ZN(n10996) );
  NAND2_X1 U11516 ( .A1(n12562), .A2(n12558), .ZN(n10997) );
  NAND2_X1 U11517 ( .A1(n12571), .A2(n12570), .ZN(n12962) );
  NOR2_X1 U11518 ( .A1(n15578), .A2(n10998), .ZN(n15799) );
  OR2_X1 U11519 ( .A1(n15634), .A2(n15707), .ZN(n10998) );
  NOR2_X2 U11520 ( .A1(n18266), .A2(n18254), .ZN(n18253) );
  NOR2_X2 U11521 ( .A1(n18296), .A2(n20736), .ZN(n18295) );
  NAND2_X1 U11522 ( .A1(n12865), .A2(n16358), .ZN(n10999) );
  NAND2_X1 U11523 ( .A1(n12865), .A2(n16358), .ZN(n11000) );
  NAND2_X1 U11524 ( .A1(n12865), .A2(n16358), .ZN(n13689) );
  NAND2_X1 U11525 ( .A1(n16566), .A2(n20182), .ZN(n11002) );
  NAND2_X1 U11526 ( .A1(n16558), .A2(n16382), .ZN(n11003) );
  NAND2_X1 U11527 ( .A1(n11002), .A2(n11003), .ZN(n16559) );
  NAND2_X2 U11529 ( .A1(n14074), .A2(n13998), .ZN(n17318) );
  NOR2_X2 U11530 ( .A1(n20937), .A2(n20896), .ZN(n20902) );
  NOR2_X2 U11531 ( .A1(n20928), .A2(n20929), .ZN(n20927) );
  NOR2_X2 U11532 ( .A1(n20965), .A2(n20952), .ZN(n20951) );
  NOR2_X2 U11533 ( .A1(n13759), .A2(n13758), .ZN(n13842) );
  INV_X1 U11534 ( .A(n15444), .ZN(n11004) );
  OAI21_X2 U11535 ( .B1(n16633), .B2(n16632), .A(n16631), .ZN(n16712) );
  NOR2_X4 U11536 ( .A1(n15190), .A2(n14134), .ZN(n15183) );
  AND2_X1 U11537 ( .A1(n15986), .A2(n14502), .ZN(n16652) );
  AND2_X1 U11538 ( .A1(n11360), .A2(n11359), .ZN(n11363) );
  NAND2_X2 U11539 ( .A1(n16988), .A2(n11740), .ZN(n11745) );
  NAND2_X1 U11540 ( .A1(n12667), .A2(n12641), .ZN(n13128) );
  NOR2_X2 U11541 ( .A1(n12281), .A2(n12273), .ZN(n12269) );
  NOR3_X2 U11542 ( .A1(n12262), .A2(n12261), .A3(n11116), .ZN(n12291) );
  AOI211_X1 U11543 ( .C1(n18297), .C2(n20763), .A(n18285), .B(n18284), .ZN(
        n18286) );
  INV_X4 U11544 ( .A(n18236), .ZN(n18380) );
  OAI22_X2 U11545 ( .A1(n21445), .A2(n21437), .B1(n21443), .B2(n21102), .ZN(
        n21446) );
  NAND2_X1 U11546 ( .A1(n15624), .A2(n13007), .ZN(n15794) );
  AND2_X2 U11547 ( .A1(n12611), .A2(n12562), .ZN(n12569) );
  OAI21_X1 U11548 ( .B1(n16145), .B2(n16215), .A(n16214), .ZN(n21778) );
  NOR2_X2 U11549 ( .A1(n18807), .A2(n18808), .ZN(n18806) );
  NAND2_X2 U11550 ( .A1(n11166), .A2(n11165), .ZN(n11383) );
  BUF_X8 U11551 ( .A(n11383), .Z(n11969) );
  AOI21_X2 U11552 ( .B1(n10994), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n11465), .ZN(n11828) );
  CLKBUF_X1 U11553 ( .A(n14300), .Z(n14484) );
  NAND2_X1 U11554 ( .A1(n11113), .A2(n11112), .ZN(n15986) );
  OR2_X2 U11555 ( .A1(n14962), .A2(n11110), .ZN(n15188) );
  NOR2_X2 U11556 ( .A1(n18410), .A2(n18411), .ZN(n18409) );
  XNOR2_X2 U11557 ( .A(n11142), .B(n11141), .ZN(n18410) );
  NOR2_X2 U11558 ( .A1(n18394), .A2(n13866), .ZN(n13867) );
  NOR2_X2 U11559 ( .A1(n18396), .A2(n18395), .ZN(n18394) );
  NOR2_X2 U11560 ( .A1(n11969), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12010) );
  INV_X2 U11561 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12445) );
  NAND2_X1 U11562 ( .A1(n10995), .A2(n12609), .ZN(n15082) );
  NOR2_X2 U11563 ( .A1(n14971), .A2(n15073), .ZN(n15074) );
  NAND2_X1 U11564 ( .A1(n13079), .A2(n13078), .ZN(n13081) );
  CLKBUF_X1 U11565 ( .A(n20145), .Z(n11005) );
  CLKBUF_X1 U11566 ( .A(n15490), .Z(n11006) );
  NAND2_X1 U11567 ( .A1(n12594), .A2(n12593), .ZN(n12643) );
  NAND2_X2 U11568 ( .A1(n12590), .A2(n12586), .ZN(n12673) );
  NOR2_X4 U11569 ( .A1(n16808), .A2(n13712), .ZN(n14498) );
  NAND2_X2 U11570 ( .A1(n16807), .A2(n13750), .ZN(n16808) );
  NAND2_X4 U11571 ( .A1(n11034), .A2(n12502), .ZN(n12562) );
  INV_X1 U11572 ( .A(n13813), .ZN(n11009) );
  INV_X1 U11573 ( .A(n10970), .ZN(n11012) );
  INV_X1 U11574 ( .A(n10970), .ZN(n11013) );
  NOR2_X1 U11575 ( .A1(n13759), .A2(n13760), .ZN(n13813) );
  NAND2_X2 U11576 ( .A1(n12573), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12590) );
  NOR2_X2 U11577 ( .A1(n16693), .A2(n16692), .ZN(n16616) );
  BUF_X8 U11579 ( .A(n11983), .Z(n11015) );
  NAND2_X1 U11580 ( .A1(n11416), .A2(n11417), .ZN(n11466) );
  OAI211_X2 U11581 ( .C1(n11944), .C2(n11411), .A(P2_STATE2_REG_0__SCAN_IN), 
        .B(n11413), .ZN(n11417) );
  NAND2_X2 U11582 ( .A1(n11103), .A2(n12859), .ZN(n16366) );
  INV_X2 U11583 ( .A(n12465), .ZN(n11016) );
  NOR3_X4 U11584 ( .A1(n20981), .A2(n20799), .A3(n20798), .ZN(n20970) );
  AND2_X1 U11585 ( .A1(n12453), .A2(n12455), .ZN(n11017) );
  NOR2_X2 U11586 ( .A1(n15789), .A2(n11217), .ZN(n15861) );
  NAND2_X2 U11587 ( .A1(n13235), .A2(n13234), .ZN(n15789) );
  NOR3_X4 U11588 ( .A1(n16671), .A2(n16670), .A3(n11114), .ZN(n16655) );
  NAND2_X2 U11589 ( .A1(n15612), .A2(n12849), .ZN(n15887) );
  NAND2_X1 U11590 ( .A1(n15082), .A2(n12672), .ZN(n15382) );
  NOR2_X2 U11591 ( .A1(n16157), .A2(n16160), .ZN(n16143) );
  AND2_X2 U11592 ( .A1(n16143), .A2(n13461), .ZN(n16145) );
  XNOR2_X2 U11593 ( .A(n12726), .B(n12725), .ZN(n14897) );
  NAND2_X2 U11594 ( .A1(n12724), .A2(n12723), .ZN(n12726) );
  AND2_X4 U11595 ( .A1(n12454), .A2(n11091), .ZN(n13419) );
  XNOR2_X2 U11596 ( .A(n14772), .B(n12721), .ZN(n11111) );
  NAND2_X1 U11597 ( .A1(n12720), .A2(n12719), .ZN(n12721) );
  OAI21_X2 U11598 ( .B1(n16113), .B2(n16115), .A(n16114), .ZN(n16337) );
  NOR2_X4 U11599 ( .A1(n16127), .A2(n16128), .ZN(n16113) );
  INV_X1 U11600 ( .A(n11022), .ZN(n11023) );
  XNOR2_X2 U11601 ( .A(n11105), .B(n12643), .ZN(n13136) );
  NOR2_X1 U11602 ( .A1(n11215), .A2(n16104), .ZN(n11214) );
  INV_X1 U11603 ( .A(n13687), .ZN(n11215) );
  AND2_X1 U11604 ( .A1(n13987), .A2(n14977), .ZN(n13988) );
  AND2_X1 U11605 ( .A1(n20793), .A2(n20801), .ZN(n13987) );
  NAND2_X1 U11606 ( .A1(n11440), .A2(n11441), .ZN(n11454) );
  OR2_X1 U11607 ( .A1(n21471), .A2(n21876), .ZN(n17300) );
  NAND2_X1 U11608 ( .A1(n12888), .A2(n12887), .ZN(n12899) );
  NAND2_X1 U11609 ( .A1(n12966), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12683) );
  NAND2_X1 U11610 ( .A1(n14099), .A2(n19674), .ZN(n11101) );
  INV_X1 U11611 ( .A(n19674), .ZN(n11100) );
  AND2_X1 U11612 ( .A1(n11969), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14106) );
  INV_X2 U11613 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15266) );
  NAND2_X2 U11614 ( .A1(n12684), .A2(n12683), .ZN(n12943) );
  NAND2_X1 U11615 ( .A1(n11225), .A2(n11223), .ZN(n15566) );
  NAND2_X1 U11616 ( .A1(n11227), .A2(n15568), .ZN(n11226) );
  INV_X1 U11617 ( .A(n11057), .ZN(n11227) );
  AND2_X2 U11618 ( .A1(n12559), .A2(n15096), .ZN(n15215) );
  INV_X1 U11619 ( .A(n12561), .ZN(n12611) );
  AND2_X1 U11620 ( .A1(n11777), .A2(n11776), .ZN(n15316) );
  NAND2_X1 U11621 ( .A1(n12191), .A2(n11026), .ZN(n12194) );
  INV_X1 U11622 ( .A(n14417), .ZN(n14346) );
  OR2_X1 U11623 ( .A1(n14127), .A2(n14918), .ZN(n14942) );
  CLKBUF_X1 U11624 ( .A(n12021), .Z(n12418) );
  NAND2_X1 U11625 ( .A1(n14720), .A2(n11992), .ZN(n11999) );
  INV_X1 U11626 ( .A(n18157), .ZN(n11133) );
  NOR2_X1 U11627 ( .A1(n21020), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n14002) );
  AOI21_X1 U11628 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n17316), .A(
        n13901), .ZN(n14003) );
  AND2_X1 U11629 ( .A1(n22106), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13604) );
  NAND2_X1 U11630 ( .A1(n11216), .A2(n11214), .ZN(n11213) );
  INV_X1 U11631 ( .A(n13620), .ZN(n11216) );
  NAND2_X1 U11632 ( .A1(n15469), .A2(n15499), .ZN(n15497) );
  AND2_X1 U11633 ( .A1(n14770), .A2(n15755), .ZN(n11155) );
  NAND2_X1 U11634 ( .A1(n14120), .A2(n14119), .ZN(n14733) );
  NAND2_X1 U11635 ( .A1(n18600), .A2(n14116), .ZN(n14120) );
  AOI22_X1 U11636 ( .A1(n17909), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17920), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13893) );
  AOI22_X1 U11637 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n18054), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13894) );
  AOI211_X1 U11638 ( .C1(n18047), .C2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A(
        n13891), .B(n13890), .ZN(n13892) );
  NAND2_X1 U11639 ( .A1(n14150), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n11098) );
  OR3_X2 U11640 ( .A1(n11487), .A2(n16033), .A3(n11497), .ZN(n11629) );
  AOI21_X1 U11641 ( .B1(n12899), .B2(n12890), .A(n12889), .ZN(n12897) );
  OR2_X1 U11642 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n22105), .ZN(
        n12890) );
  AND2_X1 U11643 ( .A1(n12447), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12453) );
  INV_X1 U11644 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11209) );
  NAND2_X1 U11645 ( .A1(n11716), .A2(n11715), .ZN(n11735) );
  INV_X1 U11646 ( .A(n12231), .ZN(n11716) );
  OAI21_X1 U11647 ( .B1(n14715), .B2(n11977), .A(n19459), .ZN(n11978) );
  NOR2_X1 U11648 ( .A1(n20845), .A2(n14022), .ZN(n14019) );
  NOR2_X1 U11649 ( .A1(n20971), .A2(n19133), .ZN(n14061) );
  NAND2_X1 U11650 ( .A1(n16186), .A2(n11221), .ZN(n16157) );
  AND2_X1 U11651 ( .A1(n11222), .A2(n16172), .ZN(n11221) );
  AND2_X1 U11652 ( .A1(n16229), .A2(n13379), .ZN(n11222) );
  NAND2_X1 U11653 ( .A1(n11220), .A2(n15936), .ZN(n11219) );
  INV_X1 U11654 ( .A(n13299), .ZN(n11220) );
  INV_X1 U11655 ( .A(n15660), .ZN(n13234) );
  INV_X1 U11656 ( .A(n15446), .ZN(n13179) );
  INV_X1 U11657 ( .A(n13597), .ZN(n13600) );
  AND2_X1 U11658 ( .A1(n16343), .A2(n12868), .ZN(n11108) );
  INV_X1 U11659 ( .A(n12853), .ZN(n12854) );
  INV_X1 U11660 ( .A(n15613), .ZN(n12847) );
  INV_X1 U11661 ( .A(n15614), .ZN(n12848) );
  OR2_X1 U11662 ( .A1(n12966), .A2(n21804), .ZN(n12913) );
  INV_X1 U11663 ( .A(n11107), .ZN(n11106) );
  OR2_X1 U11664 ( .A1(n12684), .A2(n12665), .ZN(n12838) );
  AND2_X1 U11665 ( .A1(n15240), .A2(n15239), .ZN(n17365) );
  AND2_X1 U11666 ( .A1(n15210), .A2(n15209), .ZN(n15246) );
  NOR2_X1 U11667 ( .A1(n13707), .A2(n13706), .ZN(n11115) );
  NAND2_X1 U11668 ( .A1(n12192), .A2(n12193), .ZN(n12246) );
  INV_X1 U11669 ( .A(n12194), .ZN(n12192) );
  INV_X1 U11670 ( .A(n12198), .ZN(n12191) );
  NOR2_X1 U11671 ( .A1(n11575), .A2(n11238), .ZN(n11576) );
  NOR2_X1 U11672 ( .A1(n11572), .A2(n11571), .ZN(n11577) );
  NAND2_X1 U11673 ( .A1(n15313), .A2(n11772), .ZN(n12171) );
  OAI211_X1 U11674 ( .C1(n16639), .C2(n16650), .A(n14463), .B(n16647), .ZN(
        n14461) );
  AND2_X1 U11675 ( .A1(n14372), .A2(n11170), .ZN(n11168) );
  NAND2_X1 U11676 ( .A1(n15950), .A2(n11160), .ZN(n11159) );
  INV_X1 U11677 ( .A(n15929), .ZN(n11160) );
  INV_X1 U11678 ( .A(n16798), .ZN(n11121) );
  OR2_X1 U11679 ( .A1(n18804), .A2(n12202), .ZN(n13709) );
  INV_X1 U11680 ( .A(n11745), .ZN(n16930) );
  AND3_X1 U11681 ( .A1(n12071), .A2(n12070), .A3(n12069), .ZN(n14567) );
  AND3_X1 U11682 ( .A1(n11697), .A2(n11248), .A3(n11696), .ZN(n12184) );
  NOR2_X1 U11683 ( .A1(n11704), .A2(n11701), .ZN(n11700) );
  NAND2_X1 U11684 ( .A1(n11704), .A2(n11703), .ZN(n11709) );
  INV_X1 U11685 ( .A(n11702), .ZN(n11703) );
  NAND2_X1 U11686 ( .A1(n11582), .A2(n11581), .ZN(n11612) );
  AND2_X1 U11687 ( .A1(n11804), .A2(n14715), .ZN(n11384) );
  NAND2_X1 U11688 ( .A1(n11035), .A2(n11408), .ZN(n11409) );
  INV_X1 U11689 ( .A(n11476), .ZN(n11492) );
  AOI21_X1 U11690 ( .B1(n11365), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n11374), .ZN(n11277) );
  NAND3_X1 U11691 ( .A1(n11487), .A2(n11477), .A3(n14791), .ZN(n11627) );
  NAND2_X1 U11692 ( .A1(n19571), .A2(n19564), .ZN(n19391) );
  AND2_X1 U11693 ( .A1(n11407), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14116) );
  INV_X1 U11694 ( .A(n13838), .ZN(n13961) );
  NOR2_X1 U11695 ( .A1(n21022), .A2(n20343), .ZN(n13838) );
  NAND2_X1 U11696 ( .A1(n18025), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11090) );
  INV_X1 U11697 ( .A(n13847), .ZN(n11087) );
  NAND2_X1 U11698 ( .A1(n20351), .A2(n13986), .ZN(n20284) );
  OAI21_X1 U11699 ( .B1(n18384), .B2(n18383), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n14037) );
  NAND2_X1 U11700 ( .A1(n18406), .A2(n14031), .ZN(n14033) );
  NOR3_X1 U11701 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21020), .A3(
        n21028), .ZN(n13790) );
  AND2_X1 U11702 ( .A1(n13643), .A2(n17346), .ZN(n13648) );
  OR2_X1 U11703 ( .A1(n12941), .A2(n12940), .ZN(n12946) );
  INV_X1 U11704 ( .A(n15443), .ZN(n11225) );
  XNOR2_X1 U11705 ( .A(n13614), .B(n13613), .ZN(n15161) );
  INV_X1 U11706 ( .A(n11214), .ZN(n11212) );
  NAND2_X1 U11707 ( .A1(n13517), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13553) );
  CLKBUF_X1 U11708 ( .A(n15566), .Z(n15567) );
  NOR2_X1 U11709 ( .A1(n13173), .A2(n21643), .ZN(n13181) );
  AND2_X1 U11710 ( .A1(n15175), .A2(n13120), .ZN(n17371) );
  NAND2_X1 U11711 ( .A1(n16366), .A2(n12860), .ZN(n11104) );
  INV_X1 U11712 ( .A(n15792), .ZN(n13014) );
  NAND2_X1 U11713 ( .A1(n13136), .A2(n21804), .ZN(n12660) );
  INV_X1 U11714 ( .A(n15415), .ZN(n21961) );
  NOR2_X1 U11715 ( .A1(n12956), .A2(n12955), .ZN(n14803) );
  INV_X1 U11716 ( .A(n21813), .ZN(n15174) );
  NAND2_X1 U11717 ( .A1(n16583), .A2(n22013), .ZN(n21988) );
  NAND2_X1 U11718 ( .A1(n21956), .A2(n15080), .ZN(n15124) );
  NAND2_X1 U11719 ( .A1(n15087), .A2(n15123), .ZN(n22054) );
  NAND2_X1 U11720 ( .A1(n15087), .A2(n13134), .ZN(n22085) );
  NAND2_X1 U11721 ( .A1(n13715), .A2(n13716), .ZN(n13722) );
  AND2_X1 U11722 ( .A1(n11246), .A2(n12158), .ZN(n11164) );
  AND4_X1 U11723 ( .A1(n12017), .A2(n12016), .A3(n12015), .A4(n12014), .ZN(
        n15498) );
  AND2_X1 U11724 ( .A1(n14947), .A2(n14946), .ZN(n14131) );
  NAND2_X1 U11725 ( .A1(n14462), .A2(n16632), .ZN(n11187) );
  NAND2_X1 U11726 ( .A1(n14369), .A2(n10959), .ZN(n11174) );
  NOR2_X2 U11727 ( .A1(n14797), .A2(n14567), .ZN(n14937) );
  AND3_X1 U11728 ( .A1(n12057), .A2(n12056), .A3(n12055), .ZN(n14795) );
  NAND2_X1 U11729 ( .A1(n11184), .A2(n14108), .ZN(n14945) );
  AND2_X1 U11730 ( .A1(n14713), .A2(n14712), .ZN(n15264) );
  NAND2_X1 U11731 ( .A1(n10984), .A2(n10983), .ZN(n12363) );
  AND2_X1 U11732 ( .A1(n11745), .A2(n17130), .ZN(n16924) );
  NAND2_X1 U11733 ( .A1(n11934), .A2(n11052), .ZN(n11185) );
  AND2_X1 U11734 ( .A1(n11467), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11422) );
  NAND2_X1 U11735 ( .A1(n16702), .A2(n12430), .ZN(n13663) );
  AND4_X1 U11736 ( .A1(n11726), .A2(n11725), .A3(n11724), .A4(n11723), .ZN(
        n11733) );
  NAND2_X1 U11737 ( .A1(n11199), .A2(n11051), .ZN(n11198) );
  INV_X1 U11738 ( .A(n13705), .ZN(n11199) );
  OR2_X1 U11739 ( .A1(n12322), .A2(n12321), .ZN(n13704) );
  CLKBUF_X1 U11740 ( .A(n15735), .Z(n15736) );
  OR2_X1 U11741 ( .A1(n11737), .A2(n17252), .ZN(n11738) );
  INV_X1 U11742 ( .A(n11147), .ZN(n11146) );
  OAI21_X1 U11743 ( .B1(n17246), .B2(n11148), .A(n16989), .ZN(n11147) );
  INV_X1 U11744 ( .A(n11738), .ZN(n11148) );
  AND2_X1 U11745 ( .A1(n13735), .A2(n11007), .ZN(n12020) );
  AND2_X1 U11746 ( .A1(n11665), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11149) );
  AND2_X1 U11747 ( .A1(n11947), .A2(n15312), .ZN(n17103) );
  AND2_X1 U11748 ( .A1(n11947), .A2(n11935), .ZN(n17104) );
  OR2_X1 U11749 ( .A1(n17103), .A2(n17104), .ZN(n17262) );
  INV_X1 U11750 ( .A(n15471), .ZN(n11161) );
  AND2_X1 U11751 ( .A1(n14785), .A2(n14122), .ZN(n14789) );
  NAND2_X1 U11752 ( .A1(n14788), .A2(n14789), .ZN(n14941) );
  NAND2_X1 U11753 ( .A1(n11364), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11165) );
  NAND2_X1 U11754 ( .A1(n11375), .A2(n11374), .ZN(n11166) );
  AND2_X1 U11755 ( .A1(n11481), .A2(n11476), .ZN(n11474) );
  NAND2_X1 U11756 ( .A1(n19521), .A2(n19502), .ZN(n19402) );
  AND2_X1 U11757 ( .A1(n17328), .A2(n17327), .ZN(n19837) );
  NAND2_X1 U11758 ( .A1(n18906), .A2(n11407), .ZN(n17328) );
  INV_X1 U11759 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19459) );
  NOR2_X1 U11760 ( .A1(n20666), .A2(n20765), .ZN(n20667) );
  INV_X1 U11761 ( .A(n20639), .ZN(n11123) );
  NOR2_X1 U11762 ( .A1(n21500), .A2(n21471), .ZN(n18073) );
  AND2_X1 U11763 ( .A1(n21041), .A2(n21180), .ZN(n18317) );
  NOR2_X1 U11764 ( .A1(n18137), .A2(n11129), .ZN(n11128) );
  INV_X1 U11765 ( .A(n18126), .ZN(n11130) );
  NAND2_X1 U11766 ( .A1(n21296), .A2(n11137), .ZN(n11136) );
  NOR2_X1 U11767 ( .A1(n21102), .A2(n21297), .ZN(n11137) );
  NAND2_X1 U11768 ( .A1(n13833), .A2(n14085), .ZN(n21308) );
  OAI211_X1 U11769 ( .C1(n13907), .C2(n13906), .A(n14003), .B(n14005), .ZN(
        n21445) );
  OAI211_X1 U11770 ( .C1(n17389), .C2(n13997), .A(n13996), .B(n13995), .ZN(
        n21007) );
  INV_X1 U11771 ( .A(n21500), .ZN(n21475) );
  NAND2_X1 U11772 ( .A1(n14532), .A2(n14530), .ZN(n13607) );
  AND2_X1 U11773 ( .A1(n13608), .A2(n22059), .ZN(n20186) );
  NAND2_X1 U11774 ( .A1(n14536), .A2(n14537), .ZN(n13078) );
  NAND2_X1 U11775 ( .A1(n13100), .A2(n13083), .ZN(n21560) );
  AND2_X1 U11777 ( .A1(n16924), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17124) );
  INV_X1 U11778 ( .A(n17647), .ZN(n17631) );
  OR2_X1 U11779 ( .A1(n18917), .A2(n11969), .ZN(n17648) );
  AOI21_X1 U11780 ( .B1(n16779), .B2(n18879), .A(n11250), .ZN(n16047) );
  XNOR2_X1 U11781 ( .A(n13740), .B(n13739), .ZN(n16008) );
  AND2_X1 U11782 ( .A1(n17124), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n17107) );
  INV_X1 U11783 ( .A(n18876), .ZN(n17229) );
  OR2_X1 U11784 ( .A1(n12325), .A2(n11915), .ZN(n18885) );
  INV_X1 U11785 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n20337) );
  INV_X1 U11786 ( .A(n20762), .ZN(n20776) );
  NOR2_X1 U11787 ( .A1(n20707), .A2(n20706), .ZN(n20752) );
  NOR2_X1 U11788 ( .A1(n20971), .A2(n20985), .ZN(n20959) );
  AND2_X1 U11789 ( .A1(n12611), .A2(n14811), .ZN(n12576) );
  INV_X1 U11790 ( .A(n11612), .ZN(n11200) );
  NAND2_X1 U11791 ( .A1(n11341), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11327) );
  NAND2_X1 U11792 ( .A1(n11366), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11326) );
  NAND2_X1 U11793 ( .A1(n11748), .A2(n11747), .ZN(n11757) );
  INV_X1 U11794 ( .A(n11764), .ZN(n11758) );
  OR2_X1 U11795 ( .A1(n13904), .A2(n13905), .ZN(n13896) );
  AOI21_X1 U11796 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n21450), .A(
        n13895), .ZN(n13905) );
  AND2_X1 U11797 ( .A1(n14001), .A2(n14002), .ZN(n13895) );
  NAND2_X1 U11798 ( .A1(n12935), .A2(n12904), .ZN(n12939) );
  INV_X1 U11799 ( .A(n12817), .ZN(n12815) );
  OR2_X1 U11800 ( .A1(n12786), .A2(n12785), .ZN(n12797) );
  OR2_X1 U11801 ( .A1(n12764), .A2(n12763), .ZN(n12794) );
  OAI21_X1 U11802 ( .B1(n12608), .B2(n15401), .A(n13095), .ZN(n11107) );
  INV_X1 U11803 ( .A(n12716), .ZN(n12636) );
  OR2_X1 U11804 ( .A1(n12699), .A2(n12698), .ZN(n12703) );
  NAND2_X1 U11805 ( .A1(n12582), .A2(n16585), .ZN(n12608) );
  AND2_X1 U11806 ( .A1(n12561), .A2(n14811), .ZN(n12565) );
  AND2_X1 U11807 ( .A1(n12269), .A2(n12270), .ZN(n12268) );
  AND3_X1 U11808 ( .A1(n11658), .A2(n11240), .A3(n11657), .ZN(n12011) );
  AND2_X1 U11809 ( .A1(n11809), .A2(n11433), .ZN(n11389) );
  AND2_X1 U11810 ( .A1(n11699), .A2(n11698), .ZN(n11715) );
  NAND2_X1 U11811 ( .A1(n11200), .A2(n12006), .ZN(n11663) );
  INV_X1 U11812 ( .A(n11431), .ZN(n11205) );
  NAND2_X1 U11813 ( .A1(n11466), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11203) );
  NAND2_X1 U11814 ( .A1(n11913), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11201) );
  AND2_X1 U11815 ( .A1(n11975), .A2(n11527), .ZN(n11922) );
  AND2_X1 U11816 ( .A1(n11774), .A2(n11773), .ZN(n11789) );
  INV_X1 U11817 ( .A(n11789), .ZN(n11791) );
  NAND2_X1 U11818 ( .A1(n13834), .A2(n14011), .ZN(n13864) );
  NOR2_X1 U11819 ( .A1(n20840), .A2(n13858), .ZN(n13834) );
  NOR2_X1 U11820 ( .A1(n14027), .A2(n14012), .ZN(n14022) );
  INV_X1 U11821 ( .A(n14061), .ZN(n13999) );
  AND2_X1 U11822 ( .A1(n12896), .A2(n12895), .ZN(n12908) );
  AND2_X1 U11823 ( .A1(n12931), .A2(n12937), .ZN(n12934) );
  NAND2_X1 U11824 ( .A1(n12893), .A2(n12892), .ZN(n12942) );
  NOR2_X1 U11825 ( .A1(n12939), .A2(n12942), .ZN(n12940) );
  OR2_X1 U11826 ( .A1(n15835), .A2(n15833), .ZN(n13299) );
  OR2_X1 U11827 ( .A1(n13218), .A2(n13217), .ZN(n13236) );
  NOR2_X1 U11828 ( .A1(n13147), .A2(n15167), .ZN(n13166) );
  AND2_X1 U11829 ( .A1(n12988), .A2(n12987), .ZN(n15145) );
  OR2_X1 U11830 ( .A1(n12656), .A2(n12655), .ZN(n12715) );
  OR2_X1 U11831 ( .A1(n12635), .A2(n12634), .ZN(n12841) );
  INV_X1 U11832 ( .A(n13129), .ZN(n11210) );
  NAND3_X2 U11833 ( .A1(n12556), .A2(n12555), .A3(n12554), .ZN(n12601) );
  AOI21_X1 U11834 ( .B1(n12650), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A(
        n12549), .ZN(n12555) );
  NAND2_X1 U11835 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12531) );
  NAND2_X1 U11836 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12526) );
  AND2_X1 U11837 ( .A1(n12473), .A2(n12472), .ZN(n12477) );
  INV_X1 U11838 ( .A(n13134), .ZN(n15123) );
  NAND2_X1 U11839 ( .A1(n12745), .A2(n12744), .ZN(n21955) );
  NAND2_X1 U11840 ( .A1(n22015), .A2(n21804), .ZN(n12745) );
  INV_X1 U11841 ( .A(n22013), .ZN(n21956) );
  NAND2_X1 U11842 ( .A1(n11376), .A2(n11527), .ZN(n11785) );
  INV_X1 U11843 ( .A(n14636), .ZN(n11376) );
  NOR2_X1 U11844 ( .A1(n12314), .A2(n12313), .ZN(n12404) );
  INV_X1 U11845 ( .A(n12288), .ZN(n11116) );
  NAND2_X1 U11846 ( .A1(n12268), .A2(n12283), .ZN(n12267) );
  NAND2_X1 U11847 ( .A1(n11095), .A2(n11094), .ZN(n12177) );
  NAND2_X1 U11848 ( .A1(n15313), .A2(n11773), .ZN(n11094) );
  NAND2_X1 U11849 ( .A1(n12002), .A2(n11394), .ZN(n11095) );
  NAND2_X1 U11850 ( .A1(n11204), .A2(n11205), .ZN(n11449) );
  NAND2_X1 U11851 ( .A1(n11179), .A2(n11178), .ZN(n11177) );
  INV_X1 U11852 ( .A(n16659), .ZN(n11178) );
  AND2_X1 U11853 ( .A1(n14325), .A2(n14324), .ZN(n14369) );
  INV_X1 U11854 ( .A(n11397), .ZN(n11925) );
  NOR2_X2 U11855 ( .A1(n12357), .A2(n16888), .ZN(n12338) );
  NOR2_X2 U11856 ( .A1(n12347), .A2(n17645), .ZN(n12343) );
  NOR2_X1 U11857 ( .A1(n16816), .A2(n11196), .ZN(n11195) );
  INV_X1 U11858 ( .A(n13704), .ZN(n11196) );
  AND2_X1 U11859 ( .A1(n18790), .A2(n13735), .ZN(n12320) );
  NAND2_X1 U11860 ( .A1(n15134), .A2(n17145), .ZN(n15423) );
  AND2_X1 U11861 ( .A1(n16978), .A2(n12241), .ZN(n12237) );
  NAND2_X1 U11862 ( .A1(n11469), .A2(n11468), .ZN(n11827) );
  NAND2_X1 U11863 ( .A1(n11466), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11120) );
  INV_X1 U11864 ( .A(n12170), .ZN(n11993) );
  NAND2_X1 U11865 ( .A1(n11007), .A2(n11974), .ZN(n11152) );
  AND2_X1 U11866 ( .A1(n11762), .A2(n11761), .ZN(n11795) );
  CLKBUF_X1 U11867 ( .A(n11271), .Z(n15283) );
  OR2_X1 U11868 ( .A1(n19521), .A2(n17692), .ZN(n19491) );
  NAND2_X1 U11869 ( .A1(n14300), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11092) );
  NAND2_X1 U11870 ( .A1(n11369), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11093) );
  NAND2_X1 U11871 ( .A1(n11304), .A2(n11374), .ZN(n11311) );
  NAND2_X1 U11872 ( .A1(n11309), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11310) );
  AND2_X1 U11873 ( .A1(n17676), .A2(n18909), .ZN(n19382) );
  CLKBUF_X1 U11874 ( .A(n15266), .Z(n15291) );
  AOI21_X1 U11875 ( .B1(n11765), .B2(n11781), .A(n11795), .ZN(n15319) );
  OR2_X1 U11876 ( .A1(n11247), .A2(n21329), .ZN(n11140) );
  INV_X1 U11877 ( .A(n21315), .ZN(n11134) );
  NAND2_X1 U11878 ( .A1(n18084), .A2(n13880), .ZN(n18151) );
  OR2_X1 U11879 ( .A1(n18086), .A2(n18121), .ZN(n18090) );
  NAND2_X1 U11880 ( .A1(n14008), .A2(n21308), .ZN(n18105) );
  NOR2_X1 U11881 ( .A1(n20832), .A2(n13864), .ZN(n13833) );
  OR2_X2 U11882 ( .A1(n18424), .A2(n13860), .ZN(n11142) );
  NOR2_X1 U11883 ( .A1(n13990), .A2(n20803), .ZN(n14067) );
  AOI21_X1 U11884 ( .B1(n14068), .B2(n14060), .A(n14059), .ZN(n13994) );
  AND2_X1 U11885 ( .A1(n12947), .A2(n15178), .ZN(n14695) );
  NAND2_X1 U11886 ( .A1(n21656), .A2(P1_REIP_REG_7__SCAN_IN), .ZN(n21666) );
  INV_X1 U11887 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n15167) );
  AND2_X1 U11888 ( .A1(n13054), .A2(n13053), .ZN(n16162) );
  AOI22_X1 U11889 ( .A1(n12527), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        P1_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n13238), .ZN(n12488) );
  INV_X1 U11890 ( .A(n15942), .ZN(n15865) );
  AND2_X1 U11891 ( .A1(n15177), .A2(n17347), .ZN(n20017) );
  AOI21_X1 U11892 ( .B1(n13603), .B2(n13602), .A(n13601), .ZN(n14530) );
  NAND2_X1 U11893 ( .A1(n13555), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13612) );
  AOI21_X1 U11894 ( .B1(n13600), .B2(n16097), .A(n13552), .ZN(n13687) );
  OAI21_X1 U11895 ( .B1(n13597), .B2(n16329), .A(n13536), .ZN(n16104) );
  AND2_X1 U11896 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n13479), .ZN(
        n13480) );
  INV_X1 U11897 ( .A(n13478), .ZN(n13479) );
  AOI21_X1 U11898 ( .B1(n13600), .B2(n21781), .A(n13477), .ZN(n16215) );
  NOR2_X1 U11899 ( .A1(n13434), .A2(n13433), .ZN(n13435) );
  NOR2_X1 U11900 ( .A1(n13409), .A2(n21763), .ZN(n13410) );
  NAND2_X1 U11901 ( .A1(n13410), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13434) );
  CLKBUF_X1 U11902 ( .A(n16157), .Z(n16158) );
  AND2_X1 U11903 ( .A1(n21768), .A2(n13600), .ZN(n13393) );
  AND2_X1 U11904 ( .A1(n13375), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13376) );
  NAND2_X1 U11905 ( .A1(n13376), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13409) );
  NOR2_X1 U11906 ( .A1(n13343), .A2(n16195), .ZN(n13375) );
  CLKBUF_X1 U11907 ( .A(n16186), .Z(n16187) );
  NAND2_X1 U11908 ( .A1(n13330), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13343) );
  NAND2_X1 U11909 ( .A1(n11218), .A2(n15863), .ZN(n11217) );
  INV_X1 U11910 ( .A(n11219), .ZN(n11218) );
  NAND2_X1 U11911 ( .A1(n13300), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13315) );
  NOR2_X1 U11912 ( .A1(n13253), .A2(n15914), .ZN(n13300) );
  NAND2_X1 U11913 ( .A1(n13237), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13253) );
  INV_X1 U11914 ( .A(n13281), .ZN(n13237) );
  NOR2_X1 U11915 ( .A1(n13236), .A2(n13219), .ZN(n13280) );
  NAND2_X1 U11916 ( .A1(n13280), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13281) );
  NAND2_X1 U11917 ( .A1(n13203), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13218) );
  AND2_X1 U11918 ( .A1(n13181), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13203) );
  AOI21_X1 U11919 ( .B1(n13178), .B2(n13312), .A(n13177), .ZN(n15446) );
  CLKBUF_X1 U11920 ( .A(n15443), .Z(n15444) );
  AND2_X1 U11921 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n13166), .ZN(
        n13167) );
  NAND2_X1 U11922 ( .A1(n13167), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13173) );
  AOI21_X1 U11923 ( .B1(n13161), .B2(n13312), .A(n13160), .ZN(n15198) );
  NAND2_X1 U11924 ( .A1(n15114), .A2(n13145), .ZN(n15107) );
  OAI21_X1 U11925 ( .B1(n13126), .B2(n13163), .A(n13125), .ZN(n13127) );
  NAND2_X1 U11926 ( .A1(n16304), .A2(n11108), .ZN(n11109) );
  OAI21_X1 U11927 ( .B1(n13689), .B2(n13690), .A(n16382), .ZN(n16334) );
  AND3_X1 U11928 ( .A1(n21530), .A2(n13106), .A3(n13105), .ZN(n21598) );
  AND2_X1 U11929 ( .A1(n13046), .A2(n13045), .ZN(n16231) );
  AND2_X1 U11930 ( .A1(n15622), .A2(n15623), .ZN(n13007) );
  OAI21_X1 U11931 ( .B1(n15583), .B2(n15584), .A(n12846), .ZN(n15614) );
  OR2_X1 U11932 ( .A1(n12845), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12846) );
  INV_X1 U11933 ( .A(n15145), .ZN(n12989) );
  INV_X1 U11934 ( .A(n15144), .ZN(n12990) );
  NAND2_X1 U11935 ( .A1(n14898), .A2(n14930), .ZN(n15144) );
  INV_X1 U11936 ( .A(n15616), .ZN(n21530) );
  NOR2_X1 U11937 ( .A1(n21531), .A2(n14881), .ZN(n21533) );
  INV_X1 U11938 ( .A(n16453), .ZN(n21544) );
  NOR2_X1 U11939 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n16468), .ZN(
        n14881) );
  NAND2_X1 U11940 ( .A1(n14535), .A2(n13070), .ZN(n14777) );
  INV_X1 U11941 ( .A(n12642), .ZN(n11105) );
  NAND2_X1 U11942 ( .A1(n12672), .A2(n12671), .ZN(n12681) );
  NAND2_X1 U11943 ( .A1(n12679), .A2(n12678), .ZN(n12680) );
  INV_X1 U11944 ( .A(n12583), .ZN(n16585) );
  AND2_X1 U11945 ( .A1(n12569), .A2(n15156), .ZN(n12570) );
  NAND2_X1 U11946 ( .A1(n14865), .A2(n14864), .ZN(n17356) );
  NAND2_X1 U11947 ( .A1(n20186), .A2(n15942), .ZN(n15414) );
  INV_X1 U11948 ( .A(n21992), .ZN(n22113) );
  INV_X1 U11949 ( .A(n15175), .ZN(n14870) );
  AND2_X1 U11950 ( .A1(n12406), .A2(n13721), .ZN(n13731) );
  NOR2_X1 U11951 ( .A1(n13711), .A2(n12405), .ZN(n13715) );
  NAND2_X1 U11952 ( .A1(n11115), .A2(n11058), .ZN(n13711) );
  INV_X1 U11953 ( .A(n11115), .ZN(n13714) );
  NOR2_X1 U11954 ( .A1(n18796), .A2(n18795), .ZN(n18794) );
  NAND2_X1 U11955 ( .A1(n12312), .A2(n12311), .ZN(n12314) );
  NAND2_X1 U11956 ( .A1(n18752), .A2(n18783), .ZN(n18781) );
  NAND2_X1 U11957 ( .A1(n11119), .A2(n11118), .ZN(n12281) );
  INV_X1 U11958 ( .A(n12278), .ZN(n11118) );
  INV_X1 U11959 ( .A(n12279), .ZN(n11119) );
  OR2_X1 U11960 ( .A1(n12257), .A2(n12258), .ZN(n12279) );
  NAND2_X1 U11961 ( .A1(n12191), .A2(n12199), .ZN(n12197) );
  NAND2_X1 U11962 ( .A1(n12220), .A2(n12233), .ZN(n12186) );
  MUX2_X1 U11963 ( .A(n12177), .B(n15684), .S(n19633), .Z(n12205) );
  MUX2_X1 U11964 ( .A(n12174), .B(n12173), .S(n19633), .Z(n12213) );
  NAND2_X1 U11965 ( .A1(n12213), .A2(n12212), .ZN(n12211) );
  NAND2_X1 U11966 ( .A1(n12427), .A2(n11163), .ZN(n11162) );
  NOR2_X1 U11967 ( .A1(n11179), .A2(n14397), .ZN(n11176) );
  OR2_X2 U11968 ( .A1(n16660), .A2(n16659), .ZN(n11181) );
  OAI211_X1 U11969 ( .C1(n11171), .C2(n14372), .A(n11169), .B(n11167), .ZN(
        n16665) );
  NAND2_X1 U11970 ( .A1(n16675), .A2(n11172), .ZN(n11169) );
  NAND2_X1 U11971 ( .A1(n11171), .A2(n11168), .ZN(n11167) );
  OR2_X1 U11972 ( .A1(n11159), .A2(n16762), .ZN(n11158) );
  CLKBUF_X1 U11973 ( .A(n16679), .Z(n16684) );
  INV_X1 U11974 ( .A(n15882), .ZN(n11189) );
  INV_X1 U11975 ( .A(n15638), .ZN(n11190) );
  AND3_X1 U11976 ( .A1(n12144), .A2(n12143), .A3(n12142), .ZN(n15424) );
  CLKBUF_X1 U11977 ( .A(n15423), .Z(n17144) );
  INV_X1 U11978 ( .A(n14795), .ZN(n11156) );
  INV_X1 U11979 ( .A(n14794), .ZN(n11157) );
  INV_X1 U11980 ( .A(n11975), .ZN(n14719) );
  INV_X1 U11981 ( .A(n15647), .ZN(n19376) );
  NAND2_X1 U11982 ( .A1(n12374), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12333) );
  INV_X1 U11983 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16947) );
  OAI21_X1 U11984 ( .B1(n13727), .B2(n13726), .A(n14497), .ZN(n13728) );
  INV_X1 U11985 ( .A(n14501), .ZN(n11112) );
  INV_X1 U11986 ( .A(n14500), .ZN(n11113) );
  XNOR2_X1 U11987 ( .A(n13713), .B(n13712), .ZN(n16795) );
  NAND2_X1 U11988 ( .A1(n18828), .A2(n13735), .ZN(n13713) );
  NOR2_X1 U11989 ( .A1(n16671), .A2(n16670), .ZN(n16672) );
  AOI21_X1 U11990 ( .B1(n12295), .B2(n11041), .A(n11025), .ZN(n11207) );
  NOR2_X1 U11991 ( .A1(n15642), .A2(n15929), .ZN(n15949) );
  INV_X1 U11992 ( .A(n15958), .ZN(n11898) );
  CLKBUF_X1 U11993 ( .A(n15878), .Z(n15879) );
  AND2_X1 U11994 ( .A1(n12146), .A2(n12145), .ZN(n15734) );
  INV_X1 U11995 ( .A(n15394), .ZN(n11867) );
  AND2_X1 U11996 ( .A1(n12306), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16942) );
  OR2_X1 U11997 ( .A1(n14963), .A2(n14958), .ZN(n11110) );
  NOR2_X2 U11998 ( .A1(n15188), .A2(n15189), .ZN(n15187) );
  AND2_X1 U11999 ( .A1(n15760), .A2(n12254), .ZN(n17215) );
  OR2_X1 U12000 ( .A1(n16991), .A2(n16994), .ZN(n17210) );
  OR2_X1 U12001 ( .A1(n11739), .A2(n17232), .ZN(n11740) );
  INV_X1 U12002 ( .A(n14770), .ZN(n11153) );
  INV_X1 U12003 ( .A(n14771), .ZN(n11154) );
  AND2_X1 U12004 ( .A1(n17251), .A2(n17231), .ZN(n17218) );
  OR2_X1 U12005 ( .A1(n17245), .A2(n17242), .ZN(n16991) );
  CLKBUF_X1 U12006 ( .A(n14962), .Z(n15151) );
  AND2_X1 U12007 ( .A1(n12023), .A2(n12022), .ZN(n14767) );
  AND2_X1 U12008 ( .A1(n11007), .A2(n12018), .ZN(n12019) );
  NAND2_X1 U12009 ( .A1(n11150), .A2(n11241), .ZN(n17260) );
  NAND2_X1 U12010 ( .A1(n11710), .A2(n11700), .ZN(n11150) );
  NAND2_X1 U12011 ( .A1(n17260), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17259) );
  NAND2_X1 U12012 ( .A1(n14105), .A2(n11182), .ZN(n14109) );
  NOR2_X1 U12013 ( .A1(n11183), .A2(n14108), .ZN(n11182) );
  INV_X1 U12014 ( .A(n14104), .ZN(n11183) );
  INV_X1 U12015 ( .A(n19558), .ZN(n19539) );
  AND2_X1 U12016 ( .A1(n19408), .A2(n19467), .ZN(n19538) );
  INV_X1 U12017 ( .A(n19491), .ZN(n19489) );
  NAND2_X2 U12018 ( .A1(n11287), .A2(n11286), .ZN(n19753) );
  NAND2_X1 U12019 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19571), .ZN(n19839) );
  OR2_X1 U12020 ( .A1(n19402), .A2(n19408), .ZN(n19381) );
  AND3_X1 U12021 ( .A1(n15265), .A2(n15264), .A3(n15263), .ZN(n15784) );
  NOR2_X1 U12022 ( .A1(n20735), .A2(n11037), .ZN(n20750) );
  NAND2_X1 U12023 ( .A1(n11127), .A2(n20723), .ZN(n11126) );
  OR2_X1 U12024 ( .A1(n20724), .A2(n20765), .ZN(n11127) );
  AND2_X1 U12025 ( .A1(n11122), .A2(n20592), .ZN(n20681) );
  NOR2_X1 U12026 ( .A1(n20681), .A2(n20682), .ZN(n20695) );
  NOR2_X1 U12027 ( .A1(n20654), .A2(n20765), .ZN(n20655) );
  NOR2_X1 U12028 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n20620), .ZN(n20630) );
  NOR2_X1 U12029 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n20580), .ZN(n20600) );
  INV_X1 U12030 ( .A(n20614), .ZN(n20598) );
  NAND2_X1 U12031 ( .A1(n20341), .A2(n20340), .ZN(n20349) );
  AND2_X1 U12032 ( .A1(n13846), .A2(n11090), .ZN(n11088) );
  INV_X1 U12033 ( .A(n18515), .ZN(n18516) );
  XNOR2_X1 U12034 ( .A(n11132), .B(n11131), .ZN(n20615) );
  NAND2_X1 U12035 ( .A1(n18295), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11132) );
  AOI21_X1 U12036 ( .B1(n21275), .B2(n21274), .A(n18468), .ZN(n18293) );
  NAND2_X1 U12037 ( .A1(n18267), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n18266) );
  NOR2_X1 U12038 ( .A1(n18210), .A2(n21246), .ZN(n21275) );
  NOR2_X2 U12039 ( .A1(n18303), .A2(n18307), .ZN(n20584) );
  INV_X1 U12040 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n20519) );
  NAND2_X1 U12041 ( .A1(n14043), .A2(n20414), .ZN(n18126) );
  INV_X1 U12042 ( .A(n20451), .ZN(n18358) );
  NAND2_X1 U12043 ( .A1(n14039), .A2(n18369), .ZN(n21041) );
  INV_X1 U12044 ( .A(n14037), .ZN(n14035) );
  NAND2_X1 U12045 ( .A1(n18105), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18327) );
  INV_X1 U12046 ( .A(n18421), .ZN(n18428) );
  NAND2_X1 U12047 ( .A1(n18218), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n21269) );
  NOR2_X1 U12048 ( .A1(n21102), .A2(n21308), .ZN(n11138) );
  NOR2_X1 U12049 ( .A1(n21319), .A2(n14041), .ZN(n18211) );
  NAND2_X1 U12050 ( .A1(n18211), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n18210) );
  NAND2_X1 U12051 ( .A1(n21207), .A2(n14040), .ZN(n21320) );
  NAND2_X1 U12052 ( .A1(n13879), .A2(n18152), .ZN(n18225) );
  NOR2_X1 U12053 ( .A1(n18225), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18224) );
  NOR2_X2 U12054 ( .A1(n21368), .A2(n21231), .ZN(n21215) );
  NOR2_X1 U12055 ( .A1(n13877), .A2(n11143), .ZN(n18311) );
  NAND2_X1 U12056 ( .A1(n11145), .A2(n11144), .ZN(n11143) );
  NAND2_X1 U12057 ( .A1(n18258), .A2(n21398), .ZN(n11144) );
  NAND2_X1 U12058 ( .A1(n13875), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11145) );
  INV_X1 U12059 ( .A(n21308), .ZN(n18258) );
  NAND2_X1 U12060 ( .A1(n18317), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n21200) );
  NOR2_X1 U12061 ( .A1(n21200), .A2(n21213), .ZN(n21360) );
  INV_X1 U12062 ( .A(n18327), .ZN(n21362) );
  INV_X1 U12063 ( .A(n21345), .ZN(n21361) );
  INV_X1 U12064 ( .A(n21041), .ZN(n21155) );
  NAND3_X1 U12065 ( .A1(n13832), .A2(n13831), .A3(n13830), .ZN(n14085) );
  NAND2_X1 U12066 ( .A1(n18401), .A2(n14034), .ZN(n18384) );
  XNOR2_X1 U12067 ( .A(n13867), .B(n13868), .ZN(n18390) );
  NOR2_X1 U12068 ( .A1(n18390), .A2(n21135), .ZN(n18389) );
  INV_X1 U12069 ( .A(n13861), .ZN(n11141) );
  NAND2_X1 U12070 ( .A1(n11086), .A2(n14030), .ZN(n18407) );
  NAND2_X1 U12071 ( .A1(n18419), .A2(n18420), .ZN(n11086) );
  NAND2_X1 U12072 ( .A1(n18407), .A2(n18408), .ZN(n18406) );
  NAND2_X1 U12073 ( .A1(n18443), .A2(n14028), .ZN(n18436) );
  NAND2_X1 U12074 ( .A1(n18437), .A2(n18436), .ZN(n18435) );
  XNOR2_X1 U12075 ( .A(n14026), .B(n21083), .ZN(n18445) );
  NAND2_X1 U12076 ( .A1(n18445), .A2(n18444), .ZN(n18443) );
  OAI21_X1 U12077 ( .B1(n14005), .B2(n14004), .A(n14003), .ZN(n21471) );
  NOR2_X1 U12078 ( .A1(n13959), .A2(n13958), .ZN(n14057) );
  NOR2_X2 U12079 ( .A1(n20275), .A2(n17299), .ZN(n21368) );
  NAND2_X1 U12080 ( .A1(n14024), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18462) );
  INV_X2 U12081 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21006) );
  INV_X1 U12082 ( .A(n21007), .ZN(n21025) );
  NOR2_X1 U12083 ( .A1(n13918), .A2(n13917), .ZN(n19262) );
  INV_X1 U12084 ( .A(n19259), .ZN(n19173) );
  NAND2_X1 U12085 ( .A1(n19216), .A2(n13986), .ZN(n21476) );
  OR2_X1 U12086 ( .A1(n13644), .A2(n13648), .ZN(n21761) );
  NOR2_X1 U12087 ( .A1(n20070), .A2(n21737), .ZN(n21759) );
  NOR2_X1 U12088 ( .A1(n20067), .A2(n21717), .ZN(n21739) );
  INV_X1 U12089 ( .A(n21777), .ZN(n21754) );
  AND2_X1 U12090 ( .A1(n13647), .A2(n13641), .ZN(n21724) );
  NAND2_X1 U12091 ( .A1(n16136), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21776) );
  AND2_X1 U12092 ( .A1(n16136), .A2(n15162), .ZN(n21782) );
  AND2_X1 U12093 ( .A1(n15161), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15162) );
  INV_X1 U12094 ( .A(n21776), .ZN(n21748) );
  INV_X1 U12095 ( .A(n16415), .ZN(n13632) );
  OAI21_X1 U12096 ( .B1(n15175), .B2(n13626), .A(n13625), .ZN(n16246) );
  OR2_X1 U12097 ( .A1(n14807), .A2(n11020), .ZN(n13625) );
  OR2_X1 U12098 ( .A1(n15216), .A2(n21813), .ZN(n13626) );
  CLKBUF_X1 U12099 ( .A(n15868), .Z(n16298) );
  INV_X1 U12100 ( .A(n16265), .ZN(n16295) );
  NOR2_X1 U12101 ( .A1(n15509), .A2(n11057), .ZN(n11224) );
  NOR2_X1 U12102 ( .A1(n16248), .A2(n14812), .ZN(n15920) );
  NAND2_X1 U12103 ( .A1(n14809), .A2(n14808), .ZN(n16273) );
  INV_X1 U12104 ( .A(n15920), .ZN(n15944) );
  NAND2_X1 U12105 ( .A1(n11038), .A2(n13620), .ZN(n13621) );
  OAI21_X1 U12106 ( .B1(n15908), .B2(n15907), .A(n15906), .ZN(n16403) );
  INV_X1 U12107 ( .A(n16504), .ZN(n21600) );
  NAND2_X1 U12108 ( .A1(n13100), .A2(n14862), .ZN(n16453) );
  INV_X1 U12109 ( .A(n16526), .ZN(n16468) );
  INV_X1 U12110 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n22076) );
  INV_X1 U12111 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n22039) );
  INV_X1 U12112 ( .A(n13146), .ZN(n16583) );
  INV_X1 U12113 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14894) );
  OAI211_X1 U12114 ( .C1(n21967), .C2(n22106), .A(n22045), .B(n21966), .ZN(
        n22311) );
  INV_X1 U12115 ( .A(n22321), .ZN(n22323) );
  OAI211_X1 U12116 ( .C1(n21983), .C2(n21982), .A(n22045), .B(n21981), .ZN(
        n22324) );
  OAI21_X1 U12117 ( .B1(n15812), .B2(n15811), .A(n22094), .ZN(n15853) );
  OR2_X1 U12118 ( .A1(n15124), .A2(n22082), .ZN(n22010) );
  INV_X1 U12119 ( .A(n22010), .ZN(n22335) );
  OAI211_X1 U12120 ( .C1(n22343), .C2(n22072), .A(n22045), .B(n22022), .ZN(
        n22345) );
  AND2_X1 U12121 ( .A1(n22033), .A2(n22029), .ZN(n22354) );
  OAI211_X1 U12122 ( .C1(n22368), .C2(n22072), .A(n22094), .B(n22071), .ZN(
        n22370) );
  INV_X1 U12123 ( .A(n22380), .ZN(n22367) );
  OAI211_X1 U12124 ( .C1(n22382), .C2(n22095), .A(n22094), .B(n22093), .ZN(
        n22385) );
  NOR2_X2 U12125 ( .A1(n22112), .A2(n22082), .ZN(n22384) );
  INV_X1 U12126 ( .A(n22075), .ZN(n22108) );
  INV_X1 U12127 ( .A(n22141), .ZN(n22147) );
  INV_X1 U12128 ( .A(n22172), .ZN(n22179) );
  INV_X1 U12129 ( .A(n22236), .ZN(n22242) );
  INV_X1 U12130 ( .A(n22267), .ZN(n22273) );
  NOR2_X2 U12131 ( .A1(n22112), .A2(n22054), .ZN(n22393) );
  INV_X1 U12132 ( .A(n22373), .ZN(n22389) );
  NOR2_X1 U12133 ( .A1(n14870), .A2(n22072), .ZN(n21807) );
  AND2_X1 U12134 ( .A1(n17379), .A2(n17378), .ZN(n21814) );
  AND2_X1 U12135 ( .A1(n21798), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21800) );
  INV_X1 U12136 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n21798) );
  INV_X1 U12137 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n21804) );
  INV_X1 U12138 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21847) );
  INV_X1 U12139 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19470) );
  XNOR2_X1 U12140 ( .A(n13722), .B(n13721), .ZN(n18838) );
  NOR2_X1 U12141 ( .A1(n18822), .A2(n12364), .ZN(n18833) );
  INV_X1 U12142 ( .A(n18803), .ZN(n18853) );
  OR2_X1 U12143 ( .A1(n18850), .A2(n19459), .ZN(n18621) );
  INV_X1 U12144 ( .A(n18897), .ZN(n18861) );
  AND2_X1 U12145 ( .A1(n12409), .A2(n12402), .ZN(n18811) );
  OR2_X1 U12146 ( .A1(n12068), .A2(n12067), .ZN(n15184) );
  INV_X1 U12147 ( .A(n11487), .ZN(n15682) );
  AND2_X1 U12148 ( .A1(n14494), .A2(n18592), .ZN(n16651) );
  OR2_X1 U12149 ( .A1(n16689), .A2(n19380), .ZN(n16698) );
  XNOR2_X1 U12150 ( .A(n11188), .B(n14492), .ZN(n16077) );
  NAND2_X1 U12151 ( .A1(n11187), .A2(n14464), .ZN(n11188) );
  NAND2_X1 U12152 ( .A1(n11186), .A2(n14464), .ZN(n16631) );
  INV_X1 U12153 ( .A(n11187), .ZN(n11186) );
  INV_X1 U12154 ( .A(n11171), .ZN(n16676) );
  AND2_X1 U12155 ( .A1(n16771), .A2(n16765), .ZN(n19367) );
  AOI21_X2 U12156 ( .B1(n15264), .B2(n14714), .A(n18914), .ZN(n19374) );
  INV_X1 U12157 ( .A(n16765), .ZN(n19585) );
  INV_X1 U12158 ( .A(n19374), .ZN(n19579) );
  BUF_X1 U12159 ( .A(n17721), .Z(n17735) );
  CLKBUF_X1 U12160 ( .A(n17727), .Z(n17736) );
  OR2_X1 U12161 ( .A1(n14522), .A2(n17648), .ZN(n14528) );
  INV_X1 U12162 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17645) );
  INV_X1 U12163 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17622) );
  INV_X1 U12164 ( .A(n17648), .ZN(n17668) );
  NAND2_X1 U12165 ( .A1(n17658), .A2(n17324), .ZN(n17651) );
  AND2_X1 U12166 ( .A1(n17658), .A2(n17660), .ZN(n17647) );
  INV_X1 U12167 ( .A(n17658), .ZN(n17661) );
  NAND2_X1 U12168 ( .A1(n15994), .A2(n18876), .ZN(n16003) );
  NAND2_X1 U12169 ( .A1(n15993), .A2(n17204), .ZN(n16004) );
  NAND2_X1 U12170 ( .A1(n11198), .A2(n13704), .ZN(n16820) );
  AOI21_X1 U12171 ( .B1(n16840), .B2(n12321), .A(n16807), .ZN(n16832) );
  INV_X1 U12172 ( .A(n18885), .ZN(n17204) );
  AND2_X1 U12173 ( .A1(n17227), .A2(n11938), .ZN(n17222) );
  NAND2_X1 U12174 ( .A1(n17641), .A2(n11738), .ZN(n16990) );
  NAND2_X1 U12175 ( .A1(n17247), .A2(n17246), .ZN(n17641) );
  AND2_X1 U12176 ( .A1(n11711), .A2(n11665), .ZN(n15765) );
  INV_X1 U12177 ( .A(n15521), .ZN(n11589) );
  AND2_X1 U12178 ( .A1(n11947), .A2(n11824), .ZN(n18879) );
  INV_X1 U12179 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19424) );
  OR2_X1 U12180 ( .A1(n14733), .A2(n14732), .ZN(n19455) );
  INV_X1 U12181 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19518) );
  INV_X1 U12182 ( .A(n19549), .ZN(n19564) );
  NAND2_X1 U12183 ( .A1(n19470), .A2(n19459), .ZN(n19549) );
  NAND2_X1 U12184 ( .A1(n15363), .A2(n12001), .ZN(n15470) );
  AOI221_X1 U12185 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n17329), .C1(n18901), .C2(
        n17329), .A(n19571), .ZN(n17696) );
  INV_X1 U12186 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17330) );
  CLKBUF_X1 U12187 ( .A(n11913), .Z(n15786) );
  OR2_X1 U12188 ( .A1(n14788), .A2(n14789), .ZN(n14790) );
  AND2_X1 U12189 ( .A1(n15781), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n18906) );
  CLKBUF_X1 U12190 ( .A(n11809), .Z(n18870) );
  NAND2_X1 U12191 ( .A1(n19539), .A2(n19538), .ZN(n19933) );
  INV_X1 U12192 ( .A(n19933), .ZN(n19936) );
  NOR2_X1 U12193 ( .A1(n19558), .A2(n19517), .ZN(n19929) );
  OAI22_X1 U12194 ( .A1(n19514), .A2(n19510), .B1(n19567), .B2(n19509), .ZN(
        n19916) );
  NAND2_X1 U12195 ( .A1(n19489), .A2(n19538), .ZN(n19818) );
  INV_X1 U12196 ( .A(n19899), .ZN(n19813) );
  INV_X1 U12197 ( .A(n19808), .ZN(n19881) );
  OAI21_X1 U12198 ( .B1(n19442), .B2(n19441), .A(n19440), .ZN(n19875) );
  OAI22_X1 U12199 ( .A1(n19442), .A2(n19438), .B1(n19567), .B2(n19437), .ZN(
        n19876) );
  INV_X1 U12200 ( .A(n19706), .ZN(n19708) );
  AOI21_X1 U12201 ( .B1(n19848), .B2(n19571), .A(n19393), .ZN(n19851) );
  INV_X1 U12202 ( .A(n19826), .ZN(n19832) );
  INV_X1 U12203 ( .A(n19791), .ZN(n19783) );
  INV_X1 U12204 ( .A(n19666), .ZN(n19668) );
  INV_X1 U12205 ( .A(n19950), .ZN(n19845) );
  INV_X1 U12206 ( .A(n19622), .ZN(n19626) );
  INV_X1 U12207 ( .A(n19854), .ZN(n19796) );
  INV_X1 U12208 ( .A(n19533), .ZN(n19563) );
  OR2_X1 U12209 ( .A1(n19381), .A2(n19455), .ZN(n19950) );
  OR4_X1 U12210 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), 
        .A3(P2_STATEBS16_REG_SCAN_IN), .A4(n17326), .ZN(n18897) );
  INV_X1 U12211 ( .A(n18592), .ZN(n18914) );
  OR2_X1 U12212 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n17321), .ZN(n17770) );
  INV_X1 U12213 ( .A(n20339), .ZN(n20341) );
  OAI21_X1 U12214 ( .B1(n21439), .B2(n21440), .A(n18073), .ZN(n20339) );
  INV_X1 U12215 ( .A(n11122), .ZN(n20680) );
  INV_X1 U12216 ( .A(n11124), .ZN(n20638) );
  INV_X1 U12217 ( .A(n11125), .ZN(n20637) );
  AND2_X1 U12218 ( .A1(n20614), .A2(n20613), .ZN(n20626) );
  AOI21_X1 U12219 ( .B1(n20616), .B2(n20617), .A(n20615), .ZN(n20618) );
  NOR2_X2 U12220 ( .A1(n21477), .A2(n20349), .ZN(n20614) );
  NAND2_X1 U12221 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n20612), .ZN(n20770) );
  AND2_X1 U12222 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n18012), .ZN(n18042) );
  AOI211_X1 U12223 ( .C1(n13919), .C2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n13967), .B(n13966), .ZN(n13968) );
  INV_X1 U12224 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17835) );
  NAND2_X1 U12225 ( .A1(n20902), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n20928) );
  NOR2_X1 U12226 ( .A1(n20944), .A2(n20943), .ZN(n20942) );
  NOR2_X1 U12227 ( .A1(n20802), .A2(n20817), .ZN(n20815) );
  INV_X1 U12228 ( .A(n14012), .ZN(n20850) );
  INV_X1 U12229 ( .A(n20959), .ZN(n20966) );
  INV_X1 U12230 ( .A(n14024), .ZN(n20991) );
  OAI21_X1 U12231 ( .B1(n20797), .B2(n20796), .A(n21475), .ZN(n20985) );
  INV_X1 U12232 ( .A(n20792), .ZN(n20795) );
  NAND2_X1 U12233 ( .A1(n20804), .A2(n20828), .ZN(n20990) );
  INV_X1 U12234 ( .A(n20853), .ZN(n20986) );
  NOR2_X1 U12237 ( .A1(n20297), .A2(n20285), .ZN(n20328) );
  CLKBUF_X2 U12239 ( .A(n20297), .Z(n20333) );
  INV_X1 U12240 ( .A(n18185), .ZN(n18165) );
  NOR3_X2 U12241 ( .A1(P3_STATEBS16_REG_SCAN_IN), .A2(n18439), .A3(n20997), 
        .ZN(n18297) );
  INV_X1 U12242 ( .A(n18238), .ZN(n18240) );
  INV_X1 U12243 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18307) );
  INV_X1 U12244 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18375) );
  NOR2_X2 U12245 ( .A1(n21297), .A2(n18467), .ZN(n18379) );
  INV_X1 U12246 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20436) );
  NAND2_X1 U12247 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18421) );
  NAND2_X1 U12248 ( .A1(n19259), .A2(n18979), .ZN(n19054) );
  NAND2_X1 U12249 ( .A1(n18305), .A2(n18304), .ZN(n18450) );
  INV_X1 U12250 ( .A(n18450), .ZN(n18460) );
  OAI21_X1 U12251 ( .B1(n18079), .B2(P3_STATE2_REG_0__SCAN_IN), .A(n21505), 
        .ZN(n18463) );
  INV_X1 U12252 ( .A(n18423), .ZN(n18468) );
  INV_X1 U12253 ( .A(n18457), .ZN(n18467) );
  NOR2_X1 U12254 ( .A1(n14076), .A2(n14075), .ZN(n21372) );
  NOR2_X1 U12255 ( .A1(n21430), .A2(n21437), .ZN(n21271) );
  INV_X1 U12256 ( .A(n21410), .ZN(n21383) );
  INV_X1 U12257 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21450) );
  INV_X1 U12258 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18968) );
  INV_X1 U12259 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17316) );
  AOI21_X1 U12260 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n20337), .A(n17306), 
        .ZN(n21040) );
  INV_X1 U12261 ( .A(n21040), .ZN(n21038) );
  INV_X1 U12262 ( .A(n20606), .ZN(n21485) );
  INV_X1 U12263 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n21488) );
  INV_X1 U12264 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n21881) );
  NOR2_X1 U12265 ( .A1(n21871), .A2(n18561), .ZN(n18571) );
  AOI21_X1 U12267 ( .B1(n16412), .B2(n13631), .A(n14539), .ZN(n14540) );
  OAI21_X1 U12268 ( .B1(n13119), .B2(n21789), .A(n11027), .ZN(P1_U2968) );
  OAI21_X1 U12269 ( .B1(n16431), .B2(n21789), .A(n13701), .ZN(n13702) );
  NOR2_X1 U12270 ( .A1(n13700), .A2(n13699), .ZN(n13701) );
  NOR2_X1 U12271 ( .A1(n13117), .A2(n13116), .ZN(n13118) );
  NAND2_X1 U12272 ( .A1(n11230), .A2(n13115), .ZN(n13116) );
  AOI21_X1 U12273 ( .B1(n15993), .B2(n17672), .A(n13748), .ZN(n13751) );
  INV_X1 U12274 ( .A(n16049), .ZN(n16050) );
  AOI211_X1 U12275 ( .C1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n17115), .A(
        n17114), .B(n17113), .ZN(n17116) );
  AOI21_X1 U12276 ( .B1(n20776), .B2(n20775), .A(n20774), .ZN(n20780) );
  AND2_X1 U12277 ( .A1(n14095), .A2(n14094), .ZN(n14096) );
  INV_X1 U12278 ( .A(n11383), .ZN(n11527) );
  BUF_X2 U12279 ( .A(n13919), .Z(n18046) );
  INV_X2 U12280 ( .A(n11832), .ZN(n12398) );
  OR2_X1 U12281 ( .A1(n11173), .A2(n14372), .ZN(n11024) );
  OR2_X1 U12282 ( .A1(n12310), .A2(n12309), .ZN(n11025) );
  NAND3_X1 U12283 ( .A1(n11200), .A2(n11661), .A3(n12006), .ZN(n12231) );
  XNOR2_X1 U12284 ( .A(n12753), .B(n21955), .ZN(n13146) );
  AND2_X1 U12285 ( .A1(n12199), .A2(n12196), .ZN(n11026) );
  AND2_X1 U12286 ( .A1(n13619), .A2(n13618), .ZN(n11027) );
  AND2_X1 U12287 ( .A1(n11528), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n11028) );
  AND2_X2 U12288 ( .A1(n14467), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11559) );
  NOR2_X1 U12289 ( .A1(n21021), .A2(n13761), .ZN(n13841) );
  NAND2_X1 U12290 ( .A1(n11194), .A2(n16817), .ZN(n16794) );
  OR2_X1 U12291 ( .A1(n12262), .A2(n12261), .ZN(n11029) );
  AND2_X1 U12292 ( .A1(n16186), .A2(n13379), .ZN(n16228) );
  XOR2_X1 U12293 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n13884), .Z(
        n11030) );
  NAND2_X1 U12294 ( .A1(n18310), .A2(n21308), .ZN(n18152) );
  NAND2_X1 U12295 ( .A1(n12159), .A2(n12158), .ZN(n12415) );
  AND2_X1 U12296 ( .A1(n11980), .A2(n11979), .ZN(n11031) );
  NOR3_X1 U12297 ( .A1(n18224), .A2(n18151), .A3(n21329), .ZN(n11032) );
  AND2_X1 U12298 ( .A1(n15887), .A2(n12854), .ZN(n11033) );
  AND2_X1 U12299 ( .A1(n16186), .A2(n11222), .ZN(n16171) );
  NAND2_X1 U12300 ( .A1(n12159), .A2(n11164), .ZN(n16737) );
  AND3_X1 U12301 ( .A1(n11102), .A2(n11800), .A3(n19753), .ZN(n11035) );
  NAND2_X1 U12302 ( .A1(n11618), .A2(n11617), .ZN(n11666) );
  AND3_X1 U12303 ( .A1(n11269), .A2(n11259), .A3(n11098), .ZN(n11036) );
  XNOR2_X1 U12304 ( .A(n14916), .B(n14126), .ZN(n14788) );
  INV_X1 U12305 ( .A(n12562), .ZN(n12574) );
  NAND2_X1 U12306 ( .A1(n11207), .A2(n11206), .ZN(n16835) );
  AND2_X1 U12307 ( .A1(n14109), .A2(n14945), .ZN(n14918) );
  OR2_X1 U12308 ( .A1(n16103), .A2(n11212), .ZN(n11038) );
  AND3_X1 U12309 ( .A1(n11400), .A2(n11401), .A3(n11185), .ZN(n11039) );
  OR2_X1 U12310 ( .A1(n15992), .A2(n17648), .ZN(n11040) );
  AND2_X1 U12311 ( .A1(n12294), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11041) );
  INV_X1 U12312 ( .A(n11173), .ZN(n16674) );
  NAND2_X1 U12313 ( .A1(n11171), .A2(n11170), .ZN(n11173) );
  NAND2_X1 U12314 ( .A1(n16304), .A2(n16343), .ZN(n16302) );
  NAND2_X1 U12315 ( .A1(n16501), .A2(n13084), .ZN(n11042) );
  AND2_X1 U12316 ( .A1(n12854), .A2(n11042), .ZN(n11043) );
  NAND2_X1 U12317 ( .A1(n12702), .A2(n12701), .ZN(n12753) );
  NOR2_X1 U12318 ( .A1(n16737), .A2(n16738), .ZN(n16728) );
  INV_X1 U12319 ( .A(n14397), .ZN(n11180) );
  AND2_X1 U12320 ( .A1(n14396), .A2(n11228), .ZN(n14397) );
  AND2_X1 U12321 ( .A1(n12291), .A2(n12292), .ZN(n12312) );
  NAND2_X1 U12322 ( .A1(n16655), .A2(n16656), .ZN(n14500) );
  AND2_X1 U12323 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11044) );
  OR2_X1 U12324 ( .A1(n21307), .A2(n21306), .ZN(n11045) );
  OR2_X1 U12325 ( .A1(n14510), .A2(n16060), .ZN(n11046) );
  AND2_X1 U12326 ( .A1(n12001), .A2(n11161), .ZN(n11047) );
  INV_X1 U12327 ( .A(n13165), .ZN(n13137) );
  INV_X1 U12328 ( .A(n13137), .ZN(n13599) );
  AND2_X1 U12329 ( .A1(n15183), .A2(n15184), .ZN(n15396) );
  NAND2_X1 U12330 ( .A1(n12010), .A2(n12181), .ZN(n11973) );
  NAND2_X1 U12331 ( .A1(n14967), .A2(n14965), .ZN(n11048) );
  NOR2_X2 U12332 ( .A1(n12349), .A2(n17659), .ZN(n12342) );
  NAND2_X1 U12333 ( .A1(n16691), .A2(n16690), .ZN(n16683) );
  NAND2_X1 U12334 ( .A1(n15396), .A2(n14195), .ZN(n15638) );
  NOR2_X1 U12335 ( .A1(n15789), .A2(n11219), .ZN(n15862) );
  NOR2_X1 U12336 ( .A1(n15789), .A2(n13299), .ZN(n15834) );
  NOR2_X1 U12337 ( .A1(n15509), .A2(n15443), .ZN(n11049) );
  OR2_X1 U12338 ( .A1(n18126), .A2(n18137), .ZN(n11050) );
  AND2_X1 U12339 ( .A1(n14937), .A2(n14936), .ZN(n14935) );
  NAND2_X1 U12340 ( .A1(n15861), .A2(n15964), .ZN(n15965) );
  AND2_X1 U12341 ( .A1(n14935), .A2(n15135), .ZN(n15134) );
  NAND2_X1 U12342 ( .A1(n14771), .A2(n11155), .ZN(n14794) );
  OR2_X1 U12343 ( .A1(n15642), .A2(n11159), .ZN(n15948) );
  OR2_X1 U12344 ( .A1(n15423), .A2(n15424), .ZN(n15422) );
  NOR2_X1 U12345 ( .A1(n15105), .A2(n15198), .ZN(n15197) );
  AND2_X1 U12346 ( .A1(n15486), .A2(n15456), .ZN(n15455) );
  AND2_X1 U12347 ( .A1(n12221), .A2(n12222), .ZN(n12220) );
  AND2_X1 U12348 ( .A1(n11004), .A2(n11224), .ZN(n15565) );
  BUF_X1 U12349 ( .A(n11481), .Z(n14791) );
  NAND2_X1 U12350 ( .A1(n20351), .A2(n21392), .ZN(n21102) );
  OR2_X1 U12351 ( .A1(n12320), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11051) );
  AND2_X1 U12352 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n11052) );
  OR2_X1 U12353 ( .A1(n15424), .A2(n15734), .ZN(n11053) );
  BUF_X1 U12354 ( .A(n11527), .Z(n19793) );
  OR2_X1 U12355 ( .A1(n15642), .A2(n11158), .ZN(n16619) );
  OR2_X1 U12356 ( .A1(n11048), .A2(n14956), .ZN(n11054) );
  OR2_X1 U12357 ( .A1(n12867), .A2(n20182), .ZN(n11055) );
  INV_X1 U12358 ( .A(n11974), .ZN(n17666) );
  OR2_X1 U12359 ( .A1(n11538), .A2(n11537), .ZN(n11974) );
  NAND2_X1 U12360 ( .A1(n11467), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11056) );
  OR2_X1 U12361 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n13597) );
  AND2_X2 U12362 ( .A1(n14481), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14152) );
  INV_X1 U12363 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15285) );
  OR2_X1 U12364 ( .A1(n14133), .A2(n11048), .ZN(n14955) );
  OR2_X1 U12365 ( .A1(n14962), .A2(n14963), .ZN(n14957) );
  NOR2_X1 U12366 ( .A1(n11154), .A2(n11153), .ZN(n14768) );
  INV_X1 U12367 ( .A(n14372), .ZN(n11172) );
  NAND2_X1 U12368 ( .A1(n12558), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13163) );
  INV_X1 U12369 ( .A(n13163), .ZN(n13312) );
  NAND2_X2 U12370 ( .A1(n17371), .A2(n15174), .ZN(n21789) );
  INV_X1 U12371 ( .A(n21789), .ZN(n20188) );
  INV_X1 U12372 ( .A(n16675), .ZN(n11170) );
  AND4_X1 U12373 ( .A1(n13202), .A2(n13201), .A3(n13200), .A4(n13199), .ZN(
        n11057) );
  AND2_X1 U12374 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n20344) );
  INV_X1 U12375 ( .A(n16060), .ZN(n11163) );
  NAND2_X1 U12376 ( .A1(n19633), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11058) );
  INV_X1 U12377 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11129) );
  INV_X1 U12378 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11131) );
  INV_X1 U12379 ( .A(n19837), .ZN(n19571) );
  OAI22_X2 U12380 ( .A1(n20260), .A2(n15414), .B1(n17510), .B2(n15413), .ZN(
        n22175) );
  INV_X1 U12381 ( .A(n22383), .ZN(n11059) );
  INV_X1 U12382 ( .A(n11059), .ZN(n11060) );
  INV_X1 U12383 ( .A(n22144), .ZN(n11061) );
  INV_X1 U12384 ( .A(n11061), .ZN(n11062) );
  INV_X1 U12385 ( .A(n22302), .ZN(n11063) );
  INV_X1 U12386 ( .A(n11063), .ZN(n11064) );
  INV_X1 U12387 ( .A(n22239), .ZN(n11065) );
  INV_X1 U12388 ( .A(n11065), .ZN(n11066) );
  INV_X1 U12389 ( .A(n22208), .ZN(n11067) );
  INV_X1 U12390 ( .A(n11067), .ZN(n11068) );
  INV_X1 U12391 ( .A(n22096), .ZN(n11069) );
  INV_X1 U12392 ( .A(n11069), .ZN(n11070) );
  INV_X1 U12393 ( .A(n22118), .ZN(n11071) );
  INV_X1 U12394 ( .A(n11071), .ZN(n11072) );
  INV_X1 U12395 ( .A(n22213), .ZN(n11073) );
  INV_X1 U12396 ( .A(n11073), .ZN(n11074) );
  INV_X1 U12397 ( .A(n22275), .ZN(n11075) );
  INV_X1 U12398 ( .A(n11075), .ZN(n11076) );
  INV_X1 U12399 ( .A(n22392), .ZN(n11077) );
  INV_X1 U12400 ( .A(n11077), .ZN(n11078) );
  INV_X1 U12401 ( .A(n22149), .ZN(n11079) );
  INV_X1 U12402 ( .A(n11079), .ZN(n11080) );
  INV_X1 U12403 ( .A(n22307), .ZN(n11081) );
  INV_X1 U12404 ( .A(n11081), .ZN(n11082) );
  INV_X1 U12405 ( .A(n22244), .ZN(n11083) );
  INV_X1 U12406 ( .A(n11083), .ZN(n11084) );
  CLKBUF_X1 U12407 ( .A(n21462), .Z(n11085) );
  OAI22_X2 U12408 ( .A1(n20266), .A2(n15414), .B1(n17414), .B2(n15413), .ZN(
        n22270) );
  OAI22_X2 U12409 ( .A1(n20243), .A2(n15414), .B1(n15100), .B2(n15413), .ZN(
        n22181) );
  NAND2_X1 U12410 ( .A1(n20186), .A2(n15865), .ZN(n15413) );
  NOR2_X2 U12411 ( .A1(n15412), .A2(n15096), .ZN(n22212) );
  OR3_X1 U12412 ( .A1(n22072), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n15079), 
        .ZN(n15412) );
  AND4_X1 U12413 ( .A1(n13843), .A2(n13844), .A3(n11087), .A4(n13845), .ZN(
        n11089) );
  NAND4_X1 U12414 ( .A1(n11089), .A2(n13849), .A3(n13850), .A4(n11088), .ZN(
        n14024) );
  INV_X2 U12415 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n21001) );
  AND2_X4 U12416 ( .A1(n11266), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14300) );
  AND2_X2 U12417 ( .A1(n11258), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11266) );
  NOR4_X1 U12418 ( .A1(n11273), .A2(n11097), .A3(n11044), .A4(n11028), .ZN(
        n11096) );
  NAND3_X1 U12419 ( .A1(n11260), .A2(n11274), .A3(n11270), .ZN(n11097) );
  NAND2_X1 U12420 ( .A1(n11101), .A2(n11099), .ZN(n11102) );
  NAND2_X1 U12421 ( .A1(n11100), .A2(n14715), .ZN(n11099) );
  INV_X1 U12422 ( .A(n19674), .ZN(n11804) );
  NAND2_X1 U12423 ( .A1(n11104), .A2(n20182), .ZN(n16357) );
  NOR2_X2 U12424 ( .A1(n16320), .A2(n16319), .ZN(n12877) );
  AND2_X2 U12425 ( .A1(n11109), .A2(n11055), .ZN(n16320) );
  NAND2_X1 U12426 ( .A1(n11111), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12724) );
  XNOR2_X1 U12427 ( .A(n11111), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14914) );
  NAND3_X1 U12428 ( .A1(n12880), .A2(n12878), .A3(n12879), .ZN(n13119) );
  INV_X1 U12429 ( .A(n16666), .ZN(n11114) );
  NAND2_X1 U12430 ( .A1(n14924), .A2(n14923), .ZN(n12752) );
  NAND2_X1 U12431 ( .A1(n14897), .A2(n14896), .ZN(n11117) );
  NAND2_X1 U12432 ( .A1(n16616), .A2(n16617), .ZN(n11909) );
  NAND2_X1 U12433 ( .A1(n15878), .A2(n11898), .ZN(n16693) );
  NAND2_X1 U12434 ( .A1(n15455), .A2(n15579), .ZN(n15578) );
  NOR2_X2 U12435 ( .A1(n15485), .A2(n15484), .ZN(n15486) );
  NAND2_X1 U12436 ( .A1(n11868), .A2(n11867), .ZN(n15485) );
  NAND3_X1 U12437 ( .A1(n12220), .A2(n12233), .A3(n12188), .ZN(n12198) );
  NAND3_X1 U12438 ( .A1(n11194), .A2(n16817), .A3(n11197), .ZN(n16798) );
  INV_X1 U12439 ( .A(n11127), .ZN(n20725) );
  INV_X1 U12440 ( .A(n11126), .ZN(n20734) );
  NOR2_X1 U12441 ( .A1(n20713), .A2(n20714), .ZN(n20724) );
  NOR2_X2 U12442 ( .A1(n18227), .A2(n18215), .ZN(n18267) );
  AND2_X2 U12443 ( .A1(n18185), .A2(n11133), .ZN(n18197) );
  NAND2_X1 U12444 ( .A1(n11134), .A2(n18247), .ZN(n18291) );
  NOR2_X1 U12445 ( .A1(n11134), .A2(n18248), .ZN(n18257) );
  NAND2_X1 U12446 ( .A1(n11135), .A2(n11045), .ZN(n21309) );
  NAND2_X1 U12447 ( .A1(n21296), .A2(n11138), .ZN(n11135) );
  NAND2_X1 U12448 ( .A1(n11136), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n21300) );
  AND3_X2 U12449 ( .A1(n18220), .A2(n13882), .A3(n11139), .ZN(n13883) );
  INV_X1 U12450 ( .A(n11142), .ZN(n13862) );
  NOR2_X1 U12451 ( .A1(n18426), .A2(n18425), .ZN(n18424) );
  NOR2_X1 U12452 ( .A1(n18462), .A2(n18453), .ZN(n18452) );
  NAND2_X2 U12453 ( .A1(n21006), .A2(n20344), .ZN(n21012) );
  INV_X1 U12454 ( .A(n11976), .ZN(n11151) );
  NAND2_X2 U12455 ( .A1(n15362), .A2(n15361), .ZN(n15363) );
  NOR2_X2 U12456 ( .A1(n14510), .A2(n11162), .ZN(n16702) );
  NOR2_X2 U12457 ( .A1(n15423), .A2(n11053), .ZN(n15735) );
  NAND2_X1 U12458 ( .A1(n16679), .A2(n16680), .ZN(n11175) );
  NAND2_X2 U12459 ( .A1(n11175), .A2(n11174), .ZN(n11171) );
  INV_X1 U12460 ( .A(n11181), .ZN(n16658) );
  INV_X1 U12461 ( .A(n14440), .ZN(n11179) );
  NAND2_X1 U12462 ( .A1(n14105), .A2(n14104), .ZN(n11184) );
  AND2_X1 U12463 ( .A1(n11184), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n14946) );
  NAND2_X2 U12464 ( .A1(n11934), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11464) );
  OR2_X2 U12466 ( .A1(n14133), .A2(n11054), .ZN(n15190) );
  INV_X1 U12467 ( .A(n14133), .ZN(n14966) );
  NOR2_X2 U12468 ( .A1(n15946), .A2(n15947), .ZN(n16691) );
  NAND3_X1 U12469 ( .A1(n11191), .A2(n19380), .A3(n11391), .ZN(n11397) );
  NAND2_X2 U12470 ( .A1(n11311), .A2(n11310), .ZN(n14715) );
  NAND3_X1 U12471 ( .A1(n11192), .A2(n11348), .A3(n11408), .ZN(n11410) );
  NAND4_X1 U12472 ( .A1(n11192), .A2(n11348), .A3(n11411), .A4(n11408), .ZN(
        n11809) );
  AND2_X1 U12473 ( .A1(n19674), .A2(n14715), .ZN(n11193) );
  NOR2_X1 U12474 ( .A1(n16795), .A2(n16805), .ZN(n11197) );
  AND2_X2 U12475 ( .A1(n11208), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15269) );
  NAND2_X1 U12476 ( .A1(n11210), .A2(n12641), .ZN(n11211) );
  NOR2_X1 U12477 ( .A1(n16103), .A2(n16104), .ZN(n13686) );
  NOR2_X2 U12478 ( .A1(n16103), .A2(n11213), .ZN(n14532) );
  NOR2_X1 U12479 ( .A1(n15509), .A2(n11226), .ZN(n11223) );
  INV_X1 U12480 ( .A(n15566), .ZN(n13235) );
  XNOR2_X1 U12481 ( .A(n12231), .B(n11715), .ZN(n12169) );
  AOI21_X1 U12482 ( .B1(n18613), .B2(n14116), .A(n14115), .ZN(n14782) );
  NOR2_X1 U12483 ( .A1(n11490), .A2(n18613), .ZN(n11638) );
  NAND2_X1 U12484 ( .A1(n12564), .A2(n12563), .ZN(n12568) );
  NAND2_X1 U12485 ( .A1(n12560), .A2(n12559), .ZN(n12564) );
  XNOR2_X2 U12486 ( .A(n21083), .B(n13853), .ZN(n21077) );
  NOR2_X2 U12487 ( .A1(n21078), .A2(n21077), .ZN(n18447) );
  AND3_X4 U12488 ( .A1(n15229), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n12447), .ZN(n13238) );
  NAND2_X1 U12489 ( .A1(n12954), .A2(n12580), .ZN(n13096) );
  AOI22_X1 U12490 ( .A1(n12685), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12518), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12487) );
  OAI21_X1 U12491 ( .B1(n11801), .B2(n11969), .A(n11377), .ZN(n11386) );
  AOI211_X2 U12492 ( .C1(n17007), .C2(n18876), .A(n17006), .B(n17005), .ZN(
        n17010) );
  NAND2_X1 U12493 ( .A1(n14461), .A2(n14460), .ZN(n14462) );
  OAI211_X1 U12494 ( .C1(n16777), .C2(n18885), .A(n16048), .B(n16047), .ZN(
        n16049) );
  AND2_X1 U12495 ( .A1(n15977), .A2(n15976), .ZN(n15978) );
  AND4_X1 U12496 ( .A1(n12506), .A2(n12505), .A3(n12504), .A4(n12503), .ZN(
        n12512) );
  NAND2_X1 U12497 ( .A1(n14453), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11276) );
  NAND2_X1 U12498 ( .A1(n11464), .A2(n11418), .ZN(n11419) );
  AND3_X1 U12499 ( .A1(n11331), .A2(n11330), .A3(n11374), .ZN(n11334) );
  AND3_X1 U12500 ( .A1(n14398), .A2(n14417), .A3(n14393), .ZN(n11228) );
  AOI21_X1 U12501 ( .B1(n16044), .B2(n18763), .A(n13670), .ZN(n13671) );
  AND2_X1 U12502 ( .A1(n16003), .A2(n16002), .ZN(n11229) );
  OR3_X1 U12503 ( .A1(n16410), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n16310), .ZN(n11230) );
  INV_X1 U12504 ( .A(n11968), .ZN(n11982) );
  OR2_X1 U12505 ( .A1(n13668), .A2(n13680), .ZN(n11231) );
  AND2_X1 U12506 ( .A1(n14496), .A2(n14495), .ZN(n11232) );
  AND2_X1 U12507 ( .A1(n14528), .A2(n14527), .ZN(n11233) );
  NAND3_X2 U12508 ( .A1(n13894), .A2(n13893), .A3(n13892), .ZN(n20351) );
  INV_X1 U12509 ( .A(n11528), .ZN(n14230) );
  AND2_X1 U12510 ( .A1(n13286), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11234) );
  AND4_X1 U12511 ( .A1(n16484), .A2(n16367), .A3(n16456), .A4(n20183), .ZN(
        n11235) );
  AND2_X1 U12512 ( .A1(n12871), .A2(n12870), .ZN(n11236) );
  NOR2_X1 U12513 ( .A1(n12229), .A2(n15694), .ZN(n11237) );
  NAND2_X1 U12514 ( .A1(n20137), .A2(n15867), .ZN(n16247) );
  INV_X1 U12515 ( .A(n16247), .ZN(n13631) );
  AND2_X1 U12516 ( .A1(n11574), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11238) );
  AND3_X1 U12517 ( .A1(n11278), .A2(n11277), .A3(n11276), .ZN(n11239) );
  AND4_X1 U12518 ( .A1(n11656), .A2(n11655), .A3(n11654), .A4(n11653), .ZN(
        n11240) );
  AND2_X1 U12519 ( .A1(n11709), .A2(n11708), .ZN(n11241) );
  NOR2_X1 U12520 ( .A1(n12442), .A2(n12441), .ZN(n11242) );
  OR2_X1 U12521 ( .A1(n12702), .A2(n12701), .ZN(n11243) );
  INV_X1 U12522 ( .A(n16863), .ZN(n12294) );
  INV_X1 U12523 ( .A(n18561), .ZN(n21831) );
  AND2_X1 U12524 ( .A1(n11586), .A2(n11993), .ZN(n11244) );
  INV_X1 U12525 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12331) );
  INV_X1 U12526 ( .A(n11705), .ZN(n11664) );
  AND2_X1 U12527 ( .A1(n21279), .A2(n21275), .ZN(n11245) );
  INV_X1 U12528 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n13871) );
  INV_X1 U12529 ( .A(n16382), .ZN(n12866) );
  NAND2_X1 U12530 ( .A1(n20137), .A2(n14811), .ZN(n16237) );
  NAND2_X1 U12531 ( .A1(n12417), .A2(n12416), .ZN(n11246) );
  OR2_X1 U12532 ( .A1(n21246), .A2(n21247), .ZN(n11247) );
  AND4_X1 U12533 ( .A1(n11695), .A2(n11694), .A3(n11693), .A4(n11692), .ZN(
        n11248) );
  AND2_X1 U12534 ( .A1(n11312), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11249) );
  INV_X1 U12535 ( .A(n18881), .ZN(n12326) );
  AND2_X1 U12536 ( .A1(n12562), .A2(n14745), .ZN(n12904) );
  NOR2_X1 U12537 ( .A1(n16611), .A2(n12202), .ZN(n15976) );
  INV_X1 U12538 ( .A(n15976), .ZN(n13720) );
  INV_X1 U12539 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12330) );
  AND2_X1 U12540 ( .A1(n16046), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11250) );
  INV_X1 U12541 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13712) );
  INV_X1 U12542 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15914) );
  AND3_X1 U12543 ( .A1(n14052), .A2(n14051), .A3(n14050), .ZN(n11251) );
  NAND2_X1 U12544 ( .A1(n18196), .A2(n11018), .ZN(n18305) );
  INV_X1 U12545 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n14101) );
  NAND2_X1 U12546 ( .A1(n14125), .A2(n14124), .ZN(n11252) );
  INV_X1 U12547 ( .A(n13757), .ZN(n15053) );
  NOR2_X1 U12548 ( .A1(n21021), .A2(n20343), .ZN(n13757) );
  INV_X2 U12549 ( .A(n13801), .ZN(n17865) );
  INV_X1 U12550 ( .A(n16187), .ZN(n16235) );
  INV_X1 U12551 ( .A(n16143), .ZN(n16159) );
  INV_X1 U12552 ( .A(n12161), .ZN(n16970) );
  AND2_X1 U12553 ( .A1(n14519), .A2(n14518), .ZN(n11253) );
  INV_X1 U12554 ( .A(n15879), .ZN(n15959) );
  NAND2_X1 U12555 ( .A1(n12240), .A2(n16979), .ZN(n11254) );
  OR3_X2 U12556 ( .A1(n11486), .A2(n11487), .A3(n18613), .ZN(n11632) );
  INV_X1 U12557 ( .A(n11701), .ZN(n11712) );
  AND4_X1 U12558 ( .A1(n12459), .A2(n12458), .A3(n12457), .A4(n12456), .ZN(
        n11255) );
  AND4_X1 U12559 ( .A1(n12511), .A2(n12510), .A3(n12509), .A4(n12508), .ZN(
        n11256) );
  NAND2_X1 U12560 ( .A1(n14273), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n11565) );
  NAND2_X1 U12561 ( .A1(n11638), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11522) );
  OAI22_X1 U12562 ( .A1(n11471), .A2(n11632), .B1(n11633), .B2(n14196), .ZN(
        n11480) );
  NAND2_X1 U12563 ( .A1(n14806), .A2(n12910), .ZN(n12927) );
  AND2_X1 U12564 ( .A1(n12887), .A2(n12886), .ZN(n12901) );
  AOI22_X1 U12565 ( .A1(n12527), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        P1_INSTQUEUE_REG_14__2__SCAN_IN), .B2(n13238), .ZN(n12448) );
  OR2_X1 U12566 ( .A1(n12894), .A2(n12911), .ZN(n12896) );
  NAND2_X1 U12567 ( .A1(n12569), .A2(n14860), .ZN(n12563) );
  INV_X1 U12568 ( .A(n12841), .ZN(n12665) );
  NAND2_X1 U12569 ( .A1(n11750), .A2(n11749), .ZN(n11755) );
  AOI22_X1 U12570 ( .A1(n11341), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11366), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11330) );
  INV_X1 U12571 ( .A(n12187), .ZN(n12188) );
  AND2_X1 U12572 ( .A1(n11660), .A2(n11659), .ZN(n11661) );
  INV_X1 U12573 ( .A(n12767), .ZN(n12765) );
  INV_X1 U12574 ( .A(n16234), .ZN(n13379) );
  OAI21_X1 U12575 ( .B1(n16382), .B2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n15889), .ZN(n12853) );
  OR2_X1 U12576 ( .A1(n12814), .A2(n12813), .ZN(n12829) );
  OR2_X1 U12577 ( .A1(n12622), .A2(n12621), .ZN(n12716) );
  OR2_X1 U12578 ( .A1(n12684), .A2(n12636), .ZN(n12623) );
  AOI21_X1 U12579 ( .B1(n11755), .B2(n11753), .A(n11751), .ZN(n11760) );
  OR2_X1 U12580 ( .A1(n14944), .A2(n14940), .ZN(n14129) );
  NOR2_X1 U12581 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14303) );
  AOI22_X1 U12582 ( .A1(n11369), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11332) );
  AOI22_X1 U12583 ( .A1(n11369), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11307) );
  INV_X1 U12584 ( .A(n11453), .ZN(n11447) );
  INV_X1 U12585 ( .A(n11978), .ZN(n11979) );
  NAND2_X1 U12586 ( .A1(n14791), .A2(n14116), .ZN(n14113) );
  AOI22_X1 U12587 ( .A1(n11369), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11345) );
  INV_X1 U12588 ( .A(n11923), .ZN(n11808) );
  NOR2_X1 U12589 ( .A1(n11020), .A2(n13074), .ZN(n13066) );
  INV_X1 U12590 ( .A(n16144), .ZN(n13461) );
  AND2_X1 U12591 ( .A1(n13554), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13555) );
  INV_X1 U12592 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n13217) );
  AND2_X1 U12593 ( .A1(n13043), .A2(n13042), .ZN(n16238) );
  NOR2_X1 U12594 ( .A1(n16390), .A2(n16392), .ZN(n15889) );
  AND2_X1 U12595 ( .A1(n12598), .A2(n12597), .ZN(n13098) );
  AND2_X1 U12596 ( .A1(n12569), .A2(n13074), .ZN(n12596) );
  INV_X1 U12597 ( .A(n11574), .ZN(n12099) );
  AND4_X1 U12598 ( .A1(n11730), .A2(n11729), .A3(n11728), .A4(n11727), .ZN(
        n11732) );
  NAND2_X1 U12599 ( .A1(n11254), .A2(n12241), .ZN(n12242) );
  INV_X1 U12600 ( .A(n11512), .ZN(n11620) );
  NAND2_X1 U12601 ( .A1(n19055), .A2(n20856), .ZN(n14060) );
  NOR2_X1 U12602 ( .A1(n14060), .A2(n21004), .ZN(n14977) );
  NOR2_X1 U12603 ( .A1(n20351), .A2(n20340), .ZN(n20793) );
  NOR2_X1 U12604 ( .A1(n14078), .A2(n21269), .ZN(n14010) );
  AND2_X1 U12605 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13865), .ZN(
        n13866) );
  AOI211_X1 U12606 ( .C1(n14055), .C2(n14064), .A(n14067), .B(n13992), .ZN(
        n13996) );
  NOR2_X1 U12607 ( .A1(n13516), .A2(n16336), .ZN(n13517) );
  NAND2_X1 U12608 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13147) );
  NAND2_X1 U12609 ( .A1(n12583), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13573) );
  OR2_X1 U12610 ( .A1(n13612), .A2(n16314), .ZN(n13614) );
  NAND2_X1 U12611 ( .A1(n13172), .A2(n13171), .ZN(n15449) );
  NAND2_X1 U12612 ( .A1(n10992), .A2(n16305), .ZN(n16306) );
  NAND2_X1 U12613 ( .A1(n16239), .A2(n16238), .ZN(n16241) );
  NAND2_X1 U12614 ( .A1(n13014), .A2(n15662), .ZN(n13015) );
  OR2_X1 U12615 ( .A1(n12743), .A2(n12742), .ZN(n12747) );
  NAND2_X1 U12616 ( .A1(n12733), .A2(n12732), .ZN(n15081) );
  INV_X1 U12617 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n22066) );
  INV_X1 U12618 ( .A(n14636), .ZN(n11411) );
  NAND2_X1 U12619 ( .A1(n13669), .A2(n11231), .ZN(n13670) );
  INV_X1 U12620 ( .A(n11015), .ZN(n12009) );
  NAND2_X1 U12621 ( .A1(n12247), .A2(n12248), .ZN(n12257) );
  INV_X1 U12622 ( .A(n15192), .ZN(n14134) );
  NAND2_X1 U12623 ( .A1(n14100), .A2(n19459), .ZN(n14118) );
  AND2_X1 U12624 ( .A1(n14106), .A2(n19592), .ZN(n14417) );
  INV_X1 U12625 ( .A(n12099), .ZN(n14295) );
  INV_X1 U12626 ( .A(n13728), .ZN(n13729) );
  NOR2_X2 U12627 ( .A1(n15986), .A2(n15985), .ZN(n16635) );
  INV_X1 U12628 ( .A(n14515), .ZN(n13750) );
  AND2_X1 U12629 ( .A1(n16883), .A2(n12300), .ZN(n16862) );
  INV_X1 U12630 ( .A(n11627), .ZN(n19383) );
  INV_X1 U12631 ( .A(n19174), .ZN(n13982) );
  INV_X1 U12632 ( .A(n17317), .ZN(n17302) );
  INV_X1 U12633 ( .A(n20793), .ZN(n20794) );
  OR3_X1 U12634 ( .A1(n21308), .A2(n18091), .A3(n18090), .ZN(n18178) );
  NOR2_X1 U12635 ( .A1(n20850), .A2(n13851), .ZN(n14023) );
  INV_X1 U12636 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n21720) );
  NOR2_X1 U12637 ( .A1(n20063), .A2(n21712), .ZN(n15915) );
  INV_X1 U12638 ( .A(n16273), .ZN(n16248) );
  NAND2_X1 U12639 ( .A1(n14805), .A2(n14804), .ZN(n14863) );
  INV_X1 U12640 ( .A(n14530), .ZN(n14531) );
  NAND2_X1 U12641 ( .A1(n13480), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13516) );
  NOR2_X1 U12642 ( .A1(n13315), .A2(n21720), .ZN(n13330) );
  INV_X1 U12643 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n21643) );
  NOR2_X1 U12644 ( .A1(n13114), .A2(n13615), .ZN(n13115) );
  OAI21_X1 U12645 ( .B1(n16302), .B2(n16307), .A(n16306), .ZN(n16309) );
  NOR2_X2 U12646 ( .A1(n10955), .A2(n16196), .ZN(n16198) );
  AND2_X1 U12647 ( .A1(n12850), .A2(n16551), .ZN(n16398) );
  INV_X1 U12648 ( .A(n15618), .ZN(n21531) );
  OR2_X1 U12649 ( .A1(n21794), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13609) );
  INV_X1 U12650 ( .A(n15805), .ZN(n15856) );
  INV_X1 U12651 ( .A(n15201), .ZN(n15438) );
  OR2_X1 U12652 ( .A1(n15124), .A2(n22085), .ZN(n21999) );
  NOR2_X1 U12653 ( .A1(n22064), .A2(n21961), .ZN(n22045) );
  INV_X1 U12654 ( .A(n22033), .ZN(n22055) );
  AOI21_X1 U12655 ( .B1(n21511), .B2(n21803), .A(n21807), .ZN(n15079) );
  NOR2_X1 U12656 ( .A1(n22037), .A2(n21961), .ZN(n22094) );
  NOR2_X1 U12657 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n22117) );
  INV_X1 U12658 ( .A(n19581), .ZN(n16766) );
  OAI21_X1 U12659 ( .B1(n14564), .B2(n14563), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n15647) );
  INV_X1 U12660 ( .A(n16788), .ZN(n15983) );
  AND2_X1 U12661 ( .A1(n18720), .A2(n12301), .ZN(n16900) );
  AND2_X1 U12662 ( .A1(n16917), .A2(n16954), .ZN(n16946) );
  NOR2_X1 U12663 ( .A1(n16930), .A2(n17141), .ZN(n16957) );
  OR2_X1 U12664 ( .A1(n11735), .A2(n12202), .ZN(n11739) );
  AND2_X1 U12665 ( .A1(n11937), .A2(n14503), .ZN(n17227) );
  AND2_X1 U12666 ( .A1(n11823), .A2(n18592), .ZN(n11947) );
  INV_X1 U12667 ( .A(n14918), .ZN(n14919) );
  OR2_X1 U12668 ( .A1(n19521), .A2(n19502), .ZN(n19558) );
  INV_X1 U12669 ( .A(n14007), .ZN(n14005) );
  INV_X1 U12670 ( .A(n20771), .ZN(n20772) );
  NOR2_X1 U12671 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n20640), .ZN(n20657) );
  NOR2_X1 U12672 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n20496), .ZN(n20508) );
  INV_X1 U12673 ( .A(n20615), .ZN(n20592) );
  INV_X1 U12674 ( .A(n20787), .ZN(n20757) );
  OAI21_X1 U12675 ( .B1(n17299), .B2(n21445), .A(n14978), .ZN(n20792) );
  NAND2_X1 U12676 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .ZN(n20798) );
  NOR2_X1 U12677 ( .A1(n20795), .A2(n20794), .ZN(n20796) );
  OR2_X1 U12678 ( .A1(n21301), .A2(n21361), .ZN(n21304) );
  AOI21_X1 U12679 ( .B1(n14000), .B2(n14076), .A(n21007), .ZN(n21217) );
  NOR2_X1 U12680 ( .A1(n13877), .A2(n13876), .ZN(n18121) );
  INV_X1 U12681 ( .A(n21334), .ZN(n21392) );
  NOR2_X1 U12682 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n17388), .ZN(n19259) );
  INV_X1 U12683 ( .A(n19016), .ZN(n19261) );
  AND2_X1 U12684 ( .A1(n14695), .A2(n15174), .ZN(n13635) );
  INV_X1 U12685 ( .A(n21761), .ZN(n21773) );
  INV_X1 U12686 ( .A(n21738), .ZN(n21710) );
  INV_X1 U12687 ( .A(n16237), .ZN(n13627) );
  NAND2_X1 U12688 ( .A1(n16161), .A2(n16147), .ZN(n16217) );
  INV_X1 U12689 ( .A(n16246), .ZN(n15926) );
  OR2_X1 U12690 ( .A1(n13686), .A2(n13687), .ZN(n13688) );
  NAND2_X1 U12691 ( .A1(n14863), .A2(n15174), .ZN(n14809) );
  INV_X1 U12692 ( .A(n21951), .ZN(n14854) );
  INV_X1 U12693 ( .A(n21949), .ZN(n21945) );
  INV_X1 U12694 ( .A(n21886), .ZN(n21943) );
  NAND2_X1 U12695 ( .A1(n13435), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13478) );
  INV_X1 U12696 ( .A(n20155), .ZN(n20192) );
  AND2_X1 U12697 ( .A1(n20155), .A2(n20138), .ZN(n20172) );
  OR2_X1 U12698 ( .A1(n14775), .A2(n16468), .ZN(n16513) );
  INV_X1 U12699 ( .A(n21600), .ZN(n21585) );
  INV_X1 U12700 ( .A(n16575), .ZN(n21596) );
  OR2_X1 U12701 ( .A1(n13101), .A2(n16529), .ZN(n15616) );
  INV_X1 U12702 ( .A(n21560), .ZN(n21595) );
  AOI21_X1 U12703 ( .B1(n12961), .B2(n12960), .A(n21813), .ZN(n13100) );
  NAND2_X1 U12704 ( .A1(n21798), .A2(n22072), .ZN(n21794) );
  NOR2_X2 U12705 ( .A1(n21988), .A2(n22058), .ZN(n22317) );
  OR2_X1 U12706 ( .A1(n15087), .A2(n13134), .ZN(n22082) );
  NOR2_X2 U12707 ( .A1(n21988), .A2(n22085), .ZN(n22330) );
  NOR2_X1 U12708 ( .A1(n15124), .A2(n22058), .ZN(n15805) );
  INV_X1 U12709 ( .A(n21999), .ZN(n22337) );
  INV_X1 U12710 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n22105) );
  INV_X1 U12711 ( .A(n22366), .ZN(n22356) );
  AND2_X1 U12712 ( .A1(n13146), .A2(n22013), .ZN(n22033) );
  NOR2_X2 U12713 ( .A1(n22055), .A2(n22054), .ZN(n22369) );
  NOR2_X1 U12714 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15079), .ZN(n15415) );
  OR2_X1 U12715 ( .A1(n15087), .A2(n15123), .ZN(n22058) );
  INV_X1 U12716 ( .A(n22205), .ZN(n22211) );
  INV_X1 U12717 ( .A(n22299), .ZN(n22305) );
  NAND2_X1 U12718 ( .A1(n21956), .A2(n21955), .ZN(n22112) );
  NAND2_X1 U12719 ( .A1(n11799), .A2(n11796), .ZN(n15781) );
  NOR2_X1 U12720 ( .A1(n12410), .A2(n18803), .ZN(n12411) );
  INV_X1 U12721 ( .A(n12404), .ZN(n12319) );
  AND2_X1 U12722 ( .A1(n18589), .A2(n12413), .ZN(n18850) );
  NOR2_X1 U12723 ( .A1(n18589), .A2(n15338), .ZN(n18763) );
  INV_X1 U12724 ( .A(n19408), .ZN(n19423) );
  INV_X1 U12725 ( .A(n16698), .ZN(n16686) );
  INV_X1 U12726 ( .A(n18600), .ZN(n18884) );
  INV_X1 U12727 ( .A(n15427), .ZN(n19369) );
  INV_X1 U12728 ( .A(n14690), .ZN(n14616) );
  INV_X1 U12729 ( .A(n14644), .ZN(n14686) );
  INV_X1 U12730 ( .A(n17651), .ZN(n17672) );
  INV_X1 U12731 ( .A(n15980), .ZN(n15981) );
  OR2_X1 U12732 ( .A1(n18734), .A2(n12202), .ZN(n16893) );
  NOR2_X1 U12733 ( .A1(n16850), .A2(n16851), .ZN(n16956) );
  XNOR2_X1 U12734 ( .A(n11739), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16989) );
  AND2_X1 U12735 ( .A1(n11947), .A2(n11946), .ZN(n18876) );
  XNOR2_X1 U12736 ( .A(n14920), .B(n14919), .ZN(n19521) );
  AND2_X1 U12737 ( .A1(n14941), .A2(n14790), .ZN(n19502) );
  OAI21_X1 U12738 ( .B1(n19942), .B2(n19572), .A(n19571), .ZN(n19947) );
  NOR2_X1 U12739 ( .A1(n19558), .A2(n19557), .ZN(n19943) );
  INV_X1 U12740 ( .A(n19925), .ZN(n19658) );
  OAI21_X1 U12741 ( .B1(n19514), .B2(n19513), .A(n19512), .ZN(n19915) );
  INV_X1 U12742 ( .A(n19912), .ZN(n19914) );
  INV_X1 U12743 ( .A(n19818), .ZN(n19907) );
  NAND2_X1 U12744 ( .A1(n19489), .A2(n19423), .ZN(n19473) );
  OAI21_X1 U12745 ( .B1(n19887), .B2(n19461), .A(n19571), .ZN(n19890) );
  NAND2_X1 U12746 ( .A1(n19408), .A2(n19455), .ZN(n19557) );
  INV_X1 U12747 ( .A(n19879), .ZN(n19870) );
  NAND2_X1 U12748 ( .A1(n19521), .A2(n17692), .ZN(n19445) );
  INV_X1 U12749 ( .A(n19750), .ZN(n19742) );
  INV_X1 U12750 ( .A(n19538), .ZN(n19432) );
  INV_X1 U12751 ( .A(n19926), .ZN(n19944) );
  INV_X1 U12752 ( .A(n19455), .ZN(n19467) );
  AND3_X1 U12753 ( .A1(n17326), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n18592) );
  INV_X1 U12754 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n17321) );
  NAND2_X1 U12755 ( .A1(n20773), .A2(n20772), .ZN(n20774) );
  NAND2_X1 U12756 ( .A1(n20742), .A2(n20741), .ZN(n20743) );
  INV_X1 U12757 ( .A(n20646), .ZN(n20665) );
  NOR2_X1 U12758 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n20548), .ZN(n20576) );
  NOR2_X1 U12759 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n20517), .ZN(n20541) );
  NOR2_X1 U12760 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n20464), .ZN(n20487) );
  NOR2_X1 U12761 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n20439), .ZN(n20459) );
  NOR2_X1 U12762 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n20411), .ZN(n20432) );
  INV_X1 U12763 ( .A(n20770), .ZN(n20708) );
  AND2_X1 U12764 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n18010), .ZN(n17936) );
  NAND4_X1 U12765 ( .A1(n21475), .A2(n20340), .A3(n20351), .A4(n20792), .ZN(
        n18069) );
  INV_X1 U12766 ( .A(n20922), .ZN(n20918) );
  NOR2_X1 U12767 ( .A1(n20861), .A2(n20889), .ZN(n20880) );
  INV_X1 U12768 ( .A(n20934), .ZN(n20949) );
  OR2_X1 U12769 ( .A1(n13788), .A2(n13787), .ZN(n14012) );
  INV_X1 U12770 ( .A(n20990), .ZN(n20978) );
  INV_X1 U12771 ( .A(n19262), .ZN(n20340) );
  INV_X1 U12772 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18397) );
  INV_X1 U12773 ( .A(n18463), .ZN(n18439) );
  NAND2_X2 U12774 ( .A1(n21215), .A2(n21217), .ZN(n21334) );
  INV_X1 U12775 ( .A(n21337), .ZN(n21432) );
  NOR2_X1 U12776 ( .A1(n21102), .A2(n14085), .ZN(n21345) );
  NOR2_X1 U12777 ( .A1(n21430), .A2(n21102), .ZN(n21131) );
  NOR2_X1 U12778 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21488), .ZN(
        n21490) );
  INV_X1 U12779 ( .A(n18573), .ZN(n18567) );
  INV_X1 U12780 ( .A(n19376), .ZN(n19375) );
  INV_X1 U12781 ( .A(n13657), .ZN(n13658) );
  INV_X1 U12782 ( .A(n21724), .ZN(n21788) );
  INV_X1 U12783 ( .A(n21782), .ZN(n21702) );
  INV_X1 U12784 ( .A(n15926), .ZN(n20137) );
  INV_X1 U12785 ( .A(n20164), .ZN(n21716) );
  NAND2_X1 U12786 ( .A1(n20017), .A2(n15178), .ZN(n15555) );
  INV_X1 U12787 ( .A(n20017), .ZN(n20044) );
  NOR2_X1 U12788 ( .A1(n14744), .A2(n14743), .ZN(n21949) );
  INV_X1 U12789 ( .A(n20172), .ZN(n20200) );
  NAND2_X1 U12790 ( .A1(n21789), .A2(n13610), .ZN(n20155) );
  NAND2_X1 U12791 ( .A1(n13100), .A2(n12970), .ZN(n16575) );
  AOI22_X1 U12792 ( .A1(n21965), .A2(n21962), .B1(n22037), .B2(n21967), .ZN(
        n22314) );
  OR2_X1 U12793 ( .A1(n21988), .A2(n22082), .ZN(n22321) );
  AOI22_X1 U12794 ( .A1(n21979), .A2(n21982), .B1(n22037), .B2(n22003), .ZN(
        n22327) );
  AOI22_X1 U12795 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21990), .B1(n21995), 
        .B2(n21991), .ZN(n22334) );
  AOI22_X1 U12796 ( .A1(n22004), .A2(n22008), .B1(n22003), .B2(n22064), .ZN(
        n22341) );
  NAND2_X1 U12797 ( .A1(n22033), .A2(n22014), .ZN(n22353) );
  AOI22_X1 U12798 ( .A1(n22043), .A2(n22040), .B1(n22038), .B2(n22037), .ZN(
        n22360) );
  NAND2_X1 U12799 ( .A1(n22033), .A2(n22032), .ZN(n22366) );
  AOI22_X1 U12800 ( .A1(n22070), .A2(n22067), .B1(n22065), .B2(n22064), .ZN(
        n22374) );
  OR2_X1 U12801 ( .A1(n22112), .A2(n22058), .ZN(n22380) );
  OR2_X1 U12802 ( .A1(n22112), .A2(n22085), .ZN(n22397) );
  INV_X1 U12803 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n22072) );
  OR2_X1 U12804 ( .A1(n15328), .A2(n18914), .ZN(n18589) );
  INV_X1 U12805 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n21819) );
  NAND2_X1 U12806 ( .A1(n16630), .A2(n18811), .ZN(n13684) );
  INV_X1 U12807 ( .A(n18811), .ZN(n18857) );
  INV_X1 U12808 ( .A(n18763), .ZN(n18855) );
  INV_X1 U12809 ( .A(n19502), .ZN(n17692) );
  AND2_X1 U12810 ( .A1(n14785), .A2(n14784), .ZN(n19408) );
  NOR2_X1 U12811 ( .A1(n17710), .A2(n17736), .ZN(n17721) );
  INV_X1 U12812 ( .A(n17710), .ZN(n17738) );
  OR2_X1 U12813 ( .A1(n14581), .A2(n11969), .ZN(n14690) );
  INV_X1 U12814 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17659) );
  NAND2_X1 U12815 ( .A1(n18917), .A2(n13744), .ZN(n17658) );
  INV_X1 U12816 ( .A(n18879), .ZN(n17277) );
  OR2_X1 U12817 ( .A1(n12325), .A2(n12324), .ZN(n18881) );
  INV_X1 U12818 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19523) );
  INV_X1 U12819 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18873) );
  INV_X1 U12820 ( .A(n19943), .ZN(n19940) );
  INV_X1 U12821 ( .A(n19929), .ZN(n19782) );
  NAND2_X1 U12822 ( .A1(n19539), .A2(n19503), .ZN(n19925) );
  NAND2_X1 U12823 ( .A1(n19489), .A2(n19488), .ZN(n19912) );
  OR2_X1 U12824 ( .A1(n19473), .A2(n19467), .ZN(n19905) );
  OR2_X1 U12825 ( .A1(n19473), .A2(n19455), .ZN(n19899) );
  OR2_X1 U12826 ( .A1(n19445), .A2(n19557), .ZN(n19886) );
  OR2_X1 U12827 ( .A1(n19445), .A2(n19432), .ZN(n19808) );
  OR2_X1 U12828 ( .A1(n19445), .A2(n19517), .ZN(n19879) );
  OR2_X1 U12829 ( .A1(n19445), .A2(n19409), .ZN(n19873) );
  OR2_X1 U12830 ( .A1(n19402), .A2(n19432), .ZN(n19860) );
  OR2_X1 U12831 ( .A1(n19381), .A2(n19467), .ZN(n19854) );
  INV_X1 U12832 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n17326) );
  INV_X1 U12833 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n21823) );
  AOI21_X1 U12834 ( .B1(n20745), .B2(n20744), .A(n20743), .ZN(n20748) );
  INV_X1 U12835 ( .A(n20788), .ZN(n20768) );
  NOR2_X1 U12836 ( .A1(n20659), .A2(n17974), .ZN(n17980) );
  INV_X1 U12837 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17818) );
  NAND2_X1 U12838 ( .A1(n20918), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n20917) );
  NOR2_X1 U12839 ( .A1(n13767), .A2(n13766), .ZN(n20832) );
  NOR2_X1 U12840 ( .A1(n13777), .A2(n13776), .ZN(n20840) );
  NOR2_X1 U12841 ( .A1(n21489), .A2(n18516), .ZN(n18525) );
  NAND3_X1 U12842 ( .A1(n17317), .A2(n20348), .A3(n18073), .ZN(n18515) );
  INV_X1 U12843 ( .A(n18379), .ZN(n18287) );
  NOR2_X1 U12844 ( .A1(n18439), .A2(n18329), .ZN(n18459) );
  NAND2_X1 U12845 ( .A1(n14085), .A2(n21131), .ZN(n21337) );
  INV_X1 U12846 ( .A(n14092), .ZN(n21379) );
  INV_X1 U12847 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21435) );
  INV_X1 U12848 ( .A(n21403), .ZN(n21430) );
  INV_X1 U12849 ( .A(n21271), .ZN(n21239) );
  INV_X1 U12850 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21449) );
  AND4_X1 U12851 ( .A1(n21503), .A2(n21474), .A3(n21473), .A4(n21472), .ZN(
        n21499) );
  INV_X1 U12852 ( .A(n21826), .ZN(n17312) );
  INV_X1 U12853 ( .A(n20013), .ZN(n20002) );
  NAND2_X1 U12854 ( .A1(n13634), .A2(n13633), .ZN(P1_U2843) );
  OAI21_X1 U12855 ( .B1(n13119), .B2(n16575), .A(n13118), .ZN(P1_U3000) );
  OAI211_X1 U12856 ( .C1(n16008), .C2(n17670), .A(n13751), .B(n11040), .ZN(
        P2_U2984) );
  INV_X1 U12857 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11258) );
  AND2_X1 U12858 ( .A1(n14484), .A2(n11374), .ZN(n11528) );
  AND2_X4 U12859 ( .A1(n15269), .A2(n11418), .ZN(n11370) );
  AND2_X2 U12861 ( .A1(n14483), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14150) );
  AND2_X4 U12862 ( .A1(n11266), .A2(n15266), .ZN(n11369) );
  NAND2_X1 U12863 ( .A1(n14151), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11260) );
  AND2_X4 U12864 ( .A1(n11261), .A2(n15266), .ZN(n11366) );
  NAND2_X1 U12865 ( .A1(n14152), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11259) );
  AND2_X2 U12866 ( .A1(n10962), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14269) );
  NAND2_X1 U12867 ( .A1(n14269), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11265) );
  NAND2_X1 U12868 ( .A1(n14270), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n11264) );
  NAND2_X1 U12869 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11263) );
  AOI22_X1 U12870 ( .A1(n14273), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11262) );
  AND4_X1 U12871 ( .A1(n11265), .A2(n11264), .A3(n11263), .A4(n11262), .ZN(
        n11275) );
  AND2_X1 U12872 ( .A1(n11266), .A2(n14303), .ZN(n14210) );
  NOR2_X1 U12873 ( .A1(n11418), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11267) );
  AOI22_X1 U12874 ( .A1(n14210), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n14288), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11270) );
  AND2_X4 U12875 ( .A1(n11271), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11365) );
  NAND2_X1 U12876 ( .A1(n14480), .A2(n11374), .ZN(n15306) );
  NAND2_X1 U12877 ( .A1(n14287), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n11269) );
  AND2_X4 U12878 ( .A1(n11268), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14467) );
  AND2_X4 U12879 ( .A1(n11271), .A2(n15266), .ZN(n14453) );
  NAND2_X1 U12880 ( .A1(n14253), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n11272) );
  OAI21_X1 U12881 ( .B1(n14107), .B2(n14285), .A(n11272), .ZN(n11273) );
  NAND3_X1 U12882 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11768) );
  NOR2_X1 U12883 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n11768), .ZN(
        n11574) );
  NAND2_X1 U12884 ( .A1(n11574), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11274) );
  INV_X1 U12885 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11471) );
  AOI22_X1 U12886 ( .A1(n11369), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11280) );
  AOI22_X1 U12887 ( .A1(n11341), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11366), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11279) );
  AOI22_X1 U12888 ( .A1(n11370), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14467), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11278) );
  NAND3_X1 U12889 ( .A1(n11280), .A2(n11279), .A3(n11239), .ZN(n11287) );
  AOI22_X1 U12890 ( .A1(n14453), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11365), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11282) );
  AOI22_X1 U12891 ( .A1(n11370), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14467), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11281) );
  AND3_X1 U12892 ( .A1(n11282), .A2(n11281), .A3(n11374), .ZN(n11285) );
  AOI22_X1 U12893 ( .A1(n10961), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11366), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11284) );
  AOI22_X1 U12894 ( .A1(n11369), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11283) );
  NAND3_X1 U12895 ( .A1(n11285), .A2(n11284), .A3(n11283), .ZN(n11286) );
  INV_X1 U12896 ( .A(n19753), .ZN(n11798) );
  AOI22_X1 U12897 ( .A1(n14453), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11365), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11290) );
  AOI22_X1 U12898 ( .A1(n14452), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11366), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11289) );
  AOI22_X1 U12899 ( .A1(n11370), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14467), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11288) );
  NAND3_X1 U12900 ( .A1(n11290), .A2(n11289), .A3(n11288), .ZN(n11292) );
  AOI22_X1 U12901 ( .A1(n11369), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11296) );
  AOI22_X1 U12902 ( .A1(n11370), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n14467), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11295) );
  AOI22_X1 U12903 ( .A1(n10961), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11366), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11294) );
  AOI22_X1 U12904 ( .A1(n14453), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11365), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11293) );
  NAND4_X1 U12905 ( .A1(n11296), .A2(n11295), .A3(n11294), .A4(n11293), .ZN(
        n11297) );
  NAND2_X1 U12906 ( .A1(n11297), .A2(n11374), .ZN(n11298) );
  AOI22_X1 U12907 ( .A1(n14453), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11365), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11303) );
  AOI22_X1 U12908 ( .A1(n11369), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11302) );
  AOI22_X1 U12909 ( .A1(n11341), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11366), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11301) );
  AOI22_X1 U12910 ( .A1(n11370), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n14467), .ZN(n11300) );
  NAND4_X1 U12911 ( .A1(n11303), .A2(n11302), .A3(n11301), .A4(n11300), .ZN(
        n11304) );
  AOI22_X1 U12912 ( .A1(n14453), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11365), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11308) );
  AOI22_X1 U12913 ( .A1(n11341), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11366), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11306) );
  AOI22_X1 U12914 ( .A1(n11370), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14467), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11305) );
  NAND4_X1 U12915 ( .A1(n11308), .A2(n11307), .A3(n11306), .A4(n11305), .ZN(
        n11309) );
  AOI22_X1 U12916 ( .A1(n11370), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14467), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11312) );
  AOI22_X1 U12917 ( .A1(n10961), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11366), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11315) );
  AOI22_X1 U12918 ( .A1(n14453), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11365), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11314) );
  AOI22_X1 U12919 ( .A1(n11369), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11313) );
  NAND4_X1 U12920 ( .A1(n11249), .A2(n11315), .A3(n11314), .A4(n11313), .ZN(
        n11322) );
  AOI22_X1 U12921 ( .A1(n14453), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11365), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11317) );
  AOI22_X1 U12922 ( .A1(n11370), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14467), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11316) );
  AND3_X1 U12923 ( .A1(n11317), .A2(n11316), .A3(n11374), .ZN(n11320) );
  AOI22_X1 U12924 ( .A1(n11369), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11319) );
  AOI22_X1 U12925 ( .A1(n11341), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11366), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11318) );
  NAND3_X1 U12926 ( .A1(n11320), .A2(n11319), .A3(n11318), .ZN(n11321) );
  AOI22_X1 U12927 ( .A1(n11370), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14467), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11325) );
  AOI22_X1 U12928 ( .A1(n14453), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11365), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11324) );
  AOI22_X1 U12929 ( .A1(n11369), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11323) );
  NAND3_X1 U12930 ( .A1(n11329), .A2(n11328), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11336) );
  AOI22_X1 U12931 ( .A1(n11370), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14467), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11331) );
  AOI22_X1 U12932 ( .A1(n14453), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11365), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11333) );
  NAND3_X1 U12933 ( .A1(n11334), .A2(n11333), .A3(n11332), .ZN(n11335) );
  AND2_X2 U12934 ( .A1(n11336), .A2(n11335), .ZN(n11916) );
  AOI22_X1 U12935 ( .A1(n11369), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11340) );
  AOI22_X1 U12936 ( .A1(n11370), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14467), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11339) );
  AOI22_X1 U12937 ( .A1(n10961), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11366), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11338) );
  AOI22_X1 U12938 ( .A1(n14453), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11365), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11337) );
  NAND4_X1 U12939 ( .A1(n11340), .A2(n11339), .A3(n11338), .A4(n11337), .ZN(
        n11347) );
  AOI22_X1 U12940 ( .A1(n11370), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14467), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11344) );
  AOI22_X1 U12941 ( .A1(n11341), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11366), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11343) );
  AOI22_X1 U12942 ( .A1(n14453), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11365), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11342) );
  NAND4_X1 U12943 ( .A1(n11345), .A2(n11344), .A3(n11343), .A4(n11342), .ZN(
        n11346) );
  MUX2_X2 U12944 ( .A(n11347), .B(n11346), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11392) );
  AOI22_X1 U12945 ( .A1(n11369), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11352) );
  AOI22_X1 U12946 ( .A1(n11370), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14467), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11351) );
  AOI22_X1 U12947 ( .A1(n14452), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11366), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11350) );
  AOI22_X1 U12948 ( .A1(n14453), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11365), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11349) );
  NAND4_X1 U12949 ( .A1(n11352), .A2(n11351), .A3(n11350), .A4(n11349), .ZN(
        n11358) );
  AOI22_X1 U12950 ( .A1(n10961), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11366), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11356) );
  AOI22_X1 U12951 ( .A1(n11370), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14467), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11355) );
  AOI22_X1 U12952 ( .A1(n11369), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11354) );
  AOI22_X1 U12953 ( .A1(n14453), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11365), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11353) );
  NAND4_X1 U12954 ( .A1(n11356), .A2(n11355), .A3(n11354), .A4(n11353), .ZN(
        n11357) );
  MUX2_X2 U12955 ( .A(n11358), .B(n11357), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n14636) );
  AOI22_X1 U12956 ( .A1(n14453), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11365), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11360) );
  AOI22_X1 U12957 ( .A1(n11370), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14467), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11359) );
  AOI22_X1 U12958 ( .A1(n11369), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11362) );
  AOI22_X1 U12959 ( .A1(n14452), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11366), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11361) );
  NAND3_X1 U12960 ( .A1(n11363), .A2(n11362), .A3(n11361), .ZN(n11364) );
  AOI22_X1 U12961 ( .A1(n14453), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11365), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11368) );
  AOI22_X1 U12962 ( .A1(n14452), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11366), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11367) );
  AND2_X1 U12963 ( .A1(n11368), .A2(n11367), .ZN(n11373) );
  AOI22_X1 U12964 ( .A1(n11369), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11372) );
  AOI22_X1 U12965 ( .A1(n11370), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14467), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11371) );
  NAND3_X1 U12966 ( .A1(n11373), .A2(n11372), .A3(n11371), .ZN(n11375) );
  INV_X1 U12967 ( .A(n11785), .ZN(n11378) );
  INV_X2 U12968 ( .A(n11392), .ZN(n11377) );
  NAND2_X1 U12969 ( .A1(n11391), .A2(n14715), .ZN(n11967) );
  NOR2_X1 U12970 ( .A1(n11967), .A2(n19592), .ZN(n11380) );
  NAND2_X1 U12971 ( .A1(n11926), .A2(n11380), .ZN(n11433) );
  NAND4_X1 U12972 ( .A1(n19674), .A2(n11392), .A3(n14715), .A4(n19753), .ZN(
        n11402) );
  NOR2_X2 U12973 ( .A1(n11402), .A2(n11801), .ZN(n11404) );
  NAND2_X1 U12974 ( .A1(n11404), .A2(n14636), .ZN(n12436) );
  INV_X1 U12975 ( .A(n12436), .ZN(n11382) );
  NAND2_X1 U12976 ( .A1(n11382), .A2(n10958), .ZN(n11388) );
  NAND3_X1 U12977 ( .A1(n11386), .A2(n11921), .A3(n11385), .ZN(n11420) );
  INV_X1 U12978 ( .A(n11420), .ZN(n11387) );
  NAND2_X1 U12979 ( .A1(n11387), .A2(n11923), .ZN(n11912) );
  NAND3_X1 U12980 ( .A1(n11389), .A2(n11388), .A3(n11912), .ZN(n11390) );
  INV_X1 U12981 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n17662) );
  NAND3_X1 U12982 ( .A1(n11801), .A2(n19674), .A3(n11800), .ZN(n11807) );
  NAND2_X1 U12983 ( .A1(n11975), .A2(n11804), .ZN(n11810) );
  NAND3_X1 U12984 ( .A1(n11807), .A2(n14715), .A3(n11810), .ZN(n11919) );
  MUX2_X1 U12985 ( .A(n11397), .B(n11919), .S(n11392), .Z(n11415) );
  INV_X1 U12986 ( .A(n11412), .ZN(n11393) );
  NAND3_X1 U12987 ( .A1(n11415), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n11393), 
        .ZN(n11401) );
  NOR2_X1 U12988 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11467) );
  INV_X1 U12989 ( .A(n11467), .ZN(n18891) );
  NAND2_X1 U12990 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11395) );
  NAND2_X1 U12991 ( .A1(n18891), .A2(n11395), .ZN(n11396) );
  AOI21_X1 U12992 ( .B1(n11461), .B2(P2_REIP_REG_0__SCAN_IN), .A(n11396), .ZN(
        n11400) );
  INV_X1 U12993 ( .A(n11923), .ZN(n11398) );
  INV_X1 U12994 ( .A(n11402), .ZN(n11403) );
  NAND3_X1 U12995 ( .A1(n13741), .A2(n19753), .A3(n11969), .ZN(n11406) );
  INV_X1 U12996 ( .A(n11404), .ZN(n11405) );
  INV_X1 U12997 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n11407) );
  NAND2_X1 U12998 ( .A1(n11410), .A2(n11409), .ZN(n11930) );
  NAND3_X1 U12999 ( .A1(n11412), .A2(n11930), .A3(n11411), .ZN(n11413) );
  NAND2_X1 U13000 ( .A1(n11415), .A2(n11414), .ZN(n11416) );
  NAND2_X1 U13001 ( .A1(n11466), .A2(n11419), .ZN(n11426) );
  NAND2_X1 U13002 ( .A1(n11419), .A2(n11394), .ZN(n11421) );
  NAND2_X1 U13003 ( .A1(n11421), .A2(n15280), .ZN(n11424) );
  NOR2_X1 U13004 ( .A1(n11808), .A2(n11407), .ZN(n11423) );
  AOI21_X1 U13005 ( .B1(n11424), .B2(n11423), .A(n11422), .ZN(n11425) );
  NAND2_X1 U13006 ( .A1(n11426), .A2(n11425), .ZN(n11441) );
  INV_X1 U13007 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n11430) );
  NAND2_X1 U13008 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11429) );
  NAND2_X1 U13009 ( .A1(n11461), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11428) );
  OAI211_X1 U13010 ( .C1(n11464), .C2(n11430), .A(n11429), .B(n11428), .ZN(
        n11431) );
  NAND2_X1 U13011 ( .A1(n12436), .A2(n11809), .ZN(n11943) );
  INV_X1 U13012 ( .A(n11943), .ZN(n11432) );
  NAND2_X1 U13013 ( .A1(n11433), .A2(n11432), .ZN(n11913) );
  XNOR2_X2 U13014 ( .A(n11449), .B(n11450), .ZN(n11472) );
  OAI21_X2 U13015 ( .B1(n11470), .B2(n11472), .A(n11446), .ZN(n11439) );
  AOI21_X1 U13016 ( .B1(n11407), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n11434) );
  INV_X1 U13017 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n12173) );
  NAND2_X1 U13018 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11436) );
  NAND2_X1 U13019 ( .A1(n11461), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11435) );
  OAI211_X1 U13020 ( .C1(n11464), .C2(n12173), .A(n11436), .B(n11435), .ZN(
        n11437) );
  XNOR2_X1 U13021 ( .A(n11453), .B(n11451), .ZN(n11438) );
  XNOR2_X2 U13022 ( .A(n11439), .B(n11438), .ZN(n11481) );
  INV_X1 U13023 ( .A(n11440), .ZN(n11443) );
  INV_X1 U13024 ( .A(n11441), .ZN(n11442) );
  NAND2_X1 U13025 ( .A1(n11443), .A2(n11442), .ZN(n11444) );
  NAND2_X1 U13026 ( .A1(n11481), .A2(n18884), .ZN(n11486) );
  NAND2_X1 U13027 ( .A1(n11446), .A2(n11453), .ZN(n11445) );
  NAND2_X1 U13028 ( .A1(n11445), .A2(n11451), .ZN(n11459) );
  INV_X1 U13029 ( .A(n11446), .ZN(n11448) );
  NAND2_X1 U13030 ( .A1(n11448), .A2(n11447), .ZN(n11458) );
  NAND2_X1 U13031 ( .A1(n11450), .A2(n11449), .ZN(n11456) );
  INV_X1 U13032 ( .A(n11451), .ZN(n11452) );
  NAND2_X1 U13033 ( .A1(n11453), .A2(n11452), .ZN(n11455) );
  NAND3_X1 U13034 ( .A1(n11456), .A2(n11455), .A3(n11454), .ZN(n11457) );
  INV_X1 U13035 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n15684) );
  NAND2_X1 U13036 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11463) );
  BUF_X4 U13037 ( .A(n11461), .Z(n12390) );
  NAND2_X1 U13038 ( .A1(n12390), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11462) );
  OAI211_X1 U13039 ( .C1(n11464), .C2(n15684), .A(n11462), .B(n11463), .ZN(
        n11465) );
  NAND2_X1 U13040 ( .A1(n11466), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11469) );
  NAND2_X1 U13041 ( .A1(n11467), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11468) );
  XNOR2_X2 U13042 ( .A(n11828), .B(n11827), .ZN(n11825) );
  XNOR2_X2 U13043 ( .A(n11826), .B(n11825), .ZN(n11491) );
  BUF_X4 U13044 ( .A(n11491), .Z(n11487) );
  XNOR2_X2 U13045 ( .A(n11472), .B(n11470), .ZN(n18613) );
  OR3_X2 U13046 ( .A1(n11486), .A2(n11487), .A3(n11489), .ZN(n11633) );
  INV_X1 U13047 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14196) );
  INV_X2 U13048 ( .A(n11481), .ZN(n16033) );
  INV_X1 U13049 ( .A(n11472), .ZN(n11473) );
  NAND2_X1 U13050 ( .A1(n11473), .A2(n18600), .ZN(n11497) );
  INV_X1 U13051 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11475) );
  AND2_X1 U13052 ( .A1(n11472), .A2(n18600), .ZN(n11476) );
  NAND2_X2 U13053 ( .A1(n11487), .A2(n11474), .ZN(n11628) );
  INV_X1 U13054 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14376) );
  OAI22_X1 U13055 ( .A1(n11629), .A2(n11475), .B1(n11628), .B2(n14376), .ZN(
        n11479) );
  OR3_X4 U13056 ( .A1(n16033), .A2(n11487), .A3(n11492), .ZN(n19494) );
  INV_X1 U13057 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14382) );
  INV_X1 U13058 ( .A(n11497), .ZN(n11477) );
  INV_X1 U13059 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14373) );
  OAI22_X1 U13060 ( .A1(n19494), .A2(n14382), .B1(n11627), .B2(n14373), .ZN(
        n11478) );
  OR2_X2 U13061 ( .A1(n11491), .A2(n11481), .ZN(n11498) );
  NOR2_X2 U13062 ( .A1(n11498), .A2(n11492), .ZN(n19550) );
  OR2_X1 U13063 ( .A1(n18613), .A2(n18600), .ZN(n11495) );
  NOR2_X2 U13064 ( .A1(n11498), .A2(n11495), .ZN(n11517) );
  AOI22_X1 U13065 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19550), .B1(
        n11517), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11485) );
  AND2_X1 U13066 ( .A1(n18613), .A2(n18884), .ZN(n11482) );
  INV_X1 U13067 ( .A(n11482), .ZN(n11483) );
  NOR2_X2 U13068 ( .A1(n11498), .A2(n11483), .ZN(n11621) );
  AOI22_X1 U13069 ( .A1(n19439), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11621), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11484) );
  AND2_X1 U13070 ( .A1(n11485), .A2(n11484), .ZN(n11505) );
  INV_X1 U13071 ( .A(n11486), .ZN(n11488) );
  NAND2_X1 U13072 ( .A1(n11488), .A2(n11487), .ZN(n11490) );
  NOR2_X2 U13073 ( .A1(n11490), .A2(n11489), .ZN(n19395) );
  AOI22_X1 U13074 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19395), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11504) );
  INV_X1 U13075 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11494) );
  NAND2_X2 U13076 ( .A1(n11487), .A2(n16033), .ZN(n11496) );
  INV_X1 U13077 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11493) );
  OAI22_X1 U13078 ( .A1(n11494), .A2(n11624), .B1(n19447), .B2(n11493), .ZN(
        n11502) );
  INV_X1 U13080 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11500) );
  NOR2_X2 U13081 ( .A1(n11498), .A2(n11497), .ZN(n11619) );
  NAND2_X1 U13082 ( .A1(n11619), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11499) );
  OAI21_X1 U13083 ( .B1(n11512), .B2(n11500), .A(n11499), .ZN(n11501) );
  NOR2_X1 U13084 ( .A1(n11502), .A2(n11501), .ZN(n11503) );
  NAND4_X1 U13085 ( .A1(n11506), .A2(n11505), .A3(n11504), .A4(n11503), .ZN(
        n11507) );
  MUX2_X2 U13086 ( .A(n12002), .B(n11507), .S(n11969), .Z(n11582) );
  INV_X1 U13087 ( .A(n11582), .ZN(n11580) );
  AOI22_X1 U13088 ( .A1(n19450), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11619), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11516) );
  INV_X1 U13089 ( .A(n11624), .ZN(n11508) );
  INV_X1 U13090 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14335) );
  INV_X1 U13091 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14326) );
  OAI22_X1 U13092 ( .A1(n19494), .A2(n14335), .B1(n11627), .B2(n14326), .ZN(
        n11511) );
  INV_X1 U13093 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11509) );
  NOR2_X1 U13094 ( .A1(n11632), .A2(n11509), .ZN(n11510) );
  NOR2_X1 U13095 ( .A1(n11511), .A2(n11510), .ZN(n11514) );
  INV_X1 U13096 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14135) );
  INV_X1 U13097 ( .A(n11633), .ZN(n19478) );
  AOI22_X1 U13098 ( .A1(n11620), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n19478), .ZN(n11513) );
  NAND4_X1 U13099 ( .A1(n11516), .A2(n11515), .A3(n11514), .A4(n11513), .ZN(
        n11526) );
  INV_X1 U13100 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11519) );
  INV_X1 U13101 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14329) );
  OAI211_X1 U13102 ( .C1(n11629), .C2(n11519), .A(n11969), .B(n11518), .ZN(
        n11520) );
  AOI21_X1 U13103 ( .B1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n11517), .A(
        n11520), .ZN(n11524) );
  AOI22_X1 U13104 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19550), .B1(
        n11621), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11523) );
  NAND2_X1 U13105 ( .A1(n19395), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11521) );
  NAND4_X1 U13106 ( .A1(n11524), .A2(n11523), .A3(n11522), .A4(n11521), .ZN(
        n11525) );
  AOI22_X1 U13107 ( .A1(n14288), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14273), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11532) );
  AOI22_X1 U13108 ( .A1(n14210), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11531) );
  AOI22_X1 U13109 ( .A1(n14269), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14150), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11530) );
  AOI22_X1 U13110 ( .A1(n11528), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14151), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11529) );
  NAND4_X1 U13111 ( .A1(n11532), .A2(n11531), .A3(n11530), .A4(n11529), .ZN(
        n11538) );
  AOI22_X1 U13112 ( .A1(n14152), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11559), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11536) );
  AOI22_X1 U13113 ( .A1(n11574), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14271), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11535) );
  AOI22_X1 U13114 ( .A1(n14287), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14253), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11534) );
  INV_X2 U13115 ( .A(n14285), .ZN(n14254) );
  AOI22_X1 U13116 ( .A1(n14270), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11533) );
  NAND4_X1 U13117 ( .A1(n11536), .A2(n11535), .A3(n11534), .A4(n11533), .ZN(
        n11537) );
  AOI22_X1 U13118 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n14210), .B1(
        n14288), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11541) );
  NAND2_X1 U13119 ( .A1(n14287), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11540) );
  NAND2_X1 U13120 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11539) );
  NAND3_X1 U13121 ( .A1(n11541), .A2(n11540), .A3(n11539), .ZN(n11545) );
  INV_X1 U13122 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11543) );
  NAND2_X1 U13123 ( .A1(n14253), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11542) );
  OAI21_X1 U13124 ( .B1(n14285), .B2(n11543), .A(n11542), .ZN(n11544) );
  NOR2_X1 U13125 ( .A1(n11545), .A2(n11544), .ZN(n11557) );
  NAND2_X1 U13126 ( .A1(n14269), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11549) );
  NAND2_X1 U13127 ( .A1(n14270), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11548) );
  NAND2_X1 U13128 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11547) );
  AOI22_X1 U13129 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n14273), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11546) );
  AND4_X1 U13130 ( .A1(n11549), .A2(n11548), .A3(n11547), .A4(n11546), .ZN(
        n11556) );
  NAND2_X1 U13131 ( .A1(n11528), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11553) );
  NAND2_X1 U13132 ( .A1(n14150), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11552) );
  NAND2_X1 U13133 ( .A1(n14151), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11551) );
  NAND2_X1 U13134 ( .A1(n14152), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11550) );
  AND4_X1 U13135 ( .A1(n11553), .A2(n11552), .A3(n11551), .A4(n11550), .ZN(
        n11555) );
  NAND2_X1 U13136 ( .A1(n11574), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11554) );
  NAND4_X1 U13137 ( .A1(n11557), .A2(n11556), .A3(n11555), .A4(n11554), .ZN(
        n12176) );
  AND2_X1 U13138 ( .A1(n11974), .A2(n12176), .ZN(n11558) );
  NAND2_X1 U13139 ( .A1(n11527), .A2(n11558), .ZN(n11586) );
  AOI22_X1 U13140 ( .A1(n14269), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14271), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11563) );
  AOI22_X1 U13141 ( .A1(n14254), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14270), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11562) );
  AOI22_X1 U13142 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11528), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11561) );
  AOI22_X1 U13143 ( .A1(n14152), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14150), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11560) );
  NAND4_X1 U13144 ( .A1(n11563), .A2(n11562), .A3(n11561), .A4(n11560), .ZN(
        n11572) );
  NAND2_X1 U13145 ( .A1(n14151), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11570) );
  AOI22_X1 U13146 ( .A1(n14210), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n14288), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11564) );
  INV_X1 U13147 ( .A(n11564), .ZN(n11568) );
  NAND2_X1 U13148 ( .A1(n14272), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11566) );
  NAND2_X1 U13149 ( .A1(n11566), .A2(n11565), .ZN(n11567) );
  NOR2_X1 U13150 ( .A1(n11568), .A2(n11567), .ZN(n11569) );
  NAND2_X1 U13151 ( .A1(n11570), .A2(n11569), .ZN(n11571) );
  AOI22_X1 U13152 ( .A1(n14287), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14253), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11573) );
  INV_X1 U13153 ( .A(n11573), .ZN(n11575) );
  NOR2_X2 U13154 ( .A1(n11578), .A2(n11244), .ZN(n11581) );
  INV_X1 U13155 ( .A(n11581), .ZN(n11579) );
  NAND2_X1 U13156 ( .A1(n11580), .A2(n11579), .ZN(n11583) );
  AND2_X2 U13157 ( .A1(n11583), .A2(n11612), .ZN(n12203) );
  INV_X1 U13158 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n16028) );
  NAND2_X1 U13159 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17666), .ZN(
        n17665) );
  NOR2_X1 U13160 ( .A1(n11988), .A2(n17665), .ZN(n11585) );
  INV_X1 U13161 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14624) );
  NAND2_X1 U13162 ( .A1(n17662), .A2(n17666), .ZN(n11584) );
  XNOR2_X1 U13163 ( .A(n12176), .B(n11584), .ZN(n14623) );
  NOR2_X1 U13164 ( .A1(n14624), .A2(n14623), .ZN(n14622) );
  NOR2_X1 U13165 ( .A1(n11585), .A2(n14622), .ZN(n11587) );
  XOR2_X1 U13166 ( .A(n16028), .B(n11587), .Z(n16010) );
  XNOR2_X1 U13167 ( .A(n11586), .B(n11993), .ZN(n16011) );
  NAND2_X1 U13168 ( .A1(n16010), .A2(n16011), .ZN(n16009) );
  OR2_X1 U13169 ( .A1(n11587), .A2(n16028), .ZN(n11588) );
  NAND2_X1 U13170 ( .A1(n16009), .A2(n11588), .ZN(n11590) );
  XNOR2_X1 U13171 ( .A(n11590), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15521) );
  NAND2_X1 U13172 ( .A1(n11590), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11591) );
  AOI22_X1 U13173 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n14210), .B1(
        n14288), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11594) );
  NAND2_X1 U13174 ( .A1(n14287), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11593) );
  NAND2_X1 U13175 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11592) );
  NAND3_X1 U13176 ( .A1(n11594), .A2(n11593), .A3(n11592), .ZN(n11598) );
  INV_X1 U13177 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11596) );
  NAND2_X1 U13178 ( .A1(n14253), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11595) );
  OAI21_X1 U13179 ( .B1(n11596), .B2(n14285), .A(n11595), .ZN(n11597) );
  NOR2_X1 U13180 ( .A1(n11598), .A2(n11597), .ZN(n11610) );
  NAND2_X1 U13181 ( .A1(n14269), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11602) );
  NAND2_X1 U13182 ( .A1(n14270), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11601) );
  NAND2_X1 U13183 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11600) );
  AOI22_X1 U13184 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n14273), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11599) );
  AND4_X1 U13185 ( .A1(n11602), .A2(n11601), .A3(n11600), .A4(n11599), .ZN(
        n11609) );
  NAND2_X1 U13186 ( .A1(n11528), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11606) );
  NAND2_X1 U13187 ( .A1(n14150), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11605) );
  NAND2_X1 U13188 ( .A1(n14151), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11604) );
  NAND2_X1 U13189 ( .A1(n14152), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11603) );
  AND4_X1 U13190 ( .A1(n11606), .A2(n11605), .A3(n11604), .A4(n11603), .ZN(
        n11608) );
  NAND2_X1 U13191 ( .A1(n11574), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11607) );
  NAND4_X1 U13192 ( .A1(n11610), .A2(n11609), .A3(n11608), .A4(n11607), .ZN(
        n12006) );
  INV_X1 U13193 ( .A(n12006), .ZN(n11611) );
  NAND2_X1 U13194 ( .A1(n11612), .A2(n11611), .ZN(n11613) );
  NAND2_X1 U13195 ( .A1(n11663), .A2(n11613), .ZN(n11615) );
  INV_X1 U13196 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15770) );
  NAND2_X1 U13197 ( .A1(n15692), .A2(n15770), .ZN(n11618) );
  INV_X1 U13198 ( .A(n11614), .ZN(n11616) );
  NAND2_X1 U13199 ( .A1(n11616), .A2(n11615), .ZN(n11617) );
  AOI22_X1 U13200 ( .A1(n19439), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11619), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11623) );
  AOI22_X1 U13201 ( .A1(n11620), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11621), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11622) );
  AND2_X1 U13202 ( .A1(n11623), .A2(n11622), .ZN(n11642) );
  AOI22_X1 U13203 ( .A1(n11508), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n19550), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11626) );
  AOI22_X1 U13204 ( .A1(n19450), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11517), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11625) );
  AND2_X1 U13205 ( .A1(n11626), .A2(n11625), .ZN(n11641) );
  INV_X1 U13206 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14421) );
  INV_X1 U13207 ( .A(n11628), .ZN(n19400) );
  AOI22_X1 U13208 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19383), .B1(
        n19400), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11631) );
  INV_X1 U13209 ( .A(n11629), .ZN(n19468) );
  NAND2_X1 U13210 ( .A1(n19468), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11630) );
  OAI211_X1 U13211 ( .C1(n19494), .C2(n14421), .A(n11631), .B(n11630), .ZN(
        n11637) );
  INV_X1 U13212 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11635) );
  INV_X1 U13213 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11634) );
  OAI22_X1 U13214 ( .A1(n11635), .A2(n11632), .B1(n11633), .B2(n11634), .ZN(
        n11636) );
  NOR2_X1 U13215 ( .A1(n11637), .A2(n11636), .ZN(n11640) );
  AOI22_X1 U13216 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19395), .B1(
        n19417), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11639) );
  NAND4_X1 U13217 ( .A1(n11642), .A2(n11641), .A3(n11640), .A4(n11639), .ZN(
        n11660) );
  NAND2_X1 U13218 ( .A1(n14270), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11646) );
  NAND2_X1 U13219 ( .A1(n14269), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11645) );
  NAND2_X1 U13220 ( .A1(n14150), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11644) );
  AOI22_X1 U13221 ( .A1(n14210), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11643) );
  NAND4_X1 U13222 ( .A1(n11646), .A2(n11645), .A3(n11644), .A4(n11643), .ZN(
        n11652) );
  NAND2_X1 U13223 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11650) );
  NAND2_X1 U13224 ( .A1(n14278), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11649) );
  NAND2_X1 U13225 ( .A1(n14151), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11648) );
  NAND2_X1 U13226 ( .A1(n14152), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11647) );
  NAND4_X1 U13227 ( .A1(n11650), .A2(n11649), .A3(n11648), .A4(n11647), .ZN(
        n11651) );
  NOR2_X1 U13228 ( .A1(n11652), .A2(n11651), .ZN(n11658) );
  AOI22_X1 U13229 ( .A1(n14254), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14253), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11656) );
  AOI22_X1 U13230 ( .A1(n14288), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14273), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11655) );
  NAND2_X1 U13231 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11654) );
  NAND2_X1 U13232 ( .A1(n14287), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11653) );
  NAND2_X1 U13233 ( .A1(n14295), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11657) );
  NAND2_X1 U13234 ( .A1(n12011), .A2(n10959), .ZN(n11659) );
  INV_X1 U13235 ( .A(n11661), .ZN(n11662) );
  NAND2_X1 U13236 ( .A1(n11663), .A2(n11662), .ZN(n12232) );
  NAND2_X1 U13237 ( .A1(n12231), .A2(n12232), .ZN(n11705) );
  NAND2_X1 U13238 ( .A1(n11666), .A2(n11705), .ZN(n11665) );
  INV_X1 U13239 ( .A(n11666), .ZN(n11704) );
  AOI22_X1 U13240 ( .A1(n11620), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n19550), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11668) );
  AOI22_X1 U13241 ( .A1(n19450), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11621), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11667) );
  AND2_X1 U13242 ( .A1(n11668), .A2(n11667), .ZN(n11681) );
  INV_X1 U13243 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14442) );
  AOI22_X1 U13244 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19383), .B1(
        n19400), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11670) );
  INV_X1 U13245 ( .A(n19494), .ZN(n19497) );
  NAND2_X1 U13246 ( .A1(n19497), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n11669) );
  OAI211_X1 U13247 ( .C1(n11629), .C2(n14442), .A(n11670), .B(n11669), .ZN(
        n11672) );
  INV_X1 U13248 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14249) );
  INV_X1 U13249 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14258) );
  OAI22_X1 U13250 ( .A1(n14249), .A2(n11632), .B1(n11633), .B2(n14258), .ZN(
        n11671) );
  NOR2_X1 U13251 ( .A1(n11672), .A2(n11671), .ZN(n11680) );
  INV_X1 U13252 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14257) );
  INV_X1 U13253 ( .A(n19439), .ZN(n11674) );
  INV_X1 U13254 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11673) );
  OAI22_X1 U13255 ( .A1(n14257), .A2(n11674), .B1(n11624), .B2(n11673), .ZN(
        n11677) );
  INV_X1 U13256 ( .A(n11619), .ZN(n19525) );
  INV_X1 U13257 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14261) );
  NAND2_X1 U13258 ( .A1(n11517), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11675) );
  OAI21_X1 U13259 ( .B1(n19525), .B2(n14261), .A(n11675), .ZN(n11676) );
  NOR2_X1 U13260 ( .A1(n11677), .A2(n11676), .ZN(n11679) );
  AOI22_X1 U13261 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19395), .B1(
        n19417), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11678) );
  NAND4_X1 U13262 ( .A1(n11681), .A2(n11680), .A3(n11679), .A4(n11678), .ZN(
        n11699) );
  NAND2_X1 U13263 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11685) );
  NAND2_X1 U13264 ( .A1(n14269), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11684) );
  NAND2_X1 U13265 ( .A1(n14270), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n11683) );
  AOI22_X1 U13266 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n14210), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11682) );
  NAND4_X1 U13267 ( .A1(n11685), .A2(n11684), .A3(n11683), .A4(n11682), .ZN(
        n11691) );
  NAND2_X1 U13268 ( .A1(n14278), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11689) );
  NAND2_X1 U13269 ( .A1(n14150), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11688) );
  NAND2_X1 U13270 ( .A1(n14151), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11687) );
  NAND2_X1 U13271 ( .A1(n14152), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11686) );
  NAND4_X1 U13272 ( .A1(n11689), .A2(n11688), .A3(n11687), .A4(n11686), .ZN(
        n11690) );
  NOR2_X1 U13273 ( .A1(n11691), .A2(n11690), .ZN(n11697) );
  AOI22_X1 U13274 ( .A1(n14254), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14253), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U13275 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n14273), .B1(
        n14288), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11694) );
  NAND2_X1 U13276 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11693) );
  NAND2_X1 U13277 ( .A1(n14287), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11692) );
  NAND2_X1 U13278 ( .A1(n14295), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11696) );
  NAND2_X1 U13279 ( .A1(n12184), .A2(n10959), .ZN(n11698) );
  INV_X1 U13280 ( .A(n12169), .ZN(n11701) );
  OAI21_X1 U13281 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n11664), .A(
        n11701), .ZN(n11702) );
  INV_X1 U13282 ( .A(n11715), .ZN(n11706) );
  INV_X1 U13283 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15771) );
  MUX2_X1 U13284 ( .A(n11706), .B(n15771), .S(n11705), .Z(n11707) );
  OAI21_X1 U13285 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n11712), .A(
        n11707), .ZN(n11708) );
  NAND2_X1 U13286 ( .A1(n11710), .A2(n11711), .ZN(n11713) );
  NAND2_X1 U13287 ( .A1(n11713), .A2(n11712), .ZN(n11714) );
  NAND2_X2 U13288 ( .A1(n17259), .A2(n11714), .ZN(n17247) );
  AOI22_X1 U13289 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n14273), .B1(
        n14288), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11719) );
  NAND2_X1 U13290 ( .A1(n14287), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11718) );
  NAND2_X1 U13291 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11717) );
  NAND3_X1 U13292 ( .A1(n11719), .A2(n11718), .A3(n11717), .ZN(n11722) );
  INV_X1 U13293 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14098) );
  NAND2_X1 U13294 ( .A1(n14253), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11720) );
  OAI21_X1 U13295 ( .B1(n14285), .B2(n14098), .A(n11720), .ZN(n11721) );
  NOR2_X1 U13296 ( .A1(n11722), .A2(n11721), .ZN(n11734) );
  NAND2_X1 U13297 ( .A1(n14269), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11726) );
  NAND2_X1 U13298 ( .A1(n14270), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11725) );
  NAND2_X1 U13299 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11724) );
  AOI22_X1 U13300 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n14210), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11723) );
  NAND2_X1 U13301 ( .A1(n14278), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11730) );
  NAND2_X1 U13302 ( .A1(n14150), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11729) );
  NAND2_X1 U13303 ( .A1(n14151), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11728) );
  NAND2_X1 U13304 ( .A1(n14152), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11727) );
  NAND2_X1 U13305 ( .A1(n14295), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11731) );
  NAND4_X1 U13306 ( .A1(n11734), .A2(n11733), .A3(n11732), .A4(n11731), .ZN(
        n12190) );
  NAND2_X1 U13307 ( .A1(n11735), .A2(n12202), .ZN(n11736) );
  NAND2_X1 U13308 ( .A1(n11739), .A2(n11736), .ZN(n11737) );
  XNOR2_X1 U13309 ( .A(n11737), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17246) );
  INV_X1 U13310 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17252) );
  INV_X1 U13311 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17232) );
  AND2_X1 U13312 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17185) );
  NAND2_X1 U13313 ( .A1(n17185), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17141) );
  NAND3_X1 U13314 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11741) );
  NOR2_X1 U13315 ( .A1(n17141), .A2(n11741), .ZN(n17130) );
  AND3_X1 U13316 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11742) );
  AND2_X1 U13317 ( .A1(n17130), .A2(n11742), .ZN(n17067) );
  NAND2_X1 U13318 ( .A1(n17067), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17069) );
  INV_X1 U13319 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16877) );
  AND2_X1 U13320 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12164) );
  NAND2_X1 U13321 ( .A1(n16876), .A2(n12164), .ZN(n16840) );
  INV_X1 U13322 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12321) );
  NAND2_X1 U13323 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11743) );
  OR2_X1 U13324 ( .A1(n17069), .A2(n11743), .ZN(n11940) );
  NAND2_X1 U13325 ( .A1(n12164), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11744) );
  NOR2_X1 U13326 ( .A1(n11940), .A2(n11744), .ZN(n14506) );
  MUX2_X1 U13327 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n19523), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n11780) );
  INV_X1 U13328 ( .A(n11780), .ZN(n11746) );
  NAND2_X1 U13329 ( .A1(n19424), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11764) );
  NAND2_X1 U13330 ( .A1(n11746), .A2(n11758), .ZN(n11748) );
  NAND2_X1 U13331 ( .A1(n19523), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11747) );
  XNOR2_X1 U13332 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11756) );
  NAND2_X1 U13333 ( .A1(n11757), .A2(n11756), .ZN(n11750) );
  NAND2_X1 U13334 ( .A1(n19518), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11749) );
  MUX2_X1 U13335 ( .A(n14101), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11753) );
  NOR2_X1 U13336 ( .A1(n11374), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11751) );
  NOR2_X1 U13337 ( .A1(n17330), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11752) );
  NAND2_X1 U13338 ( .A1(n11760), .A2(n11752), .ZN(n11774) );
  INV_X1 U13339 ( .A(n11753), .ZN(n11754) );
  XNOR2_X1 U13340 ( .A(n11755), .B(n11754), .ZN(n11773) );
  XNOR2_X1 U13341 ( .A(n11757), .B(n11756), .ZN(n11786) );
  NOR2_X1 U13342 ( .A1(n11791), .A2(n11786), .ZN(n11765) );
  XNOR2_X1 U13343 ( .A(n11780), .B(n11758), .ZN(n11781) );
  NAND2_X1 U13344 ( .A1(n17330), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11759) );
  NAND2_X1 U13345 ( .A1(n11760), .A2(n11759), .ZN(n11762) );
  NAND2_X1 U13346 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18873), .ZN(
        n11761) );
  NAND2_X1 U13347 ( .A1(n11418), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11763) );
  NAND2_X1 U13348 ( .A1(n11764), .A2(n11763), .ZN(n11779) );
  INV_X1 U13349 ( .A(n11779), .ZN(n11782) );
  NAND2_X1 U13350 ( .A1(n11765), .A2(n11782), .ZN(n11766) );
  NAND2_X1 U13351 ( .A1(n15319), .A2(n11766), .ZN(n11767) );
  NAND2_X1 U13352 ( .A1(n11767), .A2(n17326), .ZN(n11771) );
  AND2_X1 U13353 ( .A1(n18873), .A2(n11768), .ZN(n18869) );
  INV_X1 U13354 ( .A(n18869), .ZN(n11770) );
  NOR2_X1 U13355 ( .A1(n17326), .A2(P2_FLUSH_REG_SCAN_IN), .ZN(n11769) );
  OAI21_X1 U13356 ( .B1(n14269), .B2(n11770), .A(n11769), .ZN(n17675) );
  NAND2_X1 U13357 ( .A1(n11771), .A2(n17675), .ZN(n18901) );
  MUX2_X1 U13358 ( .A(n17666), .B(n11779), .S(n15313), .Z(n12207) );
  INV_X1 U13359 ( .A(n11786), .ZN(n11772) );
  OAI21_X1 U13360 ( .B1(n12207), .B2(n11780), .A(n12171), .ZN(n11775) );
  MUX2_X1 U13361 ( .A(n11774), .B(n12006), .S(n11394), .Z(n12180) );
  NAND3_X1 U13362 ( .A1(n11775), .A2(n12177), .A3(n12180), .ZN(n11777) );
  INV_X1 U13363 ( .A(n11795), .ZN(n11776) );
  AND2_X1 U13364 ( .A1(n10959), .A2(n14636), .ZN(n12435) );
  NAND2_X1 U13365 ( .A1(n15316), .A2(n12435), .ZN(n13743) );
  OAI21_X1 U13366 ( .B1(n10959), .B2(n18901), .A(n13743), .ZN(n11778) );
  INV_X1 U13367 ( .A(n13741), .ZN(n15317) );
  NAND2_X1 U13368 ( .A1(n11778), .A2(n15317), .ZN(n11822) );
  OAI21_X1 U13369 ( .B1(n11780), .B2(n11779), .A(n11394), .ZN(n11784) );
  OAI211_X1 U13370 ( .C1(n11969), .C2(n11782), .A(n11411), .B(n11781), .ZN(
        n11783) );
  OAI211_X1 U13371 ( .C1(n11785), .C2(n11786), .A(n11784), .B(n11783), .ZN(
        n11790) );
  OAI21_X1 U13372 ( .B1(n11527), .B2(n14636), .A(n11786), .ZN(n11787) );
  NAND2_X1 U13373 ( .A1(n11787), .A2(n12171), .ZN(n11788) );
  NAND3_X1 U13374 ( .A1(n11790), .A2(n11789), .A3(n11788), .ZN(n11793) );
  AOI21_X1 U13375 ( .B1(n11394), .B2(n11791), .A(n11795), .ZN(n11792) );
  NAND2_X1 U13376 ( .A1(n11793), .A2(n11792), .ZN(n11794) );
  MUX2_X1 U13377 ( .A(n11794), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n11407), .Z(n11799) );
  NAND3_X1 U13378 ( .A1(n11795), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n14636), 
        .ZN(n11796) );
  NAND2_X1 U13379 ( .A1(n15781), .A2(n11969), .ZN(n14634) );
  INV_X1 U13380 ( .A(n14634), .ZN(n15262) );
  NAND2_X1 U13381 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n18908) );
  INV_X1 U13382 ( .A(n18908), .ZN(n21850) );
  INV_X2 U13383 ( .A(n17770), .ZN(n21855) );
  INV_X1 U13384 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n21851) );
  NAND2_X2 U13385 ( .A1(n21855), .A2(n21851), .ZN(n17765) );
  NOR2_X1 U13386 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_0__SCAN_IN), 
        .ZN(n21852) );
  NAND2_X1 U13387 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n21852), .ZN(n17740) );
  NAND2_X1 U13388 ( .A1(n17765), .A2(n17740), .ZN(n21857) );
  INV_X1 U13389 ( .A(n21857), .ZN(n11797) );
  NOR2_X1 U13390 ( .A1(n21850), .A2(n11797), .ZN(n15326) );
  NAND3_X1 U13391 ( .A1(n15262), .A2(n15326), .A3(n11798), .ZN(n11820) );
  AOI21_X1 U13392 ( .B1(n11799), .B2(n11411), .A(n19674), .ZN(n11818) );
  NAND3_X1 U13393 ( .A1(n15319), .A2(n15340), .A3(n15326), .ZN(n11814) );
  NAND2_X1 U13394 ( .A1(n11801), .A2(n11800), .ZN(n11802) );
  NAND2_X1 U13395 ( .A1(n11802), .A2(n14715), .ZN(n11803) );
  NAND2_X1 U13396 ( .A1(n11803), .A2(n12435), .ZN(n11920) );
  AOI21_X1 U13397 ( .B1(n10959), .B2(n11804), .A(n14636), .ZN(n11805) );
  OAI21_X1 U13398 ( .B1(n11805), .B2(n19380), .A(n19753), .ZN(n11806) );
  AND4_X1 U13399 ( .A1(n11920), .A2(n11808), .A3(n11807), .A4(n11806), .ZN(
        n11813) );
  NAND2_X1 U13400 ( .A1(n11810), .A2(n19753), .ZN(n11811) );
  NAND2_X1 U13401 ( .A1(n18870), .A2(n11811), .ZN(n11812) );
  AND3_X1 U13402 ( .A1(n11814), .A2(n11813), .A3(n11812), .ZN(n15259) );
  MUX2_X1 U13403 ( .A(n15340), .B(n11798), .S(n10959), .Z(n11815) );
  NAND3_X1 U13404 ( .A1(n11815), .A2(n15319), .A3(n18908), .ZN(n11816) );
  NAND2_X1 U13405 ( .A1(n15259), .A2(n11816), .ZN(n11817) );
  AOI21_X1 U13406 ( .B1(n14634), .B2(n11818), .A(n11817), .ZN(n11819) );
  AND2_X1 U13407 ( .A1(n11820), .A2(n11819), .ZN(n11821) );
  NAND2_X1 U13408 ( .A1(n11822), .A2(n11821), .ZN(n11823) );
  INV_X1 U13409 ( .A(n12435), .ZN(n15315) );
  NOR2_X1 U13410 ( .A1(n13741), .A2(n15315), .ZN(n11824) );
  NAND2_X1 U13411 ( .A1(n11826), .A2(n11825), .ZN(n11831) );
  INV_X1 U13412 ( .A(n11827), .ZN(n11829) );
  NAND2_X1 U13413 ( .A1(n11829), .A2(n11828), .ZN(n11830) );
  NAND2_X1 U13414 ( .A1(n11831), .A2(n11830), .ZN(n14952) );
  INV_X1 U13415 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n12179) );
  NAND2_X1 U13416 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11835) );
  NAND2_X1 U13417 ( .A1(n13678), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11834) );
  OAI211_X1 U13418 ( .C1(n11833), .C2(n12179), .A(n11835), .B(n11834), .ZN(
        n11836) );
  AOI21_X1 U13419 ( .B1(n12398), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n11836), .ZN(n14951) );
  NOR2_X2 U13420 ( .A1(n14952), .A2(n14951), .ZN(n14972) );
  NAND2_X1 U13421 ( .A1(n12398), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11841) );
  INV_X1 U13422 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n14974) );
  NAND2_X1 U13423 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11838) );
  NAND2_X1 U13424 ( .A1(n12390), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11837) );
  OAI211_X1 U13425 ( .C1(n11833), .C2(n14974), .A(n11838), .B(n11837), .ZN(
        n11839) );
  INV_X1 U13426 ( .A(n11839), .ZN(n11840) );
  NAND2_X1 U13427 ( .A1(n11841), .A2(n11840), .ZN(n14973) );
  NAND2_X1 U13428 ( .A1(n14972), .A2(n14973), .ZN(n14971) );
  INV_X1 U13429 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n11844) );
  NAND2_X1 U13430 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11843) );
  NAND2_X1 U13431 ( .A1(n13678), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11842) );
  OAI211_X1 U13432 ( .C1(n11833), .C2(n11844), .A(n11843), .B(n11842), .ZN(
        n11845) );
  AOI21_X1 U13433 ( .B1(n12398), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n11845), .ZN(n15073) );
  INV_X1 U13434 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n12189) );
  NAND2_X1 U13435 ( .A1(n12398), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11847) );
  AOI22_X1 U13436 ( .A1(n13678), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11846) );
  OAI211_X1 U13437 ( .C1(n11833), .C2(n12189), .A(n11847), .B(n11846), .ZN(
        n15152) );
  NAND2_X1 U13438 ( .A1(n15074), .A2(n15152), .ZN(n14962) );
  INV_X1 U13439 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n11850) );
  NAND2_X1 U13440 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11849) );
  NAND2_X1 U13441 ( .A1(n13678), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11848) );
  OAI211_X1 U13442 ( .C1(n11833), .C2(n11850), .A(n11849), .B(n11848), .ZN(
        n11851) );
  AOI21_X1 U13443 ( .B1(n12398), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n11851), .ZN(n14963) );
  INV_X1 U13444 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n11854) );
  NAND2_X1 U13445 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11853) );
  NAND2_X1 U13446 ( .A1(n12390), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11852) );
  OAI211_X1 U13447 ( .C1(n11833), .C2(n11854), .A(n11853), .B(n11852), .ZN(
        n11855) );
  AOI21_X1 U13448 ( .B1(n12398), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n11855), .ZN(n14958) );
  INV_X1 U13449 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n11858) );
  NAND2_X1 U13450 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11857) );
  NAND2_X1 U13451 ( .A1(n12390), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11856) );
  OAI211_X1 U13452 ( .C1(n11833), .C2(n11858), .A(n11857), .B(n11856), .ZN(
        n11859) );
  AOI21_X1 U13453 ( .B1(n12398), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n11859), .ZN(n15189) );
  INV_X1 U13454 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n11862) );
  NAND2_X1 U13455 ( .A1(n12398), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11861) );
  AOI22_X1 U13456 ( .A1(n13678), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11860) );
  OAI211_X1 U13457 ( .C1(n11833), .C2(n11862), .A(n11861), .B(n11860), .ZN(
        n14571) );
  NAND2_X1 U13458 ( .A1(n15187), .A2(n14571), .ZN(n14570) );
  INV_X1 U13459 ( .A(n14570), .ZN(n11868) );
  INV_X1 U13460 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n11865) );
  NAND2_X1 U13461 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11864) );
  NAND2_X1 U13462 ( .A1(n12390), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11863) );
  OAI211_X1 U13463 ( .C1(n11833), .C2(n11865), .A(n11864), .B(n11863), .ZN(
        n11866) );
  AOI21_X1 U13464 ( .B1(n12398), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n11866), .ZN(n15394) );
  INV_X1 U13465 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n11871) );
  NAND2_X1 U13466 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11870) );
  NAND2_X1 U13467 ( .A1(n12390), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11869) );
  OAI211_X1 U13468 ( .C1(n11833), .C2(n11871), .A(n11870), .B(n11869), .ZN(
        n11872) );
  AOI21_X1 U13469 ( .B1(n12398), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n11872), .ZN(n15484) );
  INV_X1 U13470 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n11875) );
  NAND2_X1 U13471 ( .A1(n12398), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11874) );
  AOI22_X1 U13472 ( .A1(n13678), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11873) );
  OAI211_X1 U13473 ( .C1(n11833), .C2(n11875), .A(n11874), .B(n11873), .ZN(
        n15456) );
  INV_X1 U13474 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n11878) );
  NAND2_X1 U13475 ( .A1(n12398), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11877) );
  AOI22_X1 U13476 ( .A1(n13678), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11876) );
  OAI211_X1 U13477 ( .C1(n11833), .C2(n11878), .A(n11877), .B(n11876), .ZN(
        n15579) );
  INV_X1 U13478 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n11881) );
  NAND2_X1 U13479 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11880) );
  NAND2_X1 U13480 ( .A1(n12390), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11879) );
  OAI211_X1 U13481 ( .C1(n11833), .C2(n11881), .A(n11880), .B(n11879), .ZN(
        n11882) );
  AOI21_X1 U13482 ( .B1(n12398), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n11882), .ZN(n15634) );
  INV_X1 U13483 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n11885) );
  NAND2_X1 U13484 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11884) );
  NAND2_X1 U13485 ( .A1(n12390), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11883) );
  OAI211_X1 U13486 ( .C1(n11833), .C2(n11885), .A(n11884), .B(n11883), .ZN(
        n11886) );
  AOI21_X1 U13487 ( .B1(n12398), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n11886), .ZN(n15707) );
  INV_X1 U13488 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n11889) );
  NAND2_X1 U13489 ( .A1(n12398), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11888) );
  AOI22_X1 U13490 ( .A1(n13678), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11887) );
  OAI211_X1 U13491 ( .C1(n11833), .C2(n11889), .A(n11888), .B(n11887), .ZN(
        n15798) );
  NAND2_X1 U13492 ( .A1(n15799), .A2(n15798), .ZN(n15797) );
  INV_X1 U13493 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n11892) );
  NAND2_X1 U13494 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11891) );
  NAND2_X1 U13495 ( .A1(n12390), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11890) );
  OAI211_X1 U13496 ( .C1(n11833), .C2(n11892), .A(n11891), .B(n11890), .ZN(
        n11893) );
  AOI21_X1 U13497 ( .B1(n12398), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n11893), .ZN(n15880) );
  INV_X1 U13498 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n11896) );
  NAND2_X1 U13499 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11895) );
  NAND2_X1 U13500 ( .A1(n12390), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11894) );
  OAI211_X1 U13501 ( .C1(n11833), .C2(n11896), .A(n11895), .B(n11894), .ZN(
        n11897) );
  AOI21_X1 U13502 ( .B1(n12398), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11897), .ZN(n15958) );
  INV_X1 U13503 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n11901) );
  NAND2_X1 U13504 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11900) );
  NAND2_X1 U13505 ( .A1(n12390), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11899) );
  OAI211_X1 U13506 ( .C1(n11833), .C2(n11901), .A(n11900), .B(n11899), .ZN(
        n11902) );
  AOI21_X1 U13507 ( .B1(n12398), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n11902), .ZN(n16692) );
  INV_X1 U13508 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n16624) );
  NAND2_X1 U13509 ( .A1(n12398), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11904) );
  AOI22_X1 U13510 ( .A1(n13678), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11903) );
  OAI211_X1 U13511 ( .C1(n11833), .C2(n16624), .A(n11904), .B(n11903), .ZN(
        n16617) );
  INV_X1 U13512 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n11907) );
  NAND2_X1 U13513 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n11906) );
  NAND2_X1 U13514 ( .A1(n12390), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11905) );
  OAI211_X1 U13515 ( .C1(n11833), .C2(n11907), .A(n11906), .B(n11905), .ZN(
        n11908) );
  AOI21_X1 U13516 ( .B1(n12398), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n11908), .ZN(n11910) );
  OR2_X2 U13517 ( .A1(n11909), .A2(n11910), .ZN(n16671) );
  NAND2_X1 U13518 ( .A1(n11909), .A2(n11910), .ZN(n11911) );
  NAND2_X1 U13519 ( .A1(n16671), .A2(n11911), .ZN(n18792) );
  INV_X1 U13520 ( .A(n11947), .ZN(n12325) );
  NAND2_X1 U13521 ( .A1(n15786), .A2(n10959), .ZN(n11914) );
  AND2_X1 U13522 ( .A1(n11912), .A2(n11914), .ZN(n11915) );
  NAND3_X1 U13523 ( .A1(n19753), .A2(n10959), .A3(n12181), .ZN(n11917) );
  NOR2_X1 U13524 ( .A1(n15280), .A2(n11917), .ZN(n15312) );
  NAND2_X1 U13525 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n16024) );
  NAND2_X1 U13526 ( .A1(n16028), .A2(n16024), .ZN(n16021) );
  INV_X1 U13527 ( .A(n16021), .ZN(n11918) );
  NAND2_X1 U13528 ( .A1(n17103), .A2(n11918), .ZN(n11937) );
  NAND2_X1 U13529 ( .A1(n11919), .A2(n11969), .ZN(n15279) );
  AOI21_X1 U13530 ( .B1(n15279), .B2(n11920), .A(n11377), .ZN(n11929) );
  OAI21_X1 U13531 ( .B1(n11925), .B2(n11922), .A(n11921), .ZN(n11924) );
  NAND2_X1 U13532 ( .A1(n11924), .A2(n11923), .ZN(n11927) );
  NAND2_X1 U13533 ( .A1(n11926), .A2(n11925), .ZN(n14714) );
  OAI211_X1 U13534 ( .C1(n19674), .C2(n11921), .A(n11927), .B(n14714), .ZN(
        n11928) );
  OR2_X1 U13535 ( .A1(n11929), .A2(n11928), .ZN(n11933) );
  INV_X1 U13536 ( .A(n11930), .ZN(n11931) );
  MUX2_X1 U13537 ( .A(n11931), .B(n11798), .S(n14636), .Z(n11932) );
  NOR2_X1 U13538 ( .A1(n11933), .A2(n11932), .ZN(n15281) );
  INV_X1 U13539 ( .A(n11934), .ZN(n15268) );
  NAND2_X1 U13540 ( .A1(n15281), .A2(n15268), .ZN(n11935) );
  INV_X1 U13541 ( .A(n17104), .ZN(n11936) );
  NOR2_X1 U13542 ( .A1(n16028), .A2(n16024), .ZN(n16019) );
  NOR2_X1 U13543 ( .A1(n11936), .A2(n16019), .ZN(n16026) );
  OR2_X1 U13544 ( .A1(n19549), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n17602) );
  NOR2_X1 U13545 ( .A1(n17602), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12161) );
  INV_X1 U13546 ( .A(n12161), .ZN(n18746) );
  INV_X1 U13547 ( .A(n18746), .ZN(n16976) );
  NOR2_X1 U13548 ( .A1(n11947), .A2(n16976), .ZN(n18877) );
  NOR2_X1 U13549 ( .A1(n16026), .A2(n18877), .ZN(n14503) );
  INV_X1 U13550 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17268) );
  NAND3_X1 U13551 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17263) );
  NOR2_X1 U13552 ( .A1(n17268), .A2(n17263), .ZN(n17228) );
  NOR2_X1 U13553 ( .A1(n17252), .A2(n17232), .ZN(n17231) );
  NAND2_X1 U13554 ( .A1(n17228), .A2(n17231), .ZN(n14504) );
  NAND2_X1 U13555 ( .A1(n17262), .A2(n14504), .ZN(n11938) );
  NAND2_X1 U13556 ( .A1(n17262), .A2(n11940), .ZN(n11939) );
  NAND2_X1 U13557 ( .A1(n17222), .A2(n11939), .ZN(n17058) );
  INV_X1 U13558 ( .A(n11940), .ZN(n11942) );
  AND2_X1 U13559 ( .A1(n17103), .A2(n16021), .ZN(n15515) );
  AND2_X1 U13560 ( .A1(n17104), .A2(n16019), .ZN(n11941) );
  NOR2_X1 U13561 ( .A1(n15515), .A2(n11941), .ZN(n15698) );
  NOR2_X1 U13562 ( .A1(n15698), .A2(n17263), .ZN(n17266) );
  NAND2_X1 U13563 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17266), .ZN(
        n17230) );
  INV_X1 U13564 ( .A(n17230), .ZN(n17251) );
  NAND2_X1 U13565 ( .A1(n11942), .A2(n17218), .ZN(n17044) );
  NOR2_X1 U13566 ( .A1(n17044), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n17055) );
  OR2_X1 U13567 ( .A1(n17058), .A2(n17055), .ZN(n17047) );
  AND2_X1 U13568 ( .A1(n11943), .A2(n11969), .ZN(n11945) );
  NOR2_X1 U13569 ( .A1(n11944), .A2(n15280), .ZN(n15321) );
  OR2_X1 U13570 ( .A1(n11945), .A2(n15321), .ZN(n11946) );
  NAND2_X1 U13571 ( .A1(n14269), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11951) );
  NAND2_X1 U13572 ( .A1(n14278), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11950) );
  NAND2_X1 U13573 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11949) );
  AOI22_X1 U13574 ( .A1(n14210), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11948) );
  AND4_X1 U13575 ( .A1(n11951), .A2(n11950), .A3(n11949), .A4(n11948), .ZN(
        n11966) );
  NAND2_X1 U13576 ( .A1(n14270), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11955) );
  NAND2_X1 U13577 ( .A1(n14150), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11954) );
  NAND2_X1 U13578 ( .A1(n14151), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11953) );
  NAND2_X1 U13579 ( .A1(n14152), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11952) );
  AND4_X1 U13580 ( .A1(n11955), .A2(n11954), .A3(n11953), .A4(n11952), .ZN(
        n11965) );
  INV_X1 U13581 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11956) );
  INV_X1 U13582 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14154) );
  OAI22_X1 U13583 ( .A1(n14285), .A2(n11956), .B1(n15306), .B2(n14154), .ZN(
        n11962) );
  NAND2_X1 U13584 ( .A1(n14253), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11960) );
  NAND2_X1 U13585 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11959) );
  NAND2_X1 U13586 ( .A1(n14273), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11958) );
  NAND2_X1 U13587 ( .A1(n14288), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11957) );
  NAND4_X1 U13588 ( .A1(n11960), .A2(n11959), .A3(n11958), .A4(n11957), .ZN(
        n11961) );
  NOR2_X1 U13589 ( .A1(n11962), .A2(n11961), .ZN(n11964) );
  NAND2_X1 U13590 ( .A1(n14295), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11963) );
  NAND4_X1 U13591 ( .A1(n11966), .A2(n11965), .A3(n11964), .A4(n11963), .ZN(
        n14967) );
  INV_X1 U13592 ( .A(n14967), .ZN(n11972) );
  INV_X1 U13593 ( .A(n11967), .ZN(n15644) );
  AND2_X2 U13594 ( .A1(n15644), .A2(n12010), .ZN(n12021) );
  NAND2_X1 U13595 ( .A1(n12021), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11971) );
  NOR2_X1 U13596 ( .A1(n14715), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11968) );
  AOI22_X1 U13597 ( .A1(n13660), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n11015), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11970) );
  OAI211_X1 U13598 ( .C1(n11972), .C2(n11008), .A(n11971), .B(n11970), .ZN(
        n14770) );
  NAND2_X1 U13599 ( .A1(n14719), .A2(n11983), .ZN(n11994) );
  OAI211_X1 U13600 ( .C1(n19424), .C2(n19459), .A(n11994), .B(n11982), .ZN(
        n11976) );
  NAND2_X1 U13601 ( .A1(n12021), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11981) );
  NAND2_X1 U13602 ( .A1(n11969), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11980) );
  INV_X1 U13603 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n11977) );
  NAND2_X1 U13604 ( .A1(n12021), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11985) );
  AOI22_X1 U13605 ( .A1(n11968), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n11015), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11984) );
  NOR2_X1 U13606 ( .A1(n14719), .A2(n19380), .ZN(n11987) );
  MUX2_X1 U13607 ( .A(n11987), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_STATE2_REG_3__SCAN_IN), .Z(n11990) );
  INV_X1 U13608 ( .A(n12176), .ZN(n11988) );
  NOR2_X1 U13609 ( .A1(n11008), .A2(n11988), .ZN(n11989) );
  NOR2_X1 U13610 ( .A1(n11990), .A2(n11989), .ZN(n14721) );
  NAND2_X1 U13611 ( .A1(n11991), .A2(n14734), .ZN(n11992) );
  OR2_X1 U13612 ( .A1(n11008), .A2(n11993), .ZN(n11995) );
  OAI211_X1 U13613 ( .C1(n19459), .C2(n19518), .A(n11995), .B(n11994), .ZN(
        n11998) );
  XNOR2_X1 U13614 ( .A(n11999), .B(n11998), .ZN(n15362) );
  NAND2_X1 U13615 ( .A1(n12021), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11997) );
  AOI22_X1 U13616 ( .A1(n13660), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n11015), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11996) );
  AND2_X1 U13617 ( .A1(n11997), .A2(n11996), .ZN(n15361) );
  INV_X1 U13618 ( .A(n11998), .ZN(n12000) );
  NAND2_X1 U13619 ( .A1(n12000), .A2(n11999), .ZN(n12001) );
  INV_X1 U13620 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n15699) );
  OAI22_X1 U13621 ( .A1(n12009), .A2(n15699), .B1(n14101), .B2(n19459), .ZN(
        n12005) );
  INV_X1 U13622 ( .A(n12021), .ZN(n12429) );
  INV_X1 U13623 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n17744) );
  INV_X1 U13624 ( .A(n12002), .ZN(n12003) );
  OAI22_X1 U13625 ( .A1(n12429), .A2(n17744), .B1(n12003), .B2(n11008), .ZN(
        n12004) );
  AOI211_X1 U13626 ( .C1(n13660), .C2(P2_EAX_REG_3__SCAN_IN), .A(n12005), .B(
        n12004), .ZN(n15471) );
  AOI22_X1 U13627 ( .A1(n12021), .A2(P2_REIP_REG_4__SCAN_IN), .B1(n11015), 
        .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12008) );
  AOI22_X1 U13628 ( .A1(n11007), .A2(n12006), .B1(n13660), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n12007) );
  NAND2_X1 U13629 ( .A1(n12008), .A2(n12007), .ZN(n15499) );
  NAND2_X1 U13630 ( .A1(n12418), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n12017) );
  NAND2_X1 U13631 ( .A1(n11015), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12016) );
  INV_X1 U13632 ( .A(n12010), .ZN(n12013) );
  INV_X1 U13633 ( .A(n12011), .ZN(n12012) );
  NAND2_X1 U13634 ( .A1(n12181), .A2(n12012), .ZN(n12183) );
  OR2_X1 U13635 ( .A1(n12013), .A2(n12183), .ZN(n12015) );
  NAND2_X1 U13636 ( .A1(n13660), .A2(P2_EAX_REG_5__SCAN_IN), .ZN(n12014) );
  NOR2_X2 U13637 ( .A1(n15497), .A2(n15498), .ZN(n15496) );
  INV_X1 U13638 ( .A(n12184), .ZN(n12018) );
  NOR2_X1 U13639 ( .A1(n15496), .A2(n12019), .ZN(n14717) );
  AOI222_X1 U13640 ( .A1(n12021), .A2(P2_REIP_REG_6__SCAN_IN), .B1(n13660), 
        .B2(P2_EAX_REG_6__SCAN_IN), .C1(n11015), .C2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14718) );
  NOR2_X2 U13641 ( .A1(n14717), .A2(n14718), .ZN(n14716) );
  INV_X1 U13642 ( .A(n12190), .ZN(n12202) );
  NOR2_X1 U13643 ( .A1(n14716), .A2(n12020), .ZN(n14766) );
  NAND2_X1 U13644 ( .A1(n12021), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n12023) );
  AOI22_X1 U13645 ( .A1(n13660), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n11015), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12022) );
  NOR2_X2 U13646 ( .A1(n14766), .A2(n14767), .ZN(n14771) );
  AOI22_X1 U13647 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n14270), .B1(
        n14269), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12027) );
  AOI22_X1 U13648 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n14278), .B1(
        n14150), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12026) );
  AOI22_X1 U13649 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n14152), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12025) );
  AOI22_X1 U13650 ( .A1(n14151), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12024) );
  NAND4_X1 U13651 ( .A1(n12027), .A2(n12026), .A3(n12025), .A4(n12024), .ZN(
        n12033) );
  AOI22_X1 U13652 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n14287), .B1(
        n14253), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12031) );
  AOI22_X1 U13653 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12030) );
  AOI22_X1 U13654 ( .A1(n14288), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n14295), .ZN(n12029) );
  AOI22_X1 U13655 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n14210), .B1(
        n14273), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12028) );
  NAND4_X1 U13656 ( .A1(n12031), .A2(n12030), .A3(n12029), .A4(n12028), .ZN(
        n12032) );
  NOR2_X1 U13657 ( .A1(n12033), .A2(n12032), .ZN(n14956) );
  NAND2_X1 U13658 ( .A1(n12021), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12035) );
  AOI22_X1 U13659 ( .A1(n13660), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n11015), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12034) );
  OAI211_X1 U13660 ( .C1(n14956), .C2(n11008), .A(n12035), .B(n12034), .ZN(
        n15755) );
  NAND2_X1 U13661 ( .A1(n12418), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n12057) );
  AOI22_X1 U13662 ( .A1(n13660), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n11015), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12056) );
  NAND2_X1 U13663 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n12039) );
  NAND2_X1 U13664 ( .A1(n14278), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n12038) );
  NAND2_X1 U13665 ( .A1(n14269), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n12037) );
  AOI22_X1 U13666 ( .A1(n14210), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12036) );
  AND4_X1 U13667 ( .A1(n12039), .A2(n12038), .A3(n12037), .A4(n12036), .ZN(
        n12054) );
  NAND2_X1 U13668 ( .A1(n14270), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n12043) );
  NAND2_X1 U13669 ( .A1(n14150), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n12042) );
  NAND2_X1 U13670 ( .A1(n14151), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n12041) );
  NAND2_X1 U13671 ( .A1(n14152), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12040) );
  AND4_X1 U13672 ( .A1(n12043), .A2(n12042), .A3(n12041), .A4(n12040), .ZN(
        n12053) );
  INV_X1 U13673 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12044) );
  INV_X1 U13674 ( .A(n14253), .ZN(n14284) );
  INV_X1 U13675 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14358) );
  OAI22_X1 U13676 ( .A1(n14285), .A2(n12044), .B1(n14284), .B2(n14358), .ZN(
        n12050) );
  NAND2_X1 U13677 ( .A1(n14287), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12048) );
  NAND2_X1 U13678 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12047) );
  NAND2_X1 U13679 ( .A1(n14273), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n12046) );
  NAND2_X1 U13680 ( .A1(n14288), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n12045) );
  NAND4_X1 U13681 ( .A1(n12048), .A2(n12047), .A3(n12046), .A4(n12045), .ZN(
        n12049) );
  NOR2_X1 U13682 ( .A1(n12050), .A2(n12049), .ZN(n12052) );
  NAND2_X1 U13683 ( .A1(n14295), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12051) );
  NAND4_X1 U13684 ( .A1(n12054), .A2(n12053), .A3(n12052), .A4(n12051), .ZN(
        n15192) );
  OR2_X1 U13685 ( .A1(n11008), .A2(n14134), .ZN(n12055) );
  NAND2_X1 U13686 ( .A1(n12418), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n12071) );
  AOI22_X1 U13687 ( .A1(n13660), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n11015), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12070) );
  AOI22_X1 U13688 ( .A1(n14269), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14270), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12061) );
  AOI22_X1 U13689 ( .A1(n14278), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14150), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12060) );
  AOI22_X1 U13690 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14152), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12059) );
  AOI22_X1 U13691 ( .A1(n14151), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12058) );
  NAND4_X1 U13692 ( .A1(n12061), .A2(n12060), .A3(n12059), .A4(n12058), .ZN(
        n12068) );
  AOI22_X1 U13693 ( .A1(n14253), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14287), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12066) );
  AOI22_X1 U13694 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12065) );
  NOR2_X1 U13695 ( .A1(n14107), .A2(n12099), .ZN(n12062) );
  AOI21_X1 U13696 ( .B1(n14288), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n12062), .ZN(n12064) );
  AOI22_X1 U13697 ( .A1(n14210), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14273), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12063) );
  NAND4_X1 U13698 ( .A1(n12066), .A2(n12065), .A3(n12064), .A4(n12063), .ZN(
        n12067) );
  NAND2_X1 U13699 ( .A1(n11007), .A2(n15184), .ZN(n12069) );
  NAND2_X1 U13700 ( .A1(n14270), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n12075) );
  NAND2_X1 U13701 ( .A1(n14269), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12074) );
  NAND2_X1 U13702 ( .A1(n14150), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12073) );
  AOI22_X1 U13703 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n14272), .B1(
        n14273), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12072) );
  AND4_X1 U13704 ( .A1(n12075), .A2(n12074), .A3(n12073), .A4(n12072), .ZN(
        n12091) );
  NAND2_X1 U13705 ( .A1(n14151), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n12079) );
  NAND2_X1 U13706 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12078) );
  NAND2_X1 U13707 ( .A1(n11528), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12077) );
  NAND2_X1 U13708 ( .A1(n14152), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12076) );
  AND4_X1 U13709 ( .A1(n12079), .A2(n12078), .A3(n12077), .A4(n12076), .ZN(
        n12090) );
  INV_X1 U13710 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12081) );
  INV_X1 U13711 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12080) );
  OAI22_X1 U13712 ( .A1(n12081), .A2(n14285), .B1(n15306), .B2(n12080), .ZN(
        n12087) );
  NAND2_X1 U13713 ( .A1(n14253), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n12085) );
  NAND2_X1 U13714 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12084) );
  NAND2_X1 U13715 ( .A1(n14288), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12083) );
  NAND2_X1 U13716 ( .A1(n14210), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n12082) );
  NAND4_X1 U13717 ( .A1(n12085), .A2(n12084), .A3(n12083), .A4(n12082), .ZN(
        n12086) );
  NOR2_X1 U13718 ( .A1(n12087), .A2(n12086), .ZN(n12089) );
  NAND2_X1 U13719 ( .A1(n14295), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12088) );
  NAND4_X1 U13720 ( .A1(n12091), .A2(n12090), .A3(n12089), .A4(n12088), .ZN(
        n15397) );
  INV_X1 U13721 ( .A(n15397), .ZN(n12094) );
  NAND2_X1 U13722 ( .A1(n12021), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n12093) );
  AOI22_X1 U13723 ( .A1(n13660), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n11015), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12092) );
  OAI211_X1 U13724 ( .C1(n12094), .C2(n11008), .A(n12093), .B(n12092), .ZN(
        n14936) );
  AOI22_X1 U13725 ( .A1(n14269), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14270), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12098) );
  AOI22_X1 U13726 ( .A1(n14278), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14150), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12097) );
  AOI22_X1 U13727 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14152), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12096) );
  AOI22_X1 U13728 ( .A1(n14151), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12095) );
  NAND4_X1 U13729 ( .A1(n12098), .A2(n12097), .A3(n12096), .A4(n12095), .ZN(
        n12107) );
  AOI22_X1 U13730 ( .A1(n14253), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14287), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12105) );
  AOI22_X1 U13731 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12104) );
  INV_X1 U13732 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12100) );
  NOR2_X1 U13733 ( .A1(n12100), .A2(n12099), .ZN(n12101) );
  AOI21_X1 U13734 ( .B1(n14288), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n12101), .ZN(n12103) );
  AOI22_X1 U13735 ( .A1(n14210), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14273), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12102) );
  NAND4_X1 U13736 ( .A1(n12105), .A2(n12104), .A3(n12103), .A4(n12102), .ZN(
        n12106) );
  NOR2_X1 U13737 ( .A1(n12107), .A2(n12106), .ZN(n15482) );
  NAND2_X1 U13738 ( .A1(n12418), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n12109) );
  AOI22_X1 U13739 ( .A1(n13660), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n11015), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12108) );
  OAI211_X1 U13740 ( .C1(n15482), .C2(n11008), .A(n12109), .B(n12108), .ZN(
        n15135) );
  NAND2_X1 U13741 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12113) );
  NAND2_X1 U13742 ( .A1(n14270), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12112) );
  NAND2_X1 U13743 ( .A1(n14269), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12111) );
  AOI22_X1 U13744 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n14210), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12110) );
  AND4_X1 U13745 ( .A1(n12113), .A2(n12112), .A3(n12111), .A4(n12110), .ZN(
        n12128) );
  NAND2_X1 U13746 ( .A1(n14278), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n12117) );
  NAND2_X1 U13747 ( .A1(n14150), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12116) );
  NAND2_X1 U13748 ( .A1(n14151), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n12115) );
  NAND2_X1 U13749 ( .A1(n14152), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12114) );
  AND4_X1 U13750 ( .A1(n12117), .A2(n12116), .A3(n12115), .A4(n12114), .ZN(
        n12127) );
  INV_X1 U13751 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12118) );
  INV_X1 U13752 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14450) );
  OAI22_X1 U13753 ( .A1(n12118), .A2(n14285), .B1(n14284), .B2(n14450), .ZN(
        n12124) );
  NAND2_X1 U13754 ( .A1(n14287), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n12122) );
  NAND2_X1 U13755 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n12121) );
  NAND2_X1 U13756 ( .A1(n14273), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n12120) );
  NAND2_X1 U13757 ( .A1(n14288), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n12119) );
  NAND4_X1 U13758 ( .A1(n12122), .A2(n12121), .A3(n12120), .A4(n12119), .ZN(
        n12123) );
  NOR2_X1 U13759 ( .A1(n12124), .A2(n12123), .ZN(n12126) );
  NAND2_X1 U13760 ( .A1(n14295), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12125) );
  NAND4_X1 U13761 ( .A1(n12128), .A2(n12127), .A3(n12126), .A4(n12125), .ZN(
        n15461) );
  INV_X1 U13762 ( .A(n15461), .ZN(n12131) );
  NAND2_X1 U13763 ( .A1(n12418), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n12130) );
  AOI22_X1 U13764 ( .A1(n13660), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n11015), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12129) );
  OAI211_X1 U13765 ( .C1(n12131), .C2(n11008), .A(n12130), .B(n12129), .ZN(
        n17145) );
  NAND2_X1 U13766 ( .A1(n12418), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n12144) );
  AOI22_X1 U13767 ( .A1(n13660), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n11015), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12143) );
  AOI22_X1 U13768 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n14270), .B1(
        n14269), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12135) );
  AOI22_X1 U13769 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n14150), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12134) );
  AOI22_X1 U13770 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n14152), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12133) );
  AOI22_X1 U13771 ( .A1(n14151), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12132) );
  NAND4_X1 U13772 ( .A1(n12135), .A2(n12134), .A3(n12133), .A4(n12132), .ZN(
        n12141) );
  AOI22_X1 U13773 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n14287), .B1(
        n14253), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12139) );
  AOI22_X1 U13774 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12138) );
  AOI22_X1 U13775 ( .A1(n14288), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n14295), .ZN(n12137) );
  AOI22_X1 U13776 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n14210), .B1(
        n14273), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12136) );
  NAND4_X1 U13777 ( .A1(n12139), .A2(n12138), .A3(n12137), .A4(n12136), .ZN(
        n12140) );
  OR2_X1 U13778 ( .A1(n12141), .A2(n12140), .ZN(n15576) );
  NAND2_X1 U13779 ( .A1(n11007), .A2(n15576), .ZN(n12142) );
  NAND2_X1 U13780 ( .A1(n12021), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n12146) );
  AOI22_X1 U13781 ( .A1(n13660), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n11015), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12145) );
  NAND2_X1 U13782 ( .A1(n12418), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n12148) );
  AOI22_X1 U13783 ( .A1(n13660), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n11015), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12147) );
  NAND2_X1 U13784 ( .A1(n12148), .A2(n12147), .ZN(n15749) );
  NAND2_X1 U13785 ( .A1(n12418), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n12150) );
  AOI22_X1 U13786 ( .A1(n13660), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n11015), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12149) );
  NAND2_X1 U13787 ( .A1(n12150), .A2(n12149), .ZN(n15641) );
  AOI222_X1 U13788 ( .A1(n12021), .A2(P2_REIP_REG_19__SCAN_IN), .B1(n13660), 
        .B2(P2_EAX_REG_19__SCAN_IN), .C1(n11015), .C2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15929) );
  NAND2_X1 U13789 ( .A1(n12418), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n12152) );
  AOI22_X1 U13790 ( .A1(n13660), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n11015), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12151) );
  NAND2_X1 U13791 ( .A1(n12152), .A2(n12151), .ZN(n15950) );
  NAND2_X1 U13792 ( .A1(n12418), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12154) );
  AOI22_X1 U13793 ( .A1(n13660), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n11015), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12153) );
  AND2_X1 U13794 ( .A1(n12154), .A2(n12153), .ZN(n16762) );
  NAND2_X1 U13795 ( .A1(n12021), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12156) );
  AOI22_X1 U13796 ( .A1(n13660), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n11015), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12155) );
  AND2_X1 U13797 ( .A1(n12156), .A2(n12155), .ZN(n16620) );
  NOR2_X2 U13798 ( .A1(n16619), .A2(n16620), .ZN(n12159) );
  INV_X1 U13799 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n17755) );
  AOI22_X1 U13800 ( .A1(n13660), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n11015), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12157) );
  OAI21_X1 U13801 ( .B1(n12429), .B2(n17755), .A(n12157), .ZN(n12158) );
  OR2_X1 U13802 ( .A1(n12159), .A2(n12158), .ZN(n12160) );
  NAND2_X1 U13803 ( .A1(n12415), .A2(n12160), .ZN(n18791) );
  NAND2_X1 U13804 ( .A1(n12161), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n16827) );
  INV_X1 U13805 ( .A(n17044), .ZN(n12163) );
  NAND2_X1 U13806 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12162) );
  OAI211_X1 U13807 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n12164), .A(
        n12163), .B(n12162), .ZN(n12165) );
  OAI211_X1 U13808 ( .C1(n17229), .C2(n18791), .A(n16827), .B(n12165), .ZN(
        n12166) );
  AOI21_X1 U13809 ( .B1(n17047), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n12166), .ZN(n12167) );
  OAI21_X1 U13810 ( .B1(n18792), .B2(n18885), .A(n12167), .ZN(n12168) );
  AOI21_X1 U13811 ( .B1(n16832), .B2(n18879), .A(n12168), .ZN(n12329) );
  NAND2_X1 U13812 ( .A1(n12169), .A2(n12202), .ZN(n12185) );
  NAND2_X1 U13813 ( .A1(n11394), .A2(n12170), .ZN(n12172) );
  NAND2_X1 U13814 ( .A1(n12172), .A2(n12171), .ZN(n12174) );
  NOR2_X1 U13815 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n12175) );
  MUX2_X1 U13816 ( .A(n12176), .B(n12175), .S(n19633), .Z(n12212) );
  INV_X1 U13817 ( .A(n12205), .ZN(n12178) );
  MUX2_X1 U13818 ( .A(n12180), .B(n12179), .S(n19633), .Z(n12222) );
  NAND2_X1 U13819 ( .A1(n19633), .A2(n14974), .ZN(n12182) );
  NAND2_X1 U13820 ( .A1(n12183), .A2(n12182), .ZN(n12233) );
  MUX2_X1 U13821 ( .A(n12184), .B(P2_EBX_REG_6__SCAN_IN), .S(n19633), .Z(
        n12187) );
  XNOR2_X1 U13822 ( .A(n12186), .B(n12187), .ZN(n18623) );
  NAND2_X1 U13823 ( .A1(n12185), .A2(n18623), .ZN(n12239) );
  XNOR2_X1 U13824 ( .A(n12239), .B(n17268), .ZN(n16978) );
  MUX2_X1 U13825 ( .A(n12190), .B(n12189), .S(n19633), .Z(n12199) );
  NAND2_X1 U13826 ( .A1(n19633), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12196) );
  NAND2_X1 U13827 ( .A1(n19633), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12193) );
  NAND2_X1 U13828 ( .A1(n19633), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12244) );
  XNOR2_X1 U13829 ( .A(n12246), .B(n12244), .ZN(n18658) );
  AOI21_X1 U13830 ( .B1(n18658), .B2(n13735), .A(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16982) );
  INV_X1 U13831 ( .A(n16982), .ZN(n12201) );
  XNOR2_X1 U13832 ( .A(n12194), .B(n12193), .ZN(n15760) );
  NAND2_X1 U13833 ( .A1(n15760), .A2(n13735), .ZN(n12195) );
  INV_X1 U13834 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17221) );
  NAND2_X1 U13835 ( .A1(n12195), .A2(n17221), .ZN(n17211) );
  XNOR2_X1 U13836 ( .A(n12197), .B(n12196), .ZN(n18645) );
  NAND2_X1 U13837 ( .A1(n18645), .A2(n13735), .ZN(n12238) );
  NAND2_X1 U13838 ( .A1(n12238), .A2(n17232), .ZN(n16992) );
  XNOR2_X1 U13839 ( .A(n12198), .B(n12199), .ZN(n18636) );
  INV_X1 U13840 ( .A(n18636), .ZN(n12200) );
  NAND2_X1 U13841 ( .A1(n12200), .A2(n17252), .ZN(n17241) );
  AND2_X1 U13842 ( .A1(n16992), .A2(n17241), .ZN(n17209) );
  AND2_X1 U13843 ( .A1(n17211), .A2(n17209), .ZN(n16980) );
  AND2_X1 U13844 ( .A1(n12201), .A2(n16980), .ZN(n12241) );
  NAND2_X1 U13845 ( .A1(n12203), .A2(n12202), .ZN(n12206) );
  INV_X1 U13846 ( .A(n12211), .ZN(n12204) );
  XNOR2_X1 U13847 ( .A(n12205), .B(n12204), .ZN(n15685) );
  NAND2_X1 U13848 ( .A1(n12206), .A2(n15685), .ZN(n12219) );
  XNOR2_X1 U13849 ( .A(n12219), .B(n15699), .ZN(n15514) );
  INV_X1 U13850 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n14764) );
  MUX2_X1 U13851 ( .A(n12207), .B(n14764), .S(n19633), .Z(n18598) );
  NOR2_X1 U13852 ( .A1(n18598), .A2(n17662), .ZN(n12215) );
  INV_X1 U13853 ( .A(n12215), .ZN(n17664) );
  INV_X1 U13854 ( .A(n12212), .ZN(n12210) );
  AND2_X1 U13855 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n12208) );
  NAND2_X1 U13856 ( .A1(n19633), .A2(n12208), .ZN(n12209) );
  NAND2_X1 U13857 ( .A1(n12210), .A2(n12209), .ZN(n18608) );
  NAND2_X1 U13858 ( .A1(n17664), .A2(n18608), .ZN(n16013) );
  OAI21_X1 U13859 ( .B1(n12213), .B2(n12212), .A(n12211), .ZN(n15729) );
  XNOR2_X1 U13860 ( .A(n15729), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n16014) );
  INV_X1 U13861 ( .A(n18608), .ZN(n12214) );
  NAND2_X1 U13862 ( .A1(n12215), .A2(n12214), .ZN(n14626) );
  NAND2_X1 U13863 ( .A1(n14624), .A2(n14626), .ZN(n16012) );
  AND2_X1 U13864 ( .A1(n16014), .A2(n16012), .ZN(n12216) );
  NAND2_X1 U13865 ( .A1(n16013), .A2(n12216), .ZN(n16017) );
  INV_X1 U13866 ( .A(n15729), .ZN(n12217) );
  NAND2_X1 U13867 ( .A1(n12217), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12218) );
  NAND2_X1 U13868 ( .A1(n16017), .A2(n12218), .ZN(n15513) );
  NAND2_X1 U13869 ( .A1(n12219), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15693) );
  INV_X1 U13870 ( .A(n12220), .ZN(n12226) );
  INV_X1 U13871 ( .A(n12221), .ZN(n12224) );
  INV_X1 U13872 ( .A(n12222), .ZN(n12223) );
  NAND2_X1 U13873 ( .A1(n12224), .A2(n12223), .ZN(n12225) );
  NAND2_X1 U13874 ( .A1(n12226), .A2(n12225), .ZN(n15606) );
  INV_X1 U13875 ( .A(n15606), .ZN(n12227) );
  NAND2_X1 U13876 ( .A1(n12227), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12228) );
  AND2_X1 U13877 ( .A1(n15693), .A2(n12228), .ZN(n12230) );
  INV_X1 U13878 ( .A(n12228), .ZN(n12229) );
  XNOR2_X1 U13879 ( .A(n15606), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n15694) );
  NAND3_X1 U13880 ( .A1(n12232), .A2(n12202), .A3(n12231), .ZN(n12234) );
  XNOR2_X1 U13881 ( .A(n12220), .B(n12233), .ZN(n15722) );
  NAND2_X1 U13882 ( .A1(n12234), .A2(n15722), .ZN(n12235) );
  XNOR2_X1 U13883 ( .A(n12235), .B(n15771), .ZN(n15768) );
  NAND2_X1 U13884 ( .A1(n15766), .A2(n15768), .ZN(n15767) );
  NAND2_X1 U13885 ( .A1(n12235), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12236) );
  NAND2_X1 U13886 ( .A1(n15767), .A2(n12236), .ZN(n17270) );
  NAND2_X1 U13887 ( .A1(n12237), .A2(n17270), .ZN(n12243) );
  NOR2_X1 U13888 ( .A1(n12238), .A2(n17232), .ZN(n16994) );
  AND2_X1 U13889 ( .A1(n18636), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17242) );
  NOR2_X1 U13890 ( .A1(n16994), .A2(n17242), .ZN(n12240) );
  NAND2_X1 U13891 ( .A1(n12239), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16979) );
  NAND2_X1 U13892 ( .A1(n12243), .A2(n12242), .ZN(n16966) );
  INV_X1 U13893 ( .A(n12244), .ZN(n12245) );
  NAND2_X1 U13894 ( .A1(n19633), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n12248) );
  INV_X1 U13895 ( .A(n12247), .ZN(n12250) );
  INV_X1 U13896 ( .A(n12248), .ZN(n12249) );
  NAND2_X1 U13897 ( .A1(n12250), .A2(n12249), .ZN(n12251) );
  NAND2_X1 U13898 ( .A1(n12257), .A2(n12251), .ZN(n14569) );
  OR2_X1 U13899 ( .A1(n14569), .A2(n12202), .ZN(n12252) );
  INV_X1 U13900 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17184) );
  NAND2_X1 U13901 ( .A1(n12252), .A2(n17184), .ZN(n16964) );
  AND2_X2 U13902 ( .A1(n16966), .A2(n16964), .ZN(n16850) );
  INV_X1 U13903 ( .A(n12252), .ZN(n12253) );
  NAND2_X1 U13904 ( .A1(n12253), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16965) );
  AND2_X1 U13905 ( .A1(n13735), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12254) );
  AND2_X1 U13906 ( .A1(n13735), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12255) );
  AND2_X1 U13907 ( .A1(n18658), .A2(n12255), .ZN(n16981) );
  NOR2_X1 U13908 ( .A1(n17215), .A2(n16981), .ZN(n12256) );
  NAND2_X1 U13909 ( .A1(n16965), .A2(n12256), .ZN(n16851) );
  AND2_X1 U13910 ( .A1(n19633), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12258) );
  NAND2_X1 U13911 ( .A1(n12257), .A2(n12258), .ZN(n12259) );
  NAND2_X1 U13912 ( .A1(n12279), .A2(n12259), .ZN(n18671) );
  NAND2_X1 U13913 ( .A1(n13735), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12260) );
  OR2_X1 U13914 ( .A1(n18671), .A2(n12260), .ZN(n16953) );
  NAND2_X1 U13915 ( .A1(n16956), .A2(n16953), .ZN(n16917) );
  AND2_X1 U13916 ( .A1(n19633), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n12278) );
  AND2_X1 U13917 ( .A1(n19633), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12273) );
  NAND2_X1 U13918 ( .A1(n19633), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n12270) );
  NAND2_X1 U13919 ( .A1(n19633), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12283) );
  AND2_X1 U13920 ( .A1(n19633), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n12265) );
  AND2_X1 U13921 ( .A1(n19633), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12261) );
  NAND2_X1 U13922 ( .A1(n19633), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n12288) );
  XNOR2_X1 U13923 ( .A(n11029), .B(n12288), .ZN(n18745) );
  NAND2_X1 U13924 ( .A1(n18745), .A2(n13735), .ZN(n12298) );
  INV_X1 U13925 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17072) );
  NAND2_X1 U13926 ( .A1(n12298), .A2(n17072), .ZN(n16882) );
  NAND2_X1 U13927 ( .A1(n12262), .A2(n12261), .ZN(n12263) );
  NAND2_X1 U13928 ( .A1(n11029), .A2(n12263), .ZN(n18734) );
  INV_X1 U13929 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17096) );
  NAND2_X1 U13930 ( .A1(n16893), .A2(n17096), .ZN(n12264) );
  NAND2_X1 U13931 ( .A1(n16882), .A2(n12264), .ZN(n16861) );
  INV_X1 U13932 ( .A(n12265), .ZN(n12266) );
  XNOR2_X1 U13933 ( .A(n12267), .B(n12266), .ZN(n18720) );
  AOI21_X1 U13934 ( .B1(n18720), .B2(n13735), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16901) );
  INV_X1 U13935 ( .A(n12268), .ZN(n12284) );
  INV_X1 U13936 ( .A(n12269), .ZN(n12275) );
  INV_X1 U13937 ( .A(n12270), .ZN(n12271) );
  NAND2_X1 U13938 ( .A1(n12275), .A2(n12271), .ZN(n12272) );
  AND2_X1 U13939 ( .A1(n12284), .A2(n12272), .ZN(n18694) );
  NAND2_X1 U13940 ( .A1(n18694), .A2(n13735), .ZN(n12302) );
  INV_X1 U13941 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17129) );
  NAND2_X1 U13942 ( .A1(n12302), .A2(n17129), .ZN(n16920) );
  NAND2_X1 U13943 ( .A1(n12281), .A2(n12273), .ZN(n12274) );
  NAND2_X1 U13944 ( .A1(n12275), .A2(n12274), .ZN(n18682) );
  OR2_X1 U13945 ( .A1(n18682), .A2(n12202), .ZN(n12276) );
  INV_X1 U13946 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17150) );
  NAND2_X1 U13947 ( .A1(n12276), .A2(n17150), .ZN(n16919) );
  OR2_X1 U13948 ( .A1(n18671), .A2(n12202), .ZN(n12277) );
  INV_X1 U13949 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17177) );
  NAND2_X1 U13950 ( .A1(n12277), .A2(n17177), .ZN(n16954) );
  NAND2_X1 U13951 ( .A1(n12279), .A2(n12278), .ZN(n12280) );
  AND2_X1 U13952 ( .A1(n12281), .A2(n12280), .ZN(n15671) );
  NAND2_X1 U13953 ( .A1(n15671), .A2(n13735), .ZN(n12305) );
  INV_X1 U13954 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17157) );
  NAND2_X1 U13955 ( .A1(n12305), .A2(n17157), .ZN(n16943) );
  AND3_X1 U13956 ( .A1(n16919), .A2(n16954), .A3(n16943), .ZN(n12282) );
  NAND2_X1 U13957 ( .A1(n16920), .A2(n12282), .ZN(n16848) );
  XNOR2_X1 U13958 ( .A(n12284), .B(n12283), .ZN(n18704) );
  NAND2_X1 U13959 ( .A1(n18704), .A2(n13735), .ZN(n12285) );
  INV_X1 U13960 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17112) );
  NAND2_X1 U13961 ( .A1(n12285), .A2(n17112), .ZN(n12287) );
  AND2_X1 U13962 ( .A1(n13735), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12286) );
  NAND2_X1 U13963 ( .A1(n18704), .A2(n12286), .ZN(n16858) );
  NAND2_X1 U13964 ( .A1(n12287), .A2(n16858), .ZN(n16857) );
  NOR4_X1 U13965 ( .A1(n16861), .A2(n16901), .A3(n16848), .A4(n16857), .ZN(
        n12289) );
  NAND2_X1 U13966 ( .A1(n19633), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12311) );
  NAND2_X1 U13967 ( .A1(n19633), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12292) );
  XOR2_X1 U13968 ( .A(n12311), .B(n12312), .Z(n18777) );
  NAND2_X1 U13969 ( .A1(n18777), .A2(n13735), .ZN(n12296) );
  INV_X1 U13970 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17043) );
  NAND2_X1 U13971 ( .A1(n12296), .A2(n17043), .ZN(n16866) );
  AND2_X1 U13972 ( .A1(n12289), .A2(n16866), .ZN(n12290) );
  INV_X1 U13973 ( .A(n12291), .ZN(n12293) );
  XNOR2_X1 U13974 ( .A(n12293), .B(n12292), .ZN(n18766) );
  NAND2_X1 U13975 ( .A1(n18766), .A2(n13735), .ZN(n16863) );
  NAND2_X1 U13976 ( .A1(n16863), .A2(n16877), .ZN(n12295) );
  INV_X1 U13977 ( .A(n12296), .ZN(n12297) );
  NAND2_X1 U13978 ( .A1(n12297), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16865) );
  INV_X1 U13979 ( .A(n16865), .ZN(n12310) );
  OR2_X1 U13980 ( .A1(n12298), .A2(n17072), .ZN(n16883) );
  INV_X1 U13981 ( .A(n16893), .ZN(n12299) );
  NAND2_X1 U13982 ( .A1(n12299), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12300) );
  AND2_X1 U13983 ( .A1(n13735), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12301) );
  INV_X1 U13984 ( .A(n12302), .ZN(n12303) );
  NAND2_X1 U13985 ( .A1(n12303), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16921) );
  NAND2_X1 U13986 ( .A1(n13735), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12304) );
  OR2_X1 U13987 ( .A1(n18682), .A2(n12304), .ZN(n16918) );
  NAND2_X1 U13988 ( .A1(n16921), .A2(n16918), .ZN(n16854) );
  INV_X1 U13989 ( .A(n16858), .ZN(n12307) );
  INV_X1 U13990 ( .A(n12305), .ZN(n12306) );
  NOR4_X1 U13991 ( .A1(n16900), .A2(n16854), .A3(n12307), .A4(n16942), .ZN(
        n12308) );
  NAND2_X1 U13992 ( .A1(n16862), .A2(n12308), .ZN(n12309) );
  AND2_X1 U13993 ( .A1(n19633), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12313) );
  NAND2_X1 U13994 ( .A1(n12314), .A2(n12313), .ZN(n12315) );
  NAND2_X1 U13995 ( .A1(n12319), .A2(n12315), .ZN(n16629) );
  NOR2_X1 U13996 ( .A1(n16629), .A2(n12202), .ZN(n12316) );
  AND2_X1 U13997 ( .A1(n12316), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16838) );
  INV_X1 U13998 ( .A(n12316), .ZN(n12318) );
  INV_X1 U13999 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12317) );
  NAND2_X1 U14000 ( .A1(n12318), .A2(n12317), .ZN(n16836) );
  OAI21_X2 U14001 ( .B1(n16835), .B2(n16838), .A(n16836), .ZN(n13705) );
  NAND2_X1 U14002 ( .A1(n19633), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12403) );
  XNOR2_X1 U14003 ( .A(n12319), .B(n12403), .ZN(n18790) );
  INV_X1 U14004 ( .A(n12320), .ZN(n12322) );
  NAND2_X1 U14005 ( .A1(n11051), .A2(n13704), .ZN(n12323) );
  XNOR2_X1 U14006 ( .A(n13705), .B(n12323), .ZN(n16834) );
  INV_X1 U14007 ( .A(n16834), .ZN(n12327) );
  NAND2_X1 U14008 ( .A1(n15317), .A2(n11394), .ZN(n12324) );
  NAND2_X1 U14009 ( .A1(n12327), .A2(n12326), .ZN(n12328) );
  NAND2_X1 U14010 ( .A1(n12329), .A2(n12328), .ZN(P2_U3023) );
  AND2_X2 U14011 ( .A1(n12340), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12353) );
  NAND2_X2 U14012 ( .A1(n12353), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12352) );
  NOR2_X4 U14013 ( .A1(n12352), .A2(n16947), .ZN(n12339) );
  INV_X1 U14014 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16925) );
  INV_X1 U14015 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16888) );
  INV_X1 U14016 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16828) );
  INV_X1 U14017 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16811) );
  INV_X1 U14018 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12365) );
  INV_X1 U14019 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14525) );
  AND2_X2 U14020 ( .A1(n12370), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12369) );
  AND2_X2 U14021 ( .A1(n12369), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12374) );
  INV_X1 U14022 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12332) );
  XNOR2_X2 U14023 ( .A(n12333), .B(n12332), .ZN(n16773) );
  INV_X1 U14024 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12334) );
  AOI22_X2 U14025 ( .A1(n16773), .A2(n11407), .B1(n12334), .B2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n12336) );
  BUF_X4 U14026 ( .A(n12336), .Z(n18752) );
  AOI21_X1 U14027 ( .B1(n14525), .B2(n12368), .A(n12370), .ZN(n16603) );
  OAI21_X1 U14028 ( .B1(n12335), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n12363), .ZN(n16823) );
  INV_X1 U14029 ( .A(n16823), .ZN(n18807) );
  INV_X4 U14030 ( .A(n12336), .ZN(n18717) );
  OAI21_X1 U14031 ( .B1(n12337), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n12361), .ZN(n16843) );
  INV_X1 U14032 ( .A(n16843), .ZN(n16614) );
  CLKBUF_X1 U14033 ( .A(n12338), .Z(n12359) );
  AOI21_X1 U14034 ( .B1(n16888), .B2(n12357), .A(n12359), .ZN(n18753) );
  AOI21_X1 U14035 ( .B1(n12330), .B2(n12355), .A(n12358), .ZN(n18719) );
  AOI21_X1 U14036 ( .B1(n16925), .B2(n12354), .A(n12356), .ZN(n18693) );
  AOI21_X1 U14037 ( .B1(n16947), .B2(n12352), .A(n12339), .ZN(n16949) );
  NOR2_X1 U14038 ( .A1(n12340), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12341) );
  NOR2_X1 U14039 ( .A1(n12353), .A2(n12341), .ZN(n16971) );
  AOI21_X1 U14040 ( .B1(n17659), .B2(n12349), .A(n12342), .ZN(n17646) );
  CLKBUF_X1 U14041 ( .A(n12343), .Z(n12350) );
  AOI21_X1 U14042 ( .B1(n17645), .B2(n12347), .A(n12350), .ZN(n18634) );
  AOI21_X1 U14043 ( .B1(n17622), .B2(n12345), .A(n12348), .ZN(n17624) );
  AOI21_X1 U14044 ( .B1(n15681), .B2(n12344), .A(n12346), .ZN(n15679) );
  INV_X1 U14045 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18601) );
  AOI22_X1 U14046 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n17662), .B1(n18601), 
        .B2(n11407), .ZN(n18595) );
  AOI22_X1 U14047 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14624), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n11407), .ZN(n17279) );
  NOR2_X1 U14048 ( .A1(n18595), .A2(n17279), .ZN(n17278) );
  OAI21_X1 U14049 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n12344), .ZN(n17610) );
  NAND2_X1 U14050 ( .A1(n17278), .A2(n17610), .ZN(n15677) );
  NOR2_X1 U14051 ( .A1(n15679), .A2(n15677), .ZN(n15597) );
  OAI21_X1 U14052 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12346), .A(
        n12345), .ZN(n17614) );
  NAND2_X1 U14053 ( .A1(n15597), .A2(n17614), .ZN(n15714) );
  NOR2_X1 U14054 ( .A1(n17624), .A2(n15714), .ZN(n18618) );
  OAI21_X1 U14055 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n12348), .A(
        n12347), .ZN(n18620) );
  NAND2_X1 U14056 ( .A1(n18618), .A2(n18620), .ZN(n18633) );
  NOR2_X1 U14057 ( .A1(n18634), .A2(n18633), .ZN(n18649) );
  OAI21_X1 U14058 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n12350), .A(
        n12349), .ZN(n18650) );
  NAND2_X1 U14059 ( .A1(n18649), .A2(n18650), .ZN(n15757) );
  NOR2_X1 U14060 ( .A1(n17646), .A2(n15757), .ZN(n18662) );
  NOR2_X1 U14061 ( .A1(n12342), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12351) );
  OR2_X1 U14062 ( .A1(n12340), .A2(n12351), .ZN(n18663) );
  NAND2_X1 U14063 ( .A1(n18662), .A2(n18663), .ZN(n14566) );
  NOR2_X1 U14064 ( .A1(n16971), .A2(n14566), .ZN(n18673) );
  OAI21_X1 U14065 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n12353), .A(
        n12352), .ZN(n18674) );
  NAND2_X1 U14066 ( .A1(n18673), .A2(n18674), .ZN(n15665) );
  NOR2_X1 U14067 ( .A1(n16949), .A2(n15665), .ZN(n18684) );
  OAI21_X1 U14068 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n12339), .A(
        n12354), .ZN(n18685) );
  NAND2_X1 U14069 ( .A1(n18684), .A2(n18685), .ZN(n18691) );
  NOR2_X1 U14070 ( .A1(n18693), .A2(n18691), .ZN(n18708) );
  OAI21_X1 U14071 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12356), .A(
        n12355), .ZN(n18709) );
  NAND2_X1 U14072 ( .A1(n18708), .A2(n18709), .ZN(n18718) );
  NOR2_X1 U14073 ( .A1(n18719), .A2(n18718), .ZN(n18716) );
  OAI21_X1 U14074 ( .B1(n12358), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n12357), .ZN(n18737) );
  NAND2_X1 U14075 ( .A1(n18716), .A2(n18737), .ZN(n18751) );
  NOR2_X1 U14076 ( .A1(n18753), .A2(n18751), .ZN(n18772) );
  OAI21_X1 U14077 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12359), .A(
        n12360), .ZN(n18775) );
  NAND2_X1 U14078 ( .A1(n18772), .A2(n18775), .ZN(n18783) );
  INV_X1 U14079 ( .A(n18781), .ZN(n18771) );
  AOI21_X1 U14080 ( .B1(n12360), .B2(n12331), .A(n12337), .ZN(n16870) );
  INV_X1 U14081 ( .A(n16870), .ZN(n18782) );
  NOR2_X1 U14082 ( .A1(n18782), .A2(n18717), .ZN(n18784) );
  NOR2_X1 U14083 ( .A1(n16612), .A2(n18717), .ZN(n18796) );
  AOI21_X1 U14084 ( .B1(n16828), .B2(n12361), .A(n12335), .ZN(n18795) );
  NOR2_X1 U14085 ( .A1(n18717), .A2(n18794), .ZN(n18808) );
  NOR2_X1 U14086 ( .A1(n18806), .A2(n18717), .ZN(n18822) );
  INV_X1 U14087 ( .A(n12366), .ZN(n12362) );
  AOI21_X1 U14088 ( .B1(n16811), .B2(n12363), .A(n12362), .ZN(n18823) );
  AND2_X1 U14089 ( .A1(n18752), .A2(n18823), .ZN(n12364) );
  NAND2_X1 U14090 ( .A1(n12366), .A2(n12365), .ZN(n12367) );
  NAND2_X1 U14091 ( .A1(n12368), .A2(n12367), .ZN(n18832) );
  OAI21_X1 U14092 ( .B1(n16603), .B2(n16602), .A(n18752), .ZN(n18845) );
  NOR2_X1 U14093 ( .A1(n12370), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12371) );
  OR2_X1 U14094 ( .A1(n12369), .A2(n12371), .ZN(n18844) );
  NAND2_X1 U14095 ( .A1(n18845), .A2(n18844), .ZN(n18843) );
  NAND2_X1 U14096 ( .A1(n18843), .A2(n18752), .ZN(n18863) );
  INV_X1 U14097 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12373) );
  INV_X1 U14098 ( .A(n12369), .ZN(n12372) );
  AOI21_X1 U14099 ( .B1(n12373), .B2(n12372), .A(n12374), .ZN(n16789) );
  INV_X1 U14100 ( .A(n16789), .ZN(n18862) );
  NAND2_X1 U14101 ( .A1(n18863), .A2(n18862), .ZN(n18860) );
  NAND2_X1 U14102 ( .A1(n18752), .A2(n18860), .ZN(n12375) );
  XNOR2_X1 U14103 ( .A(n12374), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13747) );
  NAND2_X1 U14104 ( .A1(n12375), .A2(n13747), .ZN(n13672) );
  OAI211_X1 U14105 ( .C1(n12375), .C2(n13747), .A(n18861), .B(n13672), .ZN(
        n12444) );
  INV_X1 U14106 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n12378) );
  NAND2_X1 U14107 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12377) );
  NAND2_X1 U14108 ( .A1(n12390), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12376) );
  OAI211_X1 U14109 ( .C1(n11833), .C2(n12378), .A(n12377), .B(n12376), .ZN(
        n12379) );
  AOI21_X1 U14110 ( .B1(n12398), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n12379), .ZN(n16670) );
  INV_X1 U14111 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n12382) );
  NAND2_X1 U14112 ( .A1(n12398), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12381) );
  AOI22_X1 U14113 ( .A1(n13678), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n12380) );
  OAI211_X1 U14114 ( .C1(n11833), .C2(n12382), .A(n12381), .B(n12380), .ZN(
        n16666) );
  INV_X1 U14115 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n12385) );
  NAND2_X1 U14116 ( .A1(n12398), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12384) );
  AOI22_X1 U14117 ( .A1(n13678), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n12383) );
  OAI211_X1 U14118 ( .C1(n11464), .C2(n12385), .A(n12384), .B(n12383), .ZN(
        n16656) );
  INV_X1 U14119 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n12388) );
  NAND2_X1 U14120 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12387) );
  NAND2_X1 U14121 ( .A1(n12390), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12386) );
  OAI211_X1 U14122 ( .C1(n11833), .C2(n12388), .A(n12387), .B(n12386), .ZN(
        n12389) );
  AOI21_X1 U14123 ( .B1(n12398), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n12389), .ZN(n14501) );
  INV_X1 U14124 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n12393) );
  NAND2_X1 U14125 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12392) );
  NAND2_X1 U14126 ( .A1(n12390), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12391) );
  OAI211_X1 U14127 ( .C1(n11833), .C2(n12393), .A(n12392), .B(n12391), .ZN(
        n12394) );
  AOI21_X1 U14128 ( .B1(n12398), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n12394), .ZN(n15985) );
  INV_X1 U14129 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n12397) );
  NAND2_X1 U14130 ( .A1(n12398), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12396) );
  AOI22_X1 U14131 ( .A1(n13678), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n12395) );
  OAI211_X1 U14132 ( .C1(n11833), .C2(n12397), .A(n12396), .B(n12395), .ZN(
        n16634) );
  NAND2_X1 U14133 ( .A1(n16635), .A2(n16634), .ZN(n13675) );
  INV_X1 U14134 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n12401) );
  NAND2_X1 U14135 ( .A1(n12398), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12400) );
  AOI22_X1 U14136 ( .A1(n13678), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n12399) );
  OAI211_X1 U14137 ( .C1(n11464), .C2(n12401), .A(n12400), .B(n12399), .ZN(
        n13676) );
  NAND2_X1 U14138 ( .A1(n11943), .A2(n15319), .ZN(n15328) );
  NOR2_X1 U14139 ( .A1(n18589), .A2(n15313), .ZN(n12409) );
  NAND2_X1 U14140 ( .A1(n21819), .A2(n18908), .ZN(n12438) );
  INV_X1 U14141 ( .A(n12438), .ZN(n12402) );
  NAND2_X1 U14142 ( .A1(n12404), .A2(n12403), .ZN(n13707) );
  AND2_X1 U14143 ( .A1(n19633), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n13706) );
  NAND2_X1 U14144 ( .A1(n19633), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n13710) );
  INV_X1 U14145 ( .A(n13710), .ZN(n12405) );
  NAND2_X1 U14146 ( .A1(n19633), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n13716) );
  INV_X1 U14147 ( .A(n13722), .ZN(n12406) );
  NAND2_X1 U14148 ( .A1(n19633), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n13721) );
  NAND2_X1 U14149 ( .A1(n19633), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n13732) );
  NAND2_X1 U14150 ( .A1(n13731), .A2(n13732), .ZN(n13664) );
  NAND2_X1 U14151 ( .A1(n19633), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12407) );
  XNOR2_X1 U14152 ( .A(n13664), .B(n12407), .ZN(n13737) );
  INV_X1 U14153 ( .A(n13737), .ZN(n12410) );
  AND2_X1 U14154 ( .A1(n12438), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n12408) );
  NAND2_X1 U14155 ( .A1(n12409), .A2(n12408), .ZN(n18803) );
  AOI21_X1 U14156 ( .B1(n15993), .B2(n18811), .A(n12411), .ZN(n12443) );
  INV_X1 U14157 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12414) );
  NAND2_X1 U14158 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19470), .ZN(n18899) );
  NOR3_X1 U14159 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n19459), .A3(n18899), 
        .ZN(n18902) );
  OR2_X1 U14160 ( .A1(n16976), .A2(n18861), .ZN(n12412) );
  NOR2_X1 U14161 ( .A1(n18902), .A2(n12412), .ZN(n12413) );
  INV_X1 U14162 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n17763) );
  INV_X1 U14163 ( .A(n18850), .ZN(n18748) );
  OAI22_X1 U14164 ( .A1(n12414), .A2(n18621), .B1(n17763), .B2(n18748), .ZN(
        n12442) );
  NAND2_X1 U14165 ( .A1(n12418), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12417) );
  AOI22_X1 U14166 ( .A1(n13660), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n11015), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12416) );
  NAND2_X1 U14167 ( .A1(n12418), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12420) );
  AOI22_X1 U14168 ( .A1(n13660), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n11015), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12419) );
  AND2_X1 U14169 ( .A1(n12420), .A2(n12419), .ZN(n16738) );
  INV_X1 U14170 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n17758) );
  AOI22_X1 U14171 ( .A1(n13660), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n11015), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12421) );
  OAI21_X1 U14172 ( .B1(n12429), .B2(n17758), .A(n12421), .ZN(n16729) );
  INV_X1 U14173 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n17759) );
  AOI22_X1 U14174 ( .A1(n13660), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n11015), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12422) );
  OAI21_X1 U14175 ( .B1(n12429), .B2(n17759), .A(n12422), .ZN(n14512) );
  NAND2_X1 U14176 ( .A1(n12021), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12424) );
  AOI22_X1 U14177 ( .A1(n13660), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n11015), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12423) );
  AND2_X1 U14178 ( .A1(n12424), .A2(n12423), .ZN(n16060) );
  NAND2_X1 U14179 ( .A1(n12021), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n12426) );
  AOI22_X1 U14180 ( .A1(n13660), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n11015), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12425) );
  AND2_X1 U14181 ( .A1(n12426), .A2(n12425), .ZN(n16701) );
  INV_X1 U14182 ( .A(n16701), .ZN(n12427) );
  AOI22_X1 U14183 ( .A1(n13660), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n11015), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12428) );
  OAI21_X1 U14184 ( .B1(n12429), .B2(n17763), .A(n12428), .ZN(n12430) );
  INV_X1 U14185 ( .A(n16702), .ZN(n12432) );
  INV_X1 U14186 ( .A(n12430), .ZN(n12431) );
  NAND2_X1 U14187 ( .A1(n12432), .A2(n12431), .ZN(n12433) );
  NAND2_X1 U14188 ( .A1(n21819), .A2(n15326), .ZN(n12437) );
  INV_X1 U14189 ( .A(n12437), .ZN(n12434) );
  NAND2_X1 U14190 ( .A1(n12435), .A2(n12434), .ZN(n15338) );
  NAND2_X1 U14191 ( .A1(n15319), .A2(n18592), .ZN(n14578) );
  OR2_X1 U14192 ( .A1(n14578), .A2(n12436), .ZN(n14581) );
  NAND2_X1 U14193 ( .A1(n14616), .A2(n12437), .ZN(n13668) );
  INV_X1 U14194 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n13680) );
  NAND2_X1 U14195 ( .A1(n12438), .A2(n13680), .ZN(n12439) );
  OR2_X1 U14196 ( .A1(n14581), .A2(n12439), .ZN(n12440) );
  NAND2_X2 U14197 ( .A1(n13668), .A2(n12440), .ZN(n18852) );
  INV_X1 U14198 ( .A(n18852), .ZN(n18733) );
  OAI22_X1 U14199 ( .A1(n16074), .A2(n18855), .B1(n12401), .B2(n18733), .ZN(
        n12441) );
  NAND3_X1 U14200 ( .A1(n12444), .A2(n12443), .A3(n11242), .ZN(P2_U2825) );
  NOR2_X4 U14201 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15211) );
  AND2_X4 U14202 ( .A1(n12452), .A2(n15211), .ZN(n12645) );
  INV_X1 U14203 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12446) );
  AOI22_X1 U14204 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12686), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12451) );
  AND2_X4 U14205 ( .A1(n12452), .A2(n12454), .ZN(n12650) );
  AOI22_X1 U14206 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12629), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12450) );
  NAND2_X2 U14207 ( .A1(n15211), .A2(n15212), .ZN(n12460) );
  AOI22_X1 U14208 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12449) );
  AOI22_X1 U14209 ( .A1(n12685), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12518), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12459) );
  AOI22_X1 U14210 ( .A1(n12507), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12687), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12458) );
  AND2_X4 U14211 ( .A1(n12454), .A2(n15212), .ZN(n13192) );
  AOI22_X1 U14212 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12808), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12457) );
  AND2_X2 U14213 ( .A1(n12455), .A2(n15213), .ZN(n12693) );
  AOI22_X1 U14214 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12693), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12456) );
  AOI22_X1 U14215 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12686), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12464) );
  AOI22_X1 U14216 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12687), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12463) );
  AOI22_X1 U14217 ( .A1(n11017), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11022), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12462) );
  AOI22_X1 U14218 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12808), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12461) );
  NAND4_X1 U14219 ( .A1(n12464), .A2(n12463), .A3(n12462), .A4(n12461), .ZN(
        n12471) );
  AOI22_X1 U14220 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12469) );
  AOI22_X1 U14221 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12629), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12468) );
  AOI22_X1 U14222 ( .A1(n12685), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13187), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12467) );
  AOI22_X1 U14223 ( .A1(n12507), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12693), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12466) );
  NAND4_X1 U14224 ( .A1(n12469), .A2(n12468), .A3(n12467), .A4(n12466), .ZN(
        n12470) );
  NAND2_X1 U14225 ( .A1(n12685), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12473) );
  NAND2_X1 U14226 ( .A1(n13286), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12472) );
  AOI22_X1 U14227 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12629), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12476) );
  AOI22_X1 U14228 ( .A1(n12687), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12808), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12475) );
  AOI22_X1 U14229 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12693), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12474) );
  AOI22_X1 U14230 ( .A1(n12686), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11022), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12482) );
  AOI22_X1 U14231 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12480) );
  AOI22_X1 U14232 ( .A1(n12518), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13192), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12479) );
  AOI22_X1 U14233 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12507), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12478) );
  AOI22_X1 U14234 ( .A1(n12507), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12687), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12486) );
  AOI22_X1 U14235 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12808), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12485) );
  AOI22_X1 U14236 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12693), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12484) );
  NAND4_X1 U14237 ( .A1(n12487), .A2(n12486), .A3(n12485), .A4(n12484), .ZN(
        n12493) );
  AOI22_X1 U14238 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12686), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12491) );
  AOI22_X1 U14239 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12629), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12490) );
  AOI22_X1 U14240 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11021), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12489) );
  NAND4_X1 U14241 ( .A1(n12491), .A2(n12490), .A3(n12489), .A4(n12488), .ZN(
        n12492) );
  AND2_X1 U14242 ( .A1(n12558), .A2(n14811), .ZN(n12513) );
  AOI22_X1 U14243 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12497) );
  AOI22_X1 U14244 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12686), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12496) );
  AOI22_X1 U14245 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12629), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12495) );
  AOI22_X1 U14246 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12693), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12494) );
  AOI22_X1 U14247 ( .A1(n12685), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12518), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12501) );
  AOI22_X1 U14248 ( .A1(n12507), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12687), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12500) );
  AOI22_X1 U14249 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12499) );
  AOI22_X1 U14250 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12808), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12498) );
  AOI22_X1 U14251 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12506) );
  AOI22_X1 U14252 ( .A1(n12518), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13192), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12505) );
  AOI22_X1 U14253 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12686), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12504) );
  AOI22_X1 U14254 ( .A1(n13286), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11021), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12503) );
  AOI22_X1 U14255 ( .A1(n12685), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12687), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12511) );
  AOI22_X1 U14256 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12629), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12510) );
  AOI22_X1 U14257 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12693), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12509) );
  AOI22_X1 U14258 ( .A1(n12507), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12808), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12508) );
  NOR2_X1 U14259 ( .A1(n12562), .A2(n12561), .ZN(n14700) );
  NAND2_X1 U14260 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12517) );
  NAND2_X1 U14261 ( .A1(n12687), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12516) );
  NAND2_X1 U14262 ( .A1(n12507), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12515) );
  NAND2_X1 U14263 ( .A1(n12808), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12514) );
  NAND2_X1 U14264 ( .A1(n12685), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12522) );
  NAND2_X1 U14265 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12521) );
  NAND2_X1 U14266 ( .A1(n11017), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12520) );
  NAND2_X1 U14267 ( .A1(n12693), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12519) );
  NAND2_X1 U14268 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12525) );
  NAND2_X1 U14269 ( .A1(n12612), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12524) );
  NAND2_X1 U14270 ( .A1(n12629), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12523) );
  NAND2_X1 U14271 ( .A1(n12686), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12530) );
  NAND2_X1 U14272 ( .A1(n12527), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12529) );
  NAND2_X1 U14273 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12528) );
  NAND2_X1 U14274 ( .A1(n12507), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12539) );
  NAND2_X1 U14275 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12538) );
  NAND2_X1 U14276 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12537) );
  NAND2_X1 U14277 ( .A1(n12687), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12536) );
  NAND2_X1 U14278 ( .A1(n12685), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12542) );
  NAND2_X1 U14279 ( .A1(n12808), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12541) );
  NAND2_X1 U14280 ( .A1(n12693), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12540) );
  NAND3_X1 U14281 ( .A1(n12542), .A2(n12541), .A3(n12540), .ZN(n12543) );
  NOR2_X1 U14282 ( .A1(n11234), .A2(n12543), .ZN(n12544) );
  NAND2_X1 U14283 ( .A1(n12527), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12548) );
  NAND2_X1 U14284 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12547) );
  NAND2_X1 U14285 ( .A1(n12629), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12546) );
  NAND3_X1 U14286 ( .A1(n12548), .A2(n12547), .A3(n12546), .ZN(n12549) );
  NAND2_X1 U14287 ( .A1(n11017), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12553) );
  NAND2_X1 U14288 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12552) );
  NAND2_X1 U14289 ( .A1(n12686), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12551) );
  NAND2_X1 U14290 ( .A1(n11022), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12550) );
  XNOR2_X1 U14291 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n12881) );
  NAND2_X1 U14292 ( .A1(n15401), .A2(n12881), .ZN(n12557) );
  NAND4_X1 U14293 ( .A1(n13121), .A2(n15156), .A3(n15215), .A4(n12574), .ZN(
        n13082) );
  INV_X1 U14294 ( .A(n13082), .ZN(n12968) );
  AND2_X2 U14295 ( .A1(n12565), .A2(n14810), .ZN(n12583) );
  NAND2_X1 U14296 ( .A1(n12562), .A2(n13623), .ZN(n12560) );
  INV_X1 U14297 ( .A(n12565), .ZN(n12566) );
  NAND2_X1 U14298 ( .A1(n15869), .A2(n12566), .ZN(n12567) );
  OAI211_X2 U14299 ( .C1(n12583), .C2(n15096), .A(n12568), .B(n12567), .ZN(
        n12595) );
  INV_X1 U14300 ( .A(n12595), .ZN(n12571) );
  NAND2_X1 U14301 ( .A1(n12572), .A2(n12962), .ZN(n12573) );
  NAND2_X1 U14302 ( .A1(n12574), .A2(n13623), .ZN(n12575) );
  NAND2_X1 U14303 ( .A1(n12576), .A2(n12575), .ZN(n12600) );
  INV_X1 U14304 ( .A(n12600), .ZN(n12577) );
  NAND2_X1 U14305 ( .A1(n12577), .A2(n10997), .ZN(n12582) );
  OAI21_X1 U14306 ( .B1(n14810), .B2(n12966), .A(n12599), .ZN(n12578) );
  NAND2_X1 U14307 ( .A1(n12582), .A2(n12578), .ZN(n12954) );
  INV_X1 U14308 ( .A(n12952), .ZN(n12579) );
  NAND2_X1 U14309 ( .A1(n12579), .A2(n15178), .ZN(n12580) );
  NOR2_X2 U14310 ( .A1(n13096), .A2(n12596), .ZN(n14869) );
  NAND2_X1 U14311 ( .A1(n15228), .A2(n15401), .ZN(n12581) );
  OAI21_X1 U14312 ( .B1(n12595), .B2(n12581), .A(n12966), .ZN(n12584) );
  NAND3_X1 U14313 ( .A1(n14869), .A2(n12584), .A3(n12608), .ZN(n12585) );
  NAND2_X1 U14314 ( .A1(n12585), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12586) );
  NAND2_X1 U14315 ( .A1(n12673), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12589) );
  XNOR2_X1 U14316 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21978) );
  OR2_X1 U14317 ( .A1(n21800), .A2(n22066), .ZN(n12668) );
  OAI21_X1 U14318 ( .B1(n13609), .B2(n21978), .A(n12668), .ZN(n12587) );
  INV_X1 U14319 ( .A(n12587), .ZN(n12588) );
  NAND2_X1 U14320 ( .A1(n12589), .A2(n12588), .ZN(n12591) );
  INV_X1 U14321 ( .A(n12590), .ZN(n12669) );
  NAND2_X1 U14322 ( .A1(n12673), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12594) );
  INV_X1 U14323 ( .A(n21800), .ZN(n17348) );
  INV_X1 U14324 ( .A(n13609), .ZN(n12731) );
  MUX2_X1 U14325 ( .A(n17348), .B(n12731), .S(n22076), .Z(n12592) );
  INV_X1 U14326 ( .A(n12592), .ZN(n12593) );
  NAND2_X1 U14327 ( .A1(n12956), .A2(n15156), .ZN(n13095) );
  INV_X1 U14328 ( .A(n12596), .ZN(n12598) );
  NAND2_X1 U14329 ( .A1(n15215), .A2(n12558), .ZN(n12597) );
  NAND2_X1 U14330 ( .A1(n12600), .A2(n21510), .ZN(n12606) );
  NAND2_X1 U14331 ( .A1(n12966), .A2(n14745), .ZN(n15164) );
  OR2_X1 U14332 ( .A1(n21794), .A2(n21804), .ZN(n20204) );
  INV_X1 U14333 ( .A(n20204), .ZN(n12602) );
  OAI211_X1 U14334 ( .C1(n12559), .C2(n12966), .A(n15164), .B(n12602), .ZN(
        n12603) );
  INV_X1 U14335 ( .A(n12603), .ZN(n12605) );
  AND2_X1 U14336 ( .A1(n14806), .A2(n14535), .ZN(n14693) );
  OAI21_X1 U14337 ( .B1(n15096), .B2(n14810), .A(n14693), .ZN(n12604) );
  NAND2_X1 U14338 ( .A1(n12643), .A2(n12642), .ZN(n12609) );
  INV_X1 U14339 ( .A(n12609), .ZN(n12610) );
  NAND2_X1 U14340 ( .A1(n15125), .A2(n12610), .ZN(n12672) );
  AOI22_X1 U14341 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13419), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12616) );
  AOI22_X1 U14342 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12615) );
  AOI22_X1 U14343 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12614) );
  AOI22_X1 U14344 ( .A1(n13418), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12613) );
  NAND4_X1 U14345 ( .A1(n12616), .A2(n12615), .A3(n12614), .A4(n12613), .ZN(
        n12622) );
  AOI22_X1 U14346 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12620) );
  AOI22_X1 U14347 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12619) );
  INV_X1 U14348 ( .A(n12629), .ZN(n12692) );
  AOI22_X1 U14349 ( .A1(n13578), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12808), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12618) );
  BUF_X1 U14350 ( .A(n12685), .Z(n12644) );
  AOI22_X1 U14351 ( .A1(n12644), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12624), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12617) );
  NAND4_X1 U14352 ( .A1(n12620), .A2(n12619), .A3(n12618), .A4(n12617), .ZN(
        n12621) );
  OAI21_X2 U14353 ( .B1(n15382), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n12623), 
        .ZN(n12714) );
  NAND2_X1 U14354 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12639) );
  AOI22_X1 U14355 ( .A1(n12644), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12628) );
  AOI22_X1 U14356 ( .A1(n12507), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12627) );
  AOI22_X1 U14357 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12808), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12626) );
  BUF_X1 U14358 ( .A(n12693), .Z(n12624) );
  AOI22_X1 U14359 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12624), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12625) );
  NAND4_X1 U14360 ( .A1(n12628), .A2(n12627), .A3(n12626), .A4(n12625), .ZN(
        n12635) );
  AOI22_X1 U14361 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12633) );
  AOI22_X1 U14362 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13578), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12632) );
  AOI22_X1 U14363 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11022), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12631) );
  AOI22_X1 U14364 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12630) );
  NAND4_X1 U14365 ( .A1(n12633), .A2(n12632), .A3(n12631), .A4(n12630), .ZN(
        n12634) );
  OAI22_X1 U14366 ( .A1(n12684), .A2(n12841), .B1(n12683), .B2(n12636), .ZN(
        n12637) );
  INV_X1 U14367 ( .A(n12637), .ZN(n12638) );
  NAND2_X1 U14368 ( .A1(n12639), .A2(n12638), .ZN(n12640) );
  NAND2_X1 U14369 ( .A1(n12714), .A2(n12640), .ZN(n12641) );
  INV_X1 U14370 ( .A(n12684), .ZN(n12658) );
  AOI22_X1 U14371 ( .A1(n12644), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12649) );
  AOI22_X1 U14372 ( .A1(n12507), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12648) );
  AOI22_X1 U14373 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13578), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12647) );
  AOI22_X1 U14374 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12624), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12646) );
  NAND4_X1 U14375 ( .A1(n12649), .A2(n12648), .A3(n12647), .A4(n12646), .ZN(
        n12656) );
  AOI22_X1 U14376 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13192), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12654) );
  AOI22_X1 U14377 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11022), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12653) );
  AOI22_X1 U14378 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12652) );
  AOI22_X1 U14379 ( .A1(n13584), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12808), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12651) );
  NAND4_X1 U14380 ( .A1(n12654), .A2(n12653), .A3(n12652), .A4(n12651), .ZN(
        n12655) );
  XNOR2_X1 U14381 ( .A(n12665), .B(n12715), .ZN(n12657) );
  NAND2_X1 U14382 ( .A1(n12658), .A2(n12657), .ZN(n12659) );
  NAND2_X2 U14383 ( .A1(n12660), .A2(n12659), .ZN(n12710) );
  NAND2_X1 U14384 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12664) );
  INV_X1 U14385 ( .A(n12715), .ZN(n12661) );
  NAND2_X1 U14386 ( .A1(n12661), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12662) );
  AOI22_X1 U14387 ( .A1(n12913), .A2(n12662), .B1(n15411), .B2(n12841), .ZN(
        n12663) );
  NAND2_X1 U14388 ( .A1(n12664), .A2(n12663), .ZN(n12709) );
  NAND2_X1 U14389 ( .A1(n12710), .A2(n12709), .ZN(n12666) );
  INV_X1 U14390 ( .A(n12668), .ZN(n12670) );
  OAI21_X1 U14391 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n12670), .A(
        n12669), .ZN(n12671) );
  NAND2_X1 U14392 ( .A1(n12673), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12679) );
  NAND2_X1 U14393 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n12674) );
  NAND2_X1 U14394 ( .A1(n22039), .A2(n12674), .ZN(n12676) );
  NAND2_X1 U14395 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n22104) );
  INV_X1 U14396 ( .A(n22104), .ZN(n12675) );
  NAND2_X1 U14397 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12675), .ZN(
        n12729) );
  NAND2_X1 U14398 ( .A1(n12676), .A2(n12729), .ZN(n15809) );
  OAI22_X1 U14399 ( .A1(n13609), .A2(n15809), .B1(n21800), .B2(n22039), .ZN(
        n12677) );
  INV_X1 U14400 ( .A(n12677), .ZN(n12678) );
  AOI22_X1 U14401 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11016), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12691) );
  AOI22_X1 U14402 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12644), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12690) );
  AOI22_X1 U14403 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12689) );
  AOI22_X1 U14404 ( .A1(n13564), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12688) );
  NAND4_X1 U14405 ( .A1(n12691), .A2(n12690), .A3(n12689), .A4(n12688), .ZN(
        n12699) );
  INV_X2 U14406 ( .A(n12692), .ZN(n13578) );
  AOI22_X1 U14407 ( .A1(n13418), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13578), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12697) );
  AOI22_X1 U14408 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12624), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12696) );
  AOI22_X1 U14409 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12695) );
  AOI22_X1 U14410 ( .A1(n11022), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12808), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12694) );
  NAND4_X1 U14411 ( .A1(n12697), .A2(n12696), .A3(n12695), .A4(n12694), .ZN(
        n12698) );
  AOI22_X1 U14412 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12943), .B2(n12703), .ZN(n12700) );
  NAND2_X1 U14413 ( .A1(n12753), .A2(n11243), .ZN(n13126) );
  INV_X1 U14414 ( .A(n12904), .ZN(n12837) );
  INV_X1 U14415 ( .A(n12703), .ZN(n12705) );
  NAND2_X1 U14416 ( .A1(n12716), .A2(n12715), .ZN(n12704) );
  NAND2_X1 U14417 ( .A1(n12704), .A2(n12705), .ZN(n12746) );
  OAI21_X1 U14418 ( .B1(n12705), .B2(n12704), .A(n12746), .ZN(n12707) );
  NAND2_X1 U14419 ( .A1(n12966), .A2(n12971), .ZN(n12711) );
  INV_X1 U14420 ( .A(n12711), .ZN(n12706) );
  AOI21_X1 U14421 ( .B1(n12707), .B2(n21510), .A(n12706), .ZN(n12708) );
  OAI21_X1 U14422 ( .B1(n13126), .B2(n12837), .A(n12708), .ZN(n14896) );
  XNOR2_X2 U14423 ( .A(n12710), .B(n12709), .ZN(n13134) );
  OAI21_X1 U14424 ( .B1(n12599), .B2(n12715), .A(n12711), .ZN(n12712) );
  INV_X1 U14425 ( .A(n12712), .ZN(n12713) );
  OAI21_X2 U14426 ( .B1(n13134), .B2(n12837), .A(n12713), .ZN(n14773) );
  NAND2_X2 U14427 ( .A1(n14773), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14772) );
  OR2_X1 U14428 ( .A1(n12714), .A2(n12837), .ZN(n12720) );
  XNOR2_X1 U14429 ( .A(n12716), .B(n12715), .ZN(n12717) );
  OAI211_X1 U14430 ( .C1(n12717), .C2(n12599), .A(n12559), .B(n12562), .ZN(
        n12718) );
  INV_X1 U14431 ( .A(n12718), .ZN(n12719) );
  INV_X1 U14432 ( .A(n12721), .ZN(n12722) );
  OR2_X1 U14433 ( .A1(n12722), .A2(n14772), .ZN(n12723) );
  INV_X1 U14434 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12725) );
  NAND2_X1 U14435 ( .A1(n12726), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12727) );
  INV_X1 U14436 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12728) );
  NAND2_X1 U14437 ( .A1(n12673), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12733) );
  INV_X1 U14438 ( .A(n12729), .ZN(n22099) );
  NAND2_X1 U14439 ( .A1(n22099), .A2(n22105), .ZN(n15421) );
  NAND2_X1 U14440 ( .A1(n12729), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12730) );
  NAND2_X1 U14441 ( .A1(n15421), .A2(n12730), .ZN(n22016) );
  AOI22_X1 U14442 ( .A1(n12731), .A2(n22016), .B1(n17348), .B2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12732) );
  AOI22_X1 U14443 ( .A1(n12644), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12737) );
  AOI22_X1 U14444 ( .A1(n13418), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12736) );
  INV_X1 U14445 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13500) );
  AOI22_X1 U14446 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12808), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12735) );
  AOI22_X1 U14447 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12624), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12734) );
  NAND4_X1 U14448 ( .A1(n12737), .A2(n12736), .A3(n12735), .A4(n12734), .ZN(
        n12743) );
  AOI22_X1 U14449 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12741) );
  AOI22_X1 U14450 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13578), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12740) );
  AOI22_X1 U14451 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12739) );
  AOI22_X1 U14452 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12738) );
  NAND4_X1 U14453 ( .A1(n12741), .A2(n12740), .A3(n12739), .A4(n12738), .ZN(
        n12742) );
  AOI22_X1 U14454 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12943), .B2(n12747), .ZN(n12744) );
  NAND2_X1 U14455 ( .A1(n13146), .A2(n12904), .ZN(n12749) );
  NAND2_X1 U14456 ( .A1(n12746), .A2(n12747), .ZN(n12796) );
  OAI211_X1 U14457 ( .C1(n12747), .C2(n12746), .A(n12796), .B(n21510), .ZN(
        n12748) );
  NAND2_X1 U14458 ( .A1(n12749), .A2(n12748), .ZN(n14923) );
  NAND2_X1 U14459 ( .A1(n12750), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12751) );
  NAND2_X1 U14460 ( .A1(n12752), .A2(n12751), .ZN(n15139) );
  INV_X1 U14461 ( .A(n12753), .ZN(n12754) );
  NAND2_X1 U14462 ( .A1(n12754), .A2(n21955), .ZN(n12768) );
  INV_X1 U14463 ( .A(n12768), .ZN(n12766) );
  AOI22_X1 U14464 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n12644), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12758) );
  AOI22_X1 U14465 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n13192), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12757) );
  AOI22_X1 U14466 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12650), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12756) );
  AOI22_X1 U14467 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n13419), .B1(
        n12624), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12755) );
  NAND4_X1 U14468 ( .A1(n12758), .A2(n12757), .A3(n12756), .A4(n12755), .ZN(
        n12764) );
  AOI22_X1 U14469 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12762) );
  AOI22_X1 U14470 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13578), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12761) );
  AOI22_X1 U14471 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12760) );
  AOI22_X1 U14472 ( .A1(n13418), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12808), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12759) );
  NAND4_X1 U14473 ( .A1(n12762), .A2(n12761), .A3(n12760), .A4(n12759), .ZN(
        n12763) );
  AOI22_X1 U14474 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12943), .B2(n12794), .ZN(n12767) );
  NAND2_X1 U14475 ( .A1(n12768), .A2(n12767), .ZN(n12769) );
  AND2_X1 U14476 ( .A1(n12792), .A2(n12769), .ZN(n13161) );
  NAND2_X1 U14477 ( .A1(n13161), .A2(n12904), .ZN(n12772) );
  XNOR2_X1 U14478 ( .A(n12796), .B(n12794), .ZN(n12770) );
  NAND2_X1 U14479 ( .A1(n12770), .A2(n21510), .ZN(n12771) );
  NAND2_X1 U14480 ( .A1(n12772), .A2(n12771), .ZN(n12774) );
  INV_X1 U14481 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12773) );
  XNOR2_X1 U14482 ( .A(n12774), .B(n12773), .ZN(n15140) );
  NAND2_X1 U14483 ( .A1(n15139), .A2(n15140), .ZN(n12776) );
  NAND2_X1 U14484 ( .A1(n12774), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12775) );
  NAND2_X1 U14485 ( .A1(n12776), .A2(n12775), .ZN(n20145) );
  INV_X1 U14486 ( .A(n12792), .ZN(n12789) );
  NAND2_X1 U14487 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12788) );
  AOI22_X1 U14488 ( .A1(n12644), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12780) );
  AOI22_X1 U14489 ( .A1(n13418), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12779) );
  AOI22_X1 U14490 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13526), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12778) );
  AOI22_X1 U14491 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12624), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12777) );
  NAND4_X1 U14492 ( .A1(n12780), .A2(n12779), .A3(n12778), .A4(n12777), .ZN(
        n12786) );
  AOI22_X1 U14493 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12784) );
  AOI22_X1 U14494 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13578), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12783) );
  AOI22_X1 U14495 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12782) );
  AOI22_X1 U14496 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12781) );
  NAND4_X1 U14497 ( .A1(n12784), .A2(n12783), .A3(n12782), .A4(n12781), .ZN(
        n12785) );
  NAND2_X1 U14498 ( .A1(n12943), .A2(n12797), .ZN(n12787) );
  NAND2_X1 U14499 ( .A1(n12788), .A2(n12787), .ZN(n12790) );
  INV_X1 U14500 ( .A(n12790), .ZN(n12791) );
  NAND2_X1 U14501 ( .A1(n12792), .A2(n12791), .ZN(n12793) );
  NAND2_X1 U14502 ( .A1(n12818), .A2(n12793), .ZN(n13162) );
  OR2_X1 U14503 ( .A1(n13162), .A2(n12837), .ZN(n12800) );
  INV_X1 U14504 ( .A(n12794), .ZN(n12795) );
  NOR2_X1 U14505 ( .A1(n12796), .A2(n12795), .ZN(n12798) );
  NAND2_X1 U14506 ( .A1(n12798), .A2(n12797), .ZN(n12828) );
  OAI211_X1 U14507 ( .C1(n12798), .C2(n12797), .A(n12828), .B(n21510), .ZN(
        n12799) );
  NAND2_X1 U14508 ( .A1(n12800), .A2(n12799), .ZN(n12801) );
  INV_X1 U14509 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21552) );
  XNOR2_X1 U14510 ( .A(n12801), .B(n21552), .ZN(n20146) );
  NAND2_X1 U14511 ( .A1(n20145), .A2(n20146), .ZN(n12803) );
  NAND2_X1 U14512 ( .A1(n12801), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12802) );
  NAND2_X1 U14513 ( .A1(n12803), .A2(n12802), .ZN(n15490) );
  INV_X1 U14514 ( .A(n12818), .ZN(n12816) );
  AOI22_X1 U14515 ( .A1(n13564), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13192), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12807) );
  AOI22_X1 U14516 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12806) );
  AOI22_X1 U14517 ( .A1(n13418), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12805) );
  AOI22_X1 U14518 ( .A1(n12644), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12624), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12804) );
  NAND4_X1 U14519 ( .A1(n12807), .A2(n12806), .A3(n12805), .A4(n12804), .ZN(
        n12814) );
  AOI22_X1 U14520 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11016), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12812) );
  AOI22_X1 U14521 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12811) );
  AOI22_X1 U14522 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12810) );
  AOI22_X1 U14523 ( .A1(n13578), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12808), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12809) );
  NAND4_X1 U14524 ( .A1(n12812), .A2(n12811), .A3(n12810), .A4(n12809), .ZN(
        n12813) );
  AOI22_X1 U14525 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12943), .B2(n12829), .ZN(n12817) );
  NAND2_X1 U14526 ( .A1(n12818), .A2(n12817), .ZN(n13178) );
  NAND3_X1 U14527 ( .A1(n12840), .A2(n13178), .A3(n12904), .ZN(n12821) );
  XNOR2_X1 U14528 ( .A(n12828), .B(n12829), .ZN(n12819) );
  NAND2_X1 U14529 ( .A1(n12819), .A2(n21510), .ZN(n12820) );
  NAND2_X1 U14530 ( .A1(n12821), .A2(n12820), .ZN(n12822) );
  INV_X1 U14531 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21541) );
  XNOR2_X1 U14532 ( .A(n12822), .B(n21541), .ZN(n15491) );
  NAND2_X1 U14533 ( .A1(n15490), .A2(n15491), .ZN(n12824) );
  NAND2_X1 U14534 ( .A1(n12822), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12823) );
  INV_X1 U14535 ( .A(n12935), .ZN(n12925) );
  INV_X1 U14536 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12826) );
  NAND2_X1 U14537 ( .A1(n12943), .A2(n12841), .ZN(n12825) );
  OAI21_X1 U14538 ( .B1(n12925), .B2(n12826), .A(n12825), .ZN(n12827) );
  NAND2_X1 U14539 ( .A1(n13186), .A2(n12904), .ZN(n12833) );
  INV_X1 U14540 ( .A(n12828), .ZN(n12830) );
  NAND2_X1 U14541 ( .A1(n12830), .A2(n12829), .ZN(n12843) );
  XNOR2_X1 U14542 ( .A(n12843), .B(n12841), .ZN(n12831) );
  NAND2_X1 U14543 ( .A1(n12831), .A2(n21510), .ZN(n12832) );
  NAND2_X1 U14544 ( .A1(n12833), .A2(n12832), .ZN(n12834) );
  INV_X1 U14545 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15591) );
  XNOR2_X1 U14546 ( .A(n12834), .B(n15591), .ZN(n15557) );
  NAND2_X1 U14547 ( .A1(n15556), .A2(n15557), .ZN(n12836) );
  NAND2_X1 U14548 ( .A1(n12834), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12835) );
  NOR2_X1 U14549 ( .A1(n12838), .A2(n12837), .ZN(n12839) );
  NAND2_X1 U14550 ( .A1(n21510), .A2(n12841), .ZN(n12842) );
  OR2_X1 U14551 ( .A1(n12843), .A2(n12842), .ZN(n12844) );
  NAND2_X1 U14552 ( .A1(n12850), .A2(n12844), .ZN(n12845) );
  XNOR2_X1 U14553 ( .A(n12845), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15584) );
  INV_X1 U14554 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16569) );
  XNOR2_X1 U14555 ( .A(n12850), .B(n16569), .ZN(n15613) );
  NAND2_X1 U14556 ( .A1(n12848), .A2(n12847), .ZN(n15612) );
  NAND2_X1 U14557 ( .A1(n16382), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12849) );
  NAND2_X1 U14558 ( .A1(n16382), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15891) );
  INV_X1 U14559 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21521) );
  NAND2_X1 U14560 ( .A1(n12850), .A2(n21521), .ZN(n12851) );
  NAND2_X1 U14561 ( .A1(n15891), .A2(n12851), .ZN(n16395) );
  INV_X1 U14562 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16551) );
  NAND2_X1 U14563 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12852) );
  INV_X1 U14564 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21565) );
  NAND2_X1 U14565 ( .A1(n16382), .A2(n21565), .ZN(n16501) );
  AND2_X1 U14566 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n21555) );
  NAND2_X1 U14567 ( .A1(n21555), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13084) );
  OAI21_X1 U14568 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(n16382), .ZN(n12856) );
  NOR2_X1 U14569 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16391) );
  NAND2_X1 U14570 ( .A1(n16391), .A2(n16551), .ZN(n12855) );
  NAND2_X1 U14571 ( .A1(n16382), .A2(n12855), .ZN(n15888) );
  NAND2_X1 U14572 ( .A1(n12856), .A2(n15888), .ZN(n16381) );
  INV_X1 U14573 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16522) );
  NAND2_X1 U14574 ( .A1(n16522), .A2(n21565), .ZN(n21556) );
  NOR2_X1 U14575 ( .A1(n21556), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12857) );
  NOR2_X1 U14576 ( .A1(n12866), .A2(n12857), .ZN(n12858) );
  NOR2_X1 U14577 ( .A1(n16381), .A2(n12858), .ZN(n12859) );
  NAND4_X1 U14578 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16458) );
  INV_X1 U14579 ( .A(n16458), .ZN(n12860) );
  INV_X1 U14580 ( .A(n16366), .ZN(n12861) );
  INV_X1 U14581 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16484) );
  INV_X1 U14582 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16367) );
  INV_X1 U14583 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16456) );
  INV_X1 U14584 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n20183) );
  NAND2_X1 U14585 ( .A1(n12861), .A2(n11235), .ZN(n12862) );
  NAND2_X1 U14586 ( .A1(n12862), .A2(n16382), .ZN(n16358) );
  AND2_X1 U14587 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n13107) );
  NAND2_X1 U14588 ( .A1(n13107), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13691) );
  NAND2_X1 U14589 ( .A1(n10999), .A2(n13691), .ZN(n12863) );
  NAND2_X1 U14590 ( .A1(n12863), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12864) );
  INV_X1 U14591 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21603) );
  INV_X1 U14592 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n13057) );
  INV_X1 U14593 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16433) );
  NAND3_X1 U14594 ( .A1(n21603), .A2(n13057), .A3(n16433), .ZN(n13690) );
  NAND2_X1 U14595 ( .A1(n12865), .A2(n12866), .ZN(n16343) );
  NAND2_X1 U14596 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16424) );
  NAND2_X1 U14597 ( .A1(n20182), .A2(n16424), .ZN(n12868) );
  INV_X1 U14598 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21580) );
  INV_X1 U14599 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13696) );
  NAND2_X1 U14600 ( .A1(n21580), .A2(n13696), .ZN(n16425) );
  INV_X1 U14601 ( .A(n16425), .ZN(n12867) );
  NOR2_X1 U14602 ( .A1(n16382), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16319) );
  INV_X1 U14603 ( .A(n12877), .ZN(n12872) );
  XNOR2_X1 U14604 ( .A(n12866), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12876) );
  INV_X1 U14605 ( .A(n12876), .ZN(n12871) );
  NOR2_X1 U14606 ( .A1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12869) );
  OR2_X1 U14607 ( .A1(n12866), .A2(n12869), .ZN(n12870) );
  NAND2_X1 U14608 ( .A1(n12872), .A2(n11236), .ZN(n12880) );
  INV_X1 U14609 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16419) );
  NOR2_X1 U14610 ( .A1(n20182), .A2(n16419), .ZN(n16318) );
  INV_X1 U14611 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16310) );
  NAND2_X1 U14612 ( .A1(n12866), .A2(n16310), .ZN(n12875) );
  INV_X1 U14613 ( .A(n12875), .ZN(n12873) );
  AOI211_X1 U14614 ( .C1(n16382), .C2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n16318), .B(n12873), .ZN(n12874) );
  OR2_X1 U14615 ( .A1(n12874), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12879) );
  NAND3_X1 U14616 ( .A1(n12877), .A2(n12876), .A3(n12875), .ZN(n12878) );
  INV_X1 U14617 ( .A(n12881), .ZN(n12882) );
  NAND2_X1 U14618 ( .A1(n12882), .A2(n21847), .ZN(n21842) );
  INV_X1 U14619 ( .A(n21842), .ZN(n17347) );
  NAND2_X1 U14620 ( .A1(n22066), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12885) );
  NAND2_X1 U14621 ( .A1(n12883), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12884) );
  NAND2_X1 U14622 ( .A1(n12885), .A2(n12884), .ZN(n12894) );
  NAND2_X1 U14623 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n22076), .ZN(
        n12911) );
  NAND2_X1 U14624 ( .A1(n12896), .A2(n12885), .ZN(n12900) );
  NAND2_X1 U14625 ( .A1(n22039), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12887) );
  NAND2_X1 U14626 ( .A1(n12445), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12886) );
  NAND2_X1 U14627 ( .A1(n12900), .A2(n12901), .ZN(n12888) );
  NOR2_X1 U14628 ( .A1(n11209), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12889) );
  INV_X1 U14629 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17385) );
  NAND2_X1 U14630 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17385), .ZN(
        n12891) );
  NAND2_X1 U14631 ( .A1(n12897), .A2(n12891), .ZN(n12893) );
  NAND2_X1 U14632 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n14894), .ZN(
        n12892) );
  NAND2_X1 U14633 ( .A1(n12894), .A2(n12911), .ZN(n12895) );
  NAND3_X1 U14634 ( .A1(n12897), .A2(n14894), .A3(
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n12931) );
  XNOR2_X1 U14635 ( .A(n11209), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12898) );
  XNOR2_X1 U14636 ( .A(n12899), .B(n12898), .ZN(n12937) );
  XOR2_X1 U14637 ( .A(n12901), .B(n12900), .Z(n12924) );
  AND2_X1 U14638 ( .A1(n12934), .A2(n12924), .ZN(n12902) );
  NAND2_X1 U14639 ( .A1(n12908), .A2(n12902), .ZN(n12903) );
  NAND2_X1 U14640 ( .A1(n12942), .A2(n12903), .ZN(n14705) );
  NAND2_X1 U14641 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21834) );
  INV_X1 U14642 ( .A(n21834), .ZN(n21841) );
  NOR2_X1 U14643 ( .A1(n14705), .A2(n21841), .ZN(n14802) );
  OAI21_X1 U14644 ( .B1(n15401), .B2(n17347), .A(n14802), .ZN(n12951) );
  NAND2_X1 U14645 ( .A1(n12574), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12907) );
  INV_X1 U14646 ( .A(n12907), .ZN(n12905) );
  NOR3_X1 U14647 ( .A1(n12943), .A2(n12905), .A3(n15401), .ZN(n12906) );
  INV_X1 U14648 ( .A(n12906), .ZN(n12932) );
  NOR2_X1 U14649 ( .A1(n12906), .A2(n12908), .ZN(n12923) );
  OAI21_X1 U14650 ( .B1(n12925), .B2(n12908), .A(n12907), .ZN(n12909) );
  AOI21_X1 U14651 ( .B1(n12943), .B2(n14745), .A(n12909), .ZN(n12922) );
  NOR3_X1 U14652 ( .A1(n12909), .A2(n12908), .A3(n14745), .ZN(n12921) );
  NAND2_X1 U14653 ( .A1(n15401), .A2(n12562), .ZN(n12910) );
  INV_X1 U14654 ( .A(n12569), .ZN(n12914) );
  INV_X1 U14655 ( .A(n12911), .ZN(n12912) );
  AOI21_X1 U14656 ( .B1(n12447), .B2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n12912), .ZN(n12915) );
  INV_X1 U14657 ( .A(n12943), .ZN(n12917) );
  INV_X1 U14658 ( .A(n12915), .ZN(n12916) );
  OAI21_X1 U14659 ( .B1(n12917), .B2(n12916), .A(n12939), .ZN(n12918) );
  OAI21_X1 U14660 ( .B1(n12927), .B2(n12919), .A(n12918), .ZN(n12920) );
  OAI22_X1 U14661 ( .A1(n12923), .A2(n12922), .B1(n12921), .B2(n12920), .ZN(
        n12926) );
  OAI211_X1 U14662 ( .C1(n12926), .C2(n12927), .A(n12943), .B(n12924), .ZN(
        n12930) );
  NOR2_X1 U14663 ( .A1(n12925), .A2(n12924), .ZN(n12928) );
  OAI21_X1 U14664 ( .B1(n12928), .B2(n12927), .A(n12926), .ZN(n12929) );
  OAI211_X1 U14665 ( .C1(n12932), .C2(n12931), .A(n12930), .B(n12929), .ZN(
        n12933) );
  OAI21_X1 U14666 ( .B1(n12935), .B2(n12934), .A(n12933), .ZN(n12936) );
  OAI21_X1 U14667 ( .B1(n12939), .B2(n12937), .A(n12936), .ZN(n12938) );
  AOI21_X1 U14668 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n21804), .A(
        n12938), .ZN(n12941) );
  INV_X1 U14669 ( .A(n12942), .ZN(n12944) );
  NAND2_X1 U14670 ( .A1(n12944), .A2(n12943), .ZN(n12945) );
  AND2_X4 U14671 ( .A1(n12946), .A2(n12945), .ZN(n15175) );
  NAND2_X1 U14672 ( .A1(n15401), .A2(n21842), .ZN(n13643) );
  NAND3_X1 U14673 ( .A1(n12947), .A2(n21834), .A3(n13643), .ZN(n12948) );
  NAND3_X1 U14674 ( .A1(n12948), .A2(n15178), .A3(n15869), .ZN(n12949) );
  NAND2_X1 U14675 ( .A1(n15175), .A2(n12949), .ZN(n12950) );
  MUX2_X1 U14676 ( .A(n12951), .B(n12950), .S(n12559), .Z(n12961) );
  NAND2_X1 U14677 ( .A1(n12583), .A2(n14745), .ZN(n12958) );
  NAND2_X1 U14678 ( .A1(n12952), .A2(n12583), .ZN(n12964) );
  NAND3_X1 U14679 ( .A1(n15178), .A2(n12559), .A3(n12971), .ZN(n14702) );
  NAND2_X1 U14680 ( .A1(n14810), .A2(n15411), .ZN(n12953) );
  NAND2_X1 U14681 ( .A1(n12953), .A2(n14811), .ZN(n13092) );
  AOI21_X1 U14682 ( .B1(n12964), .B2(n14702), .A(n13092), .ZN(n12963) );
  AND2_X1 U14683 ( .A1(n12954), .A2(n12963), .ZN(n12957) );
  NAND2_X1 U14684 ( .A1(n12569), .A2(n12966), .ZN(n12955) );
  OR2_X1 U14685 ( .A1(n12957), .A2(n14803), .ZN(n14858) );
  OAI21_X1 U14686 ( .B1(n15175), .B2(n12958), .A(n14858), .ZN(n12959) );
  INV_X1 U14687 ( .A(n12959), .ZN(n12960) );
  NAND2_X1 U14688 ( .A1(n21800), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n21813) );
  AND2_X1 U14689 ( .A1(n12963), .A2(n12569), .ZN(n13120) );
  OR2_X1 U14690 ( .A1(n12964), .A2(n14806), .ZN(n15217) );
  INV_X1 U14691 ( .A(n15217), .ZN(n12965) );
  NOR2_X1 U14692 ( .A1(n13120), .A2(n12965), .ZN(n14704) );
  OR2_X2 U14693 ( .A1(n12967), .A2(n12966), .ZN(n12973) );
  NAND2_X1 U14694 ( .A1(n12947), .A2(n14886), .ZN(n14800) );
  NAND2_X1 U14695 ( .A1(n12968), .A2(n12561), .ZN(n12969) );
  NAND4_X1 U14696 ( .A1(n10996), .A2(n14704), .A3(n14800), .A4(n12969), .ZN(
        n12970) );
  OR2_X1 U14697 ( .A1(n12971), .A2(n12966), .ZN(n12979) );
  MUX2_X1 U14698 ( .A(n13071), .B(n12979), .S(P1_EBX_REG_1__SCAN_IN), .Z(
        n12976) );
  INV_X1 U14699 ( .A(n12979), .ZN(n12972) );
  NAND2_X1 U14700 ( .A1(n11020), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12974) );
  AND2_X1 U14701 ( .A1(n13052), .A2(n12974), .ZN(n12975) );
  NAND2_X1 U14702 ( .A1(n12979), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12977) );
  OAI21_X1 U14703 ( .B1(n13074), .B2(P1_EBX_REG_0__SCAN_IN), .A(n12977), .ZN(
        n14776) );
  XNOR2_X1 U14704 ( .A(n12978), .B(n14776), .ZN(n14887) );
  NAND2_X1 U14705 ( .A1(n14887), .A2(n14886), .ZN(n14885) );
  NAND2_X1 U14706 ( .A1(n14885), .A2(n12978), .ZN(n14899) );
  MUX2_X1 U14707 ( .A(n13071), .B(n13070), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n12982) );
  NAND2_X1 U14708 ( .A1(n11020), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12980) );
  AND2_X1 U14709 ( .A1(n13052), .A2(n12980), .ZN(n12981) );
  INV_X1 U14710 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n20122) );
  NAND2_X1 U14711 ( .A1(n13066), .A2(n20122), .ZN(n12985) );
  NAND2_X1 U14712 ( .A1(n14535), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12983) );
  OAI211_X1 U14713 ( .C1(n11020), .C2(P1_EBX_REG_3__SCAN_IN), .A(n12983), .B(
        n13070), .ZN(n12984) );
  AND2_X1 U14714 ( .A1(n12985), .A2(n12984), .ZN(n14930) );
  MUX2_X1 U14715 ( .A(n13071), .B(n13070), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n12988) );
  NAND2_X1 U14716 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n11020), .ZN(
        n12986) );
  AND2_X1 U14717 ( .A1(n13052), .A2(n12986), .ZN(n12987) );
  INV_X1 U14718 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20136) );
  NAND2_X1 U14719 ( .A1(n13066), .A2(n20136), .ZN(n12993) );
  NAND2_X1 U14720 ( .A1(n14535), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12991) );
  OAI211_X1 U14721 ( .C1(n11020), .C2(P1_EBX_REG_5__SCAN_IN), .A(n12991), .B(
        n13070), .ZN(n12992) );
  NAND2_X1 U14722 ( .A1(n12993), .A2(n12992), .ZN(n20131) );
  MUX2_X1 U14723 ( .A(n13071), .B(n13070), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n12996) );
  NAND2_X1 U14724 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n11020), .ZN(
        n12994) );
  AND2_X1 U14725 ( .A1(n13052), .A2(n12994), .ZN(n12995) );
  NAND2_X1 U14726 ( .A1(n12996), .A2(n12995), .ZN(n15507) );
  MUX2_X1 U14727 ( .A(n13066), .B(n13074), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n12998) );
  NOR2_X1 U14728 ( .A1(n14777), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12997) );
  NOR2_X1 U14729 ( .A1(n12998), .A2(n12997), .ZN(n15506) );
  AND2_X1 U14730 ( .A1(n15507), .A2(n15506), .ZN(n12999) );
  NAND2_X1 U14731 ( .A1(n13066), .A2(n21676), .ZN(n13002) );
  NAND2_X1 U14732 ( .A1(n14535), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13000) );
  OAI211_X1 U14733 ( .C1(n11020), .C2(P1_EBX_REG_9__SCAN_IN), .A(n13000), .B(
        n13070), .ZN(n13001) );
  AND2_X1 U14734 ( .A1(n13002), .A2(n13001), .ZN(n15622) );
  INV_X1 U14735 ( .A(n13071), .ZN(n13075) );
  INV_X1 U14736 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n20130) );
  NAND2_X1 U14737 ( .A1(n13075), .A2(n20130), .ZN(n13006) );
  INV_X1 U14738 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n13003) );
  NAND2_X1 U14739 ( .A1(n13070), .A2(n13003), .ZN(n13004) );
  OAI211_X1 U14740 ( .C1(n11020), .C2(P1_EBX_REG_8__SCAN_IN), .A(n13004), .B(
        n14535), .ZN(n13005) );
  NAND2_X1 U14741 ( .A1(n13006), .A2(n13005), .ZN(n15623) );
  MUX2_X1 U14742 ( .A(n13066), .B(n13074), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n13008) );
  INV_X1 U14743 ( .A(n13008), .ZN(n13010) );
  INV_X1 U14744 ( .A(n14777), .ZN(n13048) );
  INV_X1 U14745 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16560) );
  NAND2_X1 U14746 ( .A1(n13048), .A2(n16560), .ZN(n13009) );
  NAND2_X1 U14747 ( .A1(n13010), .A2(n13009), .ZN(n15792) );
  MUX2_X1 U14748 ( .A(n13071), .B(n13070), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n13013) );
  NAND2_X1 U14749 ( .A1(n11020), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13011) );
  AND2_X1 U14750 ( .A1(n13052), .A2(n13011), .ZN(n13012) );
  NAND2_X1 U14751 ( .A1(n13013), .A2(n13012), .ZN(n15662) );
  INV_X1 U14752 ( .A(n15662), .ZN(n15793) );
  MUX2_X1 U14753 ( .A(n13066), .B(n13074), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n13017) );
  NOR2_X1 U14754 ( .A1(n14777), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13016) );
  NOR2_X1 U14755 ( .A1(n13017), .A2(n13016), .ZN(n15909) );
  MUX2_X1 U14756 ( .A(n13071), .B(n13070), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n13020) );
  NAND2_X1 U14757 ( .A1(n11020), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13018) );
  AND2_X1 U14758 ( .A1(n13052), .A2(n13018), .ZN(n13019) );
  NAND2_X1 U14759 ( .A1(n13020), .A2(n13019), .ZN(n15924) );
  NAND2_X1 U14760 ( .A1(n15909), .A2(n15924), .ZN(n13021) );
  INV_X1 U14761 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n21719) );
  NAND2_X1 U14762 ( .A1(n13066), .A2(n21719), .ZN(n13024) );
  NAND2_X1 U14763 ( .A1(n14535), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13022) );
  OAI211_X1 U14764 ( .C1(n11020), .C2(P1_EBX_REG_15__SCAN_IN), .A(n13022), .B(
        n13070), .ZN(n13023) );
  AND2_X1 U14765 ( .A1(n13024), .A2(n13023), .ZN(n16518) );
  INV_X1 U14766 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n15839) );
  NAND2_X1 U14767 ( .A1(n13075), .A2(n15839), .ZN(n13028) );
  INV_X1 U14768 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n13025) );
  NAND2_X1 U14769 ( .A1(n13070), .A2(n13025), .ZN(n13026) );
  OAI211_X1 U14770 ( .C1(n11020), .C2(P1_EBX_REG_14__SCAN_IN), .A(n13026), .B(
        n14535), .ZN(n13027) );
  NAND2_X1 U14771 ( .A1(n13028), .A2(n13027), .ZN(n15836) );
  AND2_X1 U14772 ( .A1(n16518), .A2(n15836), .ZN(n13029) );
  MUX2_X1 U14773 ( .A(n13071), .B(n13070), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n13032) );
  NAND2_X1 U14774 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n11020), .ZN(
        n13030) );
  AND2_X1 U14775 ( .A1(n13052), .A2(n13030), .ZN(n13031) );
  NAND2_X1 U14776 ( .A1(n13032), .A2(n13031), .ZN(n15885) );
  INV_X1 U14777 ( .A(n15885), .ZN(n13033) );
  INV_X1 U14778 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n20125) );
  NAND2_X1 U14779 ( .A1(n13066), .A2(n20125), .ZN(n13037) );
  INV_X1 U14780 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n13035) );
  NAND2_X1 U14781 ( .A1(n14886), .A2(n20125), .ZN(n13034) );
  OAI211_X1 U14782 ( .C1(n13074), .C2(n13035), .A(n13034), .B(n13070), .ZN(
        n13036) );
  NAND2_X1 U14783 ( .A1(n13037), .A2(n13036), .ZN(n16196) );
  MUX2_X1 U14784 ( .A(n13071), .B(n13070), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n13040) );
  NAND2_X1 U14785 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n11020), .ZN(
        n13038) );
  AND2_X1 U14786 ( .A1(n13052), .A2(n13038), .ZN(n13039) );
  NAND2_X1 U14787 ( .A1(n13040), .A2(n13039), .ZN(n16189) );
  AND2_X2 U14788 ( .A1(n16198), .A2(n16189), .ZN(n16239) );
  INV_X1 U14789 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n16242) );
  NAND2_X1 U14790 ( .A1(n13066), .A2(n16242), .ZN(n13043) );
  NAND2_X1 U14791 ( .A1(n14535), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13041) );
  OAI211_X1 U14792 ( .C1(n11020), .C2(P1_EBX_REG_19__SCAN_IN), .A(n13041), .B(
        n13070), .ZN(n13042) );
  MUX2_X1 U14793 ( .A(n13071), .B(n13070), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n13046) );
  NAND2_X1 U14794 ( .A1(n11020), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13044) );
  AND2_X1 U14795 ( .A1(n13052), .A2(n13044), .ZN(n13045) );
  OR2_X2 U14796 ( .A1(n16241), .A2(n16231), .ZN(n16233) );
  MUX2_X1 U14797 ( .A(n13066), .B(n13074), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n13047) );
  INV_X1 U14798 ( .A(n13047), .ZN(n13050) );
  NAND2_X1 U14799 ( .A1(n13048), .A2(n16456), .ZN(n13049) );
  NAND2_X1 U14800 ( .A1(n13050), .A2(n13049), .ZN(n16173) );
  MUX2_X1 U14801 ( .A(n13071), .B(n13070), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n13054) );
  NAND2_X1 U14802 ( .A1(n11020), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13051) );
  AND2_X1 U14803 ( .A1(n13052), .A2(n13051), .ZN(n13053) );
  MUX2_X1 U14804 ( .A(n13066), .B(n13074), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n13056) );
  NOR2_X1 U14805 ( .A1(n14777), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13055) );
  NOR2_X1 U14806 ( .A1(n13056), .A2(n13055), .ZN(n16147) );
  INV_X1 U14807 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n16220) );
  NAND2_X1 U14808 ( .A1(n13075), .A2(n16220), .ZN(n13060) );
  NAND2_X1 U14809 ( .A1(n13070), .A2(n13057), .ZN(n13058) );
  OAI211_X1 U14810 ( .C1(n11020), .C2(P1_EBX_REG_24__SCAN_IN), .A(n13058), .B(
        n14535), .ZN(n13059) );
  AND2_X1 U14811 ( .A1(n13060), .A2(n13059), .ZN(n16216) );
  OR2_X2 U14812 ( .A1(n16217), .A2(n16216), .ZN(n16219) );
  INV_X1 U14813 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n16213) );
  NAND2_X1 U14814 ( .A1(n13066), .A2(n16213), .ZN(n13063) );
  NAND2_X1 U14815 ( .A1(n14535), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13061) );
  OAI211_X1 U14816 ( .C1(P1_EBX_REG_25__SCAN_IN), .C2(n11020), .A(n13061), .B(
        n13070), .ZN(n13062) );
  NAND2_X1 U14817 ( .A1(n13063), .A2(n13062), .ZN(n16130) );
  INV_X1 U14818 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16432) );
  NAND2_X1 U14819 ( .A1(n13070), .A2(n16432), .ZN(n13064) );
  OAI211_X1 U14820 ( .C1(n11020), .C2(P1_EBX_REG_26__SCAN_IN), .A(n13064), .B(
        n14535), .ZN(n13065) );
  OAI21_X1 U14821 ( .B1(n13071), .B2(P1_EBX_REG_26__SCAN_IN), .A(n13065), .ZN(
        n16117) );
  INV_X1 U14822 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n16210) );
  NAND2_X1 U14823 ( .A1(n13066), .A2(n16210), .ZN(n13069) );
  NAND2_X1 U14824 ( .A1(n14535), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13067) );
  OAI211_X1 U14825 ( .C1(P1_EBX_REG_27__SCAN_IN), .C2(n11020), .A(n13067), .B(
        n13070), .ZN(n13068) );
  NAND2_X1 U14826 ( .A1(n13069), .A2(n13068), .ZN(n16100) );
  MUX2_X1 U14827 ( .A(n13071), .B(n13070), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n13073) );
  NAND2_X1 U14828 ( .A1(n11020), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13072) );
  AND2_X1 U14829 ( .A1(n13073), .A2(n13072), .ZN(n16087) );
  NOR2_X4 U14830 ( .A1(n16102), .A2(n16087), .ZN(n16088) );
  OAI22_X1 U14831 ( .A1(n14777), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        P1_EBX_REG_29__SCAN_IN), .B2(n11020), .ZN(n14533) );
  OR2_X1 U14832 ( .A1(n14533), .A2(n13074), .ZN(n13077) );
  INV_X1 U14833 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n16078) );
  NAND2_X1 U14834 ( .A1(n13075), .A2(n16078), .ZN(n13076) );
  NAND2_X1 U14835 ( .A1(n13077), .A2(n13076), .ZN(n13628) );
  AND2_X2 U14836 ( .A1(n16088), .A2(n13628), .ZN(n14536) );
  OR2_X1 U14837 ( .A1(n14536), .A2(n13074), .ZN(n13079) );
  OAI22_X1 U14838 ( .A1(n14777), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(n11020), .ZN(n14537) );
  OAI22_X1 U14839 ( .A1(n14777), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        P1_EBX_REG_31__SCAN_IN), .B2(n11020), .ZN(n13080) );
  XNOR2_X2 U14840 ( .A(n13081), .B(n13080), .ZN(n16208) );
  NAND2_X1 U14841 ( .A1(n14695), .A2(n15401), .ZN(n17344) );
  OAI21_X1 U14842 ( .B1(n13082), .B2(n12561), .A(n17344), .ZN(n13083) );
  NOR2_X1 U14843 ( .A1(n16208), .A2(n21560), .ZN(n13117) );
  NAND3_X1 U14844 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n13085) );
  NAND2_X1 U14845 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16512) );
  NOR2_X1 U14846 ( .A1(n13084), .A2(n16512), .ZN(n16489) );
  NAND2_X1 U14847 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16489), .ZN(
        n16455) );
  NOR3_X1 U14848 ( .A1(n10990), .A2(n13085), .A3(n16455), .ZN(n13090) );
  NOR2_X1 U14849 ( .A1(n16560), .A2(n16551), .ZN(n16454) );
  INV_X1 U14850 ( .A(n16454), .ZN(n13086) );
  NAND3_X1 U14851 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15621) );
  AOI21_X1 U14852 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14929) );
  NAND2_X1 U14853 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n15141) );
  NOR2_X1 U14854 ( .A1(n14929), .A2(n15141), .ZN(n21543) );
  NAND2_X1 U14855 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n21543), .ZN(
        n21542) );
  NOR2_X1 U14856 ( .A1(n15621), .A2(n21542), .ZN(n15620) );
  NAND3_X1 U14857 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n15620), .ZN(n16546) );
  NOR2_X1 U14858 ( .A1(n13086), .A2(n16546), .ZN(n16467) );
  NAND2_X1 U14859 ( .A1(n13090), .A2(n16467), .ZN(n13102) );
  NOR2_X1 U14860 ( .A1(n14702), .A2(n15401), .ZN(n13087) );
  NAND2_X1 U14861 ( .A1(n13087), .A2(n12583), .ZN(n15216) );
  INV_X1 U14862 ( .A(n15216), .ZN(n14862) );
  INV_X1 U14863 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n13089) );
  NAND4_X1 U14864 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21529) );
  NOR2_X1 U14865 ( .A1(n21552), .A2(n21529), .ZN(n15560) );
  INV_X1 U14866 ( .A(n15621), .ZN(n13088) );
  NAND2_X1 U14867 ( .A1(n15560), .A2(n13088), .ZN(n15617) );
  NOR3_X1 U14868 ( .A1(n16569), .A2(n13089), .A3(n15617), .ZN(n16548) );
  NAND3_X1 U14869 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n16548), .ZN(n16525) );
  INV_X1 U14870 ( .A(n16525), .ZN(n16527) );
  AND2_X1 U14871 ( .A1(n13090), .A2(n16527), .ZN(n13103) );
  AND2_X1 U14872 ( .A1(n14803), .A2(n14745), .ZN(n17352) );
  NAND2_X1 U14873 ( .A1(n13100), .A2(n17352), .ZN(n16526) );
  INV_X1 U14874 ( .A(n14811), .ZN(n15867) );
  AOI21_X1 U14875 ( .B1(n12558), .B2(n14860), .A(n15867), .ZN(n13091) );
  OAI211_X1 U14876 ( .C1(n12569), .C2(n15178), .A(n13091), .B(n15228), .ZN(
        n13093) );
  AOI21_X1 U14877 ( .B1(n13093), .B2(n14745), .A(n13092), .ZN(n13094) );
  AND2_X1 U14878 ( .A1(n13095), .A2(n13094), .ZN(n14868) );
  INV_X1 U14879 ( .A(n13096), .ZN(n13097) );
  OAI211_X1 U14880 ( .C1(n13098), .C2(n15178), .A(n14868), .B(n13097), .ZN(
        n13099) );
  NAND2_X1 U14881 ( .A1(n13100), .A2(n13099), .ZN(n16466) );
  NAND2_X1 U14882 ( .A1(n16526), .A2(n16466), .ZN(n15618) );
  NAND2_X1 U14883 ( .A1(n13103), .A2(n21533), .ZN(n16442) );
  OAI21_X1 U14884 ( .B1(n13102), .B2(n16453), .A(n16442), .ZN(n21602) );
  NAND2_X1 U14885 ( .A1(n21602), .A2(n13107), .ZN(n21592) );
  NAND2_X1 U14886 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16435) );
  NOR2_X1 U14887 ( .A1(n21592), .A2(n16435), .ZN(n21581) );
  NOR2_X1 U14888 ( .A1(n16424), .A2(n16419), .ZN(n16303) );
  NAND2_X1 U14889 ( .A1(n21581), .A2(n16303), .ZN(n16410) );
  NOR2_X1 U14890 ( .A1(n16466), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13101) );
  NOR2_X1 U14891 ( .A1(n13609), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16504) );
  NOR2_X1 U14892 ( .A1(n13100), .A2(n21585), .ZN(n16529) );
  OAI21_X1 U14893 ( .B1(n21603), .B2(n13102), .A(n21544), .ZN(n13106) );
  INV_X1 U14894 ( .A(n13103), .ZN(n13104) );
  NAND2_X1 U14895 ( .A1(n15618), .A2(n13104), .ZN(n13105) );
  INV_X1 U14896 ( .A(n13107), .ZN(n16342) );
  NAND2_X1 U14897 ( .A1(n15618), .A2(n16342), .ZN(n13108) );
  OAI21_X1 U14898 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n16453), .A(
        n13108), .ZN(n13109) );
  INV_X1 U14899 ( .A(n13109), .ZN(n13110) );
  NAND2_X1 U14900 ( .A1(n21598), .A2(n13110), .ZN(n21586) );
  OR2_X1 U14901 ( .A1(n21586), .A2(n16435), .ZN(n13112) );
  NAND2_X1 U14902 ( .A1(n16453), .A2(n16466), .ZN(n14775) );
  NOR2_X1 U14903 ( .A1(n15616), .A2(n16513), .ZN(n16451) );
  INV_X1 U14904 ( .A(n16451), .ZN(n13111) );
  AND2_X1 U14905 ( .A1(n13112), .A2(n13111), .ZN(n21582) );
  INV_X1 U14906 ( .A(n21582), .ZN(n16405) );
  NAND2_X1 U14907 ( .A1(n16405), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16404) );
  INV_X1 U14908 ( .A(n16513), .ZN(n16490) );
  NOR2_X1 U14909 ( .A1(n16490), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16406) );
  NOR3_X1 U14910 ( .A1(n16404), .A2(n16406), .A3(n16424), .ZN(n13113) );
  INV_X1 U14911 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16589) );
  NOR3_X1 U14912 ( .A1(n13113), .A2(n16451), .A3(n16589), .ZN(n13114) );
  INV_X1 U14913 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20091) );
  NOR2_X1 U14914 ( .A1(n21600), .A2(n20091), .ZN(n13615) );
  NAND2_X1 U14915 ( .A1(n13121), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13151) );
  XNOR2_X1 U14916 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15360) );
  INV_X2 U14917 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n22106) );
  AOI21_X1 U14918 ( .B1(n13600), .B2(n15360), .A(n13604), .ZN(n13123) );
  NOR2_X2 U14919 ( .A1(n14811), .A2(n22106), .ZN(n13165) );
  NAND2_X1 U14920 ( .A1(n13599), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n13122) );
  OAI211_X1 U14921 ( .C1(n13151), .C2(n12445), .A(n13123), .B(n13122), .ZN(
        n13124) );
  INV_X1 U14922 ( .A(n13124), .ZN(n13125) );
  NAND2_X1 U14923 ( .A1(n13604), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13145) );
  NAND2_X1 U14924 ( .A1(n13127), .A2(n13145), .ZN(n15117) );
  INV_X1 U14925 ( .A(n15117), .ZN(n13144) );
  XNOR2_X2 U14926 ( .A(n13128), .B(n13129), .ZN(n15087) );
  NAND2_X1 U14927 ( .A1(n15087), .A2(n13312), .ZN(n13133) );
  AOI22_X1 U14928 ( .A1(n13165), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n22106), .ZN(n13131) );
  INV_X1 U14929 ( .A(n13151), .ZN(n13155) );
  NAND2_X1 U14930 ( .A1(n13155), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13130) );
  AND2_X1 U14931 ( .A1(n13131), .A2(n13130), .ZN(n13132) );
  NAND2_X1 U14932 ( .A1(n13134), .A2(n12558), .ZN(n13135) );
  NAND2_X1 U14933 ( .A1(n13135), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14814) );
  NAND2_X1 U14934 ( .A1(n22106), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13139) );
  NAND2_X1 U14935 ( .A1(n13599), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n13138) );
  OAI211_X1 U14936 ( .C1(n13151), .C2(n12447), .A(n13139), .B(n13138), .ZN(
        n13140) );
  AOI21_X1 U14937 ( .B1(n13136), .B2(n13312), .A(n13140), .ZN(n14813) );
  OR2_X1 U14938 ( .A1(n14814), .A2(n14813), .ZN(n14816) );
  INV_X1 U14939 ( .A(n14813), .ZN(n13141) );
  OR2_X1 U14940 ( .A1(n13141), .A2(n13597), .ZN(n13142) );
  NAND2_X1 U14941 ( .A1(n14816), .A2(n13142), .ZN(n14908) );
  NAND2_X1 U14942 ( .A1(n14909), .A2(n14908), .ZN(n15116) );
  INV_X1 U14943 ( .A(n15116), .ZN(n13143) );
  NAND2_X1 U14944 ( .A1(n13143), .A2(n13144), .ZN(n15114) );
  NAND2_X1 U14945 ( .A1(n13146), .A2(n13312), .ZN(n13154) );
  INV_X1 U14946 ( .A(n13147), .ZN(n13148) );
  INV_X1 U14947 ( .A(n13166), .ZN(n13157) );
  OAI21_X1 U14948 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n13148), .A(
        n13157), .ZN(n15160) );
  AOI22_X1 U14949 ( .A1(n13600), .A2(n15160), .B1(n13604), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13150) );
  NAND2_X1 U14950 ( .A1(n13599), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n13149) );
  OAI211_X1 U14951 ( .C1(n13151), .C2(n11209), .A(n13150), .B(n13149), .ZN(
        n13152) );
  INV_X1 U14952 ( .A(n13152), .ZN(n13153) );
  NAND2_X1 U14953 ( .A1(n13154), .A2(n13153), .ZN(n15106) );
  NAND2_X1 U14954 ( .A1(n15107), .A2(n15106), .ZN(n15105) );
  NAND2_X1 U14955 ( .A1(n13155), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13159) );
  INV_X1 U14956 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n21616) );
  AOI21_X1 U14957 ( .B1(n21616), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13156) );
  AOI21_X1 U14958 ( .B1(n13599), .B2(P1_EAX_REG_4__SCAN_IN), .A(n13156), .ZN(
        n13158) );
  XNOR2_X1 U14959 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B(n13157), .ZN(
        n21608) );
  AOI22_X1 U14960 ( .A1(n13159), .A2(n13158), .B1(n13600), .B2(n21608), .ZN(
        n13160) );
  INV_X1 U14961 ( .A(n13162), .ZN(n13164) );
  NAND2_X1 U14962 ( .A1(n13164), .A2(n13312), .ZN(n13172) );
  INV_X1 U14963 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n13169) );
  OAI21_X1 U14964 ( .B1(n13167), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n13173), .ZN(n21635) );
  AOI22_X1 U14965 ( .A1(n21635), .A2(n13600), .B1(n13604), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13168) );
  OAI21_X1 U14966 ( .B1(n13137), .B2(n13169), .A(n13168), .ZN(n13170) );
  INV_X1 U14967 ( .A(n13170), .ZN(n13171) );
  NAND2_X1 U14968 ( .A1(n15197), .A2(n15449), .ZN(n15445) );
  INV_X1 U14969 ( .A(n15445), .ZN(n13180) );
  INV_X1 U14970 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n13176) );
  AND2_X1 U14971 ( .A1(n13173), .A2(n21643), .ZN(n13174) );
  OR2_X1 U14972 ( .A1(n13174), .A2(n13181), .ZN(n21650) );
  AOI22_X1 U14973 ( .A1(n21650), .A2(n13600), .B1(n13604), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n13175) );
  OAI21_X1 U14974 ( .B1(n13137), .B2(n13176), .A(n13175), .ZN(n13177) );
  NAND2_X1 U14975 ( .A1(n13180), .A2(n13179), .ZN(n15443) );
  INV_X1 U14976 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n13184) );
  NOR2_X1 U14977 ( .A1(n13181), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13182) );
  OR2_X1 U14978 ( .A1(n13203), .A2(n13182), .ZN(n21661) );
  AOI22_X1 U14979 ( .A1(n21661), .A2(n13600), .B1(n13604), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n13183) );
  OAI21_X1 U14980 ( .B1(n13137), .B2(n13184), .A(n13183), .ZN(n13185) );
  AOI21_X1 U14981 ( .B1(n13186), .B2(n13312), .A(n13185), .ZN(n15509) );
  AOI22_X1 U14982 ( .A1(n12644), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11016), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13191) );
  AOI22_X1 U14983 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13190) );
  AOI22_X1 U14984 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13189) );
  AOI22_X1 U14985 ( .A1(n13418), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12624), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13188) );
  NAND4_X1 U14986 ( .A1(n13191), .A2(n13190), .A3(n13189), .A4(n13188), .ZN(
        n13198) );
  AOI22_X1 U14987 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13419), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13196) );
  AOI22_X1 U14988 ( .A1(n13584), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13195) );
  AOI22_X1 U14989 ( .A1(n13578), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13194) );
  AOI22_X1 U14990 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13526), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13193) );
  NAND4_X1 U14991 ( .A1(n13196), .A2(n13195), .A3(n13194), .A4(n13193), .ZN(
        n13197) );
  OAI21_X1 U14992 ( .B1(n13198), .B2(n13197), .A(n13312), .ZN(n13202) );
  NAND2_X1 U14993 ( .A1(n13599), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n13201) );
  XNOR2_X1 U14994 ( .A(n13203), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n21663) );
  NAND2_X1 U14995 ( .A1(n21663), .A2(n13600), .ZN(n13200) );
  NAND2_X1 U14996 ( .A1(n13604), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13199) );
  XNOR2_X1 U14997 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n13218), .ZN(
        n21674) );
  AOI22_X1 U14998 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12650), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13207) );
  AOI22_X1 U14999 ( .A1(n12644), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13419), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13206) );
  AOI22_X1 U15000 ( .A1(n13585), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13526), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13205) );
  AOI22_X1 U15001 ( .A1(n13584), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12624), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13204) );
  NAND4_X1 U15002 ( .A1(n13207), .A2(n13206), .A3(n13205), .A4(n13204), .ZN(
        n13213) );
  AOI22_X1 U15003 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13418), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13211) );
  AOI22_X1 U15004 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13578), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13210) );
  AOI22_X1 U15005 ( .A1(n13564), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11022), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13209) );
  AOI22_X1 U15006 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13208) );
  NAND4_X1 U15007 ( .A1(n13211), .A2(n13210), .A3(n13209), .A4(n13208), .ZN(
        n13212) );
  OR2_X1 U15008 ( .A1(n13213), .A2(n13212), .ZN(n13214) );
  AOI22_X1 U15009 ( .A1(n13312), .A2(n13214), .B1(n13604), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n13216) );
  NAND2_X1 U15010 ( .A1(n13599), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n13215) );
  OAI211_X1 U15011 ( .C1(n21674), .C2(n13597), .A(n13216), .B(n13215), .ZN(
        n15568) );
  INV_X1 U15012 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n13219) );
  XNOR2_X1 U15013 ( .A(n13236), .B(n13219), .ZN(n20156) );
  AOI22_X1 U15014 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13418), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13223) );
  AOI22_X1 U15015 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13578), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13222) );
  AOI22_X1 U15016 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13221) );
  AOI22_X1 U15017 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13526), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13220) );
  NAND4_X1 U15018 ( .A1(n13223), .A2(n13222), .A3(n13221), .A4(n13220), .ZN(
        n13229) );
  AOI22_X1 U15019 ( .A1(n12644), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13227) );
  AOI22_X1 U15020 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13226) );
  AOI22_X1 U15021 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13225) );
  AOI22_X1 U15022 ( .A1(n13584), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12624), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13224) );
  NAND4_X1 U15023 ( .A1(n13227), .A2(n13226), .A3(n13225), .A4(n13224), .ZN(
        n13228) );
  OAI21_X1 U15024 ( .B1(n13229), .B2(n13228), .A(n13312), .ZN(n13232) );
  NAND2_X1 U15025 ( .A1(n13599), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n13231) );
  NAND2_X1 U15026 ( .A1(n13604), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13230) );
  NAND3_X1 U15027 ( .A1(n13232), .A2(n13231), .A3(n13230), .ZN(n13233) );
  AOI21_X1 U15028 ( .B1(n13600), .B2(n20156), .A(n13233), .ZN(n15660) );
  XNOR2_X1 U15029 ( .A(n13300), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15896) );
  AOI22_X1 U15030 ( .A1(n12644), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13578), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13242) );
  AOI22_X1 U15031 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11021), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13241) );
  AOI22_X1 U15032 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13240) );
  AOI22_X1 U15033 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13526), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13239) );
  NAND4_X1 U15034 ( .A1(n13242), .A2(n13241), .A3(n13240), .A4(n13239), .ZN(
        n13248) );
  AOI22_X1 U15035 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13418), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13246) );
  AOI22_X1 U15036 ( .A1(n13564), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13192), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13245) );
  AOI22_X1 U15037 ( .A1(n13584), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13244) );
  AOI22_X1 U15038 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12624), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13243) );
  NAND4_X1 U15039 ( .A1(n13246), .A2(n13245), .A3(n13244), .A4(n13243), .ZN(
        n13247) );
  OAI21_X1 U15040 ( .B1(n13248), .B2(n13247), .A(n13312), .ZN(n13251) );
  NAND2_X1 U15041 ( .A1(n13599), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n13250) );
  NAND2_X1 U15042 ( .A1(n13604), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13249) );
  NAND3_X1 U15043 ( .A1(n13251), .A2(n13250), .A3(n13249), .ZN(n13252) );
  AOI21_X1 U15044 ( .B1(n15896), .B2(n13600), .A(n13252), .ZN(n15835) );
  XNOR2_X1 U15045 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n13253), .ZN(
        n16400) );
  AOI22_X1 U15046 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13418), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13257) );
  AOI22_X1 U15047 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13256) );
  AOI22_X1 U15048 ( .A1(n12644), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13255) );
  AOI22_X1 U15049 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13526), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13254) );
  NAND4_X1 U15050 ( .A1(n13257), .A2(n13256), .A3(n13255), .A4(n13254), .ZN(
        n13263) );
  AOI22_X1 U15051 ( .A1(n13564), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13261) );
  AOI22_X1 U15052 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13578), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13260) );
  AOI22_X1 U15053 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12624), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13259) );
  AOI22_X1 U15054 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13258) );
  NAND4_X1 U15055 ( .A1(n13261), .A2(n13260), .A3(n13259), .A4(n13258), .ZN(
        n13262) );
  OR2_X1 U15056 ( .A1(n13263), .A2(n13262), .ZN(n13264) );
  AOI22_X1 U15057 ( .A1(n13312), .A2(n13264), .B1(n13604), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n13266) );
  NAND2_X1 U15058 ( .A1(n13599), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n13265) );
  OAI211_X1 U15059 ( .C1(n16400), .C2(n13597), .A(n13266), .B(n13265), .ZN(
        n15907) );
  INV_X1 U15060 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n21929) );
  AOI22_X1 U15061 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13419), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13270) );
  AOI22_X1 U15062 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12645), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13269) );
  AOI22_X1 U15063 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13268) );
  AOI22_X1 U15064 ( .A1(n11021), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13526), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13267) );
  NAND4_X1 U15065 ( .A1(n13270), .A2(n13269), .A3(n13268), .A4(n13267), .ZN(
        n13276) );
  AOI22_X1 U15066 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13274) );
  AOI22_X1 U15067 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12644), .B1(
        n13418), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13273) );
  AOI22_X1 U15068 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13578), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13272) );
  AOI22_X1 U15069 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n13584), .B1(
        n12624), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13271) );
  NAND4_X1 U15070 ( .A1(n13274), .A2(n13273), .A3(n13272), .A4(n13271), .ZN(
        n13275) );
  OAI21_X1 U15071 ( .B1(n13276), .B2(n13275), .A(n13312), .ZN(n13279) );
  XNOR2_X1 U15072 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n13281), .ZN(
        n21713) );
  INV_X1 U15073 ( .A(n21713), .ZN(n13277) );
  AOI22_X1 U15074 ( .A1(n13604), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n13600), .B2(n13277), .ZN(n13278) );
  OAI211_X1 U15075 ( .C1(n13137), .C2(n21929), .A(n13279), .B(n13278), .ZN(
        n15922) );
  OR2_X1 U15076 ( .A1(n13280), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13282) );
  NAND2_X1 U15077 ( .A1(n13282), .A2(n13281), .ZN(n21701) );
  INV_X1 U15078 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n21919) );
  INV_X1 U15079 ( .A(n13604), .ZN(n13284) );
  INV_X1 U15080 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n13283) );
  OAI22_X1 U15081 ( .A1(n13137), .A2(n21919), .B1(n13284), .B2(n13283), .ZN(
        n13285) );
  AOI21_X1 U15082 ( .B1(n21701), .B2(n13600), .A(n13285), .ZN(n15901) );
  AOI22_X1 U15083 ( .A1(n12644), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11016), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13290) );
  AOI22_X1 U15084 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13289) );
  AOI22_X1 U15085 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13578), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13288) );
  AOI22_X1 U15086 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13526), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13287) );
  NAND4_X1 U15087 ( .A1(n13290), .A2(n13289), .A3(n13288), .A4(n13287), .ZN(
        n13296) );
  AOI22_X1 U15088 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13294) );
  AOI22_X1 U15089 ( .A1(n13585), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13293) );
  AOI22_X1 U15090 ( .A1(n13418), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12624), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13292) );
  AOI22_X1 U15091 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13291) );
  NAND4_X1 U15092 ( .A1(n13294), .A2(n13293), .A3(n13292), .A4(n13291), .ZN(
        n13295) );
  OR2_X1 U15093 ( .A1(n13296), .A2(n13295), .ZN(n13297) );
  NAND2_X1 U15094 ( .A1(n13312), .A2(n13297), .ZN(n15791) );
  NAND2_X1 U15095 ( .A1(n15901), .A2(n15791), .ZN(n13298) );
  NAND3_X1 U15096 ( .A1(n15907), .A2(n15922), .A3(n13298), .ZN(n15833) );
  XNOR2_X1 U15097 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n13315), .ZN(
        n21722) );
  AOI22_X1 U15098 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12650), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13304) );
  AOI22_X1 U15099 ( .A1(n12644), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13419), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13303) );
  AOI22_X1 U15100 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13302) );
  AOI22_X1 U15101 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13526), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13301) );
  NAND4_X1 U15102 ( .A1(n13304), .A2(n13303), .A3(n13302), .A4(n13301), .ZN(
        n13310) );
  AOI22_X1 U15103 ( .A1(n13564), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11022), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13308) );
  AOI22_X1 U15104 ( .A1(n13418), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13578), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13307) );
  AOI22_X1 U15105 ( .A1(n13584), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12624), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13306) );
  AOI22_X1 U15106 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13305) );
  NAND4_X1 U15107 ( .A1(n13308), .A2(n13307), .A3(n13306), .A4(n13305), .ZN(
        n13309) );
  OR2_X1 U15108 ( .A1(n13310), .A2(n13309), .ZN(n13311) );
  AOI22_X1 U15109 ( .A1(n13312), .A2(n13311), .B1(n13604), .B2(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n13314) );
  NAND2_X1 U15110 ( .A1(n13165), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n13313) );
  OAI211_X1 U15111 ( .C1(n21722), .C2(n13597), .A(n13314), .B(n13313), .ZN(
        n15936) );
  INV_X1 U15112 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16386) );
  XNOR2_X1 U15113 ( .A(n13330), .B(n16386), .ZN(n21732) );
  AOI22_X1 U15114 ( .A1(n13165), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n22106), .ZN(n13329) );
  AOI22_X1 U15115 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13192), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13319) );
  AOI22_X1 U15116 ( .A1(n13418), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11021), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13318) );
  AOI22_X1 U15117 ( .A1(n13564), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13238), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13317) );
  AOI22_X1 U15118 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13526), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13316) );
  NAND4_X1 U15119 ( .A1(n13319), .A2(n13318), .A3(n13317), .A4(n13316), .ZN(
        n13327) );
  AOI22_X1 U15120 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13325) );
  AOI22_X1 U15121 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13324) );
  AOI22_X1 U15122 ( .A1(n12644), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13578), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13323) );
  AOI21_X1 U15123 ( .B1(n13579), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A(
        n13600), .ZN(n13321) );
  NAND2_X1 U15124 ( .A1(n12624), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n13320) );
  AND2_X1 U15125 ( .A1(n13321), .A2(n13320), .ZN(n13322) );
  NAND4_X1 U15126 ( .A1(n13325), .A2(n13324), .A3(n13323), .A4(n13322), .ZN(
        n13326) );
  NAND2_X1 U15127 ( .A1(n13573), .A2(n13597), .ZN(n13426) );
  OAI21_X1 U15128 ( .B1(n13327), .B2(n13326), .A(n13426), .ZN(n13328) );
  AOI22_X1 U15129 ( .A1(n21732), .A2(n13600), .B1(n13329), .B2(n13328), .ZN(
        n15863) );
  XNOR2_X1 U15130 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n13343), .ZN(
        n20171) );
  AOI22_X1 U15131 ( .A1(n13165), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n13604), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n13342) );
  AOI22_X1 U15132 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13334) );
  AOI22_X1 U15133 ( .A1(n13578), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13333) );
  AOI22_X1 U15134 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13332) );
  AOI22_X1 U15135 ( .A1(n12693), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13526), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13331) );
  NAND4_X1 U15136 ( .A1(n13334), .A2(n13333), .A3(n13332), .A4(n13331), .ZN(
        n13340) );
  AOI22_X1 U15137 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13338) );
  AOI22_X1 U15138 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12650), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13337) );
  AOI22_X1 U15139 ( .A1(n12685), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13336) );
  AOI22_X1 U15140 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13418), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13335) );
  NAND4_X1 U15141 ( .A1(n13338), .A2(n13337), .A3(n13336), .A4(n13335), .ZN(
        n13339) );
  INV_X1 U15142 ( .A(n13573), .ZN(n13594) );
  OAI21_X1 U15143 ( .B1(n13340), .B2(n13339), .A(n13594), .ZN(n13341) );
  OAI211_X1 U15144 ( .C1(n20171), .C2(n13597), .A(n13342), .B(n13341), .ZN(
        n15964) );
  INV_X1 U15145 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16195) );
  INV_X1 U15146 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n13344) );
  XNOR2_X1 U15147 ( .A(n13375), .B(n13344), .ZN(n16375) );
  NAND2_X1 U15148 ( .A1(n16375), .A2(n13600), .ZN(n13360) );
  AOI22_X1 U15149 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12650), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13348) );
  AOI22_X1 U15150 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13192), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13347) );
  AOI22_X1 U15151 ( .A1(n11021), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13238), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13346) );
  AOI22_X1 U15152 ( .A1(n13584), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12693), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13345) );
  NAND4_X1 U15153 ( .A1(n13348), .A2(n13347), .A3(n13346), .A4(n13345), .ZN(
        n13356) );
  AOI22_X1 U15154 ( .A1(n12685), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13418), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13354) );
  AOI22_X1 U15155 ( .A1(n13585), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13578), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13353) );
  AOI22_X1 U15156 ( .A1(n13564), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13526), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13352) );
  NAND2_X1 U15157 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n13350) );
  AOI21_X1 U15158 ( .B1(n13579), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A(
        n13600), .ZN(n13349) );
  AND2_X1 U15159 ( .A1(n13350), .A2(n13349), .ZN(n13351) );
  NAND4_X1 U15160 ( .A1(n13354), .A2(n13353), .A3(n13352), .A4(n13351), .ZN(
        n13355) );
  OAI21_X1 U15161 ( .B1(n13356), .B2(n13355), .A(n13426), .ZN(n13358) );
  AOI22_X1 U15162 ( .A1(n13165), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n22106), .ZN(n13357) );
  NAND2_X1 U15163 ( .A1(n13358), .A2(n13357), .ZN(n13359) );
  NAND2_X1 U15164 ( .A1(n13360), .A2(n13359), .ZN(n16188) );
  NOR2_X2 U15165 ( .A1(n15965), .A2(n16188), .ZN(n16186) );
  AOI22_X1 U15166 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12650), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13364) );
  AOI22_X1 U15167 ( .A1(n12685), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13363) );
  AOI22_X1 U15168 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11022), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13362) );
  AOI22_X1 U15169 ( .A1(n13418), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13526), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13361) );
  NAND4_X1 U15170 ( .A1(n13364), .A2(n13363), .A3(n13362), .A4(n13361), .ZN(
        n13370) );
  AOI22_X1 U15171 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13368) );
  AOI22_X1 U15172 ( .A1(n13564), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13578), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13367) );
  AOI22_X1 U15173 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12693), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13366) );
  AOI22_X1 U15174 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13365) );
  NAND4_X1 U15175 ( .A1(n13368), .A2(n13367), .A3(n13366), .A4(n13365), .ZN(
        n13369) );
  NOR2_X1 U15176 ( .A1(n13370), .A2(n13369), .ZN(n13374) );
  NAND2_X1 U15177 ( .A1(n22106), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13371) );
  NAND2_X1 U15178 ( .A1(n13597), .A2(n13371), .ZN(n13372) );
  AOI21_X1 U15179 ( .B1(n13599), .B2(P1_EAX_REG_19__SCAN_IN), .A(n13372), .ZN(
        n13373) );
  OAI21_X1 U15180 ( .B1(n13573), .B2(n13374), .A(n13373), .ZN(n13378) );
  OAI21_X1 U15181 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n13376), .A(
        n13409), .ZN(n21746) );
  OR2_X1 U15182 ( .A1(n13597), .A2(n21746), .ZN(n13377) );
  NAND2_X1 U15183 ( .A1(n13378), .A2(n13377), .ZN(n16234) );
  AOI22_X1 U15184 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12644), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13385) );
  AOI22_X1 U15185 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n13585), .B1(
        n11021), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13384) );
  AOI22_X1 U15186 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13526), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13383) );
  NAND2_X1 U15187 ( .A1(n12624), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n13381) );
  NAND2_X1 U15188 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n13380) );
  AND3_X1 U15189 ( .A1(n13381), .A2(n13380), .A3(n13597), .ZN(n13382) );
  NAND4_X1 U15190 ( .A1(n13385), .A2(n13384), .A3(n13383), .A4(n13382), .ZN(
        n13391) );
  AOI22_X1 U15191 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13418), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13389) );
  AOI22_X1 U15192 ( .A1(n13584), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13192), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13388) );
  AOI22_X1 U15193 ( .A1(n13564), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13578), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13387) );
  AOI22_X1 U15194 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13386) );
  NAND4_X1 U15195 ( .A1(n13389), .A2(n13388), .A3(n13387), .A4(n13386), .ZN(
        n13390) );
  OR2_X1 U15196 ( .A1(n13391), .A2(n13390), .ZN(n13392) );
  NAND2_X1 U15197 ( .A1(n13426), .A2(n13392), .ZN(n13395) );
  AOI22_X1 U15198 ( .A1(n13165), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n22106), .ZN(n13394) );
  XNOR2_X1 U15199 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n13409), .ZN(
        n21768) );
  AOI21_X1 U15200 ( .B1(n13395), .B2(n13394), .A(n13393), .ZN(n16229) );
  AOI22_X1 U15201 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13399) );
  AOI22_X1 U15202 ( .A1(n12685), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13398) );
  AOI22_X1 U15203 ( .A1(n13418), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12693), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13397) );
  AOI22_X1 U15204 ( .A1(n13564), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11021), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13396) );
  NAND4_X1 U15205 ( .A1(n13399), .A2(n13398), .A3(n13397), .A4(n13396), .ZN(
        n13405) );
  AOI22_X1 U15206 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12650), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13403) );
  AOI22_X1 U15207 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13578), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13402) );
  AOI22_X1 U15208 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13401) );
  AOI22_X1 U15209 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13526), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13400) );
  NAND4_X1 U15210 ( .A1(n13403), .A2(n13402), .A3(n13401), .A4(n13400), .ZN(
        n13404) );
  NOR2_X1 U15211 ( .A1(n13405), .A2(n13404), .ZN(n13406) );
  OR2_X1 U15212 ( .A1(n13573), .A2(n13406), .ZN(n13413) );
  NAND2_X1 U15213 ( .A1(n22106), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13407) );
  NAND2_X1 U15214 ( .A1(n13597), .A2(n13407), .ZN(n13408) );
  AOI21_X1 U15215 ( .B1(n13599), .B2(P1_EAX_REG_21__SCAN_IN), .A(n13408), .ZN(
        n13412) );
  INV_X1 U15216 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n21763) );
  OAI21_X1 U15217 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n13410), .A(
        n13434), .ZN(n20191) );
  NOR2_X1 U15218 ( .A1(n20191), .A2(n13597), .ZN(n13411) );
  AOI21_X1 U15219 ( .B1(n13413), .B2(n13412), .A(n13411), .ZN(n16172) );
  AOI22_X1 U15220 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12650), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13417) );
  AOI22_X1 U15221 ( .A1(n13585), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13578), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13416) );
  AOI22_X1 U15222 ( .A1(n12685), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12693), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13415) );
  AOI22_X1 U15223 ( .A1(n12612), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13238), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13414) );
  NAND4_X1 U15224 ( .A1(n13417), .A2(n13416), .A3(n13415), .A4(n13414), .ZN(
        n13428) );
  AOI22_X1 U15225 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13425) );
  AOI22_X1 U15226 ( .A1(n13584), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13192), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13424) );
  AOI22_X1 U15227 ( .A1(n13418), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13526), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13423) );
  NAND2_X1 U15228 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n13421) );
  AOI21_X1 U15229 ( .B1(n13579), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n13600), .ZN(n13420) );
  AND2_X1 U15230 ( .A1(n13421), .A2(n13420), .ZN(n13422) );
  NAND4_X1 U15231 ( .A1(n13425), .A2(n13424), .A3(n13423), .A4(n13422), .ZN(
        n13427) );
  OAI21_X1 U15232 ( .B1(n13428), .B2(n13427), .A(n13426), .ZN(n13430) );
  AOI22_X1 U15233 ( .A1(n13165), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n22106), .ZN(n13429) );
  NAND2_X1 U15234 ( .A1(n13430), .A2(n13429), .ZN(n13432) );
  XNOR2_X1 U15235 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B(n13434), .ZN(
        n16360) );
  NAND2_X1 U15236 ( .A1(n13600), .A2(n16360), .ZN(n13431) );
  NAND2_X1 U15237 ( .A1(n13432), .A2(n13431), .ZN(n16160) );
  INV_X1 U15238 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n13433) );
  OR2_X1 U15239 ( .A1(n13435), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13436) );
  NAND2_X1 U15240 ( .A1(n13436), .A2(n13478), .ZN(n20199) );
  AOI22_X1 U15241 ( .A1(n12644), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13419), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13440) );
  AOI22_X1 U15242 ( .A1(n13418), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13578), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13439) );
  AOI22_X1 U15243 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11022), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13438) );
  AOI22_X1 U15244 ( .A1(n13564), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13238), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13437) );
  NAND4_X1 U15245 ( .A1(n13440), .A2(n13439), .A3(n13438), .A4(n13437), .ZN(
        n13446) );
  AOI22_X1 U15246 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13444) );
  AOI22_X1 U15247 ( .A1(n13584), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12624), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13443) );
  AOI22_X1 U15248 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13442) );
  AOI22_X1 U15249 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13526), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13441) );
  NAND4_X1 U15250 ( .A1(n13444), .A2(n13443), .A3(n13442), .A4(n13441), .ZN(
        n13445) );
  NOR2_X1 U15251 ( .A1(n13446), .A2(n13445), .ZN(n13462) );
  AOI22_X1 U15252 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13450) );
  AOI22_X1 U15253 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13578), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13449) );
  AOI22_X1 U15254 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13238), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13448) );
  AOI22_X1 U15255 ( .A1(n12644), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13526), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13447) );
  NAND4_X1 U15256 ( .A1(n13450), .A2(n13449), .A3(n13448), .A4(n13447), .ZN(
        n13456) );
  AOI22_X1 U15257 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13454) );
  AOI22_X1 U15258 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13418), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13453) );
  AOI22_X1 U15259 ( .A1(n12612), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13452) );
  AOI22_X1 U15260 ( .A1(n13585), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12624), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13451) );
  NAND4_X1 U15261 ( .A1(n13454), .A2(n13453), .A3(n13452), .A4(n13451), .ZN(
        n13455) );
  NOR2_X1 U15262 ( .A1(n13456), .A2(n13455), .ZN(n13463) );
  XNOR2_X1 U15263 ( .A(n13462), .B(n13463), .ZN(n13457) );
  NOR2_X1 U15264 ( .A1(n13573), .A2(n13457), .ZN(n13460) );
  INV_X1 U15265 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n16272) );
  NAND2_X1 U15266 ( .A1(n22106), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13458) );
  OAI211_X1 U15267 ( .C1(n13137), .C2(n16272), .A(n13597), .B(n13458), .ZN(
        n13459) );
  OAI22_X1 U15268 ( .A1(n20199), .A2(n13597), .B1(n13460), .B2(n13459), .ZN(
        n16144) );
  XNOR2_X1 U15269 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B(n13478), .ZN(
        n21781) );
  INV_X1 U15270 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n21775) );
  OAI21_X1 U15271 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n21775), .A(n13597), 
        .ZN(n13476) );
  NOR2_X1 U15272 ( .A1(n13463), .A2(n13462), .ZN(n13482) );
  AOI22_X1 U15273 ( .A1(n12644), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13467) );
  AOI22_X1 U15274 ( .A1(n13418), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13466) );
  AOI22_X1 U15275 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13526), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13465) );
  AOI22_X1 U15276 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12624), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13464) );
  NAND4_X1 U15277 ( .A1(n13467), .A2(n13466), .A3(n13465), .A4(n13464), .ZN(
        n13473) );
  AOI22_X1 U15278 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13471) );
  AOI22_X1 U15279 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13578), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13470) );
  AOI22_X1 U15280 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11021), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13469) );
  AOI22_X1 U15281 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13468) );
  NAND4_X1 U15282 ( .A1(n13471), .A2(n13470), .A3(n13469), .A4(n13468), .ZN(
        n13472) );
  OR2_X1 U15283 ( .A1(n13473), .A2(n13472), .ZN(n13481) );
  XNOR2_X1 U15284 ( .A(n13482), .B(n13481), .ZN(n13474) );
  NOR2_X1 U15285 ( .A1(n13474), .A2(n13573), .ZN(n13475) );
  AOI211_X1 U15286 ( .C1(n13599), .C2(P1_EAX_REG_24__SCAN_IN), .A(n13476), .B(
        n13475), .ZN(n13477) );
  OAI21_X1 U15287 ( .B1(n13480), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n13516), .ZN(n16347) );
  NAND2_X1 U15288 ( .A1(n13482), .A2(n13481), .ZN(n13497) );
  AOI22_X1 U15289 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13486) );
  AOI22_X1 U15290 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13578), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13485) );
  AOI22_X1 U15291 ( .A1(n13418), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12624), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13484) );
  AOI22_X1 U15292 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13483) );
  NAND4_X1 U15293 ( .A1(n13486), .A2(n13485), .A3(n13484), .A4(n13483), .ZN(
        n13492) );
  AOI22_X1 U15294 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13490) );
  AOI22_X1 U15295 ( .A1(n12644), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13489) );
  AOI22_X1 U15296 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11022), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13488) );
  AOI22_X1 U15297 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13526), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13487) );
  NAND4_X1 U15298 ( .A1(n13490), .A2(n13489), .A3(n13488), .A4(n13487), .ZN(
        n13491) );
  NOR2_X1 U15299 ( .A1(n13492), .A2(n13491), .ZN(n13498) );
  XNOR2_X1 U15300 ( .A(n13497), .B(n13498), .ZN(n13495) );
  AOI21_X1 U15301 ( .B1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n22106), .A(
        n13600), .ZN(n13494) );
  NAND2_X1 U15302 ( .A1(n13165), .A2(P1_EAX_REG_25__SCAN_IN), .ZN(n13493) );
  OAI211_X1 U15303 ( .C1(n13495), .C2(n13573), .A(n13494), .B(n13493), .ZN(
        n13496) );
  OAI21_X1 U15304 ( .B1(n13597), .B2(n16347), .A(n13496), .ZN(n16128) );
  XNOR2_X1 U15305 ( .A(n13516), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16340) );
  INV_X1 U15306 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16336) );
  OAI21_X1 U15307 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n16336), .A(n13597), 
        .ZN(n13514) );
  NOR2_X1 U15308 ( .A1(n13498), .A2(n13497), .ZN(n13521) );
  INV_X1 U15309 ( .A(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13499) );
  NOR2_X1 U15310 ( .A1(n12692), .A2(n13499), .ZN(n13503) );
  INV_X1 U15311 ( .A(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13501) );
  OAI22_X1 U15312 ( .A1(n12465), .A2(n13501), .B1(n11023), .B2(n13500), .ZN(
        n13502) );
  AOI211_X1 U15313 ( .C1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .C2(n12650), .A(
        n13503), .B(n13502), .ZN(n13511) );
  AOI22_X1 U15314 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13510) );
  AOI22_X1 U15315 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13509) );
  AOI22_X1 U15316 ( .A1(n12644), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13507) );
  AOI22_X1 U15317 ( .A1(n13418), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13506) );
  AOI22_X1 U15318 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13526), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13505) );
  AOI22_X1 U15319 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12693), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13504) );
  AND4_X1 U15320 ( .A1(n13507), .A2(n13506), .A3(n13505), .A4(n13504), .ZN(
        n13508) );
  NAND4_X1 U15321 ( .A1(n13511), .A2(n13510), .A3(n13509), .A4(n13508), .ZN(
        n13520) );
  XNOR2_X1 U15322 ( .A(n13521), .B(n13520), .ZN(n13512) );
  NOR2_X1 U15323 ( .A1(n13512), .A2(n13573), .ZN(n13513) );
  AOI211_X1 U15324 ( .C1(n13165), .C2(P1_EAX_REG_26__SCAN_IN), .A(n13514), .B(
        n13513), .ZN(n13515) );
  AOI21_X1 U15325 ( .B1(n13600), .B2(n16340), .A(n13515), .ZN(n16115) );
  NAND2_X1 U15326 ( .A1(n16113), .A2(n16115), .ZN(n16103) );
  INV_X1 U15327 ( .A(n13517), .ZN(n13518) );
  INV_X1 U15328 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16106) );
  NAND2_X1 U15329 ( .A1(n13518), .A2(n16106), .ZN(n13519) );
  NAND2_X1 U15330 ( .A1(n13553), .A2(n13519), .ZN(n16329) );
  NAND2_X1 U15331 ( .A1(n13521), .A2(n13520), .ZN(n13537) );
  AOI22_X1 U15332 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n12645), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13525) );
  AOI22_X1 U15333 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13578), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13524) );
  AOI22_X1 U15334 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n13584), .B1(
        n12624), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13523) );
  AOI22_X1 U15335 ( .A1(n13564), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13238), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13522) );
  NAND4_X1 U15336 ( .A1(n13525), .A2(n13524), .A3(n13523), .A4(n13522), .ZN(
        n13532) );
  AOI22_X1 U15337 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n12644), .B1(
        n13419), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13530) );
  AOI22_X1 U15338 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n13585), .B1(
        n13418), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13529) );
  AOI22_X1 U15339 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13528) );
  AOI22_X1 U15340 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13526), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13527) );
  NAND4_X1 U15341 ( .A1(n13530), .A2(n13529), .A3(n13528), .A4(n13527), .ZN(
        n13531) );
  NOR2_X1 U15342 ( .A1(n13532), .A2(n13531), .ZN(n13538) );
  XNOR2_X1 U15343 ( .A(n13537), .B(n13538), .ZN(n13535) );
  AOI21_X1 U15344 ( .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n22106), .A(
        n13600), .ZN(n13534) );
  NAND2_X1 U15345 ( .A1(n13165), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n13533) );
  OAI211_X1 U15346 ( .C1(n13535), .C2(n13573), .A(n13534), .B(n13533), .ZN(
        n13536) );
  XNOR2_X1 U15347 ( .A(n13553), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16097) );
  INV_X1 U15348 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16091) );
  AOI21_X1 U15349 ( .B1(n16091), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13551) );
  NOR2_X1 U15350 ( .A1(n13538), .A2(n13537), .ZN(n13559) );
  AOI22_X1 U15351 ( .A1(n12685), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13542) );
  AOI22_X1 U15352 ( .A1(n13418), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13541) );
  AOI22_X1 U15353 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13526), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13540) );
  AOI22_X1 U15354 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12693), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13539) );
  NAND4_X1 U15355 ( .A1(n13542), .A2(n13541), .A3(n13540), .A4(n13539), .ZN(
        n13548) );
  AOI22_X1 U15356 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13546) );
  AOI22_X1 U15357 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13578), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13545) );
  AOI22_X1 U15358 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11021), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13544) );
  AOI22_X1 U15359 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13543) );
  NAND4_X1 U15360 ( .A1(n13546), .A2(n13545), .A3(n13544), .A4(n13543), .ZN(
        n13547) );
  OR2_X1 U15361 ( .A1(n13548), .A2(n13547), .ZN(n13558) );
  XNOR2_X1 U15362 ( .A(n13559), .B(n13558), .ZN(n13549) );
  NOR2_X1 U15363 ( .A1(n13549), .A2(n13573), .ZN(n13550) );
  AOI211_X1 U15364 ( .C1(n13165), .C2(P1_EAX_REG_28__SCAN_IN), .A(n13551), .B(
        n13550), .ZN(n13552) );
  INV_X1 U15365 ( .A(n13553), .ZN(n13554) );
  INV_X1 U15366 ( .A(n13555), .ZN(n13556) );
  INV_X1 U15367 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16079) );
  NAND2_X1 U15368 ( .A1(n13556), .A2(n16079), .ZN(n13557) );
  NAND2_X1 U15369 ( .A1(n13612), .A2(n13557), .ZN(n16323) );
  NAND2_X1 U15370 ( .A1(n13559), .A2(n13558), .ZN(n13576) );
  AOI22_X1 U15371 ( .A1(n12685), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13563) );
  AOI22_X1 U15372 ( .A1(n12612), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13238), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13562) );
  AOI22_X1 U15373 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12624), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13561) );
  AOI22_X1 U15374 ( .A1(n13585), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13526), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13560) );
  NAND4_X1 U15375 ( .A1(n13563), .A2(n13562), .A3(n13561), .A4(n13560), .ZN(
        n13570) );
  AOI22_X1 U15376 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12650), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13568) );
  AOI22_X1 U15377 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13418), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13567) );
  AOI22_X1 U15378 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13578), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13566) );
  AOI22_X1 U15379 ( .A1(n13564), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13565) );
  NAND4_X1 U15380 ( .A1(n13568), .A2(n13567), .A3(n13566), .A4(n13565), .ZN(
        n13569) );
  NOR2_X1 U15381 ( .A1(n13570), .A2(n13569), .ZN(n13577) );
  XNOR2_X1 U15382 ( .A(n13576), .B(n13577), .ZN(n13574) );
  AOI21_X1 U15383 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n22106), .A(
        n13600), .ZN(n13572) );
  NAND2_X1 U15384 ( .A1(n13165), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n13571) );
  OAI211_X1 U15385 ( .C1(n13574), .C2(n13573), .A(n13572), .B(n13571), .ZN(
        n13575) );
  OAI21_X1 U15386 ( .B1(n13597), .B2(n16323), .A(n13575), .ZN(n13620) );
  NOR2_X1 U15387 ( .A1(n13577), .A2(n13576), .ZN(n13593) );
  AOI22_X1 U15388 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13578), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13583) );
  AOI22_X1 U15389 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11021), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13582) );
  AOI22_X1 U15390 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13579), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13581) );
  AOI22_X1 U15391 ( .A1(n13192), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13526), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13580) );
  NAND4_X1 U15392 ( .A1(n13583), .A2(n13582), .A3(n13581), .A4(n13580), .ZN(
        n13591) );
  AOI22_X1 U15393 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13589) );
  AOI22_X1 U15394 ( .A1(n12685), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13588) );
  AOI22_X1 U15395 ( .A1(n13418), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13587) );
  AOI22_X1 U15396 ( .A1(n13419), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12693), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13586) );
  NAND4_X1 U15397 ( .A1(n13589), .A2(n13588), .A3(n13587), .A4(n13586), .ZN(
        n13590) );
  NOR2_X1 U15398 ( .A1(n13591), .A2(n13590), .ZN(n13592) );
  XNOR2_X1 U15399 ( .A(n13593), .B(n13592), .ZN(n13595) );
  NAND2_X1 U15400 ( .A1(n13595), .A2(n13594), .ZN(n13603) );
  NAND2_X1 U15401 ( .A1(n22106), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13596) );
  NAND2_X1 U15402 ( .A1(n13597), .A2(n13596), .ZN(n13598) );
  AOI21_X1 U15403 ( .B1(n13599), .B2(P1_EAX_REG_30__SCAN_IN), .A(n13598), .ZN(
        n13602) );
  XNOR2_X1 U15404 ( .A(n13612), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16312) );
  AND2_X1 U15405 ( .A1(n16312), .A2(n13600), .ZN(n13601) );
  AOI22_X1 U15406 ( .A1(n13165), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n13604), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13605) );
  INV_X1 U15407 ( .A(n13605), .ZN(n13606) );
  XNOR2_X2 U15408 ( .A(n13607), .B(n13606), .ZN(n16250) );
  NAND3_X1 U15409 ( .A1(n21804), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n21801) );
  INV_X1 U15410 ( .A(n21801), .ZN(n13608) );
  NAND2_X1 U15411 ( .A1(n16250), .A2(n20186), .ZN(n13619) );
  INV_X1 U15412 ( .A(n22117), .ZN(n22115) );
  NAND2_X1 U15413 ( .A1(n22115), .A2(n13609), .ZN(n21514) );
  NAND2_X1 U15414 ( .A1(n21514), .A2(n21804), .ZN(n13610) );
  NAND2_X1 U15415 ( .A1(n21804), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17349) );
  NAND2_X1 U15416 ( .A1(n15084), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13611) );
  NAND2_X1 U15417 ( .A1(n17349), .A2(n13611), .ZN(n20138) );
  INV_X1 U15418 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16314) );
  INV_X1 U15419 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13613) );
  AOI21_X1 U15420 ( .B1(n20192), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n13615), .ZN(n13616) );
  OAI21_X1 U15421 ( .B1(n20200), .B2(n15161), .A(n13616), .ZN(n13617) );
  INV_X1 U15422 ( .A(n13617), .ZN(n13618) );
  INV_X1 U15423 ( .A(n14532), .ZN(n13622) );
  NOR2_X1 U15424 ( .A1(n14811), .A2(n21813), .ZN(n13624) );
  NAND4_X1 U15425 ( .A1(n15215), .A2(n14700), .A3(n13624), .A4(n13623), .ZN(
        n14807) );
  NAND2_X1 U15426 ( .A1(n16325), .A2(n13627), .ZN(n13634) );
  NOR2_X1 U15427 ( .A1(n16088), .A2(n13628), .ZN(n13629) );
  NOR2_X1 U15428 ( .A1(n20137), .A2(n16078), .ZN(n13630) );
  NOR2_X1 U15429 ( .A1(n14705), .A2(n21813), .ZN(n13636) );
  NAND2_X1 U15430 ( .A1(n14803), .A2(n13636), .ZN(n14620) );
  NAND2_X2 U15431 ( .A1(n14744), .A2(n14620), .ZN(n21513) );
  OAI211_X1 U15432 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n21798), .A(n21794), 
        .B(n21804), .ZN(n13638) );
  NAND2_X1 U15433 ( .A1(n21798), .A2(n22106), .ZN(n21511) );
  OAI22_X1 U15434 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_0__SCAN_IN), .B1(n21511), .B2(n22072), .ZN(n13637) );
  AND2_X1 U15435 ( .A1(n13638), .A2(n13637), .ZN(n13639) );
  OR2_X4 U15436 ( .A1(n21513), .A2(n13639), .ZN(n16136) );
  NOR2_X1 U15437 ( .A1(n15161), .A2(n21798), .ZN(n13640) );
  NAND2_X1 U15438 ( .A1(n16136), .A2(n13640), .ZN(n21777) );
  NAND2_X1 U15439 ( .A1(n16250), .A2(n21754), .ZN(n13659) );
  NOR2_X2 U15440 ( .A1(n12966), .A2(n15163), .ZN(n13647) );
  NAND2_X1 U15441 ( .A1(n14745), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13642) );
  AND2_X1 U15442 ( .A1(n21834), .A2(n15084), .ZN(n17346) );
  NOR2_X1 U15443 ( .A1(n13642), .A2(n17346), .ZN(n13641) );
  NAND2_X1 U15444 ( .A1(n13647), .A2(n13642), .ZN(n13644) );
  INV_X1 U15445 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n16207) );
  INV_X1 U15446 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n21696) );
  INV_X1 U15447 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20074) );
  NAND4_X1 U15448 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_19__SCAN_IN), .A4(P1_REIP_REG_18__SCAN_IN), .ZN(n13646) );
  NAND4_X1 U15449 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(P1_REIP_REG_17__SCAN_IN), 
        .A3(P1_REIP_REG_13__SCAN_IN), .A4(P1_REIP_REG_12__SCAN_IN), .ZN(n13645) );
  NOR4_X1 U15450 ( .A1(n21696), .A2(n20074), .A3(n13646), .A4(n13645), .ZN(
        n16139) );
  NAND3_X1 U15451 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .A3(P1_REIP_REG_10__SCAN_IN), .ZN(n16138) );
  NAND4_X1 U15452 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_4__SCAN_IN), .ZN(n21623)
         );
  INV_X1 U15453 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21627) );
  NOR2_X1 U15454 ( .A1(n21623), .A2(n21627), .ZN(n16137) );
  INV_X1 U15455 ( .A(n16137), .ZN(n13649) );
  OR2_X2 U15456 ( .A1(n21622), .A2(n13649), .ZN(n21638) );
  INV_X1 U15457 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20053) );
  NOR2_X2 U15458 ( .A1(n21638), .A2(n20053), .ZN(n21656) );
  NOR2_X2 U15459 ( .A1(n16138), .A2(n21666), .ZN(n21707) );
  NAND2_X1 U15460 ( .A1(n16139), .A2(n21707), .ZN(n16183) );
  INV_X1 U15461 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20076) );
  NOR2_X2 U15462 ( .A1(n16183), .A2(n20076), .ZN(n16169) );
  NAND2_X1 U15463 ( .A1(n16169), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n16151) );
  INV_X1 U15464 ( .A(n16151), .ZN(n13650) );
  AND2_X2 U15465 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n13650), .ZN(n21785) );
  NAND2_X1 U15466 ( .A1(n21785), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n16133) );
  NAND2_X1 U15467 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n13651) );
  NOR2_X2 U15468 ( .A1(n16133), .A2(n13651), .ZN(n16123) );
  NAND2_X1 U15469 ( .A1(n16123), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n16110) );
  INV_X1 U15470 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n13652) );
  OR2_X2 U15471 ( .A1(n16110), .A2(n13652), .ZN(n16092) );
  INV_X1 U15472 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20089) );
  NOR2_X2 U15473 ( .A1(n16092), .A2(n20089), .ZN(n16080) );
  NAND2_X1 U15474 ( .A1(n16080), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n13653) );
  OAI22_X1 U15475 ( .A1(n21761), .A2(n16207), .B1(P1_REIP_REG_31__SCAN_IN), 
        .B2(n13653), .ZN(n13655) );
  NAND2_X1 U15476 ( .A1(n16136), .A2(n21622), .ZN(n21738) );
  AND3_X1 U15477 ( .A1(n21738), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n13653), 
        .ZN(n13654) );
  OAI21_X1 U15478 ( .B1(n16208), .B2(n21788), .A(n13656), .ZN(n13657) );
  NAND2_X1 U15479 ( .A1(n13659), .A2(n13658), .ZN(P1_U2809) );
  AOI222_X1 U15480 ( .A1(n12021), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n13660), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n11015), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13661) );
  INV_X1 U15481 ( .A(n13661), .ZN(n13662) );
  INV_X2 U15482 ( .A(n18621), .ZN(n18851) );
  NOR2_X1 U15483 ( .A1(n13664), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13665) );
  MUX2_X1 U15484 ( .A(n12198), .B(n13665), .S(n19633), .Z(n16037) );
  INV_X1 U15485 ( .A(n16037), .ZN(n13666) );
  INV_X1 U15486 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n17764) );
  OAI22_X1 U15487 ( .A1(n13666), .A2(n18803), .B1(n17764), .B2(n18748), .ZN(
        n13667) );
  AOI21_X1 U15488 ( .B1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n18851), .A(
        n13667), .ZN(n13669) );
  INV_X1 U15489 ( .A(n13672), .ZN(n13674) );
  NAND2_X1 U15490 ( .A1(n18861), .A2(n18752), .ZN(n18605) );
  INV_X1 U15491 ( .A(n18605), .ZN(n13673) );
  NAND2_X1 U15492 ( .A1(n13674), .A2(n13673), .ZN(n13685) );
  INV_X1 U15493 ( .A(n13675), .ZN(n13677) );
  NAND2_X1 U15494 ( .A1(n13677), .A2(n13676), .ZN(n13683) );
  AOI22_X1 U15495 ( .A1(n13678), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n13679) );
  OAI21_X1 U15496 ( .B1(n11464), .B2(n13680), .A(n13679), .ZN(n13681) );
  AOI21_X1 U15497 ( .B1(n12398), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n13681), .ZN(n13682) );
  XNOR2_X2 U15498 ( .A(n13683), .B(n13682), .ZN(n16777) );
  INV_X1 U15499 ( .A(n16777), .ZN(n16630) );
  NAND3_X1 U15500 ( .A1(n13671), .A2(n13685), .A3(n13684), .ZN(P2_U2824) );
  INV_X1 U15501 ( .A(n20186), .ZN(n20194) );
  NOR2_X1 U15502 ( .A1(n16258), .A2(n20194), .ZN(n13703) );
  OR2_X1 U15503 ( .A1(n13690), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13693) );
  NAND2_X1 U15504 ( .A1(n20182), .A2(n13691), .ZN(n16333) );
  NAND3_X1 U15505 ( .A1(n10999), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n16333), .ZN(n13692) );
  OAI21_X1 U15506 ( .B1(n11000), .B2(n13693), .A(n13692), .ZN(n13695) );
  MUX2_X1 U15507 ( .A(n21580), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n12866), .Z(n13694) );
  NAND2_X1 U15508 ( .A1(n13695), .A2(n13694), .ZN(n13697) );
  XNOR2_X1 U15509 ( .A(n13697), .B(n13696), .ZN(n16431) );
  NAND2_X1 U15510 ( .A1(n21585), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n16426) );
  OAI21_X1 U15511 ( .B1(n20155), .B2(n16091), .A(n16426), .ZN(n13700) );
  INV_X1 U15512 ( .A(n16097), .ZN(n13698) );
  NOR2_X1 U15513 ( .A1(n13698), .A2(n20200), .ZN(n13699) );
  OR2_X1 U15514 ( .A1(n13703), .A2(n13702), .ZN(P1_U2971) );
  NAND2_X1 U15515 ( .A1(n13707), .A2(n13706), .ZN(n13708) );
  NAND2_X1 U15516 ( .A1(n13714), .A2(n13708), .ZN(n18804) );
  INV_X1 U15517 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17036) );
  NOR2_X1 U15518 ( .A1(n13709), .A2(n17036), .ZN(n16816) );
  NAND2_X1 U15519 ( .A1(n13709), .A2(n17036), .ZN(n16817) );
  XNOR2_X1 U15520 ( .A(n13714), .B(n11058), .ZN(n18815) );
  AOI21_X1 U15521 ( .B1(n18815), .B2(n13735), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16805) );
  INV_X1 U15522 ( .A(n13715), .ZN(n13718) );
  INV_X1 U15523 ( .A(n13716), .ZN(n13717) );
  NAND2_X1 U15524 ( .A1(n13718), .A2(n13717), .ZN(n13719) );
  NAND2_X1 U15525 ( .A1(n13722), .A2(n13719), .ZN(n16611) );
  NAND2_X1 U15526 ( .A1(n13720), .A2(n16061), .ZN(n13723) );
  NAND2_X1 U15527 ( .A1(n18838), .A2(n12190), .ZN(n13727) );
  XNOR2_X1 U15528 ( .A(n13727), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15980) );
  NOR2_X1 U15529 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13726) );
  NAND3_X1 U15530 ( .A1(n18828), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n12190), .ZN(n13725) );
  AND2_X1 U15531 ( .A1(n12190), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13724) );
  NAND2_X1 U15532 ( .A1(n18815), .A2(n13724), .ZN(n16803) );
  AND2_X1 U15533 ( .A1(n13725), .A2(n16803), .ZN(n14497) );
  NAND2_X1 U15534 ( .A1(n13730), .A2(n13729), .ZN(n16784) );
  XOR2_X1 U15535 ( .A(n13732), .B(n13731), .Z(n18854) );
  NAND2_X1 U15536 ( .A1(n18854), .A2(n12190), .ZN(n13733) );
  INV_X1 U15537 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17004) );
  NAND2_X1 U15538 ( .A1(n13733), .A2(n17004), .ZN(n16783) );
  NAND2_X1 U15539 ( .A1(n16784), .A2(n16783), .ZN(n16036) );
  INV_X1 U15540 ( .A(n13733), .ZN(n13734) );
  NAND2_X1 U15541 ( .A1(n13734), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16782) );
  NAND2_X1 U15542 ( .A1(n16036), .A2(n16782), .ZN(n13740) );
  AOI21_X1 U15543 ( .B1(n13737), .B2(n13735), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16035) );
  AND2_X1 U15544 ( .A1(n12190), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13736) );
  NAND2_X1 U15545 ( .A1(n13737), .A2(n13736), .ZN(n16034) );
  INV_X1 U15546 ( .A(n16034), .ZN(n13738) );
  NOR2_X1 U15547 ( .A1(n16035), .A2(n13738), .ZN(n13739) );
  OR2_X1 U15548 ( .A1(n18901), .A2(n15313), .ZN(n13742) );
  AOI21_X1 U15549 ( .B1(n13743), .B2(n13742), .A(n13741), .ZN(n15329) );
  NAND2_X1 U15550 ( .A1(n15329), .A2(n18592), .ZN(n18917) );
  NAND2_X1 U15551 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n17676) );
  NAND2_X1 U15552 ( .A1(n19459), .A2(n17676), .ZN(n18591) );
  OR2_X1 U15553 ( .A1(n18591), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13744) );
  AND2_X1 U15554 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n17324) );
  INV_X1 U15555 ( .A(n14116), .ZN(n15342) );
  NAND2_X1 U15556 ( .A1(n21819), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13745) );
  NAND2_X1 U15557 ( .A1(n15342), .A2(n13745), .ZN(n17660) );
  NOR2_X1 U15558 ( .A1(n16970), .A2(n17763), .ZN(n15999) );
  AOI21_X1 U15559 ( .B1(n17661), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15999), .ZN(n13746) );
  OAI21_X1 U15560 ( .B1(n17631), .B2(n13747), .A(n13746), .ZN(n13748) );
  NAND2_X1 U15561 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14515) );
  AND2_X2 U15562 ( .A1(n14498), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14499) );
  NAND2_X2 U15563 ( .A1(n14499), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16788) );
  NOR2_X2 U15564 ( .A1(n16788), .A2(n17004), .ZN(n16787) );
  AND3_X1 U15565 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15995) );
  AND2_X1 U15566 ( .A1(n15995), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16041) );
  NAND2_X1 U15567 ( .A1(n14498), .A2(n16041), .ZN(n16045) );
  BUF_X4 U15568 ( .A(n13839), .Z(n18045) );
  AOI22_X1 U15569 ( .A1(n18031), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18045), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13756) );
  INV_X1 U15570 ( .A(n13841), .ZN(n17984) );
  INV_X2 U15571 ( .A(n17984), .ZN(n18055) );
  NOR2_X2 U15572 ( .A1(n13761), .A2(n21022), .ZN(n13848) );
  AOI22_X1 U15573 ( .A1(n18055), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13755) );
  AOI22_X1 U15574 ( .A1(n18025), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10956), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13754) );
  NOR3_X1 U15575 ( .A1(n21020), .A2(n21001), .A3(n21021), .ZN(n13752) );
  INV_X1 U15576 ( .A(n13752), .ZN(n13801) );
  AOI22_X1 U15577 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17998), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13753) );
  NAND4_X1 U15578 ( .A1(n13756), .A2(n13755), .A3(n13754), .A4(n13753), .ZN(
        n13767) );
  NOR2_X2 U15579 ( .A1(n13759), .A2(n21022), .ZN(n13837) );
  CLKBUF_X3 U15580 ( .A(n13837), .Z(n18054) );
  AOI22_X1 U15581 ( .A1(n10957), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18054), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13765) );
  NOR2_X4 U15582 ( .A1(n13760), .A2(n20343), .ZN(n13919) );
  INV_X2 U15583 ( .A(n15053), .ZN(n18033) );
  AOI22_X1 U15584 ( .A1(n18046), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17890), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13764) );
  AOI22_X1 U15585 ( .A1(n18047), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13763) );
  AOI22_X1 U15586 ( .A1(n10967), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18032), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13762) );
  NAND4_X1 U15587 ( .A1(n13765), .A2(n13764), .A3(n13763), .A4(n13762), .ZN(
        n13766) );
  AOI22_X1 U15588 ( .A1(n18046), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18045), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13771) );
  AOI22_X1 U15589 ( .A1(n18047), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13770) );
  AOI22_X1 U15590 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17998), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13769) );
  AOI22_X1 U15591 ( .A1(n18025), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13835), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13768) );
  NAND4_X1 U15592 ( .A1(n13771), .A2(n13770), .A3(n13769), .A4(n13768), .ZN(
        n13777) );
  AOI22_X1 U15593 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18054), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13775) );
  AOI22_X1 U15594 ( .A1(n18055), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18032), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13774) );
  AOI22_X1 U15595 ( .A1(n18031), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13773) );
  AOI22_X1 U15596 ( .A1(n17909), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17890), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13772) );
  NAND4_X1 U15597 ( .A1(n13775), .A2(n13774), .A3(n13773), .A4(n13772), .ZN(
        n13776) );
  AOI22_X1 U15598 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13919), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13782) );
  AOI22_X1 U15599 ( .A1(n18031), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13757), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13781) );
  AOI22_X1 U15600 ( .A1(n13840), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18056), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13780) );
  AOI22_X1 U15601 ( .A1(n18055), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18045), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13779) );
  NAND4_X1 U15602 ( .A1(n13782), .A2(n13781), .A3(n13780), .A4(n13779), .ZN(
        n13788) );
  AOI22_X1 U15603 ( .A1(n18034), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13786) );
  AOI22_X1 U15604 ( .A1(n11010), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13848), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13785) );
  AOI22_X1 U15605 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17865), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13784) );
  AOI22_X1 U15606 ( .A1(n20370), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13835), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13783) );
  NAND4_X1 U15607 ( .A1(n13786), .A2(n13785), .A3(n13784), .A4(n13783), .ZN(
        n13787) );
  AOI22_X1 U15608 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18056), .B1(
        n10960), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13794) );
  AOI22_X1 U15609 ( .A1(n18034), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13838), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13793) );
  AOI22_X1 U15610 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20370), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n13835), .ZN(n13792) );
  AOI22_X1 U15611 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n13752), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n18049), .ZN(n13791) );
  NAND4_X1 U15612 ( .A1(n13794), .A2(n13793), .A3(n13792), .A4(n13791), .ZN(
        n13800) );
  AOI22_X1 U15613 ( .A1(n13840), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n13757), .ZN(n13798) );
  AOI22_X1 U15614 ( .A1(n11010), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13919), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13797) );
  AOI22_X1 U15615 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n13841), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n18045), .ZN(n13796) );
  AOI22_X1 U15616 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n13848), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13795) );
  NAND4_X1 U15617 ( .A1(n13798), .A2(n13797), .A3(n13796), .A4(n13795), .ZN(
        n13799) );
  NOR2_X2 U15618 ( .A1(n13800), .A2(n13799), .ZN(n13851) );
  AOI22_X1 U15619 ( .A1(n17909), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13811) );
  AOI22_X1 U15620 ( .A1(n18034), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18045), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13810) );
  INV_X1 U15621 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17778) );
  AOI22_X1 U15622 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18013), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13802) );
  OAI21_X1 U15623 ( .B1(n13801), .B2(n17778), .A(n13802), .ZN(n13808) );
  AOI22_X1 U15624 ( .A1(n11010), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18047), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13806) );
  AOI22_X1 U15625 ( .A1(n18055), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18032), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13805) );
  AOI22_X1 U15626 ( .A1(n18046), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13804) );
  AOI22_X1 U15627 ( .A1(n18033), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13803) );
  NAND4_X1 U15628 ( .A1(n13806), .A2(n13805), .A3(n13804), .A4(n13803), .ZN(
        n13807) );
  AOI211_X1 U15629 ( .C1(n18025), .C2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A(
        n13808), .B(n13807), .ZN(n13809) );
  NAND3_X1 U15630 ( .A1(n13811), .A2(n13810), .A3(n13809), .ZN(n13856) );
  NAND2_X1 U15631 ( .A1(n14023), .A2(n13856), .ZN(n13858) );
  AOI22_X1 U15632 ( .A1(n18046), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13822) );
  AOI22_X1 U15633 ( .A1(n18055), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13821) );
  AOI22_X1 U15634 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13835), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13812) );
  OAI21_X1 U15635 ( .B1(n13801), .B2(n17835), .A(n13812), .ZN(n13819) );
  AOI22_X1 U15636 ( .A1(n17909), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11010), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13817) );
  AOI22_X1 U15637 ( .A1(n18034), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18056), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13816) );
  AOI22_X1 U15638 ( .A1(n18045), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13815) );
  AOI22_X1 U15639 ( .A1(n18047), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17890), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13814) );
  NAND4_X1 U15640 ( .A1(n13817), .A2(n13816), .A3(n13815), .A4(n13814), .ZN(
        n13818) );
  AOI211_X1 U15641 ( .C1(n18025), .C2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A(
        n13819), .B(n13818), .ZN(n13820) );
  NAND3_X1 U15642 ( .A1(n13822), .A2(n13821), .A3(n13820), .ZN(n14011) );
  AOI22_X1 U15643 ( .A1(n18046), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18045), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13832) );
  AOI22_X1 U15644 ( .A1(n10971), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n18056), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13831) );
  AOI22_X1 U15645 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13835), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13823) );
  OAI21_X1 U15646 ( .B1(n13801), .B2(n17818), .A(n13823), .ZN(n13829) );
  AOI22_X1 U15647 ( .A1(n17909), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17890), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13827) );
  AOI22_X1 U15648 ( .A1(n10967), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18047), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13826) );
  AOI22_X1 U15649 ( .A1(n18055), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13825) );
  AOI22_X1 U15650 ( .A1(n18034), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13824) );
  NAND4_X1 U15651 ( .A1(n13827), .A2(n13826), .A3(n13825), .A4(n13824), .ZN(
        n13828) );
  AOI211_X1 U15652 ( .C1(n18025), .C2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n13829), .B(n13828), .ZN(n13830) );
  INV_X1 U15653 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21398) );
  INV_X1 U15654 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n21213) );
  INV_X1 U15655 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n21412) );
  NOR2_X1 U15656 ( .A1(n21435), .A2(n21412), .ZN(n21158) );
  NAND3_X1 U15657 ( .A1(n21158), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21166) );
  INV_X1 U15658 ( .A(n21166), .ZN(n18130) );
  NAND2_X1 U15659 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18130), .ZN(
        n21196) );
  INV_X1 U15660 ( .A(n21196), .ZN(n21180) );
  NAND2_X1 U15661 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n21180), .ZN(
        n21205) );
  NOR2_X1 U15662 ( .A1(n21213), .A2(n21205), .ZN(n21366) );
  INV_X1 U15663 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21135) );
  OAI21_X1 U15664 ( .B1(n13833), .B2(n14085), .A(n21308), .ZN(n13868) );
  INV_X1 U15665 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18411) );
  XNOR2_X1 U15666 ( .A(n14011), .B(n13834), .ZN(n13861) );
  INV_X1 U15667 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17785) );
  AOI22_X1 U15668 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13835), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13836) );
  OAI21_X1 U15669 ( .B1(n13801), .B2(n17785), .A(n13836), .ZN(n13847) );
  AOI22_X1 U15670 ( .A1(n13837), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13838), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13846) );
  AOI22_X1 U15671 ( .A1(n13840), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17908), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13845) );
  INV_X4 U15672 ( .A(n17984), .ZN(n17920) );
  AOI22_X1 U15673 ( .A1(n17920), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13842), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13844) );
  AOI22_X1 U15674 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18032), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13843) );
  AOI22_X1 U15675 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18033), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13850) );
  AOI22_X1 U15676 ( .A1(n13919), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13849) );
  XNOR2_X1 U15677 ( .A(n13851), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18453) );
  INV_X1 U15678 ( .A(n13851), .ZN(n20977) );
  INV_X1 U15679 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20995) );
  NOR2_X1 U15680 ( .A1(n20977), .A2(n20995), .ZN(n13852) );
  INV_X1 U15681 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21083) );
  XNOR2_X2 U15682 ( .A(n20977), .B(n14012), .ZN(n13853) );
  NOR2_X1 U15683 ( .A1(n21083), .A2(n13853), .ZN(n13854) );
  NOR2_X2 U15684 ( .A1(n18447), .A2(n13854), .ZN(n13855) );
  INV_X1 U15685 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21097) );
  NOR2_X1 U15686 ( .A1(n13855), .A2(n21097), .ZN(n13857) );
  XNOR2_X1 U15687 ( .A(n13855), .B(n21097), .ZN(n18434) );
  INV_X1 U15688 ( .A(n13856), .ZN(n20845) );
  XOR2_X1 U15689 ( .A(n20845), .B(n14023), .Z(n18433) );
  NOR2_X1 U15690 ( .A1(n18434), .A2(n18433), .ZN(n18432) );
  NOR2_X1 U15691 ( .A1(n13857), .A2(n18432), .ZN(n18426) );
  INV_X1 U15692 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21100) );
  XNOR2_X1 U15693 ( .A(n20840), .B(n13858), .ZN(n13859) );
  XNOR2_X1 U15694 ( .A(n21100), .B(n13859), .ZN(n18425) );
  NOR2_X1 U15695 ( .A1(n21100), .A2(n13859), .ZN(n13860) );
  NOR2_X1 U15696 ( .A1(n13862), .A2(n13861), .ZN(n13863) );
  NOR2_X2 U15697 ( .A1(n18409), .A2(n13863), .ZN(n18396) );
  XOR2_X1 U15698 ( .A(n20832), .B(n13864), .Z(n13865) );
  XNOR2_X1 U15699 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n13865), .ZN(
        n18395) );
  NOR2_X1 U15700 ( .A1(n13867), .A2(n13868), .ZN(n13869) );
  NAND2_X1 U15701 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21308), .ZN(
        n13870) );
  NOR2_X1 U15702 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21308), .ZN(
        n18371) );
  NAND2_X1 U15703 ( .A1(n21366), .A2(n18339), .ZN(n13875) );
  INV_X1 U15704 ( .A(n18339), .ZN(n13874) );
  NOR3_X1 U15705 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18107) );
  NAND3_X1 U15706 ( .A1(n18107), .A2(n21213), .A3(n13871), .ZN(n13872) );
  NAND2_X1 U15707 ( .A1(n21435), .A2(n21412), .ZN(n18351) );
  NOR2_X1 U15708 ( .A1(n13872), .A2(n18351), .ZN(n13873) );
  INV_X1 U15709 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18315) );
  INV_X1 U15710 ( .A(n13875), .ZN(n13876) );
  NOR2_X1 U15711 ( .A1(n21398), .A2(n18315), .ZN(n21364) );
  INV_X1 U15712 ( .A(n21364), .ZN(n18086) );
  INV_X1 U15713 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18091) );
  NOR2_X1 U15714 ( .A1(n18086), .A2(n18091), .ZN(n18089) );
  INV_X1 U15715 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18181) );
  INV_X1 U15716 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18177) );
  NOR2_X1 U15717 ( .A1(n18181), .A2(n18177), .ZN(n21049) );
  NAND2_X1 U15718 ( .A1(n21049), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n18149) );
  INV_X1 U15719 ( .A(n18149), .ZN(n21222) );
  AND2_X1 U15720 ( .A1(n18089), .A2(n21222), .ZN(n18150) );
  NAND3_X1 U15721 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n18150), .ZN(n14009) );
  NAND2_X1 U15722 ( .A1(n21308), .A2(n18091), .ZN(n18176) );
  NOR2_X1 U15723 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18176), .ZN(
        n13878) );
  NAND2_X1 U15724 ( .A1(n13878), .A2(n18181), .ZN(n18163) );
  NOR2_X1 U15725 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18163), .ZN(
        n18154) );
  INV_X1 U15726 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21257) );
  NAND2_X1 U15727 ( .A1(n18154), .A2(n21257), .ZN(n18193) );
  OAI22_X1 U15728 ( .A1(n18121), .A2(n14009), .B1(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18193), .ZN(n13879) );
  NAND2_X1 U15729 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21329) );
  AND2_X1 U15730 ( .A1(n21222), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13880) );
  INV_X1 U15731 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n21246) );
  INV_X1 U15732 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21247) );
  AOI21_X1 U15733 ( .B1(n21246), .B2(n21247), .A(n18258), .ZN(n13881) );
  INV_X1 U15734 ( .A(n13881), .ZN(n13882) );
  INV_X1 U15735 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21306) );
  NAND2_X1 U15736 ( .A1(n13883), .A2(n21306), .ZN(n21315) );
  NOR2_X1 U15737 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18258), .ZN(
        n18247) );
  INV_X1 U15738 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14084) );
  NAND3_X1 U15739 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18258), .A3(
        n18248), .ZN(n21299) );
  INV_X1 U15740 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21288) );
  OAI33_X1 U15741 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n18291), .B1(n14084), .B2(
        n21299), .B3(n21288), .ZN(n13884) );
  INV_X1 U15742 ( .A(n14085), .ZN(n21297) );
  INV_X1 U15743 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15032) );
  AOI22_X1 U15744 ( .A1(n18046), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n18045), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13885) );
  OAI21_X1 U15745 ( .B1(n13961), .B2(n15032), .A(n13885), .ZN(n13891) );
  AOI22_X1 U15746 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13889) );
  AOI22_X1 U15747 ( .A1(n18033), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13888) );
  AOI22_X1 U15748 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17865), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13887) );
  AOI22_X1 U15749 ( .A1(n20370), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10956), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13886) );
  NAND4_X1 U15750 ( .A1(n13889), .A2(n13888), .A3(n13887), .A4(n13886), .ZN(
        n13890) );
  NOR2_X1 U15751 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n20337), .ZN(n21481) );
  NAND2_X1 U15752 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n21481), .ZN(n21500) );
  AOI21_X1 U15753 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n21020), .A(
        n14002), .ZN(n14006) );
  INV_X1 U15754 ( .A(n14006), .ZN(n13907) );
  OAI22_X1 U15755 ( .A1(n21001), .A2(n21450), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14001) );
  AOI22_X1 U15756 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n18968), .B2(n21006), .ZN(
        n13904) );
  OAI21_X1 U15757 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n21006), .A(
        n13896), .ZN(n13897) );
  OAI22_X1 U15758 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17316), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13897), .ZN(n13899) );
  NOR2_X1 U15759 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17316), .ZN(
        n13898) );
  NAND2_X1 U15760 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13897), .ZN(
        n13900) );
  AOI22_X1 U15761 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13899), .B1(
        n13898), .B2(n13900), .ZN(n13902) );
  NAND2_X1 U15762 ( .A1(n14001), .A2(n13902), .ZN(n13906) );
  AOI21_X1 U15763 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n13900), .A(
        n13899), .ZN(n13901) );
  OAI21_X1 U15764 ( .B1(n13905), .B2(n13904), .A(n13902), .ZN(n13903) );
  AOI21_X1 U15765 ( .B1(n13905), .B2(n13904), .A(n13903), .ZN(n14007) );
  AOI22_X1 U15766 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13912) );
  AOI22_X1 U15767 ( .A1(n18047), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18056), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13911) );
  AOI22_X1 U15768 ( .A1(n10956), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17865), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13910) );
  AOI22_X1 U15769 ( .A1(n20370), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18013), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13909) );
  NAND4_X1 U15770 ( .A1(n13912), .A2(n13911), .A3(n13910), .A4(n13909), .ZN(
        n13918) );
  AOI22_X1 U15771 ( .A1(n17909), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17890), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13916) );
  INV_X2 U15772 ( .A(n13961), .ZN(n17991) );
  AOI22_X1 U15773 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13919), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13915) );
  AOI22_X1 U15774 ( .A1(n17920), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13914) );
  AOI22_X1 U15775 ( .A1(n10967), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18045), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13913) );
  NAND4_X1 U15776 ( .A1(n13916), .A2(n13915), .A3(n13914), .A4(n13913), .ZN(
        n13917) );
  NAND2_X1 U15777 ( .A1(n20340), .A2(n19216), .ZN(n13990) );
  NAND2_X1 U15778 ( .A1(n19262), .A2(n20351), .ZN(n13989) );
  NAND2_X1 U15779 ( .A1(n13990), .A2(n13989), .ZN(n20275) );
  AOI22_X1 U15780 ( .A1(n18034), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n18046), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13923) );
  AOI22_X1 U15781 ( .A1(n18031), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13922) );
  AOI22_X1 U15782 ( .A1(n18025), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17998), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13921) );
  AOI22_X1 U15783 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13835), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13920) );
  NAND4_X1 U15784 ( .A1(n13923), .A2(n13922), .A3(n13921), .A4(n13920), .ZN(
        n13929) );
  AOI22_X1 U15785 ( .A1(n10957), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18056), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13927) );
  AOI22_X1 U15786 ( .A1(n10967), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13926) );
  AOI22_X1 U15787 ( .A1(n18055), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18047), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13925) );
  AOI22_X1 U15788 ( .A1(n18045), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17890), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13924) );
  NAND4_X1 U15789 ( .A1(n13927), .A2(n13926), .A3(n13925), .A4(n13924), .ZN(
        n13928) );
  AOI22_X1 U15790 ( .A1(n17909), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13933) );
  AOI22_X1 U15791 ( .A1(n11010), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13932) );
  AOI22_X1 U15792 ( .A1(n10956), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17865), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13931) );
  AOI22_X1 U15793 ( .A1(n20370), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13835), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13930) );
  NAND4_X1 U15794 ( .A1(n13933), .A2(n13932), .A3(n13931), .A4(n13930), .ZN(
        n13939) );
  AOI22_X1 U15795 ( .A1(n17920), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17890), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13937) );
  AOI22_X1 U15796 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13936) );
  AOI22_X1 U15797 ( .A1(n18046), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18056), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13935) );
  AOI22_X1 U15798 ( .A1(n18047), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18045), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13934) );
  NAND4_X1 U15799 ( .A1(n13937), .A2(n13936), .A3(n13935), .A4(n13934), .ZN(
        n13938) );
  INV_X1 U15800 ( .A(n17389), .ZN(n13981) );
  NOR2_X1 U15801 ( .A1(n13982), .A2(n13981), .ZN(n14068) );
  AOI22_X1 U15802 ( .A1(n18047), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13919), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13949) );
  AOI22_X1 U15803 ( .A1(n17920), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17890), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13948) );
  AOI22_X1 U15804 ( .A1(n18045), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13940) );
  OAI21_X1 U15805 ( .B1(n13961), .B2(n17835), .A(n13940), .ZN(n13946) );
  AOI22_X1 U15806 ( .A1(n10967), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18054), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13944) );
  AOI22_X1 U15807 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13943) );
  AOI22_X1 U15808 ( .A1(n10956), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13835), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13942) );
  AOI22_X1 U15809 ( .A1(n20370), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17865), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13941) );
  NAND4_X1 U15810 ( .A1(n13944), .A2(n13943), .A3(n13942), .A4(n13941), .ZN(
        n13945) );
  AOI211_X1 U15811 ( .C1(n13840), .C2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n13946), .B(n13945), .ZN(n13947) );
  NAND3_X1 U15812 ( .A1(n13949), .A2(n13948), .A3(n13947), .ZN(n20855) );
  AOI22_X1 U15813 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13953) );
  AOI22_X1 U15814 ( .A1(n18033), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18056), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13952) );
  AOI22_X1 U15815 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17865), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13951) );
  AOI22_X1 U15816 ( .A1(n20370), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10956), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13950) );
  NAND4_X1 U15817 ( .A1(n13953), .A2(n13952), .A3(n13951), .A4(n13950), .ZN(
        n13959) );
  AOI22_X1 U15818 ( .A1(n17920), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18054), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13957) );
  AOI22_X1 U15819 ( .A1(n18045), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13956) );
  AOI22_X1 U15820 ( .A1(n13840), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18047), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13955) );
  AOI22_X1 U15821 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n18046), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13954) );
  NAND4_X1 U15822 ( .A1(n13957), .A2(n13956), .A3(n13955), .A4(n13954), .ZN(
        n13958) );
  NOR2_X1 U15823 ( .A1(n19055), .A2(n13982), .ZN(n14059) );
  AOI22_X1 U15824 ( .A1(n17920), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17890), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13970) );
  AOI22_X1 U15825 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13969) );
  AOI22_X1 U15826 ( .A1(n18045), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18056), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13960) );
  OAI21_X1 U15827 ( .B1(n13961), .B2(n17818), .A(n13960), .ZN(n13967) );
  AOI22_X1 U15828 ( .A1(n18047), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13848), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13965) );
  AOI22_X1 U15829 ( .A1(n13840), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10967), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13964) );
  AOI22_X1 U15830 ( .A1(n20370), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17865), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13963) );
  AOI22_X1 U15831 ( .A1(n10956), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13835), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13962) );
  NAND4_X1 U15832 ( .A1(n13965), .A2(n13964), .A3(n13963), .A4(n13962), .ZN(
        n13966) );
  AOI22_X1 U15833 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n18045), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13974) );
  AOI22_X1 U15834 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13973) );
  AOI22_X1 U15835 ( .A1(n10956), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13835), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13972) );
  AOI22_X1 U15836 ( .A1(n20370), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17865), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13971) );
  NAND4_X1 U15837 ( .A1(n13974), .A2(n13973), .A3(n13972), .A4(n13971), .ZN(
        n13980) );
  AOI22_X1 U15838 ( .A1(n17909), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13919), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13978) );
  AOI22_X1 U15839 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18056), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13977) );
  AOI22_X1 U15840 ( .A1(n17920), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13976) );
  AOI22_X1 U15841 ( .A1(n18047), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17890), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13975) );
  NAND4_X1 U15842 ( .A1(n13978), .A2(n13977), .A3(n13976), .A4(n13975), .ZN(
        n13979) );
  NOR2_X1 U15843 ( .A1(n13994), .A2(n13999), .ZN(n13984) );
  NOR2_X1 U15844 ( .A1(n17389), .A2(n20856), .ZN(n13983) );
  NAND2_X1 U15845 ( .A1(n13984), .A2(n13983), .ZN(n17299) );
  NAND3_X1 U15846 ( .A1(n19262), .A2(n19133), .A3(n20801), .ZN(n13993) );
  NAND2_X1 U15847 ( .A1(n20855), .A2(n20856), .ZN(n14055) );
  NOR3_X2 U15848 ( .A1(n13981), .A2(n13993), .A3(n14055), .ZN(n14074) );
  NAND2_X1 U15849 ( .A1(n14074), .A2(n13982), .ZN(n14062) );
  INV_X1 U15850 ( .A(n20804), .ZN(n20992) );
  OAI21_X1 U15851 ( .B1(n20340), .B2(n13982), .A(n20992), .ZN(n14069) );
  INV_X1 U15852 ( .A(n13983), .ZN(n21005) );
  NAND3_X1 U15853 ( .A1(n14060), .A2(n14069), .A3(n21005), .ZN(n13991) );
  NAND3_X1 U15854 ( .A1(n13984), .A2(n19055), .A3(n13991), .ZN(n13985) );
  INV_X1 U15855 ( .A(n13985), .ZN(n13986) );
  NAND2_X1 U15856 ( .A1(n19174), .A2(n19133), .ZN(n21004) );
  NOR2_X2 U15857 ( .A1(n21440), .A2(n13988), .ZN(n14000) );
  AND2_X1 U15858 ( .A1(n20801), .A2(n14055), .ZN(n13997) );
  NAND2_X1 U15859 ( .A1(n19174), .A2(n13989), .ZN(n14064) );
  NOR2_X1 U15860 ( .A1(n20971), .A2(n20804), .ZN(n20803) );
  INV_X1 U15861 ( .A(n13991), .ZN(n13992) );
  OAI21_X1 U15862 ( .B1(n19133), .B2(n13994), .A(n13993), .ZN(n13995) );
  NAND2_X2 U15863 ( .A1(n14000), .A2(n17318), .ZN(n21231) );
  NAND2_X1 U15864 ( .A1(n20351), .A2(n13999), .ZN(n21002) );
  NAND2_X1 U15865 ( .A1(n21004), .A2(n21002), .ZN(n14076) );
  NOR2_X4 U15866 ( .A1(n20351), .A2(n21334), .ZN(n21343) );
  XNOR2_X1 U15867 ( .A(n14002), .B(n14001), .ZN(n14004) );
  AOI21_X1 U15868 ( .B1(n14007), .B2(n14006), .A(n21471), .ZN(n14054) );
  INV_X1 U15869 ( .A(n14054), .ZN(n21443) );
  NOR2_X4 U15870 ( .A1(n19216), .A2(n21505), .ZN(n18457) );
  NAND2_X1 U15871 ( .A1(n11030), .A2(n18379), .ZN(n14053) );
  NAND2_X1 U15872 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21268) );
  NOR2_X1 U15873 ( .A1(n21268), .A2(n21288), .ZN(n21274) );
  NAND2_X1 U15874 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n21274), .ZN(
        n14078) );
  INV_X1 U15875 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21423) );
  NAND2_X1 U15876 ( .A1(n21170), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18321) );
  INV_X1 U15877 ( .A(n21208), .ZN(n18113) );
  NOR2_X4 U15878 ( .A1(n18113), .A2(n21213), .ZN(n21207) );
  INV_X1 U15879 ( .A(n14009), .ZN(n14040) );
  INV_X1 U15880 ( .A(n21320), .ZN(n18206) );
  NAND2_X1 U15881 ( .A1(n18206), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18219) );
  XNOR2_X1 U15882 ( .A(n14010), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14086) );
  NAND2_X2 U15883 ( .A1(n21297), .A2(n18457), .ZN(n18236) );
  OR2_X1 U15884 ( .A1(n14086), .A2(n18236), .ZN(n14052) );
  INV_X1 U15885 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14041) );
  INV_X1 U15886 ( .A(n14011), .ZN(n20836) );
  NOR2_X1 U15887 ( .A1(n13851), .A2(n20991), .ZN(n14027) );
  INV_X1 U15888 ( .A(n20840), .ZN(n14013) );
  NAND2_X1 U15889 ( .A1(n14019), .A2(n14013), .ZN(n14017) );
  NOR2_X1 U15890 ( .A1(n20836), .A2(n14017), .ZN(n14016) );
  INV_X1 U15891 ( .A(n20832), .ZN(n14014) );
  NAND2_X1 U15892 ( .A1(n14016), .A2(n14014), .ZN(n14015) );
  NOR2_X1 U15893 ( .A1(n21297), .A2(n14015), .ZN(n14038) );
  XNOR2_X1 U15894 ( .A(n14085), .B(n14015), .ZN(n18383) );
  XNOR2_X1 U15895 ( .A(n20832), .B(n14016), .ZN(n14032) );
  XOR2_X1 U15896 ( .A(n20836), .B(n14017), .Z(n14018) );
  NAND2_X1 U15897 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14018), .ZN(
        n14031) );
  XNOR2_X1 U15898 ( .A(n18411), .B(n14018), .ZN(n18408) );
  XNOR2_X1 U15899 ( .A(n20840), .B(n14019), .ZN(n14020) );
  NAND2_X1 U15900 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n14020), .ZN(
        n14030) );
  XNOR2_X1 U15901 ( .A(n21100), .B(n14020), .ZN(n18420) );
  XOR2_X1 U15902 ( .A(n20845), .B(n14022), .Z(n14021) );
  NAND2_X1 U15903 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n14021), .ZN(
        n14029) );
  XNOR2_X1 U15904 ( .A(n21097), .B(n14021), .ZN(n18437) );
  AOI21_X1 U15905 ( .B1(n14024), .B2(n14023), .A(n14022), .ZN(n14025) );
  INV_X1 U15906 ( .A(n14025), .ZN(n14026) );
  NAND2_X1 U15907 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14026), .ZN(
        n14028) );
  INV_X1 U15908 ( .A(n18453), .ZN(n18455) );
  INV_X1 U15909 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21071) );
  NAND2_X1 U15910 ( .A1(n20991), .A2(n21071), .ZN(n18461) );
  NOR2_X1 U15911 ( .A1(n18455), .A2(n18461), .ZN(n18454) );
  AOI211_X1 U15912 ( .C1(n13851), .C2(n20995), .A(n14027), .B(n18454), .ZN(
        n18444) );
  NAND2_X1 U15913 ( .A1(n14029), .A2(n18435), .ZN(n18419) );
  NAND2_X1 U15914 ( .A1(n14032), .A2(n14033), .ZN(n14034) );
  XOR2_X1 U15915 ( .A(n14033), .B(n14032), .Z(n18402) );
  NAND2_X1 U15916 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18402), .ZN(
        n18401) );
  NAND2_X1 U15917 ( .A1(n14038), .A2(n14035), .ZN(n14039) );
  NAND2_X1 U15918 ( .A1(n18383), .A2(n18384), .ZN(n18382) );
  NAND2_X1 U15919 ( .A1(n14038), .A2(n14037), .ZN(n14036) );
  OAI211_X1 U15920 ( .C1(n14038), .C2(n14037), .A(n18382), .B(n14036), .ZN(
        n18370) );
  NAND2_X1 U15921 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18370), .ZN(
        n18369) );
  NAND2_X1 U15922 ( .A1(n14040), .A2(n21360), .ZN(n21319) );
  INV_X1 U15923 ( .A(n21275), .ZN(n21248) );
  OR2_X1 U15924 ( .A1(n21248), .A2(n14078), .ZN(n14042) );
  XNOR2_X1 U15925 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n14042), .ZN(
        n14090) );
  NOR2_X2 U15926 ( .A1(n20351), .A2(n21505), .ZN(n18423) );
  NAND2_X1 U15927 ( .A1(n14090), .A2(n18423), .ZN(n14051) );
  NAND2_X1 U15928 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18215) );
  NAND2_X1 U15929 ( .A1(n18373), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n20451) );
  NAND2_X1 U15930 ( .A1(n20480), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n20492) );
  INV_X1 U15931 ( .A(n20492), .ZN(n14043) );
  NAND2_X1 U15932 ( .A1(n18428), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18412) );
  NAND2_X1 U15933 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18137) );
  INV_X1 U15934 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n20545) );
  INV_X1 U15935 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n20554) );
  NOR2_X1 U15936 ( .A1(n20545), .A2(n20554), .ZN(n20562) );
  INV_X1 U15937 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18187) );
  NOR2_X4 U15938 ( .A1(n18186), .A2(n18187), .ZN(n18185) );
  NAND2_X1 U15939 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18157) );
  INV_X1 U15940 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n18254) );
  INV_X1 U15941 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n20736) );
  NAND2_X1 U15942 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18076) );
  NAND2_X1 U15943 ( .A1(n21488), .A2(n18076), .ZN(n18079) );
  INV_X1 U15944 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n20997) );
  NOR2_X1 U15945 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n21491) );
  NAND2_X1 U15946 ( .A1(n21491), .A2(n21488), .ZN(n18075) );
  NOR2_X1 U15947 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18075), .ZN(n14092) );
  INV_X1 U15948 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n20761) );
  NOR2_X1 U15949 ( .A1(n21379), .A2(n20761), .ZN(n14093) );
  INV_X1 U15950 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14044) );
  NOR2_X1 U15951 ( .A1(n11050), .A2(n20519), .ZN(n18102) );
  NAND2_X1 U15952 ( .A1(n20562), .A2(n18102), .ZN(n18308) );
  NOR2_X1 U15953 ( .A1(n18307), .A2(n18308), .ZN(n18080) );
  NAND2_X1 U15954 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18080), .ZN(
        n20594) );
  NOR2_X1 U15955 ( .A1(n14044), .A2(n20594), .ZN(n20617) );
  NAND2_X1 U15956 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n20617), .ZN(
        n18166) );
  NOR2_X1 U15957 ( .A1(n18157), .A2(n18166), .ZN(n18203) );
  NAND2_X1 U15958 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18203), .ZN(
        n18214) );
  NOR2_X1 U15959 ( .A1(n18215), .A2(n18214), .ZN(n18268) );
  NAND2_X1 U15960 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18268), .ZN(
        n18242) );
  NOR2_X1 U15961 ( .A1(n18254), .A2(n18242), .ZN(n18239) );
  NAND2_X1 U15962 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18239), .ZN(
        n18288) );
  NOR2_X1 U15963 ( .A1(n20736), .A2(n18288), .ZN(n14045) );
  INV_X1 U15964 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n21352) );
  NOR2_X1 U15965 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n21352), .ZN(n18196) );
  INV_X1 U15966 ( .A(n21491), .ZN(n20276) );
  AOI21_X1 U15967 ( .B1(n20276), .B2(n18076), .A(n21490), .ZN(n17388) );
  NOR3_X2 U15968 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n21823), .ZN(n18979) );
  OAI21_X1 U15969 ( .B1(n11129), .B2(n18305), .A(n19054), .ZN(n18238) );
  NAND2_X1 U15970 ( .A1(n14045), .A2(n18238), .ZN(n18279) );
  XOR2_X1 U15971 ( .A(n11131), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n14048) );
  NOR2_X1 U15972 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18305), .ZN(
        n18298) );
  INV_X1 U15973 ( .A(n14045), .ZN(n14046) );
  AOI22_X1 U15974 ( .A1(n18196), .A2(n18296), .B1(n19215), .B2(n14046), .ZN(
        n14047) );
  NAND2_X1 U15975 ( .A1(n14047), .A2(n11018), .ZN(n18290) );
  NOR2_X1 U15976 ( .A1(n18298), .A2(n18290), .ZN(n18278) );
  OAI22_X1 U15977 ( .A1(n18279), .A2(n14048), .B1(n18278), .B2(n11131), .ZN(
        n14049) );
  AOI211_X1 U15978 ( .C1(n20592), .C2(n18297), .A(n14093), .B(n14049), .ZN(
        n14050) );
  NAND2_X1 U15979 ( .A1(n14053), .A2(n11251), .ZN(P3_U2799) );
  NAND2_X1 U15980 ( .A1(n14054), .A2(n20351), .ZN(n14056) );
  OAI22_X1 U15981 ( .A1(n14057), .A2(n14056), .B1(n21445), .B2(n14055), .ZN(
        n14072) );
  XOR2_X1 U15982 ( .A(n19216), .B(n19174), .Z(n14058) );
  INV_X1 U15983 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n21871) );
  INV_X1 U15984 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n21870) );
  NAND2_X2 U15985 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n21881), .ZN(n18561) );
  AOI211_X1 U15986 ( .C1(n21871), .C2(n21870), .A(n18571), .B(
        P3_STATE_REG_0__SCAN_IN), .ZN(n20348) );
  NAND2_X1 U15987 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n21478) );
  OAI21_X1 U15988 ( .B1(n14058), .B2(n20348), .A(n21478), .ZN(n21468) );
  NOR3_X1 U15989 ( .A1(n14059), .A2(n21471), .A3(n21468), .ZN(n14071) );
  OAI211_X1 U15990 ( .C1(n20804), .C2(n17389), .A(n14061), .B(n14060), .ZN(
        n14063) );
  OAI21_X1 U15991 ( .B1(n14064), .B2(n14063), .A(n14062), .ZN(n14065) );
  INV_X1 U15992 ( .A(n14065), .ZN(n14066) );
  AOI211_X1 U15993 ( .C1(n14069), .C2(n14068), .A(n14067), .B(n14066), .ZN(
        n14070) );
  INV_X1 U15994 ( .A(n14070), .ZN(n17303) );
  AOI211_X1 U15995 ( .C1(n19174), .C2(n14072), .A(n14071), .B(n17303), .ZN(
        n14073) );
  AOI221_X4 U15996 ( .B1(n17389), .B2(n14073), .C1(n21445), .C2(n14073), .A(
        n21500), .ZN(n21403) );
  NAND2_X1 U15997 ( .A1(n11030), .A2(n21432), .ZN(n14097) );
  NAND3_X1 U15998 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21235) );
  NOR2_X1 U15999 ( .A1(n11247), .A2(n21235), .ZN(n18237) );
  NAND2_X1 U16000 ( .A1(n21366), .A2(n18089), .ZN(n21043) );
  INV_X1 U16001 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21132) );
  NAND2_X1 U16002 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21108) );
  NOR2_X1 U16003 ( .A1(n18411), .A2(n21108), .ZN(n14077) );
  OAI21_X1 U16004 ( .B1(n20995), .B2(n21071), .A(n21083), .ZN(n21086) );
  NAND2_X1 U16005 ( .A1(n14077), .A2(n21086), .ZN(n21109) );
  NOR2_X1 U16006 ( .A1(n21132), .A2(n21109), .ZN(n21138) );
  NAND3_X1 U16007 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n21138), .ZN(n21194) );
  NOR2_X1 U16008 ( .A1(n21043), .A2(n21194), .ZN(n14081) );
  NOR2_X1 U16009 ( .A1(n21003), .A2(n14074), .ZN(n21029) );
  INV_X1 U16010 ( .A(n21029), .ZN(n14075) );
  NOR2_X1 U16011 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21231), .ZN(
        n21063) );
  NOR2_X1 U16012 ( .A1(n21372), .A2(n21063), .ZN(n21085) );
  INV_X1 U16013 ( .A(n14077), .ZN(n21133) );
  NAND2_X1 U16014 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21089) );
  NOR2_X1 U16015 ( .A1(n21133), .A2(n21089), .ZN(n21111) );
  NAND2_X1 U16016 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21111), .ZN(
        n21136) );
  NOR2_X1 U16017 ( .A1(n21135), .A2(n21136), .ZN(n21426) );
  NAND2_X1 U16018 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21426), .ZN(
        n21195) );
  NOR2_X1 U16019 ( .A1(n21043), .A2(n21195), .ZN(n21050) );
  AOI22_X1 U16020 ( .A1(n21368), .A2(n14081), .B1(n21085), .B2(n21050), .ZN(
        n21042) );
  NOR2_X1 U16021 ( .A1(n21042), .A2(n18149), .ZN(n21228) );
  NAND2_X1 U16022 ( .A1(n18237), .A2(n21228), .ZN(n21270) );
  NOR3_X1 U16023 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n14078), .A3(
        n21270), .ZN(n14089) );
  INV_X1 U16024 ( .A(n21274), .ZN(n18281) );
  INV_X1 U16025 ( .A(n21217), .ZN(n21422) );
  AND2_X1 U16026 ( .A1(n21050), .A2(n21222), .ZN(n21216) );
  NAND2_X1 U16027 ( .A1(n21216), .A2(n18237), .ZN(n14080) );
  NAND2_X1 U16028 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14079) );
  AOI222_X1 U16029 ( .A1(n21422), .A2(n14080), .B1(n21422), .B2(n14079), .C1(
        n14080), .C2(n21231), .ZN(n21278) );
  NAND2_X1 U16030 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21233) );
  NOR2_X1 U16031 ( .A1(n11247), .A2(n21233), .ZN(n21259) );
  INV_X1 U16032 ( .A(n21259), .ZN(n14083) );
  INV_X1 U16033 ( .A(n14081), .ZN(n21045) );
  NOR2_X1 U16034 ( .A1(n21045), .A2(n18149), .ZN(n14082) );
  INV_X1 U16035 ( .A(n21368), .ZN(n21438) );
  AOI21_X1 U16036 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n14082), .A(
        n21438), .ZN(n21323) );
  AOI21_X1 U16037 ( .B1(n21368), .B2(n14083), .A(n21323), .ZN(n21258) );
  NAND2_X1 U16038 ( .A1(n21278), .A2(n21258), .ZN(n21302) );
  AOI211_X1 U16039 ( .C1(n21334), .C2(n18281), .A(n21302), .B(n14084), .ZN(
        n21286) );
  NAND2_X1 U16040 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n21334), .ZN(
        n14087) );
  OAI22_X1 U16041 ( .A1(n21286), .A2(n14087), .B1(n21361), .B2(n14086), .ZN(
        n14088) );
  AOI211_X1 U16042 ( .C1(n14090), .C2(n21343), .A(n14089), .B(n14088), .ZN(
        n14091) );
  OR2_X1 U16043 ( .A1(n14091), .A2(n21430), .ZN(n14095) );
  INV_X1 U16044 ( .A(n14092), .ZN(n21428) );
  INV_X2 U16045 ( .A(n21428), .ZN(n21401) );
  NOR2_X2 U16046 ( .A1(n21401), .A2(n21403), .ZN(n21410) );
  AOI21_X1 U16047 ( .B1(n21410), .B2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n14093), .ZN(n14094) );
  NAND2_X1 U16048 ( .A1(n14097), .A2(n14096), .ZN(P3_U2831) );
  NAND2_X1 U16049 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15070) );
  NOR2_X1 U16050 ( .A1(n14098), .A2(n15070), .ZN(n14965) );
  NAND2_X1 U16051 ( .A1(n14099), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14124) );
  INV_X1 U16052 ( .A(n14124), .ZN(n14127) );
  NAND2_X1 U16053 ( .A1(n11487), .A2(n14116), .ZN(n14105) );
  NAND2_X1 U16054 ( .A1(n14099), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14100) );
  AND2_X1 U16055 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19458) );
  NAND2_X1 U16056 ( .A1(n19458), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n14111) );
  AOI21_X1 U16057 ( .B1(n14101), .B2(n14111), .A(n19549), .ZN(n14103) );
  INV_X1 U16058 ( .A(n14111), .ZN(n14102) );
  NAND2_X1 U16059 ( .A1(n14102), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19570) );
  AND2_X1 U16060 ( .A1(n14103), .A2(n19570), .ZN(n19410) );
  AOI21_X1 U16061 ( .B1(n14118), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19410), .ZN(n14104) );
  INV_X1 U16062 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14107) );
  NOR2_X1 U16063 ( .A1(n14346), .A2(n14107), .ZN(n14108) );
  INV_X1 U16064 ( .A(n19458), .ZN(n19519) );
  NAND2_X1 U16065 ( .A1(n19519), .A2(n19518), .ZN(n14110) );
  NAND2_X1 U16066 ( .A1(n14111), .A2(n14110), .ZN(n19411) );
  NOR2_X1 U16067 ( .A1(n19411), .A2(n19549), .ZN(n14112) );
  AOI21_X1 U16068 ( .B1(n14118), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n14112), .ZN(n14125) );
  NAND2_X1 U16069 ( .A1(n14417), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n14126) );
  NAND2_X1 U16070 ( .A1(n14118), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14114) );
  NAND2_X1 U16071 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19424), .ZN(
        n19534) );
  NAND2_X1 U16072 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19523), .ZN(
        n19547) );
  AND2_X1 U16073 ( .A1(n19534), .A2(n19547), .ZN(n19481) );
  OR2_X1 U16074 ( .A1(n19549), .A2(n19481), .ZN(n19535) );
  NAND2_X1 U16075 ( .A1(n14114), .A2(n19535), .ZN(n14115) );
  NOR2_X1 U16076 ( .A1(n19549), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n14117) );
  AOI21_X1 U16077 ( .B1(n14118), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n14117), .ZN(n14119) );
  NAND2_X1 U16078 ( .A1(n14417), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n14121) );
  XNOR2_X1 U16079 ( .A(n14733), .B(n14121), .ZN(n14783) );
  NAND2_X1 U16080 ( .A1(n14782), .A2(n14783), .ZN(n14785) );
  INV_X1 U16081 ( .A(n14733), .ZN(n15782) );
  NAND2_X1 U16082 ( .A1(n15782), .A2(n14121), .ZN(n14122) );
  NOR2_X1 U16083 ( .A1(n14346), .A2(n11596), .ZN(n14947) );
  AND2_X1 U16084 ( .A1(n14789), .A2(n14947), .ZN(n14123) );
  NAND2_X1 U16085 ( .A1(n14788), .A2(n14123), .ZN(n14130) );
  INV_X1 U16086 ( .A(n14947), .ZN(n14944) );
  INV_X1 U16087 ( .A(n14126), .ZN(n14915) );
  OR2_X1 U16088 ( .A1(n14127), .A2(n14915), .ZN(n14128) );
  NAND2_X1 U16089 ( .A1(n11252), .A2(n14128), .ZN(n14940) );
  NAND2_X1 U16090 ( .A1(n14130), .A2(n14129), .ZN(n14132) );
  AOI21_X1 U16091 ( .B1(n14942), .B2(n14132), .A(n14131), .ZN(n14133) );
  AOI22_X1 U16092 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n14270), .B1(
        n14271), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14140) );
  AOI22_X1 U16093 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n14151), .B1(
        n14150), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14139) );
  INV_X1 U16094 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14337) );
  INV_X1 U16095 ( .A(n14272), .ZN(n14260) );
  INV_X1 U16096 ( .A(n14273), .ZN(n14259) );
  OAI22_X1 U16097 ( .A1(n14337), .A2(n14260), .B1(n14259), .B2(n14135), .ZN(
        n14136) );
  AOI21_X1 U16098 ( .B1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n14269), .A(
        n14136), .ZN(n14138) );
  AOI22_X1 U16099 ( .A1(n14278), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14152), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14137) );
  NAND4_X1 U16100 ( .A1(n14140), .A2(n14139), .A3(n14138), .A4(n14137), .ZN(
        n14146) );
  AOI22_X1 U16101 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n14254), .B1(
        n14253), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14144) );
  AOI22_X1 U16102 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n14210), .B1(
        n14288), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14143) );
  NAND2_X1 U16103 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n14142) );
  NAND2_X1 U16104 ( .A1(n14287), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n14141) );
  NAND4_X1 U16105 ( .A1(n14144), .A2(n14143), .A3(n14142), .A4(n14141), .ZN(
        n14145) );
  NOR2_X1 U16106 ( .A1(n14146), .A2(n14145), .ZN(n14148) );
  NAND2_X1 U16107 ( .A1(n14295), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n14147) );
  AND2_X1 U16108 ( .A1(n14148), .A2(n14147), .ZN(n15710) );
  INV_X1 U16109 ( .A(n15710), .ZN(n14173) );
  INV_X1 U16110 ( .A(n15482), .ZN(n14149) );
  AND2_X1 U16111 ( .A1(n14149), .A2(n15397), .ZN(n15458) );
  AND2_X1 U16112 ( .A1(n15461), .A2(n15458), .ZN(n15459) );
  AND2_X1 U16113 ( .A1(n15576), .A2(n15459), .ZN(n15629) );
  INV_X1 U16114 ( .A(n14150), .ZN(n14227) );
  INV_X1 U16115 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14301) );
  INV_X1 U16116 ( .A(n14151), .ZN(n14225) );
  INV_X1 U16117 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14307) );
  OAI22_X1 U16118 ( .A1(n14227), .A2(n14301), .B1(n14225), .B2(n14307), .ZN(
        n14156) );
  INV_X1 U16119 ( .A(n14152), .ZN(n14228) );
  INV_X1 U16120 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14153) );
  OAI22_X1 U16121 ( .A1(n14230), .A2(n14154), .B1(n14228), .B2(n14153), .ZN(
        n14155) );
  NOR2_X1 U16122 ( .A1(n14156), .A2(n14155), .ZN(n14172) );
  INV_X1 U16123 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14158) );
  INV_X1 U16124 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14157) );
  OAI22_X1 U16125 ( .A1(n14285), .A2(n14158), .B1(n14284), .B2(n14157), .ZN(
        n14164) );
  NAND2_X1 U16126 ( .A1(n14287), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n14162) );
  NAND2_X1 U16127 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n14161) );
  NAND2_X1 U16128 ( .A1(n14288), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n14160) );
  NAND2_X1 U16129 ( .A1(n14210), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n14159) );
  NAND4_X1 U16130 ( .A1(n14162), .A2(n14161), .A3(n14160), .A4(n14159), .ZN(
        n14163) );
  NOR2_X1 U16131 ( .A1(n14164), .A2(n14163), .ZN(n14171) );
  NAND2_X1 U16132 ( .A1(n14269), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n14168) );
  NAND2_X1 U16133 ( .A1(n14270), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n14167) );
  NAND2_X1 U16134 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n14166) );
  AOI22_X1 U16135 ( .A1(n14273), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14165) );
  AND4_X1 U16136 ( .A1(n14168), .A2(n14167), .A3(n14166), .A4(n14165), .ZN(
        n14170) );
  NAND2_X1 U16137 ( .A1(n14295), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n14169) );
  NAND4_X1 U16138 ( .A1(n14172), .A2(n14171), .A3(n14170), .A4(n14169), .ZN(
        n15631) );
  AND2_X1 U16139 ( .A1(n15629), .A2(n15631), .ZN(n15630) );
  AND2_X1 U16140 ( .A1(n14173), .A2(n15630), .ZN(n15637) );
  INV_X1 U16141 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14174) );
  OAI22_X1 U16142 ( .A1(n14227), .A2(n14174), .B1(n14225), .B2(n14358), .ZN(
        n14178) );
  INV_X1 U16143 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14176) );
  INV_X1 U16144 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14175) );
  OAI22_X1 U16145 ( .A1(n14230), .A2(n14176), .B1(n14228), .B2(n14175), .ZN(
        n14177) );
  NOR2_X1 U16146 ( .A1(n14178), .A2(n14177), .ZN(n14194) );
  INV_X1 U16147 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14180) );
  INV_X1 U16148 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14179) );
  OAI22_X1 U16149 ( .A1(n14285), .A2(n14180), .B1(n14284), .B2(n14179), .ZN(
        n14186) );
  NAND2_X1 U16150 ( .A1(n14287), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n14184) );
  NAND2_X1 U16151 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n14183) );
  NAND2_X1 U16152 ( .A1(n14288), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n14182) );
  NAND2_X1 U16153 ( .A1(n14210), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n14181) );
  NAND4_X1 U16154 ( .A1(n14184), .A2(n14183), .A3(n14182), .A4(n14181), .ZN(
        n14185) );
  NOR2_X1 U16155 ( .A1(n14186), .A2(n14185), .ZN(n14193) );
  NAND2_X1 U16156 ( .A1(n14269), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n14190) );
  NAND2_X1 U16157 ( .A1(n14270), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n14189) );
  NAND2_X1 U16158 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n14188) );
  AOI22_X1 U16159 ( .A1(n14273), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14187) );
  AND4_X1 U16160 ( .A1(n14190), .A2(n14189), .A3(n14188), .A4(n14187), .ZN(
        n14192) );
  NAND2_X1 U16161 ( .A1(n14295), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n14191) );
  NAND4_X1 U16162 ( .A1(n14194), .A2(n14193), .A3(n14192), .A4(n14191), .ZN(
        n15639) );
  AND2_X1 U16163 ( .A1(n15637), .A2(n15639), .ZN(n14195) );
  AOI22_X1 U16164 ( .A1(n14270), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14271), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14201) );
  AOI22_X1 U16165 ( .A1(n14150), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14151), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14200) );
  INV_X1 U16166 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14384) );
  OAI22_X1 U16167 ( .A1(n14260), .A2(n14384), .B1(n14259), .B2(n14196), .ZN(
        n14197) );
  AOI21_X1 U16168 ( .B1(n14269), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A(
        n14197), .ZN(n14199) );
  AOI22_X1 U16169 ( .A1(n14278), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14152), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14198) );
  NAND4_X1 U16170 ( .A1(n14201), .A2(n14200), .A3(n14199), .A4(n14198), .ZN(
        n14207) );
  AOI22_X1 U16171 ( .A1(n14254), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n14253), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14205) );
  AOI22_X1 U16172 ( .A1(n14210), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14288), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14204) );
  NAND2_X1 U16173 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n14203) );
  NAND2_X1 U16174 ( .A1(n14287), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n14202) );
  NAND4_X1 U16175 ( .A1(n14205), .A2(n14204), .A3(n14203), .A4(n14202), .ZN(
        n14206) );
  NOR2_X1 U16176 ( .A1(n14207), .A2(n14206), .ZN(n14209) );
  NAND2_X1 U16177 ( .A1(n14295), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n14208) );
  AND2_X1 U16178 ( .A1(n14209), .A2(n14208), .ZN(n15882) );
  INV_X1 U16179 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14215) );
  INV_X1 U16180 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14399) );
  INV_X1 U16181 ( .A(n14210), .ZN(n14251) );
  INV_X1 U16182 ( .A(n14288), .ZN(n14250) );
  INV_X1 U16183 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14211) );
  OAI22_X1 U16184 ( .A1(n14399), .A2(n14251), .B1(n14250), .B2(n14211), .ZN(
        n14212) );
  AOI21_X1 U16185 ( .B1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B2(n11559), .A(
        n14212), .ZN(n14214) );
  AOI22_X1 U16186 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n14254), .B1(
        n14253), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14213) );
  OAI211_X1 U16187 ( .C1(n14215), .C2(n15306), .A(n14214), .B(n14213), .ZN(
        n14224) );
  INV_X1 U16188 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14409) );
  NOR2_X1 U16189 ( .A1(n14228), .A2(n14409), .ZN(n14218) );
  INV_X1 U16190 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14216) );
  INV_X1 U16191 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14407) );
  OAI22_X1 U16192 ( .A1(n14216), .A2(n14227), .B1(n14225), .B2(n14407), .ZN(
        n14217) );
  AOI211_X1 U16193 ( .C1(n14278), .C2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A(
        n14218), .B(n14217), .ZN(n14222) );
  AOI22_X1 U16194 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n14273), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14221) );
  AOI22_X1 U16195 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n14270), .B1(
        n14271), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14220) );
  NAND2_X1 U16196 ( .A1(n14269), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14219) );
  NAND4_X1 U16197 ( .A1(n14222), .A2(n14221), .A3(n14220), .A4(n14219), .ZN(
        n14223) );
  AOI211_X1 U16198 ( .C1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .C2(n14295), .A(
        n14224), .B(n14223), .ZN(n15947) );
  INV_X1 U16199 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14226) );
  INV_X1 U16200 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14429) );
  OAI22_X1 U16201 ( .A1(n14227), .A2(n14226), .B1(n14225), .B2(n14429), .ZN(
        n14232) );
  INV_X1 U16202 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14229) );
  INV_X1 U16203 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14432) );
  OAI22_X1 U16204 ( .A1(n14230), .A2(n14229), .B1(n14228), .B2(n14432), .ZN(
        n14231) );
  NOR2_X1 U16205 ( .A1(n14232), .A2(n14231), .ZN(n14248) );
  INV_X1 U16206 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14234) );
  INV_X1 U16207 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14233) );
  OAI22_X1 U16208 ( .A1(n14285), .A2(n14234), .B1(n14284), .B2(n14233), .ZN(
        n14240) );
  NAND2_X1 U16209 ( .A1(n14287), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n14238) );
  NAND2_X1 U16210 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n14237) );
  NAND2_X1 U16211 ( .A1(n14288), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n14236) );
  NAND2_X1 U16212 ( .A1(n14210), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n14235) );
  NAND4_X1 U16213 ( .A1(n14238), .A2(n14237), .A3(n14236), .A4(n14235), .ZN(
        n14239) );
  NOR2_X1 U16214 ( .A1(n14240), .A2(n14239), .ZN(n14247) );
  NAND2_X1 U16215 ( .A1(n14269), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n14244) );
  NAND2_X1 U16216 ( .A1(n14270), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n14243) );
  NAND2_X1 U16217 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n14242) );
  AOI22_X1 U16218 ( .A1(n14273), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14241) );
  AND4_X1 U16219 ( .A1(n14244), .A2(n14243), .A3(n14242), .A4(n14241), .ZN(
        n14246) );
  NAND2_X1 U16220 ( .A1(n14295), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n14245) );
  NAND4_X1 U16221 ( .A1(n14248), .A2(n14247), .A3(n14246), .A4(n14245), .ZN(
        n16690) );
  INV_X1 U16222 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14441) );
  OAI22_X1 U16223 ( .A1(n14441), .A2(n14251), .B1(n14250), .B2(n14249), .ZN(
        n14252) );
  AOI21_X1 U16224 ( .B1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B2(n11559), .A(
        n14252), .ZN(n14256) );
  AOI22_X1 U16225 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n14254), .B1(
        n14253), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14255) );
  OAI211_X1 U16226 ( .C1(n14257), .C2(n15306), .A(n14256), .B(n14255), .ZN(
        n14268) );
  AOI22_X1 U16227 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n14270), .B1(
        n14271), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14266) );
  AOI22_X1 U16228 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n14150), .B1(
        n14151), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14265) );
  OAI22_X1 U16229 ( .A1(n14261), .A2(n14260), .B1(n14259), .B2(n14258), .ZN(
        n14262) );
  AOI21_X1 U16230 ( .B1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n14269), .A(
        n14262), .ZN(n14264) );
  AOI22_X1 U16231 ( .A1(n14278), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14152), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14263) );
  NAND4_X1 U16232 ( .A1(n14266), .A2(n14265), .A3(n14264), .A4(n14263), .ZN(
        n14267) );
  AOI211_X1 U16233 ( .C1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .C2(n14295), .A(
        n14268), .B(n14267), .ZN(n16685) );
  NOR2_X2 U16234 ( .A1(n16683), .A2(n16685), .ZN(n16679) );
  NAND2_X1 U16235 ( .A1(n14269), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n14277) );
  NAND2_X1 U16236 ( .A1(n14270), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n14276) );
  NAND2_X1 U16237 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n14275) );
  AOI22_X1 U16238 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n14273), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14274) );
  AND4_X1 U16239 ( .A1(n14277), .A2(n14276), .A3(n14275), .A4(n14274), .ZN(
        n14299) );
  NAND2_X1 U16240 ( .A1(n14278), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n14282) );
  NAND2_X1 U16241 ( .A1(n14150), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n14281) );
  NAND2_X1 U16242 ( .A1(n14151), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n14280) );
  NAND2_X1 U16243 ( .A1(n14152), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n14279) );
  AND4_X1 U16244 ( .A1(n14282), .A2(n14281), .A3(n14280), .A4(n14279), .ZN(
        n14298) );
  INV_X1 U16245 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14286) );
  INV_X1 U16246 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14283) );
  OAI22_X1 U16247 ( .A1(n14286), .A2(n14285), .B1(n14284), .B2(n14283), .ZN(
        n14294) );
  NAND2_X1 U16248 ( .A1(n14287), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n14292) );
  NAND2_X1 U16249 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n14291) );
  NAND2_X1 U16250 ( .A1(n14288), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n14290) );
  NAND2_X1 U16251 ( .A1(n14210), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n14289) );
  NAND4_X1 U16252 ( .A1(n14292), .A2(n14291), .A3(n14290), .A4(n14289), .ZN(
        n14293) );
  NOR2_X1 U16253 ( .A1(n14294), .A2(n14293), .ZN(n14297) );
  NAND2_X1 U16254 ( .A1(n14295), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n14296) );
  NAND4_X1 U16255 ( .A1(n14299), .A2(n14298), .A3(n14297), .A4(n14296), .ZN(
        n14325) );
  INV_X1 U16256 ( .A(n14484), .ZN(n14444) );
  INV_X1 U16257 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14302) );
  INV_X1 U16258 ( .A(n14453), .ZN(n14475) );
  OAI22_X1 U16259 ( .A1(n14444), .A2(n14302), .B1(n14475), .B2(n14301), .ZN(
        n14309) );
  INV_X1 U16260 ( .A(n14467), .ZN(n14473) );
  NAND2_X1 U16261 ( .A1(n14480), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n14306) );
  INV_X1 U16262 ( .A(n14303), .ZN(n14305) );
  NAND2_X1 U16263 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14304) );
  AND2_X1 U16264 ( .A1(n14305), .A2(n14304), .ZN(n14431) );
  OAI211_X1 U16265 ( .C1(n14473), .C2(n14307), .A(n14306), .B(n14431), .ZN(
        n14308) );
  NOR2_X1 U16266 ( .A1(n14309), .A2(n14308), .ZN(n14312) );
  AOI22_X1 U16267 ( .A1(n14483), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10962), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14311) );
  AOI22_X1 U16268 ( .A1(n14482), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14481), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14310) );
  NAND3_X1 U16269 ( .A1(n14312), .A2(n14311), .A3(n14310), .ZN(n14322) );
  AOI22_X1 U16270 ( .A1(n14483), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10962), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14320) );
  AOI22_X1 U16271 ( .A1(n14482), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14481), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14319) );
  AOI22_X1 U16272 ( .A1(n14484), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14453), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14318) );
  INV_X1 U16273 ( .A(n14480), .ZN(n15297) );
  INV_X1 U16274 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14315) );
  INV_X1 U16275 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14313) );
  OR2_X1 U16276 ( .A1(n14473), .A2(n14313), .ZN(n14314) );
  INV_X1 U16277 ( .A(n14431), .ZN(n14471) );
  OAI211_X1 U16278 ( .C1(n15297), .C2(n14315), .A(n14314), .B(n14471), .ZN(
        n14316) );
  INV_X1 U16279 ( .A(n14316), .ZN(n14317) );
  NAND4_X1 U16280 ( .A1(n14320), .A2(n14319), .A3(n14318), .A4(n14317), .ZN(
        n14321) );
  NAND2_X1 U16281 ( .A1(n14322), .A2(n14321), .ZN(n14323) );
  XNOR2_X1 U16282 ( .A(n14325), .B(n14323), .ZN(n16680) );
  INV_X1 U16283 ( .A(n14323), .ZN(n14324) );
  INV_X1 U16284 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14327) );
  OAI22_X1 U16285 ( .A1(n14444), .A2(n14327), .B1(n14475), .B2(n14326), .ZN(
        n14331) );
  NAND2_X1 U16286 ( .A1(n14480), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n14328) );
  OAI211_X1 U16287 ( .C1(n14473), .C2(n14329), .A(n14328), .B(n14431), .ZN(
        n14330) );
  NOR2_X1 U16288 ( .A1(n14331), .A2(n14330), .ZN(n14334) );
  AOI22_X1 U16289 ( .A1(n14483), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10962), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14333) );
  AOI22_X1 U16290 ( .A1(n14482), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14481), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14332) );
  NAND3_X1 U16291 ( .A1(n14334), .A2(n14333), .A3(n14332), .ZN(n14344) );
  AOI22_X1 U16292 ( .A1(n14483), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10962), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14342) );
  AOI22_X1 U16293 ( .A1(n14482), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14481), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14341) );
  AOI22_X1 U16294 ( .A1(n14484), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n14453), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14340) );
  OR2_X1 U16295 ( .A1(n14473), .A2(n14335), .ZN(n14336) );
  OAI211_X1 U16296 ( .C1(n15297), .C2(n14337), .A(n14336), .B(n14471), .ZN(
        n14338) );
  INV_X1 U16297 ( .A(n14338), .ZN(n14339) );
  NAND4_X1 U16298 ( .A1(n14342), .A2(n14341), .A3(n14340), .A4(n14339), .ZN(
        n14343) );
  NAND2_X1 U16299 ( .A1(n14344), .A2(n14343), .ZN(n14367) );
  INV_X1 U16300 ( .A(n14367), .ZN(n14345) );
  NAND2_X1 U16301 ( .A1(n11969), .A2(n14345), .ZN(n14348) );
  INV_X1 U16302 ( .A(n14369), .ZN(n14366) );
  OAI21_X1 U16303 ( .B1(n14346), .B2(n14366), .A(n14367), .ZN(n14347) );
  OAI21_X1 U16304 ( .B1(n14348), .B2(n14366), .A(n14347), .ZN(n16675) );
  AOI22_X1 U16305 ( .A1(n14483), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10962), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14356) );
  AOI22_X1 U16306 ( .A1(n14482), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14481), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14355) );
  AOI22_X1 U16307 ( .A1(n14484), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n14453), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14354) );
  INV_X1 U16308 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14351) );
  INV_X1 U16309 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14349) );
  OR2_X1 U16310 ( .A1(n14473), .A2(n14349), .ZN(n14350) );
  OAI211_X1 U16311 ( .C1(n15297), .C2(n14351), .A(n14350), .B(n14471), .ZN(
        n14352) );
  INV_X1 U16312 ( .A(n14352), .ZN(n14353) );
  NAND4_X1 U16313 ( .A1(n14356), .A2(n14355), .A3(n14354), .A4(n14353), .ZN(
        n14365) );
  AOI22_X1 U16314 ( .A1(n14483), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10962), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14363) );
  AOI22_X1 U16315 ( .A1(n14482), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14481), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14362) );
  AOI22_X1 U16316 ( .A1(n14484), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14453), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14361) );
  NAND2_X1 U16317 ( .A1(n14480), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n14357) );
  OAI211_X1 U16318 ( .C1(n14473), .C2(n14358), .A(n14357), .B(n14431), .ZN(
        n14359) );
  INV_X1 U16319 ( .A(n14359), .ZN(n14360) );
  NAND4_X1 U16320 ( .A1(n14363), .A2(n14362), .A3(n14361), .A4(n14360), .ZN(
        n14364) );
  NAND2_X1 U16321 ( .A1(n14365), .A2(n14364), .ZN(n14371) );
  OAI21_X1 U16322 ( .B1(n14366), .B2(n14367), .A(n14371), .ZN(n14370) );
  NOR2_X1 U16323 ( .A1(n14367), .A2(n14371), .ZN(n14368) );
  NAND2_X1 U16324 ( .A1(n14369), .A2(n14368), .ZN(n14392) );
  NAND3_X1 U16325 ( .A1(n14417), .A2(n14370), .A3(n14392), .ZN(n14372) );
  NOR2_X1 U16326 ( .A1(n11969), .A2(n14371), .ZN(n16664) );
  INV_X1 U16327 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14374) );
  OAI22_X1 U16328 ( .A1(n14444), .A2(n14374), .B1(n14475), .B2(n14373), .ZN(
        n14378) );
  NAND2_X1 U16329 ( .A1(n14480), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n14375) );
  OAI211_X1 U16330 ( .C1(n14473), .C2(n14376), .A(n14375), .B(n14431), .ZN(
        n14377) );
  NOR2_X1 U16331 ( .A1(n14378), .A2(n14377), .ZN(n14381) );
  AOI22_X1 U16332 ( .A1(n14483), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10962), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14380) );
  AOI22_X1 U16333 ( .A1(n14482), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14481), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14379) );
  NAND3_X1 U16334 ( .A1(n14381), .A2(n14380), .A3(n14379), .ZN(n14391) );
  AOI22_X1 U16335 ( .A1(n14483), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10962), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14389) );
  AOI22_X1 U16336 ( .A1(n14482), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14481), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14388) );
  AOI22_X1 U16337 ( .A1(n14484), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n14453), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14387) );
  OR2_X1 U16338 ( .A1(n14473), .A2(n14382), .ZN(n14383) );
  OAI211_X1 U16339 ( .C1(n15297), .C2(n14384), .A(n14383), .B(n14471), .ZN(
        n14385) );
  INV_X1 U16340 ( .A(n14385), .ZN(n14386) );
  NAND4_X1 U16341 ( .A1(n14389), .A2(n14388), .A3(n14387), .A4(n14386), .ZN(
        n14390) );
  NAND2_X1 U16342 ( .A1(n14391), .A2(n14390), .ZN(n14394) );
  OR2_X1 U16343 ( .A1(n14392), .A2(n14394), .ZN(n14398) );
  NAND2_X1 U16344 ( .A1(n14392), .A2(n14394), .ZN(n14393) );
  INV_X1 U16346 ( .A(n14394), .ZN(n14395) );
  NAND2_X1 U16347 ( .A1(n10959), .A2(n14395), .ZN(n16659) );
  INV_X1 U16348 ( .A(n14398), .ZN(n14418) );
  AOI22_X1 U16349 ( .A1(n14482), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10962), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14406) );
  AOI22_X1 U16350 ( .A1(n14483), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14481), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14405) );
  AOI22_X1 U16351 ( .A1(n14484), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n14453), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14404) );
  INV_X1 U16352 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14401) );
  OR2_X1 U16353 ( .A1(n14473), .A2(n14399), .ZN(n14400) );
  OAI211_X1 U16354 ( .C1(n15297), .C2(n14401), .A(n14400), .B(n14471), .ZN(
        n14402) );
  INV_X1 U16355 ( .A(n14402), .ZN(n14403) );
  NAND4_X1 U16356 ( .A1(n14406), .A2(n14405), .A3(n14404), .A4(n14403), .ZN(
        n14416) );
  AOI22_X1 U16357 ( .A1(n14482), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14483), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14414) );
  AOI22_X1 U16358 ( .A1(n10961), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14481), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14413) );
  AOI22_X1 U16359 ( .A1(n14484), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14453), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14412) );
  OR2_X1 U16360 ( .A1(n14473), .A2(n14407), .ZN(n14408) );
  OAI211_X1 U16361 ( .C1(n15297), .C2(n14409), .A(n14431), .B(n14408), .ZN(
        n14410) );
  INV_X1 U16362 ( .A(n14410), .ZN(n14411) );
  NAND4_X1 U16363 ( .A1(n14414), .A2(n14413), .A3(n14412), .A4(n14411), .ZN(
        n14415) );
  AND2_X1 U16364 ( .A1(n14416), .A2(n14415), .ZN(n14419) );
  NAND2_X1 U16365 ( .A1(n14418), .A2(n14419), .ZN(n16640) );
  OAI211_X1 U16366 ( .C1(n14418), .C2(n14419), .A(n16640), .B(n14417), .ZN(
        n14440) );
  INV_X1 U16367 ( .A(n14419), .ZN(n14420) );
  NOR2_X1 U16368 ( .A1(n11969), .A2(n14420), .ZN(n16650) );
  AOI22_X1 U16369 ( .A1(n14483), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10961), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14428) );
  AOI22_X1 U16370 ( .A1(n14482), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14481), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14427) );
  AOI22_X1 U16371 ( .A1(n14484), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14453), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14426) );
  INV_X1 U16372 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14423) );
  OR2_X1 U16373 ( .A1(n14473), .A2(n14421), .ZN(n14422) );
  OAI211_X1 U16374 ( .C1(n15297), .C2(n14423), .A(n14422), .B(n14471), .ZN(
        n14424) );
  INV_X1 U16375 ( .A(n14424), .ZN(n14425) );
  NAND4_X1 U16376 ( .A1(n14428), .A2(n14427), .A3(n14426), .A4(n14425), .ZN(
        n14439) );
  AOI22_X1 U16377 ( .A1(n14483), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10961), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14437) );
  AOI22_X1 U16378 ( .A1(n14482), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14481), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14436) );
  AOI22_X1 U16379 ( .A1(n14484), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14453), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14435) );
  OR2_X1 U16380 ( .A1(n14473), .A2(n14429), .ZN(n14430) );
  OAI211_X1 U16381 ( .C1(n15297), .C2(n14432), .A(n14431), .B(n14430), .ZN(
        n14433) );
  INV_X1 U16382 ( .A(n14433), .ZN(n14434) );
  NAND4_X1 U16383 ( .A1(n14437), .A2(n14436), .A3(n14435), .A4(n14434), .ZN(
        n14438) );
  AND2_X1 U16384 ( .A1(n14439), .A2(n14438), .ZN(n14463) );
  OAI21_X1 U16385 ( .B1(n14473), .B2(n14441), .A(n14471), .ZN(n14446) );
  INV_X1 U16386 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14443) );
  OAI22_X1 U16387 ( .A1(n14444), .A2(n14443), .B1(n14475), .B2(n14442), .ZN(
        n14445) );
  AOI211_X1 U16388 ( .C1(n14480), .C2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n14446), .B(n14445), .ZN(n14449) );
  AOI22_X1 U16389 ( .A1(n14483), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14481), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14448) );
  AOI22_X1 U16390 ( .A1(n14482), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10962), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14447) );
  NAND3_X1 U16391 ( .A1(n14449), .A2(n14448), .A3(n14447), .ZN(n14459) );
  NOR2_X1 U16392 ( .A1(n14473), .A2(n14450), .ZN(n14451) );
  AOI211_X1 U16393 ( .C1(n14480), .C2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n14471), .B(n14451), .ZN(n14457) );
  AOI22_X1 U16394 ( .A1(n14482), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10961), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14456) );
  AOI22_X1 U16395 ( .A1(n14484), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14483), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14455) );
  AOI22_X1 U16396 ( .A1(n14481), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14453), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14454) );
  NAND4_X1 U16397 ( .A1(n14457), .A2(n14456), .A3(n14455), .A4(n14454), .ZN(
        n14458) );
  NAND2_X1 U16398 ( .A1(n14459), .A2(n14458), .ZN(n14460) );
  INV_X1 U16400 ( .A(n14463), .ZN(n16642) );
  NOR3_X1 U16401 ( .A1(n16640), .A2(n10959), .A3(n16642), .ZN(n16632) );
  AOI22_X1 U16402 ( .A1(n14482), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14483), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14466) );
  AOI22_X1 U16403 ( .A1(n11341), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14481), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14465) );
  NAND2_X1 U16404 ( .A1(n14466), .A2(n14465), .ZN(n14490) );
  INV_X1 U16405 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14470) );
  AOI22_X1 U16406 ( .A1(n14484), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14480), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14469) );
  AOI21_X1 U16407 ( .B1(n14467), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n14471), .ZN(n14468) );
  OAI211_X1 U16408 ( .C1(n14475), .C2(n14470), .A(n14469), .B(n14468), .ZN(
        n14489) );
  INV_X1 U16409 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14472) );
  OAI21_X1 U16410 ( .B1(n14473), .B2(n14472), .A(n14471), .ZN(n14479) );
  INV_X1 U16411 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14476) );
  INV_X1 U16412 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14474) );
  OAI22_X1 U16413 ( .A1(n10963), .A2(n14476), .B1(n14475), .B2(n14474), .ZN(
        n14478) );
  AOI211_X1 U16414 ( .C1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .C2(n14480), .A(
        n14479), .B(n14478), .ZN(n14487) );
  AOI22_X1 U16415 ( .A1(n14482), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14481), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14486) );
  AOI22_X1 U16416 ( .A1(n14484), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n14483), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14485) );
  NAND3_X1 U16417 ( .A1(n14487), .A2(n14486), .A3(n14485), .ZN(n14488) );
  OAI21_X1 U16418 ( .B1(n14490), .B2(n14489), .A(n14488), .ZN(n14491) );
  INV_X1 U16419 ( .A(n14491), .ZN(n14492) );
  INV_X1 U16420 ( .A(n15781), .ZN(n14493) );
  NAND2_X1 U16421 ( .A1(n14493), .A2(n15321), .ZN(n15260) );
  NAND2_X1 U16422 ( .A1(n15260), .A2(n15268), .ZN(n14494) );
  NAND2_X1 U16423 ( .A1(n15993), .A2(n16651), .ZN(n14496) );
  NAND2_X1 U16424 ( .A1(n16689), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14495) );
  OAI21_X1 U16425 ( .B1(n16077), .B2(n16698), .A(n11232), .ZN(P2_U2857) );
  NAND2_X1 U16426 ( .A1(n16798), .A2(n14497), .ZN(n15977) );
  INV_X1 U16427 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16061) );
  XNOR2_X1 U16428 ( .A(n15979), .B(n16061), .ZN(n14521) );
  NAND2_X1 U16429 ( .A1(n14521), .A2(n12326), .ZN(n14520) );
  INV_X1 U16430 ( .A(n14499), .ZN(n15984) );
  OAI21_X1 U16431 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14498), .A(
        n15984), .ZN(n14522) );
  OR2_X1 U16432 ( .A1(n14522), .A2(n17277), .ZN(n14519) );
  NAND2_X1 U16433 ( .A1(n14500), .A2(n14501), .ZN(n14502) );
  NAND2_X1 U16434 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14509) );
  INV_X1 U16435 ( .A(n17262), .ZN(n18890) );
  AND2_X1 U16436 ( .A1(n18890), .A2(n14503), .ZN(n14507) );
  INV_X1 U16437 ( .A(n14507), .ZN(n14508) );
  INV_X1 U16438 ( .A(n14504), .ZN(n14505) );
  NAND2_X1 U16439 ( .A1(n14506), .A2(n14505), .ZN(n14514) );
  INV_X1 U16440 ( .A(n17227), .ZN(n17261) );
  AOI211_X1 U16441 ( .C1(n17262), .C2(n14514), .A(n17036), .B(n17261), .ZN(
        n17034) );
  NOR2_X1 U16442 ( .A1(n17034), .A2(n14507), .ZN(n17026) );
  AOI21_X1 U16443 ( .B1(n14509), .B2(n14508), .A(n17026), .ZN(n16065) );
  NOR2_X1 U16444 ( .A1(n16065), .A2(n16061), .ZN(n14517) );
  OR2_X1 U16445 ( .A1(n14511), .A2(n14512), .ZN(n14513) );
  NAND2_X1 U16446 ( .A1(n14510), .A2(n14513), .ZN(n16722) );
  OR2_X1 U16447 ( .A1(n15698), .A2(n14514), .ZN(n17035) );
  NOR2_X1 U16448 ( .A1(n17035), .A2(n14515), .ZN(n17017) );
  NAND2_X1 U16449 ( .A1(n17017), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17001) );
  INV_X1 U16450 ( .A(n17001), .ZN(n15996) );
  NAND2_X1 U16451 ( .A1(n15996), .A2(n16061), .ZN(n16064) );
  NAND2_X1 U16452 ( .A1(n12161), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n14523) );
  OAI211_X1 U16453 ( .C1(n17229), .C2(n16722), .A(n16064), .B(n14523), .ZN(
        n14516) );
  AOI211_X1 U16454 ( .C1(n16652), .C2(n17204), .A(n14517), .B(n14516), .ZN(
        n14518) );
  NAND2_X1 U16455 ( .A1(n14520), .A2(n11253), .ZN(P2_U3019) );
  INV_X1 U16456 ( .A(n17670), .ZN(n17617) );
  NAND2_X1 U16457 ( .A1(n14521), .A2(n17617), .ZN(n14529) );
  NAND2_X1 U16458 ( .A1(n17647), .A2(n16603), .ZN(n14524) );
  OAI211_X1 U16459 ( .C1(n17658), .C2(n14525), .A(n14524), .B(n14523), .ZN(
        n14526) );
  AOI21_X1 U16460 ( .B1(n16652), .B2(n17672), .A(n14526), .ZN(n14527) );
  NAND2_X1 U16461 ( .A1(n14529), .A2(n11233), .ZN(P2_U2987) );
  XNOR2_X1 U16462 ( .A(n14532), .B(n14531), .ZN(n16316) );
  NAND2_X1 U16463 ( .A1(n16316), .A2(n13627), .ZN(n14541) );
  INV_X1 U16464 ( .A(n16088), .ZN(n14534) );
  OAI22_X1 U16465 ( .A1(n14536), .A2(n14535), .B1(n14534), .B2(n14533), .ZN(
        n14538) );
  XNOR2_X1 U16466 ( .A(n14538), .B(n14537), .ZN(n16412) );
  INV_X1 U16467 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n16051) );
  NOR2_X1 U16468 ( .A1(n20137), .A2(n16051), .ZN(n14539) );
  NAND2_X1 U16469 ( .A1(n14541), .A2(n14540), .ZN(P1_U2842) );
  NOR2_X1 U16470 ( .A1(P2_BE_N_REG_3__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .ZN(n14543) );
  NOR4_X1 U16471 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_0__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n14542) );
  NAND4_X1 U16472 ( .A1(n14543), .A2(P2_M_IO_N_REG_SCAN_IN), .A3(
        P2_W_R_N_REG_SCAN_IN), .A4(n14542), .ZN(n14565) );
  NOR2_X1 U16473 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n14565), .ZN(n19095)
         );
  NOR4_X1 U16474 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n14547) );
  NOR4_X1 U16475 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n14546) );
  NOR4_X1 U16476 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n14545) );
  NOR4_X1 U16477 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n14544) );
  AND4_X1 U16478 ( .A1(n14547), .A2(n14546), .A3(n14545), .A4(n14544), .ZN(
        n14552) );
  NOR4_X1 U16479 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n14550) );
  NOR4_X1 U16480 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n14549) );
  NOR4_X1 U16481 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n14548) );
  INV_X1 U16482 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20046) );
  AND4_X1 U16483 ( .A1(n14550), .A2(n14549), .A3(n14548), .A4(n20046), .ZN(
        n14551) );
  NAND2_X1 U16484 ( .A1(n14552), .A2(n14551), .ZN(n14553) );
  INV_X1 U16485 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20273) );
  INV_X1 U16486 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n22399) );
  NOR4_X1 U16487 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n20273), .A4(n22399), .ZN(n14555) );
  NOR4_X1 U16488 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_D_C_N_REG_SCAN_IN), .A3(
        P1_BE_N_REG_1__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n14554) );
  NAND3_X1 U16489 ( .A1(n15942), .A2(n14555), .A3(n14554), .ZN(U214) );
  NOR4_X1 U16490 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n14559) );
  NOR4_X1 U16491 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n14558) );
  NOR4_X1 U16492 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n14557) );
  NOR4_X1 U16493 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n14556) );
  NAND4_X1 U16494 ( .A1(n14559), .A2(n14558), .A3(n14557), .A4(n14556), .ZN(
        n14564) );
  NOR4_X1 U16495 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n14562) );
  NOR4_X1 U16496 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n14561) );
  NOR4_X1 U16497 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n14560) );
  INV_X1 U16498 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19954) );
  NAND4_X1 U16499 ( .A1(n14562), .A2(n14561), .A3(n14560), .A4(n19954), .ZN(
        n14563) );
  OR2_X1 U16500 ( .A1(n19375), .A2(n14565), .ZN(n20207) );
  INV_X2 U16501 ( .A(U214), .ZN(n20258) );
  OR2_X1 U16502 ( .A1(n20207), .A2(n20258), .ZN(U212) );
  AOI211_X1 U16503 ( .C1(n16971), .C2(n14566), .A(n18673), .B(n18605), .ZN(
        n14577) );
  AOI21_X1 U16504 ( .B1(n14567), .B2(n14797), .A(n14937), .ZN(n17188) );
  INV_X1 U16505 ( .A(n17188), .ZN(n19366) );
  AOI22_X1 U16506 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n18851), .B1(
        P2_REIP_REG_11__SCAN_IN), .B2(n18850), .ZN(n14568) );
  OAI211_X1 U16507 ( .C1(n19366), .C2(n18855), .A(n14568), .B(n18746), .ZN(
        n14576) );
  OAI22_X1 U16508 ( .A1(n14569), .A2(n18803), .B1(n18733), .B2(n11862), .ZN(
        n14575) );
  OR2_X1 U16509 ( .A1(n15187), .A2(n14571), .ZN(n14572) );
  NAND2_X1 U16510 ( .A1(n14570), .A2(n14572), .ZN(n17190) );
  NAND2_X1 U16511 ( .A1(n18717), .A2(n18861), .ZN(n18776) );
  INV_X1 U16512 ( .A(n16971), .ZN(n14573) );
  OAI22_X1 U16513 ( .A1(n17190), .A2(n18857), .B1(n18776), .B2(n14573), .ZN(
        n14574) );
  OR4_X1 U16514 ( .A1(n14577), .A2(n14576), .A3(n14575), .A4(n14574), .ZN(
        P2_U2844) );
  NOR2_X1 U16515 ( .A1(n14578), .A2(n18870), .ZN(n18614) );
  INV_X1 U16516 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n17706) );
  OAI211_X1 U16517 ( .C1(n18614), .C2(n17706), .A(n17602), .B(n14581), .ZN(
        P2_U2814) );
  INV_X1 U16518 ( .A(n11921), .ZN(n18585) );
  INV_X1 U16519 ( .A(n17602), .ZN(n14579) );
  OAI21_X1 U16520 ( .B1(n14579), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n18589), 
        .ZN(n14580) );
  OAI21_X1 U16521 ( .B1(n18585), .B2(n18589), .A(n14580), .ZN(P2_U3612) );
  OAI21_X2 U16522 ( .B1(n14581), .B2(n21850), .A(n14690), .ZN(n14644) );
  INV_X1 U16523 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n14584) );
  INV_X1 U16524 ( .A(n14581), .ZN(n14582) );
  NAND3_X1 U16525 ( .A1(n14582), .A2(n11969), .A3(n18908), .ZN(n14642) );
  AOI22_X1 U16526 ( .A1(n19376), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n19375), .ZN(n19378) );
  NOR2_X1 U16527 ( .A1(n14642), .A2(n19378), .ZN(n14589) );
  AOI21_X1 U16528 ( .B1(n14616), .B2(P2_EAX_REG_23__SCAN_IN), .A(n14589), .ZN(
        n14583) );
  OAI21_X1 U16529 ( .B1(n14644), .B2(n14584), .A(n14583), .ZN(P2_U2959) );
  INV_X1 U16530 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n14586) );
  AOI22_X1 U16531 ( .A1(n19376), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n19375), .ZN(n19631) );
  NOR2_X1 U16532 ( .A1(n14642), .A2(n19631), .ZN(n14592) );
  AOI21_X1 U16533 ( .B1(n14616), .B2(P2_EAX_REG_21__SCAN_IN), .A(n14592), .ZN(
        n14585) );
  OAI21_X1 U16534 ( .B1(n14644), .B2(n14586), .A(n14585), .ZN(P2_U2957) );
  INV_X1 U16535 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n14588) );
  AOI22_X1 U16536 ( .A1(n19376), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n19375), .ZN(n19751) );
  NOR2_X1 U16537 ( .A1(n14642), .A2(n19751), .ZN(n14606) );
  AOI21_X1 U16538 ( .B1(n14616), .B2(P2_EAX_REG_18__SCAN_IN), .A(n14606), .ZN(
        n14587) );
  OAI21_X1 U16539 ( .B1(n14644), .B2(n14588), .A(n14587), .ZN(P2_U2954) );
  INV_X1 U16540 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n14591) );
  AOI21_X1 U16541 ( .B1(n14616), .B2(P2_EAX_REG_7__SCAN_IN), .A(n14589), .ZN(
        n14590) );
  OAI21_X1 U16542 ( .B1(n14644), .B2(n14591), .A(n14590), .ZN(P2_U2974) );
  INV_X1 U16543 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n14594) );
  AOI21_X1 U16544 ( .B1(n14616), .B2(P2_EAX_REG_5__SCAN_IN), .A(n14592), .ZN(
        n14593) );
  OAI21_X1 U16545 ( .B1(n14644), .B2(n14594), .A(n14593), .ZN(P2_U2972) );
  INV_X1 U16546 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n14596) );
  AOI22_X1 U16547 ( .A1(n19376), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19375), .ZN(n19838) );
  NOR2_X1 U16548 ( .A1(n14642), .A2(n19838), .ZN(n14603) );
  AOI21_X1 U16549 ( .B1(n14616), .B2(P2_EAX_REG_16__SCAN_IN), .A(n14603), .ZN(
        n14595) );
  OAI21_X1 U16550 ( .B1(n14644), .B2(n14596), .A(n14595), .ZN(P2_U2952) );
  INV_X1 U16551 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n14598) );
  AOI22_X1 U16552 ( .A1(n19376), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19375), .ZN(n19712) );
  NOR2_X1 U16553 ( .A1(n14642), .A2(n19712), .ZN(n14612) );
  AOI21_X1 U16554 ( .B1(n14616), .B2(P2_EAX_REG_19__SCAN_IN), .A(n14612), .ZN(
        n14597) );
  OAI21_X1 U16555 ( .B1(n14644), .B2(n14598), .A(n14597), .ZN(P2_U2955) );
  INV_X1 U16556 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n14600) );
  AOI22_X1 U16557 ( .A1(n19376), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19375), .ZN(n19792) );
  NOR2_X1 U16558 ( .A1(n14642), .A2(n19792), .ZN(n14615) );
  AOI21_X1 U16559 ( .B1(n14616), .B2(P2_EAX_REG_17__SCAN_IN), .A(n14615), .ZN(
        n14599) );
  OAI21_X1 U16560 ( .B1(n14644), .B2(n14600), .A(n14599), .ZN(P2_U2953) );
  INV_X1 U16561 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n14602) );
  AOI22_X1 U16562 ( .A1(n19376), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n19375), .ZN(n19672) );
  NOR2_X1 U16563 ( .A1(n14642), .A2(n19672), .ZN(n14609) );
  AOI21_X1 U16564 ( .B1(n14616), .B2(P2_EAX_REG_20__SCAN_IN), .A(n14609), .ZN(
        n14601) );
  OAI21_X1 U16565 ( .B1(n14644), .B2(n14602), .A(n14601), .ZN(P2_U2956) );
  INV_X1 U16566 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n14605) );
  AOI21_X1 U16567 ( .B1(P2_EAX_REG_0__SCAN_IN), .B2(n14616), .A(n14603), .ZN(
        n14604) );
  OAI21_X1 U16568 ( .B1(n14644), .B2(n14605), .A(n14604), .ZN(P2_U2967) );
  INV_X1 U16569 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n14608) );
  AOI21_X1 U16570 ( .B1(P2_EAX_REG_2__SCAN_IN), .B2(n14616), .A(n14606), .ZN(
        n14607) );
  OAI21_X1 U16571 ( .B1(n14644), .B2(n14608), .A(n14607), .ZN(P2_U2969) );
  INV_X1 U16572 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n14611) );
  AOI21_X1 U16573 ( .B1(P2_EAX_REG_4__SCAN_IN), .B2(n14616), .A(n14609), .ZN(
        n14610) );
  OAI21_X1 U16574 ( .B1(n14644), .B2(n14611), .A(n14610), .ZN(P2_U2971) );
  INV_X1 U16575 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n14614) );
  AOI21_X1 U16576 ( .B1(P2_EAX_REG_3__SCAN_IN), .B2(n14616), .A(n14612), .ZN(
        n14613) );
  OAI21_X1 U16577 ( .B1(n14644), .B2(n14614), .A(n14613), .ZN(P2_U2970) );
  INV_X1 U16578 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n14618) );
  AOI21_X1 U16579 ( .B1(P2_EAX_REG_1__SCAN_IN), .B2(n14616), .A(n14615), .ZN(
        n14617) );
  OAI21_X1 U16580 ( .B1(n14644), .B2(n14618), .A(n14617), .ZN(P2_U2968) );
  AOI22_X1 U16581 ( .A1(n19376), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19375), .ZN(n15426) );
  INV_X1 U16582 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n14619) );
  INV_X1 U16583 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n17739) );
  OAI222_X1 U16584 ( .A1(n14642), .A2(n15426), .B1(n14644), .B2(n14619), .C1(
        n14690), .C2(n17739), .ZN(P2_U2982) );
  NOR2_X1 U16585 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n22115), .ZN(n15837) );
  AOI21_X1 U16586 ( .B1(P1_MEMORYFETCH_REG_SCAN_IN), .B2(n14620), .A(n15837), 
        .ZN(n14621) );
  NAND2_X1 U16587 ( .A1(n14744), .A2(n14621), .ZN(P1_U2801) );
  INV_X1 U16588 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14631) );
  AOI21_X1 U16589 ( .B1(n14624), .B2(n14623), .A(n14622), .ZN(n14724) );
  INV_X1 U16590 ( .A(n14724), .ZN(n14625) );
  NAND2_X1 U16591 ( .A1(n16976), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n14723) );
  OAI21_X1 U16592 ( .B1(n17648), .B2(n14625), .A(n14723), .ZN(n14630) );
  NAND2_X1 U16593 ( .A1(n16013), .A2(n14626), .ZN(n14628) );
  INV_X1 U16594 ( .A(n16012), .ZN(n14627) );
  AOI22_X1 U16595 ( .A1(n14628), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n16013), .B2(n14627), .ZN(n14727) );
  OAI22_X1 U16596 ( .A1(n14727), .A2(n17670), .B1(n17658), .B2(n14631), .ZN(
        n14629) );
  AOI211_X1 U16597 ( .C1(n17647), .C2(n14631), .A(n14630), .B(n14629), .ZN(
        n14632) );
  OAI21_X1 U16598 ( .B1(n11489), .B2(n17651), .A(n14632), .ZN(P2_U3013) );
  INV_X1 U16599 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n16748) );
  INV_X1 U16600 ( .A(n18870), .ZN(n15261) );
  NAND2_X1 U16601 ( .A1(n15261), .A2(n18592), .ZN(n14633) );
  OAI21_X1 U16602 ( .B1(n14634), .B2(n14633), .A(n14690), .ZN(n14635) );
  AND2_X1 U16603 ( .A1(n14635), .A2(n21857), .ZN(n17710) );
  NAND2_X1 U16604 ( .A1(n17710), .A2(n14636), .ZN(n14763) );
  NOR2_X1 U16605 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n17676), .ZN(n17727) );
  AOI22_X1 U16606 ( .A1(n17736), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n17721), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n14637) );
  OAI21_X1 U16607 ( .B1(n16748), .B2(n14763), .A(n14637), .ZN(P2_U2927) );
  INV_X1 U16608 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n14682) );
  AOI22_X1 U16609 ( .A1(n17736), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n17721), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n14638) );
  OAI21_X1 U16610 ( .B1(n14682), .B2(n14763), .A(n14638), .ZN(P2_U2929) );
  INV_X1 U16611 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14679) );
  AOI22_X1 U16612 ( .A1(n17736), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n17721), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n14639) );
  OAI21_X1 U16613 ( .B1(n14679), .B2(n14763), .A(n14639), .ZN(P2_U2926) );
  INV_X1 U16614 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n16764) );
  AOI22_X1 U16615 ( .A1(n17736), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n17721), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n14640) );
  OAI21_X1 U16616 ( .B1(n16764), .B2(n14763), .A(n14640), .ZN(P2_U2930) );
  INV_X1 U16617 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n16756) );
  AOI22_X1 U16618 ( .A1(n17736), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n17721), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n14641) );
  OAI21_X1 U16619 ( .B1(n16756), .B2(n14763), .A(n14641), .ZN(P2_U2928) );
  INV_X1 U16620 ( .A(n14642), .ZN(n14675) );
  AOI22_X1 U16621 ( .A1(n19376), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n19375), .ZN(n16749) );
  INV_X1 U16622 ( .A(n16749), .ZN(n14643) );
  NAND2_X1 U16623 ( .A1(n14675), .A2(n14643), .ZN(n14688) );
  NAND2_X1 U16624 ( .A1(n14686), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n14645) );
  OAI211_X1 U16625 ( .C1(n14690), .C2(n16748), .A(n14688), .B(n14645), .ZN(
        P2_U2960) );
  INV_X1 U16626 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19373) );
  INV_X1 U16627 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n20227) );
  OR2_X1 U16628 ( .A1(n15647), .A2(n20227), .ZN(n14647) );
  NAND2_X1 U16629 ( .A1(n15647), .A2(BUF2_REG_9__SCAN_IN), .ZN(n14646) );
  NAND2_X1 U16630 ( .A1(n14647), .A2(n14646), .ZN(n19368) );
  NAND2_X1 U16631 ( .A1(n14675), .A2(n19368), .ZN(n14678) );
  NAND2_X1 U16632 ( .A1(n14686), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n14648) );
  OAI211_X1 U16633 ( .C1(n19373), .C2(n14690), .A(n14678), .B(n14648), .ZN(
        P2_U2976) );
  INV_X1 U16634 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n14652) );
  INV_X1 U16635 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n20234) );
  OR2_X1 U16636 ( .A1(n15647), .A2(n20234), .ZN(n14650) );
  NAND2_X1 U16637 ( .A1(n19375), .A2(BUF2_REG_13__SCAN_IN), .ZN(n14649) );
  NAND2_X1 U16638 ( .A1(n14650), .A2(n14649), .ZN(n16705) );
  NAND2_X1 U16639 ( .A1(n14675), .A2(n16705), .ZN(n14666) );
  NAND2_X1 U16640 ( .A1(n14686), .A2(P2_LWORD_REG_13__SCAN_IN), .ZN(n14651) );
  OAI211_X1 U16641 ( .C1(n14690), .C2(n14652), .A(n14666), .B(n14651), .ZN(
        P2_U2980) );
  INV_X1 U16642 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n17730) );
  INV_X1 U16643 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n20230) );
  OR2_X1 U16644 ( .A1(n15647), .A2(n20230), .ZN(n14654) );
  NAND2_X1 U16645 ( .A1(n15647), .A2(BUF2_REG_11__SCAN_IN), .ZN(n14653) );
  NAND2_X1 U16646 ( .A1(n14654), .A2(n14653), .ZN(n19364) );
  NAND2_X1 U16647 ( .A1(n14675), .A2(n19364), .ZN(n14670) );
  NAND2_X1 U16648 ( .A1(n14686), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n14655) );
  OAI211_X1 U16649 ( .C1(n17730), .C2(n14690), .A(n14670), .B(n14655), .ZN(
        P2_U2978) );
  INV_X1 U16650 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n14657) );
  AOI22_X1 U16651 ( .A1(n19376), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n19375), .ZN(n14939) );
  INV_X1 U16652 ( .A(n14939), .ZN(n16713) );
  NAND2_X1 U16653 ( .A1(n14675), .A2(n16713), .ZN(n14668) );
  NAND2_X1 U16654 ( .A1(n14686), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n14656) );
  OAI211_X1 U16655 ( .C1(n14690), .C2(n14657), .A(n14668), .B(n14656), .ZN(
        P2_U2979) );
  INV_X1 U16656 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n14659) );
  OAI22_X1 U16657 ( .A1(n19375), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n19376), .ZN(n19591) );
  INV_X1 U16658 ( .A(n19591), .ZN(n19580) );
  NAND2_X1 U16659 ( .A1(n14675), .A2(n19580), .ZN(n14681) );
  NAND2_X1 U16660 ( .A1(n14686), .A2(P2_LWORD_REG_6__SCAN_IN), .ZN(n14658) );
  OAI211_X1 U16661 ( .C1(n14690), .C2(n14659), .A(n14681), .B(n14658), .ZN(
        P2_U2973) );
  INV_X1 U16662 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n17734) );
  INV_X1 U16663 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n20236) );
  OR2_X1 U16664 ( .A1(n15647), .A2(n20236), .ZN(n14661) );
  NAND2_X1 U16665 ( .A1(n15647), .A2(BUF2_REG_14__SCAN_IN), .ZN(n14660) );
  NAND2_X1 U16666 ( .A1(n14661), .A2(n14660), .ZN(n19361) );
  NAND2_X1 U16667 ( .A1(n14675), .A2(n19361), .ZN(n14664) );
  NAND2_X1 U16668 ( .A1(n14686), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n14662) );
  OAI211_X1 U16669 ( .C1(n17734), .C2(n14690), .A(n14664), .B(n14662), .ZN(
        P2_U2981) );
  INV_X1 U16670 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n14759) );
  NAND2_X1 U16671 ( .A1(n14686), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n14663) );
  OAI211_X1 U16672 ( .C1(n14759), .C2(n14690), .A(n14664), .B(n14663), .ZN(
        P2_U2966) );
  INV_X1 U16673 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n16704) );
  NAND2_X1 U16674 ( .A1(n14686), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n14665) );
  OAI211_X1 U16675 ( .C1(n14690), .C2(n16704), .A(n14666), .B(n14665), .ZN(
        P2_U2965) );
  INV_X1 U16676 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n14753) );
  NAND2_X1 U16677 ( .A1(n14686), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n14667) );
  OAI211_X1 U16678 ( .C1(n14690), .C2(n14753), .A(n14668), .B(n14667), .ZN(
        P2_U2964) );
  INV_X1 U16679 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14751) );
  NAND2_X1 U16680 ( .A1(n14686), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n14669) );
  OAI211_X1 U16681 ( .C1(n14751), .C2(n14690), .A(n14670), .B(n14669), .ZN(
        P2_U2963) );
  INV_X1 U16682 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n16731) );
  INV_X1 U16683 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n14671) );
  OR2_X1 U16684 ( .A1(n15647), .A2(n14671), .ZN(n14673) );
  NAND2_X1 U16685 ( .A1(n15647), .A2(BUF2_REG_10__SCAN_IN), .ZN(n14672) );
  AND2_X1 U16686 ( .A1(n14673), .A2(n14672), .ZN(n16727) );
  INV_X1 U16687 ( .A(n16727), .ZN(n14674) );
  NAND2_X1 U16688 ( .A1(n14675), .A2(n14674), .ZN(n14684) );
  NAND2_X1 U16689 ( .A1(n14686), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n14676) );
  OAI211_X1 U16690 ( .C1(n14690), .C2(n16731), .A(n14684), .B(n14676), .ZN(
        P2_U2962) );
  NAND2_X1 U16691 ( .A1(n14686), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n14677) );
  OAI211_X1 U16692 ( .C1(n14679), .C2(n14690), .A(n14678), .B(n14677), .ZN(
        P2_U2961) );
  NAND2_X1 U16693 ( .A1(n14686), .A2(P2_UWORD_REG_6__SCAN_IN), .ZN(n14680) );
  OAI211_X1 U16694 ( .C1(n14690), .C2(n14682), .A(n14681), .B(n14680), .ZN(
        P2_U2958) );
  INV_X1 U16695 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n14685) );
  NAND2_X1 U16696 ( .A1(n14686), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n14683) );
  OAI211_X1 U16697 ( .C1(n14690), .C2(n14685), .A(n14684), .B(n14683), .ZN(
        P2_U2977) );
  INV_X1 U16698 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n14689) );
  NAND2_X1 U16699 ( .A1(n14686), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n14687) );
  OAI211_X1 U16700 ( .C1(n14690), .C2(n14689), .A(n14688), .B(n14687), .ZN(
        P2_U2975) );
  INV_X1 U16701 ( .A(n21513), .ZN(n14692) );
  OAI21_X1 U16702 ( .B1(n15837), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n14692), 
        .ZN(n14691) );
  OAI21_X1 U16703 ( .B1(n14693), .B2(n14692), .A(n14691), .ZN(P1_U3487) );
  INV_X1 U16704 ( .A(n14705), .ZN(n14694) );
  NAND2_X1 U16705 ( .A1(n14803), .A2(n14694), .ZN(n14697) );
  INV_X1 U16706 ( .A(n14695), .ZN(n14696) );
  NAND2_X1 U16707 ( .A1(n14697), .A2(n14696), .ZN(n14698) );
  OAI21_X1 U16708 ( .B1(n15175), .B2(n15156), .A(n14698), .ZN(n20201) );
  NAND3_X1 U16709 ( .A1(n14806), .A2(n21842), .A3(n11020), .ZN(n14699) );
  AND2_X1 U16710 ( .A1(n14699), .A2(n21834), .ZN(n21508) );
  OR2_X1 U16711 ( .A1(n20201), .A2(n21508), .ZN(n17375) );
  AND2_X1 U16712 ( .A1(n17375), .A2(n15174), .ZN(n21791) );
  INV_X1 U16713 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n17370) );
  NAND2_X1 U16714 ( .A1(n14700), .A2(n12558), .ZN(n14701) );
  OR2_X1 U16715 ( .A1(n14702), .A2(n14701), .ZN(n14703) );
  AND2_X1 U16716 ( .A1(n14704), .A2(n14703), .ZN(n14708) );
  NAND2_X1 U16717 ( .A1(n15175), .A2(n14862), .ZN(n14707) );
  NAND2_X1 U16718 ( .A1(n14803), .A2(n14705), .ZN(n14706) );
  OAI211_X1 U16719 ( .C1(n15175), .C2(n14708), .A(n14707), .B(n14706), .ZN(
        n14709) );
  NAND2_X1 U16720 ( .A1(n14709), .A2(n14811), .ZN(n17372) );
  INV_X1 U16721 ( .A(n17372), .ZN(n14710) );
  NAND2_X1 U16722 ( .A1(n21791), .A2(n14710), .ZN(n14711) );
  OAI21_X1 U16723 ( .B1(n21791), .B2(n17370), .A(n14711), .ZN(P1_U3484) );
  NAND2_X1 U16724 ( .A1(n15781), .A2(n15312), .ZN(n14713) );
  NAND2_X1 U16725 ( .A1(n11921), .A2(n18908), .ZN(n15325) );
  OR2_X1 U16726 ( .A1(n15328), .A2(n15325), .ZN(n14712) );
  NAND2_X1 U16727 ( .A1(n19374), .A2(n14715), .ZN(n15646) );
  OR2_X1 U16728 ( .A1(n15646), .A2(n14719), .ZN(n15427) );
  AOI21_X1 U16729 ( .B1(n14718), .B2(n14717), .A(n14716), .ZN(n17275) );
  INV_X1 U16730 ( .A(n17275), .ZN(n18628) );
  NAND2_X1 U16731 ( .A1(n19374), .A2(n14719), .ZN(n16771) );
  NAND2_X1 U16732 ( .A1(n19374), .A2(n19380), .ZN(n16765) );
  OAI222_X1 U16733 ( .A1(n15427), .A2(n19591), .B1(n18628), .B2(n19367), .C1(
        n14659), .C2(n19374), .ZN(P2_U2913) );
  OAI21_X1 U16734 ( .B1(n14722), .B2(n14721), .A(n14720), .ZN(n17687) );
  INV_X1 U16735 ( .A(n17687), .ZN(n18611) );
  OAI21_X1 U16736 ( .B1(n17229), .B2(n18611), .A(n14723), .ZN(n14729) );
  OAI211_X1 U16737 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n17262), .B(n16024), .ZN(n14726) );
  NAND2_X1 U16738 ( .A1(n18879), .A2(n14724), .ZN(n14725) );
  OAI211_X1 U16739 ( .C1(n14727), .C2(n18881), .A(n14726), .B(n14725), .ZN(
        n14728) );
  AOI211_X1 U16740 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n18877), .A(
        n14729), .B(n14728), .ZN(n14730) );
  OAI21_X1 U16741 ( .B1(n11489), .B2(n18885), .A(n14730), .ZN(P2_U3045) );
  NAND2_X1 U16742 ( .A1(n11969), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n14731) );
  AND4_X1 U16743 ( .A1(n14731), .A2(n19592), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n19459), .ZN(n14732) );
  OAI21_X1 U16744 ( .B1(n14736), .B2(n14735), .A(n14734), .ZN(n14737) );
  INV_X1 U16745 ( .A(n14737), .ZN(n18875) );
  NOR2_X1 U16746 ( .A1(n19455), .A2(n14737), .ZN(n14876) );
  INV_X1 U16747 ( .A(n14876), .ZN(n14738) );
  INV_X1 U16748 ( .A(n16771), .ZN(n19586) );
  OAI211_X1 U16749 ( .C1(n19467), .C2(n18875), .A(n14738), .B(n19586), .ZN(
        n14740) );
  AOI22_X1 U16750 ( .A1(n19585), .A2(n18875), .B1(n19579), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n14739) );
  OAI211_X1 U16751 ( .C1(n19838), .C2(n15427), .A(n14740), .B(n14739), .ZN(
        P2_U2919) );
  INV_X1 U16752 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n15738) );
  AOI22_X1 U16753 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n17735), .B1(n17736), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n14741) );
  OAI21_X1 U16754 ( .B1(n15738), .B2(n14763), .A(n14741), .ZN(P2_U2935) );
  INV_X1 U16755 ( .A(n14744), .ZN(n14742) );
  NAND2_X1 U16756 ( .A1(n14742), .A2(n15401), .ZN(n21951) );
  INV_X1 U16757 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n20045) );
  AND2_X1 U16758 ( .A1(n12599), .A2(n21841), .ZN(n14743) );
  NAND2_X1 U16759 ( .A1(n21949), .A2(n14745), .ZN(n21886) );
  INV_X1 U16760 ( .A(DATAI_15_), .ZN(n14747) );
  INV_X1 U16761 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n14746) );
  MUX2_X1 U16762 ( .A(n14747), .B(n14746), .S(n15942), .Z(n15939) );
  INV_X1 U16763 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n14748) );
  OAI222_X1 U16764 ( .A1(n21951), .A2(n20045), .B1(n21886), .B2(n15939), .C1(
        n21949), .C2(n14748), .ZN(P1_U2967) );
  AOI22_X1 U16765 ( .A1(n17736), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n17735), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n14749) );
  OAI21_X1 U16766 ( .B1(n16704), .B2(n14763), .A(n14749), .ZN(P2_U2922) );
  AOI22_X1 U16767 ( .A1(n17736), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n17735), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n14750) );
  OAI21_X1 U16768 ( .B1(n14751), .B2(n14763), .A(n14750), .ZN(P2_U2924) );
  AOI22_X1 U16769 ( .A1(n17736), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n17735), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n14752) );
  OAI21_X1 U16770 ( .B1(n14753), .B2(n14763), .A(n14752), .ZN(P2_U2923) );
  INV_X1 U16771 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n14755) );
  AOI22_X1 U16772 ( .A1(n17736), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n17735), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n14754) );
  OAI21_X1 U16773 ( .B1(n14755), .B2(n14763), .A(n14754), .ZN(P2_U2931) );
  AOI22_X1 U16774 ( .A1(n17736), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n17735), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n14756) );
  OAI21_X1 U16775 ( .B1(n16731), .B2(n14763), .A(n14756), .ZN(P2_U2925) );
  INV_X1 U16776 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n15747) );
  AOI22_X1 U16777 ( .A1(n17727), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n17735), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n14757) );
  OAI21_X1 U16778 ( .B1(n15747), .B2(n14763), .A(n14757), .ZN(P2_U2934) );
  AOI22_X1 U16779 ( .A1(n17727), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n17735), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n14758) );
  OAI21_X1 U16780 ( .B1(n14759), .B2(n14763), .A(n14758), .ZN(P2_U2921) );
  INV_X1 U16781 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n14761) );
  AOI22_X1 U16782 ( .A1(n17727), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n17735), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n14760) );
  OAI21_X1 U16783 ( .B1(n14761), .B2(n14763), .A(n14760), .ZN(P2_U2933) );
  INV_X1 U16784 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n15930) );
  AOI22_X1 U16785 ( .A1(n17727), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n17735), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n14762) );
  OAI21_X1 U16786 ( .B1(n15930), .B2(n14763), .A(n14762), .ZN(P2_U2932) );
  MUX2_X1 U16787 ( .A(n18884), .B(n14764), .S(n16689), .Z(n14765) );
  OAI21_X1 U16788 ( .B1(n19455), .B2(n16698), .A(n14765), .ZN(P2_U2887) );
  XOR2_X1 U16789 ( .A(n14767), .B(n14766), .Z(n17256) );
  INV_X1 U16790 ( .A(n17256), .ZN(n18640) );
  INV_X1 U16791 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n17724) );
  OAI222_X1 U16792 ( .A1(n15427), .A2(n19378), .B1(n18640), .B2(n19367), .C1(
        n17724), .C2(n19374), .ZN(P2_U2912) );
  INV_X1 U16793 ( .A(n14768), .ZN(n14769) );
  OAI21_X1 U16794 ( .B1(n14771), .B2(n14770), .A(n14769), .ZN(n18657) );
  OAI222_X1 U16795 ( .A1(n15427), .A2(n16749), .B1(n18657), .B2(n19367), .C1(
        n14689), .C2(n19374), .ZN(P2_U2911) );
  OAI21_X1 U16796 ( .B1(n14773), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n14772), .ZN(n20139) );
  INV_X1 U16797 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n16591) );
  AOI21_X1 U16798 ( .B1(n16591), .B2(n14775), .A(n16529), .ZN(n14774) );
  INV_X1 U16799 ( .A(n14774), .ZN(n14882) );
  OAI22_X1 U16800 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n14775), .B1(
        n16468), .B2(n14882), .ZN(n14781) );
  OAI21_X1 U16801 ( .B1(n14777), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n14776), .ZN(n15454) );
  INV_X1 U16802 ( .A(n15454), .ZN(n14779) );
  NAND2_X1 U16803 ( .A1(n21585), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n20142) );
  INV_X1 U16804 ( .A(n20142), .ZN(n14778) );
  AOI21_X1 U16805 ( .B1(n21595), .B2(n14779), .A(n14778), .ZN(n14780) );
  OAI211_X1 U16806 ( .C1(n16575), .C2(n20139), .A(n14781), .B(n14780), .ZN(
        P1_U3031) );
  OR2_X1 U16807 ( .A1(n14783), .A2(n14782), .ZN(n14784) );
  NOR2_X1 U16808 ( .A1(n11489), .A2(n16689), .ZN(n14786) );
  AOI21_X1 U16809 ( .B1(P2_EBX_REG_1__SCAN_IN), .B2(n16689), .A(n14786), .ZN(
        n14787) );
  OAI21_X1 U16810 ( .B1(n19408), .B2(n16698), .A(n14787), .ZN(P2_U2886) );
  MUX2_X1 U16811 ( .A(P2_EBX_REG_2__SCAN_IN), .B(n14791), .S(n16651), .Z(
        n14792) );
  AOI21_X1 U16812 ( .B1(n19502), .B2(n16686), .A(n14792), .ZN(n14793) );
  INV_X1 U16813 ( .A(n14793), .ZN(P2_U2885) );
  NAND2_X1 U16814 ( .A1(n14794), .A2(n14795), .ZN(n14796) );
  NAND2_X1 U16815 ( .A1(n14797), .A2(n14796), .ZN(n18669) );
  OAI222_X1 U16816 ( .A1(n15427), .A2(n16727), .B1(n18669), .B2(n19367), .C1(
        n14685), .C2(n19374), .ZN(P2_U2909) );
  INV_X1 U16817 ( .A(DATAI_0_), .ZN(n17455) );
  NAND2_X1 U16818 ( .A1(n15865), .A2(n17455), .ZN(n14799) );
  INV_X1 U16819 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n20209) );
  NAND2_X1 U16820 ( .A1(n15942), .A2(n20209), .ZN(n14798) );
  AND2_X1 U16821 ( .A1(n14799), .A2(n14798), .ZN(n15871) );
  INV_X1 U16822 ( .A(n15871), .ZN(n14817) );
  OAI21_X1 U16823 ( .B1(n14800), .B2(n21841), .A(n15217), .ZN(n14801) );
  NAND2_X1 U16824 ( .A1(n15175), .A2(n14801), .ZN(n14805) );
  NAND3_X1 U16825 ( .A1(n14803), .A2(n15401), .A3(n14802), .ZN(n14804) );
  OR2_X1 U16826 ( .A1(n14807), .A2(n14806), .ZN(n14808) );
  NAND2_X1 U16827 ( .A1(n10997), .A2(n14811), .ZN(n14812) );
  INV_X1 U16828 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20019) );
  NAND2_X2 U16829 ( .A1(n16273), .A2(n14812), .ZN(n16280) );
  NAND2_X1 U16830 ( .A1(n14814), .A2(n14813), .ZN(n14815) );
  NAND2_X1 U16831 ( .A1(n14816), .A2(n14815), .ZN(n20144) );
  OAI222_X1 U16832 ( .A1(n14817), .A2(n15944), .B1(n16273), .B2(n20019), .C1(
        n16280), .C2(n20144), .ZN(P1_U2904) );
  AOI22_X1 U16833 ( .A1(P1_EAX_REG_20__SCAN_IN), .A2(n14854), .B1(n21945), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n14820) );
  INV_X1 U16834 ( .A(DATAI_4_), .ZN(n17550) );
  NAND2_X1 U16835 ( .A1(n15865), .A2(n17550), .ZN(n14819) );
  INV_X1 U16836 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n20217) );
  NAND2_X1 U16837 ( .A1(n15942), .A2(n20217), .ZN(n14818) );
  AND2_X1 U16838 ( .A1(n14819), .A2(n14818), .ZN(n16288) );
  NAND2_X1 U16839 ( .A1(n21943), .A2(n16288), .ZN(n14833) );
  NAND2_X1 U16840 ( .A1(n14820), .A2(n14833), .ZN(P1_U2941) );
  AOI22_X1 U16841 ( .A1(P1_EAX_REG_16__SCAN_IN), .A2(n14854), .B1(n21945), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n14821) );
  NAND2_X1 U16842 ( .A1(n21943), .A2(n15871), .ZN(n14846) );
  NAND2_X1 U16843 ( .A1(n14821), .A2(n14846), .ZN(P1_U2937) );
  AOI22_X1 U16844 ( .A1(P1_EAX_REG_19__SCAN_IN), .A2(n14854), .B1(n21945), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n14824) );
  INV_X1 U16845 ( .A(DATAI_3_), .ZN(n17546) );
  NAND2_X1 U16846 ( .A1(n15865), .A2(n17546), .ZN(n14823) );
  INV_X1 U16847 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n20215) );
  NAND2_X1 U16848 ( .A1(n15942), .A2(n20215), .ZN(n14822) );
  AND2_X1 U16849 ( .A1(n14823), .A2(n14822), .ZN(n16291) );
  NAND2_X1 U16850 ( .A1(n21943), .A2(n16291), .ZN(n14831) );
  NAND2_X1 U16851 ( .A1(n14824), .A2(n14831), .ZN(P1_U2940) );
  AOI22_X1 U16852 ( .A1(P1_EAX_REG_1__SCAN_IN), .A2(n14854), .B1(n21945), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n14827) );
  INV_X1 U16853 ( .A(DATAI_1_), .ZN(n17453) );
  NAND2_X1 U16854 ( .A1(n15865), .A2(n17453), .ZN(n14826) );
  INV_X1 U16855 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n20211) );
  NAND2_X1 U16856 ( .A1(n15942), .A2(n20211), .ZN(n14825) );
  AND2_X1 U16857 ( .A1(n14826), .A2(n14825), .ZN(n15967) );
  NAND2_X1 U16858 ( .A1(n21943), .A2(n15967), .ZN(n14841) );
  NAND2_X1 U16859 ( .A1(n14827), .A2(n14841), .ZN(P1_U2953) );
  AOI22_X1 U16860 ( .A1(P1_EAX_REG_21__SCAN_IN), .A2(n14854), .B1(n21945), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n14830) );
  INV_X1 U16861 ( .A(DATAI_5_), .ZN(n17447) );
  NAND2_X1 U16862 ( .A1(n15865), .A2(n17447), .ZN(n14829) );
  INV_X1 U16863 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n20219) );
  NAND2_X1 U16864 ( .A1(n15942), .A2(n20219), .ZN(n14828) );
  AND2_X1 U16865 ( .A1(n14829), .A2(n14828), .ZN(n16285) );
  NAND2_X1 U16866 ( .A1(n21943), .A2(n16285), .ZN(n14850) );
  NAND2_X1 U16867 ( .A1(n14830), .A2(n14850), .ZN(P1_U2942) );
  AOI22_X1 U16868 ( .A1(P1_EAX_REG_3__SCAN_IN), .A2(n14854), .B1(n21945), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n14832) );
  NAND2_X1 U16869 ( .A1(n14832), .A2(n14831), .ZN(P1_U2955) );
  AOI22_X1 U16870 ( .A1(P1_EAX_REG_4__SCAN_IN), .A2(n14854), .B1(n21945), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n14834) );
  NAND2_X1 U16871 ( .A1(n14834), .A2(n14833), .ZN(P1_U2956) );
  AOI22_X1 U16872 ( .A1(P1_EAX_REG_18__SCAN_IN), .A2(n14854), .B1(n21945), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n14837) );
  INV_X1 U16873 ( .A(DATAI_2_), .ZN(n17452) );
  NAND2_X1 U16874 ( .A1(n15865), .A2(n17452), .ZN(n14836) );
  INV_X1 U16875 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n20213) );
  NAND2_X1 U16876 ( .A1(n15942), .A2(n20213), .ZN(n14835) );
  AND2_X1 U16877 ( .A1(n14836), .A2(n14835), .ZN(n16297) );
  NAND2_X1 U16878 ( .A1(n21943), .A2(n16297), .ZN(n14855) );
  NAND2_X1 U16879 ( .A1(n14837), .A2(n14855), .ZN(P1_U2939) );
  AOI22_X1 U16880 ( .A1(P1_EAX_REG_22__SCAN_IN), .A2(n14854), .B1(n21945), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n14840) );
  INV_X1 U16881 ( .A(DATAI_6_), .ZN(n17543) );
  NAND2_X1 U16882 ( .A1(n15865), .A2(n17543), .ZN(n14839) );
  INV_X1 U16883 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n20221) );
  NAND2_X1 U16884 ( .A1(n15942), .A2(n20221), .ZN(n14838) );
  AND2_X1 U16885 ( .A1(n14839), .A2(n14838), .ZN(n16281) );
  NAND2_X1 U16886 ( .A1(n21943), .A2(n16281), .ZN(n14852) );
  NAND2_X1 U16887 ( .A1(n14840), .A2(n14852), .ZN(P1_U2943) );
  AOI22_X1 U16888 ( .A1(P1_EAX_REG_17__SCAN_IN), .A2(n14854), .B1(n21945), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n14842) );
  NAND2_X1 U16889 ( .A1(n14842), .A2(n14841), .ZN(P1_U2938) );
  AOI22_X1 U16890 ( .A1(P1_EAX_REG_23__SCAN_IN), .A2(n14854), .B1(n21945), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n14845) );
  INV_X1 U16891 ( .A(DATAI_7_), .ZN(n17541) );
  NAND2_X1 U16892 ( .A1(n15865), .A2(n17541), .ZN(n14844) );
  INV_X1 U16893 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n20223) );
  NAND2_X1 U16894 ( .A1(n15942), .A2(n20223), .ZN(n14843) );
  AND2_X1 U16895 ( .A1(n14844), .A2(n14843), .ZN(n15531) );
  NAND2_X1 U16896 ( .A1(n21943), .A2(n15531), .ZN(n14848) );
  NAND2_X1 U16897 ( .A1(n14845), .A2(n14848), .ZN(P1_U2944) );
  AOI22_X1 U16898 ( .A1(P1_EAX_REG_0__SCAN_IN), .A2(n14854), .B1(n21945), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n14847) );
  NAND2_X1 U16899 ( .A1(n14847), .A2(n14846), .ZN(P1_U2952) );
  AOI22_X1 U16900 ( .A1(P1_EAX_REG_7__SCAN_IN), .A2(n14854), .B1(n21945), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n14849) );
  NAND2_X1 U16901 ( .A1(n14849), .A2(n14848), .ZN(P1_U2959) );
  AOI22_X1 U16902 ( .A1(P1_EAX_REG_5__SCAN_IN), .A2(n14854), .B1(n21945), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n14851) );
  NAND2_X1 U16903 ( .A1(n14851), .A2(n14850), .ZN(P1_U2957) );
  AOI22_X1 U16904 ( .A1(P1_EAX_REG_6__SCAN_IN), .A2(n14854), .B1(n21945), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n14853) );
  NAND2_X1 U16905 ( .A1(n14853), .A2(n14852), .ZN(P1_U2958) );
  AOI22_X1 U16906 ( .A1(P1_EAX_REG_2__SCAN_IN), .A2(n14854), .B1(n21945), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n14856) );
  NAND2_X1 U16907 ( .A1(n14856), .A2(n14855), .ZN(P1_U2954) );
  INV_X1 U16908 ( .A(n21794), .ZN(n14892) );
  AND2_X1 U16909 ( .A1(n15175), .A2(n17347), .ZN(n14857) );
  OAI211_X1 U16910 ( .C1(n17352), .C2(n12947), .A(n14857), .B(n21834), .ZN(
        n14859) );
  OAI211_X1 U16911 ( .C1(n15164), .C2(n14860), .A(n14859), .B(n14858), .ZN(
        n14861) );
  AOI21_X1 U16912 ( .B1(n14870), .B2(n14862), .A(n14861), .ZN(n14865) );
  INV_X1 U16913 ( .A(n14863), .ZN(n14864) );
  INV_X1 U16914 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n21790) );
  NAND2_X1 U16915 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n21803) );
  NOR3_X1 U16916 ( .A1(n21804), .A2(n21790), .A3(n21803), .ZN(n14867) );
  NOR2_X1 U16917 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n22072), .ZN(n14866) );
  AOI21_X1 U16918 ( .B1(n17352), .B2(n14892), .A(n21796), .ZN(n14873) );
  INV_X1 U16919 ( .A(n13136), .ZN(n15253) );
  NAND4_X1 U16920 ( .A1(n14869), .A2(n14868), .A3(n12562), .A4(n10996), .ZN(
        n15238) );
  INV_X1 U16921 ( .A(n15238), .ZN(n16586) );
  OAI22_X1 U16922 ( .A1(n15253), .A2(n16586), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n16585), .ZN(n17353) );
  INV_X1 U16923 ( .A(n21807), .ZN(n21792) );
  OAI22_X1 U16924 ( .A1(n21798), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21792), .ZN(n14871) );
  AOI21_X1 U16925 ( .B1(n17353), .B2(n14892), .A(n14871), .ZN(n14872) );
  OAI22_X1 U16926 ( .A1(n14873), .A2(n12447), .B1(n21796), .B2(n14872), .ZN(
        P1_U3474) );
  NOR2_X1 U16927 ( .A1(n19423), .A2(n17687), .ZN(n15366) );
  INV_X1 U16928 ( .A(n15366), .ZN(n14874) );
  OAI21_X1 U16929 ( .B1(n19408), .B2(n18611), .A(n14874), .ZN(n14875) );
  NOR2_X1 U16930 ( .A1(n14875), .A2(n14876), .ZN(n15365) );
  AOI21_X1 U16931 ( .B1(n14876), .B2(n14875), .A(n15365), .ZN(n14880) );
  AOI22_X1 U16932 ( .A1(n19585), .A2(n17687), .B1(n19579), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n14879) );
  INV_X1 U16933 ( .A(n19792), .ZN(n14877) );
  NAND2_X1 U16934 ( .A1(n19369), .A2(n14877), .ZN(n14878) );
  OAI211_X1 U16935 ( .C1(n14880), .C2(n16771), .A(n14879), .B(n14878), .ZN(
        P2_U2918) );
  NOR2_X1 U16936 ( .A1(n16490), .A2(n14881), .ZN(n14883) );
  MUX2_X1 U16937 ( .A(n14883), .B(n14882), .S(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n14884) );
  INV_X1 U16938 ( .A(n14884), .ZN(n14889) );
  OAI21_X1 U16939 ( .B1(n14887), .B2(n14886), .A(n14885), .ZN(n15534) );
  AOI22_X1 U16940 ( .A1(n21595), .A2(n15534), .B1(n16504), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n14888) );
  OAI211_X1 U16941 ( .C1(n14914), .C2(n16575), .A(n14889), .B(n14888), .ZN(
        P1_U3030) );
  INV_X1 U16942 ( .A(n21796), .ZN(n14895) );
  INV_X1 U16943 ( .A(n10996), .ZN(n15205) );
  INV_X1 U16944 ( .A(n15081), .ZN(n22062) );
  OR2_X1 U16945 ( .A1(n14890), .A2(n22062), .ZN(n14891) );
  XNOR2_X1 U16946 ( .A(n14891), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n21610) );
  NAND4_X1 U16947 ( .A1(n14895), .A2(n14892), .A3(n15205), .A4(n21610), .ZN(
        n14893) );
  OAI21_X1 U16948 ( .B1(n14895), .B2(n14894), .A(n14893), .ZN(P1_U3468) );
  XNOR2_X1 U16949 ( .A(n14897), .B(n14896), .ZN(n15122) );
  NAND3_X1 U16950 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21533), .A3(
        n12725), .ZN(n14902) );
  NAND2_X1 U16951 ( .A1(n16504), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n15119) );
  NAND2_X1 U16952 ( .A1(n21544), .A2(n14929), .ZN(n14925) );
  CLKBUF_X1 U16953 ( .A(n14898), .Z(n14931) );
  AOI21_X1 U16954 ( .B1(n14900), .B2(n14899), .A(n14931), .ZN(n15466) );
  NAND2_X1 U16955 ( .A1(n21595), .A2(n15466), .ZN(n14901) );
  AND4_X1 U16956 ( .A1(n14902), .A2(n15119), .A3(n14925), .A4(n14901), .ZN(
        n14906) );
  NAND2_X1 U16957 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14903) );
  OAI22_X1 U16958 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21531), .B1(
        n14903), .B2(n16453), .ZN(n14904) );
  OAI21_X1 U16959 ( .B1(n14904), .B2(n15616), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14905) );
  OAI211_X1 U16960 ( .C1(n15122), .C2(n16575), .A(n14906), .B(n14905), .ZN(
        P1_U3029) );
  INV_X1 U16961 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14912) );
  INV_X1 U16962 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n14907) );
  OAI22_X1 U16963 ( .A1(n20155), .A2(n14912), .B1(n21600), .B2(n14907), .ZN(
        n14911) );
  XNOR2_X1 U16964 ( .A(n14909), .B(n14908), .ZN(n15536) );
  NOR2_X1 U16965 ( .A1(n15536), .A2(n20194), .ZN(n14910) );
  AOI211_X1 U16966 ( .C1(n20172), .C2(n14912), .A(n14911), .B(n14910), .ZN(
        n14913) );
  OAI21_X1 U16967 ( .B1(n14914), .B2(n21789), .A(n14913), .ZN(P1_U2998) );
  NAND2_X1 U16968 ( .A1(n14916), .A2(n14915), .ZN(n14917) );
  NAND2_X1 U16969 ( .A1(n14941), .A2(n14917), .ZN(n14920) );
  INV_X1 U16970 ( .A(n19521), .ZN(n19426) );
  NOR2_X1 U16971 ( .A1(n15682), .A2(n16689), .ZN(n14921) );
  AOI21_X1 U16972 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n16689), .A(n14921), .ZN(
        n14922) );
  OAI21_X1 U16973 ( .B1(n19426), .B2(n16698), .A(n14922), .ZN(P2_U2884) );
  XNOR2_X1 U16974 ( .A(n10981), .B(n14923), .ZN(n15113) );
  INV_X1 U16975 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n16590) );
  NOR2_X1 U16976 ( .A1(n12725), .A2(n16590), .ZN(n14926) );
  OAI211_X1 U16977 ( .C1(n21531), .C2(n14926), .A(n21530), .B(n14925), .ZN(
        n15147) );
  INV_X1 U16978 ( .A(n14926), .ZN(n14928) );
  INV_X1 U16979 ( .A(n21533), .ZN(n14927) );
  OAI22_X1 U16980 ( .A1(n14929), .A2(n16453), .B1(n14928), .B2(n14927), .ZN(
        n15142) );
  AOI22_X1 U16981 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15147), .B1(
        n15142), .B2(n12728), .ZN(n14934) );
  OAI21_X1 U16982 ( .B1(n14931), .B2(n14930), .A(n15144), .ZN(n14932) );
  INV_X1 U16983 ( .A(n14932), .ZN(n20119) );
  AND2_X1 U16984 ( .A1(n21585), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n15109) );
  AOI21_X1 U16985 ( .B1(n21595), .B2(n20119), .A(n15109), .ZN(n14933) );
  OAI211_X1 U16986 ( .C1(n16575), .C2(n15113), .A(n14934), .B(n14933), .ZN(
        P1_U3028) );
  NOR2_X1 U16987 ( .A1(n14937), .A2(n14936), .ZN(n14938) );
  OR2_X1 U16988 ( .A1(n14935), .A2(n14938), .ZN(n18680) );
  OAI222_X1 U16989 ( .A1(n15427), .A2(n14939), .B1(n18680), .B2(n19367), .C1(
        n14657), .C2(n19374), .ZN(P2_U2907) );
  NAND2_X1 U16990 ( .A1(n14941), .A2(n14940), .ZN(n14943) );
  AND2_X1 U16991 ( .A1(n14943), .A2(n14942), .ZN(n14950) );
  NAND2_X1 U16992 ( .A1(n14945), .A2(n14944), .ZN(n14949) );
  OR2_X1 U16993 ( .A1(n14950), .A2(n14946), .ZN(n14948) );
  NAND2_X1 U16994 ( .A1(n14948), .A2(n14947), .ZN(n15071) );
  OAI21_X1 U16995 ( .B1(n14950), .B2(n14949), .A(n15071), .ZN(n15611) );
  XNOR2_X1 U16996 ( .A(n14952), .B(n14951), .ZN(n17621) );
  NOR2_X1 U16997 ( .A1(n17621), .A2(n16689), .ZN(n14953) );
  AOI21_X1 U16998 ( .B1(P2_EBX_REG_4__SCAN_IN), .B2(n16689), .A(n14953), .ZN(
        n14954) );
  OAI21_X1 U16999 ( .B1(n15611), .B2(n16698), .A(n14954), .ZN(P2_U2883) );
  XNOR2_X1 U17000 ( .A(n14955), .B(n14956), .ZN(n14961) );
  NAND2_X1 U17001 ( .A1(n14957), .A2(n14958), .ZN(n14959) );
  NAND2_X1 U17002 ( .A1(n15188), .A2(n14959), .ZN(n17650) );
  MUX2_X1 U17003 ( .A(n17650), .B(n11854), .S(n16689), .Z(n14960) );
  OAI21_X1 U17004 ( .B1(n14961), .B2(n16698), .A(n14960), .ZN(P2_U2878) );
  NAND2_X1 U17005 ( .A1(n15151), .A2(n14963), .ZN(n14964) );
  NAND2_X1 U17006 ( .A1(n14957), .A2(n14964), .ZN(n18652) );
  AND2_X1 U17007 ( .A1(n14966), .A2(n14965), .ZN(n14968) );
  OAI211_X1 U17008 ( .C1(n14968), .C2(n14967), .A(n14955), .B(n16686), .ZN(
        n14970) );
  NAND2_X1 U17009 ( .A1(n16689), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n14969) );
  OAI211_X1 U17010 ( .C1(n18652), .C2(n16689), .A(n14970), .B(n14969), .ZN(
        P2_U2879) );
  XOR2_X1 U17011 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n15071), .Z(n14976)
         );
  OAI21_X1 U17012 ( .B1(n14973), .B2(n14972), .A(n14971), .ZN(n17630) );
  MUX2_X1 U17013 ( .A(n14974), .B(n17630), .S(n16651), .Z(n14975) );
  OAI21_X1 U17014 ( .B1(n14976), .B2(n16698), .A(n14975), .ZN(P2_U2882) );
  NAND3_X1 U17015 ( .A1(n20971), .A2(n17389), .A3(n14977), .ZN(n14978) );
  NOR2_X1 U17016 ( .A1(n20801), .A2(n18069), .ZN(n18067) );
  INV_X1 U17017 ( .A(n18067), .ZN(n18072) );
  NOR2_X2 U17018 ( .A1(n18069), .A2(n20971), .ZN(n18070) );
  INV_X1 U17019 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n20685) );
  INV_X1 U17020 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n20659) );
  INV_X1 U17021 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n20632) );
  INV_X1 U17022 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n20579) );
  INV_X1 U17023 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n20544) );
  INV_X1 U17024 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n20518) );
  INV_X1 U17025 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n20510) );
  AND4_X1 U17026 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(P3_EBX_REG_2__SCAN_IN), 
        .A3(P3_EBX_REG_0__SCAN_IN), .A4(P3_EBX_REG_1__SCAN_IN), .ZN(n17773) );
  NAND2_X1 U17027 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17773), .ZN(n17795) );
  INV_X1 U17028 ( .A(n17795), .ZN(n17864) );
  INV_X1 U17029 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n20486) );
  INV_X1 U17030 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17901) );
  INV_X1 U17031 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n20431) );
  NAND4_X1 U17032 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(P3_EBX_REG_8__SCAN_IN), 
        .A3(P3_EBX_REG_6__SCAN_IN), .A4(P3_EBX_REG_5__SCAN_IN), .ZN(n14979) );
  NOR4_X1 U17033 ( .A1(n20486), .A2(n17901), .A3(n20431), .A4(n14979), .ZN(
        n17863) );
  NAND3_X1 U17034 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17864), .A3(n17863), 
        .ZN(n17828) );
  NOR4_X1 U17035 ( .A1(n20544), .A2(n20518), .A3(n20510), .A4(n17828), .ZN(
        n17805) );
  NAND2_X1 U17036 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17805), .ZN(n18064) );
  NOR2_X1 U17037 ( .A1(n20579), .A2(n18064), .ZN(n18063) );
  INV_X1 U17038 ( .A(n18063), .ZN(n14980) );
  NOR2_X1 U17039 ( .A1(n18069), .A2(n14980), .ZN(n18012) );
  NAND2_X1 U17040 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n18042), .ZN(n18041) );
  INV_X1 U17041 ( .A(n18041), .ZN(n18010) );
  NAND2_X1 U17042 ( .A1(n20971), .A2(n17936), .ZN(n17949) );
  NOR2_X1 U17043 ( .A1(n20632), .A2(n17949), .ZN(n17981) );
  NAND2_X1 U17044 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17981), .ZN(n17974) );
  NAND2_X1 U17045 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17980), .ZN(n15065) );
  NOR2_X1 U17046 ( .A1(n20685), .A2(n15065), .ZN(n17969) );
  NAND2_X1 U17047 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17969), .ZN(n17952) );
  NAND2_X1 U17048 ( .A1(n18043), .A2(n17952), .ZN(n17953) );
  OAI221_X1 U17049 ( .B1(n18072), .B2(P3_EBX_REG_28__SCAN_IN), .C1(n18072), 
        .C2(P3_EBX_REG_27__SCAN_IN), .A(n17953), .ZN(n15064) );
  AOI22_X1 U17050 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14984) );
  AOI22_X1 U17051 ( .A1(n11010), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17908), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14983) );
  AOI22_X1 U17052 ( .A1(n10956), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18013), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14982) );
  INV_X1 U17053 ( .A(n13801), .ZN(n17998) );
  AOI22_X1 U17054 ( .A1(n18025), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17998), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14981) );
  NAND4_X1 U17055 ( .A1(n14984), .A2(n14983), .A3(n14982), .A4(n14981), .ZN(
        n14990) );
  AOI22_X1 U17056 ( .A1(n17909), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14988) );
  AOI22_X1 U17057 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18046), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14987) );
  AOI22_X1 U17058 ( .A1(n17920), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18056), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14986) );
  AOI22_X1 U17059 ( .A1(n18033), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14985) );
  NAND4_X1 U17060 ( .A1(n14988), .A2(n14987), .A3(n14986), .A4(n14985), .ZN(
        n14989) );
  NOR2_X1 U17061 ( .A1(n14990), .A2(n14989), .ZN(n15063) );
  AOI22_X1 U17062 ( .A1(n17920), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14994) );
  AOI22_X1 U17063 ( .A1(n10957), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10967), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14993) );
  AOI22_X1 U17064 ( .A1(n18025), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17998), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14992) );
  AOI22_X1 U17065 ( .A1(n10956), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18013), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14991) );
  NAND4_X1 U17066 ( .A1(n14994), .A2(n14993), .A3(n14992), .A4(n14991), .ZN(
        n15000) );
  AOI22_X1 U17067 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17908), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14998) );
  AOI22_X1 U17068 ( .A1(n18031), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17890), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14997) );
  AOI22_X1 U17069 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18046), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14996) );
  AOI22_X1 U17070 ( .A1(n10971), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18056), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14995) );
  NAND4_X1 U17071 ( .A1(n14998), .A2(n14997), .A3(n14996), .A4(n14995), .ZN(
        n14999) );
  NOR2_X1 U17072 ( .A1(n15000), .A2(n14999), .ZN(n17950) );
  AOI22_X1 U17073 ( .A1(n18047), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15004) );
  AOI22_X1 U17074 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18032), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15003) );
  AOI22_X1 U17075 ( .A1(n18025), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17998), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15002) );
  AOI22_X1 U17076 ( .A1(n10956), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18013), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15001) );
  NAND4_X1 U17077 ( .A1(n15004), .A2(n15003), .A3(n15002), .A4(n15001), .ZN(
        n15010) );
  AOI22_X1 U17078 ( .A1(n17909), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17920), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15008) );
  AOI22_X1 U17079 ( .A1(n18031), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18046), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15007) );
  AOI22_X1 U17080 ( .A1(n18033), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15006) );
  AOI22_X1 U17081 ( .A1(n11010), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17908), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15005) );
  NAND4_X1 U17082 ( .A1(n15008), .A2(n15007), .A3(n15006), .A4(n15005), .ZN(
        n15009) );
  NOR2_X1 U17083 ( .A1(n15010), .A2(n15009), .ZN(n17966) );
  AOI22_X1 U17084 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18046), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15014) );
  AOI22_X1 U17085 ( .A1(n10957), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17890), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15013) );
  AOI22_X1 U17086 ( .A1(n10956), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18013), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15012) );
  AOI22_X1 U17087 ( .A1(n18025), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17998), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15011) );
  NAND4_X1 U17088 ( .A1(n15014), .A2(n15013), .A3(n15012), .A4(n15011), .ZN(
        n15020) );
  AOI22_X1 U17089 ( .A1(n18047), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15018) );
  AOI22_X1 U17090 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15017) );
  AOI22_X1 U17091 ( .A1(n10971), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18032), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15016) );
  AOI22_X1 U17092 ( .A1(n17920), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17908), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15015) );
  NAND4_X1 U17093 ( .A1(n15018), .A2(n15017), .A3(n15016), .A4(n15015), .ZN(
        n15019) );
  NOR2_X1 U17094 ( .A1(n15020), .A2(n15019), .ZN(n17976) );
  AOI22_X1 U17095 ( .A1(n17920), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17890), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15024) );
  AOI22_X1 U17096 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15023) );
  AOI22_X1 U17097 ( .A1(n18025), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18013), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15022) );
  AOI22_X1 U17098 ( .A1(n10956), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17998), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15021) );
  NAND4_X1 U17099 ( .A1(n15024), .A2(n15023), .A3(n15022), .A4(n15021), .ZN(
        n15030) );
  AOI22_X1 U17100 ( .A1(n17909), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n18047), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15028) );
  AOI22_X1 U17101 ( .A1(n18031), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15027) );
  AOI22_X1 U17102 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17908), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15026) );
  AOI22_X1 U17103 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18046), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15025) );
  NAND4_X1 U17104 ( .A1(n15028), .A2(n15027), .A3(n15026), .A4(n15025), .ZN(
        n15029) );
  NOR2_X1 U17105 ( .A1(n15030), .A2(n15029), .ZN(n17977) );
  NOR2_X1 U17106 ( .A1(n17976), .A2(n17977), .ZN(n17975) );
  AOI22_X1 U17107 ( .A1(n10957), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n10969), .ZN(n15041) );
  AOI22_X1 U17108 ( .A1(n18031), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n18045), .ZN(n15040) );
  AOI22_X1 U17109 ( .A1(n18047), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n18046), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15031) );
  OAI21_X1 U17110 ( .B1(n15032), .B2(n15053), .A(n15031), .ZN(n15038) );
  AOI22_X1 U17111 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n10971), .B1(
        n18054), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n15036) );
  AOI22_X1 U17112 ( .A1(n17920), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n18056), .ZN(n15035) );
  AOI22_X1 U17113 ( .A1(n18025), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17998), .ZN(n15034) );
  AOI22_X1 U17114 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n13835), .B1(
        n10956), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15033) );
  NAND4_X1 U17115 ( .A1(n15036), .A2(n15035), .A3(n15034), .A4(n15033), .ZN(
        n15037) );
  AOI211_X1 U17116 ( .C1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .C2(n11010), .A(
        n15038), .B(n15037), .ZN(n15039) );
  NAND3_X1 U17117 ( .A1(n15041), .A2(n15040), .A3(n15039), .ZN(n17971) );
  NAND2_X1 U17118 ( .A1(n17975), .A2(n17971), .ZN(n17970) );
  NOR2_X1 U17119 ( .A1(n17966), .A2(n17970), .ZN(n17965) );
  AOI22_X1 U17120 ( .A1(n18047), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15051) );
  AOI22_X1 U17121 ( .A1(n13837), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15050) );
  AOI22_X1 U17122 ( .A1(n18031), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17908), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15042) );
  OAI21_X1 U17123 ( .B1(n15053), .B2(n17778), .A(n15042), .ZN(n15048) );
  AOI22_X1 U17124 ( .A1(n10967), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18046), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15046) );
  AOI22_X1 U17125 ( .A1(n17920), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18032), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15045) );
  AOI22_X1 U17126 ( .A1(n10956), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17998), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15044) );
  AOI22_X1 U17127 ( .A1(n18025), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18013), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15043) );
  NAND4_X1 U17128 ( .A1(n15046), .A2(n15045), .A3(n15044), .A4(n15043), .ZN(
        n15047) );
  AOI211_X1 U17129 ( .C1(n10957), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n15048), .B(n15047), .ZN(n15049) );
  NAND3_X1 U17130 ( .A1(n15051), .A2(n15050), .A3(n15049), .ZN(n17962) );
  NAND2_X1 U17131 ( .A1(n17965), .A2(n17962), .ZN(n17961) );
  NOR2_X1 U17132 ( .A1(n17950), .A2(n17961), .ZN(n17958) );
  AOI22_X1 U17133 ( .A1(n17920), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15062) );
  AOI22_X1 U17134 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n18032), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15061) );
  AOI22_X1 U17135 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17908), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15052) );
  OAI21_X1 U17136 ( .B1(n15053), .B2(n17835), .A(n15052), .ZN(n15059) );
  AOI22_X1 U17137 ( .A1(n18047), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15057) );
  AOI22_X1 U17138 ( .A1(n18031), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n18046), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15056) );
  AOI22_X1 U17139 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17998), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15055) );
  AOI22_X1 U17140 ( .A1(n18025), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18013), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15054) );
  NAND4_X1 U17141 ( .A1(n15057), .A2(n15056), .A3(n15055), .A4(n15054), .ZN(
        n15058) );
  AOI211_X1 U17142 ( .C1(n17909), .C2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n15059), .B(n15058), .ZN(n15060) );
  NAND3_X1 U17143 ( .A1(n15062), .A2(n15061), .A3(n15060), .ZN(n17957) );
  NAND2_X1 U17144 ( .A1(n17958), .A2(n17957), .ZN(n17956) );
  NOR2_X1 U17145 ( .A1(n15063), .A2(n17956), .ZN(n17932) );
  AOI21_X1 U17146 ( .B1(n15063), .B2(n17956), .A(n17932), .ZN(n20916) );
  AOI22_X1 U17147 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n15064), .B1(n20916), 
        .B2(n18070), .ZN(n15069) );
  INV_X1 U17148 ( .A(n15065), .ZN(n17973) );
  INV_X1 U17149 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n15067) );
  INV_X1 U17150 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n20710) );
  INV_X1 U17151 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n20699) );
  NOR3_X1 U17152 ( .A1(n20710), .A2(n20699), .A3(n20685), .ZN(n17955) );
  NAND2_X1 U17153 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17955), .ZN(n15972) );
  INV_X1 U17154 ( .A(n15972), .ZN(n15066) );
  NAND3_X1 U17155 ( .A1(n17973), .A2(n15067), .A3(n15066), .ZN(n15068) );
  NAND2_X1 U17156 ( .A1(n15069), .A2(n15068), .ZN(P3_U2674) );
  NOR2_X1 U17157 ( .A1(n15071), .A2(n12100), .ZN(n15072) );
  OR2_X1 U17158 ( .A1(n15071), .A2(n15070), .ZN(n15150) );
  OAI211_X1 U17159 ( .C1(n15072), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n16686), .B(n15150), .ZN(n15078) );
  AND2_X1 U17160 ( .A1(n14971), .A2(n15073), .ZN(n15075) );
  OR2_X1 U17161 ( .A1(n15075), .A2(n15074), .ZN(n18627) );
  INV_X1 U17162 ( .A(n18627), .ZN(n15076) );
  NAND2_X1 U17163 ( .A1(n15076), .A2(n16651), .ZN(n15077) );
  OAI211_X1 U17164 ( .C1(n16651), .C2(n11844), .A(n15078), .B(n15077), .ZN(
        P2_U2881) );
  NAND3_X1 U17165 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n22105), .A3(
        n22066), .ZN(n15803) );
  NOR2_X1 U17166 ( .A1(n22076), .A2(n15803), .ZN(n15083) );
  INV_X1 U17167 ( .A(n15083), .ZN(n15442) );
  NOR2_X2 U17168 ( .A1(n15412), .A2(n15867), .ZN(n22391) );
  INV_X1 U17169 ( .A(n22391), .ZN(n15828) );
  INV_X1 U17170 ( .A(n15803), .ZN(n15090) );
  OAI21_X1 U17171 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n22072), .A(
        n15415), .ZN(n21992) );
  INV_X1 U17172 ( .A(n21955), .ZN(n15080) );
  INV_X1 U17173 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n15084) );
  OR2_X1 U17174 ( .A1(n22063), .A2(n15081), .ZN(n22002) );
  INV_X1 U17175 ( .A(n22002), .ZN(n15806) );
  INV_X1 U17176 ( .A(n15082), .ZN(n22077) );
  AOI21_X1 U17177 ( .B1(n15806), .B2(n22077), .A(n15083), .ZN(n15088) );
  OAI211_X1 U17178 ( .C1(n15124), .C2(n15084), .A(n22059), .B(n15088), .ZN(
        n15085) );
  OAI211_X1 U17179 ( .C1(n22059), .C2(n15090), .A(n22113), .B(n15085), .ZN(
        n15437) );
  NAND2_X1 U17180 ( .A1(n15437), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n15095) );
  INV_X1 U17181 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20270) );
  INV_X1 U17182 ( .A(DATAI_31_), .ZN(n15086) );
  OAI22_X1 U17183 ( .A1(n20270), .A2(n15414), .B1(n15086), .B2(n15413), .ZN(
        n22383) );
  INV_X1 U17184 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n20253) );
  INV_X1 U17185 ( .A(DATAI_23_), .ZN(n17495) );
  OAI22_X1 U17186 ( .A1(n20253), .A2(n15414), .B1(n17495), .B2(n15413), .ZN(
        n22392) );
  NAND2_X1 U17187 ( .A1(n15415), .A2(n15531), .ZN(n22373) );
  INV_X1 U17188 ( .A(n15088), .ZN(n15089) );
  NAND2_X1 U17189 ( .A1(n15089), .A2(n22117), .ZN(n15092) );
  NAND2_X1 U17190 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n15090), .ZN(n15091) );
  NAND2_X1 U17191 ( .A1(n15092), .A2(n15091), .ZN(n15201) );
  OAI22_X1 U17192 ( .A1(n22010), .A2(n11077), .B1(n22373), .B2(n15438), .ZN(
        n15093) );
  AOI21_X1 U17193 ( .B1(n11060), .B2(n15805), .A(n15093), .ZN(n15094) );
  OAI211_X1 U17194 ( .C1(n15442), .C2(n15828), .A(n15095), .B(n15094), .ZN(
        P1_U3080) );
  INV_X1 U17195 ( .A(n22212), .ZN(n15832) );
  NAND2_X1 U17196 ( .A1(n15437), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n15099) );
  INV_X1 U17197 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20262) );
  INV_X1 U17198 ( .A(DATAI_27_), .ZN(n17500) );
  OAI22_X1 U17199 ( .A1(n20262), .A2(n15414), .B1(n17500), .B2(n15413), .ZN(
        n22208) );
  INV_X1 U17200 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20245) );
  INV_X1 U17201 ( .A(DATAI_19_), .ZN(n17492) );
  OAI22_X1 U17202 ( .A1(n20245), .A2(n15414), .B1(n17492), .B2(n15413), .ZN(
        n22213) );
  NAND2_X1 U17203 ( .A1(n15415), .A2(n16291), .ZN(n22205) );
  OAI22_X1 U17204 ( .A1(n22010), .A2(n11073), .B1(n22205), .B2(n15438), .ZN(
        n15097) );
  AOI21_X1 U17205 ( .B1(n11068), .B2(n15805), .A(n15097), .ZN(n15098) );
  OAI211_X1 U17206 ( .C1(n15442), .C2(n15832), .A(n15099), .B(n15098), .ZN(
        P1_U3076) );
  NOR2_X2 U17207 ( .A1(n15412), .A2(n12559), .ZN(n22180) );
  INV_X1 U17208 ( .A(n22180), .ZN(n15852) );
  NAND2_X1 U17209 ( .A1(n15437), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n15103) );
  INV_X1 U17210 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20260) );
  INV_X1 U17211 ( .A(DATAI_26_), .ZN(n17510) );
  INV_X1 U17212 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20243) );
  INV_X1 U17213 ( .A(DATAI_18_), .ZN(n15100) );
  INV_X1 U17214 ( .A(n22181), .ZN(n22178) );
  NAND2_X1 U17215 ( .A1(n15415), .A2(n16297), .ZN(n22172) );
  OAI22_X1 U17216 ( .A1(n22010), .A2(n22178), .B1(n22172), .B2(n15438), .ZN(
        n15101) );
  AOI21_X1 U17217 ( .B1(n22175), .B2(n15805), .A(n15101), .ZN(n15102) );
  OAI211_X1 U17218 ( .C1(n15442), .C2(n15852), .A(n15103), .B(n15102), .ZN(
        P1_U3075) );
  AOI22_X1 U17219 ( .A1(n15920), .A2(n15967), .B1(P1_EAX_REG_1__SCAN_IN), .B2(
        n16248), .ZN(n15104) );
  OAI21_X1 U17220 ( .B1(n16280), .B2(n15536), .A(n15104), .ZN(P1_U2903) );
  OR2_X1 U17221 ( .A1(n15107), .A2(n15106), .ZN(n15108) );
  AND2_X1 U17222 ( .A1(n15105), .A2(n15108), .ZN(n20120) );
  AOI21_X1 U17223 ( .B1(n20192), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n15109), .ZN(n15110) );
  OAI21_X1 U17224 ( .B1(n20200), .B2(n15160), .A(n15110), .ZN(n15111) );
  AOI21_X1 U17225 ( .B1(n20120), .B2(n20186), .A(n15111), .ZN(n15112) );
  OAI21_X1 U17226 ( .B1(n15113), .B2(n21789), .A(n15112), .ZN(P1_U2996) );
  INV_X1 U17227 ( .A(n15114), .ZN(n15115) );
  AOI21_X1 U17228 ( .B1(n15117), .B2(n15116), .A(n15115), .ZN(n15351) );
  NAND2_X1 U17229 ( .A1(n20192), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n15118) );
  OAI211_X1 U17230 ( .C1(n20200), .C2(n15360), .A(n15119), .B(n15118), .ZN(
        n15120) );
  AOI21_X1 U17231 ( .B1(n15351), .B2(n20186), .A(n15120), .ZN(n15121) );
  OAI21_X1 U17232 ( .B1(n21789), .B2(n15122), .A(n15121), .ZN(P1_U2997) );
  NOR2_X2 U17233 ( .A1(n15412), .A2(n12966), .ZN(n22109) );
  INV_X1 U17234 ( .A(n22109), .ZN(n15860) );
  NAND2_X1 U17235 ( .A1(n15087), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n22111) );
  NOR3_X1 U17236 ( .A1(n15124), .A2(n22115), .A3(n22111), .ZN(n16579) );
  NOR2_X1 U17237 ( .A1(n22104), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n15127) );
  OAI21_X1 U17238 ( .B1(n16579), .B2(n15127), .A(n22113), .ZN(n15419) );
  NAND2_X1 U17239 ( .A1(n15419), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n15133) );
  NOR2_X2 U17240 ( .A1(n15124), .A2(n22054), .ZN(n22344) );
  INV_X1 U17241 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20239) );
  INV_X1 U17242 ( .A(DATAI_16_), .ZN(n17522) );
  OAI22_X1 U17243 ( .A1(n20239), .A2(n15414), .B1(n17522), .B2(n15413), .ZN(
        n22118) );
  INV_X1 U17244 ( .A(DATAI_24_), .ZN(n17503) );
  INV_X1 U17245 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20255) );
  OAI22_X1 U17246 ( .A1(n17503), .A2(n15413), .B1(n20255), .B2(n15414), .ZN(
        n22096) );
  NAND2_X1 U17247 ( .A1(n15415), .A2(n15871), .ZN(n22075) );
  NAND2_X1 U17248 ( .A1(n10993), .A2(n13136), .ZN(n22100) );
  OAI21_X1 U17249 ( .B1(n22002), .B2(n22100), .A(n15421), .ZN(n15126) );
  NAND2_X1 U17250 ( .A1(n15126), .A2(n22059), .ZN(n15129) );
  NAND2_X1 U17251 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n15127), .ZN(n15128) );
  NAND2_X1 U17252 ( .A1(n15129), .A2(n15128), .ZN(n15416) );
  INV_X1 U17253 ( .A(n15416), .ZN(n15130) );
  OAI22_X1 U17254 ( .A1(n21999), .A2(n11069), .B1(n22075), .B2(n15130), .ZN(
        n15131) );
  AOI21_X1 U17255 ( .B1(n22344), .B2(n11072), .A(n15131), .ZN(n15132) );
  OAI211_X1 U17256 ( .C1(n15860), .C2(n15421), .A(n15133), .B(n15132), .ZN(
        P1_U3089) );
  NOR2_X1 U17257 ( .A1(n14935), .A2(n15135), .ZN(n15136) );
  OR2_X1 U17258 ( .A1(n15134), .A2(n15136), .ZN(n17161) );
  AOI22_X1 U17259 ( .A1(n19369), .A2(n16705), .B1(P2_EAX_REG_13__SCAN_IN), 
        .B2(n19579), .ZN(n15137) );
  OAI21_X1 U17260 ( .B1(n19367), .B2(n17161), .A(n15137), .ZN(P2_U2906) );
  INV_X1 U17261 ( .A(n16297), .ZN(n15138) );
  INV_X1 U17262 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20023) );
  INV_X1 U17263 ( .A(n15351), .ZN(n15468) );
  OAI222_X1 U17264 ( .A1(n15138), .A2(n15944), .B1(n16273), .B2(n20023), .C1(
        n16280), .C2(n15468), .ZN(P1_U2902) );
  XNOR2_X1 U17265 ( .A(n15139), .B(n15140), .ZN(n15381) );
  OAI211_X1 U17266 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n15142), .B(n15141), .ZN(n15149) );
  INV_X1 U17267 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21621) );
  NOR2_X1 U17268 ( .A1(n21600), .A2(n21621), .ZN(n15376) );
  INV_X1 U17269 ( .A(n20132), .ZN(n15143) );
  AOI21_X1 U17270 ( .B1(n15145), .B2(n15144), .A(n15143), .ZN(n21611) );
  INV_X1 U17271 ( .A(n21611), .ZN(n15575) );
  NOR2_X1 U17272 ( .A1(n21560), .A2(n15575), .ZN(n15146) );
  AOI211_X1 U17273 ( .C1(n15147), .C2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n15376), .B(n15146), .ZN(n15148) );
  OAI211_X1 U17274 ( .C1(n16575), .C2(n15381), .A(n15149), .B(n15148), .ZN(
        P1_U3027) );
  XOR2_X1 U17275 ( .A(n15150), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n15154)
         );
  OAI21_X1 U17276 ( .B1(n15074), .B2(n15152), .A(n15151), .ZN(n18639) );
  MUX2_X1 U17277 ( .A(n12189), .B(n18639), .S(n16651), .Z(n15153) );
  OAI21_X1 U17278 ( .B1(n15154), .B2(n16698), .A(n15153), .ZN(P2_U2880) );
  INV_X1 U17279 ( .A(n15163), .ZN(n15155) );
  NAND2_X1 U17280 ( .A1(n15156), .A2(n15155), .ZN(n15157) );
  NAND2_X1 U17281 ( .A1(n21777), .A2(n15157), .ZN(n21631) );
  INV_X1 U17282 ( .A(n21631), .ZN(n15393) );
  INV_X1 U17283 ( .A(n20120), .ZN(n15172) );
  INV_X1 U17284 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20049) );
  INV_X1 U17285 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20047) );
  INV_X1 U17286 ( .A(n21622), .ZN(n15158) );
  NAND2_X1 U17287 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n15158), .ZN(n15354) );
  OAI22_X1 U17288 ( .A1(n21710), .A2(n20049), .B1(n20047), .B2(n15354), .ZN(
        n15159) );
  NAND4_X1 U17289 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(n15158), .ZN(n21620) );
  NAND2_X1 U17290 ( .A1(n15159), .A2(n21620), .ZN(n15171) );
  INV_X1 U17291 ( .A(n15160), .ZN(n15169) );
  AOI22_X1 U17292 ( .A1(n20119), .A2(n21724), .B1(n21773), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n15166) );
  NOR2_X1 U17293 ( .A1(n15164), .A2(n15163), .ZN(n21609) );
  NAND2_X1 U17294 ( .A1(n22015), .A2(n21609), .ZN(n15165) );
  OAI211_X1 U17295 ( .C1(n21776), .C2(n15167), .A(n15166), .B(n15165), .ZN(
        n15168) );
  AOI21_X1 U17296 ( .B1(n15169), .B2(n21782), .A(n15168), .ZN(n15170) );
  OAI211_X1 U17297 ( .C1(n15393), .C2(n15172), .A(n15171), .B(n15170), .ZN(
        P1_U2837) );
  INV_X1 U17298 ( .A(n16291), .ZN(n15173) );
  INV_X1 U17299 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20025) );
  OAI222_X1 U17300 ( .A1(n15173), .A2(n15944), .B1(n16273), .B2(n20025), .C1(
        n16280), .C2(n15172), .ZN(P1_U2901) );
  INV_X1 U17301 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n15180) );
  NAND3_X1 U17302 ( .A1(n15175), .A2(n15174), .A3(n17352), .ZN(n15176) );
  NAND2_X1 U17303 ( .A1(n21951), .A2(n15176), .ZN(n15177) );
  NOR2_X1 U17304 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21803), .ZN(n20031) );
  NOR2_X4 U17305 ( .A1(n20017), .A2(n21515), .ZN(n20034) );
  AOI22_X1 U17306 ( .A1(n20031), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n15179) );
  OAI21_X1 U17307 ( .B1(n15180), .B2(n15555), .A(n15179), .ZN(P1_U2919) );
  INV_X1 U17308 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n15182) );
  AOI22_X1 U17309 ( .A1(n21515), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n15181) );
  OAI21_X1 U17310 ( .B1(n15182), .B2(n15555), .A(n15181), .ZN(P1_U2918) );
  XNOR2_X1 U17311 ( .A(n15183), .B(n15184), .ZN(n15186) );
  MUX2_X1 U17312 ( .A(n17190), .B(n11862), .S(n16689), .Z(n15185) );
  OAI21_X1 U17313 ( .B1(n15186), .B2(n16698), .A(n15185), .ZN(P2_U2876) );
  AOI21_X1 U17314 ( .B1(n15189), .B2(n15188), .A(n15187), .ZN(n18665) );
  INV_X1 U17315 ( .A(n18665), .ZN(n15196) );
  INV_X1 U17316 ( .A(n15190), .ZN(n15193) );
  INV_X1 U17317 ( .A(n15183), .ZN(n15191) );
  OAI211_X1 U17318 ( .C1(n15193), .C2(n15192), .A(n15191), .B(n16686), .ZN(
        n15195) );
  NAND2_X1 U17319 ( .A1(n16689), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n15194) );
  OAI211_X1 U17320 ( .C1(n15196), .C2(n16689), .A(n15195), .B(n15194), .ZN(
        P2_U2877) );
  AND2_X1 U17321 ( .A1(n15105), .A2(n15198), .ZN(n15199) );
  OR2_X1 U17322 ( .A1(n15197), .A2(n15199), .ZN(n21607) );
  INV_X1 U17323 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20027) );
  INV_X1 U17324 ( .A(n16288), .ZN(n15200) );
  OAI222_X1 U17325 ( .A1(n21607), .A2(n16280), .B1(n16273), .B2(n20027), .C1(
        n15200), .C2(n15944), .ZN(P1_U2900) );
  AOI22_X1 U17326 ( .A1(n15805), .A2(n11070), .B1(n22108), .B2(n15201), .ZN(
        n15202) );
  OAI21_X1 U17327 ( .B1(n22010), .B2(n11071), .A(n15202), .ZN(n15203) );
  AOI21_X1 U17328 ( .B1(n15437), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A(
        n15203), .ZN(n15204) );
  OAI21_X1 U17329 ( .B1(n15860), .B2(n15442), .A(n15204), .ZN(P1_U3073) );
  NAND2_X1 U17330 ( .A1(n21610), .A2(n15205), .ZN(n15206) );
  NAND2_X1 U17331 ( .A1(n17356), .A2(n15206), .ZN(n15207) );
  OAI211_X1 U17332 ( .C1(n17356), .C2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n15207), .B(n21798), .ZN(n15210) );
  NAND2_X1 U17333 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21790), .ZN(n15244) );
  INV_X1 U17334 ( .A(n15244), .ZN(n15208) );
  NAND2_X1 U17335 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15208), .ZN(
        n15209) );
  INV_X1 U17336 ( .A(n15212), .ZN(n15243) );
  OR2_X1 U17337 ( .A1(n17356), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15225) );
  OR2_X1 U17338 ( .A1(n22063), .A2(n16586), .ZN(n15223) );
  INV_X1 U17339 ( .A(n15213), .ZN(n15214) );
  NAND2_X1 U17340 ( .A1(n15214), .A2(n12445), .ZN(n15231) );
  NAND2_X1 U17341 ( .A1(n15213), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15226) );
  AND2_X1 U17342 ( .A1(n15231), .A2(n15226), .ZN(n16596) );
  NAND3_X1 U17343 ( .A1(n16586), .A2(n15215), .A3(n16596), .ZN(n15221) );
  XNOR2_X1 U17344 ( .A(n12445), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15219) );
  NAND2_X1 U17345 ( .A1(n15217), .A2(n15216), .ZN(n15233) );
  INV_X1 U17346 ( .A(n16596), .ZN(n15218) );
  AOI22_X1 U17347 ( .A1(n17352), .A2(n15219), .B1(n15233), .B2(n15218), .ZN(
        n15220) );
  AND2_X1 U17348 ( .A1(n15221), .A2(n15220), .ZN(n15222) );
  AND2_X1 U17349 ( .A1(n15223), .A2(n15222), .ZN(n16600) );
  NAND2_X1 U17350 ( .A1(n17356), .A2(n16600), .ZN(n15224) );
  NAND2_X1 U17351 ( .A1(n15225), .A2(n15224), .ZN(n17363) );
  INV_X1 U17352 ( .A(n17363), .ZN(n15241) );
  OR2_X1 U17353 ( .A1(n17356), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n15240) );
  AND2_X1 U17354 ( .A1(n15226), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n15227) );
  NOR2_X1 U17355 ( .A1(n12685), .A2(n15227), .ZN(n21793) );
  OR2_X1 U17356 ( .A1(n15228), .A2(n21793), .ZN(n15236) );
  XNOR2_X1 U17357 ( .A(n15229), .B(n11209), .ZN(n15230) );
  NAND2_X1 U17358 ( .A1(n17352), .A2(n15230), .ZN(n15235) );
  XNOR2_X1 U17359 ( .A(n15231), .B(n11209), .ZN(n15232) );
  NAND2_X1 U17360 ( .A1(n15233), .A2(n15232), .ZN(n15234) );
  OAI211_X1 U17361 ( .C1(n15238), .C2(n15236), .A(n15235), .B(n15234), .ZN(
        n15237) );
  AOI21_X1 U17362 ( .B1(n22015), .B2(n15238), .A(n15237), .ZN(n21795) );
  NAND2_X1 U17363 ( .A1(n17356), .A2(n21795), .ZN(n15239) );
  NAND3_X1 U17364 ( .A1(n15241), .A2(n17365), .A3(n21798), .ZN(n15242) );
  OAI211_X1 U17365 ( .C1(n15244), .C2(n15243), .A(n15242), .B(n15246), .ZN(
        n17377) );
  INV_X1 U17366 ( .A(n17377), .ZN(n15245) );
  AOI21_X1 U17367 ( .B1(n15246), .B2(n15211), .A(n15245), .ZN(n15252) );
  NOR2_X1 U17368 ( .A1(n21804), .A2(n21803), .ZN(n15247) );
  OAI21_X1 U17369 ( .B1(n15252), .B2(P1_FLUSH_REG_SCAN_IN), .A(n15247), .ZN(
        n15248) );
  NAND2_X1 U17370 ( .A1(n15248), .A2(n21961), .ZN(n17384) );
  OAI21_X1 U17371 ( .B1(n22013), .B2(n22111), .A(n22059), .ZN(n16582) );
  AOI21_X1 U17372 ( .B1(n22013), .B2(n22111), .A(n16582), .ZN(n15250) );
  NAND2_X1 U17373 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n22072), .ZN(n16580) );
  INV_X1 U17374 ( .A(n16580), .ZN(n16577) );
  NOR2_X1 U17375 ( .A1(n22063), .A2(n16577), .ZN(n15249) );
  OAI21_X1 U17376 ( .B1(n15250), .B2(n15249), .A(n17384), .ZN(n15251) );
  OAI21_X1 U17377 ( .B1(n17384), .B2(n22039), .A(n15251), .ZN(P1_U3476) );
  NOR2_X1 U17378 ( .A1(n15252), .A2(n21803), .ZN(n21811) );
  OAI22_X1 U17379 ( .A1(n13134), .A2(n22115), .B1(n15253), .B2(n16577), .ZN(
        n15254) );
  OAI21_X1 U17380 ( .B1(n21811), .B2(n15254), .A(n17384), .ZN(n15255) );
  OAI21_X1 U17381 ( .B1(n17384), .B2(n22076), .A(n15255), .ZN(P1_U3478) );
  AOI22_X1 U17382 ( .A1(n22344), .A2(n11078), .B1(n15416), .B2(n22389), .ZN(
        n15256) );
  OAI21_X1 U17383 ( .B1(n11059), .B2(n21999), .A(n15256), .ZN(n15257) );
  AOI21_X1 U17384 ( .B1(n15419), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n15257), .ZN(n15258) );
  OAI21_X1 U17385 ( .B1(n15421), .B2(n15828), .A(n15258), .ZN(P1_U3096) );
  AND2_X1 U17386 ( .A1(n15260), .A2(n15259), .ZN(n15265) );
  NAND3_X1 U17387 ( .A1(n15262), .A2(n15261), .A3(n15326), .ZN(n15263) );
  INV_X1 U17388 ( .A(n15281), .ZN(n15309) );
  NAND2_X1 U17389 ( .A1(n14791), .A2(n15309), .ZN(n15278) );
  INV_X1 U17390 ( .A(n15283), .ZN(n15267) );
  NAND2_X1 U17391 ( .A1(n15267), .A2(n15291), .ZN(n15302) );
  AND2_X1 U17392 ( .A1(n15297), .A2(n15302), .ZN(n15273) );
  NAND2_X1 U17393 ( .A1(n11912), .A2(n15268), .ZN(n15298) );
  INV_X1 U17394 ( .A(n15269), .ZN(n15271) );
  NAND2_X1 U17395 ( .A1(n15291), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15270) );
  NAND2_X1 U17396 ( .A1(n15271), .A2(n15270), .ZN(n15272) );
  AOI22_X1 U17397 ( .A1(n15273), .A2(n15298), .B1(n15786), .B2(n15272), .ZN(
        n15276) );
  OR2_X1 U17398 ( .A1(n15321), .A2(n15312), .ZN(n15296) );
  INV_X1 U17399 ( .A(n15273), .ZN(n15274) );
  NAND2_X1 U17400 ( .A1(n15296), .A2(n15274), .ZN(n15275) );
  AND2_X1 U17401 ( .A1(n15276), .A2(n15275), .ZN(n15277) );
  NAND2_X1 U17402 ( .A1(n15278), .A2(n15277), .ZN(n17288) );
  AND2_X1 U17403 ( .A1(n15280), .A2(n15279), .ZN(n15284) );
  OAI22_X1 U17404 ( .A1(n18884), .A2(n15281), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15284), .ZN(n15783) );
  AOI21_X1 U17405 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15786), .A(
        n15783), .ZN(n15282) );
  NAND2_X1 U17406 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15282), .ZN(
        n15290) );
  NAND2_X1 U17407 ( .A1(n18613), .A2(n15309), .ZN(n15289) );
  NOR2_X1 U17408 ( .A1(n11261), .A2(n15283), .ZN(n15287) );
  INV_X1 U17409 ( .A(n15284), .ZN(n15286) );
  AOI22_X1 U17410 ( .A1(n15287), .A2(n15286), .B1(n15786), .B2(n15285), .ZN(
        n15288) );
  NAND2_X1 U17411 ( .A1(n15289), .A2(n15288), .ZN(n17281) );
  AOI222_X1 U17412 ( .A1(n19523), .A2(n15290), .B1(n19523), .B2(n17281), .C1(
        n15290), .C2(n17281), .ZN(n15294) );
  OR2_X1 U17413 ( .A1(n17288), .A2(n15784), .ZN(n15293) );
  NAND2_X1 U17414 ( .A1(n15784), .A2(n15291), .ZN(n15292) );
  NAND2_X1 U17415 ( .A1(n15293), .A2(n15292), .ZN(n15334) );
  OAI22_X1 U17416 ( .A1(n15294), .A2(n15784), .B1(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15334), .ZN(n15295) );
  OAI21_X1 U17417 ( .B1(n17288), .B2(n19518), .A(n15295), .ZN(n15311) );
  AND2_X1 U17418 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15299) );
  AOI22_X1 U17419 ( .A1(n15296), .A2(n15302), .B1(n15299), .B2(n15786), .ZN(
        n15305) );
  NAND2_X1 U17420 ( .A1(n15298), .A2(n15297), .ZN(n15303) );
  INV_X1 U17421 ( .A(n15299), .ZN(n15300) );
  NAND2_X1 U17422 ( .A1(n15786), .A2(n15300), .ZN(n15301) );
  AND3_X1 U17423 ( .A1(n15303), .A2(n15302), .A3(n15301), .ZN(n15304) );
  MUX2_X1 U17424 ( .A(n15305), .B(n15304), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n15307) );
  NAND2_X1 U17425 ( .A1(n15307), .A2(n15306), .ZN(n15308) );
  AOI21_X1 U17426 ( .B1(n11487), .B2(n15309), .A(n15308), .ZN(n17291) );
  MUX2_X1 U17427 ( .A(n17291), .B(n11374), .S(n15784), .Z(n15335) );
  OR2_X1 U17428 ( .A1(n15335), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n15310) );
  AOI221_X1 U17429 ( .B1(n15311), .B2(n15310), .C1(n15335), .C2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15337) );
  INV_X1 U17430 ( .A(n15312), .ZN(n15324) );
  INV_X1 U17431 ( .A(n18901), .ZN(n15314) );
  OAI22_X1 U17432 ( .A1(n15316), .A2(n15315), .B1(n15314), .B2(n15313), .ZN(
        n15318) );
  NAND2_X1 U17433 ( .A1(n15318), .A2(n15317), .ZN(n15323) );
  INV_X1 U17434 ( .A(n15319), .ZN(n15320) );
  AOI22_X1 U17435 ( .A1(n15321), .A2(n15781), .B1(n11943), .B2(n15320), .ZN(
        n15322) );
  OAI211_X1 U17436 ( .C1(n15324), .C2(n15781), .A(n15323), .B(n15322), .ZN(
        n18916) );
  INV_X1 U17437 ( .A(n18916), .ZN(n15333) );
  INV_X1 U17438 ( .A(n15325), .ZN(n15327) );
  NOR3_X1 U17439 ( .A1(n15328), .A2(n15327), .A3(n15326), .ZN(n18915) );
  OR2_X1 U17440 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(P2_MORE_REG_SCAN_IN), .ZN(
        n15331) );
  NOR3_X1 U17441 ( .A1(n18870), .A2(n18869), .A3(n11969), .ZN(n15330) );
  AOI211_X1 U17442 ( .C1(n18915), .C2(n15331), .A(n15330), .B(n15329), .ZN(
        n15332) );
  OAI211_X1 U17443 ( .C1(n15335), .C2(n15334), .A(n15333), .B(n15332), .ZN(
        n15336) );
  AOI211_X1 U17444 ( .C1(n15784), .C2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n15337), .B(n15336), .ZN(n18913) );
  NAND3_X1 U17445 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n18913), .A3(n17326), 
        .ZN(n15343) );
  INV_X1 U17446 ( .A(n15338), .ZN(n15339) );
  AND2_X1 U17447 ( .A1(n15340), .A2(n15339), .ZN(n15341) );
  AOI21_X1 U17448 ( .B1(n15343), .B2(n15342), .A(n15341), .ZN(n18905) );
  OAI21_X1 U17449 ( .B1(n18905), .B2(n11407), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n15344) );
  NOR2_X1 U17450 ( .A1(n11407), .A2(n17676), .ZN(n17329) );
  INV_X1 U17451 ( .A(n17329), .ZN(n18900) );
  NAND2_X1 U17452 ( .A1(n15344), .A2(n18900), .ZN(P2_U3593) );
  AOI22_X1 U17453 ( .A1(n22344), .A2(n11074), .B1(n15416), .B2(n22211), .ZN(
        n15345) );
  OAI21_X1 U17454 ( .B1(n11067), .B2(n21999), .A(n15345), .ZN(n15346) );
  AOI21_X1 U17455 ( .B1(n15419), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n15346), .ZN(n15347) );
  OAI21_X1 U17456 ( .B1(n15421), .B2(n15832), .A(n15347), .ZN(P1_U3092) );
  INV_X1 U17457 ( .A(n22175), .ZN(n22184) );
  AOI22_X1 U17458 ( .A1(n22344), .A2(n22181), .B1(n15416), .B2(n22179), .ZN(
        n15348) );
  OAI21_X1 U17459 ( .B1(n22184), .B2(n21999), .A(n15348), .ZN(n15349) );
  AOI21_X1 U17460 ( .B1(n15419), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A(
        n15349), .ZN(n15350) );
  OAI21_X1 U17461 ( .B1(n15421), .B2(n15852), .A(n15350), .ZN(P1_U3091) );
  NAND2_X1 U17462 ( .A1(n15351), .A2(n21631), .ZN(n15359) );
  INV_X1 U17463 ( .A(n21609), .ZN(n15386) );
  NAND2_X1 U17464 ( .A1(n21773), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n15353) );
  INV_X1 U17465 ( .A(n16136), .ZN(n15388) );
  NOR2_X1 U17466 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n21622), .ZN(n15383) );
  OAI21_X1 U17467 ( .B1(n15388), .B2(n15383), .A(P1_REIP_REG_2__SCAN_IN), .ZN(
        n15352) );
  OAI211_X1 U17468 ( .C1(P1_REIP_REG_2__SCAN_IN), .C2(n15354), .A(n15353), .B(
        n15352), .ZN(n15355) );
  AOI21_X1 U17469 ( .B1(n15466), .B2(n21724), .A(n15355), .ZN(n15356) );
  OAI21_X1 U17470 ( .B1(n22063), .B2(n15386), .A(n15356), .ZN(n15357) );
  AOI21_X1 U17471 ( .B1(n21748), .B2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n15357), .ZN(n15358) );
  OAI211_X1 U17472 ( .C1(n21702), .C2(n15360), .A(n15359), .B(n15358), .ZN(
        P1_U2838) );
  OR2_X1 U17473 ( .A1(n15362), .A2(n15361), .ZN(n15364) );
  NAND2_X1 U17474 ( .A1(n15364), .A2(n15363), .ZN(n17682) );
  NOR2_X1 U17475 ( .A1(n15366), .A2(n15365), .ZN(n15473) );
  XOR2_X1 U17476 ( .A(n17682), .B(n15473), .Z(n15472) );
  XNOR2_X1 U17477 ( .A(n15472), .B(n19502), .ZN(n15370) );
  INV_X1 U17478 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n15367) );
  OAI22_X1 U17479 ( .A1(n15427), .A2(n19751), .B1(n19374), .B2(n15367), .ZN(
        n15368) );
  AOI21_X1 U17480 ( .B1(n19585), .B2(n17682), .A(n15368), .ZN(n15369) );
  OAI21_X1 U17481 ( .B1(n15370), .B2(n16771), .A(n15369), .ZN(P2_U2917) );
  INV_X1 U17482 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n15371) );
  OAI22_X1 U17483 ( .A1(n21710), .A2(n15371), .B1(n21788), .B2(n15454), .ZN(
        n15375) );
  OAI21_X1 U17484 ( .B1(n21748), .B2(n21782), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15373) );
  AOI22_X1 U17485 ( .A1(n13136), .A2(n21609), .B1(P1_EBX_REG_0__SCAN_IN), .B2(
        n21773), .ZN(n15372) );
  OAI211_X1 U17486 ( .C1(n15393), .C2(n20144), .A(n15373), .B(n15372), .ZN(
        n15374) );
  OR2_X1 U17487 ( .A1(n15375), .A2(n15374), .ZN(P1_U2840) );
  AOI21_X1 U17488 ( .B1(n20192), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n15376), .ZN(n15378) );
  NAND2_X1 U17489 ( .A1(n20172), .A2(n21608), .ZN(n15377) );
  OAI211_X1 U17490 ( .C1(n21607), .C2(n20194), .A(n15378), .B(n15377), .ZN(
        n15379) );
  INV_X1 U17491 ( .A(n15379), .ZN(n15380) );
  OAI21_X1 U17492 ( .B1(n15381), .B2(n21789), .A(n15380), .ZN(P1_U2995) );
  AOI21_X1 U17493 ( .B1(n21773), .B2(P1_EBX_REG_1__SCAN_IN), .A(n15383), .ZN(
        n15385) );
  NAND2_X1 U17494 ( .A1(n15534), .A2(n21724), .ZN(n15384) );
  OAI211_X1 U17495 ( .C1(n11019), .C2(n15386), .A(n15385), .B(n15384), .ZN(
        n15387) );
  AOI21_X1 U17496 ( .B1(n15388), .B2(P1_REIP_REG_1__SCAN_IN), .A(n15387), .ZN(
        n15390) );
  NAND2_X1 U17497 ( .A1(n21748), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15389) );
  OAI211_X1 U17498 ( .C1(n21702), .C2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n15390), .B(n15389), .ZN(n15391) );
  INV_X1 U17499 ( .A(n15391), .ZN(n15392) );
  OAI21_X1 U17500 ( .B1(n15393), .B2(n15536), .A(n15392), .ZN(P1_U2839) );
  NAND2_X1 U17501 ( .A1(n14570), .A2(n15394), .ZN(n15395) );
  AND2_X1 U17502 ( .A1(n15485), .A2(n15395), .ZN(n18676) );
  INV_X1 U17503 ( .A(n18676), .ZN(n15400) );
  NAND2_X1 U17504 ( .A1(n15396), .A2(n15397), .ZN(n15483) );
  OAI211_X1 U17505 ( .C1(n15396), .C2(n15397), .A(n15483), .B(n16686), .ZN(
        n15399) );
  NAND2_X1 U17506 ( .A1(n16689), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n15398) );
  OAI211_X1 U17507 ( .C1(n15400), .C2(n16689), .A(n15399), .B(n15398), .ZN(
        P2_U2875) );
  NOR2_X2 U17508 ( .A1(n15412), .A2(n15401), .ZN(n22148) );
  INV_X1 U17509 ( .A(n22148), .ZN(n15848) );
  INV_X1 U17510 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20257) );
  INV_X1 U17511 ( .A(DATAI_25_), .ZN(n17502) );
  OAI22_X1 U17512 ( .A1(n20257), .A2(n15414), .B1(n17502), .B2(n15413), .ZN(
        n22144) );
  INV_X1 U17513 ( .A(DATAI_17_), .ZN(n17518) );
  INV_X1 U17514 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20241) );
  OAI22_X1 U17515 ( .A1(n17518), .A2(n15413), .B1(n20241), .B2(n15414), .ZN(
        n22149) );
  NAND2_X1 U17516 ( .A1(n15415), .A2(n15967), .ZN(n22141) );
  AOI22_X1 U17517 ( .A1(n22344), .A2(n11080), .B1(n15416), .B2(n22147), .ZN(
        n15402) );
  OAI21_X1 U17518 ( .B1(n11061), .B2(n21999), .A(n15402), .ZN(n15403) );
  AOI21_X1 U17519 ( .B1(n15419), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A(
        n15403), .ZN(n15404) );
  OAI21_X1 U17520 ( .B1(n15421), .B2(n15848), .A(n15404), .ZN(P1_U3090) );
  NOR2_X2 U17521 ( .A1(n15412), .A2(n12558), .ZN(n22306) );
  INV_X1 U17522 ( .A(n22306), .ZN(n15816) );
  INV_X1 U17523 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20268) );
  INV_X1 U17524 ( .A(DATAI_30_), .ZN(n17415) );
  OAI22_X1 U17525 ( .A1(n20268), .A2(n15414), .B1(n17415), .B2(n15413), .ZN(
        n22302) );
  INV_X1 U17526 ( .A(DATAI_22_), .ZN(n17494) );
  INV_X1 U17527 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20251) );
  OAI22_X1 U17528 ( .A1(n17494), .A2(n15413), .B1(n20251), .B2(n15414), .ZN(
        n22307) );
  NAND2_X1 U17529 ( .A1(n15415), .A2(n16281), .ZN(n22299) );
  AOI22_X1 U17530 ( .A1(n22344), .A2(n11082), .B1(n15416), .B2(n22305), .ZN(
        n15405) );
  OAI21_X1 U17531 ( .B1(n11063), .B2(n21999), .A(n15405), .ZN(n15406) );
  AOI21_X1 U17532 ( .B1(n15419), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A(
        n15406), .ZN(n15407) );
  OAI21_X1 U17533 ( .B1(n15421), .B2(n15816), .A(n15407), .ZN(P1_U3095) );
  NOR2_X2 U17534 ( .A1(n15412), .A2(n12574), .ZN(n22274) );
  INV_X1 U17535 ( .A(n22274), .ZN(n15824) );
  INV_X1 U17536 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20266) );
  INV_X1 U17537 ( .A(DATAI_29_), .ZN(n17414) );
  INV_X1 U17538 ( .A(n22270), .ZN(n22278) );
  INV_X1 U17539 ( .A(DATAI_21_), .ZN(n17512) );
  INV_X1 U17540 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20249) );
  OAI22_X1 U17541 ( .A1(n17512), .A2(n15413), .B1(n20249), .B2(n15414), .ZN(
        n22275) );
  NAND2_X1 U17542 ( .A1(n15415), .A2(n16285), .ZN(n22267) );
  AOI22_X1 U17543 ( .A1(n22344), .A2(n11076), .B1(n15416), .B2(n22273), .ZN(
        n15408) );
  OAI21_X1 U17544 ( .B1(n22278), .B2(n21999), .A(n15408), .ZN(n15409) );
  AOI21_X1 U17545 ( .B1(n15419), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A(
        n15409), .ZN(n15410) );
  OAI21_X1 U17546 ( .B1(n15421), .B2(n15824), .A(n15410), .ZN(P1_U3094) );
  NOR2_X2 U17547 ( .A1(n15412), .A2(n15411), .ZN(n22243) );
  INV_X1 U17548 ( .A(n22243), .ZN(n15820) );
  INV_X1 U17549 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20264) );
  INV_X1 U17550 ( .A(DATAI_28_), .ZN(n17499) );
  OAI22_X1 U17551 ( .A1(n20264), .A2(n15414), .B1(n17499), .B2(n15413), .ZN(
        n22239) );
  INV_X1 U17552 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n20247) );
  INV_X1 U17553 ( .A(DATAI_20_), .ZN(n17513) );
  OAI22_X1 U17554 ( .A1(n20247), .A2(n15414), .B1(n17513), .B2(n15413), .ZN(
        n22244) );
  NAND2_X1 U17555 ( .A1(n15415), .A2(n16288), .ZN(n22236) );
  AOI22_X1 U17556 ( .A1(n22344), .A2(n11084), .B1(n15416), .B2(n22242), .ZN(
        n15417) );
  OAI21_X1 U17557 ( .B1(n11065), .B2(n21999), .A(n15417), .ZN(n15418) );
  AOI21_X1 U17558 ( .B1(n15419), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A(
        n15418), .ZN(n15420) );
  OAI21_X1 U17559 ( .B1(n15421), .B2(n15820), .A(n15420), .ZN(P1_U3093) );
  NAND2_X1 U17560 ( .A1(n17144), .A2(n15424), .ZN(n15425) );
  NAND2_X1 U17561 ( .A1(n15422), .A2(n15425), .ZN(n18698) );
  OAI222_X1 U17562 ( .A1(n18698), .A2(n19367), .B1(n17739), .B2(n19374), .C1(
        n15427), .C2(n15426), .ZN(P2_U2904) );
  NAND2_X1 U17563 ( .A1(n15437), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n15430) );
  OAI22_X1 U17564 ( .A1(n22010), .A2(n11075), .B1(n22267), .B2(n15438), .ZN(
        n15428) );
  AOI21_X1 U17565 ( .B1(n22270), .B2(n15805), .A(n15428), .ZN(n15429) );
  OAI211_X1 U17566 ( .C1(n15442), .C2(n15824), .A(n15430), .B(n15429), .ZN(
        P1_U3078) );
  NAND2_X1 U17567 ( .A1(n15437), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n15433) );
  OAI22_X1 U17568 ( .A1(n22010), .A2(n11081), .B1(n22299), .B2(n15438), .ZN(
        n15431) );
  AOI21_X1 U17569 ( .B1(n11064), .B2(n15805), .A(n15431), .ZN(n15432) );
  OAI211_X1 U17570 ( .C1(n15442), .C2(n15816), .A(n15433), .B(n15432), .ZN(
        P1_U3079) );
  NAND2_X1 U17571 ( .A1(n15437), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n15436) );
  OAI22_X1 U17572 ( .A1(n22010), .A2(n11083), .B1(n22236), .B2(n15438), .ZN(
        n15434) );
  AOI21_X1 U17573 ( .B1(n11066), .B2(n15805), .A(n15434), .ZN(n15435) );
  OAI211_X1 U17574 ( .C1(n15442), .C2(n15820), .A(n15436), .B(n15435), .ZN(
        P1_U3077) );
  NAND2_X1 U17575 ( .A1(n15437), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n15441) );
  OAI22_X1 U17576 ( .A1(n22010), .A2(n11079), .B1(n22141), .B2(n15438), .ZN(
        n15439) );
  AOI21_X1 U17577 ( .B1(n11062), .B2(n15805), .A(n15439), .ZN(n15440) );
  OAI211_X1 U17578 ( .C1(n15442), .C2(n15848), .A(n15441), .B(n15440), .ZN(
        P1_U3074) );
  INV_X1 U17579 ( .A(n16281), .ZN(n15448) );
  NAND2_X1 U17580 ( .A1(n15445), .A2(n15446), .ZN(n15447) );
  NAND2_X1 U17581 ( .A1(n15444), .A2(n15447), .ZN(n21645) );
  OAI222_X1 U17582 ( .A1(n15944), .A2(n15448), .B1(n16273), .B2(n13176), .C1(
        n16280), .C2(n21645), .ZN(P1_U2898) );
  INV_X1 U17583 ( .A(n16285), .ZN(n15452) );
  OR2_X1 U17584 ( .A1(n15197), .A2(n15449), .ZN(n15450) );
  AND2_X1 U17585 ( .A1(n15445), .A2(n15450), .ZN(n21632) );
  INV_X1 U17586 ( .A(n21632), .ZN(n15451) );
  OAI222_X1 U17587 ( .A1(n15452), .A2(n15944), .B1(n16273), .B2(n13169), .C1(
        n16280), .C2(n15451), .ZN(P1_U2899) );
  INV_X1 U17588 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n15453) );
  OAI222_X1 U17589 ( .A1(n15454), .A2(n16247), .B1(n16246), .B2(n15453), .C1(
        n20144), .C2(n16237), .ZN(P1_U2872) );
  NOR2_X1 U17590 ( .A1(n15486), .A2(n15456), .ZN(n15457) );
  OR2_X1 U17591 ( .A1(n15455), .A2(n15457), .ZN(n17143) );
  AND2_X1 U17592 ( .A1(n15396), .A2(n15458), .ZN(n15462) );
  AND2_X1 U17593 ( .A1(n15396), .A2(n15459), .ZN(n15577) );
  INV_X1 U17594 ( .A(n15577), .ZN(n15460) );
  OAI211_X1 U17595 ( .C1(n15462), .C2(n15461), .A(n15460), .B(n16686), .ZN(
        n15464) );
  NAND2_X1 U17596 ( .A1(n16689), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n15463) );
  OAI211_X1 U17597 ( .C1(n17143), .C2(n16689), .A(n15464), .B(n15463), .ZN(
        P2_U2873) );
  XOR2_X1 U17598 ( .A(n15507), .B(n20134), .Z(n21637) );
  AOI22_X1 U17599 ( .A1(n13631), .A2(n21637), .B1(n15926), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n15465) );
  OAI21_X1 U17600 ( .B1(n21645), .B2(n16237), .A(n15465), .ZN(P1_U2866) );
  AOI22_X1 U17601 ( .A1(n13631), .A2(n15466), .B1(n15926), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n15467) );
  OAI21_X1 U17602 ( .B1(n15468), .B2(n16237), .A(n15467), .ZN(P1_U2870) );
  AOI21_X1 U17603 ( .B1(n15471), .B2(n15470), .A(n15469), .ZN(n17690) );
  XNOR2_X1 U17604 ( .A(n19521), .B(n17690), .ZN(n15477) );
  INV_X1 U17605 ( .A(n15472), .ZN(n15475) );
  NAND2_X1 U17606 ( .A1(n15473), .A2(n17682), .ZN(n15474) );
  OAI21_X1 U17607 ( .B1(n15475), .B2(n17692), .A(n15474), .ZN(n15476) );
  NOR2_X1 U17608 ( .A1(n15476), .A2(n15477), .ZN(n15501) );
  AOI21_X1 U17609 ( .B1(n15477), .B2(n15476), .A(n15501), .ZN(n15481) );
  AOI22_X1 U17610 ( .A1(n19585), .A2(n17690), .B1(n19579), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n15480) );
  INV_X1 U17611 ( .A(n19712), .ZN(n15478) );
  NAND2_X1 U17612 ( .A1(n19369), .A2(n15478), .ZN(n15479) );
  OAI211_X1 U17613 ( .C1(n15481), .C2(n16771), .A(n15480), .B(n15479), .ZN(
        P2_U2916) );
  XNOR2_X1 U17614 ( .A(n15483), .B(n15482), .ZN(n15489) );
  AND2_X1 U17615 ( .A1(n15485), .A2(n15484), .ZN(n15487) );
  OR2_X1 U17616 ( .A1(n15487), .A2(n15486), .ZN(n17162) );
  MUX2_X1 U17617 ( .A(n17162), .B(n11871), .S(n16689), .Z(n15488) );
  OAI21_X1 U17618 ( .B1(n15489), .B2(n16698), .A(n15488), .ZN(P2_U2874) );
  XOR2_X1 U17619 ( .A(n11006), .B(n15491), .Z(n21539) );
  NAND2_X1 U17620 ( .A1(n21539), .A2(n20188), .ZN(n15495) );
  INV_X1 U17621 ( .A(n21650), .ZN(n15493) );
  NAND2_X1 U17622 ( .A1(n21585), .A2(P1_REIP_REG_6__SCAN_IN), .ZN(n21535) );
  OAI21_X1 U17623 ( .B1(n20155), .B2(n21643), .A(n21535), .ZN(n15492) );
  AOI21_X1 U17624 ( .B1(n15493), .B2(n20172), .A(n15492), .ZN(n15494) );
  OAI211_X1 U17625 ( .C1(n20194), .C2(n21645), .A(n15495), .B(n15494), .ZN(
        P1_U2993) );
  AOI21_X1 U17626 ( .B1(n15498), .B2(n15497), .A(n15496), .ZN(n15716) );
  INV_X1 U17627 ( .A(n15716), .ZN(n15776) );
  NOR2_X1 U17628 ( .A1(n19521), .A2(n17690), .ZN(n15500) );
  XOR2_X1 U17629 ( .A(n15469), .B(n15499), .Z(n15601) );
  INV_X1 U17630 ( .A(n15601), .ZN(n15701) );
  OAI21_X1 U17631 ( .B1(n15501), .B2(n15500), .A(n15701), .ZN(n15569) );
  INV_X1 U17632 ( .A(n15611), .ZN(n15502) );
  NAND3_X1 U17633 ( .A1(n15569), .A2(n19586), .A3(n15502), .ZN(n15505) );
  INV_X1 U17634 ( .A(n19631), .ZN(n15503) );
  AOI22_X1 U17635 ( .A1(n19369), .A2(n15503), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n19579), .ZN(n15504) );
  OAI211_X1 U17636 ( .C1(n19367), .C2(n15776), .A(n15505), .B(n15504), .ZN(
        P2_U2914) );
  AOI21_X1 U17637 ( .B1(n20134), .B2(n15507), .A(n15506), .ZN(n15508) );
  OR2_X1 U17638 ( .A1(n15624), .A2(n15508), .ZN(n21652) );
  INV_X1 U17639 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n15511) );
  AND2_X1 U17640 ( .A1(n15509), .A2(n15444), .ZN(n15510) );
  OR2_X1 U17641 ( .A1(n15510), .A2(n11049), .ZN(n21657) );
  OAI222_X1 U17642 ( .A1(n21652), .A2(n16247), .B1(n15511), .B2(n20137), .C1(
        n21657), .C2(n16237), .ZN(P1_U2865) );
  OAI21_X1 U17643 ( .B1(n15514), .B2(n15513), .A(n15512), .ZN(n15530) );
  NAND2_X1 U17644 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n16976), .ZN(n15517) );
  OAI211_X1 U17645 ( .C1(n16019), .C2(n15515), .A(n15699), .B(n17262), .ZN(
        n15516) );
  OAI211_X1 U17646 ( .C1(n17227), .C2(n15699), .A(n15517), .B(n15516), .ZN(
        n15519) );
  INV_X1 U17647 ( .A(n17690), .ZN(n15683) );
  OAI22_X1 U17648 ( .A1(n15682), .A2(n18885), .B1(n17229), .B2(n15683), .ZN(
        n15518) );
  NOR2_X1 U17649 ( .A1(n15519), .A2(n15518), .ZN(n15524) );
  INV_X1 U17650 ( .A(n12203), .ZN(n15522) );
  NAND2_X1 U17651 ( .A1(n15522), .A2(n15521), .ZN(n15527) );
  NAND3_X1 U17652 ( .A1(n15520), .A2(n15527), .A3(n18879), .ZN(n15523) );
  OAI211_X1 U17653 ( .C1(n15530), .C2(n18881), .A(n15524), .B(n15523), .ZN(
        P2_U3043) );
  NOR2_X1 U17654 ( .A1(n15682), .A2(n17651), .ZN(n15526) );
  OAI22_X1 U17655 ( .A1(n15681), .A2(n17658), .B1(n17744), .B2(n18746), .ZN(
        n15525) );
  AOI211_X1 U17656 ( .C1(n17647), .C2(n15679), .A(n15526), .B(n15525), .ZN(
        n15529) );
  NAND3_X1 U17657 ( .A1(n15520), .A2(n15527), .A3(n17668), .ZN(n15528) );
  OAI211_X1 U17658 ( .C1(n15530), .C2(n17670), .A(n15529), .B(n15528), .ZN(
        P2_U3011) );
  INV_X1 U17659 ( .A(n15531), .ZN(n16275) );
  OAI222_X1 U17660 ( .A1(n15944), .A2(n16275), .B1(n16273), .B2(n13184), .C1(
        n16280), .C2(n21657), .ZN(P1_U2897) );
  XNOR2_X1 U17661 ( .A(n11049), .B(n11057), .ZN(n21665) );
  INV_X1 U17662 ( .A(n21665), .ZN(n15533) );
  MUX2_X1 U17663 ( .A(DATAI_8_), .B(BUF1_REG_8__SCAN_IN), .S(n15942), .Z(
        n21884) );
  AOI22_X1 U17664 ( .A1(n15920), .A2(n21884), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n16248), .ZN(n15532) );
  OAI21_X1 U17665 ( .B1(n15533), .B2(n16280), .A(n15532), .ZN(P1_U2896) );
  AOI22_X1 U17666 ( .A1(n13631), .A2(n15534), .B1(n15926), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n15535) );
  OAI21_X1 U17667 ( .B1(n16237), .B2(n15536), .A(n15535), .ZN(P1_U2871) );
  INV_X1 U17668 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n15538) );
  AOI22_X1 U17669 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n20034), .B1(n20031), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n15537) );
  OAI21_X1 U17670 ( .B1(n15538), .B2(n15555), .A(n15537), .ZN(P1_U2920) );
  AOI22_X1 U17671 ( .A1(n20031), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n15539) );
  OAI21_X1 U17672 ( .B1(n16272), .B2(n15555), .A(n15539), .ZN(P1_U2913) );
  INV_X1 U17673 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n15541) );
  AOI22_X1 U17674 ( .A1(n21515), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n15540) );
  OAI21_X1 U17675 ( .B1(n15541), .B2(n15555), .A(n15540), .ZN(P1_U2914) );
  INV_X1 U17676 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n15543) );
  AOI22_X1 U17677 ( .A1(n21515), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n15542) );
  OAI21_X1 U17678 ( .B1(n15543), .B2(n15555), .A(n15542), .ZN(P1_U2916) );
  INV_X1 U17679 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n21896) );
  AOI22_X1 U17680 ( .A1(n21515), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n15544) );
  OAI21_X1 U17681 ( .B1(n21896), .B2(n15555), .A(n15544), .ZN(P1_U2911) );
  INV_X1 U17682 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n21888) );
  AOI22_X1 U17683 ( .A1(n21515), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n15545) );
  OAI21_X1 U17684 ( .B1(n21888), .B2(n15555), .A(n15545), .ZN(P1_U2912) );
  INV_X1 U17685 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n15547) );
  AOI22_X1 U17686 ( .A1(n21515), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n15546) );
  OAI21_X1 U17687 ( .B1(n15547), .B2(n15555), .A(n15546), .ZN(P1_U2915) );
  INV_X1 U17688 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n15549) );
  AOI22_X1 U17689 ( .A1(n21515), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n15548) );
  OAI21_X1 U17690 ( .B1(n15549), .B2(n15555), .A(n15548), .ZN(P1_U2917) );
  INV_X1 U17691 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n21906) );
  AOI22_X1 U17692 ( .A1(n21515), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n15550) );
  OAI21_X1 U17693 ( .B1(n21906), .B2(n15555), .A(n15550), .ZN(P1_U2910) );
  INV_X1 U17694 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n21916) );
  AOI22_X1 U17695 ( .A1(n21515), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n15551) );
  OAI21_X1 U17696 ( .B1(n21916), .B2(n15555), .A(n15551), .ZN(P1_U2909) );
  INV_X1 U17697 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n21936) );
  AOI22_X1 U17698 ( .A1(n21515), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n15552) );
  OAI21_X1 U17699 ( .B1(n21936), .B2(n15555), .A(n15552), .ZN(P1_U2907) );
  INV_X1 U17700 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n21926) );
  AOI22_X1 U17701 ( .A1(n21515), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n15553) );
  OAI21_X1 U17702 ( .B1(n21926), .B2(n15555), .A(n15553), .ZN(P1_U2908) );
  INV_X1 U17703 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n21947) );
  AOI22_X1 U17704 ( .A1(n21515), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n15554) );
  OAI21_X1 U17705 ( .B1(n21947), .B2(n15555), .A(n15554), .ZN(P1_U2906) );
  XOR2_X1 U17706 ( .A(n15557), .B(n10987), .Z(n20151) );
  INV_X1 U17707 ( .A(n20151), .ZN(n15564) );
  AOI211_X1 U17708 ( .C1(n15618), .C2(n21529), .A(n15616), .B(n21542), .ZN(
        n15558) );
  AOI21_X1 U17709 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15558), .A(
        n16451), .ZN(n15589) );
  INV_X1 U17710 ( .A(n21542), .ZN(n15559) );
  AOI22_X1 U17711 ( .A1(n21533), .A2(n15560), .B1(n21544), .B2(n15559), .ZN(
        n21537) );
  NOR3_X1 U17712 ( .A1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n21537), .A3(
        n21541), .ZN(n15590) );
  INV_X1 U17713 ( .A(n15590), .ZN(n15561) );
  NAND2_X1 U17714 ( .A1(n21585), .A2(P1_REIP_REG_7__SCAN_IN), .ZN(n20152) );
  OAI211_X1 U17715 ( .C1(n21560), .C2(n21652), .A(n15561), .B(n20152), .ZN(
        n15562) );
  AOI21_X1 U17716 ( .B1(n15589), .B2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n15562), .ZN(n15563) );
  OAI21_X1 U17717 ( .B1(n15564), .B2(n16575), .A(n15563), .ZN(P1_U3024) );
  OAI21_X1 U17718 ( .B1(n15565), .B2(n15568), .A(n15567), .ZN(n15653) );
  INV_X1 U17719 ( .A(DATAI_9_), .ZN(n17408) );
  MUX2_X1 U17720 ( .A(n17408), .B(n20227), .S(n15942), .Z(n21892) );
  INV_X1 U17721 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n21899) );
  OAI222_X1 U17722 ( .A1(n15653), .A2(n16280), .B1(n15944), .B2(n21892), .C1(
        n21899), .C2(n16273), .ZN(P1_U2895) );
  XOR2_X1 U17723 ( .A(n15611), .B(n15569), .Z(n15573) );
  INV_X1 U17724 ( .A(n19672), .ZN(n15570) );
  AOI22_X1 U17725 ( .A1(n19369), .A2(n15570), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19579), .ZN(n15572) );
  NAND2_X1 U17726 ( .A1(n15601), .A2(n19585), .ZN(n15571) );
  OAI211_X1 U17727 ( .C1(n15573), .C2(n16771), .A(n15572), .B(n15571), .ZN(
        P2_U2915) );
  INV_X1 U17728 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n15574) );
  OAI222_X1 U17729 ( .A1(n15575), .A2(n16247), .B1(n16246), .B2(n15574), .C1(
        n16237), .C2(n21607), .ZN(P1_U2868) );
  XNOR2_X1 U17730 ( .A(n15577), .B(n15576), .ZN(n15582) );
  OR2_X1 U17731 ( .A1(n15455), .A2(n15579), .ZN(n15580) );
  NAND2_X1 U17732 ( .A1(n15578), .A2(n15580), .ZN(n18699) );
  MUX2_X1 U17733 ( .A(n18699), .B(n11878), .S(n16689), .Z(n15581) );
  OAI21_X1 U17734 ( .B1(n15582), .B2(n16698), .A(n15581), .ZN(P2_U2872) );
  XOR2_X1 U17735 ( .A(n10980), .B(n15584), .Z(n15596) );
  AOI22_X1 U17736 ( .A1(n20192), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n16504), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n15585) );
  OAI21_X1 U17737 ( .B1(n20200), .B2(n21663), .A(n15585), .ZN(n15586) );
  AOI21_X1 U17738 ( .B1(n21665), .B2(n20186), .A(n15586), .ZN(n15587) );
  OAI21_X1 U17739 ( .B1(n15596), .B2(n21789), .A(n15587), .ZN(P1_U2991) );
  INV_X1 U17740 ( .A(n15623), .ZN(n15588) );
  XNOR2_X1 U17741 ( .A(n15624), .B(n15588), .ZN(n21662) );
  INV_X1 U17742 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n21667) );
  OAI21_X1 U17743 ( .B1(n15590), .B2(n15589), .A(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15593) );
  OR4_X1 U17744 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21537), .A3(
        n15591), .A4(n21541), .ZN(n15592) );
  OAI211_X1 U17745 ( .C1(n21600), .C2(n21667), .A(n15593), .B(n15592), .ZN(
        n15594) );
  AOI21_X1 U17746 ( .B1(n21595), .B2(n21662), .A(n15594), .ZN(n15595) );
  OAI21_X1 U17747 ( .B1(n15596), .B2(n16575), .A(n15595), .ZN(P1_U3023) );
  INV_X1 U17748 ( .A(n18614), .ZN(n15733) );
  INV_X1 U17749 ( .A(n17614), .ZN(n15600) );
  NOR2_X1 U17750 ( .A1(n18717), .A2(n15597), .ZN(n15599) );
  AOI21_X1 U17751 ( .B1(n15600), .B2(n15599), .A(n18897), .ZN(n15598) );
  OAI21_X1 U17752 ( .B1(n15600), .B2(n15599), .A(n15598), .ZN(n15610) );
  INV_X1 U17753 ( .A(n17621), .ZN(n15608) );
  INV_X1 U17754 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n15603) );
  AOI22_X1 U17755 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n18852), .B1(n18763), .B2(
        n15601), .ZN(n15602) );
  OAI211_X1 U17756 ( .C1(n15603), .C2(n18621), .A(n16970), .B(n15602), .ZN(
        n15604) );
  AOI21_X1 U17757 ( .B1(n18850), .B2(P2_REIP_REG_4__SCAN_IN), .A(n15604), .ZN(
        n15605) );
  OAI21_X1 U17758 ( .B1(n18803), .B2(n15606), .A(n15605), .ZN(n15607) );
  AOI21_X1 U17759 ( .B1(n15608), .B2(n18811), .A(n15607), .ZN(n15609) );
  OAI211_X1 U17760 ( .C1(n15611), .C2(n15733), .A(n15610), .B(n15609), .ZN(
        P2_U2851) );
  NAND2_X1 U17761 ( .A1(n15614), .A2(n15613), .ZN(n15615) );
  NAND2_X1 U17762 ( .A1(n16557), .A2(n15615), .ZN(n15659) );
  AOI21_X1 U17763 ( .B1(n15618), .B2(n15617), .A(n15616), .ZN(n15619) );
  OAI21_X1 U17764 ( .B1(n15620), .B2(n16453), .A(n15619), .ZN(n16572) );
  NOR2_X1 U17765 ( .A1(n21537), .A2(n15621), .ZN(n16571) );
  AOI22_X1 U17766 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16572), .B1(
        n16571), .B2(n16569), .ZN(n15628) );
  INV_X1 U17767 ( .A(n15794), .ZN(n15626) );
  AOI21_X1 U17768 ( .B1(n15624), .B2(n15623), .A(n15622), .ZN(n15625) );
  NOR2_X1 U17769 ( .A1(n15626), .A2(n15625), .ZN(n21673) );
  AND2_X1 U17770 ( .A1(n21585), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n15654) );
  AOI21_X1 U17771 ( .B1(n21595), .B2(n21673), .A(n15654), .ZN(n15627) );
  OAI211_X1 U17772 ( .C1(n15659), .C2(n16575), .A(n15628), .B(n15627), .ZN(
        P1_U3022) );
  AND2_X1 U17773 ( .A1(n15396), .A2(n15629), .ZN(n15632) );
  NAND2_X1 U17774 ( .A1(n15396), .A2(n15630), .ZN(n15709) );
  OAI21_X1 U17775 ( .B1(n15632), .B2(n15631), .A(n15709), .ZN(n15742) );
  INV_X1 U17776 ( .A(n15706), .ZN(n15633) );
  AOI21_X1 U17777 ( .B1(n15634), .B2(n15578), .A(n15633), .ZN(n18711) );
  NOR2_X1 U17778 ( .A1(n16651), .A2(n11881), .ZN(n15635) );
  AOI21_X1 U17779 ( .B1(n18711), .B2(n16651), .A(n15635), .ZN(n15636) );
  OAI21_X1 U17780 ( .B1(n15742), .B2(n16698), .A(n15636), .ZN(P2_U2871) );
  AND2_X1 U17781 ( .A1(n15396), .A2(n15637), .ZN(n15708) );
  OAI21_X1 U17782 ( .B1(n15708), .B2(n15639), .A(n15638), .ZN(n15802) );
  OR2_X1 U17783 ( .A1(n15640), .A2(n15641), .ZN(n15643) );
  NAND2_X1 U17784 ( .A1(n15643), .A2(n15642), .ZN(n18744) );
  AND2_X1 U17785 ( .A1(n19374), .A2(n15644), .ZN(n19581) );
  INV_X1 U17786 ( .A(n19751), .ZN(n15645) );
  AOI22_X1 U17787 ( .A1(n19581), .A2(n15645), .B1(n19579), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n15650) );
  OR2_X1 U17788 ( .A1(n15646), .A2(n19592), .ZN(n15648) );
  NOR2_X2 U17789 ( .A1(n15648), .A2(n15647), .ZN(n19582) );
  AOI22_X1 U17790 ( .A1(n19583), .A2(BUF2_REG_18__SCAN_IN), .B1(n19582), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n15649) );
  OAI211_X1 U17791 ( .C1(n18744), .C2(n16765), .A(n15650), .B(n15649), .ZN(
        n15651) );
  INV_X1 U17792 ( .A(n15651), .ZN(n15652) );
  OAI21_X1 U17793 ( .B1(n15802), .B2(n16771), .A(n15652), .ZN(P2_U2901) );
  INV_X1 U17794 ( .A(n15653), .ZN(n21679) );
  INV_X1 U17795 ( .A(n21674), .ZN(n15656) );
  AOI21_X1 U17796 ( .B1(n20192), .B2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n15654), .ZN(n15655) );
  OAI21_X1 U17797 ( .B1(n20200), .B2(n15656), .A(n15655), .ZN(n15657) );
  AOI21_X1 U17798 ( .B1(n21679), .B2(n20186), .A(n15657), .ZN(n15658) );
  OAI21_X1 U17799 ( .B1(n15659), .B2(n21789), .A(n15658), .ZN(P1_U2990) );
  XOR2_X1 U17800 ( .A(n15660), .B(n15567), .Z(n21689) );
  INV_X1 U17801 ( .A(n21689), .ZN(n15664) );
  MUX2_X1 U17802 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n15942), .Z(
        n21903) );
  AOI22_X1 U17803 ( .A1(n15920), .A2(n21903), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n16248), .ZN(n15661) );
  OAI21_X1 U17804 ( .B1(n15664), .B2(n16280), .A(n15661), .ZN(P1_U2894) );
  XNOR2_X1 U17805 ( .A(n15794), .B(n15662), .ZN(n21685) );
  AOI22_X1 U17806 ( .A1(n13631), .A2(n21685), .B1(n15926), .B2(
        P1_EBX_REG_10__SCAN_IN), .ZN(n15663) );
  OAI21_X1 U17807 ( .B1(n15664), .B2(n16237), .A(n15663), .ZN(P1_U2862) );
  NAND2_X1 U17808 ( .A1(n18752), .A2(n15665), .ZN(n15666) );
  XNOR2_X1 U17809 ( .A(n16949), .B(n15666), .ZN(n15675) );
  INV_X1 U17810 ( .A(n17161), .ZN(n15670) );
  NAND2_X1 U17811 ( .A1(n18850), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n15668) );
  AOI22_X1 U17812 ( .A1(P2_EBX_REG_13__SCAN_IN), .A2(n18852), .B1(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n18851), .ZN(n15667) );
  NAND3_X1 U17813 ( .A1(n15668), .A2(n15667), .A3(n18746), .ZN(n15669) );
  AOI21_X1 U17814 ( .B1(n15670), .B2(n18763), .A(n15669), .ZN(n15673) );
  NAND2_X1 U17815 ( .A1(n15671), .A2(n18853), .ZN(n15672) );
  OAI211_X1 U17816 ( .C1(n17162), .C2(n18857), .A(n15673), .B(n15672), .ZN(
        n15674) );
  AOI21_X1 U17817 ( .B1(n15675), .B2(n18861), .A(n15674), .ZN(n15676) );
  INV_X1 U17818 ( .A(n15676), .ZN(P2_U2842) );
  NAND2_X1 U17819 ( .A1(n18752), .A2(n15677), .ZN(n15678) );
  XNOR2_X1 U17820 ( .A(n15679), .B(n15678), .ZN(n15680) );
  NAND2_X1 U17821 ( .A1(n15680), .A2(n18861), .ZN(n15691) );
  OAI22_X1 U17822 ( .A1(n15681), .A2(n18621), .B1(n17744), .B2(n18748), .ZN(
        n15689) );
  NOR2_X1 U17823 ( .A1(n15682), .A2(n18857), .ZN(n15688) );
  OAI22_X1 U17824 ( .A1(n18733), .A2(n15684), .B1(n18855), .B2(n15683), .ZN(
        n15687) );
  NOR2_X1 U17825 ( .A1(n18803), .A2(n15685), .ZN(n15686) );
  NOR4_X1 U17826 ( .A1(n15689), .A2(n15688), .A3(n15687), .A4(n15686), .ZN(
        n15690) );
  OAI211_X1 U17827 ( .C1(n19426), .C2(n15733), .A(n15691), .B(n15690), .ZN(
        P2_U2852) );
  XNOR2_X1 U17828 ( .A(n15692), .B(n15770), .ZN(n17616) );
  INV_X1 U17829 ( .A(n17616), .ZN(n15705) );
  NAND2_X1 U17830 ( .A1(n15512), .A2(n15693), .ZN(n15695) );
  OR2_X1 U17831 ( .A1(n15695), .A2(n15694), .ZN(n15697) );
  NAND2_X1 U17832 ( .A1(n15695), .A2(n15694), .ZN(n15696) );
  AND2_X1 U17833 ( .A1(n15697), .A2(n15696), .ZN(n17618) );
  OR2_X1 U17834 ( .A1(n15699), .A2(n15698), .ZN(n15769) );
  AOI21_X1 U17835 ( .B1(n15699), .B2(n17262), .A(n17261), .ZN(n15772) );
  NAND2_X1 U17836 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n12161), .ZN(n15700) );
  OAI221_X1 U17837 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n15769), .C1(
        n15770), .C2(n15772), .A(n15700), .ZN(n15703) );
  OAI22_X1 U17838 ( .A1(n15701), .A2(n17229), .B1(n17621), .B2(n18885), .ZN(
        n15702) );
  AOI211_X1 U17839 ( .C1(n17618), .C2(n12326), .A(n15703), .B(n15702), .ZN(
        n15704) );
  OAI21_X1 U17840 ( .B1(n15705), .B2(n17277), .A(n15704), .ZN(P2_U3042) );
  XOR2_X1 U17841 ( .A(n15707), .B(n15706), .Z(n18728) );
  INV_X1 U17842 ( .A(n18728), .ZN(n15713) );
  AOI21_X1 U17843 ( .B1(n15710), .B2(n15709), .A(n15708), .ZN(n15746) );
  NAND2_X1 U17844 ( .A1(n15746), .A2(n16686), .ZN(n15712) );
  NAND2_X1 U17845 ( .A1(n16689), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n15711) );
  OAI211_X1 U17846 ( .C1(n15713), .C2(n16689), .A(n15712), .B(n15711), .ZN(
        P2_U2870) );
  NAND2_X1 U17847 ( .A1(n18752), .A2(n15714), .ZN(n15715) );
  XNOR2_X1 U17848 ( .A(n17624), .B(n15715), .ZN(n15717) );
  AOI22_X1 U17849 ( .A1(n18861), .A2(n15717), .B1(n18763), .B2(n15716), .ZN(
        n15721) );
  INV_X1 U17850 ( .A(n17630), .ZN(n15774) );
  INV_X1 U17851 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n17746) );
  AOI22_X1 U17852 ( .A1(P2_EBX_REG_5__SCAN_IN), .A2(n18852), .B1(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n18851), .ZN(n15718) );
  OAI211_X1 U17853 ( .C1(n18748), .C2(n17746), .A(n15718), .B(n16970), .ZN(
        n15719) );
  AOI21_X1 U17854 ( .B1(n15774), .B2(n18811), .A(n15719), .ZN(n15720) );
  OAI211_X1 U17855 ( .C1(n15722), .C2(n18803), .A(n15721), .B(n15720), .ZN(
        P2_U2850) );
  INV_X1 U17856 ( .A(n17610), .ZN(n15725) );
  NOR2_X1 U17857 ( .A1(n18717), .A2(n17278), .ZN(n15724) );
  INV_X1 U17858 ( .A(n15724), .ZN(n15723) );
  AOI221_X1 U17859 ( .B1(n15725), .B2(n15724), .C1(n17610), .C2(n15723), .A(
        n18897), .ZN(n15726) );
  INV_X1 U17860 ( .A(n15726), .ZN(n15732) );
  AOI22_X1 U17861 ( .A1(P2_EBX_REG_2__SCAN_IN), .A2(n18852), .B1(n18763), .B2(
        n17682), .ZN(n15728) );
  AOI22_X1 U17862 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n18851), .B1(
        P2_REIP_REG_2__SCAN_IN), .B2(n18850), .ZN(n15727) );
  OAI211_X1 U17863 ( .C1(n18803), .C2(n15729), .A(n15728), .B(n15727), .ZN(
        n15730) );
  AOI21_X1 U17864 ( .B1(n14791), .B2(n18811), .A(n15730), .ZN(n15731) );
  OAI211_X1 U17865 ( .C1(n15733), .C2(n17692), .A(n15732), .B(n15731), .ZN(
        P2_U2853) );
  AND2_X1 U17866 ( .A1(n15422), .A2(n15734), .ZN(n15737) );
  OR2_X1 U17867 ( .A1(n15737), .A2(n15736), .ZN(n18715) );
  OAI22_X1 U17868 ( .A1(n18715), .A2(n16765), .B1(n19374), .B2(n15738), .ZN(
        n15739) );
  INV_X1 U17869 ( .A(n15739), .ZN(n15741) );
  NAND2_X1 U17870 ( .A1(n19582), .A2(BUF1_REG_16__SCAN_IN), .ZN(n15740) );
  OAI211_X1 U17871 ( .C1(n19838), .C2(n16766), .A(n15741), .B(n15740), .ZN(
        n15744) );
  NOR2_X1 U17872 ( .A1(n15742), .A2(n16771), .ZN(n15743) );
  AOI211_X1 U17873 ( .C1(n19583), .C2(BUF2_REG_16__SCAN_IN), .A(n15744), .B(
        n15743), .ZN(n15745) );
  INV_X1 U17874 ( .A(n15745), .ZN(P2_U2903) );
  INV_X1 U17875 ( .A(n19583), .ZN(n16755) );
  INV_X1 U17876 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n15754) );
  NAND2_X1 U17877 ( .A1(n15746), .A2(n19586), .ZN(n15753) );
  OAI22_X1 U17878 ( .A1(n16766), .A2(n19792), .B1(n19374), .B2(n15747), .ZN(
        n15751) );
  INV_X1 U17879 ( .A(n15640), .ZN(n15748) );
  OAI21_X1 U17880 ( .B1(n15736), .B2(n15749), .A(n15748), .ZN(n18726) );
  NOR2_X1 U17881 ( .A1(n18726), .A2(n16765), .ZN(n15750) );
  AOI211_X1 U17882 ( .C1(BUF1_REG_17__SCAN_IN), .C2(n19582), .A(n15751), .B(
        n15750), .ZN(n15752) );
  OAI211_X1 U17883 ( .C1(n16755), .C2(n15754), .A(n15753), .B(n15752), .ZN(
        P2_U2902) );
  OR2_X1 U17884 ( .A1(n14768), .A2(n15755), .ZN(n15756) );
  AND2_X1 U17885 ( .A1(n15756), .A2(n14794), .ZN(n19370) );
  NAND2_X1 U17886 ( .A1(n18752), .A2(n15757), .ZN(n15758) );
  XNOR2_X1 U17887 ( .A(n17646), .B(n15758), .ZN(n15759) );
  AOI22_X1 U17888 ( .A1(n19370), .A2(n18763), .B1(n18861), .B2(n15759), .ZN(
        n15764) );
  AOI22_X1 U17889 ( .A1(P2_EBX_REG_9__SCAN_IN), .A2(n18852), .B1(n18853), .B2(
        n15760), .ZN(n15761) );
  OAI21_X1 U17890 ( .B1(n17659), .B2(n18621), .A(n15761), .ZN(n15762) );
  AOI211_X1 U17891 ( .C1(n18850), .C2(P2_REIP_REG_9__SCAN_IN), .A(n16976), .B(
        n15762), .ZN(n15763) );
  OAI211_X1 U17892 ( .C1(n17650), .C2(n18857), .A(n15764), .B(n15763), .ZN(
        P2_U2846) );
  OAI21_X1 U17893 ( .B1(n15765), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n11710), .ZN(n17626) );
  OAI21_X1 U17894 ( .B1(n15766), .B2(n15768), .A(n15767), .ZN(n17625) );
  INV_X1 U17895 ( .A(n17625), .ZN(n15779) );
  AOI221_X1 U17896 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C1(n15770), .C2(n15771), .A(
        n15769), .ZN(n15778) );
  OAI22_X1 U17897 ( .A1(n18746), .A2(n17746), .B1(n15772), .B2(n15771), .ZN(
        n15773) );
  AOI21_X1 U17898 ( .B1(n17204), .B2(n15774), .A(n15773), .ZN(n15775) );
  OAI21_X1 U17899 ( .B1(n15776), .B2(n17229), .A(n15775), .ZN(n15777) );
  AOI211_X1 U17900 ( .C1(n15779), .C2(n12326), .A(n15778), .B(n15777), .ZN(
        n15780) );
  OAI21_X1 U17901 ( .B1(n17277), .B2(n17626), .A(n15780), .ZN(P2_U3041) );
  NAND2_X1 U17902 ( .A1(n17326), .A2(n19459), .ZN(n18892) );
  INV_X1 U17903 ( .A(n18892), .ZN(n17287) );
  AOI22_X1 U17904 ( .A1(n18717), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n18595), .B2(n18752), .ZN(n17280) );
  AOI222_X1 U17905 ( .A1(n15783), .A2(n17287), .B1(n15782), .B2(n18906), .C1(
        P2_STATE2_REG_1__SCAN_IN), .C2(n17280), .ZN(n15788) );
  OAI22_X1 U17906 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19459), .B1(n15784), 
        .B2(n18914), .ZN(n15785) );
  AOI21_X1 U17907 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n17329), .A(n15785), .ZN(
        n18868) );
  AOI21_X1 U17908 ( .B1(n17287), .B2(n15786), .A(n18868), .ZN(n15787) );
  OAI22_X1 U17909 ( .A1(n15788), .A2(n18868), .B1(n15787), .B2(n11418), .ZN(
        P2_U3601) );
  INV_X1 U17910 ( .A(n15901), .ZN(n15790) );
  XNOR2_X1 U17911 ( .A(n15789), .B(n15790), .ZN(n15904) );
  INV_X1 U17912 ( .A(n15791), .ZN(n15903) );
  XNOR2_X1 U17913 ( .A(n15904), .B(n15903), .ZN(n21698) );
  OAI21_X1 U17914 ( .B1(n15794), .B2(n15793), .A(n15792), .ZN(n15795) );
  AND2_X1 U17915 ( .A1(n15795), .A2(n15925), .ZN(n21693) );
  AOI22_X1 U17916 ( .A1(n13631), .A2(n21693), .B1(n15926), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n15796) );
  OAI21_X1 U17917 ( .B1(n21698), .B2(n16237), .A(n15796), .ZN(P1_U2861) );
  OR2_X1 U17918 ( .A1(n15799), .A2(n15798), .ZN(n15800) );
  NAND2_X1 U17919 ( .A1(n15797), .A2(n15800), .ZN(n18739) );
  MUX2_X1 U17920 ( .A(n18739), .B(n11889), .S(n16689), .Z(n15801) );
  OAI21_X1 U17921 ( .B1(n15802), .B2(n16698), .A(n15801), .ZN(P2_U2869) );
  NOR2_X1 U17922 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15803), .ZN(
        n15812) );
  INV_X1 U17923 ( .A(n15812), .ZN(n15859) );
  NOR2_X2 U17924 ( .A1(n21988), .A2(n22054), .ZN(n22329) );
  INV_X1 U17925 ( .A(n21978), .ZN(n22036) );
  OR2_X1 U17926 ( .A1(n22016), .A2(n22036), .ZN(n21960) );
  NOR2_X1 U17927 ( .A1(n15809), .A2(n22106), .ZN(n22064) );
  INV_X1 U17928 ( .A(n22064), .ZN(n22088) );
  NAND3_X1 U17929 ( .A1(n15806), .A2(n22117), .A3(n11019), .ZN(n15804) );
  OAI21_X1 U17930 ( .B1(n21960), .B2(n22088), .A(n15804), .ZN(n15854) );
  OAI21_X1 U17931 ( .B1(n15805), .B2(n22329), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15808) );
  NAND2_X1 U17932 ( .A1(n15806), .A2(n11019), .ZN(n15807) );
  AOI21_X1 U17933 ( .B1(n15808), .B2(n15807), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n15811) );
  INV_X1 U17934 ( .A(n15809), .ZN(n15810) );
  NOR2_X1 U17935 ( .A1(n15810), .A2(n22106), .ZN(n22037) );
  AOI22_X1 U17936 ( .A1(n15854), .A2(n22305), .B1(
        P1_INSTQUEUE_REG_4__6__SCAN_IN), .B2(n15853), .ZN(n15813) );
  OAI21_X1 U17937 ( .B1(n15856), .B2(n11081), .A(n15813), .ZN(n15814) );
  AOI21_X1 U17938 ( .B1(n11064), .B2(n22329), .A(n15814), .ZN(n15815) );
  OAI21_X1 U17939 ( .B1(n15816), .B2(n15859), .A(n15815), .ZN(P1_U3071) );
  AOI22_X1 U17940 ( .A1(n15854), .A2(n22242), .B1(
        P1_INSTQUEUE_REG_4__4__SCAN_IN), .B2(n15853), .ZN(n15817) );
  OAI21_X1 U17941 ( .B1(n15856), .B2(n11083), .A(n15817), .ZN(n15818) );
  AOI21_X1 U17942 ( .B1(n11066), .B2(n22329), .A(n15818), .ZN(n15819) );
  OAI21_X1 U17943 ( .B1(n15820), .B2(n15859), .A(n15819), .ZN(P1_U3069) );
  AOI22_X1 U17944 ( .A1(n15854), .A2(n22273), .B1(
        P1_INSTQUEUE_REG_4__5__SCAN_IN), .B2(n15853), .ZN(n15821) );
  OAI21_X1 U17945 ( .B1(n15856), .B2(n11075), .A(n15821), .ZN(n15822) );
  AOI21_X1 U17946 ( .B1(n22270), .B2(n22329), .A(n15822), .ZN(n15823) );
  OAI21_X1 U17947 ( .B1(n15824), .B2(n15859), .A(n15823), .ZN(P1_U3070) );
  AOI22_X1 U17948 ( .A1(n15854), .A2(n22389), .B1(
        P1_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n15853), .ZN(n15825) );
  OAI21_X1 U17949 ( .B1(n15856), .B2(n11077), .A(n15825), .ZN(n15826) );
  AOI21_X1 U17950 ( .B1(n11060), .B2(n22329), .A(n15826), .ZN(n15827) );
  OAI21_X1 U17951 ( .B1(n15828), .B2(n15859), .A(n15827), .ZN(P1_U3072) );
  AOI22_X1 U17952 ( .A1(n15854), .A2(n22211), .B1(
        P1_INSTQUEUE_REG_4__3__SCAN_IN), .B2(n15853), .ZN(n15829) );
  OAI21_X1 U17953 ( .B1(n15856), .B2(n11073), .A(n15829), .ZN(n15830) );
  AOI21_X1 U17954 ( .B1(n11068), .B2(n22329), .A(n15830), .ZN(n15831) );
  OAI21_X1 U17955 ( .B1(n15832), .B2(n15859), .A(n15831), .ZN(P1_U3068) );
  INV_X1 U17956 ( .A(DATAI_11_), .ZN(n17526) );
  MUX2_X1 U17957 ( .A(n17526), .B(n20230), .S(n15942), .Z(n21912) );
  OAI222_X1 U17958 ( .A1(n16273), .A2(n21919), .B1(n15944), .B2(n21912), .C1(
        n16280), .C2(n21698), .ZN(P1_U2893) );
  OR2_X1 U17959 ( .A1(n15789), .A2(n15833), .ZN(n15906) );
  AOI21_X1 U17960 ( .B1(n15835), .B2(n15906), .A(n15834), .ZN(n15898) );
  INV_X1 U17961 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20063) );
  NAND3_X1 U17962 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .A3(n21707), .ZN(n21712) );
  NAND2_X1 U17963 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n15915), .ZN(n21717) );
  OAI211_X1 U17964 ( .C1(n15915), .C2(P1_REIP_REG_14__SCAN_IN), .A(n21717), 
        .B(n21738), .ZN(n15842) );
  INV_X1 U17965 ( .A(n15836), .ZN(n16515) );
  XNOR2_X1 U17966 ( .A(n16514), .B(n16515), .ZN(n21518) );
  NAND2_X1 U17967 ( .A1(n21518), .A2(n21724), .ZN(n15838) );
  NAND2_X1 U17968 ( .A1(n15837), .A2(n16136), .ZN(n21729) );
  OAI211_X1 U17969 ( .C1(n15839), .C2(n21761), .A(n15838), .B(n21729), .ZN(
        n15840) );
  AOI21_X1 U17970 ( .B1(n21748), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n15840), .ZN(n15841) );
  OAI211_X1 U17971 ( .C1(n21702), .C2(n15896), .A(n15842), .B(n15841), .ZN(
        n15843) );
  AOI21_X1 U17972 ( .B1(n15898), .B2(n21754), .A(n15843), .ZN(n15844) );
  INV_X1 U17973 ( .A(n15844), .ZN(P1_U2826) );
  AOI22_X1 U17974 ( .A1(n15854), .A2(n22147), .B1(
        P1_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n15853), .ZN(n15845) );
  OAI21_X1 U17975 ( .B1(n15856), .B2(n11079), .A(n15845), .ZN(n15846) );
  AOI21_X1 U17976 ( .B1(n11062), .B2(n22329), .A(n15846), .ZN(n15847) );
  OAI21_X1 U17977 ( .B1(n15848), .B2(n15859), .A(n15847), .ZN(P1_U3066) );
  AOI22_X1 U17978 ( .A1(n15854), .A2(n22179), .B1(
        P1_INSTQUEUE_REG_4__2__SCAN_IN), .B2(n15853), .ZN(n15849) );
  OAI21_X1 U17979 ( .B1(n15856), .B2(n22178), .A(n15849), .ZN(n15850) );
  AOI21_X1 U17980 ( .B1(n22175), .B2(n22329), .A(n15850), .ZN(n15851) );
  OAI21_X1 U17981 ( .B1(n15852), .B2(n15859), .A(n15851), .ZN(P1_U3067) );
  AOI22_X1 U17982 ( .A1(n15854), .A2(n22108), .B1(
        P1_INSTQUEUE_REG_4__0__SCAN_IN), .B2(n15853), .ZN(n15855) );
  OAI21_X1 U17983 ( .B1(n15856), .B2(n11071), .A(n15855), .ZN(n15857) );
  AOI21_X1 U17984 ( .B1(n11070), .B2(n22329), .A(n15857), .ZN(n15858) );
  OAI21_X1 U17985 ( .B1(n15860), .B2(n15859), .A(n15858), .ZN(P1_U3065) );
  NOR2_X1 U17986 ( .A1(n15862), .A2(n15863), .ZN(n15864) );
  OR2_X1 U17987 ( .A1(n15861), .A2(n15864), .ZN(n21735) );
  NOR2_X1 U17988 ( .A1(n15869), .A2(n15865), .ZN(n15866) );
  NAND2_X1 U17989 ( .A1(n16273), .A2(n15866), .ZN(n16265) );
  AOI22_X1 U17990 ( .A1(n16295), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n16248), .ZN(n15873) );
  NOR3_X1 U17991 ( .A1(n16248), .A2(n15867), .A3(n12562), .ZN(n15868) );
  NOR3_X1 U17992 ( .A1(n16248), .A2(n15942), .A3(n15869), .ZN(n15870) );
  AOI22_X1 U17993 ( .A1(n16298), .A2(n15871), .B1(n16296), .B2(DATAI_16_), 
        .ZN(n15872) );
  OAI211_X1 U17994 ( .C1(n21735), .C2(n16280), .A(n15873), .B(n15872), .ZN(
        P1_U2888) );
  INV_X1 U17995 ( .A(n15898), .ZN(n15877) );
  AOI22_X1 U17996 ( .A1(n13631), .A2(n21518), .B1(n15926), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n15874) );
  OAI21_X1 U17997 ( .B1(n15877), .B2(n16237), .A(n15874), .ZN(P1_U2858) );
  INV_X1 U17998 ( .A(DATAI_14_), .ZN(n17410) );
  NAND2_X1 U17999 ( .A1(n15942), .A2(BUF1_REG_14__SCAN_IN), .ZN(n15875) );
  OAI21_X1 U18000 ( .B1(n15942), .B2(n17410), .A(n15875), .ZN(n21942) );
  AOI22_X1 U18001 ( .A1(n15920), .A2(n21942), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n16248), .ZN(n15876) );
  OAI21_X1 U18002 ( .B1(n15877), .B2(n16280), .A(n15876), .ZN(P1_U2890) );
  AOI21_X1 U18003 ( .B1(n15880), .B2(n15797), .A(n15879), .ZN(n18755) );
  INV_X1 U18004 ( .A(n18755), .ZN(n17084) );
  INV_X1 U18005 ( .A(n15946), .ZN(n15881) );
  AOI21_X1 U18006 ( .B1(n15882), .B2(n15638), .A(n15881), .ZN(n15928) );
  NAND2_X1 U18007 ( .A1(n15928), .A2(n16686), .ZN(n15884) );
  NAND2_X1 U18008 ( .A1(n16689), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n15883) );
  OAI211_X1 U18009 ( .C1(n17084), .C2(n16689), .A(n15884), .B(n15883), .ZN(
        P2_U2868) );
  INV_X1 U18010 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n21730) );
  INV_X1 U18011 ( .A(n16517), .ZN(n15886) );
  OAI21_X1 U18012 ( .B1(n15886), .B2(n15885), .A(n10955), .ZN(n21742) );
  OAI222_X1 U18013 ( .A1(n21735), .A2(n16237), .B1(n16246), .B2(n21730), .C1(
        n21742), .C2(n16247), .ZN(P1_U2856) );
  INV_X1 U18014 ( .A(n15888), .ZN(n15890) );
  OAI21_X1 U18015 ( .B1(n15887), .B2(n15890), .A(n15889), .ZN(n15892) );
  NAND2_X1 U18016 ( .A1(n15892), .A2(n15891), .ZN(n15894) );
  MUX2_X1 U18017 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n13025), .S(
        n12866), .Z(n15893) );
  XNOR2_X1 U18018 ( .A(n15894), .B(n15893), .ZN(n21519) );
  INV_X1 U18019 ( .A(n21519), .ZN(n15900) );
  AOI22_X1 U18020 ( .A1(n20192), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n16504), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n15895) );
  OAI21_X1 U18021 ( .B1(n20200), .B2(n15896), .A(n15895), .ZN(n15897) );
  AOI21_X1 U18022 ( .B1(n15898), .B2(n20186), .A(n15897), .ZN(n15899) );
  OAI21_X1 U18023 ( .B1(n15900), .B2(n21789), .A(n15899), .ZN(P1_U2985) );
  NOR2_X1 U18024 ( .A1(n15789), .A2(n15901), .ZN(n15902) );
  AOI21_X1 U18025 ( .B1(n15904), .B2(n15903), .A(n15902), .ZN(n15923) );
  INV_X1 U18026 ( .A(n15922), .ZN(n15905) );
  NOR2_X1 U18027 ( .A1(n15923), .A2(n15905), .ZN(n15908) );
  INV_X1 U18028 ( .A(n15925), .ZN(n15910) );
  AOI21_X1 U18029 ( .B1(n15910), .B2(n15924), .A(n15909), .ZN(n15911) );
  OR2_X1 U18030 ( .A1(n15911), .A2(n16514), .ZN(n16538) );
  INV_X1 U18031 ( .A(n16538), .ZN(n15912) );
  AOI22_X1 U18032 ( .A1(n15912), .A2(n21724), .B1(n21773), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n15913) );
  OAI211_X1 U18033 ( .C1(n21776), .C2(n15914), .A(n15913), .B(n21729), .ZN(
        n15917) );
  AOI211_X1 U18034 ( .C1(n21712), .C2(n20063), .A(n21710), .B(n15915), .ZN(
        n15916) );
  AOI211_X1 U18035 ( .C1(n16400), .C2(n21782), .A(n15917), .B(n15916), .ZN(
        n15918) );
  OAI21_X1 U18036 ( .B1(n16403), .B2(n21777), .A(n15918), .ZN(P1_U2827) );
  INV_X1 U18037 ( .A(DATAI_13_), .ZN(n17525) );
  NAND2_X1 U18038 ( .A1(n15942), .A2(BUF1_REG_13__SCAN_IN), .ZN(n15919) );
  OAI21_X1 U18039 ( .B1(n15942), .B2(n17525), .A(n15919), .ZN(n21933) );
  AOI22_X1 U18040 ( .A1(n15920), .A2(n21933), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n16248), .ZN(n15921) );
  OAI21_X1 U18041 ( .B1(n16403), .B2(n16280), .A(n15921), .ZN(P1_U2891) );
  XNOR2_X1 U18042 ( .A(n15923), .B(n15922), .ZN(n20164) );
  XNOR2_X1 U18043 ( .A(n15925), .B(n15924), .ZN(n21703) );
  AOI22_X1 U18044 ( .A1(n13631), .A2(n21703), .B1(n15926), .B2(
        P1_EBX_REG_12__SCAN_IN), .ZN(n15927) );
  OAI21_X1 U18045 ( .B1(n21716), .B2(n16237), .A(n15927), .ZN(P1_U2860) );
  INV_X1 U18046 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n15935) );
  NAND2_X1 U18047 ( .A1(n15928), .A2(n19586), .ZN(n15934) );
  XNOR2_X1 U18048 ( .A(n15929), .B(n15642), .ZN(n18759) );
  OAI22_X1 U18049 ( .A1(n16765), .A2(n18759), .B1(n19374), .B2(n15930), .ZN(
        n15932) );
  NOR2_X1 U18050 ( .A1(n16766), .A2(n19712), .ZN(n15931) );
  AOI211_X1 U18051 ( .C1(BUF1_REG_19__SCAN_IN), .C2(n19582), .A(n15932), .B(
        n15931), .ZN(n15933) );
  OAI211_X1 U18052 ( .C1(n16755), .C2(n15935), .A(n15934), .B(n15933), .ZN(
        P2_U2900) );
  INV_X1 U18053 ( .A(n15936), .ZN(n15938) );
  INV_X1 U18054 ( .A(n15834), .ZN(n15937) );
  AOI21_X1 U18055 ( .B1(n15938), .B2(n15937), .A(n15862), .ZN(n21725) );
  INV_X1 U18056 ( .A(n21725), .ZN(n15940) );
  OAI222_X1 U18057 ( .A1(n15940), .A2(n16280), .B1(n15944), .B2(n15939), .C1(
        n16273), .C2(n20045), .ZN(P1_U2889) );
  INV_X1 U18058 ( .A(DATAI_12_), .ZN(n17529) );
  NAND2_X1 U18059 ( .A1(n15942), .A2(BUF1_REG_12__SCAN_IN), .ZN(n15941) );
  OAI21_X1 U18060 ( .B1(n15942), .B2(n17529), .A(n15941), .ZN(n21923) );
  INV_X1 U18061 ( .A(n21923), .ZN(n15943) );
  OAI222_X1 U18062 ( .A1(n21716), .A2(n16280), .B1(n15944), .B2(n15943), .C1(
        n21929), .C2(n16273), .ZN(P1_U2892) );
  INV_X1 U18063 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n15945) );
  OAI222_X1 U18064 ( .A1(n16538), .A2(n16247), .B1(n15945), .B2(n20137), .C1(
        n16403), .C2(n16237), .ZN(P1_U2859) );
  INV_X1 U18065 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n15956) );
  AOI21_X1 U18066 ( .B1(n15947), .B2(n15946), .A(n16691), .ZN(n15957) );
  NAND2_X1 U18067 ( .A1(n15957), .A2(n19586), .ZN(n15955) );
  OR2_X1 U18068 ( .A1(n15950), .A2(n15949), .ZN(n15951) );
  AND2_X1 U18069 ( .A1(n15948), .A2(n15951), .ZN(n18762) );
  AOI22_X1 U18070 ( .A1(n19585), .A2(n18762), .B1(n19579), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n15952) );
  OAI21_X1 U18071 ( .B1(n19672), .B2(n16766), .A(n15952), .ZN(n15953) );
  AOI21_X1 U18072 ( .B1(n19582), .B2(BUF1_REG_20__SCAN_IN), .A(n15953), .ZN(
        n15954) );
  OAI211_X1 U18073 ( .C1(n16755), .C2(n15956), .A(n15955), .B(n15954), .ZN(
        P2_U2899) );
  NAND2_X1 U18074 ( .A1(n15957), .A2(n16686), .ZN(n15963) );
  NAND2_X1 U18075 ( .A1(n15959), .A2(n15958), .ZN(n15960) );
  NAND2_X1 U18076 ( .A1(n16693), .A2(n15960), .ZN(n18769) );
  INV_X1 U18077 ( .A(n18769), .ZN(n15961) );
  NAND2_X1 U18078 ( .A1(n15961), .A2(n16651), .ZN(n15962) );
  OAI211_X1 U18079 ( .C1(n16651), .C2(n11896), .A(n15963), .B(n15962), .ZN(
        P2_U2867) );
  OR2_X1 U18080 ( .A1(n15861), .A2(n15964), .ZN(n15966) );
  AND2_X1 U18081 ( .A1(n15966), .A2(n15965), .ZN(n20173) );
  INV_X1 U18082 ( .A(n20173), .ZN(n15970) );
  AOI22_X1 U18083 ( .A1(n16295), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n16248), .ZN(n15969) );
  AOI22_X1 U18084 ( .A1(n16298), .A2(n15967), .B1(n16296), .B2(DATAI_17_), 
        .ZN(n15968) );
  OAI211_X1 U18085 ( .C1(n15970), .C2(n16280), .A(n15969), .B(n15968), .ZN(
        P1_U2887) );
  INV_X1 U18086 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n20641) );
  NAND4_X1 U18087 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_24__SCAN_IN), 
        .A3(P3_EBX_REG_21__SCAN_IN), .A4(n17936), .ZN(n15971) );
  NOR4_X1 U18088 ( .A1(n20659), .A2(n20641), .A3(n15972), .A4(n15971), .ZN(
        n17933) );
  NAND2_X1 U18089 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n17933), .ZN(n15973) );
  NOR2_X1 U18090 ( .A1(n20801), .A2(n15973), .ZN(n15975) );
  NAND2_X1 U18091 ( .A1(n18043), .A2(n15973), .ZN(n17934) );
  INV_X1 U18092 ( .A(n17934), .ZN(n15974) );
  MUX2_X1 U18093 ( .A(n15975), .B(n15974), .S(P3_EBX_REG_31__SCAN_IN), .Z(
        P3_U2672) );
  XNOR2_X1 U18094 ( .A(n15982), .B(n15981), .ZN(n16071) );
  INV_X1 U18095 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17003) );
  AOI21_X1 U18096 ( .B1(n17003), .B2(n15984), .A(n15983), .ZN(n16069) );
  AND2_X1 U18097 ( .A1(n15986), .A2(n15985), .ZN(n15987) );
  OR2_X1 U18098 ( .A1(n15987), .A2(n16635), .ZN(n18841) );
  INV_X1 U18099 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n17760) );
  NOR2_X1 U18100 ( .A1(n16970), .A2(n17760), .ZN(n16063) );
  NOR2_X1 U18101 ( .A1(n17631), .A2(n18844), .ZN(n15988) );
  AOI211_X1 U18102 ( .C1(n17661), .C2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16063), .B(n15988), .ZN(n15989) );
  OAI21_X1 U18103 ( .B1(n18841), .B2(n17651), .A(n15989), .ZN(n15990) );
  AOI21_X1 U18104 ( .B1(n16069), .B2(n17668), .A(n15990), .ZN(n15991) );
  OAI21_X1 U18105 ( .B1(n16071), .B2(n17670), .A(n15991), .ZN(P2_U2986) );
  NOR2_X1 U18106 ( .A1(n15992), .A2(n17277), .ZN(n16006) );
  INV_X1 U18107 ( .A(n16074), .ZN(n15994) );
  OAI21_X1 U18108 ( .B1(n18890), .B2(n16041), .A(n16065), .ZN(n16046) );
  INV_X1 U18109 ( .A(n16046), .ZN(n15998) );
  AOI21_X1 U18110 ( .B1(n15996), .B2(n15995), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15997) );
  OR2_X1 U18111 ( .A1(n15998), .A2(n15997), .ZN(n16001) );
  INV_X1 U18112 ( .A(n15999), .ZN(n16000) );
  AND2_X1 U18113 ( .A1(n16001), .A2(n16000), .ZN(n16002) );
  NAND2_X1 U18114 ( .A1(n16004), .A2(n11229), .ZN(n16005) );
  OAI21_X1 U18115 ( .B1(n16008), .B2(n18881), .A(n16007), .ZN(P2_U3016) );
  OAI21_X1 U18116 ( .B1(n16011), .B2(n16010), .A(n16009), .ZN(n17605) );
  NAND2_X1 U18117 ( .A1(n16013), .A2(n16012), .ZN(n16016) );
  INV_X1 U18118 ( .A(n16014), .ZN(n16015) );
  NAND2_X1 U18119 ( .A1(n16016), .A2(n16015), .ZN(n16018) );
  AND2_X1 U18120 ( .A1(n16018), .A2(n16017), .ZN(n17606) );
  INV_X1 U18121 ( .A(n16019), .ZN(n16020) );
  NAND2_X1 U18122 ( .A1(n16021), .A2(n16020), .ZN(n16022) );
  AOI22_X1 U18123 ( .A1(n12326), .A2(n17606), .B1(n17103), .B2(n16022), .ZN(
        n16023) );
  NAND2_X1 U18124 ( .A1(n12161), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n17609) );
  OAI211_X1 U18125 ( .C1(n17277), .C2(n17605), .A(n16023), .B(n17609), .ZN(
        n16031) );
  AOI21_X1 U18126 ( .B1(n17104), .B2(n16024), .A(n18877), .ZN(n16029) );
  INV_X1 U18127 ( .A(n16024), .ZN(n16025) );
  NAND2_X1 U18128 ( .A1(n16026), .A2(n16025), .ZN(n16027) );
  OAI21_X1 U18129 ( .B1(n16029), .B2(n16028), .A(n16027), .ZN(n16030) );
  AOI211_X1 U18130 ( .C1(n18876), .C2(n17682), .A(n16031), .B(n16030), .ZN(
        n16032) );
  OAI21_X1 U18131 ( .B1(n16033), .B2(n18885), .A(n16032), .ZN(P2_U3044) );
  OAI211_X2 U18132 ( .C1(n16036), .C2(n16035), .A(n16034), .B(n16782), .ZN(
        n16040) );
  NAND2_X1 U18133 ( .A1(n16037), .A2(n12190), .ZN(n16038) );
  XNOR2_X1 U18134 ( .A(n16038), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16039) );
  XNOR2_X1 U18135 ( .A(n16040), .B(n16039), .ZN(n16781) );
  NOR2_X1 U18136 ( .A1(n16970), .A2(n17764), .ZN(n16775) );
  INV_X1 U18137 ( .A(n16041), .ZN(n16042) );
  NOR3_X1 U18138 ( .A1(n17001), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n16042), .ZN(n16043) );
  XNOR2_X1 U18139 ( .A(n16045), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16779) );
  OAI21_X1 U18140 ( .B1(n16781), .B2(n18881), .A(n16050), .ZN(P2_U3015) );
  INV_X1 U18141 ( .A(n16316), .ZN(n16059) );
  OAI22_X1 U18142 ( .A1(n21776), .A2(n16314), .B1(n21761), .B2(n16051), .ZN(
        n16055) );
  INV_X1 U18143 ( .A(n16312), .ZN(n16053) );
  XNOR2_X1 U18144 ( .A(n16080), .B(P1_REIP_REG_30__SCAN_IN), .ZN(n16052) );
  OAI22_X1 U18145 ( .A1(n21702), .A2(n16053), .B1(n21710), .B2(n16052), .ZN(
        n16054) );
  AOI211_X1 U18146 ( .C1(n16412), .C2(n21724), .A(n16055), .B(n16054), .ZN(
        n16056) );
  OAI21_X1 U18147 ( .B1(n16059), .B2(n21777), .A(n16056), .ZN(P1_U2810) );
  AOI22_X1 U18148 ( .A1(n16295), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n16248), .ZN(n16058) );
  AOI22_X1 U18149 ( .A1(n16298), .A2(n21942), .B1(n16296), .B2(DATAI_30_), 
        .ZN(n16057) );
  OAI211_X1 U18150 ( .C1(n16059), .C2(n16280), .A(n16058), .B(n16057), .ZN(
        P1_U2874) );
  XNOR2_X1 U18151 ( .A(n14510), .B(n11163), .ZN(n18839) );
  NOR3_X1 U18152 ( .A1(n17001), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n16061), .ZN(n16062) );
  AOI211_X1 U18153 ( .C1(n18876), .C2(n18839), .A(n16063), .B(n16062), .ZN(
        n16067) );
  NAND2_X1 U18154 ( .A1(n16065), .A2(n16064), .ZN(n17008) );
  NAND2_X1 U18155 ( .A1(n17008), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16066) );
  OAI211_X1 U18156 ( .C1(n18841), .C2(n18885), .A(n16067), .B(n16066), .ZN(
        n16068) );
  AOI21_X1 U18157 ( .B1(n16069), .B2(n18879), .A(n16068), .ZN(n16070) );
  OAI21_X1 U18158 ( .B1(n16071), .B2(n18881), .A(n16070), .ZN(P2_U3018) );
  AOI22_X1 U18159 ( .A1(n19581), .A2(n19361), .B1(n19579), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n16073) );
  NAND2_X1 U18160 ( .A1(n19582), .A2(BUF1_REG_30__SCAN_IN), .ZN(n16072) );
  OAI211_X1 U18161 ( .C1(n16074), .C2(n16765), .A(n16073), .B(n16072), .ZN(
        n16075) );
  AOI21_X1 U18162 ( .B1(n19583), .B2(BUF2_REG_30__SCAN_IN), .A(n16075), .ZN(
        n16076) );
  OAI21_X1 U18163 ( .B1(n16077), .B2(n16771), .A(n16076), .ZN(P2_U2889) );
  NAND2_X1 U18164 ( .A1(n16325), .A2(n21754), .ZN(n16086) );
  INV_X1 U18165 ( .A(n16323), .ZN(n16084) );
  OAI22_X1 U18166 ( .A1(n21776), .A2(n16079), .B1(n21761), .B2(n16078), .ZN(
        n16083) );
  NAND2_X1 U18167 ( .A1(n21738), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n16081) );
  AOI21_X1 U18168 ( .B1(n16081), .B2(n16092), .A(n16080), .ZN(n16082) );
  AOI211_X1 U18169 ( .C1(n21782), .C2(n16084), .A(n16083), .B(n16082), .ZN(
        n16085) );
  OAI211_X1 U18170 ( .C1(n21788), .C2(n16415), .A(n16086), .B(n16085), .ZN(
        P1_U2811) );
  AND2_X1 U18171 ( .A1(n16102), .A2(n16087), .ZN(n16089) );
  OR2_X1 U18172 ( .A1(n16089), .A2(n16088), .ZN(n16427) );
  INV_X1 U18173 ( .A(n16258), .ZN(n16090) );
  NAND2_X1 U18174 ( .A1(n16090), .A2(n21754), .ZN(n16099) );
  INV_X1 U18175 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n16209) );
  OAI22_X1 U18176 ( .A1(n21776), .A2(n16091), .B1(n21761), .B2(n16209), .ZN(
        n16096) );
  NAND2_X1 U18177 ( .A1(n21738), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n16094) );
  INV_X1 U18178 ( .A(n16092), .ZN(n16093) );
  AOI21_X1 U18179 ( .B1(n16094), .B2(n16110), .A(n16093), .ZN(n16095) );
  AOI211_X1 U18180 ( .C1(n21782), .C2(n16097), .A(n16096), .B(n16095), .ZN(
        n16098) );
  OAI211_X1 U18181 ( .C1(n21788), .C2(n16427), .A(n16099), .B(n16098), .ZN(
        P1_U2812) );
  NAND2_X1 U18182 ( .A1(n16116), .A2(n16100), .ZN(n16101) );
  NAND2_X1 U18183 ( .A1(n16102), .A2(n16101), .ZN(n21575) );
  AOI21_X1 U18184 ( .B1(n16104), .B2(n16114), .A(n13686), .ZN(n16331) );
  NAND2_X1 U18185 ( .A1(n16331), .A2(n21754), .ZN(n16112) );
  INV_X1 U18186 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21578) );
  INV_X1 U18187 ( .A(n16123), .ZN(n16105) );
  OAI21_X1 U18188 ( .B1(n21710), .B2(n21578), .A(n16105), .ZN(n16109) );
  OAI22_X1 U18189 ( .A1(n21776), .A2(n16106), .B1(n21761), .B2(n16210), .ZN(
        n16108) );
  NOR2_X1 U18190 ( .A1(n21702), .A2(n16329), .ZN(n16107) );
  AOI211_X1 U18191 ( .C1(n16110), .C2(n16109), .A(n16108), .B(n16107), .ZN(
        n16111) );
  OAI211_X1 U18192 ( .C1(n21788), .C2(n21575), .A(n16112), .B(n16111), .ZN(
        P1_U2813) );
  OAI21_X1 U18193 ( .B1(n16129), .B2(n16117), .A(n16116), .ZN(n16438) );
  INV_X1 U18194 ( .A(n16438), .ZN(n16125) );
  INV_X1 U18195 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20082) );
  INV_X1 U18196 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n16118) );
  NOR2_X1 U18197 ( .A1(n20082), .A2(n16118), .ZN(n16119) );
  AOI22_X1 U18198 ( .A1(n21738), .A2(P1_REIP_REG_26__SCAN_IN), .B1(n21785), 
        .B2(n16119), .ZN(n16122) );
  AOI22_X1 U18199 ( .A1(n21748), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(
        n21773), .B2(P1_EBX_REG_26__SCAN_IN), .ZN(n16121) );
  NAND2_X1 U18200 ( .A1(n21782), .A2(n16340), .ZN(n16120) );
  OAI211_X1 U18201 ( .C1(n16123), .C2(n16122), .A(n16121), .B(n16120), .ZN(
        n16124) );
  AOI21_X1 U18202 ( .B1(n16125), .B2(n21724), .A(n16124), .ZN(n16126) );
  OAI21_X1 U18203 ( .B1(n16337), .B2(n21777), .A(n16126), .ZN(P1_U2814) );
  AOI21_X1 U18204 ( .B1(n16128), .B2(n16214), .A(n16113), .ZN(n16349) );
  INV_X1 U18205 ( .A(n16349), .ZN(n16269) );
  INV_X1 U18206 ( .A(n16129), .ZN(n16132) );
  NAND2_X1 U18207 ( .A1(n16219), .A2(n16130), .ZN(n16131) );
  NAND2_X1 U18208 ( .A1(n16132), .A2(n16131), .ZN(n16212) );
  INV_X1 U18209 ( .A(n16212), .ZN(n21588) );
  OAI22_X1 U18210 ( .A1(n21761), .A2(n16213), .B1(P1_REIP_REG_25__SCAN_IN), 
        .B2(n16133), .ZN(n16134) );
  AOI21_X1 U18211 ( .B1(n21748), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16134), .ZN(n16135) );
  OAI21_X1 U18212 ( .B1(n16347), .B2(n21702), .A(n16135), .ZN(n16141) );
  INV_X1 U18213 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20078) );
  INV_X1 U18214 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n21599) );
  INV_X1 U18215 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21655) );
  NAND3_X1 U18216 ( .A1(n16137), .A2(P1_REIP_REG_6__SCAN_IN), .A3(n16136), 
        .ZN(n21636) );
  NOR3_X1 U18217 ( .A1(n16138), .A2(n21655), .A3(n21636), .ZN(n21684) );
  NAND2_X1 U18218 ( .A1(n16139), .A2(n21684), .ZN(n16176) );
  NOR4_X1 U18219 ( .A1(n20076), .A2(n20078), .A3(n21599), .A4(n16176), .ZN(
        n16150) );
  AOI211_X1 U18220 ( .C1(n16150), .C2(P1_REIP_REG_24__SCAN_IN), .A(n21710), 
        .B(n20082), .ZN(n16140) );
  AOI211_X1 U18221 ( .C1(n21724), .C2(n21588), .A(n16141), .B(n16140), .ZN(
        n16142) );
  OAI21_X1 U18222 ( .B1(n16269), .B2(n21777), .A(n16142), .ZN(P1_U2815) );
  AND2_X1 U18223 ( .A1(n16159), .A2(n16144), .ZN(n16146) );
  OR2_X1 U18224 ( .A1(n16146), .A2(n16145), .ZN(n20195) );
  OR2_X1 U18225 ( .A1(n10972), .A2(n16147), .ZN(n16148) );
  NAND2_X1 U18226 ( .A1(n16217), .A2(n16148), .ZN(n16223) );
  INV_X1 U18227 ( .A(n16223), .ZN(n21594) );
  INV_X1 U18228 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16149) );
  NOR2_X1 U18229 ( .A1(n21776), .A2(n16149), .ZN(n16155) );
  NOR2_X1 U18230 ( .A1(n21710), .A2(n16150), .ZN(n21772) );
  NAND2_X1 U18231 ( .A1(n16151), .A2(n21599), .ZN(n16152) );
  AOI22_X1 U18232 ( .A1(n21773), .A2(P1_EBX_REG_23__SCAN_IN), .B1(n21772), 
        .B2(n16152), .ZN(n16153) );
  OAI21_X1 U18233 ( .B1(n21702), .B2(n20199), .A(n16153), .ZN(n16154) );
  AOI211_X1 U18234 ( .C1(n21594), .C2(n21724), .A(n16155), .B(n16154), .ZN(
        n16156) );
  OAI21_X1 U18235 ( .B1(n20195), .B2(n21777), .A(n16156), .ZN(P1_U2817) );
  AOI21_X1 U18236 ( .B1(n16160), .B2(n16158), .A(n16143), .ZN(n16364) );
  INV_X1 U18237 ( .A(n16364), .ZN(n16284) );
  NAND2_X1 U18238 ( .A1(n16175), .A2(n16162), .ZN(n16163) );
  NAND2_X1 U18239 ( .A1(n10973), .A2(n16163), .ZN(n16459) );
  NOR2_X1 U18240 ( .A1(n16459), .A2(n21788), .ZN(n16168) );
  NAND2_X1 U18241 ( .A1(n21782), .A2(n16360), .ZN(n16166) );
  NOR3_X1 U18242 ( .A1(n16169), .A2(n21710), .A3(n20078), .ZN(n16164) );
  AOI21_X1 U18243 ( .B1(n21773), .B2(P1_EBX_REG_22__SCAN_IN), .A(n16164), .ZN(
        n16165) );
  OAI211_X1 U18244 ( .C1(n21776), .C2(n13433), .A(n16166), .B(n16165), .ZN(
        n16167) );
  AOI211_X1 U18245 ( .C1(n16169), .C2(n20078), .A(n16168), .B(n16167), .ZN(
        n16170) );
  OAI21_X1 U18246 ( .B1(n16284), .B2(n21777), .A(n16170), .ZN(P1_U2818) );
  OAI21_X1 U18247 ( .B1(n16171), .B2(n16172), .A(n16158), .ZN(n20185) );
  NAND2_X1 U18248 ( .A1(n16233), .A2(n16173), .ZN(n16174) );
  NAND2_X1 U18249 ( .A1(n16175), .A2(n16174), .ZN(n16226) );
  INV_X1 U18250 ( .A(n16226), .ZN(n21569) );
  NAND2_X1 U18251 ( .A1(n21738), .A2(n16176), .ZN(n21770) );
  INV_X1 U18252 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16180) );
  INV_X1 U18253 ( .A(n20191), .ZN(n16177) );
  NAND2_X1 U18254 ( .A1(n21782), .A2(n16177), .ZN(n16179) );
  NAND2_X1 U18255 ( .A1(n21773), .A2(P1_EBX_REG_21__SCAN_IN), .ZN(n16178) );
  OAI211_X1 U18256 ( .C1(n16180), .C2(n21776), .A(n16179), .B(n16178), .ZN(
        n16181) );
  INV_X1 U18257 ( .A(n16181), .ZN(n16182) );
  OAI221_X1 U18258 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n16183), .C1(n20076), 
        .C2(n21770), .A(n16182), .ZN(n16184) );
  AOI21_X1 U18259 ( .B1(n21569), .B2(n21724), .A(n16184), .ZN(n16185) );
  OAI21_X1 U18260 ( .B1(n20185), .B2(n21777), .A(n16185), .ZN(P1_U2819) );
  AOI21_X1 U18261 ( .B1(n16188), .B2(n15965), .A(n16187), .ZN(n16379) );
  INV_X1 U18262 ( .A(n16379), .ZN(n16301) );
  INV_X1 U18263 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20070) );
  INV_X1 U18264 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20067) );
  NAND2_X1 U18265 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n21739), .ZN(n21737) );
  NOR2_X1 U18266 ( .A1(n21759), .A2(n21710), .ZN(n21753) );
  INV_X1 U18267 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21743) );
  NOR2_X1 U18268 ( .A1(n16198), .A2(n16189), .ZN(n16190) );
  OR2_X1 U18269 ( .A1(n16239), .A2(n16190), .ZN(n16495) );
  INV_X1 U18270 ( .A(n21729), .ZN(n21745) );
  AOI21_X1 U18271 ( .B1(n21748), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n21745), .ZN(n16192) );
  AOI22_X1 U18272 ( .A1(n21782), .A2(n16375), .B1(P1_EBX_REG_18__SCAN_IN), 
        .B2(n21773), .ZN(n16191) );
  OAI211_X1 U18273 ( .C1(n21788), .C2(n16495), .A(n16192), .B(n16191), .ZN(
        n16193) );
  AOI221_X1 U18274 ( .B1(n21753), .B2(P1_REIP_REG_18__SCAN_IN), .C1(n21759), 
        .C2(n21743), .A(n16193), .ZN(n16194) );
  OAI21_X1 U18275 ( .B1(n16301), .B2(n21777), .A(n16194), .ZN(P1_U2822) );
  NOR2_X1 U18276 ( .A1(n21776), .A2(n16195), .ZN(n16203) );
  AND2_X1 U18277 ( .A1(n10955), .A2(n16196), .ZN(n16197) );
  NOR2_X1 U18278 ( .A1(n16198), .A2(n16197), .ZN(n20123) );
  NAND2_X1 U18279 ( .A1(n20123), .A2(n21724), .ZN(n16201) );
  NAND2_X1 U18280 ( .A1(n21782), .A2(n20171), .ZN(n16200) );
  NAND2_X1 U18281 ( .A1(n21773), .A2(P1_EBX_REG_17__SCAN_IN), .ZN(n16199) );
  NAND4_X1 U18282 ( .A1(n16201), .A2(n21729), .A3(n16200), .A4(n16199), .ZN(
        n16202) );
  AOI211_X1 U18283 ( .C1(n20173), .C2(n21754), .A(n16203), .B(n16202), .ZN(
        n16206) );
  NAND2_X1 U18284 ( .A1(n20070), .A2(n21737), .ZN(n16204) );
  NAND2_X1 U18285 ( .A1(n21753), .A2(n16204), .ZN(n16205) );
  NAND2_X1 U18286 ( .A1(n16206), .A2(n16205), .ZN(P1_U2823) );
  OAI22_X1 U18287 ( .A1(n16208), .A2(n16247), .B1(n16207), .B2(n20137), .ZN(
        P1_U2841) );
  OAI222_X1 U18288 ( .A1(n16209), .A2(n20137), .B1(n16247), .B2(n16427), .C1(
        n16258), .C2(n16237), .ZN(P1_U2844) );
  INV_X1 U18289 ( .A(n16331), .ZN(n16262) );
  OAI222_X1 U18290 ( .A1(n16210), .A2(n20137), .B1(n16247), .B2(n21575), .C1(
        n16262), .C2(n16237), .ZN(P1_U2845) );
  INV_X1 U18291 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n16211) );
  OAI222_X1 U18292 ( .A1(n16211), .A2(n20137), .B1(n16247), .B2(n16438), .C1(
        n16337), .C2(n16237), .ZN(P1_U2846) );
  OAI222_X1 U18293 ( .A1(n16213), .A2(n20137), .B1(n16247), .B2(n16212), .C1(
        n16269), .C2(n16237), .ZN(P1_U2847) );
  NAND2_X1 U18294 ( .A1(n16217), .A2(n16216), .ZN(n16218) );
  NAND2_X1 U18295 ( .A1(n16219), .A2(n16218), .ZN(n21787) );
  OAI22_X1 U18296 ( .A1(n21787), .A2(n16247), .B1(n16220), .B2(n20137), .ZN(
        n16221) );
  INV_X1 U18297 ( .A(n16221), .ZN(n16222) );
  OAI21_X1 U18298 ( .B1(n21778), .B2(n16237), .A(n16222), .ZN(P1_U2848) );
  INV_X1 U18299 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n16224) );
  OAI222_X1 U18300 ( .A1(n16224), .A2(n20137), .B1(n16247), .B2(n16223), .C1(
        n20195), .C2(n16237), .ZN(P1_U2849) );
  INV_X1 U18301 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n16225) );
  OAI222_X1 U18302 ( .A1(n16237), .A2(n16284), .B1(n16246), .B2(n16225), .C1(
        n16459), .C2(n16247), .ZN(P1_U2850) );
  INV_X1 U18303 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n16227) );
  OAI222_X1 U18304 ( .A1(n16227), .A2(n20137), .B1(n16237), .B2(n20185), .C1(
        n16226), .C2(n16247), .ZN(P1_U2851) );
  NOR2_X1 U18305 ( .A1(n16228), .A2(n16229), .ZN(n16230) );
  OR2_X1 U18306 ( .A1(n16171), .A2(n16230), .ZN(n21765) );
  INV_X1 U18307 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n21762) );
  NAND2_X1 U18308 ( .A1(n16241), .A2(n16231), .ZN(n16232) );
  AND2_X1 U18309 ( .A1(n16233), .A2(n16232), .ZN(n16473) );
  INV_X1 U18310 ( .A(n16473), .ZN(n21764) );
  OAI222_X1 U18311 ( .A1(n16237), .A2(n21765), .B1(n16246), .B2(n21762), .C1(
        n21764), .C2(n16247), .ZN(P1_U2852) );
  AND2_X1 U18312 ( .A1(n16235), .A2(n16234), .ZN(n16236) );
  NOR2_X1 U18313 ( .A1(n16228), .A2(n16236), .ZN(n21755) );
  OR2_X1 U18314 ( .A1(n16239), .A2(n16238), .ZN(n16240) );
  NAND2_X1 U18315 ( .A1(n16241), .A2(n16240), .ZN(n21751) );
  OAI22_X1 U18316 ( .A1(n21751), .A2(n16247), .B1(n16242), .B2(n20137), .ZN(
        n16243) );
  AOI21_X1 U18317 ( .B1(n21755), .B2(n13627), .A(n16243), .ZN(n16244) );
  INV_X1 U18318 ( .A(n16244), .ZN(P1_U2853) );
  INV_X1 U18319 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n16245) );
  OAI222_X1 U18320 ( .A1(n16495), .A2(n16247), .B1(n16246), .B2(n16245), .C1(
        n16237), .C2(n16301), .ZN(P1_U2854) );
  NOR2_X1 U18321 ( .A1(n16248), .A2(n14811), .ZN(n16249) );
  NAND2_X1 U18322 ( .A1(n16250), .A2(n16249), .ZN(n16252) );
  AOI22_X1 U18323 ( .A1(n16296), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n16248), .ZN(n16251) );
  OAI211_X1 U18324 ( .C1(n16265), .C2(n20270), .A(n16252), .B(n16251), .ZN(
        P1_U2873) );
  INV_X1 U18325 ( .A(n16325), .ZN(n16255) );
  AOI22_X1 U18326 ( .A1(n16295), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n16248), .ZN(n16254) );
  AOI22_X1 U18327 ( .A1(n16298), .A2(n21933), .B1(n16296), .B2(DATAI_29_), 
        .ZN(n16253) );
  OAI211_X1 U18328 ( .C1(n16255), .C2(n16280), .A(n16254), .B(n16253), .ZN(
        P1_U2875) );
  AOI22_X1 U18329 ( .A1(n16295), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n16248), .ZN(n16257) );
  AOI22_X1 U18330 ( .A1(n16298), .A2(n21923), .B1(n16296), .B2(DATAI_28_), 
        .ZN(n16256) );
  OAI211_X1 U18331 ( .C1(n16258), .C2(n16280), .A(n16257), .B(n16256), .ZN(
        P1_U2876) );
  NOR2_X1 U18332 ( .A1(n16265), .A2(n20262), .ZN(n16260) );
  INV_X1 U18333 ( .A(n16298), .ZN(n16276) );
  INV_X1 U18334 ( .A(n16296), .ZN(n16274) );
  OAI22_X1 U18335 ( .A1(n16276), .A2(n21912), .B1(n16274), .B2(n17500), .ZN(
        n16259) );
  AOI211_X1 U18336 ( .C1(n16248), .C2(P1_EAX_REG_27__SCAN_IN), .A(n16260), .B(
        n16259), .ZN(n16261) );
  OAI21_X1 U18337 ( .B1(n16262), .B2(n16280), .A(n16261), .ZN(P1_U2877) );
  AOI22_X1 U18338 ( .A1(n16295), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n16248), .ZN(n16264) );
  AOI22_X1 U18339 ( .A1(n16298), .A2(n21903), .B1(n16296), .B2(DATAI_26_), 
        .ZN(n16263) );
  OAI211_X1 U18340 ( .C1(n16337), .C2(n16280), .A(n16264), .B(n16263), .ZN(
        P1_U2878) );
  OAI22_X1 U18341 ( .A1(n16265), .A2(n20257), .B1(n21896), .B2(n16273), .ZN(
        n16267) );
  NOR2_X1 U18342 ( .A1(n16276), .A2(n21892), .ZN(n16266) );
  AOI211_X1 U18343 ( .C1(n16296), .C2(DATAI_25_), .A(n16267), .B(n16266), .ZN(
        n16268) );
  OAI21_X1 U18344 ( .B1(n16269), .B2(n16280), .A(n16268), .ZN(P1_U2879) );
  AOI22_X1 U18345 ( .A1(n16295), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n16248), .ZN(n16271) );
  AOI22_X1 U18346 ( .A1(n16298), .A2(n21884), .B1(n16296), .B2(DATAI_24_), 
        .ZN(n16270) );
  OAI211_X1 U18347 ( .C1(n21778), .C2(n16280), .A(n16271), .B(n16270), .ZN(
        P1_U2880) );
  NOR2_X1 U18348 ( .A1(n16273), .A2(n16272), .ZN(n16278) );
  OAI22_X1 U18349 ( .A1(n16276), .A2(n16275), .B1(n16274), .B2(n17495), .ZN(
        n16277) );
  AOI211_X1 U18350 ( .C1(BUF1_REG_23__SCAN_IN), .C2(n16295), .A(n16278), .B(
        n16277), .ZN(n16279) );
  OAI21_X1 U18351 ( .B1(n20195), .B2(n16280), .A(n16279), .ZN(P1_U2881) );
  AOI22_X1 U18352 ( .A1(n16295), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n16248), .ZN(n16283) );
  AOI22_X1 U18353 ( .A1(n16298), .A2(n16281), .B1(n16296), .B2(DATAI_22_), 
        .ZN(n16282) );
  OAI211_X1 U18354 ( .C1(n16284), .C2(n16280), .A(n16283), .B(n16282), .ZN(
        P1_U2882) );
  AOI22_X1 U18355 ( .A1(n16295), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n16248), .ZN(n16287) );
  AOI22_X1 U18356 ( .A1(n16298), .A2(n16285), .B1(n16296), .B2(DATAI_21_), 
        .ZN(n16286) );
  OAI211_X1 U18357 ( .C1(n20185), .C2(n16280), .A(n16287), .B(n16286), .ZN(
        P1_U2883) );
  AOI22_X1 U18358 ( .A1(n16295), .A2(BUF1_REG_20__SCAN_IN), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(n16248), .ZN(n16290) );
  AOI22_X1 U18359 ( .A1(n16298), .A2(n16288), .B1(n16296), .B2(DATAI_20_), 
        .ZN(n16289) );
  OAI211_X1 U18360 ( .C1(n21765), .C2(n16280), .A(n16290), .B(n16289), .ZN(
        P1_U2884) );
  INV_X1 U18361 ( .A(n21755), .ZN(n16294) );
  AOI22_X1 U18362 ( .A1(n16295), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n16248), .ZN(n16293) );
  AOI22_X1 U18363 ( .A1(n16298), .A2(n16291), .B1(n16296), .B2(DATAI_19_), 
        .ZN(n16292) );
  OAI211_X1 U18364 ( .C1(n16294), .C2(n16280), .A(n16293), .B(n16292), .ZN(
        P1_U2885) );
  AOI22_X1 U18365 ( .A1(n16295), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n16248), .ZN(n16300) );
  AOI22_X1 U18366 ( .A1(n16298), .A2(n16297), .B1(n16296), .B2(DATAI_18_), 
        .ZN(n16299) );
  OAI211_X1 U18367 ( .C1(n16301), .C2(n16280), .A(n16300), .B(n16299), .ZN(
        P1_U2886) );
  INV_X1 U18368 ( .A(n16303), .ZN(n16307) );
  NOR2_X1 U18369 ( .A1(n20182), .A2(n16425), .ZN(n16305) );
  INV_X1 U18370 ( .A(n16318), .ZN(n16308) );
  NAND2_X1 U18371 ( .A1(n16309), .A2(n16308), .ZN(n16311) );
  XNOR2_X1 U18372 ( .A(n16311), .B(n16310), .ZN(n16414) );
  NAND2_X1 U18373 ( .A1(n20172), .A2(n16312), .ZN(n16313) );
  NAND2_X1 U18374 ( .A1(n21585), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n16407) );
  OAI211_X1 U18375 ( .C1(n16314), .C2(n20155), .A(n16313), .B(n16407), .ZN(
        n16315) );
  AOI21_X1 U18376 ( .B1(n16316), .B2(n20186), .A(n16315), .ZN(n16317) );
  OAI21_X1 U18377 ( .B1(n16414), .B2(n21789), .A(n16317), .ZN(P1_U2969) );
  NOR2_X1 U18378 ( .A1(n16319), .A2(n16318), .ZN(n16321) );
  XOR2_X1 U18379 ( .A(n16321), .B(n16320), .Z(n16423) );
  NOR2_X1 U18380 ( .A1(n21600), .A2(n20089), .ZN(n16417) );
  AOI21_X1 U18381 ( .B1(n20192), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n16417), .ZN(n16322) );
  OAI21_X1 U18382 ( .B1(n20200), .B2(n16323), .A(n16322), .ZN(n16324) );
  AOI21_X1 U18383 ( .B1(n16325), .B2(n20186), .A(n16324), .ZN(n16326) );
  OAI21_X1 U18384 ( .B1(n16423), .B2(n21789), .A(n16326), .ZN(P1_U2970) );
  XNOR2_X1 U18385 ( .A(n20182), .B(n21580), .ZN(n16327) );
  XNOR2_X1 U18386 ( .A(n16302), .B(n16327), .ZN(n21574) );
  AOI22_X1 U18387 ( .A1(n20192), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B1(
        n16504), .B2(P1_REIP_REG_27__SCAN_IN), .ZN(n16328) );
  OAI21_X1 U18388 ( .B1(n20200), .B2(n16329), .A(n16328), .ZN(n16330) );
  AOI21_X1 U18389 ( .B1(n16331), .B2(n20186), .A(n16330), .ZN(n16332) );
  OAI21_X1 U18390 ( .B1(n21789), .B2(n21574), .A(n16332), .ZN(P1_U2972) );
  NAND3_X1 U18391 ( .A1(n16334), .A2(n16343), .A3(n16333), .ZN(n16335) );
  XNOR2_X1 U18392 ( .A(n16335), .B(n16432), .ZN(n16441) );
  NAND2_X1 U18393 ( .A1(n21585), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n16437) );
  OAI21_X1 U18394 ( .B1(n20155), .B2(n16336), .A(n16437), .ZN(n16339) );
  NOR2_X1 U18395 ( .A1(n16337), .A2(n20194), .ZN(n16338) );
  AOI211_X1 U18396 ( .C1(n20172), .C2(n16340), .A(n16339), .B(n16338), .ZN(
        n16341) );
  OAI21_X1 U18397 ( .B1(n21789), .B2(n16441), .A(n16341), .ZN(P1_U2973) );
  OAI21_X1 U18398 ( .B1(n11000), .B2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n16342), .ZN(n16344) );
  OAI211_X1 U18399 ( .C1(n21603), .C2(n20182), .A(n16344), .B(n16343), .ZN(
        n16345) );
  XNOR2_X1 U18400 ( .A(n16345), .B(n16433), .ZN(n21587) );
  AOI22_X1 U18401 ( .A1(n20192), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B1(
        n16504), .B2(P1_REIP_REG_25__SCAN_IN), .ZN(n16346) );
  OAI21_X1 U18402 ( .B1(n20200), .B2(n16347), .A(n16346), .ZN(n16348) );
  AOI21_X1 U18403 ( .B1(n16349), .B2(n20186), .A(n16348), .ZN(n16350) );
  OAI21_X1 U18404 ( .B1(n21789), .B2(n21587), .A(n16350), .ZN(P1_U2974) );
  OR2_X1 U18405 ( .A1(n20182), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16352) );
  NAND3_X1 U18406 ( .A1(n11000), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n20182), .ZN(n16351) );
  OAI21_X1 U18407 ( .B1(n11000), .B2(n16352), .A(n16351), .ZN(n16353) );
  XNOR2_X1 U18408 ( .A(n16353), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16449) );
  NAND2_X1 U18409 ( .A1(n21585), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n16444) );
  OAI21_X1 U18410 ( .B1(n20155), .B2(n21775), .A(n16444), .ZN(n16355) );
  NOR2_X1 U18411 ( .A1(n21778), .A2(n20194), .ZN(n16354) );
  AOI211_X1 U18412 ( .C1(n20172), .C2(n21781), .A(n16355), .B(n16354), .ZN(
        n16356) );
  OAI21_X1 U18413 ( .B1(n16449), .B2(n21789), .A(n16356), .ZN(P1_U2975) );
  NAND2_X1 U18414 ( .A1(n16358), .A2(n16357), .ZN(n16359) );
  XOR2_X1 U18415 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n16359), .Z(
        n16464) );
  INV_X1 U18416 ( .A(n16360), .ZN(n16362) );
  AOI22_X1 U18417 ( .A1(n20192), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n16504), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n16361) );
  OAI21_X1 U18418 ( .B1(n20200), .B2(n16362), .A(n16361), .ZN(n16363) );
  AOI21_X1 U18419 ( .B1(n16364), .B2(n20186), .A(n16363), .ZN(n16365) );
  OAI21_X1 U18420 ( .B1(n21789), .B2(n16464), .A(n16365), .ZN(P1_U2977) );
  MUX2_X1 U18421 ( .A(n16367), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .S(
        n12866), .Z(n16374) );
  NAND2_X1 U18422 ( .A1(n16366), .A2(n16374), .ZN(n16373) );
  OAI21_X1 U18423 ( .B1(n16367), .B2(n20182), .A(n16373), .ZN(n16479) );
  AOI22_X1 U18424 ( .A1(n16479), .A2(n16484), .B1(n20182), .B2(n16373), .ZN(
        n20181) );
  OAI21_X1 U18425 ( .B1(n20182), .B2(n16484), .A(n20181), .ZN(n16368) );
  XNOR2_X1 U18426 ( .A(n16368), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16465) );
  NAND2_X1 U18427 ( .A1(n16465), .A2(n20188), .ZN(n16372) );
  NOR2_X1 U18428 ( .A1(n21600), .A2(n20074), .ZN(n16472) );
  INV_X1 U18429 ( .A(n21768), .ZN(n16369) );
  NOR2_X1 U18430 ( .A1(n20200), .A2(n16369), .ZN(n16370) );
  AOI211_X1 U18431 ( .C1(n20192), .C2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16472), .B(n16370), .ZN(n16371) );
  OAI211_X1 U18432 ( .C1(n20194), .C2(n21765), .A(n16372), .B(n16371), .ZN(
        P1_U2979) );
  OAI21_X1 U18433 ( .B1(n16366), .B2(n16374), .A(n16373), .ZN(n16498) );
  INV_X1 U18434 ( .A(n16375), .ZN(n16377) );
  NAND2_X1 U18435 ( .A1(n16504), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n16494) );
  NAND2_X1 U18436 ( .A1(n20192), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16376) );
  OAI211_X1 U18437 ( .C1(n20200), .C2(n16377), .A(n16494), .B(n16376), .ZN(
        n16378) );
  AOI21_X1 U18438 ( .B1(n16379), .B2(n20186), .A(n16378), .ZN(n16380) );
  OAI21_X1 U18439 ( .B1(n21789), .B2(n16498), .A(n16380), .ZN(P1_U2981) );
  OAI21_X1 U18440 ( .B1(n16382), .B2(n21565), .A(n16501), .ZN(n16384) );
  OAI21_X1 U18441 ( .B1(n20182), .B2(n16522), .A(n16510), .ZN(n16502) );
  OAI21_X1 U18442 ( .B1(n16382), .B2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n16502), .ZN(n16383) );
  XOR2_X1 U18443 ( .A(n16384), .B(n16383), .Z(n21554) );
  INV_X1 U18444 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n16385) );
  OAI22_X1 U18445 ( .A1(n20155), .A2(n16386), .B1(n21600), .B2(n16385), .ZN(
        n16388) );
  NOR2_X1 U18446 ( .A1(n21735), .A2(n20194), .ZN(n16387) );
  AOI211_X1 U18447 ( .C1(n20172), .C2(n21732), .A(n16388), .B(n16387), .ZN(
        n16389) );
  OAI21_X1 U18448 ( .B1(n21554), .B2(n21789), .A(n16389), .ZN(P1_U2983) );
  INV_X1 U18449 ( .A(n16390), .ZN(n16396) );
  INV_X1 U18450 ( .A(n15887), .ZN(n16393) );
  OAI22_X1 U18451 ( .A1(n16393), .A2(n16392), .B1(n16391), .B2(n20182), .ZN(
        n16545) );
  INV_X1 U18452 ( .A(n16398), .ZN(n16394) );
  OAI21_X1 U18453 ( .B1(n20182), .B2(n16551), .A(n16394), .ZN(n16544) );
  NOR2_X1 U18454 ( .A1(n16545), .A2(n16544), .ZN(n16543) );
  MUX2_X1 U18455 ( .A(n16396), .B(n16395), .S(n16543), .Z(n16397) );
  AOI21_X1 U18456 ( .B1(n16398), .B2(n21521), .A(n16397), .ZN(n16541) );
  NAND2_X1 U18457 ( .A1(n16541), .A2(n20188), .ZN(n16402) );
  NAND2_X1 U18458 ( .A1(n16504), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n16536) );
  OAI21_X1 U18459 ( .B1(n20155), .B2(n15914), .A(n16536), .ZN(n16399) );
  AOI21_X1 U18460 ( .B1(n20172), .B2(n16400), .A(n16399), .ZN(n16401) );
  OAI211_X1 U18461 ( .C1(n20194), .C2(n16403), .A(n16402), .B(n16401), .ZN(
        P1_U2986) );
  INV_X1 U18462 ( .A(n16404), .ZN(n16409) );
  INV_X1 U18463 ( .A(n16424), .ZN(n16420) );
  OAI21_X1 U18464 ( .B1(n16420), .B2(n16451), .A(n16405), .ZN(n16418) );
  OAI21_X1 U18465 ( .B1(n16418), .B2(n16406), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16408) );
  OAI211_X1 U18466 ( .C1(n16410), .C2(n16409), .A(n16408), .B(n16407), .ZN(
        n16411) );
  AOI21_X1 U18467 ( .B1(n16412), .B2(n21595), .A(n16411), .ZN(n16413) );
  OAI21_X1 U18468 ( .B1(n16414), .B2(n16575), .A(n16413), .ZN(P1_U3001) );
  NOR2_X1 U18469 ( .A1(n16415), .A2(n21560), .ZN(n16416) );
  AOI211_X1 U18470 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16418), .A(
        n16417), .B(n16416), .ZN(n16422) );
  NAND3_X1 U18471 ( .A1(n21581), .A2(n16420), .A3(n16419), .ZN(n16421) );
  OAI211_X1 U18472 ( .C1(n16423), .C2(n16575), .A(n16422), .B(n16421), .ZN(
        P1_U3002) );
  AND3_X1 U18473 ( .A1(n21581), .A2(n16425), .A3(n16424), .ZN(n16429) );
  OAI21_X1 U18474 ( .B1(n16427), .B2(n21560), .A(n16426), .ZN(n16428) );
  AOI211_X1 U18475 ( .C1(n21582), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16429), .B(n16428), .ZN(n16430) );
  OAI21_X1 U18476 ( .B1(n16431), .B2(n16575), .A(n16430), .ZN(P1_U3003) );
  AOI21_X1 U18477 ( .B1(n16433), .B2(n16432), .A(n21592), .ZN(n16434) );
  NAND2_X1 U18478 ( .A1(n16435), .A2(n16434), .ZN(n16436) );
  OAI211_X1 U18479 ( .C1(n16438), .C2(n21560), .A(n16437), .B(n16436), .ZN(
        n16439) );
  AOI21_X1 U18480 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n21586), .A(
        n16439), .ZN(n16440) );
  OAI21_X1 U18481 ( .B1(n16441), .B2(n16575), .A(n16440), .ZN(P1_U3005) );
  NOR2_X1 U18482 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n21603), .ZN(
        n16447) );
  OAI21_X1 U18483 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n16442), .A(
        n21598), .ZN(n16443) );
  NAND2_X1 U18484 ( .A1(n16443), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16445) );
  OAI211_X1 U18485 ( .C1(n21560), .C2(n21787), .A(n16445), .B(n16444), .ZN(
        n16446) );
  AOI21_X1 U18486 ( .B1(n21602), .B2(n16447), .A(n16446), .ZN(n16448) );
  OAI21_X1 U18487 ( .B1(n16449), .B2(n16575), .A(n16448), .ZN(P1_U3007) );
  INV_X1 U18488 ( .A(n16467), .ZN(n16450) );
  NAND2_X1 U18489 ( .A1(n21544), .A2(n16450), .ZN(n16533) );
  OAI211_X1 U18490 ( .C1(n21531), .C2(n16527), .A(n21530), .B(n16533), .ZN(
        n16511) );
  AOI21_X1 U18491 ( .B1(n16513), .B2(n16455), .A(n16511), .ZN(n16480) );
  NOR2_X1 U18492 ( .A1(n20183), .A2(n16484), .ZN(n16452) );
  AOI21_X1 U18493 ( .B1(n16480), .B2(n16452), .A(n16451), .ZN(n21567) );
  NAND2_X1 U18494 ( .A1(n16548), .A2(n21533), .ZN(n16549) );
  OAI21_X1 U18495 ( .B1(n16546), .B2(n16453), .A(n16549), .ZN(n16561) );
  NAND2_X1 U18496 ( .A1(n16454), .A2(n16561), .ZN(n21520) );
  NOR2_X1 U18497 ( .A1(n16455), .A2(n21520), .ZN(n16485) );
  NAND4_X1 U18498 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(n16485), .A4(n16456), .ZN(
        n21570) );
  INV_X1 U18499 ( .A(n21570), .ZN(n16457) );
  OAI21_X1 U18500 ( .B1(n21567), .B2(n16457), .A(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16463) );
  INV_X1 U18501 ( .A(n16489), .ZN(n16491) );
  NOR4_X1 U18502 ( .A1(n21520), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n16458), .A4(n16491), .ZN(n16461) );
  OAI22_X1 U18503 ( .A1(n16459), .A2(n21560), .B1(n20078), .B2(n21600), .ZN(
        n16460) );
  NOR2_X1 U18504 ( .A1(n16461), .A2(n16460), .ZN(n16462) );
  OAI211_X1 U18505 ( .C1(n16464), .C2(n16575), .A(n16463), .B(n16462), .ZN(
        P1_U3009) );
  INV_X1 U18506 ( .A(n16465), .ZN(n16477) );
  INV_X1 U18507 ( .A(n16466), .ZN(n16532) );
  NOR2_X1 U18508 ( .A1(n16591), .A2(n16525), .ZN(n16530) );
  AOI22_X1 U18509 ( .A1(n21544), .A2(n16467), .B1(n16532), .B2(n16530), .ZN(
        n21522) );
  INV_X1 U18510 ( .A(n21522), .ZN(n16469) );
  OAI21_X1 U18511 ( .B1(n16469), .B2(n16468), .A(n16484), .ZN(n16470) );
  AOI21_X1 U18512 ( .B1(n16480), .B2(n16470), .A(n20183), .ZN(n16471) );
  AOI211_X1 U18513 ( .C1(n21595), .C2(n16473), .A(n16472), .B(n16471), .ZN(
        n16476) );
  NOR2_X1 U18514 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n16484), .ZN(
        n16474) );
  NAND2_X1 U18515 ( .A1(n16485), .A2(n16474), .ZN(n16475) );
  OAI211_X1 U18516 ( .C1(n16477), .C2(n16575), .A(n16476), .B(n16475), .ZN(
        P1_U3011) );
  XNOR2_X1 U18517 ( .A(n12866), .B(n16484), .ZN(n16478) );
  XNOR2_X1 U18518 ( .A(n16479), .B(n16478), .ZN(n20177) );
  INV_X1 U18519 ( .A(n20177), .ZN(n16487) );
  INV_X1 U18520 ( .A(n16480), .ZN(n16481) );
  AOI22_X1 U18521 ( .A1(n21585), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n16481), .ZN(n16482) );
  OAI21_X1 U18522 ( .B1(n21751), .B2(n21560), .A(n16482), .ZN(n16483) );
  AOI21_X1 U18523 ( .B1(n16485), .B2(n16484), .A(n16483), .ZN(n16486) );
  OAI21_X1 U18524 ( .B1(n16487), .B2(n16575), .A(n16486), .ZN(P1_U3012) );
  INV_X1 U18525 ( .A(n16511), .ZN(n16488) );
  OAI21_X1 U18526 ( .B1(n16490), .B2(n16489), .A(n16488), .ZN(n16505) );
  NOR2_X1 U18527 ( .A1(n16491), .A2(n21520), .ZN(n16492) );
  NAND2_X1 U18528 ( .A1(n16367), .A2(n16492), .ZN(n16493) );
  OAI211_X1 U18529 ( .C1(n16495), .C2(n21560), .A(n16494), .B(n16493), .ZN(
        n16496) );
  AOI21_X1 U18530 ( .B1(n16505), .B2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n16496), .ZN(n16497) );
  OAI21_X1 U18531 ( .B1(n16498), .B2(n16575), .A(n16497), .ZN(P1_U3013) );
  INV_X1 U18532 ( .A(n16510), .ZN(n16499) );
  NAND3_X1 U18533 ( .A1(n16499), .A2(n21555), .A3(n12866), .ZN(n16500) );
  OAI21_X1 U18534 ( .B1(n16502), .B2(n16501), .A(n16500), .ZN(n16503) );
  XNOR2_X1 U18535 ( .A(n16503), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n20176) );
  AOI22_X1 U18536 ( .A1(n21595), .A2(n20123), .B1(n16504), .B2(
        P1_REIP_REG_17__SCAN_IN), .ZN(n16508) );
  NOR2_X1 U18537 ( .A1(n16512), .A2(n21520), .ZN(n21558) );
  AND2_X1 U18538 ( .A1(n21558), .A2(n21555), .ZN(n16506) );
  OAI21_X1 U18539 ( .B1(n16506), .B2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n16505), .ZN(n16507) );
  OAI211_X1 U18540 ( .C1(n20176), .C2(n16575), .A(n16508), .B(n16507), .ZN(
        P1_U3014) );
  XNOR2_X1 U18541 ( .A(n12866), .B(n16522), .ZN(n16509) );
  XNOR2_X1 U18542 ( .A(n16510), .B(n16509), .ZN(n20170) );
  AOI21_X1 U18543 ( .B1(n16513), .B2(n16512), .A(n16511), .ZN(n21566) );
  INV_X1 U18544 ( .A(n21566), .ZN(n16521) );
  INV_X1 U18545 ( .A(n16514), .ZN(n16516) );
  NOR2_X1 U18546 ( .A1(n16516), .A2(n16515), .ZN(n16519) );
  OAI21_X1 U18547 ( .B1(n16519), .B2(n16518), .A(n16517), .ZN(n20126) );
  OAI22_X1 U18548 ( .A1(n21560), .A2(n20126), .B1(n21600), .B2(n20067), .ZN(
        n16520) );
  AOI21_X1 U18549 ( .B1(n16521), .B2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n16520), .ZN(n16524) );
  NAND2_X1 U18550 ( .A1(n21558), .A2(n16522), .ZN(n16523) );
  OAI211_X1 U18551 ( .C1(n20170), .C2(n16575), .A(n16524), .B(n16523), .ZN(
        P1_U3016) );
  AOI221_X1 U18552 ( .B1(n16525), .B2(n21522), .C1(n16526), .C2(n21522), .A(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16540) );
  AOI21_X1 U18553 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16527), .A(
        n16526), .ZN(n16528) );
  NOR2_X1 U18554 ( .A1(n16529), .A2(n16528), .ZN(n16535) );
  INV_X1 U18555 ( .A(n16530), .ZN(n16531) );
  NAND2_X1 U18556 ( .A1(n16532), .A2(n16531), .ZN(n16534) );
  NAND3_X1 U18557 ( .A1(n16535), .A2(n16534), .A3(n16533), .ZN(n21523) );
  NAND2_X1 U18558 ( .A1(n21523), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16537) );
  OAI211_X1 U18559 ( .C1(n21560), .C2(n16538), .A(n16537), .B(n16536), .ZN(
        n16539) );
  AOI211_X1 U18560 ( .C1(n16541), .C2(n21596), .A(n16540), .B(n16539), .ZN(
        n16542) );
  INV_X1 U18561 ( .A(n16542), .ZN(P1_U3018) );
  AOI21_X1 U18562 ( .B1(n16545), .B2(n16544), .A(n16543), .ZN(n20167) );
  OAI21_X1 U18563 ( .B1(n16560), .B2(n16546), .A(n21544), .ZN(n16547) );
  OAI211_X1 U18564 ( .C1(n21531), .C2(n16548), .A(n21530), .B(n16547), .ZN(
        n16562) );
  INV_X1 U18565 ( .A(n16562), .ZN(n16550) );
  AOI221_X1 U18566 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16550), 
        .C1(n16549), .C2(n16550), .A(n16551), .ZN(n16555) );
  INV_X1 U18567 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n21709) );
  NAND3_X1 U18568 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16551), .A3(
        n16561), .ZN(n16553) );
  NAND2_X1 U18569 ( .A1(n21595), .A2(n21703), .ZN(n16552) );
  OAI211_X1 U18570 ( .C1(n21709), .C2(n21600), .A(n16553), .B(n16552), .ZN(
        n16554) );
  NOR2_X1 U18571 ( .A1(n16555), .A2(n16554), .ZN(n16556) );
  OAI21_X1 U18572 ( .B1(n20167), .B2(n16575), .A(n16556), .ZN(P1_U3019) );
  MUX2_X1 U18573 ( .A(n15887), .B(n16557), .S(n20182), .Z(n16565) );
  NOR2_X2 U18574 ( .A1(n16565), .A2(n13089), .ZN(n16566) );
  NOR2_X1 U18575 ( .A1(n16566), .A2(n15887), .ZN(n16558) );
  AOI22_X1 U18576 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16562), .B1(
        n16561), .B2(n16560), .ZN(n16564) );
  NOR2_X1 U18577 ( .A1(n21600), .A2(n21696), .ZN(n20162) );
  AOI21_X1 U18578 ( .B1(n21595), .B2(n21693), .A(n20162), .ZN(n16563) );
  OAI211_X1 U18579 ( .C1(n20160), .C2(n16575), .A(n16564), .B(n16563), .ZN(
        P1_U3020) );
  INV_X1 U18580 ( .A(n16565), .ZN(n16568) );
  INV_X1 U18581 ( .A(n16566), .ZN(n16567) );
  OAI21_X1 U18582 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16568), .A(
        n16567), .ZN(n20159) );
  XNOR2_X1 U18583 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n16569), .ZN(
        n16570) );
  AOI22_X1 U18584 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n16572), .B1(
        n16571), .B2(n16570), .ZN(n16574) );
  AOI22_X1 U18585 ( .A1(n21595), .A2(n21685), .B1(n21585), .B2(
        P1_REIP_REG_10__SCAN_IN), .ZN(n16573) );
  OAI211_X1 U18586 ( .C1(n20159), .C2(n16575), .A(n16574), .B(n16573), .ZN(
        P1_U3021) );
  OAI211_X1 U18587 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n15087), .A(n22111), 
        .B(n22059), .ZN(n16576) );
  OAI21_X1 U18588 ( .B1(n16577), .B2(n11019), .A(n16576), .ZN(n16578) );
  MUX2_X1 U18589 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n16578), .S(
        n17384), .Z(P1_U3477) );
  AOI21_X1 U18590 ( .B1(n16580), .B2(n22015), .A(n16579), .ZN(n16581) );
  OAI21_X1 U18591 ( .B1(n16583), .B2(n16582), .A(n16581), .ZN(n16584) );
  MUX2_X1 U18592 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n16584), .S(
        n17384), .Z(P1_U3475) );
  NOR3_X1 U18593 ( .A1(n16585), .A2(n15211), .A3(n15213), .ZN(n16588) );
  NOR2_X1 U18594 ( .A1(n11019), .A2(n16586), .ZN(n16587) );
  AOI211_X1 U18595 ( .C1(n17352), .C2(n12883), .A(n16588), .B(n16587), .ZN(
        n17358) );
  AOI22_X1 U18596 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n16590), .B2(n16589), .ZN(
        n16598) );
  INV_X1 U18597 ( .A(n16598), .ZN(n16593) );
  NOR2_X1 U18598 ( .A1(n21798), .A2(n16591), .ZN(n16597) );
  NOR3_X1 U18599 ( .A1(n15211), .A2(n15213), .A3(n21792), .ZN(n16592) );
  AOI21_X1 U18600 ( .B1(n16593), .B2(n16597), .A(n16592), .ZN(n16594) );
  OAI21_X1 U18601 ( .B1(n17358), .B2(n21794), .A(n16594), .ZN(n16595) );
  MUX2_X1 U18602 ( .A(n16595), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n21796), .Z(P1_U3473) );
  AOI22_X1 U18603 ( .A1(n16598), .A2(n16597), .B1(n16596), .B2(n21807), .ZN(
        n16599) );
  OAI21_X1 U18604 ( .B1(n16600), .B2(n21794), .A(n16599), .ZN(n16601) );
  MUX2_X1 U18605 ( .A(n16601), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n21796), .Z(P1_U3472) );
  NAND2_X1 U18606 ( .A1(n16602), .A2(n18752), .ZN(n16604) );
  XNOR2_X1 U18607 ( .A(n16604), .B(n16603), .ZN(n16605) );
  NAND2_X1 U18608 ( .A1(n16605), .A2(n18861), .ZN(n16610) );
  AOI22_X1 U18609 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n18851), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n18850), .ZN(n16607) );
  NAND2_X1 U18610 ( .A1(n18852), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n16606) );
  OAI211_X1 U18611 ( .C1(n16722), .C2(n18855), .A(n16607), .B(n16606), .ZN(
        n16608) );
  AOI21_X1 U18612 ( .B1(n16652), .B2(n18811), .A(n16608), .ZN(n16609) );
  OAI211_X1 U18613 ( .C1(n18803), .C2(n16611), .A(n16610), .B(n16609), .ZN(
        P2_U2828) );
  AOI21_X1 U18614 ( .B1(n16614), .B2(n16613), .A(n16612), .ZN(n16615) );
  NAND2_X1 U18615 ( .A1(n16615), .A2(n18861), .ZN(n16628) );
  OR2_X1 U18616 ( .A1(n16616), .A2(n16617), .ZN(n16618) );
  NAND2_X1 U18617 ( .A1(n11909), .A2(n16618), .ZN(n17050) );
  INV_X1 U18618 ( .A(n17050), .ZN(n16626) );
  AOI22_X1 U18619 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18851), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n18850), .ZN(n16623) );
  INV_X1 U18620 ( .A(n16620), .ZN(n16621) );
  XNOR2_X1 U18621 ( .A(n16619), .B(n16621), .ZN(n19584) );
  NAND2_X1 U18622 ( .A1(n18763), .A2(n19584), .ZN(n16622) );
  OAI211_X1 U18623 ( .C1(n18733), .C2(n16624), .A(n16623), .B(n16622), .ZN(
        n16625) );
  AOI21_X1 U18624 ( .B1(n16626), .B2(n18811), .A(n16625), .ZN(n16627) );
  OAI211_X1 U18625 ( .C1(n18803), .C2(n16629), .A(n16628), .B(n16627), .ZN(
        P2_U2833) );
  MUX2_X1 U18626 ( .A(P2_EBX_REG_31__SCAN_IN), .B(n16630), .S(n16651), .Z(
        P2_U2856) );
  OR2_X1 U18627 ( .A1(n16635), .A2(n16634), .ZN(n16636) );
  NAND2_X1 U18628 ( .A1(n13675), .A2(n16636), .ZN(n18858) );
  NOR2_X1 U18629 ( .A1(n18858), .A2(n16689), .ZN(n16637) );
  AOI21_X1 U18630 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(n16689), .A(n16637), .ZN(
        n16638) );
  OAI21_X1 U18631 ( .B1(n16712), .B2(n16698), .A(n16638), .ZN(P2_U2858) );
  INV_X1 U18632 ( .A(n16640), .ZN(n16641) );
  NOR2_X1 U18633 ( .A1(n16646), .A2(n16641), .ZN(n16643) );
  XNOR2_X1 U18634 ( .A(n16643), .B(n16642), .ZN(n16719) );
  NOR2_X1 U18635 ( .A1(n18841), .A2(n16689), .ZN(n16644) );
  AOI21_X1 U18636 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n16689), .A(n16644), .ZN(
        n16645) );
  OAI21_X1 U18637 ( .B1(n16719), .B2(n16698), .A(n16645), .ZN(P2_U2859) );
  INV_X1 U18638 ( .A(n16646), .ZN(n16648) );
  NAND2_X1 U18639 ( .A1(n16648), .A2(n16647), .ZN(n16649) );
  XOR2_X1 U18640 ( .A(n16650), .B(n16649), .Z(n16725) );
  NAND2_X1 U18641 ( .A1(n16689), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n16654) );
  NAND2_X1 U18642 ( .A1(n16652), .A2(n16651), .ZN(n16653) );
  OAI211_X1 U18643 ( .C1(n16725), .C2(n16698), .A(n16654), .B(n16653), .ZN(
        P2_U2860) );
  OR2_X1 U18644 ( .A1(n16655), .A2(n16656), .ZN(n16657) );
  NAND2_X1 U18645 ( .A1(n14500), .A2(n16657), .ZN(n18830) );
  AOI21_X1 U18646 ( .B1(n16660), .B2(n16659), .A(n16658), .ZN(n16726) );
  NAND2_X1 U18647 ( .A1(n16726), .A2(n16686), .ZN(n16662) );
  NAND2_X1 U18648 ( .A1(n16689), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n16661) );
  OAI211_X1 U18649 ( .C1(n18830), .C2(n16689), .A(n16662), .B(n16661), .ZN(
        P2_U2861) );
  OAI21_X1 U18650 ( .B1(n16665), .B2(n16664), .A(n16663), .ZN(n16745) );
  NOR2_X1 U18651 ( .A1(n16672), .A2(n16666), .ZN(n16667) );
  OR2_X1 U18652 ( .A1(n16655), .A2(n16667), .ZN(n18818) );
  NOR2_X1 U18653 ( .A1(n18818), .A2(n16689), .ZN(n16668) );
  AOI21_X1 U18654 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n16689), .A(n16668), .ZN(
        n16669) );
  OAI21_X1 U18655 ( .B1(n16745), .B2(n16698), .A(n16669), .ZN(P2_U2862) );
  AND2_X1 U18656 ( .A1(n16671), .A2(n16670), .ZN(n16673) );
  OR2_X1 U18657 ( .A1(n16673), .A2(n16672), .ZN(n16821) );
  AOI21_X1 U18658 ( .B1(n16676), .B2(n16675), .A(n16674), .ZN(n16746) );
  NAND2_X1 U18659 ( .A1(n16746), .A2(n16686), .ZN(n16678) );
  NAND2_X1 U18660 ( .A1(n16689), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n16677) );
  OAI211_X1 U18661 ( .C1(n16821), .C2(n16689), .A(n16678), .B(n16677), .ZN(
        P2_U2863) );
  XNOR2_X1 U18662 ( .A(n16684), .B(n16680), .ZN(n16761) );
  NOR2_X1 U18663 ( .A1(n18792), .A2(n16689), .ZN(n16681) );
  AOI21_X1 U18664 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n16689), .A(n16681), .ZN(
        n16682) );
  OAI21_X1 U18665 ( .B1(n16761), .B2(n16698), .A(n16682), .ZN(P2_U2864) );
  AOI21_X1 U18666 ( .B1(n16685), .B2(n16683), .A(n16684), .ZN(n19587) );
  NAND2_X1 U18667 ( .A1(n19587), .A2(n16686), .ZN(n16688) );
  NAND2_X1 U18668 ( .A1(n16689), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n16687) );
  OAI211_X1 U18669 ( .C1(n17050), .C2(n16689), .A(n16688), .B(n16687), .ZN(
        P2_U2865) );
  OAI21_X1 U18670 ( .B1(n16691), .B2(n16690), .A(n16683), .ZN(n16772) );
  INV_X1 U18671 ( .A(n16616), .ZN(n16695) );
  NAND2_X1 U18672 ( .A1(n16693), .A2(n16692), .ZN(n16694) );
  NAND2_X1 U18673 ( .A1(n16695), .A2(n16694), .ZN(n18779) );
  NOR2_X1 U18674 ( .A1(n18779), .A2(n16689), .ZN(n16696) );
  AOI21_X1 U18675 ( .B1(P2_EBX_REG_21__SCAN_IN), .B2(n16689), .A(n16696), .ZN(
        n16697) );
  OAI21_X1 U18676 ( .B1(n16772), .B2(n16698), .A(n16697), .ZN(P2_U2866) );
  INV_X1 U18677 ( .A(n19582), .ZN(n16742) );
  NAND2_X1 U18678 ( .A1(n16044), .A2(n19585), .ZN(n16700) );
  AOI22_X1 U18679 ( .A1(n19583), .A2(BUF2_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19579), .ZN(n16699) );
  OAI211_X1 U18680 ( .C1(n20270), .C2(n16742), .A(n16700), .B(n16699), .ZN(
        P2_U2888) );
  AND2_X1 U18681 ( .A1(n11046), .A2(n16701), .ZN(n16703) );
  OR2_X1 U18682 ( .A1(n19374), .A2(n16704), .ZN(n16707) );
  NAND2_X1 U18683 ( .A1(n19581), .A2(n16705), .ZN(n16706) );
  OAI211_X1 U18684 ( .C1(n18856), .C2(n16765), .A(n16707), .B(n16706), .ZN(
        n16709) );
  AND2_X1 U18685 ( .A1(n19582), .A2(BUF1_REG_29__SCAN_IN), .ZN(n16708) );
  NOR2_X1 U18686 ( .A1(n16709), .A2(n16708), .ZN(n16711) );
  NAND2_X1 U18687 ( .A1(n19583), .A2(BUF2_REG_29__SCAN_IN), .ZN(n16710) );
  OAI211_X1 U18688 ( .C1(n16712), .C2(n16771), .A(n16711), .B(n16710), .ZN(
        P2_U2890) );
  NAND2_X1 U18689 ( .A1(n18839), .A2(n19585), .ZN(n16716) );
  AOI22_X1 U18690 ( .A1(n19581), .A2(n16713), .B1(n19579), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n16715) );
  NAND2_X1 U18691 ( .A1(n19582), .A2(BUF1_REG_28__SCAN_IN), .ZN(n16714) );
  NAND3_X1 U18692 ( .A1(n16716), .A2(n16715), .A3(n16714), .ZN(n16717) );
  AOI21_X1 U18693 ( .B1(n19583), .B2(BUF2_REG_28__SCAN_IN), .A(n16717), .ZN(
        n16718) );
  OAI21_X1 U18694 ( .B1(n16719), .B2(n16771), .A(n16718), .ZN(P2_U2891) );
  NAND2_X1 U18695 ( .A1(n19582), .A2(BUF1_REG_27__SCAN_IN), .ZN(n16721) );
  AOI22_X1 U18696 ( .A1(n19581), .A2(n19364), .B1(n19579), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n16720) );
  OAI211_X1 U18697 ( .C1(n16722), .C2(n16765), .A(n16721), .B(n16720), .ZN(
        n16723) );
  AOI21_X1 U18698 ( .B1(n19583), .B2(BUF2_REG_27__SCAN_IN), .A(n16723), .ZN(
        n16724) );
  OAI21_X1 U18699 ( .B1(n16725), .B2(n16771), .A(n16724), .ZN(P2_U2892) );
  INV_X1 U18700 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n16736) );
  NAND2_X1 U18701 ( .A1(n16726), .A2(n19586), .ZN(n16735) );
  NOR2_X1 U18702 ( .A1(n16766), .A2(n16727), .ZN(n16733) );
  NOR2_X1 U18703 ( .A1(n16728), .A2(n16729), .ZN(n16730) );
  OR2_X1 U18704 ( .A1(n14511), .A2(n16730), .ZN(n18829) );
  OAI22_X1 U18705 ( .A1(n18829), .A2(n16765), .B1(n19374), .B2(n16731), .ZN(
        n16732) );
  AOI211_X1 U18706 ( .C1(BUF1_REG_26__SCAN_IN), .C2(n19582), .A(n16733), .B(
        n16732), .ZN(n16734) );
  OAI211_X1 U18707 ( .C1(n16755), .C2(n16736), .A(n16735), .B(n16734), .ZN(
        P2_U2893) );
  AND2_X1 U18708 ( .A1(n16737), .A2(n16738), .ZN(n16739) );
  NOR2_X1 U18709 ( .A1(n16728), .A2(n16739), .ZN(n18816) );
  AOI22_X1 U18710 ( .A1(n18816), .A2(n19585), .B1(P2_EAX_REG_25__SCAN_IN), 
        .B2(n19579), .ZN(n16741) );
  NAND2_X1 U18711 ( .A1(n19581), .A2(n19368), .ZN(n16740) );
  OAI211_X1 U18712 ( .C1(n16742), .C2(n20257), .A(n16741), .B(n16740), .ZN(
        n16743) );
  AOI21_X1 U18713 ( .B1(n19583), .B2(BUF2_REG_25__SCAN_IN), .A(n16743), .ZN(
        n16744) );
  OAI21_X1 U18714 ( .B1(n16745), .B2(n16771), .A(n16744), .ZN(P2_U2894) );
  INV_X1 U18715 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n16754) );
  NAND2_X1 U18716 ( .A1(n16746), .A2(n19586), .ZN(n16753) );
  INV_X1 U18717 ( .A(n12415), .ZN(n16747) );
  OAI21_X1 U18718 ( .B1(n16747), .B2(n11246), .A(n16737), .ZN(n18814) );
  OAI22_X1 U18719 ( .A1(n16765), .A2(n18814), .B1(n19374), .B2(n16748), .ZN(
        n16751) );
  NOR2_X1 U18720 ( .A1(n16766), .A2(n16749), .ZN(n16750) );
  AOI211_X1 U18721 ( .C1(BUF1_REG_24__SCAN_IN), .C2(n19582), .A(n16751), .B(
        n16750), .ZN(n16752) );
  OAI211_X1 U18722 ( .C1(n16755), .C2(n16754), .A(n16753), .B(n16752), .ZN(
        P2_U2895) );
  OAI22_X1 U18723 ( .A1(n16765), .A2(n18791), .B1(n19374), .B2(n16756), .ZN(
        n16758) );
  NOR2_X1 U18724 ( .A1(n16766), .A2(n19378), .ZN(n16757) );
  AOI211_X1 U18725 ( .C1(BUF1_REG_23__SCAN_IN), .C2(n19582), .A(n16758), .B(
        n16757), .ZN(n16760) );
  NAND2_X1 U18726 ( .A1(n19583), .A2(BUF2_REG_23__SCAN_IN), .ZN(n16759) );
  OAI211_X1 U18727 ( .C1(n16761), .C2(n16771), .A(n16760), .B(n16759), .ZN(
        P2_U2896) );
  NAND2_X1 U18728 ( .A1(n15948), .A2(n16762), .ZN(n16763) );
  AND2_X1 U18729 ( .A1(n16619), .A2(n16763), .ZN(n17057) );
  INV_X1 U18730 ( .A(n17057), .ZN(n18778) );
  OAI22_X1 U18731 ( .A1(n16765), .A2(n18778), .B1(n19374), .B2(n16764), .ZN(
        n16768) );
  NOR2_X1 U18732 ( .A1(n16766), .A2(n19631), .ZN(n16767) );
  AOI211_X1 U18733 ( .C1(BUF1_REG_21__SCAN_IN), .C2(n19582), .A(n16768), .B(
        n16767), .ZN(n16770) );
  NAND2_X1 U18734 ( .A1(n19583), .A2(BUF2_REG_21__SCAN_IN), .ZN(n16769) );
  OAI211_X1 U18735 ( .C1(n16772), .C2(n16771), .A(n16770), .B(n16769), .ZN(
        P2_U2898) );
  NOR2_X1 U18736 ( .A1(n17631), .A2(n16773), .ZN(n16774) );
  AOI211_X1 U18737 ( .C1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n17661), .A(
        n16775), .B(n16774), .ZN(n16776) );
  OAI21_X1 U18738 ( .B1(n16777), .B2(n17651), .A(n16776), .ZN(n16778) );
  OAI21_X1 U18739 ( .B1(n16781), .B2(n17670), .A(n16780), .ZN(P2_U2983) );
  NAND2_X1 U18740 ( .A1(n16783), .A2(n16782), .ZN(n16786) );
  XOR2_X1 U18741 ( .A(n16786), .B(n16785), .Z(n17014) );
  AOI21_X1 U18742 ( .B1(n17004), .B2(n16788), .A(n16787), .ZN(n17012) );
  INV_X1 U18743 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n17761) );
  NOR2_X1 U18744 ( .A1(n16970), .A2(n17761), .ZN(n17006) );
  AOI21_X1 U18745 ( .B1(n17661), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n17006), .ZN(n16791) );
  NAND2_X1 U18746 ( .A1(n17647), .A2(n16789), .ZN(n16790) );
  OAI211_X1 U18747 ( .C1(n18858), .C2(n17651), .A(n16791), .B(n16790), .ZN(
        n16792) );
  AOI21_X1 U18748 ( .B1(n17012), .B2(n17668), .A(n16792), .ZN(n16793) );
  OAI21_X1 U18749 ( .B1(n17014), .B2(n17670), .A(n16793), .ZN(P2_U2985) );
  AOI21_X1 U18750 ( .B1(n16794), .B2(n16803), .A(n16805), .ZN(n16796) );
  MUX2_X1 U18751 ( .A(n16803), .B(n16796), .S(n16795), .Z(n16797) );
  NAND2_X1 U18752 ( .A1(n16798), .A2(n16797), .ZN(n17023) );
  AOI21_X1 U18753 ( .B1(n13712), .B2(n16808), .A(n14498), .ZN(n17021) );
  NOR2_X1 U18754 ( .A1(n16970), .A2(n17758), .ZN(n17015) );
  NOR2_X1 U18755 ( .A1(n17631), .A2(n18832), .ZN(n16799) );
  AOI211_X1 U18756 ( .C1(n17661), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n17015), .B(n16799), .ZN(n16800) );
  OAI21_X1 U18757 ( .B1(n18830), .B2(n17651), .A(n16800), .ZN(n16801) );
  AOI21_X1 U18758 ( .B1(n17021), .B2(n17668), .A(n16801), .ZN(n16802) );
  OAI21_X1 U18759 ( .B1(n17023), .B2(n17670), .A(n16802), .ZN(P2_U2988) );
  INV_X1 U18760 ( .A(n16803), .ZN(n16804) );
  NOR2_X1 U18761 ( .A1(n16805), .A2(n16804), .ZN(n16806) );
  XOR2_X1 U18762 ( .A(n16806), .B(n16794), .Z(n17032) );
  AOI21_X1 U18763 ( .B1(n16807), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16810) );
  INV_X1 U18764 ( .A(n16808), .ZN(n16809) );
  NOR2_X1 U18765 ( .A1(n16810), .A2(n16809), .ZN(n17030) );
  AND2_X1 U18766 ( .A1(n12161), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n17025) );
  NOR2_X1 U18767 ( .A1(n17658), .A2(n16811), .ZN(n16812) );
  AOI211_X1 U18768 ( .C1(n18823), .C2(n17647), .A(n17025), .B(n16812), .ZN(
        n16813) );
  OAI21_X1 U18769 ( .B1(n18818), .B2(n17651), .A(n16813), .ZN(n16814) );
  AOI21_X1 U18770 ( .B1(n17030), .B2(n17668), .A(n16814), .ZN(n16815) );
  OAI21_X1 U18771 ( .B1(n17032), .B2(n17670), .A(n16815), .ZN(P2_U2989) );
  XNOR2_X1 U18772 ( .A(n13749), .B(n17036), .ZN(n17042) );
  INV_X1 U18773 ( .A(n16816), .ZN(n16818) );
  NAND2_X1 U18774 ( .A1(n16818), .A2(n16817), .ZN(n16819) );
  XNOR2_X1 U18775 ( .A(n16820), .B(n16819), .ZN(n17033) );
  NAND2_X1 U18776 ( .A1(n17033), .A2(n17617), .ZN(n16826) );
  INV_X1 U18777 ( .A(n16821), .ZN(n18810) );
  NAND2_X1 U18778 ( .A1(n12161), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n17037) );
  NAND2_X1 U18779 ( .A1(n17661), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16822) );
  OAI211_X1 U18780 ( .C1(n17631), .C2(n16823), .A(n17037), .B(n16822), .ZN(
        n16824) );
  AOI21_X1 U18781 ( .B1(n18810), .B2(n17672), .A(n16824), .ZN(n16825) );
  OAI211_X1 U18782 ( .C1(n17042), .C2(n17648), .A(n16826), .B(n16825), .ZN(
        P2_U2990) );
  OAI21_X1 U18783 ( .B1(n17658), .B2(n16828), .A(n16827), .ZN(n16829) );
  AOI21_X1 U18784 ( .B1(n17647), .B2(n18795), .A(n16829), .ZN(n16830) );
  OAI21_X1 U18785 ( .B1(n18792), .B2(n17651), .A(n16830), .ZN(n16831) );
  AOI21_X1 U18786 ( .B1(n16832), .B2(n17668), .A(n16831), .ZN(n16833) );
  OAI21_X1 U18787 ( .B1(n16834), .B2(n17670), .A(n16833), .ZN(P2_U2991) );
  INV_X1 U18788 ( .A(n16836), .ZN(n16837) );
  NOR2_X1 U18789 ( .A1(n16838), .A2(n16837), .ZN(n16839) );
  XNOR2_X1 U18790 ( .A(n16835), .B(n16839), .ZN(n17054) );
  INV_X1 U18791 ( .A(n16840), .ZN(n16842) );
  AOI21_X1 U18792 ( .B1(n16876), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16841) );
  NOR2_X1 U18793 ( .A1(n16842), .A2(n16841), .ZN(n17052) );
  INV_X1 U18794 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n17754) );
  NOR2_X1 U18795 ( .A1(n16970), .A2(n17754), .ZN(n17046) );
  NOR2_X1 U18796 ( .A1(n17631), .A2(n16843), .ZN(n16844) );
  AOI211_X1 U18797 ( .C1(n17661), .C2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n17046), .B(n16844), .ZN(n16845) );
  OAI21_X1 U18798 ( .B1(n17050), .B2(n17651), .A(n16845), .ZN(n16846) );
  AOI21_X1 U18799 ( .B1(n17052), .B2(n17668), .A(n16846), .ZN(n16847) );
  OAI21_X1 U18800 ( .B1(n17054), .B2(n17670), .A(n16847), .ZN(P2_U2992) );
  INV_X1 U18801 ( .A(n16848), .ZN(n16849) );
  NAND2_X1 U18802 ( .A1(n16850), .A2(n16849), .ZN(n16856) );
  INV_X1 U18803 ( .A(n16953), .ZN(n16852) );
  OR3_X1 U18804 ( .A1(n16942), .A2(n16852), .A3(n16851), .ZN(n16853) );
  NOR2_X1 U18805 ( .A1(n16854), .A2(n16853), .ZN(n16855) );
  NAND2_X1 U18806 ( .A1(n16856), .A2(n16855), .ZN(n16911) );
  INV_X1 U18807 ( .A(n16857), .ZN(n16910) );
  NAND2_X1 U18808 ( .A1(n16911), .A2(n16910), .ZN(n16912) );
  NAND2_X1 U18809 ( .A1(n16912), .A2(n16858), .ZN(n16903) );
  INV_X1 U18810 ( .A(n16901), .ZN(n16859) );
  NAND2_X1 U18811 ( .A1(n16860), .A2(n16859), .ZN(n16884) );
  AOI21_X1 U18812 ( .B1(n16884), .B2(n16862), .A(n16861), .ZN(n16864) );
  XNOR2_X1 U18813 ( .A(n16864), .B(n16863), .ZN(n16875) );
  AOI22_X1 U18814 ( .A1(n16875), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n12294), .B2(n16864), .ZN(n16868) );
  NAND2_X1 U18815 ( .A1(n16866), .A2(n16865), .ZN(n16867) );
  XNOR2_X1 U18816 ( .A(n16868), .B(n16867), .ZN(n17064) );
  XNOR2_X1 U18817 ( .A(n16876), .B(n17043), .ZN(n17062) );
  INV_X1 U18818 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n16869) );
  NOR2_X1 U18819 ( .A1(n16970), .A2(n16869), .ZN(n17056) );
  AOI21_X1 U18820 ( .B1(n17661), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n17056), .ZN(n16872) );
  NAND2_X1 U18821 ( .A1(n17647), .A2(n16870), .ZN(n16871) );
  OAI211_X1 U18822 ( .C1(n18779), .C2(n17651), .A(n16872), .B(n16871), .ZN(
        n16873) );
  AOI21_X1 U18823 ( .B1(n17062), .B2(n17668), .A(n16873), .ZN(n16874) );
  OAI21_X1 U18824 ( .B1(n17064), .B2(n17670), .A(n16874), .ZN(P2_U2993) );
  XNOR2_X1 U18825 ( .A(n16875), .B(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17079) );
  AOI21_X1 U18826 ( .B1(n16877), .B2(n16889), .A(n16876), .ZN(n17077) );
  INV_X1 U18827 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n17753) );
  NOR2_X1 U18828 ( .A1(n16970), .A2(n17753), .ZN(n17066) );
  NOR2_X1 U18829 ( .A1(n17631), .A2(n18775), .ZN(n16878) );
  AOI211_X1 U18830 ( .C1(n17661), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n17066), .B(n16878), .ZN(n16879) );
  OAI21_X1 U18831 ( .B1(n18769), .B2(n17651), .A(n16879), .ZN(n16880) );
  AOI21_X1 U18832 ( .B1(n17077), .B2(n17668), .A(n16880), .ZN(n16881) );
  OAI21_X1 U18833 ( .B1(n17079), .B2(n17670), .A(n16881), .ZN(P2_U2994) );
  NAND2_X1 U18834 ( .A1(n16883), .A2(n16882), .ZN(n16886) );
  XNOR2_X1 U18835 ( .A(n16884), .B(n17096), .ZN(n16894) );
  OAI22_X1 U18836 ( .A1(n16894), .A2(n16893), .B1(n17096), .B2(n16884), .ZN(
        n16885) );
  XOR2_X1 U18837 ( .A(n16886), .B(n16885), .Z(n17080) );
  NAND2_X1 U18838 ( .A1(n17647), .A2(n18753), .ZN(n16887) );
  NAND2_X1 U18839 ( .A1(n12161), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n17083) );
  OAI211_X1 U18840 ( .C1(n17658), .C2(n16888), .A(n16887), .B(n17083), .ZN(
        n16891) );
  OAI21_X1 U18841 ( .B1(n16895), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n16889), .ZN(n17090) );
  NOR2_X1 U18842 ( .A1(n17090), .A2(n17648), .ZN(n16890) );
  AOI211_X1 U18843 ( .C1(n17672), .C2(n18755), .A(n16891), .B(n16890), .ZN(
        n16892) );
  OAI21_X1 U18844 ( .B1(n17080), .B2(n17670), .A(n16892), .ZN(P2_U2995) );
  XNOR2_X1 U18845 ( .A(n16894), .B(n16893), .ZN(n17102) );
  NAND2_X1 U18846 ( .A1(n11745), .A2(n17067), .ZN(n16904) );
  AOI21_X1 U18847 ( .B1(n17096), .B2(n16904), .A(n16895), .ZN(n17100) );
  INV_X1 U18848 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n18732) );
  NOR2_X1 U18849 ( .A1(n16970), .A2(n18732), .ZN(n17093) );
  NOR2_X1 U18850 ( .A1(n17631), .A2(n18737), .ZN(n16896) );
  AOI211_X1 U18851 ( .C1(n17661), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n17093), .B(n16896), .ZN(n16897) );
  OAI21_X1 U18852 ( .B1(n18739), .B2(n17651), .A(n16897), .ZN(n16898) );
  AOI21_X1 U18853 ( .B1(n17100), .B2(n17668), .A(n16898), .ZN(n16899) );
  OAI21_X1 U18854 ( .B1(n17102), .B2(n17670), .A(n16899), .ZN(P2_U2996) );
  NOR2_X1 U18855 ( .A1(n16901), .A2(n16900), .ZN(n16902) );
  XNOR2_X1 U18856 ( .A(n16903), .B(n16902), .ZN(n17117) );
  OAI211_X1 U18857 ( .C1(n17107), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n17668), .B(n16904), .ZN(n16908) );
  NAND2_X1 U18858 ( .A1(n17647), .A2(n18719), .ZN(n16905) );
  NAND2_X1 U18859 ( .A1(n16976), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n17108) );
  OAI211_X1 U18860 ( .C1(n17658), .C2(n12330), .A(n16905), .B(n17108), .ZN(
        n16906) );
  AOI21_X1 U18861 ( .B1(n18728), .B2(n17672), .A(n16906), .ZN(n16907) );
  OAI211_X1 U18862 ( .C1(n17117), .C2(n17670), .A(n16908), .B(n16907), .ZN(
        P2_U2997) );
  OAI21_X1 U18863 ( .B1(n17124), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n17668), .ZN(n16916) );
  NAND2_X1 U18864 ( .A1(n16976), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n17118) );
  NAND2_X1 U18865 ( .A1(n17661), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16909) );
  OAI211_X1 U18866 ( .C1(n17631), .C2(n18709), .A(n17118), .B(n16909), .ZN(
        n16914) );
  NOR2_X1 U18867 ( .A1(n16911), .A2(n16910), .ZN(n17120) );
  INV_X1 U18868 ( .A(n16912), .ZN(n17119) );
  NOR3_X1 U18869 ( .A1(n17120), .A2(n17119), .A3(n17670), .ZN(n16913) );
  AOI211_X1 U18870 ( .C1(n18711), .C2(n17672), .A(n16914), .B(n16913), .ZN(
        n16915) );
  OAI21_X1 U18871 ( .B1(n17107), .B2(n16916), .A(n16915), .ZN(P2_U2998) );
  AOI21_X1 U18872 ( .B1(n16943), .B2(n16946), .A(n16942), .ZN(n16935) );
  AND2_X1 U18873 ( .A1(n16919), .A2(n16918), .ZN(n16934) );
  NAND2_X1 U18874 ( .A1(n16935), .A2(n16934), .ZN(n16933) );
  NAND2_X1 U18875 ( .A1(n16933), .A2(n16919), .ZN(n16923) );
  NAND2_X1 U18876 ( .A1(n16921), .A2(n16920), .ZN(n16922) );
  XNOR2_X1 U18877 ( .A(n16923), .B(n16922), .ZN(n17139) );
  INV_X1 U18878 ( .A(n16924), .ZN(n16931) );
  AOI21_X1 U18879 ( .B1(n17129), .B2(n16931), .A(n17124), .ZN(n17137) );
  NAND2_X1 U18880 ( .A1(n16976), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n17132) );
  OAI21_X1 U18881 ( .B1(n17658), .B2(n16925), .A(n17132), .ZN(n16926) );
  AOI21_X1 U18882 ( .B1(n17647), .B2(n18693), .A(n16926), .ZN(n16927) );
  OAI21_X1 U18883 ( .B1(n18699), .B2(n17651), .A(n16927), .ZN(n16928) );
  AOI21_X1 U18884 ( .B1(n17137), .B2(n17668), .A(n16928), .ZN(n16929) );
  OAI21_X1 U18885 ( .B1(n17139), .B2(n17670), .A(n16929), .ZN(P2_U2999) );
  NAND2_X1 U18886 ( .A1(n16957), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17169) );
  OAI21_X1 U18887 ( .B1(n17169), .B2(n17157), .A(n17150), .ZN(n16932) );
  NAND2_X1 U18888 ( .A1(n16932), .A2(n16931), .ZN(n17155) );
  OAI21_X1 U18889 ( .B1(n16935), .B2(n16934), .A(n16933), .ZN(n17153) );
  INV_X1 U18890 ( .A(n18685), .ZN(n16938) );
  INV_X1 U18891 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16936) );
  NAND2_X1 U18892 ( .A1(n16976), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n17146) );
  OAI21_X1 U18893 ( .B1(n17658), .B2(n16936), .A(n17146), .ZN(n16937) );
  AOI21_X1 U18894 ( .B1(n17647), .B2(n16938), .A(n16937), .ZN(n16939) );
  OAI21_X1 U18895 ( .B1(n17143), .B2(n17651), .A(n16939), .ZN(n16940) );
  AOI21_X1 U18896 ( .B1(n17153), .B2(n17617), .A(n16940), .ZN(n16941) );
  OAI21_X1 U18897 ( .B1(n17648), .B2(n17155), .A(n16941), .ZN(P2_U3000) );
  XNOR2_X1 U18898 ( .A(n17169), .B(n17157), .ZN(n17168) );
  INV_X1 U18899 ( .A(n16942), .ZN(n16944) );
  NAND2_X1 U18900 ( .A1(n16944), .A2(n16943), .ZN(n16945) );
  XNOR2_X1 U18901 ( .A(n16946), .B(n16945), .ZN(n17156) );
  NAND2_X1 U18902 ( .A1(n16976), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n17160) );
  OAI21_X1 U18903 ( .B1(n17658), .B2(n16947), .A(n17160), .ZN(n16948) );
  AOI21_X1 U18904 ( .B1(n17647), .B2(n16949), .A(n16948), .ZN(n16950) );
  OAI21_X1 U18905 ( .B1(n17162), .B2(n17651), .A(n16950), .ZN(n16951) );
  AOI21_X1 U18906 ( .B1(n17156), .B2(n17617), .A(n16951), .ZN(n16952) );
  OAI21_X1 U18907 ( .B1(n17648), .B2(n17168), .A(n16952), .ZN(P2_U3001) );
  NAND2_X1 U18908 ( .A1(n16954), .A2(n16953), .ZN(n16955) );
  XNOR2_X1 U18909 ( .A(n16956), .B(n16955), .ZN(n17182) );
  INV_X1 U18910 ( .A(n16957), .ZN(n16963) );
  NAND2_X1 U18911 ( .A1(n16963), .A2(n17177), .ZN(n17170) );
  NAND3_X1 U18912 ( .A1(n17170), .A2(n17668), .A3(n17169), .ZN(n16961) );
  NAND2_X1 U18913 ( .A1(n16976), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n17172) );
  NAND2_X1 U18914 ( .A1(n17661), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16958) );
  OAI211_X1 U18915 ( .C1(n17631), .C2(n18674), .A(n17172), .B(n16958), .ZN(
        n16959) );
  AOI21_X1 U18916 ( .B1(n18676), .B2(n17672), .A(n16959), .ZN(n16960) );
  OAI211_X1 U18917 ( .C1(n17182), .C2(n17670), .A(n16961), .B(n16960), .ZN(
        P2_U3002) );
  NAND2_X1 U18918 ( .A1(n11745), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17654) );
  INV_X1 U18919 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17200) );
  OAI21_X1 U18920 ( .B1(n17654), .B2(n17200), .A(n17184), .ZN(n16962) );
  NAND2_X1 U18921 ( .A1(n16963), .A2(n16962), .ZN(n17195) );
  NAND2_X1 U18922 ( .A1(n16965), .A2(n16964), .ZN(n16968) );
  NOR3_X1 U18923 ( .A1(n16966), .A2(n16981), .A3(n17215), .ZN(n16967) );
  XOR2_X1 U18924 ( .A(n16968), .B(n16967), .Z(n17193) );
  INV_X1 U18925 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n16969) );
  NOR2_X1 U18926 ( .A1(n16970), .A2(n16969), .ZN(n17187) );
  AOI21_X1 U18927 ( .B1(n17661), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n17187), .ZN(n16973) );
  NAND2_X1 U18928 ( .A1(n17647), .A2(n16971), .ZN(n16972) );
  OAI211_X1 U18929 ( .C1(n17190), .C2(n17651), .A(n16973), .B(n16972), .ZN(
        n16974) );
  AOI21_X1 U18930 ( .B1(n17193), .B2(n17617), .A(n16974), .ZN(n16975) );
  OAI21_X1 U18931 ( .B1(n17648), .B2(n17195), .A(n16975), .ZN(P2_U3003) );
  XNOR2_X1 U18932 ( .A(n17654), .B(n17200), .ZN(n17208) );
  NAND2_X1 U18933 ( .A1(n16976), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n17198) );
  NAND2_X1 U18934 ( .A1(n17661), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16977) );
  OAI211_X1 U18935 ( .C1(n17631), .C2(n18663), .A(n17198), .B(n16977), .ZN(
        n16986) );
  NAND2_X1 U18936 ( .A1(n17270), .A2(n16978), .ZN(n17272) );
  NAND2_X1 U18937 ( .A1(n17272), .A2(n16979), .ZN(n17245) );
  NAND2_X1 U18938 ( .A1(n17210), .A2(n16980), .ZN(n17216) );
  INV_X1 U18939 ( .A(n17215), .ZN(n17212) );
  NAND2_X1 U18940 ( .A1(n17216), .A2(n17212), .ZN(n16984) );
  NOR2_X1 U18941 ( .A1(n16982), .A2(n16981), .ZN(n16983) );
  XNOR2_X1 U18942 ( .A(n16984), .B(n16983), .ZN(n17205) );
  NOR2_X1 U18943 ( .A1(n17205), .A2(n17670), .ZN(n16985) );
  AOI211_X1 U18944 ( .C1(n17672), .C2(n18665), .A(n16986), .B(n16985), .ZN(
        n16987) );
  OAI21_X1 U18945 ( .B1(n17648), .B2(n17208), .A(n16987), .ZN(P2_U3004) );
  OAI21_X1 U18946 ( .B1(n16990), .B2(n16989), .A(n10976), .ZN(n17240) );
  NAND2_X1 U18947 ( .A1(n16991), .A2(n17241), .ZN(n16996) );
  INV_X1 U18948 ( .A(n16992), .ZN(n16993) );
  NOR2_X1 U18949 ( .A1(n16994), .A2(n16993), .ZN(n16995) );
  XNOR2_X1 U18950 ( .A(n16996), .B(n16995), .ZN(n17237) );
  INV_X1 U18951 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n18647) );
  OAI22_X1 U18952 ( .A1(n18647), .A2(n18746), .B1(n17631), .B2(n18650), .ZN(
        n16999) );
  INV_X1 U18953 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16997) );
  OAI22_X1 U18954 ( .A1(n18652), .A2(n17651), .B1(n16997), .B2(n17658), .ZN(
        n16998) );
  AOI211_X1 U18955 ( .C1(n17237), .C2(n17617), .A(n16999), .B(n16998), .ZN(
        n17000) );
  OAI21_X1 U18956 ( .B1(n17240), .B2(n17648), .A(n17000), .ZN(P2_U3006) );
  INV_X1 U18957 ( .A(n18856), .ZN(n17007) );
  AOI21_X1 U18958 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17004), .A(
        n17003), .ZN(n17002) );
  AOI211_X1 U18959 ( .C1(n17004), .C2(n17003), .A(n17002), .B(n17001), .ZN(
        n17005) );
  NAND2_X1 U18960 ( .A1(n17008), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17009) );
  OAI211_X1 U18961 ( .C1(n18858), .C2(n18885), .A(n17010), .B(n17009), .ZN(
        n17011) );
  AOI21_X1 U18962 ( .B1(n17012), .B2(n18879), .A(n17011), .ZN(n17013) );
  OAI21_X1 U18963 ( .B1(n17014), .B2(n18881), .A(n17013), .ZN(P2_U3017) );
  NOR2_X1 U18964 ( .A1(n17229), .A2(n18829), .ZN(n17016) );
  AOI211_X1 U18965 ( .C1(n17017), .C2(n13712), .A(n17016), .B(n17015), .ZN(
        n17019) );
  NOR3_X1 U18966 ( .A1(n17035), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n17036), .ZN(n17024) );
  OAI21_X1 U18967 ( .B1(n17026), .B2(n17024), .A(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17018) );
  OAI211_X1 U18968 ( .C1(n18830), .C2(n18885), .A(n17019), .B(n17018), .ZN(
        n17020) );
  AOI21_X1 U18969 ( .B1(n17021), .B2(n18879), .A(n17020), .ZN(n17022) );
  OAI21_X1 U18970 ( .B1(n17023), .B2(n18881), .A(n17022), .ZN(P2_U3020) );
  AOI211_X1 U18971 ( .C1(n18876), .C2(n18816), .A(n17025), .B(n17024), .ZN(
        n17028) );
  NAND2_X1 U18972 ( .A1(n17026), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17027) );
  OAI211_X1 U18973 ( .C1(n18818), .C2(n18885), .A(n17028), .B(n17027), .ZN(
        n17029) );
  AOI21_X1 U18974 ( .B1(n17030), .B2(n18879), .A(n17029), .ZN(n17031) );
  OAI21_X1 U18975 ( .B1(n17032), .B2(n18881), .A(n17031), .ZN(P2_U3021) );
  NAND2_X1 U18976 ( .A1(n17033), .A2(n12326), .ZN(n17041) );
  AOI21_X1 U18977 ( .B1(n17036), .B2(n17035), .A(n17034), .ZN(n17039) );
  OAI21_X1 U18978 ( .B1(n17229), .B2(n18814), .A(n17037), .ZN(n17038) );
  AOI211_X1 U18979 ( .C1(n18810), .C2(n17204), .A(n17039), .B(n17038), .ZN(
        n17040) );
  OAI211_X1 U18980 ( .C1(n17277), .C2(n17042), .A(n17041), .B(n17040), .ZN(
        P2_U3022) );
  NOR3_X1 U18981 ( .A1(n17044), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n17043), .ZN(n17045) );
  AOI211_X1 U18982 ( .C1(n18876), .C2(n19584), .A(n17046), .B(n17045), .ZN(
        n17049) );
  NAND2_X1 U18983 ( .A1(n17047), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17048) );
  OAI211_X1 U18984 ( .C1(n17050), .C2(n18885), .A(n17049), .B(n17048), .ZN(
        n17051) );
  AOI21_X1 U18985 ( .B1(n17052), .B2(n18879), .A(n17051), .ZN(n17053) );
  OAI21_X1 U18986 ( .B1(n17054), .B2(n18881), .A(n17053), .ZN(P2_U3024) );
  AOI211_X1 U18987 ( .C1(n18876), .C2(n17057), .A(n17056), .B(n17055), .ZN(
        n17060) );
  NAND2_X1 U18988 ( .A1(n17058), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n17059) );
  OAI211_X1 U18989 ( .C1(n18779), .C2(n18885), .A(n17060), .B(n17059), .ZN(
        n17061) );
  AOI21_X1 U18990 ( .B1(n17062), .B2(n18879), .A(n17061), .ZN(n17063) );
  OAI21_X1 U18991 ( .B1(n17064), .B2(n18881), .A(n17063), .ZN(P2_U3025) );
  NAND2_X1 U18992 ( .A1(n17067), .A2(n17218), .ZN(n17091) );
  NOR4_X1 U18993 ( .A1(n17091), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n17072), .A4(n17096), .ZN(n17065) );
  AOI211_X1 U18994 ( .C1(n18876), .C2(n18762), .A(n17066), .B(n17065), .ZN(
        n17075) );
  INV_X1 U18995 ( .A(n17103), .ZN(n17071) );
  INV_X1 U18996 ( .A(n17067), .ZN(n17068) );
  AOI22_X1 U18997 ( .A1(n17104), .A2(n17069), .B1(n17103), .B2(n17068), .ZN(
        n17070) );
  AND2_X1 U18998 ( .A1(n17222), .A2(n17070), .ZN(n17097) );
  OAI21_X1 U18999 ( .B1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n17071), .A(
        n17097), .ZN(n17087) );
  NAND2_X1 U19000 ( .A1(n17072), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17073) );
  NOR2_X1 U19001 ( .A1(n17091), .A2(n17073), .ZN(n17081) );
  OAI21_X1 U19002 ( .B1(n17087), .B2(n17081), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17074) );
  OAI211_X1 U19003 ( .C1(n18769), .C2(n18885), .A(n17075), .B(n17074), .ZN(
        n17076) );
  AOI21_X1 U19004 ( .B1(n17077), .B2(n18879), .A(n17076), .ZN(n17078) );
  OAI21_X1 U19005 ( .B1(n17079), .B2(n18881), .A(n17078), .ZN(P2_U3026) );
  OR2_X1 U19006 ( .A1(n17080), .A2(n18881), .ZN(n17089) );
  INV_X1 U19007 ( .A(n17081), .ZN(n17082) );
  OAI211_X1 U19008 ( .C1(n17229), .C2(n18759), .A(n17083), .B(n17082), .ZN(
        n17086) );
  NOR2_X1 U19009 ( .A1(n17084), .A2(n18885), .ZN(n17085) );
  AOI211_X1 U19010 ( .C1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17087), .A(
        n17086), .B(n17085), .ZN(n17088) );
  OAI211_X1 U19011 ( .C1(n17090), .C2(n17277), .A(n17089), .B(n17088), .ZN(
        P2_U3027) );
  NOR2_X1 U19012 ( .A1(n18739), .A2(n18885), .ZN(n17099) );
  INV_X1 U19013 ( .A(n18744), .ZN(n17094) );
  NOR2_X1 U19014 ( .A1(n17091), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17092) );
  AOI211_X1 U19015 ( .C1(n17094), .C2(n18876), .A(n17093), .B(n17092), .ZN(
        n17095) );
  OAI21_X1 U19016 ( .B1(n17097), .B2(n17096), .A(n17095), .ZN(n17098) );
  AOI211_X1 U19017 ( .C1(n17100), .C2(n18879), .A(n17099), .B(n17098), .ZN(
        n17101) );
  OAI21_X1 U19018 ( .B1(n17102), .B2(n18881), .A(n17101), .ZN(P2_U3028) );
  NOR2_X1 U19019 ( .A1(n18879), .A2(n17103), .ZN(n17123) );
  INV_X1 U19020 ( .A(n17130), .ZN(n17110) );
  AOI22_X1 U19021 ( .A1(n17262), .A2(n17110), .B1(n17104), .B2(n17129), .ZN(
        n17105) );
  NAND2_X1 U19022 ( .A1(n17222), .A2(n17105), .ZN(n17134) );
  AOI21_X1 U19023 ( .B1(n17112), .B2(n17262), .A(n17134), .ZN(n17106) );
  OAI21_X1 U19024 ( .B1(n17107), .B2(n17123), .A(n17106), .ZN(n17115) );
  NAND2_X1 U19025 ( .A1(n18728), .A2(n17204), .ZN(n17109) );
  OAI211_X1 U19026 ( .C1(n17229), .C2(n18726), .A(n17109), .B(n17108), .ZN(
        n17114) );
  INV_X1 U19027 ( .A(n17218), .ZN(n17140) );
  NOR3_X1 U19028 ( .A1(n17110), .A2(n17129), .A3(n17140), .ZN(n17111) );
  AOI21_X1 U19029 ( .B1(n17124), .B2(n18879), .A(n17111), .ZN(n17128) );
  NOR3_X1 U19030 ( .A1(n17128), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n17112), .ZN(n17113) );
  OAI21_X1 U19031 ( .B1(n17117), .B2(n18881), .A(n17116), .ZN(P2_U3029) );
  OAI21_X1 U19032 ( .B1(n18715), .B2(n17229), .A(n17118), .ZN(n17122) );
  NOR3_X1 U19033 ( .A1(n17120), .A2(n17119), .A3(n18881), .ZN(n17121) );
  AOI211_X1 U19034 ( .C1(n17204), .C2(n18711), .A(n17122), .B(n17121), .ZN(
        n17127) );
  NOR2_X1 U19035 ( .A1(n17124), .A2(n17123), .ZN(n17125) );
  OAI21_X1 U19036 ( .B1(n17125), .B2(n17134), .A(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17126) );
  OAI211_X1 U19037 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n17128), .A(
        n17127), .B(n17126), .ZN(P2_U3030) );
  NAND3_X1 U19038 ( .A1(n17130), .A2(n17218), .A3(n17129), .ZN(n17131) );
  OAI211_X1 U19039 ( .C1(n17229), .C2(n18698), .A(n17132), .B(n17131), .ZN(
        n17133) );
  AOI21_X1 U19040 ( .B1(n17134), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n17133), .ZN(n17135) );
  OAI21_X1 U19041 ( .B1(n18699), .B2(n18885), .A(n17135), .ZN(n17136) );
  AOI21_X1 U19042 ( .B1(n17137), .B2(n18879), .A(n17136), .ZN(n17138) );
  OAI21_X1 U19043 ( .B1(n17139), .B2(n18881), .A(n17138), .ZN(P2_U3031) );
  NOR2_X1 U19044 ( .A1(n17141), .A2(n17140), .ZN(n17158) );
  NAND2_X1 U19045 ( .A1(n17262), .A2(n17141), .ZN(n17142) );
  AND2_X1 U19046 ( .A1(n17222), .A2(n17142), .ZN(n17178) );
  NAND2_X1 U19047 ( .A1(n17158), .A2(n17177), .ZN(n17171) );
  NAND2_X1 U19048 ( .A1(n17178), .A2(n17171), .ZN(n17165) );
  AOI21_X1 U19049 ( .B1(n17158), .B2(n17157), .A(n17165), .ZN(n17151) );
  INV_X1 U19050 ( .A(n17143), .ZN(n18687) );
  OAI21_X1 U19051 ( .B1(n15134), .B2(n17145), .A(n17144), .ZN(n19363) );
  NAND4_X1 U19052 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n17158), .A4(n17150), .ZN(
        n17147) );
  OAI211_X1 U19053 ( .C1(n17229), .C2(n19363), .A(n17147), .B(n17146), .ZN(
        n17148) );
  AOI21_X1 U19054 ( .B1(n18687), .B2(n17204), .A(n17148), .ZN(n17149) );
  OAI21_X1 U19055 ( .B1(n17151), .B2(n17150), .A(n17149), .ZN(n17152) );
  AOI21_X1 U19056 ( .B1(n17153), .B2(n12326), .A(n17152), .ZN(n17154) );
  OAI21_X1 U19057 ( .B1(n17277), .B2(n17155), .A(n17154), .ZN(P2_U3032) );
  NAND2_X1 U19058 ( .A1(n17156), .A2(n12326), .ZN(n17167) );
  NAND3_X1 U19059 ( .A1(n17158), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        n17157), .ZN(n17159) );
  OAI211_X1 U19060 ( .C1(n17229), .C2(n17161), .A(n17160), .B(n17159), .ZN(
        n17164) );
  NOR2_X1 U19061 ( .A1(n17162), .A2(n18885), .ZN(n17163) );
  AOI211_X1 U19062 ( .C1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n17165), .A(
        n17164), .B(n17163), .ZN(n17166) );
  OAI211_X1 U19063 ( .C1(n17168), .C2(n17277), .A(n17167), .B(n17166), .ZN(
        P2_U3033) );
  NAND3_X1 U19064 ( .A1(n17170), .A2(n18879), .A3(n17169), .ZN(n17181) );
  NAND2_X1 U19065 ( .A1(n18676), .A2(n17204), .ZN(n17176) );
  INV_X1 U19066 ( .A(n18680), .ZN(n17174) );
  NAND2_X1 U19067 ( .A1(n17172), .A2(n17171), .ZN(n17173) );
  AOI21_X1 U19068 ( .B1(n18876), .B2(n17174), .A(n17173), .ZN(n17175) );
  OAI211_X1 U19069 ( .C1(n17178), .C2(n17177), .A(n17176), .B(n17175), .ZN(
        n17179) );
  INV_X1 U19070 ( .A(n17179), .ZN(n17180) );
  OAI211_X1 U19071 ( .C1(n17182), .C2(n18881), .A(n17181), .B(n17180), .ZN(
        P2_U3034) );
  INV_X1 U19072 ( .A(n17222), .ZN(n17183) );
  AOI21_X1 U19073 ( .B1(n17221), .B2(n17262), .A(n17183), .ZN(n17201) );
  NAND3_X1 U19074 ( .A1(n17200), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n17218), .ZN(n17197) );
  AOI21_X1 U19075 ( .B1(n17201), .B2(n17197), .A(n17184), .ZN(n17192) );
  AND3_X1 U19076 ( .A1(n17185), .A2(n17218), .A3(n17184), .ZN(n17186) );
  AOI211_X1 U19077 ( .C1(n18876), .C2(n17188), .A(n17187), .B(n17186), .ZN(
        n17189) );
  OAI21_X1 U19078 ( .B1(n17190), .B2(n18885), .A(n17189), .ZN(n17191) );
  AOI211_X1 U19079 ( .C1(n17193), .C2(n12326), .A(n17192), .B(n17191), .ZN(
        n17194) );
  OAI21_X1 U19080 ( .B1(n17277), .B2(n17195), .A(n17194), .ZN(P2_U3035) );
  INV_X1 U19081 ( .A(n18669), .ZN(n17196) );
  NAND2_X1 U19082 ( .A1(n18876), .A2(n17196), .ZN(n17199) );
  NAND3_X1 U19083 ( .A1(n17199), .A2(n17198), .A3(n17197), .ZN(n17203) );
  NOR2_X1 U19084 ( .A1(n17201), .A2(n17200), .ZN(n17202) );
  AOI211_X1 U19085 ( .C1(n18665), .C2(n17204), .A(n17203), .B(n17202), .ZN(
        n17207) );
  OR2_X1 U19086 ( .A1(n17205), .A2(n18881), .ZN(n17206) );
  OAI211_X1 U19087 ( .C1(n17208), .C2(n17277), .A(n17207), .B(n17206), .ZN(
        P2_U3036) );
  AND2_X1 U19088 ( .A1(n17210), .A2(n17209), .ZN(n17214) );
  AND2_X1 U19089 ( .A1(n17212), .A2(n17211), .ZN(n17213) );
  OAI22_X1 U19090 ( .A1(n17216), .A2(n17215), .B1(n17214), .B2(n17213), .ZN(
        n17652) );
  NOR2_X1 U19091 ( .A1(n11745), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17649) );
  INV_X1 U19092 ( .A(n17649), .ZN(n17217) );
  NAND3_X1 U19093 ( .A1(n17217), .A2(n18879), .A3(n17654), .ZN(n17226) );
  NAND2_X1 U19094 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n12161), .ZN(n17220) );
  NAND2_X1 U19095 ( .A1(n17221), .A2(n17218), .ZN(n17219) );
  OAI211_X1 U19096 ( .C1(n17650), .C2(n18885), .A(n17220), .B(n17219), .ZN(
        n17224) );
  NOR2_X1 U19097 ( .A1(n17222), .A2(n17221), .ZN(n17223) );
  AOI211_X1 U19098 ( .C1(n18876), .C2(n19370), .A(n17224), .B(n17223), .ZN(
        n17225) );
  OAI211_X1 U19099 ( .C1(n17652), .C2(n18881), .A(n17226), .B(n17225), .ZN(
        P2_U3037) );
  OAI21_X1 U19100 ( .B1(n18890), .B2(n17228), .A(n17227), .ZN(n17249) );
  NOR2_X1 U19101 ( .A1(n17229), .A2(n18657), .ZN(n17236) );
  AOI211_X1 U19102 ( .C1(n17252), .C2(n17232), .A(n17231), .B(n17230), .ZN(
        n17233) );
  AOI21_X1 U19103 ( .B1(n12161), .B2(P2_REIP_REG_8__SCAN_IN), .A(n17233), .ZN(
        n17234) );
  OAI21_X1 U19104 ( .B1(n18652), .B2(n18885), .A(n17234), .ZN(n17235) );
  AOI211_X1 U19105 ( .C1(n17249), .C2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n17236), .B(n17235), .ZN(n17239) );
  NAND2_X1 U19106 ( .A1(n17237), .A2(n12326), .ZN(n17238) );
  OAI211_X1 U19107 ( .C1(n17240), .C2(n17277), .A(n17239), .B(n17238), .ZN(
        P2_U3038) );
  INV_X1 U19108 ( .A(n17241), .ZN(n17243) );
  NOR2_X1 U19109 ( .A1(n17243), .A2(n17242), .ZN(n17244) );
  XNOR2_X1 U19110 ( .A(n17245), .B(n17244), .ZN(n17639) );
  NOR2_X1 U19111 ( .A1(n17247), .A2(n17246), .ZN(n17638) );
  INV_X1 U19112 ( .A(n17638), .ZN(n17248) );
  NAND3_X1 U19113 ( .A1(n17248), .A2(n18879), .A3(n17641), .ZN(n17258) );
  NAND2_X1 U19114 ( .A1(n17249), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17254) );
  INV_X1 U19115 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n18638) );
  NOR2_X1 U19116 ( .A1(n18638), .A2(n18746), .ZN(n17250) );
  AOI21_X1 U19117 ( .B1(n17252), .B2(n17251), .A(n17250), .ZN(n17253) );
  OAI211_X1 U19118 ( .C1(n18639), .C2(n18885), .A(n17254), .B(n17253), .ZN(
        n17255) );
  AOI21_X1 U19119 ( .B1(n17256), .B2(n18876), .A(n17255), .ZN(n17257) );
  OAI211_X1 U19120 ( .C1(n17639), .C2(n18881), .A(n17258), .B(n17257), .ZN(
        P2_U3039) );
  OAI21_X1 U19121 ( .B1(n17260), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n17259), .ZN(n17634) );
  AOI21_X1 U19122 ( .B1(n17263), .B2(n17262), .A(n17261), .ZN(n17269) );
  INV_X1 U19123 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n18626) );
  NOR2_X1 U19124 ( .A1(n18626), .A2(n18746), .ZN(n17265) );
  NOR2_X1 U19125 ( .A1(n18885), .A2(n18627), .ZN(n17264) );
  AOI211_X1 U19126 ( .C1(n17266), .C2(n17268), .A(n17265), .B(n17264), .ZN(
        n17267) );
  OAI21_X1 U19127 ( .B1(n17269), .B2(n17268), .A(n17267), .ZN(n17274) );
  OR2_X1 U19128 ( .A1(n17270), .A2(n16978), .ZN(n17271) );
  NAND2_X1 U19129 ( .A1(n17272), .A2(n17271), .ZN(n17633) );
  NOR2_X1 U19130 ( .A1(n17633), .A2(n18881), .ZN(n17273) );
  AOI211_X1 U19131 ( .C1(n18876), .C2(n17275), .A(n17274), .B(n17273), .ZN(
        n17276) );
  OAI21_X1 U19132 ( .B1(n17277), .B2(n17634), .A(n17276), .ZN(P2_U3040) );
  INV_X1 U19133 ( .A(n18906), .ZN(n17292) );
  AOI211_X1 U19134 ( .C1(n18595), .C2(n17279), .A(n18717), .B(n17278), .ZN(
        n18615) );
  AOI21_X1 U19135 ( .B1(n18717), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n18615), .ZN(n17284) );
  NOR2_X1 U19136 ( .A1(n17280), .A2(n17326), .ZN(n17285) );
  AOI22_X1 U19137 ( .A1(n17281), .A2(n17287), .B1(n17284), .B2(n17285), .ZN(
        n17282) );
  OAI21_X1 U19138 ( .B1(n19408), .B2(n17292), .A(n17282), .ZN(n17283) );
  MUX2_X1 U19139 ( .A(n17283), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n18868), .Z(P2_U3600) );
  INV_X1 U19140 ( .A(n17284), .ZN(n17286) );
  AOI222_X1 U19141 ( .A1(n17288), .A2(n17287), .B1(n18906), .B2(n19502), .C1(
        n17286), .C2(n17285), .ZN(n17290) );
  NAND2_X1 U19142 ( .A1(n18868), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n17289) );
  OAI21_X1 U19143 ( .B1(n17290), .B2(n18868), .A(n17289), .ZN(P2_U3599) );
  OAI22_X1 U19144 ( .A1(n19426), .A2(n17292), .B1(n17291), .B2(n18892), .ZN(
        n17293) );
  MUX2_X1 U19145 ( .A(n17293), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n18868), .Z(P2_U3596) );
  NAND2_X1 U19146 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18944) );
  INV_X1 U19147 ( .A(n18076), .ZN(n17294) );
  NOR2_X1 U19148 ( .A1(n20997), .A2(n21823), .ZN(n18329) );
  OAI21_X1 U19149 ( .B1(n17294), .B2(n18329), .A(n21488), .ZN(n17296) );
  NOR2_X1 U19150 ( .A1(n20337), .A2(n18076), .ZN(n17314) );
  INV_X1 U19151 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17309) );
  OAI21_X1 U19152 ( .B1(n21021), .B2(n21001), .A(n17309), .ZN(n17295) );
  INV_X1 U19153 ( .A(n17295), .ZN(n17307) );
  NAND2_X1 U19154 ( .A1(n17307), .A2(n17984), .ZN(n18077) );
  AOI221_X1 U19155 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(n17314), .C1(n18077), .C2(
        n17314), .A(n19259), .ZN(n18474) );
  NAND2_X1 U19156 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n21449), .ZN(n18974) );
  INV_X1 U19157 ( .A(n18974), .ZN(n18475) );
  AOI211_X1 U19158 ( .C1(n18944), .C2(n17296), .A(n18474), .B(n18475), .ZN(
        n18471) );
  INV_X1 U19159 ( .A(n18079), .ZN(n20278) );
  INV_X1 U19160 ( .A(n18329), .ZN(n18427) );
  NAND2_X1 U19161 ( .A1(n20278), .A2(n18427), .ZN(n17297) );
  OAI21_X1 U19162 ( .B1(n21449), .B2(n21488), .A(n17297), .ZN(n18472) );
  INV_X1 U19163 ( .A(n18474), .ZN(n18473) );
  OAI221_X1 U19164 ( .B1(n18979), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18979), .C2(n18472), .A(n18473), .ZN(n17298) );
  AOI22_X1 U19165 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18471), .B1(
        n17298), .B2(n18968), .ZN(P3_U2865) );
  NOR2_X1 U19166 ( .A1(n21445), .A2(n17299), .ZN(n17305) );
  INV_X1 U19167 ( .A(n21478), .ZN(n21876) );
  INV_X1 U19168 ( .A(n20348), .ZN(n17301) );
  NOR4_X1 U19169 ( .A1(n21876), .A2(n17302), .A3(n21471), .A4(n17301), .ZN(
        n17304) );
  NOR4_X1 U19170 ( .A1(n17305), .A2(n20797), .A3(n17304), .A4(n17303), .ZN(
        n21462) );
  INV_X1 U19171 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n21506) );
  INV_X1 U19172 ( .A(n17314), .ZN(n21486) );
  OAI22_X1 U19173 ( .A1(n11085), .A2(n21500), .B1(n21506), .B2(n21486), .ZN(
        n17306) );
  NOR2_X1 U19174 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n21036) );
  NOR2_X1 U19175 ( .A1(n17307), .A2(n17318), .ZN(n21447) );
  NAND3_X1 U19176 ( .A1(n21038), .A2(n21036), .A3(n21447), .ZN(n17308) );
  OAI21_X1 U19177 ( .B1(n21038), .B2(n17309), .A(n17308), .ZN(P3_U3284) );
  INV_X1 U19178 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17311) );
  OAI21_X1 U19179 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(n21870), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n18535) );
  AND2_X1 U19180 ( .A1(n18561), .A2(n18535), .ZN(n21826) );
  NOR2_X1 U19181 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n21827) );
  OAI21_X1 U19182 ( .B1(BS16), .B2(n21827), .A(n21826), .ZN(n21824) );
  INV_X1 U19183 ( .A(n21824), .ZN(n17310) );
  AOI21_X1 U19184 ( .B1(n17311), .B2(n17312), .A(n17310), .ZN(P3_U3280) );
  AND2_X1 U19185 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n17312), .ZN(P3_U3028) );
  AND2_X1 U19186 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n17312), .ZN(P3_U3027) );
  AND2_X1 U19187 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n17312), .ZN(P3_U3026) );
  AND2_X1 U19188 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n17312), .ZN(P3_U3025) );
  AND2_X1 U19189 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n17312), .ZN(P3_U3024) );
  AND2_X1 U19190 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n17312), .ZN(P3_U3023) );
  AND2_X1 U19191 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n17312), .ZN(P3_U3022) );
  AND2_X1 U19192 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n17312), .ZN(P3_U3021) );
  AND2_X1 U19193 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n17312), .ZN(
        P3_U3020) );
  AND2_X1 U19194 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n17312), .ZN(
        P3_U3019) );
  AND2_X1 U19195 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n17312), .ZN(
        P3_U3018) );
  AND2_X1 U19196 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n17312), .ZN(
        P3_U3017) );
  AND2_X1 U19197 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n17312), .ZN(
        P3_U3016) );
  AND2_X1 U19198 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n17312), .ZN(
        P3_U3015) );
  AND2_X1 U19199 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n17312), .ZN(
        P3_U3014) );
  AND2_X1 U19200 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n17312), .ZN(
        P3_U3013) );
  AND2_X1 U19201 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n17312), .ZN(
        P3_U3012) );
  AND2_X1 U19202 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n17312), .ZN(
        P3_U3011) );
  AND2_X1 U19203 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n17312), .ZN(
        P3_U3010) );
  AND2_X1 U19204 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n17312), .ZN(
        P3_U3009) );
  AND2_X1 U19205 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n17312), .ZN(
        P3_U3008) );
  AND2_X1 U19206 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n17312), .ZN(
        P3_U3007) );
  AND2_X1 U19207 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n17312), .ZN(
        P3_U3006) );
  AND2_X1 U19208 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n17312), .ZN(
        P3_U3005) );
  AND2_X1 U19209 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n17312), .ZN(
        P3_U3004) );
  AND2_X1 U19210 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n17312), .ZN(
        P3_U3003) );
  AND2_X1 U19211 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n17312), .ZN(
        P3_U3002) );
  AND2_X1 U19212 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n17312), .ZN(
        P3_U3001) );
  AND2_X1 U19213 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n17312), .ZN(
        P3_U3000) );
  AND2_X1 U19214 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n17312), .ZN(
        P3_U2999) );
  AOI21_X1 U19215 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n17315)
         );
  NAND4_X1 U19216 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(n21876), .A4(n21352), .ZN(n21483) );
  INV_X1 U19217 ( .A(n21483), .ZN(n17313) );
  AOI211_X1 U19218 ( .C1(n18427), .C2(n17315), .A(n17314), .B(n17313), .ZN(
        P3_U2998) );
  NOR2_X1 U19219 ( .A1(n17316), .A2(n18473), .ZN(P3_U2867) );
  INV_X1 U19220 ( .A(n18196), .ZN(n18464) );
  AND2_X1 U19221 ( .A1(n18525), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U19222 ( .A(n17318), .ZN(n21439) );
  AND2_X1 U19223 ( .A1(n18075), .A2(n20339), .ZN(n17320) );
  INV_X1 U19224 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n17319) );
  AOI22_X1 U19225 ( .A1(n17320), .A2(n17319), .B1(n20341), .B2(n20275), .ZN(
        P3_U3298) );
  INV_X1 U19226 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18496) );
  NAND2_X1 U19227 ( .A1(n19262), .A2(n20341), .ZN(n20791) );
  INV_X1 U19228 ( .A(n20791), .ZN(n20390) );
  AOI21_X1 U19229 ( .B1(n17320), .B2(n18496), .A(n20390), .ZN(P3_U3299) );
  NOR2_X1 U19230 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n17321), .ZN(n21859) );
  AOI21_X1 U19231 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21859), .A(n21852), 
        .ZN(n17323) );
  INV_X1 U19232 ( .A(n17323), .ZN(n21822) );
  INV_X1 U19233 ( .A(n21822), .ZN(n17708) );
  INV_X1 U19234 ( .A(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17341) );
  INV_X1 U19235 ( .A(BS16), .ZN(n17556) );
  NAND2_X1 U19236 ( .A1(n21851), .A2(n17321), .ZN(n17322) );
  AOI21_X1 U19237 ( .B1(n17556), .B2(n17322), .A(n17708), .ZN(n21818) );
  AOI21_X1 U19238 ( .B1(n17708), .B2(n17341), .A(n21818), .ZN(P2_U3591) );
  AND2_X1 U19239 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n17708), .ZN(P2_U3208) );
  AND2_X1 U19240 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n17323), .ZN(P2_U3207) );
  AND2_X1 U19241 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n17708), .ZN(P2_U3206) );
  AND2_X1 U19242 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n17708), .ZN(P2_U3205) );
  AND2_X1 U19243 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n17708), .ZN(P2_U3204) );
  AND2_X1 U19244 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n17708), .ZN(P2_U3203) );
  AND2_X1 U19245 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n17323), .ZN(P2_U3202) );
  AND2_X1 U19246 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n17323), .ZN(P2_U3201) );
  AND2_X1 U19247 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n17323), .ZN(
        P2_U3200) );
  AND2_X1 U19248 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n17323), .ZN(
        P2_U3199) );
  AND2_X1 U19249 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n17323), .ZN(
        P2_U3198) );
  AND2_X1 U19250 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n17323), .ZN(
        P2_U3197) );
  AND2_X1 U19251 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n17323), .ZN(
        P2_U3196) );
  AND2_X1 U19252 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n17323), .ZN(
        P2_U3195) );
  AND2_X1 U19253 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n17323), .ZN(
        P2_U3194) );
  AND2_X1 U19254 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n17323), .ZN(
        P2_U3193) );
  AND2_X1 U19255 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n17323), .ZN(
        P2_U3192) );
  AND2_X1 U19256 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n17323), .ZN(
        P2_U3191) );
  AND2_X1 U19257 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n17708), .ZN(
        P2_U3190) );
  AND2_X1 U19258 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n17708), .ZN(
        P2_U3189) );
  AND2_X1 U19259 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n17708), .ZN(
        P2_U3188) );
  AND2_X1 U19260 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n17708), .ZN(
        P2_U3187) );
  AND2_X1 U19261 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n17323), .ZN(
        P2_U3186) );
  AND2_X1 U19262 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n17708), .ZN(
        P2_U3185) );
  AND2_X1 U19263 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n17708), .ZN(
        P2_U3184) );
  AND2_X1 U19264 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n17708), .ZN(
        P2_U3183) );
  AND2_X1 U19265 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n17708), .ZN(
        P2_U3182) );
  AND2_X1 U19266 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n17708), .ZN(
        P2_U3181) );
  AND2_X1 U19267 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n17708), .ZN(
        P2_U3180) );
  AND2_X1 U19268 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n17708), .ZN(
        P2_U3179) );
  NAND2_X1 U19269 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n18908), .ZN(n18893) );
  AOI21_X1 U19270 ( .B1(n17324), .B2(n11407), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17325) );
  AOI221_X1 U19271 ( .B1(n18893), .B2(n17325), .C1(n17326), .C2(n17325), .A(
        n17329), .ZN(P2_U3178) );
  AOI21_X1 U19272 ( .B1(n19470), .B2(n17326), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n18909) );
  INV_X1 U19273 ( .A(n19382), .ZN(n17327) );
  INV_X1 U19274 ( .A(n17696), .ZN(n17688) );
  NOR2_X1 U19275 ( .A1(n17330), .A2(n17688), .ZN(P2_U3047) );
  AND2_X1 U19276 ( .A1(n17721), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  NOR4_X1 U19277 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n17334) );
  NOR4_X1 U19278 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n17333) );
  NOR4_X1 U19279 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n17332) );
  NOR4_X1 U19280 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n17331) );
  NAND4_X1 U19281 ( .A1(n17334), .A2(n17333), .A3(n17332), .A4(n17331), .ZN(
        n17340) );
  NOR4_X1 U19282 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n17338) );
  AOI211_X1 U19283 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_31__SCAN_IN), .B(
        P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n17337) );
  NOR4_X1 U19284 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n17336) );
  NOR4_X1 U19285 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n17335) );
  NAND4_X1 U19286 ( .A1(n17338), .A2(n17337), .A3(n17336), .A4(n17335), .ZN(
        n17339) );
  NOR2_X1 U19287 ( .A1(n17340), .A2(n17339), .ZN(n17704) );
  INV_X1 U19288 ( .A(n17704), .ZN(n17703) );
  NOR2_X1 U19289 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n17703), .ZN(n17697) );
  INV_X1 U19290 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n17698) );
  INV_X1 U19291 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21821) );
  NAND3_X1 U19292 ( .A1(n17698), .A2(n21821), .A3(n17341), .ZN(n17702) );
  INV_X1 U19293 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n17769) );
  AOI22_X1 U19294 ( .A1(n17697), .A2(n17702), .B1(n17703), .B2(n17769), .ZN(
        P2_U2821) );
  INV_X1 U19295 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n17767) );
  AOI22_X1 U19296 ( .A1(n17697), .A2(n17698), .B1(n17703), .B2(n17767), .ZN(
        P2_U2820) );
  INV_X1 U19297 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17342) );
  INV_X1 U19298 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n21840) );
  AOI21_X1 U19299 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21840), .A(n21847), 
        .ZN(n21835) );
  NAND2_X1 U19300 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n21847), .ZN(n22398) );
  NAND2_X1 U19301 ( .A1(n21840), .A2(n21847), .ZN(n20206) );
  AOI21_X1 U19302 ( .B1(n17556), .B2(n20206), .A(n17343), .ZN(n21816) );
  AOI21_X1 U19303 ( .B1(n17342), .B2(n17343), .A(n21816), .ZN(P1_U3464) );
  AND2_X1 U19304 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n17343), .ZN(P1_U3193) );
  AND2_X1 U19305 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n17343), .ZN(P1_U3192) );
  AND2_X1 U19306 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n17343), .ZN(P1_U3191) );
  AND2_X1 U19307 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n17343), .ZN(P1_U3190) );
  AND2_X1 U19308 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n17343), .ZN(P1_U3189) );
  AND2_X1 U19309 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n17343), .ZN(P1_U3188) );
  AND2_X1 U19310 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n17343), .ZN(P1_U3187) );
  AND2_X1 U19311 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n17343), .ZN(P1_U3186) );
  AND2_X1 U19312 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n17343), .ZN(
        P1_U3185) );
  AND2_X1 U19313 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n17343), .ZN(
        P1_U3184) );
  AND2_X1 U19314 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n17343), .ZN(
        P1_U3183) );
  AND2_X1 U19315 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n17343), .ZN(
        P1_U3182) );
  AND2_X1 U19316 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n17343), .ZN(
        P1_U3181) );
  AND2_X1 U19317 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n17343), .ZN(
        P1_U3180) );
  AND2_X1 U19318 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n17343), .ZN(
        P1_U3179) );
  AND2_X1 U19319 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n17343), .ZN(
        P1_U3178) );
  AND2_X1 U19320 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n17343), .ZN(
        P1_U3177) );
  AND2_X1 U19321 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n17343), .ZN(
        P1_U3176) );
  AND2_X1 U19322 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n17343), .ZN(
        P1_U3175) );
  AND2_X1 U19323 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n17343), .ZN(
        P1_U3174) );
  AND2_X1 U19324 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n17343), .ZN(
        P1_U3173) );
  AND2_X1 U19325 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n17343), .ZN(
        P1_U3172) );
  AND2_X1 U19326 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n17343), .ZN(
        P1_U3171) );
  AND2_X1 U19327 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n17343), .ZN(
        P1_U3170) );
  AND2_X1 U19328 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n17343), .ZN(
        P1_U3169) );
  AND2_X1 U19329 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n17343), .ZN(
        P1_U3168) );
  AND2_X1 U19330 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n17343), .ZN(
        P1_U3167) );
  AND2_X1 U19331 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n17343), .ZN(
        P1_U3166) );
  AND2_X1 U19332 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n17343), .ZN(
        P1_U3165) );
  AND2_X1 U19333 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n17343), .ZN(
        P1_U3164) );
  OAI221_X1 U19334 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n15084), .C1(n21804), 
        .C2(n21841), .A(n22106), .ZN(n17383) );
  INV_X1 U19335 ( .A(n17344), .ZN(n17345) );
  NAND3_X1 U19336 ( .A1(n17347), .A2(n17346), .A3(n17345), .ZN(n17351) );
  OAI21_X1 U19337 ( .B1(n21834), .B2(n17349), .A(n17348), .ZN(n17350) );
  NAND2_X1 U19338 ( .A1(n17351), .A2(n17350), .ZN(n17382) );
  INV_X1 U19339 ( .A(n17352), .ZN(n17355) );
  INV_X1 U19340 ( .A(n17353), .ZN(n17354) );
  OAI211_X1 U19341 ( .C1(n12447), .C2(n17355), .A(n17354), .B(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n17361) );
  INV_X1 U19342 ( .A(n17356), .ZN(n17359) );
  INV_X1 U19343 ( .A(n17361), .ZN(n17357) );
  OAI22_X1 U19344 ( .A1(n17359), .A2(n17358), .B1(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n17357), .ZN(n17360) );
  OAI21_X1 U19345 ( .B1(n22066), .B2(n17361), .A(n17360), .ZN(n17362) );
  AOI222_X1 U19346 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n17363), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n17362), .C1(n17363), 
        .C2(n17362), .ZN(n17366) );
  OR2_X1 U19347 ( .A1(n17366), .A2(n17365), .ZN(n17364) );
  NAND2_X1 U19348 ( .A1(n17364), .A2(n22105), .ZN(n17368) );
  NAND2_X1 U19349 ( .A1(n17366), .A2(n17365), .ZN(n17367) );
  NAND2_X1 U19350 ( .A1(n17368), .A2(n17367), .ZN(n17369) );
  NAND2_X1 U19351 ( .A1(n17369), .A2(n17385), .ZN(n17379) );
  AND2_X1 U19352 ( .A1(n17370), .A2(n21790), .ZN(n17374) );
  INV_X1 U19353 ( .A(n17371), .ZN(n17373) );
  OAI211_X1 U19354 ( .C1(n17375), .C2(n17374), .A(n17373), .B(n17372), .ZN(
        n17376) );
  NOR2_X1 U19355 ( .A1(n17377), .A2(n17376), .ZN(n17378) );
  INV_X1 U19356 ( .A(n21814), .ZN(n17380) );
  AOI221_X1 U19357 ( .B1(n21804), .B2(n21798), .C1(n17380), .C2(n21798), .A(
        n17382), .ZN(n21806) );
  NOR2_X1 U19358 ( .A1(n21806), .A2(n21804), .ZN(n21805) );
  INV_X1 U19359 ( .A(n21511), .ZN(n21808) );
  NAND2_X1 U19360 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21808), .ZN(n17381) );
  OAI211_X1 U19361 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n21834), .A(n21805), 
        .B(n17381), .ZN(n21810) );
  OAI222_X1 U19362 ( .A1(n21798), .A2(n17383), .B1(n21798), .B2(n17382), .C1(
        P1_STATE2_REG_1__SCAN_IN), .C2(n21810), .ZN(P1_U3162) );
  NOR2_X1 U19363 ( .A1(n17385), .A2(n17384), .ZN(P1_U3032) );
  AND2_X1 U19364 ( .A1(n20034), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  INV_X1 U19365 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n17557) );
  AOI21_X1 U19366 ( .B1(n21835), .B2(n17557), .A(n22401), .ZN(P1_U2802) );
  NOR2_X1 U19367 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18944), .ZN(
        n18972) );
  NOR2_X1 U19368 ( .A1(n19173), .A2(n18475), .ZN(n18958) );
  AND2_X1 U19369 ( .A1(n21450), .A2(n18958), .ZN(n19002) );
  INV_X1 U19370 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21465) );
  NOR2_X1 U19371 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n21465), .ZN(
        n18959) );
  AOI22_X1 U19372 ( .A1(n19215), .A2(n18972), .B1(n19002), .B2(n18959), .ZN(
        n19297) );
  NAND2_X1 U19373 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18972), .ZN(
        n19300) );
  INV_X1 U19374 ( .A(n19300), .ZN(n19308) );
  NAND2_X1 U19375 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n19215), .ZN(n19123) );
  INV_X1 U19376 ( .A(n19123), .ZN(n19127) );
  INV_X1 U19377 ( .A(n18959), .ZN(n17386) );
  NOR2_X1 U19378 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n21488), .ZN(n20338) );
  INV_X1 U19379 ( .A(n20338), .ZN(n21479) );
  NAND2_X1 U19380 ( .A1(n21450), .A2(n21479), .ZN(n19000) );
  NOR2_X1 U19381 ( .A1(n17386), .A2(n19000), .ZN(n19295) );
  INV_X1 U19382 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n20843) );
  NOR2_X2 U19383 ( .A1(n20843), .A2(n19173), .ZN(n19126) );
  AOI22_X1 U19384 ( .A1(n19308), .A2(n19127), .B1(n19295), .B2(n19126), .ZN(
        n17387) );
  INV_X1 U19385 ( .A(n17387), .ZN(n17392) );
  NAND2_X1 U19386 ( .A1(n18972), .A2(n21449), .ZN(n19306) );
  NAND2_X1 U19387 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19215), .ZN(n19131) );
  NOR2_X1 U19388 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21449), .ZN(
        n18987) );
  NAND2_X1 U19389 ( .A1(n18959), .A2(n18987), .ZN(n19283) );
  NOR3_X1 U19390 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n17388), .A3(n21488), 
        .ZN(n19016) );
  NOR2_X2 U19391 ( .A1(n19261), .A2(n17389), .ZN(n19128) );
  INV_X1 U19392 ( .A(n19128), .ZN(n17390) );
  OAI22_X1 U19393 ( .A1(n19306), .A2(n19131), .B1(n19283), .B2(n17390), .ZN(
        n17391) );
  AOI211_X1 U19394 ( .C1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .C2(n19297), .A(
        n17392), .B(n17391), .ZN(n17601) );
  OAI22_X1 U19395 ( .A1(n20076), .A2(keyinput_62), .B1(keyinput_63), .B2(
        P1_REIP_REG_20__SCAN_IN), .ZN(n17393) );
  AOI221_X1 U19396 ( .B1(n20076), .B2(keyinput_62), .C1(
        P1_REIP_REG_20__SCAN_IN), .C2(keyinput_63), .A(n17393), .ZN(n17599) );
  INV_X1 U19397 ( .A(keyinput_61), .ZN(n17487) );
  INV_X1 U19398 ( .A(keyinput_60), .ZN(n17485) );
  INV_X1 U19399 ( .A(keyinput_59), .ZN(n17483) );
  INV_X1 U19400 ( .A(keyinput_58), .ZN(n17481) );
  INV_X1 U19401 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n20093) );
  INV_X1 U19402 ( .A(keyinput_53), .ZN(n17474) );
  OAI22_X1 U19403 ( .A1(n15084), .A2(keyinput_44), .B1(keyinput_45), .B2(
        P1_MORE_REG_SCAN_IN), .ZN(n17394) );
  AOI221_X1 U19404 ( .B1(n15084), .B2(keyinput_44), .C1(P1_MORE_REG_SCAN_IN), 
        .C2(keyinput_45), .A(n17394), .ZN(n17472) );
  INV_X1 U19405 ( .A(NA), .ZN(n21833) );
  INV_X1 U19406 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n20202) );
  OAI22_X1 U19407 ( .A1(n21833), .A2(keyinput_34), .B1(n20202), .B2(
        keyinput_40), .ZN(n17395) );
  AOI221_X1 U19408 ( .B1(n21833), .B2(keyinput_34), .C1(keyinput_40), .C2(
        n20202), .A(n17395), .ZN(n17462) );
  OAI22_X1 U19409 ( .A1(n22399), .A2(keyinput_41), .B1(keyinput_42), .B2(
        P1_D_C_N_REG_SCAN_IN), .ZN(n17396) );
  AOI221_X1 U19410 ( .B1(n22399), .B2(keyinput_41), .C1(P1_D_C_N_REG_SCAN_IN), 
        .C2(keyinput_42), .A(n17396), .ZN(n17461) );
  INV_X1 U19411 ( .A(READY2), .ZN(n17561) );
  AOI22_X1 U19412 ( .A1(n17556), .A2(keyinput_35), .B1(n17561), .B2(
        keyinput_37), .ZN(n17397) );
  OAI221_X1 U19413 ( .B1(n17556), .B2(keyinput_35), .C1(n17561), .C2(
        keyinput_37), .A(n17397), .ZN(n17405) );
  INV_X1 U19414 ( .A(READY1), .ZN(n17399) );
  AOI22_X1 U19415 ( .A1(n17557), .A2(keyinput_39), .B1(n17399), .B2(
        keyinput_36), .ZN(n17398) );
  OAI221_X1 U19416 ( .B1(n17557), .B2(keyinput_39), .C1(n17399), .C2(
        keyinput_36), .A(n17398), .ZN(n17404) );
  INV_X1 U19417 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n17402) );
  INV_X1 U19418 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n17401) );
  AOI22_X1 U19419 ( .A1(n17402), .A2(keyinput_43), .B1(keyinput_38), .B2(
        n17401), .ZN(n17400) );
  OAI221_X1 U19420 ( .B1(n17402), .B2(keyinput_43), .C1(n17401), .C2(
        keyinput_38), .A(n17400), .ZN(n17403) );
  NOR3_X1 U19421 ( .A1(n17405), .A2(n17404), .A3(n17403), .ZN(n17460) );
  INV_X1 U19422 ( .A(keyinput_26), .ZN(n17445) );
  INV_X1 U19423 ( .A(keyinput_25), .ZN(n17443) );
  INV_X1 U19424 ( .A(keyinput_24), .ZN(n17441) );
  INV_X1 U19425 ( .A(DATAI_8_), .ZN(n17538) );
  AOI22_X1 U19426 ( .A1(n17529), .A2(keyinput_20), .B1(n17525), .B2(
        keyinput_19), .ZN(n17406) );
  OAI221_X1 U19427 ( .B1(n17529), .B2(keyinput_20), .C1(n17525), .C2(
        keyinput_19), .A(n17406), .ZN(n17439) );
  INV_X1 U19428 ( .A(DATAI_10_), .ZN(n17528) );
  AOI22_X1 U19429 ( .A1(n17408), .A2(keyinput_23), .B1(n17528), .B2(
        keyinput_22), .ZN(n17407) );
  OAI221_X1 U19430 ( .B1(n17408), .B2(keyinput_23), .C1(n17528), .C2(
        keyinput_22), .A(n17407), .ZN(n17438) );
  AOI22_X1 U19431 ( .A1(n14747), .A2(keyinput_17), .B1(n17410), .B2(
        keyinput_18), .ZN(n17409) );
  OAI221_X1 U19432 ( .B1(n14747), .B2(keyinput_17), .C1(n17410), .C2(
        keyinput_18), .A(n17409), .ZN(n17436) );
  INV_X1 U19433 ( .A(keyinput_16), .ZN(n17433) );
  AOI22_X1 U19434 ( .A1(DATAI_18_), .A2(keyinput_14), .B1(DATAI_19_), .B2(
        keyinput_13), .ZN(n17411) );
  OAI221_X1 U19435 ( .B1(DATAI_18_), .B2(keyinput_14), .C1(DATAI_19_), .C2(
        keyinput_13), .A(n17411), .ZN(n17430) );
  OAI22_X1 U19436 ( .A1(DATAI_23_), .A2(keyinput_9), .B1(DATAI_22_), .B2(
        keyinput_10), .ZN(n17412) );
  AOI221_X1 U19437 ( .B1(DATAI_23_), .B2(keyinput_9), .C1(keyinput_10), .C2(
        DATAI_22_), .A(n17412), .ZN(n17428) );
  AOI22_X1 U19438 ( .A1(n17415), .A2(keyinput_2), .B1(keyinput_3), .B2(n17414), 
        .ZN(n17413) );
  OAI221_X1 U19439 ( .B1(n17415), .B2(keyinput_2), .C1(n17414), .C2(keyinput_3), .A(n17413), .ZN(n17424) );
  AOI22_X1 U19440 ( .A1(P1_MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_0), .B1(
        DATAI_31_), .B2(keyinput_1), .ZN(n17416) );
  OAI221_X1 U19441 ( .B1(P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_0), .C1(
        DATAI_31_), .C2(keyinput_1), .A(n17416), .ZN(n17423) );
  OAI22_X1 U19442 ( .A1(n17502), .A2(keyinput_7), .B1(DATAI_26_), .B2(
        keyinput_6), .ZN(n17417) );
  AOI221_X1 U19443 ( .B1(n17502), .B2(keyinput_7), .C1(keyinput_6), .C2(
        DATAI_26_), .A(n17417), .ZN(n17420) );
  OAI22_X1 U19444 ( .A1(DATAI_27_), .A2(keyinput_5), .B1(keyinput_8), .B2(
        DATAI_24_), .ZN(n17418) );
  AOI221_X1 U19445 ( .B1(DATAI_27_), .B2(keyinput_5), .C1(DATAI_24_), .C2(
        keyinput_8), .A(n17418), .ZN(n17419) );
  OAI211_X1 U19446 ( .C1(DATAI_28_), .C2(keyinput_4), .A(n17420), .B(n17419), 
        .ZN(n17421) );
  AOI21_X1 U19447 ( .B1(DATAI_28_), .B2(keyinput_4), .A(n17421), .ZN(n17422)
         );
  OAI21_X1 U19448 ( .B1(n17424), .B2(n17423), .A(n17422), .ZN(n17427) );
  AOI22_X1 U19449 ( .A1(DATAI_21_), .A2(keyinput_11), .B1(n17513), .B2(
        keyinput_12), .ZN(n17425) );
  OAI221_X1 U19450 ( .B1(DATAI_21_), .B2(keyinput_11), .C1(n17513), .C2(
        keyinput_12), .A(n17425), .ZN(n17426) );
  AOI21_X1 U19451 ( .B1(n17428), .B2(n17427), .A(n17426), .ZN(n17429) );
  OAI22_X1 U19452 ( .A1(n17430), .A2(n17429), .B1(keyinput_15), .B2(DATAI_17_), 
        .ZN(n17431) );
  AOI21_X1 U19453 ( .B1(keyinput_15), .B2(DATAI_17_), .A(n17431), .ZN(n17432)
         );
  AOI221_X1 U19454 ( .B1(DATAI_16_), .B2(n17433), .C1(n17522), .C2(keyinput_16), .A(n17432), .ZN(n17435) );
  NAND2_X1 U19455 ( .A1(keyinput_21), .A2(DATAI_11_), .ZN(n17434) );
  OAI221_X1 U19456 ( .B1(n17436), .B2(n17435), .C1(keyinput_21), .C2(DATAI_11_), .A(n17434), .ZN(n17437) );
  NOR3_X1 U19457 ( .A1(n17439), .A2(n17438), .A3(n17437), .ZN(n17440) );
  AOI221_X1 U19458 ( .B1(DATAI_8_), .B2(n17441), .C1(n17538), .C2(keyinput_24), 
        .A(n17440), .ZN(n17442) );
  AOI221_X1 U19459 ( .B1(DATAI_7_), .B2(n17443), .C1(n17541), .C2(keyinput_25), 
        .A(n17442), .ZN(n17444) );
  AOI221_X1 U19460 ( .B1(DATAI_6_), .B2(n17445), .C1(n17543), .C2(keyinput_26), 
        .A(n17444), .ZN(n17450) );
  OAI22_X1 U19461 ( .A1(n17447), .A2(keyinput_27), .B1(keyinput_29), .B2(
        DATAI_3_), .ZN(n17446) );
  AOI221_X1 U19462 ( .B1(n17447), .B2(keyinput_27), .C1(DATAI_3_), .C2(
        keyinput_29), .A(n17446), .ZN(n17448) );
  OAI21_X1 U19463 ( .B1(keyinput_28), .B2(n17550), .A(n17448), .ZN(n17449) );
  AOI211_X1 U19464 ( .C1(keyinput_28), .C2(n17550), .A(n17450), .B(n17449), 
        .ZN(n17458) );
  AOI22_X1 U19465 ( .A1(n17453), .A2(keyinput_31), .B1(n17452), .B2(
        keyinput_30), .ZN(n17451) );
  OAI221_X1 U19466 ( .B1(n17453), .B2(keyinput_31), .C1(n17452), .C2(
        keyinput_30), .A(n17451), .ZN(n17457) );
  OAI22_X1 U19467 ( .A1(n17455), .A2(keyinput_32), .B1(keyinput_33), .B2(HOLD), 
        .ZN(n17454) );
  AOI221_X1 U19468 ( .B1(n17455), .B2(keyinput_32), .C1(HOLD), .C2(keyinput_33), .A(n17454), .ZN(n17456) );
  OAI21_X1 U19469 ( .B1(n17458), .B2(n17457), .A(n17456), .ZN(n17459) );
  NAND4_X1 U19470 ( .A1(n17462), .A2(n17461), .A3(n17460), .A4(n17459), .ZN(
        n17471) );
  INV_X1 U19471 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20114) );
  AOI22_X1 U19472 ( .A1(n20091), .A2(keyinput_52), .B1(keyinput_49), .B2(
        n20114), .ZN(n17463) );
  OAI221_X1 U19473 ( .B1(n20091), .B2(keyinput_52), .C1(n20114), .C2(
        keyinput_49), .A(n17463), .ZN(n17470) );
  OAI22_X1 U19474 ( .A1(P1_BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput_51), .B1(
        keyinput_48), .B2(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n17464) );
  AOI221_X1 U19475 ( .B1(P1_BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_51), .C1(
        P1_BYTEENABLE_REG_0__SCAN_IN), .C2(keyinput_48), .A(n17464), .ZN(
        n17468) );
  INV_X1 U19476 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20110) );
  AOI22_X1 U19477 ( .A1(n20110), .A2(keyinput_50), .B1(n21790), .B2(
        keyinput_46), .ZN(n17465) );
  OAI221_X1 U19478 ( .B1(n20110), .B2(keyinput_50), .C1(n21790), .C2(
        keyinput_46), .A(n17465), .ZN(n17466) );
  AOI21_X1 U19479 ( .B1(keyinput_47), .B2(n20273), .A(n17466), .ZN(n17467) );
  OAI211_X1 U19480 ( .C1(keyinput_47), .C2(n20273), .A(n17468), .B(n17467), 
        .ZN(n17469) );
  AOI211_X1 U19481 ( .C1(n17472), .C2(n17471), .A(n17470), .B(n17469), .ZN(
        n17473) );
  AOI221_X1 U19482 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(keyinput_53), .C1(
        n20093), .C2(n17474), .A(n17473), .ZN(n17479) );
  AOI22_X1 U19483 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(keyinput_54), .B1(n13652), .B2(keyinput_55), .ZN(n17475) );
  OAI221_X1 U19484 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(keyinput_54), .C1(
        n13652), .C2(keyinput_55), .A(n17475), .ZN(n17478) );
  INV_X1 U19485 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20085) );
  OAI22_X1 U19486 ( .A1(n20085), .A2(keyinput_57), .B1(P1_REIP_REG_27__SCAN_IN), .B2(keyinput_56), .ZN(n17476) );
  AOI221_X1 U19487 ( .B1(n20085), .B2(keyinput_57), .C1(keyinput_56), .C2(
        P1_REIP_REG_27__SCAN_IN), .A(n17476), .ZN(n17477) );
  OAI21_X1 U19488 ( .B1(n17479), .B2(n17478), .A(n17477), .ZN(n17480) );
  OAI221_X1 U19489 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(n17481), .C1(n20082), 
        .C2(keyinput_58), .A(n17480), .ZN(n17482) );
  OAI221_X1 U19490 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(keyinput_59), .C1(
        n16118), .C2(n17483), .A(n17482), .ZN(n17484) );
  OAI221_X1 U19491 ( .B1(P1_REIP_REG_23__SCAN_IN), .B2(keyinput_60), .C1(
        n21599), .C2(n17485), .A(n17484), .ZN(n17486) );
  OAI221_X1 U19492 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(keyinput_61), .C1(
        n20078), .C2(n17487), .A(n17486), .ZN(n17598) );
  INV_X1 U19493 ( .A(keyinput_125), .ZN(n17594) );
  INV_X1 U19494 ( .A(keyinput_124), .ZN(n17592) );
  INV_X1 U19495 ( .A(keyinput_123), .ZN(n17590) );
  INV_X1 U19496 ( .A(keyinput_122), .ZN(n17588) );
  OAI22_X1 U19497 ( .A1(n20089), .A2(keyinput_118), .B1(n13652), .B2(
        keyinput_119), .ZN(n17488) );
  AOI221_X1 U19498 ( .B1(n20089), .B2(keyinput_118), .C1(keyinput_119), .C2(
        n13652), .A(n17488), .ZN(n17586) );
  INV_X1 U19499 ( .A(keyinput_117), .ZN(n17582) );
  OAI22_X1 U19500 ( .A1(DATAI_2_), .A2(keyinput_94), .B1(DATAI_1_), .B2(
        keyinput_95), .ZN(n17489) );
  AOI221_X1 U19501 ( .B1(DATAI_2_), .B2(keyinput_94), .C1(keyinput_95), .C2(
        DATAI_1_), .A(n17489), .ZN(n17554) );
  INV_X1 U19502 ( .A(keyinput_90), .ZN(n17544) );
  INV_X1 U19503 ( .A(keyinput_89), .ZN(n17540) );
  INV_X1 U19504 ( .A(keyinput_88), .ZN(n17537) );
  OAI22_X1 U19505 ( .A1(n14747), .A2(keyinput_81), .B1(keyinput_82), .B2(
        DATAI_14_), .ZN(n17490) );
  AOI221_X1 U19506 ( .B1(n14747), .B2(keyinput_81), .C1(DATAI_14_), .C2(
        keyinput_82), .A(n17490), .ZN(n17533) );
  INV_X1 U19507 ( .A(keyinput_80), .ZN(n17523) );
  AOI22_X1 U19508 ( .A1(DATAI_18_), .A2(keyinput_78), .B1(n17492), .B2(
        keyinput_77), .ZN(n17491) );
  OAI221_X1 U19509 ( .B1(DATAI_18_), .B2(keyinput_78), .C1(n17492), .C2(
        keyinput_77), .A(n17491), .ZN(n17520) );
  OAI22_X1 U19510 ( .A1(n17495), .A2(keyinput_73), .B1(n17494), .B2(
        keyinput_74), .ZN(n17493) );
  AOI221_X1 U19511 ( .B1(n17495), .B2(keyinput_73), .C1(keyinput_74), .C2(
        n17494), .A(n17493), .ZN(n17516) );
  OAI22_X1 U19512 ( .A1(DATAI_29_), .A2(keyinput_67), .B1(keyinput_64), .B2(
        P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n17496) );
  AOI221_X1 U19513 ( .B1(DATAI_29_), .B2(keyinput_67), .C1(
        P1_MEMORYFETCH_REG_SCAN_IN), .C2(keyinput_64), .A(n17496), .ZN(n17507)
         );
  OAI22_X1 U19514 ( .A1(DATAI_31_), .A2(keyinput_65), .B1(keyinput_66), .B2(
        DATAI_30_), .ZN(n17497) );
  AOI221_X1 U19515 ( .B1(DATAI_31_), .B2(keyinput_65), .C1(DATAI_30_), .C2(
        keyinput_66), .A(n17497), .ZN(n17506) );
  AOI22_X1 U19516 ( .A1(n17500), .A2(keyinput_69), .B1(n17499), .B2(
        keyinput_68), .ZN(n17498) );
  OAI221_X1 U19517 ( .B1(n17500), .B2(keyinput_69), .C1(n17499), .C2(
        keyinput_68), .A(n17498), .ZN(n17505) );
  AOI22_X1 U19518 ( .A1(n17503), .A2(keyinput_72), .B1(n17502), .B2(
        keyinput_71), .ZN(n17501) );
  OAI221_X1 U19519 ( .B1(n17503), .B2(keyinput_72), .C1(n17502), .C2(
        keyinput_71), .A(n17501), .ZN(n17504) );
  AOI211_X1 U19520 ( .C1(n17507), .C2(n17506), .A(n17505), .B(n17504), .ZN(
        n17509) );
  NAND2_X1 U19521 ( .A1(keyinput_70), .A2(n17510), .ZN(n17508) );
  OAI211_X1 U19522 ( .C1(keyinput_70), .C2(n17510), .A(n17509), .B(n17508), 
        .ZN(n17515) );
  AOI22_X1 U19523 ( .A1(n17513), .A2(keyinput_76), .B1(n17512), .B2(
        keyinput_75), .ZN(n17511) );
  OAI221_X1 U19524 ( .B1(n17513), .B2(keyinput_76), .C1(n17512), .C2(
        keyinput_75), .A(n17511), .ZN(n17514) );
  AOI21_X1 U19525 ( .B1(n17516), .B2(n17515), .A(n17514), .ZN(n17519) );
  NAND2_X1 U19526 ( .A1(n17518), .A2(keyinput_79), .ZN(n17517) );
  OAI221_X1 U19527 ( .B1(n17520), .B2(n17519), .C1(n17518), .C2(keyinput_79), 
        .A(n17517), .ZN(n17521) );
  OAI221_X1 U19528 ( .B1(DATAI_16_), .B2(n17523), .C1(n17522), .C2(keyinput_80), .A(n17521), .ZN(n17532) );
  AOI22_X1 U19529 ( .A1(n17526), .A2(keyinput_85), .B1(n17525), .B2(
        keyinput_83), .ZN(n17524) );
  OAI221_X1 U19530 ( .B1(n17526), .B2(keyinput_85), .C1(n17525), .C2(
        keyinput_83), .A(n17524), .ZN(n17531) );
  AOI22_X1 U19531 ( .A1(n17529), .A2(keyinput_84), .B1(keyinput_86), .B2(
        n17528), .ZN(n17527) );
  OAI221_X1 U19532 ( .B1(n17529), .B2(keyinput_84), .C1(n17528), .C2(
        keyinput_86), .A(n17527), .ZN(n17530) );
  AOI211_X1 U19533 ( .C1(n17533), .C2(n17532), .A(n17531), .B(n17530), .ZN(
        n17534) );
  OAI21_X1 U19534 ( .B1(DATAI_9_), .B2(keyinput_87), .A(n17534), .ZN(n17535)
         );
  AOI21_X1 U19535 ( .B1(DATAI_9_), .B2(keyinput_87), .A(n17535), .ZN(n17536)
         );
  AOI221_X1 U19536 ( .B1(DATAI_8_), .B2(keyinput_88), .C1(n17538), .C2(n17537), 
        .A(n17536), .ZN(n17539) );
  AOI221_X1 U19537 ( .B1(DATAI_7_), .B2(keyinput_89), .C1(n17541), .C2(n17540), 
        .A(n17539), .ZN(n17542) );
  AOI221_X1 U19538 ( .B1(DATAI_6_), .B2(n17544), .C1(n17543), .C2(keyinput_90), 
        .A(n17542), .ZN(n17548) );
  AOI22_X1 U19539 ( .A1(DATAI_5_), .A2(keyinput_91), .B1(n17546), .B2(
        keyinput_93), .ZN(n17545) );
  OAI221_X1 U19540 ( .B1(DATAI_5_), .B2(keyinput_91), .C1(n17546), .C2(
        keyinput_93), .A(n17545), .ZN(n17547) );
  AOI211_X1 U19541 ( .C1(n17550), .C2(keyinput_92), .A(n17548), .B(n17547), 
        .ZN(n17549) );
  OAI21_X1 U19542 ( .B1(n17550), .B2(keyinput_92), .A(n17549), .ZN(n17553) );
  AOI22_X1 U19543 ( .A1(HOLD), .A2(keyinput_97), .B1(DATAI_0_), .B2(
        keyinput_96), .ZN(n17551) );
  OAI221_X1 U19544 ( .B1(HOLD), .B2(keyinput_97), .C1(DATAI_0_), .C2(
        keyinput_96), .A(n17551), .ZN(n17552) );
  AOI21_X1 U19545 ( .B1(n17554), .B2(n17553), .A(n17552), .ZN(n17569) );
  AOI22_X1 U19546 ( .A1(n17557), .A2(keyinput_103), .B1(keyinput_99), .B2(
        n17556), .ZN(n17555) );
  OAI221_X1 U19547 ( .B1(n17557), .B2(keyinput_103), .C1(n17556), .C2(
        keyinput_99), .A(n17555), .ZN(n17568) );
  OAI22_X1 U19548 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(keyinput_104), .B1(
        P1_D_C_N_REG_SCAN_IN), .B2(keyinput_106), .ZN(n17558) );
  AOI221_X1 U19549 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_104), .C1(
        keyinput_106), .C2(P1_D_C_N_REG_SCAN_IN), .A(n17558), .ZN(n17566) );
  OAI22_X1 U19550 ( .A1(READY1), .A2(keyinput_100), .B1(keyinput_98), .B2(NA), 
        .ZN(n17559) );
  AOI221_X1 U19551 ( .B1(READY1), .B2(keyinput_100), .C1(NA), .C2(keyinput_98), 
        .A(n17559), .ZN(n17565) );
  OAI22_X1 U19552 ( .A1(n17561), .A2(keyinput_101), .B1(keyinput_102), .B2(
        P1_READREQUEST_REG_SCAN_IN), .ZN(n17560) );
  AOI221_X1 U19553 ( .B1(n17561), .B2(keyinput_101), .C1(
        P1_READREQUEST_REG_SCAN_IN), .C2(keyinput_102), .A(n17560), .ZN(n17564) );
  OAI22_X1 U19554 ( .A1(n22399), .A2(keyinput_105), .B1(
        P1_REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_107), .ZN(n17562) );
  AOI221_X1 U19555 ( .B1(n22399), .B2(keyinput_105), .C1(keyinput_107), .C2(
        P1_REQUESTPENDING_REG_SCAN_IN), .A(n17562), .ZN(n17563) );
  NAND4_X1 U19556 ( .A1(n17566), .A2(n17565), .A3(n17564), .A4(n17563), .ZN(
        n17567) );
  NOR3_X1 U19557 ( .A1(n17569), .A2(n17568), .A3(n17567), .ZN(n17580) );
  AOI22_X1 U19558 ( .A1(P1_MORE_REG_SCAN_IN), .A2(keyinput_109), .B1(n15084), 
        .B2(keyinput_108), .ZN(n17570) );
  OAI221_X1 U19559 ( .B1(P1_MORE_REG_SCAN_IN), .B2(keyinput_109), .C1(n15084), 
        .C2(keyinput_108), .A(n17570), .ZN(n17579) );
  OAI22_X1 U19560 ( .A1(n20091), .A2(keyinput_116), .B1(n20273), .B2(
        keyinput_111), .ZN(n17571) );
  AOI221_X1 U19561 ( .B1(n20091), .B2(keyinput_116), .C1(keyinput_111), .C2(
        n20273), .A(n17571), .ZN(n17578) );
  OAI22_X1 U19562 ( .A1(n20110), .A2(keyinput_114), .B1(
        P1_BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_113), .ZN(n17572) );
  AOI221_X1 U19563 ( .B1(n20110), .B2(keyinput_114), .C1(keyinput_113), .C2(
        P1_BYTEENABLE_REG_1__SCAN_IN), .A(n17572), .ZN(n17575) );
  INV_X1 U19564 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20095) );
  INV_X1 U19565 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20117) );
  OAI22_X1 U19566 ( .A1(n20095), .A2(keyinput_115), .B1(n20117), .B2(
        keyinput_112), .ZN(n17573) );
  AOI221_X1 U19567 ( .B1(n20095), .B2(keyinput_115), .C1(keyinput_112), .C2(
        n20117), .A(n17573), .ZN(n17574) );
  OAI211_X1 U19568 ( .C1(P1_FLUSH_REG_SCAN_IN), .C2(keyinput_110), .A(n17575), 
        .B(n17574), .ZN(n17576) );
  AOI21_X1 U19569 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(keyinput_110), .A(n17576), 
        .ZN(n17577) );
  OAI211_X1 U19570 ( .C1(n17580), .C2(n17579), .A(n17578), .B(n17577), .ZN(
        n17581) );
  OAI221_X1 U19571 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n17582), .C1(n20093), 
        .C2(keyinput_117), .A(n17581), .ZN(n17585) );
  AOI22_X1 U19572 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(keyinput_120), .B1(
        n20085), .B2(keyinput_121), .ZN(n17583) );
  OAI221_X1 U19573 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(keyinput_120), .C1(
        n20085), .C2(keyinput_121), .A(n17583), .ZN(n17584) );
  AOI21_X1 U19574 ( .B1(n17586), .B2(n17585), .A(n17584), .ZN(n17587) );
  AOI221_X1 U19575 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(n17588), .C1(n20082), 
        .C2(keyinput_122), .A(n17587), .ZN(n17589) );
  AOI221_X1 U19576 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n17590), .C1(n16118), 
        .C2(keyinput_123), .A(n17589), .ZN(n17591) );
  AOI221_X1 U19577 ( .B1(P1_REIP_REG_23__SCAN_IN), .B2(keyinput_124), .C1(
        n21599), .C2(n17592), .A(n17591), .ZN(n17593) );
  AOI221_X1 U19578 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(n17594), .C1(n20078), 
        .C2(keyinput_125), .A(n17593), .ZN(n17597) );
  AOI22_X1 U19579 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(keyinput_127), .B1(
        n20076), .B2(keyinput_126), .ZN(n17595) );
  OAI221_X1 U19580 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(keyinput_127), .C1(
        n20076), .C2(keyinput_126), .A(n17595), .ZN(n17596) );
  AOI211_X1 U19581 ( .C1(n17599), .C2(n17598), .A(n17597), .B(n17596), .ZN(
        n17600) );
  XNOR2_X1 U19582 ( .A(n17601), .B(n17600), .ZN(P3_U2944) );
  INV_X1 U19583 ( .A(n18589), .ZN(n17604) );
  INV_X1 U19584 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n17603) );
  OAI22_X1 U19585 ( .A1(n17604), .A2(n17603), .B1(n11407), .B2(n17602), .ZN(
        P2_U2816) );
  INV_X1 U19586 ( .A(n17605), .ZN(n17607) );
  AOI22_X1 U19587 ( .A1(n17607), .A2(n17668), .B1(n17617), .B2(n17606), .ZN(
        n17613) );
  NAND2_X1 U19588 ( .A1(n17661), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n17608) );
  OAI211_X1 U19589 ( .C1(n17631), .C2(n17610), .A(n17609), .B(n17608), .ZN(
        n17611) );
  AOI21_X1 U19590 ( .B1(n14791), .B2(n17672), .A(n17611), .ZN(n17612) );
  NAND2_X1 U19591 ( .A1(n17613), .A2(n17612), .ZN(P2_U3012) );
  INV_X1 U19592 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n17745) );
  OAI22_X1 U19593 ( .A1(n17745), .A2(n18746), .B1(n17631), .B2(n17614), .ZN(
        n17615) );
  AOI21_X1 U19594 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17661), .A(
        n17615), .ZN(n17620) );
  AOI22_X1 U19595 ( .A1(n17618), .A2(n17617), .B1(n17668), .B2(n17616), .ZN(
        n17619) );
  OAI211_X1 U19596 ( .C1(n17651), .C2(n17621), .A(n17620), .B(n17619), .ZN(
        P2_U3010) );
  OAI22_X1 U19597 ( .A1(n17622), .A2(n17658), .B1(n17746), .B2(n18746), .ZN(
        n17623) );
  AOI21_X1 U19598 ( .B1(n17647), .B2(n17624), .A(n17623), .ZN(n17629) );
  OAI22_X1 U19599 ( .A1(n17626), .A2(n17648), .B1(n17625), .B2(n17670), .ZN(
        n17627) );
  INV_X1 U19600 ( .A(n17627), .ZN(n17628) );
  OAI211_X1 U19601 ( .C1(n17651), .C2(n17630), .A(n17629), .B(n17628), .ZN(
        P2_U3009) );
  OAI22_X1 U19602 ( .A1(n18626), .A2(n18746), .B1(n17631), .B2(n18620), .ZN(
        n17632) );
  AOI21_X1 U19603 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17661), .A(
        n17632), .ZN(n17637) );
  OAI22_X1 U19604 ( .A1(n17634), .A2(n17648), .B1(n17670), .B2(n17633), .ZN(
        n17635) );
  INV_X1 U19605 ( .A(n17635), .ZN(n17636) );
  OAI211_X1 U19606 ( .C1(n17651), .C2(n18627), .A(n17637), .B(n17636), .ZN(
        P2_U3008) );
  AOI22_X1 U19607 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n16976), .B1(n17647), 
        .B2(n18634), .ZN(n17644) );
  NOR2_X1 U19608 ( .A1(n17638), .A2(n17648), .ZN(n17642) );
  OAI22_X1 U19609 ( .A1(n17639), .A2(n17670), .B1(n17651), .B2(n18639), .ZN(
        n17640) );
  AOI21_X1 U19610 ( .B1(n17642), .B2(n17641), .A(n17640), .ZN(n17643) );
  OAI211_X1 U19611 ( .C1(n17645), .C2(n17658), .A(n17644), .B(n17643), .ZN(
        P2_U3007) );
  AOI22_X1 U19612 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n16976), .B1(n17647), 
        .B2(n17646), .ZN(n17657) );
  NOR2_X1 U19613 ( .A1(n17649), .A2(n17648), .ZN(n17655) );
  OAI22_X1 U19614 ( .A1(n17652), .A2(n17670), .B1(n17651), .B2(n17650), .ZN(
        n17653) );
  AOI21_X1 U19615 ( .B1(n17655), .B2(n17654), .A(n17653), .ZN(n17656) );
  OAI211_X1 U19616 ( .C1(n17659), .C2(n17658), .A(n17657), .B(n17656), .ZN(
        P2_U3005) );
  NOR2_X1 U19617 ( .A1(n17661), .A2(n17660), .ZN(n17674) );
  NAND2_X1 U19618 ( .A1(n18598), .A2(n17662), .ZN(n17663) );
  NAND2_X1 U19619 ( .A1(n17664), .A2(n17663), .ZN(n18882) );
  OAI21_X1 U19620 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n17666), .A(
        n17665), .ZN(n17667) );
  INV_X1 U19621 ( .A(n17667), .ZN(n18878) );
  NAND2_X1 U19622 ( .A1(n17668), .A2(n18878), .ZN(n17669) );
  NAND2_X1 U19623 ( .A1(n16976), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n18883) );
  OAI211_X1 U19624 ( .C1(n18882), .C2(n17670), .A(n17669), .B(n18883), .ZN(
        n17671) );
  AOI21_X1 U19625 ( .B1(n18600), .B2(n17672), .A(n17671), .ZN(n17673) );
  OAI21_X1 U19626 ( .B1(n17674), .B2(n18601), .A(n17673), .ZN(P2_U3014) );
  INV_X1 U19627 ( .A(n17675), .ZN(n17677) );
  OAI22_X1 U19628 ( .A1(n19455), .A2(n18591), .B1(n17677), .B2(n17676), .ZN(
        n17678) );
  AOI21_X1 U19629 ( .B1(n19424), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n17678), 
        .ZN(n17679) );
  OAI22_X1 U19630 ( .A1(n19424), .A2(n17688), .B1(n17696), .B2(n17679), .ZN(
        P2_U3605) );
  NOR2_X1 U19631 ( .A1(n19408), .A2(n21819), .ZN(n17680) );
  OR2_X1 U19632 ( .A1(n17680), .A2(n19549), .ZN(n17684) );
  NAND2_X1 U19633 ( .A1(n18892), .A2(n17684), .ZN(n17691) );
  NAND2_X1 U19634 ( .A1(n17692), .A2(n17680), .ZN(n19522) );
  INV_X1 U19635 ( .A(n19522), .ZN(n17681) );
  AOI222_X1 U19636 ( .A1(n17682), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n19502), 
        .B2(n17691), .C1(n19564), .C2(n17681), .ZN(n17683) );
  AOI22_X1 U19637 ( .A1(n17696), .A2(n19518), .B1(n17683), .B2(n17688), .ZN(
        P2_U3603) );
  AND2_X1 U19638 ( .A1(n17684), .A2(n18892), .ZN(n17685) );
  OAI22_X1 U19639 ( .A1(n17685), .A2(n19408), .B1(n21819), .B2(n17684), .ZN(
        n17686) );
  AOI21_X1 U19640 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n17687), .A(n17686), 
        .ZN(n17689) );
  AOI22_X1 U19641 ( .A1(n17696), .A2(n19523), .B1(n17689), .B2(n17688), .ZN(
        P2_U3604) );
  AOI22_X1 U19642 ( .A1(n19521), .A2(n17691), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n17690), .ZN(n17695) );
  AOI211_X1 U19643 ( .C1(n19445), .C2(n19473), .A(n21819), .B(n19549), .ZN(
        n17693) );
  NOR2_X1 U19644 ( .A1(n17696), .A2(n17693), .ZN(n17694) );
  AOI22_X1 U19645 ( .A1(n14101), .A2(n17696), .B1(n17695), .B2(n17694), .ZN(
        P2_U3602) );
  NAND2_X1 U19646 ( .A1(n17697), .A2(n21821), .ZN(n17701) );
  INV_X1 U19647 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n17742) );
  OAI21_X1 U19648 ( .B1(n17698), .B2(n17742), .A(n17704), .ZN(n17699) );
  OAI21_X1 U19649 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n17704), .A(n17699), 
        .ZN(n17700) );
  OAI221_X1 U19650 ( .B1(n17701), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n17701), .C2(P2_REIP_REG_0__SCAN_IN), .A(n17700), .ZN(P2_U2822) );
  INV_X1 U19651 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17772) );
  OAI221_X1 U19652 ( .B1(n17704), .B2(n17772), .C1(n17703), .C2(n17702), .A(
        n17701), .ZN(P2_U2823) );
  INV_X1 U19653 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n17705) );
  AOI22_X1 U19654 ( .A1(n21855), .A2(n17706), .B1(n17705), .B2(n17770), .ZN(
        P2_U3611) );
  INV_X1 U19655 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n17707) );
  AOI22_X1 U19656 ( .A1(n21855), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n17707), 
        .B2(n17770), .ZN(P2_U3608) );
  INV_X1 U19657 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n21867) );
  INV_X1 U19658 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n17709) );
  OAI21_X1 U19659 ( .B1(n21867), .B2(n17709), .A(n17708), .ZN(P2_U2815) );
  AOI22_X1 U19660 ( .A1(n17736), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n17735), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n17711) );
  OAI21_X1 U19661 ( .B1(n11977), .B2(n17738), .A(n17711), .ZN(P2_U2951) );
  INV_X1 U19662 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n17713) );
  AOI22_X1 U19663 ( .A1(n17736), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n17735), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n17712) );
  OAI21_X1 U19664 ( .B1(n17713), .B2(n17738), .A(n17712), .ZN(P2_U2950) );
  AOI22_X1 U19665 ( .A1(n17736), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n17721), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n17714) );
  OAI21_X1 U19666 ( .B1(n15367), .B2(n17738), .A(n17714), .ZN(P2_U2949) );
  INV_X1 U19667 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n17716) );
  AOI22_X1 U19668 ( .A1(n17727), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n17721), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n17715) );
  OAI21_X1 U19669 ( .B1(n17716), .B2(n17738), .A(n17715), .ZN(P2_U2948) );
  INV_X1 U19670 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n17718) );
  AOI22_X1 U19671 ( .A1(n17736), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n17721), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n17717) );
  OAI21_X1 U19672 ( .B1(n17718), .B2(n17738), .A(n17717), .ZN(P2_U2947) );
  INV_X1 U19673 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n17720) );
  AOI22_X1 U19674 ( .A1(n17727), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n17721), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n17719) );
  OAI21_X1 U19675 ( .B1(n17720), .B2(n17738), .A(n17719), .ZN(P2_U2946) );
  AOI22_X1 U19676 ( .A1(n17727), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n17721), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n17722) );
  OAI21_X1 U19677 ( .B1(n14659), .B2(n17738), .A(n17722), .ZN(P2_U2945) );
  AOI22_X1 U19678 ( .A1(n17727), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n17735), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n17723) );
  OAI21_X1 U19679 ( .B1(n17724), .B2(n17738), .A(n17723), .ZN(P2_U2944) );
  AOI22_X1 U19680 ( .A1(n17727), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n17735), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n17725) );
  OAI21_X1 U19681 ( .B1(n14689), .B2(n17738), .A(n17725), .ZN(P2_U2943) );
  AOI22_X1 U19682 ( .A1(n17736), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n17735), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n17726) );
  OAI21_X1 U19683 ( .B1(n19373), .B2(n17738), .A(n17726), .ZN(P2_U2942) );
  AOI22_X1 U19684 ( .A1(n17727), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n17735), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n17728) );
  OAI21_X1 U19685 ( .B1(n14685), .B2(n17738), .A(n17728), .ZN(P2_U2941) );
  AOI22_X1 U19686 ( .A1(n17736), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n17735), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n17729) );
  OAI21_X1 U19687 ( .B1(n17730), .B2(n17738), .A(n17729), .ZN(P2_U2940) );
  AOI22_X1 U19688 ( .A1(n17736), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n17735), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n17731) );
  OAI21_X1 U19689 ( .B1(n14657), .B2(n17738), .A(n17731), .ZN(P2_U2939) );
  AOI22_X1 U19690 ( .A1(n17736), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n17735), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n17732) );
  OAI21_X1 U19691 ( .B1(n14652), .B2(n17738), .A(n17732), .ZN(P2_U2938) );
  AOI22_X1 U19692 ( .A1(n17736), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n17735), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n17733) );
  OAI21_X1 U19693 ( .B1(n17734), .B2(n17738), .A(n17733), .ZN(P2_U2937) );
  AOI22_X1 U19694 ( .A1(n17736), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n17735), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n17737) );
  OAI21_X1 U19695 ( .B1(n17739), .B2(n17738), .A(n17737), .ZN(P2_U2936) );
  AOI21_X1 U19696 ( .B1(n21867), .B2(n17740), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n17741) );
  AOI21_X1 U19697 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n21855), .A(n17741), 
        .ZN(P2_U2817) );
  INV_X1 U19698 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n17743) );
  OAI222_X1 U19699 ( .A1(n17762), .A2(n17742), .B1(n19954), .B2(n21855), .C1(
        n17743), .C2(n17765), .ZN(P2_U3212) );
  INV_X1 U19700 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19956) );
  OAI222_X1 U19701 ( .A1(n17762), .A2(n17743), .B1(n19956), .B2(n21855), .C1(
        n17744), .C2(n17765), .ZN(P2_U3213) );
  INV_X1 U19702 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19958) );
  OAI222_X1 U19703 ( .A1(n17762), .A2(n17744), .B1(n19958), .B2(n21855), .C1(
        n17745), .C2(n17765), .ZN(P2_U3214) );
  INV_X1 U19704 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19960) );
  OAI222_X1 U19705 ( .A1(n17765), .A2(n17746), .B1(n19960), .B2(n21855), .C1(
        n17745), .C2(n17762), .ZN(P2_U3215) );
  INV_X1 U19706 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19962) );
  OAI222_X1 U19707 ( .A1(n17765), .A2(n18626), .B1(n19962), .B2(n21855), .C1(
        n17746), .C2(n17762), .ZN(P2_U3216) );
  INV_X1 U19708 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19964) );
  OAI222_X1 U19709 ( .A1(n17765), .A2(n18638), .B1(n19964), .B2(n21855), .C1(
        n18626), .C2(n17762), .ZN(P2_U3217) );
  INV_X1 U19710 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19966) );
  OAI222_X1 U19711 ( .A1(n17765), .A2(n18647), .B1(n19966), .B2(n21855), .C1(
        n18638), .C2(n17762), .ZN(P2_U3218) );
  INV_X1 U19712 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n17747) );
  INV_X1 U19713 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19968) );
  OAI222_X1 U19714 ( .A1(n17765), .A2(n17747), .B1(n19968), .B2(n21855), .C1(
        n18647), .C2(n17762), .ZN(P2_U3219) );
  INV_X1 U19715 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19970) );
  INV_X1 U19716 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n18660) );
  OAI222_X1 U19717 ( .A1(n17762), .A2(n17747), .B1(n19970), .B2(n21855), .C1(
        n18660), .C2(n17765), .ZN(P2_U3220) );
  INV_X1 U19718 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19972) );
  OAI222_X1 U19719 ( .A1(n17762), .A2(n18660), .B1(n19972), .B2(n21855), .C1(
        n16969), .C2(n17765), .ZN(P2_U3221) );
  INV_X1 U19720 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19974) );
  INV_X1 U19721 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n17748) );
  OAI222_X1 U19722 ( .A1(n17762), .A2(n16969), .B1(n19974), .B2(n21855), .C1(
        n17748), .C2(n17765), .ZN(P2_U3222) );
  INV_X1 U19723 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19976) );
  INV_X1 U19724 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n17749) );
  OAI222_X1 U19725 ( .A1(n17762), .A2(n17748), .B1(n19976), .B2(n21855), .C1(
        n17749), .C2(n17765), .ZN(P2_U3223) );
  INV_X1 U19726 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19978) );
  INV_X1 U19727 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n17750) );
  OAI222_X1 U19728 ( .A1(n17762), .A2(n17749), .B1(n19978), .B2(n21855), .C1(
        n17750), .C2(n17765), .ZN(P2_U3224) );
  INV_X1 U19729 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19980) );
  INV_X1 U19730 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n17751) );
  OAI222_X1 U19731 ( .A1(n17762), .A2(n17750), .B1(n19980), .B2(n21855), .C1(
        n17751), .C2(n17765), .ZN(P2_U3225) );
  INV_X1 U19732 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19982) );
  INV_X1 U19733 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n18706) );
  OAI222_X1 U19734 ( .A1(n17762), .A2(n17751), .B1(n19982), .B2(n21855), .C1(
        n18706), .C2(n17765), .ZN(P2_U3226) );
  INV_X1 U19735 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19984) );
  INV_X1 U19736 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n17752) );
  OAI222_X1 U19737 ( .A1(n17762), .A2(n18706), .B1(n19984), .B2(n21855), .C1(
        n17752), .C2(n17765), .ZN(P2_U3227) );
  INV_X1 U19738 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19986) );
  OAI222_X1 U19739 ( .A1(n17762), .A2(n17752), .B1(n19986), .B2(n21855), .C1(
        n18732), .C2(n17765), .ZN(P2_U3228) );
  INV_X1 U19740 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n18749) );
  INV_X1 U19741 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19988) );
  OAI222_X1 U19742 ( .A1(n17765), .A2(n18749), .B1(n19988), .B2(n21855), .C1(
        n18732), .C2(n17762), .ZN(P2_U3229) );
  INV_X1 U19743 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19990) );
  OAI222_X1 U19744 ( .A1(n17762), .A2(n18749), .B1(n19990), .B2(n21855), .C1(
        n17753), .C2(n17765), .ZN(P2_U3230) );
  INV_X1 U19745 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19992) );
  OAI222_X1 U19746 ( .A1(n17765), .A2(n16869), .B1(n19992), .B2(n21855), .C1(
        n17753), .C2(n17762), .ZN(P2_U3231) );
  INV_X1 U19747 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19994) );
  OAI222_X1 U19748 ( .A1(n17765), .A2(n17754), .B1(n19994), .B2(n21855), .C1(
        n16869), .C2(n17762), .ZN(P2_U3232) );
  INV_X1 U19749 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19996) );
  OAI222_X1 U19750 ( .A1(n17765), .A2(n17755), .B1(n19996), .B2(n21855), .C1(
        n17754), .C2(n17762), .ZN(P2_U3233) );
  INV_X1 U19751 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n17756) );
  INV_X1 U19752 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19998) );
  OAI222_X1 U19753 ( .A1(n17765), .A2(n17756), .B1(n19998), .B2(n21855), .C1(
        n17755), .C2(n17762), .ZN(P2_U3234) );
  INV_X1 U19754 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n17757) );
  INV_X1 U19755 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20000) );
  OAI222_X1 U19756 ( .A1(n17765), .A2(n17757), .B1(n20000), .B2(n21855), .C1(
        n17756), .C2(n17762), .ZN(P2_U3235) );
  INV_X1 U19757 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20003) );
  OAI222_X1 U19758 ( .A1(n17762), .A2(n17757), .B1(n20003), .B2(n21855), .C1(
        n17758), .C2(n17765), .ZN(P2_U3236) );
  INV_X1 U19759 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20005) );
  OAI222_X1 U19760 ( .A1(n17765), .A2(n17759), .B1(n20005), .B2(n21855), .C1(
        n17758), .C2(n17762), .ZN(P2_U3237) );
  INV_X1 U19761 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20007) );
  OAI222_X1 U19762 ( .A1(n17762), .A2(n17759), .B1(n20007), .B2(n21855), .C1(
        n17760), .C2(n17765), .ZN(P2_U3238) );
  INV_X1 U19763 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20009) );
  OAI222_X1 U19764 ( .A1(n17762), .A2(n17760), .B1(n20009), .B2(n21855), .C1(
        n17761), .C2(n17765), .ZN(P2_U3239) );
  INV_X1 U19765 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20011) );
  OAI222_X1 U19766 ( .A1(n17762), .A2(n17761), .B1(n20011), .B2(n21855), .C1(
        n17763), .C2(n17765), .ZN(P2_U3240) );
  INV_X1 U19767 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20014) );
  OAI222_X1 U19768 ( .A1(n17765), .A2(n17764), .B1(n20014), .B2(n21855), .C1(
        n17763), .C2(n17762), .ZN(P2_U3241) );
  INV_X1 U19769 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n17766) );
  AOI22_X1 U19770 ( .A1(n21855), .A2(n17767), .B1(n17766), .B2(n17770), .ZN(
        P2_U3588) );
  INV_X1 U19771 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n17768) );
  AOI22_X1 U19772 ( .A1(n21855), .A2(n17769), .B1(n17768), .B2(n17770), .ZN(
        P2_U3587) );
  MUX2_X1 U19773 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n21855), .Z(P2_U3586) );
  INV_X1 U19774 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n17771) );
  AOI22_X1 U19775 ( .A1(n21855), .A2(n17772), .B1(n17771), .B2(n17770), .ZN(
        P2_U3585) );
  NOR2_X1 U19776 ( .A1(n18072), .A2(n17795), .ZN(n17776) );
  AOI22_X1 U19777 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n18043), .B1(n18067), .B2(
        n17773), .ZN(n17775) );
  INV_X1 U19778 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17774) );
  OAI22_X1 U19779 ( .A1(n17776), .A2(n17775), .B1(n17774), .B2(n18043), .ZN(
        P3_U2699) );
  NAND4_X1 U19780 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .A4(n18067), .ZN(n17780) );
  NAND3_X1 U19781 ( .A1(n17780), .A2(P3_EBX_REG_3__SCAN_IN), .A3(n18043), .ZN(
        n17777) );
  OAI221_X1 U19782 ( .B1(n17780), .B2(P3_EBX_REG_3__SCAN_IN), .C1(n18043), 
        .C2(n17778), .A(n17777), .ZN(P3_U2700) );
  INV_X1 U19783 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17783) );
  NAND2_X1 U19784 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17779) );
  NOR2_X1 U19785 ( .A1(n18069), .A2(n17779), .ZN(n17781) );
  OAI211_X1 U19786 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17781), .A(n17780), .B(
        n18043), .ZN(n17782) );
  OAI21_X1 U19787 ( .B1(n18043), .B2(n17783), .A(n17782), .ZN(P3_U2701) );
  AOI22_X1 U19788 ( .A1(n11010), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18056), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17794) );
  AOI22_X1 U19789 ( .A1(n18033), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17793) );
  AOI22_X1 U19790 ( .A1(n13919), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18045), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17784) );
  OAI21_X1 U19791 ( .B1(n17850), .B2(n17785), .A(n17784), .ZN(n17791) );
  AOI22_X1 U19792 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17789) );
  AOI22_X1 U19793 ( .A1(n17920), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18047), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17788) );
  AOI22_X1 U19794 ( .A1(n20370), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10956), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17787) );
  AOI22_X1 U19795 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17865), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17786) );
  NAND4_X1 U19796 ( .A1(n17789), .A2(n17788), .A3(n17787), .A4(n17786), .ZN(
        n17790) );
  AOI211_X1 U19797 ( .C1(n17991), .C2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n17791), .B(n17790), .ZN(n17792) );
  NAND3_X1 U19798 ( .A1(n17794), .A2(n17793), .A3(n17792), .ZN(n20972) );
  INV_X1 U19799 ( .A(n20972), .ZN(n17798) );
  NOR2_X1 U19800 ( .A1(n18069), .A2(n17795), .ZN(n17803) );
  AND3_X1 U19801 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .A3(n17803), .ZN(n17799) );
  NAND2_X1 U19802 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n17799), .ZN(n17916) );
  INV_X1 U19803 ( .A(n17916), .ZN(n17796) );
  INV_X1 U19804 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n20443) );
  AOI22_X1 U19805 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17916), .B1(n17796), .B2(
        n20443), .ZN(n17797) );
  AOI22_X1 U19806 ( .A1(n18070), .A2(n17798), .B1(n17797), .B2(n18043), .ZN(
        P3_U2695) );
  OAI21_X1 U19807 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17799), .A(n17916), .ZN(
        n17800) );
  AOI22_X1 U19808 ( .A1(n18070), .A2(n17818), .B1(n17800), .B2(n18043), .ZN(
        P3_U2696) );
  NAND3_X1 U19809 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n18067), .A3(n17864), .ZN(
        n17802) );
  INV_X1 U19810 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17983) );
  NAND3_X1 U19811 ( .A1(n17802), .A2(P3_EBX_REG_6__SCAN_IN), .A3(n18043), .ZN(
        n17801) );
  OAI221_X1 U19812 ( .B1(n17802), .B2(P3_EBX_REG_6__SCAN_IN), .C1(n18043), 
        .C2(n17983), .A(n17801), .ZN(P3_U2697) );
  OAI211_X1 U19813 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n17803), .A(n17802), .B(
        n18043), .ZN(n17804) );
  OAI21_X1 U19814 ( .B1(n18043), .B2(n17835), .A(n17804), .ZN(P3_U2698) );
  NAND2_X1 U19815 ( .A1(n18067), .A2(n17805), .ZN(n17830) );
  AOI22_X1 U19816 ( .A1(n17909), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17809) );
  AOI22_X1 U19817 ( .A1(n17920), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18056), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17808) );
  AOI22_X1 U19818 ( .A1(n20370), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10956), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17807) );
  AOI22_X1 U19819 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17865), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17806) );
  NAND4_X1 U19820 ( .A1(n17809), .A2(n17808), .A3(n17807), .A4(n17806), .ZN(
        n17815) );
  AOI22_X1 U19821 ( .A1(n18045), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17813) );
  AOI22_X1 U19822 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17890), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17812) );
  AOI22_X1 U19823 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18047), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17811) );
  AOI22_X1 U19824 ( .A1(n11010), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n18046), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17810) );
  NAND4_X1 U19825 ( .A1(n17813), .A2(n17812), .A3(n17811), .A4(n17810), .ZN(
        n17814) );
  NOR2_X1 U19826 ( .A1(n17815), .A2(n17814), .ZN(n20956) );
  NAND3_X1 U19827 ( .A1(n17830), .A2(P3_EBX_REG_16__SCAN_IN), .A3(n18043), 
        .ZN(n17816) );
  OAI221_X1 U19828 ( .B1(n17830), .B2(P3_EBX_REG_16__SCAN_IN), .C1(n18043), 
        .C2(n20956), .A(n17816), .ZN(P3_U2687) );
  AOI22_X1 U19829 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17890), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17827) );
  AOI22_X1 U19830 ( .A1(n17920), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n18047), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17826) );
  AOI22_X1 U19831 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18046), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17817) );
  OAI21_X1 U19832 ( .B1(n17850), .B2(n17818), .A(n17817), .ZN(n17824) );
  AOI22_X1 U19833 ( .A1(n18045), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17822) );
  AOI22_X1 U19834 ( .A1(n10971), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18056), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17821) );
  AOI22_X1 U19835 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17865), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17820) );
  AOI22_X1 U19836 ( .A1(n18025), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10956), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17819) );
  NAND4_X1 U19837 ( .A1(n17822), .A2(n17821), .A3(n17820), .A4(n17819), .ZN(
        n17823) );
  AOI211_X1 U19838 ( .C1(n10967), .C2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n17824), .B(n17823), .ZN(n17825) );
  NAND3_X1 U19839 ( .A1(n17827), .A2(n17826), .A3(n17825), .ZN(n20964) );
  INV_X1 U19840 ( .A(n20964), .ZN(n17833) );
  NOR2_X1 U19841 ( .A1(n20518), .A2(n20510), .ZN(n17829) );
  NOR2_X1 U19842 ( .A1(n18069), .A2(n17828), .ZN(n17848) );
  AOI21_X1 U19843 ( .B1(n17829), .B2(n17848), .A(P3_EBX_REG_15__SCAN_IN), .ZN(
        n17832) );
  NAND2_X1 U19844 ( .A1(n18043), .A2(n17830), .ZN(n17831) );
  OAI22_X1 U19845 ( .A1(n17833), .A2(n18043), .B1(n17832), .B2(n17831), .ZN(
        P3_U2688) );
  AOI22_X1 U19846 ( .A1(n18033), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18056), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17844) );
  AOI22_X1 U19847 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17908), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17843) );
  AOI22_X1 U19848 ( .A1(n18046), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17834) );
  OAI21_X1 U19849 ( .B1(n17850), .B2(n17835), .A(n17834), .ZN(n17841) );
  AOI22_X1 U19850 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17839) );
  AOI22_X1 U19851 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17838) );
  AOI22_X1 U19852 ( .A1(n10956), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18013), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17837) );
  AOI22_X1 U19853 ( .A1(n18025), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17865), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17836) );
  NAND4_X1 U19854 ( .A1(n17839), .A2(n17838), .A3(n17837), .A4(n17836), .ZN(
        n17840) );
  AOI211_X1 U19855 ( .C1(n17920), .C2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n17841), .B(n17840), .ZN(n17842) );
  NAND3_X1 U19856 ( .A1(n17844), .A2(n17843), .A3(n17842), .ZN(n20805) );
  INV_X1 U19857 ( .A(n17848), .ZN(n17845) );
  OAI33_X1 U19858 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n20801), .A3(n17845), 
        .B1(n20510), .B2(n18070), .B3(n17848), .ZN(n17846) );
  AOI21_X1 U19859 ( .B1(n18070), .B2(n20805), .A(n17846), .ZN(n17847) );
  INV_X1 U19860 ( .A(n17847), .ZN(P3_U2690) );
  NAND3_X1 U19861 ( .A1(n20971), .A2(P3_EBX_REG_13__SCAN_IN), .A3(n17848), 
        .ZN(n17862) );
  AOI22_X1 U19862 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17859) );
  AOI22_X1 U19863 ( .A1(n17920), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18046), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17858) );
  AOI22_X1 U19864 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17908), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17849) );
  OAI21_X1 U19865 ( .B1(n17850), .B2(n17983), .A(n17849), .ZN(n17856) );
  AOI22_X1 U19866 ( .A1(n18033), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17854) );
  AOI22_X1 U19867 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18056), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17853) );
  AOI22_X1 U19868 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17865), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17852) );
  AOI22_X1 U19869 ( .A1(n18025), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10956), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17851) );
  NAND4_X1 U19870 ( .A1(n17854), .A2(n17853), .A3(n17852), .A4(n17851), .ZN(
        n17855) );
  AOI211_X1 U19871 ( .C1(n10967), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n17856), .B(n17855), .ZN(n17857) );
  NAND3_X1 U19872 ( .A1(n17859), .A2(n17858), .A3(n17857), .ZN(n20958) );
  INV_X1 U19873 ( .A(n20958), .ZN(n17861) );
  NAND3_X1 U19874 ( .A1(n17862), .A2(P3_EBX_REG_14__SCAN_IN), .A3(n18043), 
        .ZN(n17860) );
  OAI221_X1 U19875 ( .B1(n17862), .B2(P3_EBX_REG_14__SCAN_IN), .C1(n18043), 
        .C2(n17861), .A(n17860), .ZN(P3_U2689) );
  NAND3_X1 U19876 ( .A1(n18067), .A2(n17864), .A3(n17863), .ZN(n17877) );
  AOI22_X1 U19877 ( .A1(n10957), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n18056), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17869) );
  AOI22_X1 U19878 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17890), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17868) );
  AOI22_X1 U19879 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17865), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17867) );
  AOI22_X1 U19880 ( .A1(n18025), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10956), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17866) );
  NAND4_X1 U19881 ( .A1(n17869), .A2(n17868), .A3(n17867), .A4(n17866), .ZN(
        n17875) );
  AOI22_X1 U19882 ( .A1(n17920), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18047), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17873) );
  AOI22_X1 U19883 ( .A1(n13919), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17872) );
  AOI22_X1 U19884 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17908), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17871) );
  AOI22_X1 U19885 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17870) );
  NAND4_X1 U19886 ( .A1(n17873), .A2(n17872), .A3(n17871), .A4(n17870), .ZN(
        n17874) );
  NOR2_X1 U19887 ( .A1(n17875), .A2(n17874), .ZN(n20809) );
  NAND3_X1 U19888 ( .A1(n17877), .A2(P3_EBX_REG_12__SCAN_IN), .A3(n18043), 
        .ZN(n17876) );
  OAI221_X1 U19889 ( .B1(n17877), .B2(P3_EBX_REG_12__SCAN_IN), .C1(n18043), 
        .C2(n20809), .A(n17876), .ZN(P3_U2691) );
  INV_X1 U19890 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n20462) );
  NOR3_X1 U19891 ( .A1(n20462), .A2(n20443), .A3(n17916), .ZN(n17902) );
  AOI21_X1 U19892 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17902), .A(
        P3_EBX_REG_11__SCAN_IN), .ZN(n17889) );
  NAND2_X1 U19893 ( .A1(n18043), .A2(n17877), .ZN(n17888) );
  AOI22_X1 U19894 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17881) );
  AOI22_X1 U19895 ( .A1(n18045), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17880) );
  AOI22_X1 U19896 ( .A1(n18025), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10956), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17879) );
  AOI22_X1 U19897 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17998), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17878) );
  NAND4_X1 U19898 ( .A1(n17881), .A2(n17880), .A3(n17879), .A4(n17878), .ZN(
        n17887) );
  AOI22_X1 U19899 ( .A1(n13919), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18056), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17885) );
  AOI22_X1 U19900 ( .A1(n10957), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n18054), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17884) );
  AOI22_X1 U19901 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18047), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17883) );
  AOI22_X1 U19902 ( .A1(n17920), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17890), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17882) );
  NAND4_X1 U19903 ( .A1(n17885), .A2(n17884), .A3(n17883), .A4(n17882), .ZN(
        n17886) );
  NOR2_X1 U19904 ( .A1(n17887), .A2(n17886), .ZN(n20813) );
  OAI22_X1 U19905 ( .A1(n17889), .A2(n17888), .B1(n20813), .B2(n18043), .ZN(
        P3_U2692) );
  AOI22_X1 U19906 ( .A1(n18045), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17894) );
  AOI22_X1 U19907 ( .A1(n17920), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17890), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17893) );
  AOI22_X1 U19908 ( .A1(n10956), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18013), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17892) );
  AOI22_X1 U19909 ( .A1(n18025), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17998), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17891) );
  NAND4_X1 U19910 ( .A1(n17894), .A2(n17893), .A3(n17892), .A4(n17891), .ZN(
        n17900) );
  AOI22_X1 U19911 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17898) );
  AOI22_X1 U19912 ( .A1(n18046), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18056), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17897) );
  AOI22_X1 U19913 ( .A1(n10967), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18047), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17896) );
  AOI22_X1 U19914 ( .A1(n17909), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n18054), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17895) );
  NAND4_X1 U19915 ( .A1(n17898), .A2(n17897), .A3(n17896), .A4(n17895), .ZN(
        n17899) );
  NOR2_X1 U19916 ( .A1(n17900), .A2(n17899), .ZN(n20820) );
  NOR2_X1 U19917 ( .A1(n18070), .A2(n17902), .ZN(n17917) );
  OAI222_X1 U19918 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n20971), .B1(
        P3_EBX_REG_10__SCAN_IN), .B2(n17902), .C1(n17917), .C2(n17901), .ZN(
        n17903) );
  OAI21_X1 U19919 ( .B1(n20820), .B2(n18043), .A(n17903), .ZN(P3_U2693) );
  AOI22_X1 U19920 ( .A1(n10967), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n10971), .ZN(n17907) );
  AOI22_X1 U19921 ( .A1(n13837), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n18056), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17906) );
  AOI22_X1 U19922 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n10956), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n18025), .ZN(n17905) );
  AOI22_X1 U19923 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18013), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17998), .ZN(n17904) );
  NAND4_X1 U19924 ( .A1(n17907), .A2(n17906), .A3(n17905), .A4(n17904), .ZN(
        n17915) );
  AOI22_X1 U19925 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n13919), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17913) );
  AOI22_X1 U19926 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18033), .B1(
        n17908), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17912) );
  AOI22_X1 U19927 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17991), .B1(
        n18047), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17911) );
  AOI22_X1 U19928 ( .A1(n17909), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17920), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17910) );
  NAND4_X1 U19929 ( .A1(n17913), .A2(n17912), .A3(n17911), .A4(n17910), .ZN(
        n17914) );
  NOR2_X1 U19930 ( .A1(n17915), .A2(n17914), .ZN(n20822) );
  NOR2_X1 U19931 ( .A1(n20443), .A2(n17916), .ZN(n17918) );
  OAI21_X1 U19932 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17918), .A(n17917), .ZN(
        n17919) );
  OAI21_X1 U19933 ( .B1(n20822), .B2(n18043), .A(n17919), .ZN(P3_U2694) );
  AOI22_X1 U19934 ( .A1(n18047), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13919), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17924) );
  AOI22_X1 U19935 ( .A1(n17920), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17923) );
  AOI22_X1 U19936 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17998), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17922) );
  AOI22_X1 U19937 ( .A1(n18025), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10956), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17921) );
  NAND4_X1 U19938 ( .A1(n17924), .A2(n17923), .A3(n17922), .A4(n17921), .ZN(
        n17930) );
  AOI22_X1 U19939 ( .A1(n17909), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17928) );
  AOI22_X1 U19940 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17927) );
  AOI22_X1 U19941 ( .A1(n18031), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18045), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17926) );
  AOI22_X1 U19942 ( .A1(n18034), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17890), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17925) );
  NAND4_X1 U19943 ( .A1(n17928), .A2(n17927), .A3(n17926), .A4(n17925), .ZN(
        n17929) );
  NOR2_X1 U19944 ( .A1(n17930), .A2(n17929), .ZN(n17931) );
  XOR2_X1 U19945 ( .A(n17932), .B(n17931), .Z(n20911) );
  NOR2_X1 U19946 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n17933), .ZN(n17935) );
  OAI22_X1 U19947 ( .A1(n20911), .A2(n18043), .B1(n17935), .B2(n17934), .ZN(
        P3_U2673) );
  NOR2_X1 U19948 ( .A1(n18070), .A2(n17936), .ZN(n18009) );
  AOI22_X1 U19949 ( .A1(n18045), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17940) );
  AOI22_X1 U19950 ( .A1(n10957), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17890), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17939) );
  AOI22_X1 U19951 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13835), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17938) );
  AOI22_X1 U19952 ( .A1(n18025), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17998), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17937) );
  NAND4_X1 U19953 ( .A1(n17940), .A2(n17939), .A3(n17938), .A4(n17937), .ZN(
        n17946) );
  AOI22_X1 U19954 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17944) );
  AOI22_X1 U19955 ( .A1(n18034), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17943) );
  AOI22_X1 U19956 ( .A1(n18047), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13919), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17942) );
  AOI22_X1 U19957 ( .A1(n18055), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10967), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17941) );
  NAND4_X1 U19958 ( .A1(n17944), .A2(n17943), .A3(n17942), .A4(n17941), .ZN(
        n17945) );
  NOR2_X1 U19959 ( .A1(n17946), .A2(n17945), .ZN(n20867) );
  INV_X1 U19960 ( .A(n20867), .ZN(n17947) );
  AOI22_X1 U19961 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n18009), .B1(n18070), 
        .B2(n17947), .ZN(n17948) );
  OAI21_X1 U19962 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17949), .A(n17948), .ZN(
        P3_U2682) );
  AOI21_X1 U19963 ( .B1(n17950), .B2(n17961), .A(n17958), .ZN(n20926) );
  NAND2_X1 U19964 ( .A1(n20926), .A2(n18070), .ZN(n17951) );
  OAI221_X1 U19965 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17952), .C1(n20710), 
        .C2(n17953), .A(n17951), .ZN(P3_U2676) );
  INV_X1 U19966 ( .A(n17953), .ZN(n17963) );
  INV_X1 U19967 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n17954) );
  AOI211_X1 U19968 ( .C1(n18067), .C2(n20710), .A(n17963), .B(n17954), .ZN(
        n17960) );
  AOI21_X1 U19969 ( .B1(n17973), .B2(n17955), .A(P3_EBX_REG_28__SCAN_IN), .ZN(
        n17959) );
  OAI21_X1 U19970 ( .B1(n17958), .B2(n17957), .A(n17956), .ZN(n20925) );
  OAI22_X1 U19971 ( .A1(n17960), .A2(n17959), .B1(n20925), .B2(n18043), .ZN(
        P3_U2675) );
  OAI21_X1 U19972 ( .B1(n17965), .B2(n17962), .A(n17961), .ZN(n20905) );
  AOI22_X1 U19973 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17963), .B1(n17969), 
        .B2(n20699), .ZN(n17964) );
  OAI21_X1 U19974 ( .B1(n20905), .B2(n18043), .A(n17964), .ZN(P3_U2677) );
  AOI21_X1 U19975 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n18043), .A(n17973), .ZN(
        n17968) );
  AOI21_X1 U19976 ( .B1(n17966), .B2(n17970), .A(n17965), .ZN(n20895) );
  INV_X1 U19977 ( .A(n20895), .ZN(n17967) );
  OAI22_X1 U19978 ( .A1(n17969), .A2(n17968), .B1(n17967), .B2(n18043), .ZN(
        P3_U2678) );
  AOI21_X1 U19979 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18043), .A(n17980), .ZN(
        n17972) );
  OAI21_X1 U19980 ( .B1(n17975), .B2(n17971), .A(n17970), .ZN(n20941) );
  OAI22_X1 U19981 ( .A1(n17973), .A2(n17972), .B1(n20941), .B2(n18043), .ZN(
        P3_U2679) );
  INV_X1 U19982 ( .A(n17974), .ZN(n17997) );
  AOI21_X1 U19983 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n18043), .A(n17997), .ZN(
        n17979) );
  AOI21_X1 U19984 ( .B1(n17977), .B2(n17976), .A(n17975), .ZN(n20946) );
  INV_X1 U19985 ( .A(n20946), .ZN(n17978) );
  OAI22_X1 U19986 ( .A1(n17980), .A2(n17979), .B1(n17978), .B2(n18043), .ZN(
        P3_U2680) );
  AOI21_X1 U19987 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n18043), .A(n17981), .ZN(
        n17996) );
  AOI22_X1 U19988 ( .A1(n18034), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17994) );
  AOI22_X1 U19989 ( .A1(n18047), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13919), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17993) );
  AOI22_X1 U19990 ( .A1(n18045), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17982) );
  OAI21_X1 U19991 ( .B1(n17984), .B2(n17983), .A(n17982), .ZN(n17990) );
  AOI22_X1 U19992 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18032), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17988) );
  AOI22_X1 U19993 ( .A1(n17909), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17890), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17987) );
  AOI22_X1 U19994 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17998), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17986) );
  AOI22_X1 U19995 ( .A1(n18025), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13835), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17985) );
  NAND4_X1 U19996 ( .A1(n17988), .A2(n17987), .A3(n17986), .A4(n17985), .ZN(
        n17989) );
  AOI211_X1 U19997 ( .C1(n17991), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n17990), .B(n17989), .ZN(n17992) );
  NAND3_X1 U19998 ( .A1(n17994), .A2(n17993), .A3(n17992), .ZN(n20873) );
  INV_X1 U19999 ( .A(n20873), .ZN(n17995) );
  OAI22_X1 U20000 ( .A1(n17997), .A2(n17996), .B1(n17995), .B2(n18043), .ZN(
        P3_U2681) );
  AOI22_X1 U20001 ( .A1(n18055), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18002) );
  AOI22_X1 U20002 ( .A1(n18047), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18046), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n18001) );
  AOI22_X1 U20003 ( .A1(n18025), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17998), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18000) );
  AOI22_X1 U20004 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13835), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17999) );
  NAND4_X1 U20005 ( .A1(n18002), .A2(n18001), .A3(n18000), .A4(n17999), .ZN(
        n18008) );
  AOI22_X1 U20006 ( .A1(n17890), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n18006) );
  AOI22_X1 U20007 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18032), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n18005) );
  AOI22_X1 U20008 ( .A1(n10957), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n18004) );
  AOI22_X1 U20009 ( .A1(n18034), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18045), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n18003) );
  NAND4_X1 U20010 ( .A1(n18006), .A2(n18005), .A3(n18004), .A4(n18003), .ZN(
        n18007) );
  NOR2_X1 U20011 ( .A1(n18008), .A2(n18007), .ZN(n20872) );
  OAI21_X1 U20012 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n18010), .A(n18009), .ZN(
        n18011) );
  OAI21_X1 U20013 ( .B1(n20872), .B2(n18043), .A(n18011), .ZN(P3_U2683) );
  OAI21_X1 U20014 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n18012), .A(n18043), .ZN(
        n18024) );
  AOI22_X1 U20015 ( .A1(n18034), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18017) );
  AOI22_X1 U20016 ( .A1(n18055), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17890), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18016) );
  AOI22_X1 U20017 ( .A1(n18025), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10956), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18015) );
  AOI22_X1 U20018 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17998), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18014) );
  NAND4_X1 U20019 ( .A1(n18017), .A2(n18016), .A3(n18015), .A4(n18014), .ZN(
        n18023) );
  AOI22_X1 U20020 ( .A1(n18047), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18032), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n18021) );
  AOI22_X1 U20021 ( .A1(n17909), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18020) );
  AOI22_X1 U20022 ( .A1(n10967), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18019) );
  AOI22_X1 U20023 ( .A1(n13919), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18045), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n18018) );
  NAND4_X1 U20024 ( .A1(n18021), .A2(n18020), .A3(n18019), .A4(n18018), .ZN(
        n18022) );
  NOR2_X1 U20025 ( .A1(n18023), .A2(n18022), .ZN(n20887) );
  OAI22_X1 U20026 ( .A1(n18042), .A2(n18024), .B1(n20887), .B2(n18043), .ZN(
        P3_U2685) );
  AOI22_X1 U20027 ( .A1(n18045), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18030) );
  AOI22_X1 U20028 ( .A1(n17909), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11010), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n18029) );
  AOI22_X1 U20029 ( .A1(n18025), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17865), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18028) );
  AOI22_X1 U20030 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13835), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18027) );
  NAND4_X1 U20031 ( .A1(n18030), .A2(n18029), .A3(n18028), .A4(n18027), .ZN(
        n18040) );
  AOI22_X1 U20032 ( .A1(n18031), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13919), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18038) );
  AOI22_X1 U20033 ( .A1(n18033), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18032), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n18037) );
  AOI22_X1 U20034 ( .A1(n18055), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n18047), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n18036) );
  AOI22_X1 U20035 ( .A1(n18034), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18035) );
  NAND4_X1 U20036 ( .A1(n18038), .A2(n18037), .A3(n18036), .A4(n18035), .ZN(
        n18039) );
  NOR2_X1 U20037 ( .A1(n18040), .A2(n18039), .ZN(n20883) );
  OAI21_X1 U20038 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n18042), .A(n18041), .ZN(
        n18044) );
  AOI22_X1 U20039 ( .A1(n18070), .A2(n20883), .B1(n18044), .B2(n18043), .ZN(
        P3_U2684) );
  AOI22_X1 U20040 ( .A1(n18045), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n18053) );
  AOI22_X1 U20041 ( .A1(n18047), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n18046), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n18052) );
  AOI22_X1 U20042 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20370), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n17998), .ZN(n18051) );
  AOI22_X1 U20043 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n10956), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n13835), .ZN(n18050) );
  NAND4_X1 U20044 ( .A1(n18053), .A2(n18052), .A3(n18051), .A4(n18050), .ZN(
        n18062) );
  AOI22_X1 U20045 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n10966), .B1(
        n18054), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n18060) );
  AOI22_X1 U20046 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10969), .B1(
        n17890), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18059) );
  AOI22_X1 U20047 ( .A1(n18055), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18058) );
  AOI22_X1 U20048 ( .A1(n10957), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n18056), .ZN(n18057) );
  NAND4_X1 U20049 ( .A1(n18060), .A2(n18059), .A3(n18058), .A4(n18057), .ZN(
        n18061) );
  NOR2_X1 U20050 ( .A1(n18062), .A2(n18061), .ZN(n20894) );
  AOI211_X1 U20051 ( .C1(n20579), .C2(n18064), .A(n18063), .B(n18072), .ZN(
        n18065) );
  AOI21_X1 U20052 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n18069), .A(n18065), .ZN(
        n18066) );
  OAI21_X1 U20053 ( .B1(n20894), .B2(n18043), .A(n18066), .ZN(P3_U2686) );
  NOR2_X1 U20054 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n20359) );
  AOI21_X1 U20055 ( .B1(P3_EBX_REG_1__SCAN_IN), .B2(P3_EBX_REG_0__SCAN_IN), 
        .A(n20359), .ZN(n20346) );
  AOI222_X1 U20056 ( .A1(n20346), .A2(n18067), .B1(P3_EBX_REG_1__SCAN_IN), 
        .B2(n18069), .C1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .C2(n18070), .ZN(
        n18068) );
  INV_X1 U20057 ( .A(n18068), .ZN(P3_U2702) );
  AOI22_X1 U20058 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18070), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n18069), .ZN(n18071) );
  OAI21_X1 U20059 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n18072), .A(n18071), .ZN(
        P3_U2703) );
  INV_X1 U20060 ( .A(n18073), .ZN(n20283) );
  OAI21_X1 U20061 ( .B1(n21469), .B2(n20283), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n18074) );
  OAI21_X1 U20062 ( .B1(n18075), .B2(n20337), .A(n18074), .ZN(P3_U2634) );
  AOI21_X1 U20063 ( .B1(n21506), .B2(n18077), .A(n18076), .ZN(n21494) );
  OAI21_X1 U20064 ( .B1(n21494), .B2(n18475), .A(n18473), .ZN(n18078) );
  OAI221_X1 U20065 ( .B1(n21449), .B2(n18079), .C1(n21449), .C2(n18473), .A(
        n18078), .ZN(P3_U2863) );
  AOI22_X2 U20066 ( .A1(n21362), .A2(n18380), .B1(n18423), .B2(n21041), .ZN(
        n18368) );
  INV_X1 U20067 ( .A(n21366), .ZN(n21374) );
  OAI22_X1 U20068 ( .A1(n21360), .A2(n18468), .B1(n21207), .B2(n18236), .ZN(
        n18122) );
  AOI21_X1 U20069 ( .B1(n18312), .B2(n18086), .A(n18122), .ZN(n18316) );
  INV_X1 U20070 ( .A(n18080), .ZN(n18081) );
  AOI21_X1 U20071 ( .B1(n18329), .B2(n18081), .A(n18439), .ZN(n18306) );
  OAI21_X1 U20072 ( .B1(n20584), .B2(n18464), .A(n18306), .ZN(n18094) );
  NOR3_X1 U20073 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18240), .A3(
        n18081), .ZN(n18095) );
  INV_X1 U20074 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n21378) );
  INV_X1 U20075 ( .A(n18093), .ZN(n18082) );
  OAI21_X1 U20076 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n20584), .A(
        n18082), .ZN(n20587) );
  OAI22_X1 U20077 ( .A1(n21428), .A2(n21378), .B1(n18304), .B2(n20587), .ZN(
        n18083) );
  AOI211_X1 U20078 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n18094), .A(
        n18095), .B(n18083), .ZN(n18088) );
  OAI21_X1 U20079 ( .B1(n21308), .B2(n18091), .A(n18176), .ZN(n18085) );
  XOR2_X1 U20080 ( .A(n18084), .B(n18085), .Z(n21376) );
  NOR2_X1 U20081 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18086), .ZN(
        n21375) );
  AOI22_X1 U20082 ( .A1(n18379), .A2(n21376), .B1(n18312), .B2(n21375), .ZN(
        n18087) );
  OAI211_X1 U20083 ( .C1(n18316), .C2(n18091), .A(n18088), .B(n18087), .ZN(
        P3_U2812) );
  NAND2_X1 U20084 ( .A1(n18089), .A2(n18312), .ZN(n18180) );
  NAND3_X1 U20085 ( .A1(n18089), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n21207), .ZN(n21344) );
  NAND3_X1 U20086 ( .A1(n18089), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n21360), .ZN(n21342) );
  AOI22_X1 U20087 ( .A1(n18380), .A2(n21344), .B1(n18423), .B2(n21342), .ZN(
        n18182) );
  OAI21_X1 U20088 ( .B1(n18176), .B2(n18084), .A(n18178), .ZN(n18092) );
  XNOR2_X1 U20089 ( .A(n18092), .B(n18177), .ZN(n21348) );
  NOR3_X1 U20090 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18240), .A3(
        n20594), .ZN(n18098) );
  OAI21_X1 U20091 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18093), .A(
        n18186), .ZN(n20596) );
  OAI21_X1 U20092 ( .B1(n18095), .B2(n18094), .A(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18096) );
  NAND2_X1 U20093 ( .A1(n21401), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n21349) );
  OAI211_X1 U20094 ( .C1(n18304), .C2(n20596), .A(n18096), .B(n21349), .ZN(
        n18097) );
  AOI211_X1 U20095 ( .C1(n18379), .C2(n21348), .A(n18098), .B(n18097), .ZN(
        n18099) );
  OAI221_X1 U20096 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18180), 
        .C1(n18177), .C2(n18182), .A(n18099), .ZN(P3_U2811) );
  OR2_X1 U20097 ( .A1(n18236), .A2(n21207), .ZN(n18112) );
  OAI21_X1 U20098 ( .B1(n18427), .B2(n18102), .A(n11018), .ZN(n18101) );
  INV_X1 U20099 ( .A(n18101), .ZN(n18318) );
  OAI21_X1 U20100 ( .B1(n18100), .B2(n18464), .A(n18318), .ZN(n18119) );
  INV_X1 U20101 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n20550) );
  NOR2_X1 U20102 ( .A1(n21379), .A2(n20550), .ZN(n21202) );
  NAND2_X1 U20103 ( .A1(n18102), .A2(n18238), .ZN(n18114) );
  INV_X1 U20104 ( .A(n18100), .ZN(n18115) );
  AOI22_X1 U20105 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18115), .B1(
        n18100), .B2(n20545), .ZN(n20536) );
  OAI22_X1 U20106 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18114), .B1(
        n20536), .B2(n18304), .ZN(n18103) );
  AOI211_X1 U20107 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n18119), .A(
        n21202), .B(n18103), .ZN(n18111) );
  NAND2_X1 U20108 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18104) );
  NOR3_X1 U20109 ( .A1(n13867), .A2(n21308), .A3(n18104), .ZN(n18340) );
  NAND2_X1 U20110 ( .A1(n21180), .A2(n18340), .ZN(n18322) );
  INV_X1 U20111 ( .A(n18105), .ZN(n18106) );
  NAND2_X1 U20112 ( .A1(n18106), .A2(n21423), .ZN(n18356) );
  NOR2_X1 U20113 ( .A1(n18351), .A2(n18356), .ZN(n18332) );
  NAND2_X1 U20114 ( .A1(n18107), .A2(n18332), .ZN(n18323) );
  AOI22_X1 U20115 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18322), .B1(
        n18323), .B2(n13871), .ZN(n18108) );
  XNOR2_X1 U20116 ( .A(n21213), .B(n18108), .ZN(n21203) );
  OAI21_X1 U20117 ( .B1(n21200), .B2(n18468), .A(n21213), .ZN(n18109) );
  AOI22_X1 U20118 ( .A1(n18379), .A2(n21203), .B1(n18122), .B2(n18109), .ZN(
        n18110) );
  OAI211_X1 U20119 ( .C1(n18113), .C2(n18112), .A(n18111), .B(n18110), .ZN(
        P3_U2815) );
  INV_X1 U20120 ( .A(n18312), .ZN(n18125) );
  AOI211_X1 U20121 ( .C1(n20545), .C2(n20554), .A(n20562), .B(n18114), .ZN(
        n18118) );
  INV_X1 U20122 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n20551) );
  NOR2_X1 U20123 ( .A1(n20545), .A2(n18115), .ZN(n18116) );
  OAI21_X1 U20124 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18116), .A(
        n18303), .ZN(n20547) );
  OAI22_X1 U20125 ( .A1(n21428), .A2(n20551), .B1(n18304), .B2(n20547), .ZN(
        n18117) );
  AOI211_X1 U20126 ( .C1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n18119), .A(
        n18118), .B(n18117), .ZN(n18124) );
  AOI22_X1 U20127 ( .A1(n18258), .A2(n21398), .B1(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n21308), .ZN(n18120) );
  XNOR2_X1 U20128 ( .A(n18121), .B(n18120), .ZN(n21395) );
  AOI22_X1 U20129 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18122), .B1(
        n18379), .B2(n21395), .ZN(n18123) );
  OAI211_X1 U20130 ( .C1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n18125), .A(
        n18124), .B(n18123), .ZN(P3_U2814) );
  INV_X1 U20131 ( .A(n21158), .ZN(n18352) );
  INV_X1 U20132 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18337) );
  NOR2_X1 U20133 ( .A1(n18352), .A2(n18337), .ZN(n21175) );
  INV_X1 U20134 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18144) );
  NAND2_X1 U20135 ( .A1(n21175), .A2(n18144), .ZN(n18135) );
  NOR2_X1 U20136 ( .A1(n18240), .A2(n18126), .ZN(n18138) );
  INV_X1 U20137 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18129) );
  NOR2_X1 U20138 ( .A1(n18126), .A2(n11129), .ZN(n18328) );
  AOI21_X1 U20139 ( .B1(n18329), .B2(n18126), .A(n18439), .ZN(n18127) );
  OAI21_X1 U20140 ( .B1(n18328), .B2(n18464), .A(n18127), .ZN(n18142) );
  NAND2_X1 U20141 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18328), .ZN(
        n20507) );
  OAI21_X1 U20142 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18328), .A(
        n20507), .ZN(n20494) );
  NAND2_X1 U20143 ( .A1(n21401), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n21177) );
  OAI21_X1 U20144 ( .B1(n18304), .B2(n20494), .A(n21177), .ZN(n18128) );
  AOI221_X1 U20145 ( .B1(n18138), .B2(n18129), .C1(n18142), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n18128), .ZN(n18134) );
  NAND2_X1 U20146 ( .A1(n18130), .A2(n21041), .ZN(n21168) );
  INV_X1 U20147 ( .A(n21168), .ZN(n18131) );
  OAI22_X1 U20148 ( .A1(n21170), .A2(n18236), .B1(n18131), .B2(n18468), .ZN(
        n18146) );
  INV_X1 U20149 ( .A(n18340), .ZN(n18355) );
  NOR2_X1 U20150 ( .A1(n18352), .A2(n18355), .ZN(n18132) );
  AOI22_X1 U20151 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18132), .B1(
        n18332), .B2(n18337), .ZN(n18143) );
  XNOR2_X1 U20152 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n18143), .ZN(
        n21176) );
  AOI22_X1 U20153 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18146), .B1(
        n18379), .B2(n21176), .ZN(n18133) );
  OAI211_X1 U20154 ( .C1(n18368), .C2(n18135), .A(n18134), .B(n18133), .ZN(
        P3_U2818) );
  OR2_X1 U20155 ( .A1(n21166), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n21408) );
  INV_X1 U20156 ( .A(n20507), .ZN(n18136) );
  OAI21_X1 U20157 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n18136), .A(
        n20502), .ZN(n20505) );
  OAI211_X1 U20158 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n18138), .B(n18137), .ZN(n18140) );
  NAND2_X1 U20159 ( .A1(n21401), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n18139) );
  OAI211_X1 U20160 ( .C1(n18304), .C2(n20505), .A(n18140), .B(n18139), .ZN(
        n18141) );
  AOI21_X1 U20161 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n18142), .A(
        n18141), .ZN(n18148) );
  AOI221_X1 U20162 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18337), 
        .C1(n18144), .C2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n18143), .ZN(
        n18145) );
  XOR2_X1 U20163 ( .A(n18145), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Z(
        n21400) );
  AOI22_X1 U20164 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18146), .B1(
        n18379), .B2(n21400), .ZN(n18147) );
  OAI211_X1 U20165 ( .C1(n18368), .C2(n21408), .A(n18148), .B(n18147), .ZN(
        P3_U2817) );
  NOR2_X2 U20166 ( .A1(n18149), .A2(n18180), .ZN(n18274) );
  INV_X1 U20167 ( .A(n18274), .ZN(n18162) );
  NAND2_X1 U20168 ( .A1(n18150), .A2(n21207), .ZN(n21047) );
  NAND2_X1 U20169 ( .A1(n18150), .A2(n21360), .ZN(n21046) );
  AOI22_X1 U20170 ( .A1(n18380), .A2(n21047), .B1(n18423), .B2(n21046), .ZN(
        n18170) );
  INV_X1 U20171 ( .A(n18151), .ZN(n18153) );
  OAI21_X1 U20172 ( .B1(n18154), .B2(n18153), .A(n18152), .ZN(n18192) );
  XNOR2_X1 U20173 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n18192), .ZN(
        n21225) );
  INV_X1 U20174 ( .A(n18305), .ZN(n18265) );
  AOI22_X1 U20175 ( .A1(n18196), .A2(n18186), .B1(n18329), .B2(n18166), .ZN(
        n18155) );
  NAND2_X1 U20176 ( .A1(n18155), .A2(n11018), .ZN(n18184) );
  AOI21_X1 U20177 ( .B1(n18265), .B2(n18187), .A(n18184), .ZN(n18167) );
  INV_X1 U20178 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n20642) );
  NAND2_X1 U20179 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n18185), .ZN(
        n18156) );
  AOI21_X1 U20180 ( .B1(n20642), .B2(n18156), .A(n18197), .ZN(n20639) );
  INV_X1 U20181 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18168) );
  AOI211_X1 U20182 ( .C1(n20642), .C2(n18168), .A(n18240), .B(n18166), .ZN(
        n18158) );
  AOI22_X1 U20183 ( .A1(n20639), .A2(n18297), .B1(n18158), .B2(n18157), .ZN(
        n18159) );
  NAND2_X1 U20184 ( .A1(n21401), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n21226) );
  OAI211_X1 U20185 ( .C1(n18167), .C2(n20642), .A(n18159), .B(n21226), .ZN(
        n18160) );
  AOI21_X1 U20186 ( .B1(n18379), .B2(n21225), .A(n18160), .ZN(n18161) );
  OAI221_X1 U20187 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18162), 
        .C1(n21257), .C2(n18170), .A(n18161), .ZN(P3_U2808) );
  INV_X1 U20188 ( .A(n21049), .ZN(n21051) );
  OAI22_X1 U20189 ( .A1(n21051), .A2(n18178), .B1(n18163), .B2(n18084), .ZN(
        n18164) );
  XOR2_X1 U20190 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18164), .Z(
        n21054) );
  INV_X1 U20191 ( .A(n21054), .ZN(n18174) );
  AOI22_X1 U20192 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n18185), .B1(
        n18165), .B2(n18168), .ZN(n20629) );
  OR2_X1 U20193 ( .A1(n18166), .A2(n18240), .ZN(n18169) );
  NAND2_X1 U20194 ( .A1(n21401), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n21055) );
  OAI221_X1 U20195 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n18169), .C1(
        n18168), .C2(n18167), .A(n21055), .ZN(n18172) );
  INV_X1 U20196 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n21220) );
  NAND2_X1 U20197 ( .A1(n21049), .A2(n21220), .ZN(n21057) );
  OAI22_X1 U20198 ( .A1(n18170), .A2(n21220), .B1(n18180), .B2(n21057), .ZN(
        n18171) );
  AOI211_X1 U20199 ( .C1(n18297), .C2(n20629), .A(n18172), .B(n18171), .ZN(
        n18173) );
  OAI21_X1 U20200 ( .B1(n18174), .B2(n18287), .A(n18173), .ZN(P3_U2809) );
  INV_X1 U20201 ( .A(n18152), .ZN(n18175) );
  AOI221_X1 U20202 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18178), 
        .C1(n18177), .C2(n18176), .A(n18175), .ZN(n18179) );
  XNOR2_X1 U20203 ( .A(n18179), .B(n18181), .ZN(n21351) );
  NAND2_X1 U20204 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18181), .ZN(
        n21359) );
  OAI22_X1 U20205 ( .A1(n18182), .A2(n18181), .B1(n18180), .B2(n21359), .ZN(
        n18183) );
  AOI21_X1 U20206 ( .B1(n18379), .B2(n21351), .A(n18183), .ZN(n18191) );
  NAND2_X1 U20207 ( .A1(n21401), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n18190) );
  OAI221_X1 U20208 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20617), .C1(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n19215), .A(n18184), .ZN(
        n18189) );
  AOI21_X1 U20209 ( .B1(n18187), .B2(n18186), .A(n18185), .ZN(n20619) );
  OAI21_X1 U20210 ( .B1(n18297), .B2(n18265), .A(n20619), .ZN(n18188) );
  NAND4_X1 U20211 ( .A1(n18191), .A2(n18190), .A3(n18189), .A4(n18188), .ZN(
        P3_U2810) );
  AOI221_X1 U20212 ( .B1(n21308), .B2(n18193), .C1(n21257), .C2(n18193), .A(
        n18192), .ZN(n18194) );
  XNOR2_X1 U20213 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n18194), .ZN(
        n21328) );
  AND2_X1 U20214 ( .A1(n18214), .A2(n19215), .ZN(n18202) );
  INV_X1 U20215 ( .A(n18197), .ZN(n18195) );
  AOI211_X1 U20216 ( .C1(n18196), .C2(n18195), .A(n18439), .B(n18202), .ZN(
        n18212) );
  INV_X1 U20217 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18200) );
  NAND2_X1 U20218 ( .A1(n21401), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n21327) );
  OAI21_X1 U20219 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18197), .A(
        n18227), .ZN(n18198) );
  INV_X1 U20220 ( .A(n18198), .ZN(n20656) );
  OAI21_X1 U20221 ( .B1(n18297), .B2(n18265), .A(n20656), .ZN(n18199) );
  OAI211_X1 U20222 ( .C1(n18212), .C2(n18200), .A(n21327), .B(n18199), .ZN(
        n18201) );
  AOI21_X1 U20223 ( .B1(n18203), .B2(n18202), .A(n18201), .ZN(n18209) );
  NAND2_X1 U20224 ( .A1(n18423), .A2(n21319), .ZN(n18205) );
  NAND2_X1 U20225 ( .A1(n18380), .A2(n21320), .ZN(n18204) );
  OAI22_X1 U20226 ( .A1(n21046), .A2(n18205), .B1(n21047), .B2(n18204), .ZN(
        n18207) );
  OAI21_X1 U20227 ( .B1(n18206), .B2(n18236), .A(n18205), .ZN(n18233) );
  AOI22_X1 U20228 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18207), .B1(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18233), .ZN(n18208) );
  OAI211_X1 U20229 ( .C1(n18287), .C2(n21328), .A(n18209), .B(n18208), .ZN(
        P3_U2807) );
  OAI21_X1 U20230 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n18211), .A(
        n18210), .ZN(n21238) );
  OAI21_X1 U20231 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18305), .A(
        n18212), .ZN(n18230) );
  INV_X1 U20232 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n20671) );
  NOR2_X1 U20233 ( .A1(n20671), .A2(n18227), .ZN(n18226) );
  INV_X1 U20234 ( .A(n18267), .ZN(n18213) );
  OAI21_X1 U20235 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n18226), .A(
        n18213), .ZN(n20679) );
  NOR2_X1 U20236 ( .A1(n18240), .A2(n18214), .ZN(n18231) );
  OAI211_X1 U20237 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n18231), .B(n18215), .ZN(n18216) );
  NAND2_X1 U20238 ( .A1(n21401), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n21243) );
  OAI211_X1 U20239 ( .C1(n18304), .C2(n20679), .A(n18216), .B(n21243), .ZN(
        n18217) );
  AOI21_X1 U20240 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n18230), .A(
        n18217), .ZN(n18223) );
  AOI21_X1 U20241 ( .B1(n21247), .B2(n18219), .A(n18218), .ZN(n21237) );
  OAI21_X1 U20242 ( .B1(n21308), .B2(n11032), .A(n18220), .ZN(n18221) );
  XNOR2_X1 U20243 ( .A(n18221), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n21242) );
  AOI22_X1 U20244 ( .A1(n18380), .A2(n21237), .B1(n18379), .B2(n21242), .ZN(
        n18222) );
  OAI211_X1 U20245 ( .C1(n18468), .C2(n21238), .A(n18223), .B(n18222), .ZN(
        P3_U2805) );
  AOI21_X1 U20246 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n18225), .A(
        n18224), .ZN(n21338) );
  INV_X1 U20247 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n20678) );
  AOI21_X1 U20248 ( .B1(n20671), .B2(n18227), .A(n18226), .ZN(n20668) );
  INV_X1 U20249 ( .A(n20668), .ZN(n18228) );
  OAI22_X1 U20250 ( .A1(n21428), .A2(n20678), .B1(n18304), .B2(n18228), .ZN(
        n18229) );
  AOI221_X1 U20251 ( .B1(n18231), .B2(n20671), .C1(n18230), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n18229), .ZN(n18235) );
  NOR2_X1 U20252 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n21329), .ZN(
        n18232) );
  AOI22_X1 U20253 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18233), .B1(
        n18274), .B2(n18232), .ZN(n18234) );
  OAI211_X1 U20254 ( .C1(n21338), .C2(n18287), .A(n18235), .B(n18234), .ZN(
        P3_U2806) );
  INV_X1 U20255 ( .A(n21269), .ZN(n21245) );
  OAI22_X1 U20256 ( .A1(n21275), .A2(n18468), .B1(n21245), .B2(n18236), .ZN(
        n18273) );
  NOR2_X1 U20257 ( .A1(n21306), .A2(n18273), .ZN(n18263) );
  OAI21_X1 U20258 ( .B1(n18380), .B2(n18423), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n18252) );
  NAND2_X1 U20259 ( .A1(n18237), .A2(n18274), .ZN(n18280) );
  NOR3_X1 U20260 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n21306), .A3(
        n18280), .ZN(n18246) );
  OAI21_X1 U20261 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n18253), .A(
        n18296), .ZN(n20723) );
  INV_X1 U20262 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n20732) );
  NAND3_X1 U20263 ( .A1(n18239), .A2(n20732), .A3(n18238), .ZN(n18244) );
  NOR3_X1 U20264 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n18240), .A3(
        n18242), .ZN(n18255) );
  OAI21_X1 U20265 ( .B1(n18267), .B2(n18464), .A(n11018), .ZN(n18241) );
  AOI21_X1 U20266 ( .B1(n18329), .B2(n18242), .A(n18241), .ZN(n18270) );
  OAI21_X1 U20267 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18305), .A(
        n18270), .ZN(n18259) );
  OAI21_X1 U20268 ( .B1(n18255), .B2(n18259), .A(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n18243) );
  OAI211_X1 U20269 ( .C1(n18304), .C2(n20723), .A(n18244), .B(n18243), .ZN(
        n18245) );
  AOI211_X1 U20270 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n21401), .A(n18246), 
        .B(n18245), .ZN(n18251) );
  AOI21_X1 U20271 ( .B1(n18258), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n18247), .ZN(n21314) );
  NAND2_X1 U20272 ( .A1(n18257), .A2(n18258), .ZN(n18256) );
  NAND2_X1 U20273 ( .A1(n18256), .A2(n21315), .ZN(n18249) );
  NAND2_X1 U20274 ( .A1(n18249), .A2(n21314), .ZN(n21296) );
  OAI211_X1 U20275 ( .C1(n21314), .C2(n18249), .A(n18379), .B(n21296), .ZN(
        n18250) );
  OAI211_X1 U20276 ( .C1(n18263), .C2(n18252), .A(n18251), .B(n18250), .ZN(
        P3_U2802) );
  AND2_X1 U20277 ( .A1(n21306), .A2(n18280), .ZN(n18262) );
  AOI21_X1 U20278 ( .B1(n18254), .B2(n18266), .A(n18253), .ZN(n20714) );
  INV_X1 U20279 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n20721) );
  NOR2_X1 U20280 ( .A1(n21379), .A2(n20721), .ZN(n21265) );
  AOI211_X1 U20281 ( .C1(n18297), .C2(n20714), .A(n21265), .B(n18255), .ZN(
        n18261) );
  OAI21_X1 U20282 ( .B1(n18258), .B2(n18257), .A(n18256), .ZN(n21266) );
  AOI22_X1 U20283 ( .A1(n18379), .A2(n21266), .B1(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n18259), .ZN(n18260) );
  OAI211_X1 U20284 ( .C1(n18263), .C2(n18262), .A(n18261), .B(n18260), .ZN(
        P3_U2803) );
  OAI221_X1 U20285 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n21308), 
        .C1(n21247), .C2(n11032), .A(n18220), .ZN(n18264) );
  XNOR2_X1 U20286 ( .A(n21246), .B(n18264), .ZN(n21256) );
  OAI21_X1 U20287 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18267), .A(
        n18266), .ZN(n20694) );
  AOI21_X1 U20288 ( .B1(n18304), .B2(n18305), .A(n20694), .ZN(n18272) );
  AOI21_X1 U20289 ( .B1(n18268), .B2(n19215), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n18269) );
  INV_X1 U20290 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n20707) );
  OAI22_X1 U20291 ( .A1(n18270), .A2(n18269), .B1(n21379), .B2(n20707), .ZN(
        n18271) );
  AOI211_X1 U20292 ( .C1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n18273), .A(
        n18272), .B(n18271), .ZN(n18276) );
  NOR2_X1 U20293 ( .A1(n21247), .A2(n21235), .ZN(n21252) );
  NAND3_X1 U20294 ( .A1(n18274), .A2(n21252), .A3(n21246), .ZN(n18275) );
  OAI211_X1 U20295 ( .C1(n21256), .C2(n18287), .A(n18276), .B(n18275), .ZN(
        P3_U2804) );
  AOI22_X1 U20296 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n21299), .B1(
        n18291), .B2(n21288), .ZN(n18277) );
  XNOR2_X1 U20297 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n18277), .ZN(
        n21295) );
  XOR2_X1 U20298 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n18295), .Z(
        n20763) );
  INV_X1 U20299 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n20753) );
  NAND2_X1 U20300 ( .A1(n21401), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n21293) );
  OAI221_X1 U20301 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n18279), .C1(
        n20753), .C2(n18278), .A(n21293), .ZN(n18285) );
  NOR2_X1 U20302 ( .A1(n18281), .A2(n18280), .ZN(n18283) );
  NAND2_X1 U20303 ( .A1(n21245), .A2(n21274), .ZN(n21277) );
  AOI21_X1 U20304 ( .B1(n18380), .B2(n21277), .A(n18293), .ZN(n18282) );
  INV_X1 U20305 ( .A(n18282), .ZN(n18294) );
  MUX2_X1 U20306 ( .A(n18283), .B(n18294), .S(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Z(n18284) );
  OAI21_X1 U20307 ( .B1(n21295), .B2(n18287), .A(n18286), .ZN(P3_U2800) );
  OAI21_X1 U20308 ( .B1(n18288), .B2(n19054), .A(n20736), .ZN(n18289) );
  AOI22_X1 U20309 ( .A1(n21401), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n18290), 
        .B2(n18289), .ZN(n18302) );
  INV_X1 U20310 ( .A(n21268), .ZN(n21279) );
  NAND2_X1 U20311 ( .A1(n18291), .A2(n21299), .ZN(n18292) );
  XNOR2_X1 U20312 ( .A(n18292), .B(n21288), .ZN(n21282) );
  AOI22_X1 U20313 ( .A1(n11245), .A2(n18293), .B1(n18379), .B2(n21282), .ZN(
        n18301) );
  NOR2_X1 U20314 ( .A1(n21269), .A2(n21268), .ZN(n21301) );
  OAI21_X1 U20315 ( .B1(n21301), .B2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n18294), .ZN(n18300) );
  AOI21_X1 U20316 ( .B1(n20736), .B2(n18296), .A(n18295), .ZN(n20735) );
  OAI21_X1 U20317 ( .B1(n18298), .B2(n18297), .A(n20735), .ZN(n18299) );
  NAND4_X1 U20318 ( .A1(n18302), .A2(n18301), .A3(n18300), .A4(n18299), .ZN(
        P3_U2801) );
  AOI21_X1 U20319 ( .B1(n18307), .B2(n18303), .A(n20584), .ZN(n20565) );
  INV_X1 U20320 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n20573) );
  NOR2_X1 U20321 ( .A1(n21379), .A2(n20573), .ZN(n21387) );
  AOI221_X1 U20322 ( .B1(n18308), .B2(n18307), .C1(n19054), .C2(n18307), .A(
        n18306), .ZN(n18309) );
  AOI211_X1 U20323 ( .C1(n20565), .C2(n18450), .A(n21387), .B(n18309), .ZN(
        n18314) );
  OAI21_X1 U20324 ( .B1(n18311), .B2(n18315), .A(n18310), .ZN(n21385) );
  NOR2_X1 U20325 ( .A1(n21398), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n21381) );
  AOI22_X1 U20326 ( .A1(n18379), .A2(n21385), .B1(n18312), .B2(n21381), .ZN(
        n18313) );
  OAI211_X1 U20327 ( .C1(n18316), .C2(n18315), .A(n18314), .B(n18313), .ZN(
        P3_U2813) );
  OAI21_X1 U20328 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18317), .A(
        n21200), .ZN(n21185) );
  AOI21_X1 U20329 ( .B1(n20519), .B2(n20502), .A(n18100), .ZN(n20529) );
  AOI221_X1 U20330 ( .B1(n11050), .B2(n20519), .C1(n19054), .C2(n20519), .A(
        n18318), .ZN(n18320) );
  NAND2_X1 U20331 ( .A1(n21401), .A2(P3_REIP_REG_14__SCAN_IN), .ZN(n21191) );
  INV_X1 U20332 ( .A(n21191), .ZN(n18319) );
  AOI211_X1 U20333 ( .C1(n20529), .C2(n18450), .A(n18320), .B(n18319), .ZN(
        n18326) );
  AOI21_X1 U20334 ( .B1(n13871), .B2(n18321), .A(n21208), .ZN(n21189) );
  NAND2_X1 U20335 ( .A1(n18323), .A2(n18322), .ZN(n18324) );
  XNOR2_X1 U20336 ( .A(n18324), .B(n13871), .ZN(n21190) );
  AOI22_X1 U20337 ( .A1(n18380), .A2(n21189), .B1(n18379), .B2(n21190), .ZN(
        n18325) );
  OAI211_X1 U20338 ( .C1(n18468), .C2(n21185), .A(n18326), .B(n18325), .ZN(
        P3_U2816) );
  AOI22_X1 U20339 ( .A1(n18423), .A2(n21155), .B1(n18380), .B2(n18327), .ZN(
        n18367) );
  INV_X1 U20340 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n20490) );
  INV_X1 U20341 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20456) );
  NAND2_X1 U20342 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n20414), .ZN(
        n18374) );
  NOR2_X1 U20343 ( .A1(n11129), .A2(n18374), .ZN(n18391) );
  NAND2_X1 U20344 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18391), .ZN(
        n20450) );
  NOR2_X1 U20345 ( .A1(n20456), .A2(n20450), .ZN(n18360) );
  NAND2_X1 U20346 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18360), .ZN(
        n18345) );
  AOI21_X1 U20347 ( .B1(n20490), .B2(n18345), .A(n18328), .ZN(n20482) );
  NOR3_X1 U20348 ( .A1(n18399), .A2(n18397), .A3(n19054), .ZN(n18387) );
  NAND2_X1 U20349 ( .A1(n20480), .A2(n18387), .ZN(n18344) );
  NAND2_X1 U20350 ( .A1(n18344), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18330) );
  NAND2_X1 U20351 ( .A1(n21401), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n21162) );
  OAI221_X1 U20352 ( .B1(n18344), .B2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C1(
        n18330), .C2(n18459), .A(n21162), .ZN(n18331) );
  AOI21_X1 U20353 ( .B1(n20482), .B2(n18450), .A(n18331), .ZN(n18336) );
  AOI21_X1 U20354 ( .B1(n18340), .B2(n21158), .A(n18332), .ZN(n18333) );
  XNOR2_X1 U20355 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18333), .ZN(
        n21160) );
  INV_X1 U20356 ( .A(n18368), .ZN(n18350) );
  NAND2_X1 U20357 ( .A1(n21158), .A2(n18337), .ZN(n21164) );
  OAI21_X1 U20358 ( .B1(n21158), .B2(n18337), .A(n21164), .ZN(n18334) );
  AOI22_X1 U20359 ( .A1(n18379), .A2(n21160), .B1(n18350), .B2(n18334), .ZN(
        n18335) );
  OAI211_X1 U20360 ( .C1(n18367), .C2(n18337), .A(n18336), .B(n18335), .ZN(
        P3_U2819) );
  INV_X1 U20361 ( .A(n18351), .ZN(n18343) );
  AOI21_X1 U20362 ( .B1(n21308), .B2(n21435), .A(n18340), .ZN(n18338) );
  AOI211_X1 U20363 ( .C1(n18339), .C2(n21435), .A(n18338), .B(n21412), .ZN(
        n18342) );
  NOR3_X1 U20364 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18340), .A3(
        n21435), .ZN(n18341) );
  AOI211_X1 U20365 ( .C1(n18343), .C2(n18356), .A(n18342), .B(n18341), .ZN(
        n21416) );
  NAND2_X1 U20366 ( .A1(n21401), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n21417) );
  INV_X1 U20367 ( .A(n21417), .ZN(n18349) );
  INV_X1 U20368 ( .A(n18344), .ZN(n18347) );
  INV_X1 U20369 ( .A(n18459), .ZN(n18359) );
  AOI22_X1 U20370 ( .A1(n18358), .A2(n18387), .B1(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18359), .ZN(n18346) );
  OAI21_X1 U20371 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18360), .A(
        n18345), .ZN(n20468) );
  OAI22_X1 U20372 ( .A1(n18347), .A2(n18346), .B1(n18460), .B2(n20468), .ZN(
        n18348) );
  AOI211_X1 U20373 ( .C1(n18379), .C2(n21416), .A(n18349), .B(n18348), .ZN(
        n18354) );
  NAND3_X1 U20374 ( .A1(n18352), .A2(n18351), .A3(n18350), .ZN(n18353) );
  OAI211_X1 U20375 ( .C1(n18367), .C2(n21412), .A(n18354), .B(n18353), .ZN(
        P3_U2820) );
  NAND2_X1 U20376 ( .A1(n18356), .A2(n18355), .ZN(n18357) );
  XNOR2_X1 U20377 ( .A(n18357), .B(n21435), .ZN(n21431) );
  INV_X1 U20378 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18546) );
  NOR2_X1 U20379 ( .A1(n21379), .A2(n18546), .ZN(n18365) );
  AND2_X1 U20380 ( .A1(n18358), .A2(n18387), .ZN(n18363) );
  AOI22_X1 U20381 ( .A1(n18373), .A2(n18387), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18359), .ZN(n18362) );
  AOI21_X1 U20382 ( .B1(n20456), .B2(n20450), .A(n18360), .ZN(n18361) );
  INV_X1 U20383 ( .A(n18361), .ZN(n20453) );
  OAI22_X1 U20384 ( .A1(n18363), .A2(n18362), .B1(n18460), .B2(n20453), .ZN(
        n18364) );
  AOI211_X1 U20385 ( .C1(n18379), .C2(n21431), .A(n18365), .B(n18364), .ZN(
        n18366) );
  OAI221_X1 U20386 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18368), .C1(
        n21435), .C2(n18367), .A(n18366), .ZN(P3_U2821) );
  OAI21_X1 U20387 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18370), .A(
        n18369), .ZN(n21145) );
  AOI21_X1 U20388 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n21308), .A(
        n18371), .ZN(n18372) );
  XNOR2_X1 U20389 ( .A(n18372), .B(n14008), .ZN(n21148) );
  INV_X1 U20390 ( .A(n21148), .ZN(n21147) );
  OAI21_X1 U20391 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18391), .A(
        n20450), .ZN(n20438) );
  AOI21_X1 U20392 ( .B1(n20414), .B2(n11018), .A(n18459), .ZN(n18388) );
  AOI211_X1 U20393 ( .C1(n18375), .C2(n18374), .A(n18373), .B(n19054), .ZN(
        n18376) );
  AOI21_X1 U20394 ( .B1(n18388), .B2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n18376), .ZN(n18377) );
  NAND2_X1 U20395 ( .A1(n21401), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n21149) );
  OAI211_X1 U20396 ( .C1(n18460), .C2(n20438), .A(n18377), .B(n21149), .ZN(
        n18378) );
  AOI221_X1 U20397 ( .B1(n18380), .B2(n21147), .C1(n18379), .C2(n21148), .A(
        n18378), .ZN(n18381) );
  OAI21_X1 U20398 ( .B1(n18468), .B2(n21145), .A(n18381), .ZN(P3_U2822) );
  INV_X1 U20399 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n21128) );
  OAI21_X1 U20400 ( .B1(n18384), .B2(n18383), .A(n18382), .ZN(n18385) );
  XNOR2_X1 U20401 ( .A(n18385), .B(n21135), .ZN(n21141) );
  OAI22_X1 U20402 ( .A1(n21379), .A2(n21128), .B1(n18468), .B2(n21141), .ZN(
        n18386) );
  AOI221_X1 U20403 ( .B1(n18388), .B2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C1(
        n18387), .C2(n20436), .A(n18386), .ZN(n18393) );
  AOI21_X1 U20404 ( .B1(n21135), .B2(n18390), .A(n18389), .ZN(n21130) );
  NAND2_X1 U20405 ( .A1(n20414), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18400) );
  AOI21_X1 U20406 ( .B1(n20436), .B2(n18400), .A(n18391), .ZN(n20423) );
  AOI22_X1 U20407 ( .A1(n18457), .A2(n21130), .B1(n20423), .B2(n18450), .ZN(
        n18392) );
  NAND2_X1 U20408 ( .A1(n18393), .A2(n18392), .ZN(P3_U2823) );
  INV_X1 U20409 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n20430) );
  AOI21_X1 U20410 ( .B1(n18396), .B2(n18395), .A(n18394), .ZN(n21124) );
  NOR2_X1 U20411 ( .A1(n18399), .A2(n19054), .ZN(n18398) );
  AOI22_X1 U20412 ( .A1(n18457), .A2(n21124), .B1(n18398), .B2(n18397), .ZN(
        n18405) );
  NOR2_X1 U20413 ( .A1(n18459), .A2(n18398), .ZN(n18415) );
  NOR2_X1 U20414 ( .A1(n18399), .A2(n11129), .ZN(n20412) );
  OAI21_X1 U20415 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n20412), .A(
        n18400), .ZN(n20416) );
  OAI21_X1 U20416 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18402), .A(
        n18401), .ZN(n21127) );
  OAI22_X1 U20417 ( .A1(n18460), .A2(n20416), .B1(n18468), .B2(n21127), .ZN(
        n18403) );
  AOI21_X1 U20418 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18415), .A(
        n18403), .ZN(n18404) );
  OAI211_X1 U20419 ( .C1(n21379), .C2(n20430), .A(n18405), .B(n18404), .ZN(
        P3_U2824) );
  OAI21_X1 U20420 ( .B1(n18408), .B2(n18407), .A(n18406), .ZN(n21119) );
  AOI21_X1 U20421 ( .B1(n18411), .B2(n18410), .A(n18409), .ZN(n21116) );
  AOI22_X1 U20422 ( .A1(n21401), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18457), 
        .B2(n21116), .ZN(n18417) );
  INV_X1 U20423 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20410) );
  OAI21_X1 U20424 ( .B1(n18439), .B2(n18412), .A(n20410), .ZN(n18414) );
  NAND2_X1 U20425 ( .A1(n18413), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18418) );
  AOI21_X1 U20426 ( .B1(n20410), .B2(n18418), .A(n20412), .ZN(n20402) );
  AOI22_X1 U20427 ( .A1(n18415), .A2(n18414), .B1(n20402), .B2(n18450), .ZN(
        n18416) );
  OAI211_X1 U20428 ( .C1(n18468), .C2(n21119), .A(n18417), .B(n18416), .ZN(
        P3_U2825) );
  NOR2_X1 U20429 ( .A1(n18421), .A2(n11129), .ZN(n18431) );
  OAI21_X1 U20430 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18431), .A(
        n18418), .ZN(n20385) );
  XOR2_X1 U20431 ( .A(n18420), .B(n18419), .Z(n21096) );
  INV_X1 U20432 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n20399) );
  NOR2_X1 U20433 ( .A1(n21379), .A2(n20399), .ZN(n21098) );
  NOR3_X1 U20434 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18421), .A3(
        n19054), .ZN(n18422) );
  AOI211_X1 U20435 ( .C1(n18423), .C2(n21096), .A(n21098), .B(n18422), .ZN(
        n18430) );
  AOI21_X1 U20436 ( .B1(n18426), .B2(n18425), .A(n18424), .ZN(n21103) );
  OAI21_X1 U20437 ( .B1(n18428), .B2(n18427), .A(n11018), .ZN(n18440) );
  AOI22_X1 U20438 ( .A1(n18457), .A2(n21103), .B1(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18440), .ZN(n18429) );
  OAI211_X1 U20439 ( .C1(n18460), .C2(n20385), .A(n18430), .B(n18429), .ZN(
        P3_U2826) );
  INV_X1 U20440 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n20363) );
  NOR2_X1 U20441 ( .A1(n20363), .A2(n11129), .ZN(n20366) );
  INV_X1 U20442 ( .A(n18431), .ZN(n20386) );
  OAI21_X1 U20443 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n20366), .A(
        n20386), .ZN(n20373) );
  AOI21_X1 U20444 ( .B1(n18434), .B2(n18433), .A(n18432), .ZN(n21093) );
  INV_X1 U20445 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n21090) );
  OAI21_X1 U20446 ( .B1(n18437), .B2(n18436), .A(n18435), .ZN(n21095) );
  OAI22_X1 U20447 ( .A1(n21379), .A2(n21090), .B1(n18468), .B2(n21095), .ZN(
        n18438) );
  AOI21_X1 U20448 ( .B1(n18457), .B2(n21093), .A(n18438), .ZN(n18442) );
  NOR2_X1 U20449 ( .A1(n18439), .A2(n20363), .ZN(n18446) );
  OAI21_X1 U20450 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18446), .A(
        n18440), .ZN(n18441) );
  OAI211_X1 U20451 ( .C1(n18460), .C2(n20373), .A(n18442), .B(n18441), .ZN(
        P3_U2827) );
  OAI21_X1 U20452 ( .B1(n18445), .B2(n18444), .A(n18443), .ZN(n21076) );
  AOI21_X1 U20453 ( .B1(n20363), .B2(n11129), .A(n20366), .ZN(n20358) );
  AOI21_X1 U20454 ( .B1(n20363), .B2(n19054), .A(n18446), .ZN(n18449) );
  AOI211_X1 U20455 ( .C1(n21078), .C2(n21077), .A(n18447), .B(n18467), .ZN(
        n18448) );
  AOI211_X1 U20456 ( .C1(n20358), .C2(n18450), .A(n18449), .B(n18448), .ZN(
        n18451) );
  NAND2_X1 U20457 ( .A1(n21401), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n21081) );
  OAI211_X1 U20458 ( .C1(n18468), .C2(n21076), .A(n18451), .B(n21081), .ZN(
        P3_U2828) );
  AOI21_X1 U20459 ( .B1(n18453), .B2(n18462), .A(n18452), .ZN(n21066) );
  AOI21_X1 U20460 ( .B1(n18455), .B2(n18461), .A(n18454), .ZN(n21070) );
  INV_X1 U20461 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n20357) );
  OAI22_X1 U20462 ( .A1(n21070), .A2(n18468), .B1(n21379), .B2(n20357), .ZN(
        n18456) );
  AOI21_X1 U20463 ( .B1(n18457), .B2(n21066), .A(n18456), .ZN(n18458) );
  OAI221_X1 U20464 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18460), .C1(
        n11129), .C2(n18459), .A(n18458), .ZN(P3_U2829) );
  NAND2_X1 U20465 ( .A1(n18462), .A2(n18461), .ZN(n21060) );
  INV_X1 U20466 ( .A(n21060), .ZN(n21059) );
  NAND3_X1 U20467 ( .A1(n20997), .A2(n18464), .A3(n11018), .ZN(n18465) );
  AOI22_X1 U20468 ( .A1(n21401), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18465), .ZN(n18466) );
  OAI221_X1 U20469 ( .B1(n21059), .B2(n18468), .C1(n21060), .C2(n18467), .A(
        n18466), .ZN(P3_U2830) );
  NAND3_X1 U20470 ( .A1(n18972), .A2(n18473), .A3(n18472), .ZN(n18470) );
  NAND2_X1 U20471 ( .A1(n18968), .A2(n21465), .ZN(n18999) );
  NAND2_X1 U20472 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18945) );
  NAND4_X1 U20473 ( .A1(n18979), .A2(n18999), .A3(n18473), .A4(n18945), .ZN(
        n18469) );
  OAI211_X1 U20474 ( .C1(n18471), .C2(n21465), .A(n18470), .B(n18469), .ZN(
        P3_U2866) );
  NAND2_X1 U20475 ( .A1(n18473), .A2(n18472), .ZN(n18477) );
  NOR4_X1 U20476 ( .A1(n18475), .A2(n18979), .A3(n18474), .A4(n21450), .ZN(
        n18476) );
  AOI21_X1 U20477 ( .B1(n21450), .B2(n18477), .A(n18476), .ZN(P3_U2864) );
  NOR4_X1 U20478 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18481) );
  NOR4_X1 U20479 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18480) );
  NOR4_X1 U20480 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18479) );
  NOR4_X1 U20481 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18478) );
  NAND4_X1 U20482 ( .A1(n18481), .A2(n18480), .A3(n18479), .A4(n18478), .ZN(
        n18487) );
  NOR4_X1 U20483 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18485) );
  AOI211_X1 U20484 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_31__SCAN_IN), .B(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n18484) );
  NOR4_X1 U20485 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18483) );
  NOR4_X1 U20486 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18482) );
  NAND4_X1 U20487 ( .A1(n18485), .A2(n18484), .A3(n18483), .A4(n18482), .ZN(
        n18486) );
  NOR2_X1 U20488 ( .A1(n18487), .A2(n18486), .ZN(n18495) );
  INV_X1 U20489 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18575) );
  OAI21_X1 U20490 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18495), .ZN(n18488) );
  OAI21_X1 U20491 ( .B1(n18495), .B2(n18575), .A(n18488), .ZN(P3_U3293) );
  INV_X1 U20492 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18579) );
  AOI21_X1 U20493 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18489) );
  OAI221_X1 U20494 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n18489), .C1(n20357), 
        .C2(P3_REIP_REG_0__SCAN_IN), .A(n18495), .ZN(n18490) );
  OAI21_X1 U20495 ( .B1(n18495), .B2(n18579), .A(n18490), .ZN(P3_U3292) );
  INV_X1 U20496 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18577) );
  NOR3_X1 U20497 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n18492) );
  OAI21_X1 U20498 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n18492), .A(n18495), .ZN(
        n18491) );
  OAI21_X1 U20499 ( .B1(n18495), .B2(n18577), .A(n18491), .ZN(P3_U2638) );
  INV_X1 U20500 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21825) );
  AOI21_X1 U20501 ( .B1(n20357), .B2(n21825), .A(n18492), .ZN(n18494) );
  INV_X1 U20502 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18581) );
  INV_X1 U20503 ( .A(n18495), .ZN(n18493) );
  AOI22_X1 U20504 ( .A1(n18495), .A2(n18494), .B1(n18581), .B2(n18493), .ZN(
        P3_U2639) );
  INV_X1 U20505 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n18582) );
  AOI22_X1 U20506 ( .A1(n21831), .A2(n18496), .B1(n18582), .B2(n18561), .ZN(
        P3_U3297) );
  INV_X1 U20507 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18497) );
  AOI22_X1 U20508 ( .A1(n21831), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18497), 
        .B2(n18561), .ZN(P3_U3294) );
  AOI22_X1 U20509 ( .A1(P3_D_C_N_REG_SCAN_IN), .A2(n18561), .B1(n21827), .B2(
        n21881), .ZN(n18498) );
  OAI21_X1 U20510 ( .B1(P3_CODEFETCH_REG_SCAN_IN), .B2(n18561), .A(n18498), 
        .ZN(P3_U2635) );
  INV_X1 U20511 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n20979) );
  AOI22_X1 U20512 ( .A1(n21489), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18532), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18499) );
  OAI21_X1 U20513 ( .B1(n20979), .B2(n18515), .A(n18499), .ZN(P3_U2767) );
  INV_X1 U20514 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n20829) );
  AOI22_X1 U20515 ( .A1(n21489), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18532), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18500) );
  OAI21_X1 U20516 ( .B1(n20829), .B2(n18515), .A(n18500), .ZN(P3_U2766) );
  INV_X1 U20517 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n20312) );
  AOI22_X1 U20518 ( .A1(n21489), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18525), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18501) );
  OAI21_X1 U20519 ( .B1(n20312), .B2(n18515), .A(n18501), .ZN(P3_U2765) );
  INV_X1 U20520 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n20830) );
  AOI22_X1 U20521 ( .A1(n21489), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18525), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18502) );
  OAI21_X1 U20522 ( .B1(n20830), .B2(n18515), .A(n18502), .ZN(P3_U2764) );
  INV_X1 U20523 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n20315) );
  AOI22_X1 U20524 ( .A1(n21489), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18525), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18503) );
  OAI21_X1 U20525 ( .B1(n20315), .B2(n18515), .A(n18503), .ZN(P3_U2763) );
  INV_X1 U20526 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n20831) );
  AOI22_X1 U20527 ( .A1(n21489), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18525), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18504) );
  OAI21_X1 U20528 ( .B1(n20831), .B2(n18515), .A(n18504), .ZN(P3_U2762) );
  INV_X1 U20529 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n20318) );
  AOI22_X1 U20530 ( .A1(n21489), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18525), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18505) );
  OAI21_X1 U20531 ( .B1(n20318), .B2(n18515), .A(n18505), .ZN(P3_U2761) );
  INV_X1 U20532 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n20800) );
  AOI22_X1 U20533 ( .A1(n21489), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18532), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18506) );
  OAI21_X1 U20534 ( .B1(n20800), .B2(n18515), .A(n18506), .ZN(P3_U2760) );
  INV_X1 U20535 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n20975) );
  AOI22_X1 U20536 ( .A1(n20279), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18532), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18507) );
  OAI21_X1 U20537 ( .B1(n20975), .B2(n18515), .A(n18507), .ZN(P3_U2759) );
  INV_X1 U20538 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n20322) );
  AOI22_X1 U20539 ( .A1(n20279), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18532), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18508) );
  OAI21_X1 U20540 ( .B1(n20322), .B2(n18515), .A(n18508), .ZN(P3_U2758) );
  INV_X1 U20541 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n20324) );
  AOI22_X1 U20542 ( .A1(n20279), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18532), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18509) );
  OAI21_X1 U20543 ( .B1(n20324), .B2(n18515), .A(n18509), .ZN(P3_U2757) );
  INV_X1 U20544 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n20802) );
  AOI22_X1 U20545 ( .A1(n20279), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18532), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18510) );
  OAI21_X1 U20546 ( .B1(n20802), .B2(n18515), .A(n18510), .ZN(P3_U2756) );
  INV_X1 U20547 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n20327) );
  AOI22_X1 U20548 ( .A1(n20279), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18532), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18511) );
  OAI21_X1 U20549 ( .B1(n20327), .B2(n18515), .A(n18511), .ZN(P3_U2755) );
  INV_X1 U20550 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n20330) );
  AOI22_X1 U20551 ( .A1(n20279), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18532), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18512) );
  OAI21_X1 U20552 ( .B1(n20330), .B2(n18515), .A(n18512), .ZN(P3_U2754) );
  INV_X1 U20553 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n20960) );
  AOI22_X1 U20554 ( .A1(n20279), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18532), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18513) );
  OAI21_X1 U20555 ( .B1(n20960), .B2(n18515), .A(n18513), .ZN(P3_U2753) );
  INV_X1 U20556 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n20336) );
  AOI22_X1 U20557 ( .A1(n20279), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18532), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18514) );
  OAI21_X1 U20558 ( .B1(n20336), .B2(n18515), .A(n18514), .ZN(P3_U2752) );
  INV_X1 U20559 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n20952) );
  NAND2_X1 U20560 ( .A1(n18516), .A2(n20340), .ZN(n18534) );
  AOI22_X1 U20561 ( .A1(n20279), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18532), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18517) );
  OAI21_X1 U20562 ( .B1(n20952), .B2(n18534), .A(n18517), .ZN(P3_U2751) );
  INV_X1 U20563 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n20890) );
  AOI22_X1 U20564 ( .A1(n20279), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18532), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18518) );
  OAI21_X1 U20565 ( .B1(n20890), .B2(n18534), .A(n18518), .ZN(P3_U2750) );
  INV_X1 U20566 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n20289) );
  AOI22_X1 U20567 ( .A1(n20279), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18532), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18519) );
  OAI21_X1 U20568 ( .B1(n20289), .B2(n18534), .A(n18519), .ZN(P3_U2749) );
  INV_X1 U20569 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n20291) );
  AOI22_X1 U20570 ( .A1(n20279), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18532), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18520) );
  OAI21_X1 U20571 ( .B1(n20291), .B2(n18534), .A(n18520), .ZN(P3_U2748) );
  INV_X1 U20572 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n20293) );
  AOI22_X1 U20573 ( .A1(n20279), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18525), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18521) );
  OAI21_X1 U20574 ( .B1(n20293), .B2(n18534), .A(n18521), .ZN(P3_U2747) );
  INV_X1 U20575 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n20860) );
  AOI22_X1 U20576 ( .A1(n20279), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18525), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18522) );
  OAI21_X1 U20577 ( .B1(n20860), .B2(n18534), .A(n18522), .ZN(P3_U2746) );
  INV_X1 U20578 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n20296) );
  AOI22_X1 U20579 ( .A1(n20279), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18525), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18523) );
  OAI21_X1 U20580 ( .B1(n20296), .B2(n18534), .A(n18523), .ZN(P3_U2745) );
  INV_X1 U20581 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n20943) );
  AOI22_X1 U20582 ( .A1(n20279), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18525), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18524) );
  OAI21_X1 U20583 ( .B1(n20943), .B2(n18534), .A(n18524), .ZN(P3_U2744) );
  INV_X1 U20584 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n20936) );
  AOI22_X1 U20585 ( .A1(n20279), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18525), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18526) );
  OAI21_X1 U20586 ( .B1(n20936), .B2(n18534), .A(n18526), .ZN(P3_U2743) );
  INV_X1 U20587 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n20896) );
  AOI22_X1 U20588 ( .A1(n20279), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18532), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18527) );
  OAI21_X1 U20589 ( .B1(n20896), .B2(n18534), .A(n18527), .ZN(P3_U2742) );
  INV_X1 U20590 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n20302) );
  AOI22_X1 U20591 ( .A1(n20279), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18532), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18528) );
  OAI21_X1 U20592 ( .B1(n20302), .B2(n18534), .A(n18528), .ZN(P3_U2741) );
  INV_X1 U20593 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n20929) );
  AOI22_X1 U20594 ( .A1(n20279), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18532), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18529) );
  OAI21_X1 U20595 ( .B1(n20929), .B2(n18534), .A(n18529), .ZN(P3_U2740) );
  INV_X1 U20596 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n20305) );
  AOI22_X1 U20597 ( .A1(n20279), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18532), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18530) );
  OAI21_X1 U20598 ( .B1(n20305), .B2(n18534), .A(n18530), .ZN(P3_U2739) );
  INV_X1 U20599 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n20307) );
  AOI22_X1 U20600 ( .A1(n20279), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18532), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18531) );
  OAI21_X1 U20601 ( .B1(n20307), .B2(n18534), .A(n18531), .ZN(P3_U2738) );
  INV_X1 U20602 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n20915) );
  AOI22_X1 U20603 ( .A1(n20279), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18532), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18533) );
  OAI21_X1 U20604 ( .B1(n20915), .B2(n18534), .A(n18533), .ZN(P3_U2737) );
  NOR2_X1 U20605 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(n18535), .ZN(n18536) );
  NOR2_X1 U20606 ( .A1(n21831), .A2(n18536), .ZN(P3_U2633) );
  NOR2_X1 U20607 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n18561), .ZN(n18569) );
  INV_X1 U20608 ( .A(n18569), .ZN(n18573) );
  AOI22_X1 U20609 ( .A1(n18567), .A2(P3_REIP_REG_2__SCAN_IN), .B1(
        P3_ADDRESS_REG_0__SCAN_IN), .B2(n18561), .ZN(n18537) );
  OAI21_X1 U20610 ( .B1(n18553), .B2(n20357), .A(n18537), .ZN(P3_U3032) );
  AOI22_X1 U20611 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n18571), .B1(
        P3_ADDRESS_REG_1__SCAN_IN), .B2(n18561), .ZN(n18538) );
  OAI21_X1 U20612 ( .B1(n21090), .B2(n18573), .A(n18538), .ZN(P3_U3033) );
  AOI22_X1 U20613 ( .A1(n18567), .A2(P3_REIP_REG_4__SCAN_IN), .B1(
        P3_ADDRESS_REG_2__SCAN_IN), .B2(n18561), .ZN(n18539) );
  OAI21_X1 U20614 ( .B1(n18553), .B2(n21090), .A(n18539), .ZN(P3_U3034) );
  AOI22_X1 U20615 ( .A1(n18567), .A2(P3_REIP_REG_5__SCAN_IN), .B1(
        P3_ADDRESS_REG_3__SCAN_IN), .B2(n18561), .ZN(n18540) );
  OAI21_X1 U20616 ( .B1(n18553), .B2(n20399), .A(n18540), .ZN(P3_U3035) );
  AOI22_X1 U20617 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n18571), .B1(
        P3_ADDRESS_REG_4__SCAN_IN), .B2(n18561), .ZN(n18541) );
  OAI21_X1 U20618 ( .B1(n20430), .B2(n18573), .A(n18541), .ZN(P3_U3036) );
  AOI22_X1 U20619 ( .A1(n18567), .A2(P3_REIP_REG_7__SCAN_IN), .B1(
        P3_ADDRESS_REG_5__SCAN_IN), .B2(n18561), .ZN(n18542) );
  OAI21_X1 U20620 ( .B1(n18553), .B2(n20430), .A(n18542), .ZN(P3_U3037) );
  AOI22_X1 U20621 ( .A1(n18567), .A2(P3_REIP_REG_8__SCAN_IN), .B1(
        P3_ADDRESS_REG_6__SCAN_IN), .B2(n18561), .ZN(n18543) );
  OAI21_X1 U20622 ( .B1(n18553), .B2(n21128), .A(n18543), .ZN(P3_U3038) );
  INV_X1 U20623 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n20442) );
  AOI22_X1 U20624 ( .A1(n18567), .A2(P3_REIP_REG_9__SCAN_IN), .B1(
        P3_ADDRESS_REG_7__SCAN_IN), .B2(n18561), .ZN(n18544) );
  OAI21_X1 U20625 ( .B1(n18553), .B2(n20442), .A(n18544), .ZN(P3_U3039) );
  AOI22_X1 U20626 ( .A1(n18567), .A2(P3_REIP_REG_10__SCAN_IN), .B1(
        P3_ADDRESS_REG_8__SCAN_IN), .B2(n18561), .ZN(n18545) );
  OAI21_X1 U20627 ( .B1(n18553), .B2(n18546), .A(n18545), .ZN(P3_U3040) );
  INV_X1 U20628 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n20477) );
  AOI22_X1 U20629 ( .A1(n18567), .A2(P3_REIP_REG_11__SCAN_IN), .B1(
        P3_ADDRESS_REG_9__SCAN_IN), .B2(n18561), .ZN(n18547) );
  OAI21_X1 U20630 ( .B1(n18553), .B2(n20477), .A(n18547), .ZN(P3_U3041) );
  INV_X1 U20631 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n20476) );
  AOI22_X1 U20632 ( .A1(n18567), .A2(P3_REIP_REG_12__SCAN_IN), .B1(
        P3_ADDRESS_REG_10__SCAN_IN), .B2(n18561), .ZN(n18548) );
  OAI21_X1 U20633 ( .B1(n18553), .B2(n20476), .A(n18548), .ZN(P3_U3042) );
  INV_X1 U20634 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n20524) );
  AOI22_X1 U20635 ( .A1(n18567), .A2(P3_REIP_REG_13__SCAN_IN), .B1(
        P3_ADDRESS_REG_11__SCAN_IN), .B2(n18561), .ZN(n18549) );
  OAI21_X1 U20636 ( .B1(n18553), .B2(n20524), .A(n18549), .ZN(P3_U3043) );
  INV_X1 U20637 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n20525) );
  AOI22_X1 U20638 ( .A1(n18567), .A2(P3_REIP_REG_14__SCAN_IN), .B1(
        P3_ADDRESS_REG_12__SCAN_IN), .B2(n18561), .ZN(n18550) );
  OAI21_X1 U20639 ( .B1(n18553), .B2(n20525), .A(n18550), .ZN(P3_U3044) );
  AOI22_X1 U20640 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n18571), .B1(
        P3_ADDRESS_REG_13__SCAN_IN), .B2(n18561), .ZN(n18551) );
  OAI21_X1 U20641 ( .B1(n20550), .B2(n18573), .A(n18551), .ZN(P3_U3045) );
  AOI22_X1 U20642 ( .A1(n18567), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_ADDRESS_REG_14__SCAN_IN), .B2(n18561), .ZN(n18552) );
  OAI21_X1 U20643 ( .B1(n18553), .B2(n20550), .A(n18552), .ZN(P3_U3046) );
  AOI22_X1 U20644 ( .A1(n18569), .A2(P3_REIP_REG_17__SCAN_IN), .B1(
        P3_ADDRESS_REG_15__SCAN_IN), .B2(n18561), .ZN(n18554) );
  OAI21_X1 U20645 ( .B1(n18553), .B2(n20551), .A(n18554), .ZN(P3_U3047) );
  AOI22_X1 U20646 ( .A1(n18569), .A2(P3_REIP_REG_18__SCAN_IN), .B1(
        P3_ADDRESS_REG_16__SCAN_IN), .B2(n18561), .ZN(n18555) );
  OAI21_X1 U20647 ( .B1(n18553), .B2(n20573), .A(n18555), .ZN(P3_U3048) );
  AOI22_X1 U20648 ( .A1(n18569), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_ADDRESS_REG_17__SCAN_IN), .B2(n18561), .ZN(n18556) );
  OAI21_X1 U20649 ( .B1(n18553), .B2(n21378), .A(n18556), .ZN(P3_U3049) );
  INV_X1 U20650 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n20611) );
  AOI22_X1 U20651 ( .A1(n18569), .A2(P3_REIP_REG_20__SCAN_IN), .B1(
        P3_ADDRESS_REG_18__SCAN_IN), .B2(n18561), .ZN(n18557) );
  OAI21_X1 U20652 ( .B1(n18553), .B2(n20611), .A(n18557), .ZN(P3_U3050) );
  INV_X1 U20653 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n20625) );
  AOI22_X1 U20654 ( .A1(n18569), .A2(P3_REIP_REG_21__SCAN_IN), .B1(
        P3_ADDRESS_REG_19__SCAN_IN), .B2(n18561), .ZN(n18558) );
  OAI21_X1 U20655 ( .B1(n18553), .B2(n20625), .A(n18558), .ZN(P3_U3051) );
  INV_X1 U20656 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n20636) );
  AOI22_X1 U20657 ( .A1(n18569), .A2(P3_REIP_REG_22__SCAN_IN), .B1(
        P3_ADDRESS_REG_20__SCAN_IN), .B2(n18561), .ZN(n18559) );
  OAI21_X1 U20658 ( .B1(n18553), .B2(n20636), .A(n18559), .ZN(P3_U3052) );
  INV_X1 U20659 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n20651) );
  AOI22_X1 U20660 ( .A1(n18569), .A2(P3_REIP_REG_23__SCAN_IN), .B1(
        P3_ADDRESS_REG_21__SCAN_IN), .B2(n18561), .ZN(n18560) );
  OAI21_X1 U20661 ( .B1(n18553), .B2(n20651), .A(n18560), .ZN(P3_U3053) );
  INV_X1 U20662 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n20663) );
  AOI22_X1 U20663 ( .A1(n18569), .A2(P3_REIP_REG_24__SCAN_IN), .B1(
        P3_ADDRESS_REG_22__SCAN_IN), .B2(n18561), .ZN(n18562) );
  OAI21_X1 U20664 ( .B1(n18553), .B2(n20663), .A(n18562), .ZN(P3_U3054) );
  AOI22_X1 U20665 ( .A1(n18569), .A2(P3_REIP_REG_25__SCAN_IN), .B1(
        P3_ADDRESS_REG_23__SCAN_IN), .B2(n18561), .ZN(n18563) );
  OAI21_X1 U20666 ( .B1(n18553), .B2(n20678), .A(n18563), .ZN(P3_U3055) );
  INV_X1 U20667 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n20693) );
  AOI22_X1 U20668 ( .A1(n18567), .A2(P3_REIP_REG_26__SCAN_IN), .B1(
        P3_ADDRESS_REG_24__SCAN_IN), .B2(n18561), .ZN(n18564) );
  OAI21_X1 U20669 ( .B1(n18553), .B2(n20693), .A(n18564), .ZN(P3_U3056) );
  AOI22_X1 U20670 ( .A1(n18567), .A2(P3_REIP_REG_27__SCAN_IN), .B1(
        P3_ADDRESS_REG_25__SCAN_IN), .B2(n18561), .ZN(n18565) );
  OAI21_X1 U20671 ( .B1(n18553), .B2(n20707), .A(n18565), .ZN(P3_U3057) );
  AOI22_X1 U20672 ( .A1(n18567), .A2(P3_REIP_REG_28__SCAN_IN), .B1(
        P3_ADDRESS_REG_26__SCAN_IN), .B2(n18561), .ZN(n18566) );
  OAI21_X1 U20673 ( .B1(n18553), .B2(n20721), .A(n18566), .ZN(P3_U3058) );
  INV_X1 U20674 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n21317) );
  AOI22_X1 U20675 ( .A1(n18567), .A2(P3_REIP_REG_29__SCAN_IN), .B1(
        P3_ADDRESS_REG_27__SCAN_IN), .B2(n18561), .ZN(n18568) );
  OAI21_X1 U20676 ( .B1(n18553), .B2(n21317), .A(n18568), .ZN(P3_U3059) );
  INV_X1 U20677 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n20746) );
  AOI22_X1 U20678 ( .A1(n18569), .A2(P3_REIP_REG_30__SCAN_IN), .B1(
        P3_ADDRESS_REG_28__SCAN_IN), .B2(n18561), .ZN(n18570) );
  OAI21_X1 U20679 ( .B1(n18553), .B2(n20746), .A(n18570), .ZN(P3_U3060) );
  AOI22_X1 U20680 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n18571), .B1(
        P3_ADDRESS_REG_29__SCAN_IN), .B2(n18561), .ZN(n18572) );
  OAI21_X1 U20681 ( .B1(n20761), .B2(n18573), .A(n18572), .ZN(P3_U3061) );
  INV_X1 U20682 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18574) );
  AOI22_X1 U20683 ( .A1(n21831), .A2(n18575), .B1(n18574), .B2(n18561), .ZN(
        P3_U3277) );
  INV_X1 U20684 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n18576) );
  AOI22_X1 U20685 ( .A1(n21831), .A2(n18577), .B1(n18576), .B2(n18561), .ZN(
        P3_U3276) );
  INV_X1 U20686 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n18578) );
  AOI22_X1 U20687 ( .A1(n21831), .A2(n18579), .B1(n18578), .B2(n18561), .ZN(
        P3_U3275) );
  INV_X1 U20688 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n18580) );
  AOI22_X1 U20689 ( .A1(n21831), .A2(n18581), .B1(n18580), .B2(n18561), .ZN(
        P3_U3274) );
  NOR4_X1 U20690 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_BE_N_REG_2__SCAN_IN), .A4(P3_BE_N_REG_0__SCAN_IN), .ZN(n18584)
         );
  NOR4_X1 U20691 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(P3_D_C_N_REG_SCAN_IN), .A3(
        P3_W_R_N_REG_SCAN_IN), .A4(n18582), .ZN(n18583) );
  NAND3_X1 U20692 ( .A1(n18584), .A2(n18583), .A3(U215), .ZN(U213) );
  NOR2_X1 U20693 ( .A1(n21850), .A2(n19470), .ZN(n18588) );
  OAI21_X1 U20694 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n11969), .A(n21857), 
        .ZN(n18586) );
  NAND3_X1 U20695 ( .A1(n18586), .A2(n18585), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n18587) );
  OAI21_X1 U20696 ( .B1(n18588), .B2(n18909), .A(n18587), .ZN(n18594) );
  NAND4_X1 U20697 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .A3(n11407), .A4(n18908), .ZN(n18590) );
  OAI211_X1 U20698 ( .C1(n18592), .C2(n18591), .A(n18590), .B(n18589), .ZN(
        n18593) );
  MUX2_X1 U20699 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .B(n18594), .S(n18593), 
        .Z(P2_U3610) );
  INV_X1 U20700 ( .A(n18595), .ZN(n18606) );
  AOI22_X1 U20701 ( .A1(n18763), .A2(n18875), .B1(n18850), .B2(
        P2_REIP_REG_0__SCAN_IN), .ZN(n18597) );
  NAND2_X1 U20702 ( .A1(n18852), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n18596) );
  OAI211_X1 U20703 ( .C1(n18598), .C2(n18803), .A(n18597), .B(n18596), .ZN(
        n18599) );
  AOI21_X1 U20704 ( .B1(n18600), .B2(n18811), .A(n18599), .ZN(n18604) );
  AOI21_X1 U20705 ( .B1(n18621), .B2(n18776), .A(n18601), .ZN(n18602) );
  AOI21_X1 U20706 ( .B1(n18614), .B2(n19467), .A(n18602), .ZN(n18603) );
  OAI211_X1 U20707 ( .C1(n18606), .C2(n18605), .A(n18604), .B(n18603), .ZN(
        P2_U2855) );
  AOI22_X1 U20708 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18851), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n18850), .ZN(n18607) );
  OAI21_X1 U20709 ( .B1(n18803), .B2(n18608), .A(n18607), .ZN(n18609) );
  AOI21_X1 U20710 ( .B1(P2_EBX_REG_1__SCAN_IN), .B2(n18852), .A(n18609), .ZN(
        n18610) );
  OAI21_X1 U20711 ( .B1(n18611), .B2(n18855), .A(n18610), .ZN(n18612) );
  AOI21_X1 U20712 ( .B1(n18613), .B2(n18811), .A(n18612), .ZN(n18617) );
  AOI22_X1 U20713 ( .A1(n18615), .A2(n18861), .B1(n18614), .B2(n19423), .ZN(
        n18616) );
  OAI211_X1 U20714 ( .C1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n18776), .A(
        n18617), .B(n18616), .ZN(P2_U2854) );
  NOR2_X1 U20715 ( .A1(n18717), .A2(n18618), .ZN(n18619) );
  XOR2_X1 U20716 ( .A(n18620), .B(n18619), .Z(n18632) );
  INV_X1 U20717 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18622) );
  OAI22_X1 U20718 ( .A1(n18623), .A2(n18803), .B1(n18622), .B2(n18621), .ZN(
        n18624) );
  INV_X1 U20719 ( .A(n18624), .ZN(n18625) );
  OAI211_X1 U20720 ( .C1(n18626), .C2(n18748), .A(n18625), .B(n18746), .ZN(
        n18630) );
  OAI22_X1 U20721 ( .A1(n18628), .A2(n18855), .B1(n18857), .B2(n18627), .ZN(
        n18629) );
  AOI211_X1 U20722 ( .C1(P2_EBX_REG_6__SCAN_IN), .C2(n18852), .A(n18630), .B(
        n18629), .ZN(n18631) );
  OAI21_X1 U20723 ( .B1(n18897), .B2(n18632), .A(n18631), .ZN(P2_U2849) );
  NAND2_X1 U20724 ( .A1(n18752), .A2(n18633), .ZN(n18635) );
  XOR2_X1 U20725 ( .A(n18635), .B(n18634), .Z(n18644) );
  AOI22_X1 U20726 ( .A1(n18636), .A2(n18853), .B1(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18851), .ZN(n18637) );
  OAI211_X1 U20727 ( .C1(n18638), .C2(n18748), .A(n18637), .B(n18746), .ZN(
        n18642) );
  OAI22_X1 U20728 ( .A1(n18640), .A2(n18855), .B1(n18639), .B2(n18857), .ZN(
        n18641) );
  AOI211_X1 U20729 ( .C1(P2_EBX_REG_7__SCAN_IN), .C2(n18852), .A(n18642), .B(
        n18641), .ZN(n18643) );
  OAI21_X1 U20730 ( .B1(n18644), .B2(n18897), .A(n18643), .ZN(P2_U2848) );
  AOI22_X1 U20731 ( .A1(n18645), .A2(n18853), .B1(P2_EBX_REG_8__SCAN_IN), .B2(
        n18852), .ZN(n18646) );
  OAI211_X1 U20732 ( .C1(n18647), .C2(n18748), .A(n18646), .B(n18746), .ZN(
        n18648) );
  AOI21_X1 U20733 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18851), .A(
        n18648), .ZN(n18656) );
  NOR2_X1 U20734 ( .A1(n18717), .A2(n18649), .ZN(n18651) );
  XNOR2_X1 U20735 ( .A(n18651), .B(n18650), .ZN(n18654) );
  INV_X1 U20736 ( .A(n18652), .ZN(n18653) );
  AOI22_X1 U20737 ( .A1(n18654), .A2(n18861), .B1(n18653), .B2(n18811), .ZN(
        n18655) );
  OAI211_X1 U20738 ( .C1(n18855), .C2(n18657), .A(n18656), .B(n18655), .ZN(
        P2_U2847) );
  AOI22_X1 U20739 ( .A1(n18658), .A2(n18853), .B1(P2_EBX_REG_10__SCAN_IN), 
        .B2(n18852), .ZN(n18659) );
  OAI211_X1 U20740 ( .C1(n18660), .C2(n18748), .A(n18659), .B(n18746), .ZN(
        n18661) );
  AOI21_X1 U20741 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18851), .A(
        n18661), .ZN(n18668) );
  NOR2_X1 U20742 ( .A1(n18717), .A2(n18662), .ZN(n18664) );
  XNOR2_X1 U20743 ( .A(n18664), .B(n18663), .ZN(n18666) );
  AOI22_X1 U20744 ( .A1(n18666), .A2(n18861), .B1(n18665), .B2(n18811), .ZN(
        n18667) );
  OAI211_X1 U20745 ( .C1(n18669), .C2(n18855), .A(n18668), .B(n18667), .ZN(
        P2_U2845) );
  AOI22_X1 U20746 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18851), .B1(
        P2_EBX_REG_12__SCAN_IN), .B2(n18852), .ZN(n18670) );
  OAI21_X1 U20747 ( .B1(n18671), .B2(n18803), .A(n18670), .ZN(n18672) );
  AOI211_X1 U20748 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n18850), .A(n16976), 
        .B(n18672), .ZN(n18679) );
  NOR2_X1 U20749 ( .A1(n18717), .A2(n18673), .ZN(n18675) );
  XNOR2_X1 U20750 ( .A(n18675), .B(n18674), .ZN(n18677) );
  AOI22_X1 U20751 ( .A1(n18677), .A2(n18861), .B1(n18676), .B2(n18811), .ZN(
        n18678) );
  OAI211_X1 U20752 ( .C1(n18680), .C2(n18855), .A(n18679), .B(n18678), .ZN(
        P2_U2843) );
  AOI22_X1 U20753 ( .A1(P2_EBX_REG_14__SCAN_IN), .A2(n18852), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n18851), .ZN(n18681) );
  OAI21_X1 U20754 ( .B1(n18682), .B2(n18803), .A(n18681), .ZN(n18683) );
  AOI211_X1 U20755 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n18850), .A(n16976), 
        .B(n18683), .ZN(n18690) );
  NOR2_X1 U20756 ( .A1(n18717), .A2(n18684), .ZN(n18686) );
  XNOR2_X1 U20757 ( .A(n18686), .B(n18685), .ZN(n18688) );
  AOI22_X1 U20758 ( .A1(n18688), .A2(n18861), .B1(n18687), .B2(n18811), .ZN(
        n18689) );
  OAI211_X1 U20759 ( .C1(n19363), .C2(n18855), .A(n18690), .B(n18689), .ZN(
        P2_U2841) );
  NAND2_X1 U20760 ( .A1(n18752), .A2(n18691), .ZN(n18692) );
  XOR2_X1 U20761 ( .A(n18693), .B(n18692), .Z(n18703) );
  INV_X1 U20762 ( .A(n18694), .ZN(n18696) );
  AOI22_X1 U20763 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(n18852), .B1(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18851), .ZN(n18695) );
  OAI21_X1 U20764 ( .B1(n18696), .B2(n18803), .A(n18695), .ZN(n18697) );
  AOI211_X1 U20765 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n18850), .A(n16976), 
        .B(n18697), .ZN(n18702) );
  OAI22_X1 U20766 ( .A1(n18699), .A2(n18857), .B1(n18698), .B2(n18855), .ZN(
        n18700) );
  INV_X1 U20767 ( .A(n18700), .ZN(n18701) );
  OAI211_X1 U20768 ( .C1(n18897), .C2(n18703), .A(n18702), .B(n18701), .ZN(
        P2_U2840) );
  AOI22_X1 U20769 ( .A1(n18704), .A2(n18853), .B1(P2_EBX_REG_16__SCAN_IN), 
        .B2(n18852), .ZN(n18705) );
  OAI211_X1 U20770 ( .C1(n18706), .C2(n18748), .A(n18705), .B(n18746), .ZN(
        n18707) );
  AOI21_X1 U20771 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18851), .A(
        n18707), .ZN(n18714) );
  NOR2_X1 U20772 ( .A1(n18717), .A2(n18708), .ZN(n18710) );
  XNOR2_X1 U20773 ( .A(n18710), .B(n18709), .ZN(n18712) );
  AOI22_X1 U20774 ( .A1(n18712), .A2(n18861), .B1(n18711), .B2(n18811), .ZN(
        n18713) );
  OAI211_X1 U20775 ( .C1(n18715), .C2(n18855), .A(n18714), .B(n18713), .ZN(
        P2_U2839) );
  INV_X1 U20776 ( .A(n18719), .ZN(n18731) );
  OR2_X1 U20777 ( .A1(n18717), .A2(n18716), .ZN(n18738) );
  AOI211_X1 U20778 ( .C1(n18719), .C2(n18718), .A(n18897), .B(n18738), .ZN(
        n18725) );
  NAND2_X1 U20779 ( .A1(n18720), .A2(n18853), .ZN(n18723) );
  AOI22_X1 U20780 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n18851), .B1(
        P2_REIP_REG_17__SCAN_IN), .B2(n18850), .ZN(n18722) );
  NAND2_X1 U20781 ( .A1(n18852), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n18721) );
  NAND4_X1 U20782 ( .A1(n18723), .A2(n18722), .A3(n18746), .A4(n18721), .ZN(
        n18724) );
  NOR2_X1 U20783 ( .A1(n18725), .A2(n18724), .ZN(n18730) );
  INV_X1 U20784 ( .A(n18726), .ZN(n18727) );
  AOI22_X1 U20785 ( .A1(n18728), .A2(n18811), .B1(n18763), .B2(n18727), .ZN(
        n18729) );
  OAI211_X1 U20786 ( .C1(n18731), .C2(n18776), .A(n18730), .B(n18729), .ZN(
        P2_U2838) );
  OAI21_X1 U20787 ( .B1(n18732), .B2(n18748), .A(n18746), .ZN(n18736) );
  OAI22_X1 U20788 ( .A1(n18734), .A2(n18803), .B1(n18733), .B2(n11889), .ZN(
        n18735) );
  AOI211_X1 U20789 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n18851), .A(
        n18736), .B(n18735), .ZN(n18743) );
  XOR2_X1 U20790 ( .A(n18738), .B(n18737), .Z(n18741) );
  INV_X1 U20791 ( .A(n18739), .ZN(n18740) );
  AOI22_X1 U20792 ( .A1(n18741), .A2(n18861), .B1(n18740), .B2(n18811), .ZN(
        n18742) );
  OAI211_X1 U20793 ( .C1(n18744), .C2(n18855), .A(n18743), .B(n18742), .ZN(
        P2_U2837) );
  AOI22_X1 U20794 ( .A1(n18745), .A2(n18853), .B1(P2_EBX_REG_19__SCAN_IN), 
        .B2(n18852), .ZN(n18747) );
  OAI211_X1 U20795 ( .C1(n18749), .C2(n18748), .A(n18747), .B(n18746), .ZN(
        n18750) );
  AOI21_X1 U20796 ( .B1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18851), .A(
        n18750), .ZN(n18758) );
  NAND2_X1 U20797 ( .A1(n18752), .A2(n18751), .ZN(n18754) );
  XNOR2_X1 U20798 ( .A(n18754), .B(n18753), .ZN(n18756) );
  AOI22_X1 U20799 ( .A1(n18756), .A2(n18861), .B1(n18755), .B2(n18811), .ZN(
        n18757) );
  OAI211_X1 U20800 ( .C1(n18759), .C2(n18855), .A(n18758), .B(n18757), .ZN(
        P2_U2836) );
  NAND2_X1 U20801 ( .A1(n18852), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n18765) );
  AOI22_X1 U20802 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18851), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n18850), .ZN(n18760) );
  INV_X1 U20803 ( .A(n18760), .ZN(n18761) );
  AOI21_X1 U20804 ( .B1(n18763), .B2(n18762), .A(n18761), .ZN(n18764) );
  AND2_X1 U20805 ( .A1(n18765), .A2(n18764), .ZN(n18768) );
  NAND2_X1 U20806 ( .A1(n18766), .A2(n18853), .ZN(n18767) );
  OAI211_X1 U20807 ( .C1(n18769), .C2(n18857), .A(n18768), .B(n18767), .ZN(
        n18770) );
  INV_X1 U20808 ( .A(n18770), .ZN(n18774) );
  OAI211_X1 U20809 ( .C1(n18772), .C2(n18775), .A(n18771), .B(n18861), .ZN(
        n18773) );
  OAI211_X1 U20810 ( .C1(n18776), .C2(n18775), .A(n18774), .B(n18773), .ZN(
        P2_U2835) );
  AOI22_X1 U20811 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n18851), .B1(
        P2_REIP_REG_21__SCAN_IN), .B2(n18850), .ZN(n18789) );
  AOI22_X1 U20812 ( .A1(n18777), .A2(n18853), .B1(P2_EBX_REG_21__SCAN_IN), 
        .B2(n18852), .ZN(n18788) );
  OAI22_X1 U20813 ( .A1(n18779), .A2(n18857), .B1(n18778), .B2(n18855), .ZN(
        n18780) );
  INV_X1 U20814 ( .A(n18780), .ZN(n18787) );
  AOI22_X1 U20815 ( .A1(n18784), .A2(n18783), .B1(n18782), .B2(n18781), .ZN(
        n18785) );
  NAND2_X1 U20816 ( .A1(n18861), .A2(n18785), .ZN(n18786) );
  NAND4_X1 U20817 ( .A1(n18789), .A2(n18788), .A3(n18787), .A4(n18786), .ZN(
        P2_U2834) );
  AOI22_X1 U20818 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18851), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n18850), .ZN(n18801) );
  AOI22_X1 U20819 ( .A1(n18790), .A2(n18853), .B1(P2_EBX_REG_23__SCAN_IN), 
        .B2(n18852), .ZN(n18800) );
  OAI22_X1 U20820 ( .A1(n18792), .A2(n18857), .B1(n18791), .B2(n18855), .ZN(
        n18793) );
  INV_X1 U20821 ( .A(n18793), .ZN(n18799) );
  AOI21_X1 U20822 ( .B1(n18796), .B2(n18795), .A(n18794), .ZN(n18797) );
  NAND2_X1 U20823 ( .A1(n18861), .A2(n18797), .ZN(n18798) );
  NAND4_X1 U20824 ( .A1(n18801), .A2(n18800), .A3(n18799), .A4(n18798), .ZN(
        P2_U2832) );
  AOI22_X1 U20825 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18851), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n18850), .ZN(n18802) );
  OAI21_X1 U20826 ( .B1(n18804), .B2(n18803), .A(n18802), .ZN(n18805) );
  AOI21_X1 U20827 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n18852), .A(n18805), .ZN(
        n18813) );
  AOI211_X1 U20828 ( .C1(n18808), .C2(n18807), .A(n18806), .B(n18897), .ZN(
        n18809) );
  AOI21_X1 U20829 ( .B1(n18811), .B2(n18810), .A(n18809), .ZN(n18812) );
  OAI211_X1 U20830 ( .C1(n18814), .C2(n18855), .A(n18813), .B(n18812), .ZN(
        P2_U2831) );
  AOI22_X1 U20831 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n18851), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n18850), .ZN(n18827) );
  AOI22_X1 U20832 ( .A1(n18815), .A2(n18853), .B1(P2_EBX_REG_25__SCAN_IN), 
        .B2(n18852), .ZN(n18826) );
  INV_X1 U20833 ( .A(n18816), .ZN(n18817) );
  OAI22_X1 U20834 ( .A1(n18818), .A2(n18857), .B1(n18817), .B2(n18855), .ZN(
        n18819) );
  INV_X1 U20835 ( .A(n18819), .ZN(n18825) );
  INV_X1 U20836 ( .A(n18823), .ZN(n18821) );
  INV_X1 U20837 ( .A(n18822), .ZN(n18820) );
  OAI221_X1 U20838 ( .B1(n18823), .B2(n18822), .C1(n18821), .C2(n18820), .A(
        n18861), .ZN(n18824) );
  NAND4_X1 U20839 ( .A1(n18827), .A2(n18826), .A3(n18825), .A4(n18824), .ZN(
        P2_U2830) );
  AOI22_X1 U20840 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18851), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n18850), .ZN(n18837) );
  AOI22_X1 U20841 ( .A1(n18828), .A2(n18853), .B1(P2_EBX_REG_26__SCAN_IN), 
        .B2(n18852), .ZN(n18836) );
  OAI22_X1 U20842 ( .A1(n18830), .A2(n18857), .B1(n18829), .B2(n18855), .ZN(
        n18831) );
  INV_X1 U20843 ( .A(n18831), .ZN(n18835) );
  OAI211_X1 U20844 ( .C1(n18833), .C2(n18832), .A(n18861), .B(n16602), .ZN(
        n18834) );
  NAND4_X1 U20845 ( .A1(n18837), .A2(n18836), .A3(n18835), .A4(n18834), .ZN(
        P2_U2829) );
  AOI22_X1 U20846 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18851), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n18850), .ZN(n18849) );
  AOI22_X1 U20847 ( .A1(n18838), .A2(n18853), .B1(P2_EBX_REG_28__SCAN_IN), 
        .B2(n18852), .ZN(n18848) );
  INV_X1 U20848 ( .A(n18839), .ZN(n18840) );
  OAI22_X1 U20849 ( .A1(n18841), .A2(n18857), .B1(n18840), .B2(n18855), .ZN(
        n18842) );
  INV_X1 U20850 ( .A(n18842), .ZN(n18847) );
  OAI211_X1 U20851 ( .C1(n18845), .C2(n18844), .A(n18861), .B(n18843), .ZN(
        n18846) );
  NAND4_X1 U20852 ( .A1(n18849), .A2(n18848), .A3(n18847), .A4(n18846), .ZN(
        P2_U2827) );
  AOI22_X1 U20853 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18851), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n18850), .ZN(n18867) );
  AOI22_X1 U20854 ( .A1(n18854), .A2(n18853), .B1(P2_EBX_REG_29__SCAN_IN), 
        .B2(n18852), .ZN(n18866) );
  OAI22_X1 U20855 ( .A1(n18858), .A2(n18857), .B1(n18856), .B2(n18855), .ZN(
        n18859) );
  INV_X1 U20856 ( .A(n18859), .ZN(n18865) );
  OAI211_X1 U20857 ( .C1(n18863), .C2(n18862), .A(n18861), .B(n18860), .ZN(
        n18864) );
  NAND4_X1 U20858 ( .A1(n18867), .A2(n18866), .A3(n18865), .A4(n18864), .ZN(
        P2_U2826) );
  INV_X1 U20859 ( .A(n18868), .ZN(n18874) );
  NOR4_X1 U20860 ( .A1(n18870), .A2(n18869), .A3(n11969), .A4(n18892), .ZN(
        n18871) );
  NAND2_X1 U20861 ( .A1(n18874), .A2(n18871), .ZN(n18872) );
  OAI21_X1 U20862 ( .B1(n18874), .B2(n18873), .A(n18872), .ZN(P2_U3595) );
  AOI22_X1 U20863 ( .A1(n18877), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n18876), .B2(n18875), .ZN(n18889) );
  NAND2_X1 U20864 ( .A1(n18879), .A2(n18878), .ZN(n18880) );
  OAI21_X1 U20865 ( .B1(n18882), .B2(n18881), .A(n18880), .ZN(n18887) );
  OAI21_X1 U20866 ( .B1(n18885), .B2(n18884), .A(n18883), .ZN(n18886) );
  NOR2_X1 U20867 ( .A1(n18887), .A2(n18886), .ZN(n18888) );
  OAI211_X1 U20868 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18890), .A(
        n18889), .B(n18888), .ZN(P2_U3046) );
  NAND2_X1 U20869 ( .A1(n18905), .A2(n18891), .ZN(n18907) );
  OAI21_X1 U20870 ( .B1(n18893), .B2(n18892), .A(n18914), .ZN(n18896) );
  NAND2_X1 U20871 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n21850), .ZN(n18894) );
  AOI21_X1 U20872 ( .B1(n18899), .B2(n18907), .A(n18894), .ZN(n18895) );
  AOI21_X1 U20873 ( .B1(n18907), .B2(n18896), .A(n18895), .ZN(n18898) );
  NAND2_X1 U20874 ( .A1(n18898), .A2(n18897), .ZN(P2_U3177) );
  OAI22_X1 U20875 ( .A1(n18901), .A2(n18900), .B1(n18908), .B2(n18899), .ZN(
        n18903) );
  OR2_X1 U20876 ( .A1(n18903), .A2(n18902), .ZN(n18904) );
  AOI21_X1 U20877 ( .B1(n18905), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n18904), 
        .ZN(n18912) );
  NOR2_X1 U20878 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n18906), .ZN(n18910) );
  OAI22_X1 U20879 ( .A1(n18910), .A2(n18909), .B1(n18908), .B2(n18907), .ZN(
        n18911) );
  OAI211_X1 U20880 ( .C1(n18913), .C2(n18914), .A(n18912), .B(n18911), .ZN(
        P2_U3176) );
  NOR2_X1 U20881 ( .A1(n18915), .A2(n18914), .ZN(n18919) );
  MUX2_X1 U20882 ( .A(P2_MORE_REG_SCAN_IN), .B(n18916), .S(n18919), .Z(
        P2_U3609) );
  INV_X1 U20883 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n18918) );
  OAI21_X1 U20884 ( .B1(n18919), .B2(n18918), .A(n18917), .ZN(P2_U2819) );
  INV_X1 U20885 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n20272) );
  INV_X1 U20886 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n20909) );
  AOI22_X1 U20887 ( .A1(n19257), .A2(n20272), .B1(n20909), .B2(U215), .ZN(U282) );
  INV_X1 U20888 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n18920) );
  INV_X1 U20889 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n20910) );
  AOI22_X1 U20890 ( .A1(n19257), .A2(n18920), .B1(n20910), .B2(U215), .ZN(U281) );
  INV_X1 U20891 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n18921) );
  INV_X1 U20892 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n20921) );
  AOI22_X1 U20893 ( .A1(n19257), .A2(n18921), .B1(n20921), .B2(U215), .ZN(U280) );
  OAI22_X1 U20894 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19257), .ZN(n18922) );
  INV_X1 U20895 ( .A(n18922), .ZN(U279) );
  INV_X1 U20896 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n18923) );
  INV_X1 U20897 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n20933) );
  AOI22_X1 U20898 ( .A1(n19257), .A2(n18923), .B1(n20933), .B2(U215), .ZN(U278) );
  OAI22_X1 U20899 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19257), .ZN(n18924) );
  INV_X1 U20900 ( .A(n18924), .ZN(U277) );
  OAI22_X1 U20901 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19095), .ZN(n18925) );
  INV_X1 U20902 ( .A(n18925), .ZN(U276) );
  OAI22_X1 U20903 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19095), .ZN(n18926) );
  INV_X1 U20904 ( .A(n18926), .ZN(U275) );
  OAI22_X1 U20905 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19095), .ZN(n18927) );
  INV_X1 U20906 ( .A(n18927), .ZN(U274) );
  OAI22_X1 U20907 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19095), .ZN(n18928) );
  INV_X1 U20908 ( .A(n18928), .ZN(U273) );
  OAI22_X1 U20909 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19095), .ZN(n18929) );
  INV_X1 U20910 ( .A(n18929), .ZN(U272) );
  INV_X1 U20911 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n18930) );
  AOI22_X1 U20912 ( .A1(n19095), .A2(n18930), .B1(n15956), .B2(U215), .ZN(U271) );
  OAI22_X1 U20913 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19095), .ZN(n18931) );
  INV_X1 U20914 ( .A(n18931), .ZN(U270) );
  OAI22_X1 U20915 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19257), .ZN(n18932) );
  INV_X1 U20916 ( .A(n18932), .ZN(U269) );
  OAI22_X1 U20917 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19257), .ZN(n18933) );
  INV_X1 U20918 ( .A(n18933), .ZN(U268) );
  OAI22_X1 U20919 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19257), .ZN(n18934) );
  INV_X1 U20920 ( .A(n18934), .ZN(U267) );
  OAI22_X1 U20921 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19257), .ZN(n18935) );
  INV_X1 U20922 ( .A(n18935), .ZN(U266) );
  OAI22_X1 U20923 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n19257), .ZN(n18936) );
  INV_X1 U20924 ( .A(n18936), .ZN(U265) );
  OAI22_X1 U20925 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n19257), .ZN(n18937) );
  INV_X1 U20926 ( .A(n18937), .ZN(U264) );
  INV_X1 U20927 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n18938) );
  INV_X1 U20928 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n20811) );
  AOI22_X1 U20929 ( .A1(n19257), .A2(n18938), .B1(n20811), .B2(U215), .ZN(U263) );
  INV_X1 U20930 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n18939) );
  INV_X1 U20931 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n20816) );
  AOI22_X1 U20932 ( .A1(n19257), .A2(n18939), .B1(n20816), .B2(U215), .ZN(U262) );
  OAI22_X1 U20933 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n19257), .ZN(n18940) );
  INV_X1 U20934 ( .A(n18940), .ZN(U261) );
  INV_X1 U20935 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n18941) );
  INV_X1 U20936 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n20900) );
  AOI22_X1 U20937 ( .A1(n19257), .A2(n18941), .B1(n20900), .B2(U215), .ZN(U260) );
  OAI22_X1 U20938 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n19257), .ZN(n18942) );
  INV_X1 U20939 ( .A(n18942), .ZN(U259) );
  INV_X1 U20940 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n18943) );
  INV_X1 U20941 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n20826) );
  AOI22_X1 U20942 ( .A1(n19257), .A2(n18943), .B1(n20826), .B2(U215), .ZN(U258) );
  NOR2_X1 U20943 ( .A1(n21465), .A2(n18944), .ZN(n19003) );
  NAND2_X1 U20944 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19003), .ZN(
        n19203) );
  NAND2_X1 U20945 ( .A1(n19016), .A2(n20801), .ZN(n19014) );
  NOR2_X1 U20946 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18945), .ZN(
        n18950) );
  NAND2_X1 U20947 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18950), .ZN(
        n19266) );
  INV_X1 U20948 ( .A(n19266), .ZN(n19353) );
  AND2_X1 U20949 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19215), .ZN(n19007) );
  AND2_X1 U20950 ( .A1(n21479), .A2(n19003), .ZN(n19260) );
  NOR2_X2 U20951 ( .A1(n20826), .A2(n19173), .ZN(n19006) );
  AOI22_X1 U20952 ( .A1(n19353), .A2(n19007), .B1(n19260), .B2(n19006), .ZN(
        n18947) );
  AOI22_X1 U20953 ( .A1(n19215), .A2(n18950), .B1(n18958), .B2(n19003), .ZN(
        n19263) );
  NAND2_X1 U20954 ( .A1(n21449), .A2(n18950), .ZN(n19219) );
  INV_X1 U20955 ( .A(n19219), .ZN(n19279) );
  NOR2_X2 U20956 ( .A1(n20909), .A2(n19054), .ZN(n19011) );
  AOI22_X1 U20957 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19263), .B1(
        n19279), .B2(n19011), .ZN(n18946) );
  OAI211_X1 U20958 ( .C1(n19203), .C2(n19014), .A(n18947), .B(n18946), .ZN(
        P3_U2995) );
  NAND2_X1 U20959 ( .A1(n19003), .A2(n21449), .ZN(n19360) );
  NAND2_X1 U20960 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18959), .ZN(
        n18956) );
  NOR2_X2 U20961 ( .A1(n21449), .A2(n18956), .ZN(n19285) );
  NAND2_X1 U20962 ( .A1(n19266), .A2(n19360), .ZN(n19010) );
  AND2_X1 U20963 ( .A1(n21479), .A2(n19010), .ZN(n19267) );
  AOI22_X1 U20964 ( .A1(n19011), .A2(n19285), .B1(n19006), .B2(n19267), .ZN(
        n18949) );
  INV_X1 U20965 ( .A(n19285), .ZN(n19272) );
  NAND2_X1 U20966 ( .A1(n19219), .A2(n19272), .ZN(n18953) );
  AOI21_X1 U20967 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n19173), .ZN(n19009) );
  OAI221_X1 U20968 ( .B1(n19010), .B2(n18979), .C1(n19010), .C2(n18953), .A(
        n19009), .ZN(n19269) );
  AOI22_X1 U20969 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19269), .B1(
        n19279), .B2(n19007), .ZN(n18948) );
  OAI211_X1 U20970 ( .C1(n19014), .C2(n19360), .A(n18949), .B(n18948), .ZN(
        P3_U2987) );
  NOR2_X2 U20971 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18956), .ZN(
        n19290) );
  AND2_X1 U20972 ( .A1(n21479), .A2(n18950), .ZN(n19273) );
  AOI22_X1 U20973 ( .A1(n19011), .A2(n19290), .B1(n19006), .B2(n19273), .ZN(
        n18952) );
  INV_X1 U20974 ( .A(n18956), .ZN(n18957) );
  AOI22_X1 U20975 ( .A1(n19215), .A2(n18957), .B1(n18958), .B2(n18950), .ZN(
        n19274) );
  AOI22_X1 U20976 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19274), .B1(
        n19007), .B2(n19285), .ZN(n18951) );
  OAI211_X1 U20977 ( .C1(n19014), .C2(n19266), .A(n18952), .B(n18951), .ZN(
        P3_U2979) );
  INV_X1 U20978 ( .A(n19283), .ZN(n19296) );
  AND2_X1 U20979 ( .A1(n21479), .A2(n18953), .ZN(n19278) );
  AOI22_X1 U20980 ( .A1(n19296), .A2(n19011), .B1(n19006), .B2(n19278), .ZN(
        n18955) );
  INV_X1 U20981 ( .A(n19290), .ZN(n19277) );
  NAND2_X1 U20982 ( .A1(n19283), .A2(n19277), .ZN(n18963) );
  AOI22_X1 U20983 ( .A1(n19215), .A2(n18963), .B1(n19009), .B2(n18953), .ZN(
        n19280) );
  AOI22_X1 U20984 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19280), .B1(
        n19007), .B2(n19290), .ZN(n18954) );
  OAI211_X1 U20985 ( .C1(n19219), .C2(n19014), .A(n18955), .B(n18954), .ZN(
        P3_U2971) );
  NOR2_X1 U20986 ( .A1(n20338), .A2(n18956), .ZN(n19284) );
  AOI22_X1 U20987 ( .A1(n19296), .A2(n19007), .B1(n19006), .B2(n19284), .ZN(
        n18961) );
  AOI22_X1 U20988 ( .A1(n19215), .A2(n18959), .B1(n18958), .B2(n18957), .ZN(
        n19286) );
  NOR2_X1 U20989 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21454) );
  NAND2_X1 U20990 ( .A1(n21454), .A2(n18959), .ZN(n19294) );
  INV_X1 U20991 ( .A(n19294), .ZN(n19302) );
  AOI22_X1 U20992 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19286), .B1(
        n19011), .B2(n19302), .ZN(n18960) );
  OAI211_X1 U20993 ( .C1(n19014), .C2(n19272), .A(n18961), .B(n18960), .ZN(
        P3_U2963) );
  AND2_X1 U20994 ( .A1(n21479), .A2(n18963), .ZN(n19289) );
  AOI22_X1 U20995 ( .A1(n19007), .A2(n19302), .B1(n19006), .B2(n19289), .ZN(
        n18965) );
  NAND2_X1 U20996 ( .A1(n19300), .A2(n19294), .ZN(n18969) );
  AOI21_X1 U20997 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19277), .A(n19173), 
        .ZN(n18962) );
  OAI221_X1 U20998 ( .B1(n18963), .B2(n18979), .C1(n18963), .C2(n18969), .A(
        n18962), .ZN(n19291) );
  AOI22_X1 U20999 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19291), .B1(
        n19308), .B2(n19011), .ZN(n18964) );
  OAI211_X1 U21000 ( .C1(n19014), .C2(n19277), .A(n18965), .B(n18964), .ZN(
        P3_U2955) );
  INV_X1 U21001 ( .A(n19306), .ZN(n19314) );
  AOI22_X1 U21002 ( .A1(n19314), .A2(n19011), .B1(n19295), .B2(n19006), .ZN(
        n18967) );
  AOI22_X1 U21003 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19297), .B1(
        n19308), .B2(n19007), .ZN(n18966) );
  OAI211_X1 U21004 ( .C1(n19283), .C2(n19014), .A(n18967), .B(n18966), .ZN(
        P3_U2947) );
  AND2_X1 U21005 ( .A1(n21479), .A2(n18969), .ZN(n19301) );
  AOI22_X1 U21006 ( .A1(n19314), .A2(n19007), .B1(n19006), .B2(n19301), .ZN(
        n18971) );
  NOR2_X1 U21007 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18968), .ZN(
        n18983) );
  NAND2_X1 U21008 ( .A1(n18987), .A2(n18983), .ZN(n19312) );
  NAND2_X1 U21009 ( .A1(n19306), .A2(n19312), .ZN(n18978) );
  AOI22_X1 U21010 ( .A1(n19215), .A2(n18978), .B1(n19009), .B2(n18969), .ZN(
        n19303) );
  INV_X1 U21011 ( .A(n19312), .ZN(n19320) );
  AOI22_X1 U21012 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19303), .B1(
        n19011), .B2(n19320), .ZN(n18970) );
  OAI211_X1 U21013 ( .C1(n19014), .C2(n19294), .A(n18971), .B(n18970), .ZN(
        P3_U2939) );
  NAND2_X1 U21014 ( .A1(n21454), .A2(n18983), .ZN(n19318) );
  INV_X1 U21015 ( .A(n19318), .ZN(n19326) );
  INV_X1 U21016 ( .A(n18972), .ZN(n18973) );
  NOR2_X1 U21017 ( .A1(n20338), .A2(n18973), .ZN(n19307) );
  AOI22_X1 U21018 ( .A1(n19011), .A2(n19326), .B1(n19006), .B2(n19307), .ZN(
        n18976) );
  OAI21_X1 U21019 ( .B1(n19173), .B2(n21450), .A(n19054), .ZN(n18993) );
  NAND3_X1 U21020 ( .A1(n18983), .A2(n18974), .A3(n18993), .ZN(n19309) );
  AOI22_X1 U21021 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19309), .B1(
        n19007), .B2(n19320), .ZN(n18975) );
  OAI211_X1 U21022 ( .C1(n19300), .C2(n19014), .A(n18976), .B(n18975), .ZN(
        P3_U2931) );
  AND2_X1 U21023 ( .A1(n21479), .A2(n18978), .ZN(n19313) );
  AOI22_X1 U21024 ( .A1(n19007), .A2(n19326), .B1(n19006), .B2(n19313), .ZN(
        n18981) );
  NOR2_X1 U21025 ( .A1(n21450), .A2(n18999), .ZN(n18984) );
  NAND2_X1 U21026 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18984), .ZN(
        n19240) );
  INV_X1 U21027 ( .A(n19240), .ZN(n19331) );
  OAI21_X1 U21028 ( .B1(n19326), .B2(n19331), .A(n19009), .ZN(n18977) );
  INV_X1 U21029 ( .A(n18977), .ZN(n18989) );
  AOI22_X1 U21030 ( .A1(n18979), .A2(n18989), .B1(n19009), .B2(n18978), .ZN(
        n19315) );
  AOI22_X1 U21031 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19315), .B1(
        n19011), .B2(n19331), .ZN(n18980) );
  OAI211_X1 U21032 ( .C1(n19306), .C2(n19014), .A(n18981), .B(n18980), .ZN(
        P3_U2923) );
  INV_X1 U21033 ( .A(n18984), .ZN(n18992) );
  NOR2_X2 U21034 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18992), .ZN(
        n19337) );
  INV_X1 U21035 ( .A(n18983), .ZN(n18982) );
  NOR2_X1 U21036 ( .A1(n19000), .A2(n18982), .ZN(n19319) );
  AOI22_X1 U21037 ( .A1(n19011), .A2(n19337), .B1(n19006), .B2(n19319), .ZN(
        n18986) );
  AOI22_X1 U21038 ( .A1(n19215), .A2(n18984), .B1(n19002), .B2(n18983), .ZN(
        n19321) );
  AOI22_X1 U21039 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19321), .B1(
        n19007), .B2(n19331), .ZN(n18985) );
  OAI211_X1 U21040 ( .C1(n19014), .C2(n19312), .A(n18986), .B(n18985), .ZN(
        P3_U2915) );
  INV_X1 U21041 ( .A(n18987), .ZN(n18988) );
  NOR2_X2 U21042 ( .A1(n18988), .A2(n18999), .ZN(n19345) );
  AOI21_X1 U21043 ( .B1(n19318), .B2(n19240), .A(n20338), .ZN(n19325) );
  AOI22_X1 U21044 ( .A1(n19011), .A2(n19345), .B1(n19006), .B2(n19325), .ZN(
        n18991) );
  INV_X1 U21045 ( .A(n19337), .ZN(n19324) );
  INV_X1 U21046 ( .A(n19345), .ZN(n19335) );
  NAND2_X1 U21047 ( .A1(n19324), .A2(n19335), .ZN(n18996) );
  AOI21_X1 U21048 ( .B1(n19215), .B2(n18996), .A(n18989), .ZN(n19327) );
  AOI22_X1 U21049 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19327), .B1(
        n19007), .B2(n19337), .ZN(n18990) );
  OAI211_X1 U21050 ( .C1(n19014), .C2(n19318), .A(n18991), .B(n18990), .ZN(
        P3_U2907) );
  INV_X1 U21051 ( .A(n18999), .ZN(n19001) );
  NAND2_X1 U21052 ( .A1(n21454), .A2(n19001), .ZN(n19341) );
  INV_X1 U21053 ( .A(n19341), .ZN(n19355) );
  NOR2_X1 U21054 ( .A1(n20338), .A2(n18992), .ZN(n19330) );
  AOI22_X1 U21055 ( .A1(n19011), .A2(n19355), .B1(n19006), .B2(n19330), .ZN(
        n18995) );
  OAI211_X1 U21056 ( .C1(n19331), .C2(n21488), .A(n19001), .B(n18993), .ZN(
        n19332) );
  AOI22_X1 U21057 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19332), .B1(
        n19007), .B2(n19345), .ZN(n18994) );
  OAI211_X1 U21058 ( .C1(n19014), .C2(n19240), .A(n18995), .B(n18994), .ZN(
        P3_U2899) );
  INV_X1 U21059 ( .A(n19203), .ZN(n19344) );
  AND2_X1 U21060 ( .A1(n21479), .A2(n18996), .ZN(n19336) );
  AOI22_X1 U21061 ( .A1(n19011), .A2(n19344), .B1(n19006), .B2(n19336), .ZN(
        n18998) );
  NAND2_X1 U21062 ( .A1(n19203), .A2(n19341), .ZN(n19008) );
  AOI22_X1 U21063 ( .A1(n19215), .A2(n19008), .B1(n19009), .B2(n18996), .ZN(
        n19338) );
  AOI22_X1 U21064 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19338), .B1(
        n19007), .B2(n19355), .ZN(n18997) );
  OAI211_X1 U21065 ( .C1(n19014), .C2(n19324), .A(n18998), .B(n18997), .ZN(
        P3_U2891) );
  NOR2_X1 U21066 ( .A1(n19000), .A2(n18999), .ZN(n19342) );
  AOI22_X1 U21067 ( .A1(n19344), .A2(n19007), .B1(n19006), .B2(n19342), .ZN(
        n19005) );
  AOI22_X1 U21068 ( .A1(n19215), .A2(n19003), .B1(n19002), .B2(n19001), .ZN(
        n19346) );
  INV_X1 U21069 ( .A(n19360), .ZN(n19268) );
  AOI22_X1 U21070 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19346), .B1(
        n19011), .B2(n19268), .ZN(n19004) );
  OAI211_X1 U21071 ( .C1(n19014), .C2(n19335), .A(n19005), .B(n19004), .ZN(
        P3_U2883) );
  AND2_X1 U21072 ( .A1(n21479), .A2(n19008), .ZN(n19351) );
  AOI22_X1 U21073 ( .A1(n19007), .A2(n19268), .B1(n19006), .B2(n19351), .ZN(
        n19013) );
  AOI22_X1 U21074 ( .A1(n19215), .A2(n19010), .B1(n19009), .B2(n19008), .ZN(
        n19356) );
  AOI22_X1 U21075 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19356), .B1(
        n19011), .B2(n19353), .ZN(n19012) );
  OAI211_X1 U21076 ( .C1(n19014), .C2(n19341), .A(n19013), .B(n19012), .ZN(
        P3_U2875) );
  INV_X1 U21077 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n19015) );
  INV_X1 U21078 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n20878) );
  AOI22_X1 U21079 ( .A1(n19095), .A2(n19015), .B1(n20878), .B2(U215), .ZN(U257) );
  NAND2_X1 U21080 ( .A1(n19016), .A2(n20856), .ZN(n19052) );
  AND2_X1 U21081 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n19215), .ZN(n19049) );
  NOR2_X2 U21082 ( .A1(n20878), .A2(n19173), .ZN(n19047) );
  AOI22_X1 U21083 ( .A1(n19353), .A2(n19049), .B1(n19260), .B2(n19047), .ZN(
        n19018) );
  NOR2_X2 U21084 ( .A1(n20910), .A2(n19054), .ZN(n19048) );
  AOI22_X1 U21085 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19263), .B1(
        n19279), .B2(n19048), .ZN(n19017) );
  OAI211_X1 U21086 ( .C1(n19203), .C2(n19052), .A(n19018), .B(n19017), .ZN(
        P3_U2994) );
  AOI22_X1 U21087 ( .A1(n19285), .A2(n19048), .B1(n19267), .B2(n19047), .ZN(
        n19020) );
  AOI22_X1 U21088 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19269), .B1(
        n19279), .B2(n19049), .ZN(n19019) );
  OAI211_X1 U21089 ( .C1(n19360), .C2(n19052), .A(n19020), .B(n19019), .ZN(
        P3_U2986) );
  AOI22_X1 U21090 ( .A1(n19285), .A2(n19049), .B1(n19273), .B2(n19047), .ZN(
        n19022) );
  AOI22_X1 U21091 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19274), .B1(
        n19290), .B2(n19048), .ZN(n19021) );
  OAI211_X1 U21092 ( .C1(n19266), .C2(n19052), .A(n19022), .B(n19021), .ZN(
        P3_U2978) );
  AOI22_X1 U21093 ( .A1(n19290), .A2(n19049), .B1(n19278), .B2(n19047), .ZN(
        n19024) );
  AOI22_X1 U21094 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19280), .B1(
        n19296), .B2(n19048), .ZN(n19023) );
  OAI211_X1 U21095 ( .C1(n19219), .C2(n19052), .A(n19024), .B(n19023), .ZN(
        P3_U2970) );
  AOI22_X1 U21096 ( .A1(n19302), .A2(n19048), .B1(n19284), .B2(n19047), .ZN(
        n19026) );
  AOI22_X1 U21097 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19286), .B1(
        n19296), .B2(n19049), .ZN(n19025) );
  OAI211_X1 U21098 ( .C1(n19272), .C2(n19052), .A(n19026), .B(n19025), .ZN(
        P3_U2962) );
  AOI22_X1 U21099 ( .A1(n19302), .A2(n19049), .B1(n19289), .B2(n19047), .ZN(
        n19028) );
  AOI22_X1 U21100 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19291), .B1(
        n19308), .B2(n19048), .ZN(n19027) );
  OAI211_X1 U21101 ( .C1(n19277), .C2(n19052), .A(n19028), .B(n19027), .ZN(
        P3_U2954) );
  AOI22_X1 U21102 ( .A1(n19314), .A2(n19048), .B1(n19295), .B2(n19047), .ZN(
        n19030) );
  AOI22_X1 U21103 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19297), .B1(
        n19308), .B2(n19049), .ZN(n19029) );
  OAI211_X1 U21104 ( .C1(n19283), .C2(n19052), .A(n19030), .B(n19029), .ZN(
        P3_U2946) );
  AOI22_X1 U21105 ( .A1(n19320), .A2(n19048), .B1(n19301), .B2(n19047), .ZN(
        n19032) );
  AOI22_X1 U21106 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19303), .B1(
        n19314), .B2(n19049), .ZN(n19031) );
  OAI211_X1 U21107 ( .C1(n19294), .C2(n19052), .A(n19032), .B(n19031), .ZN(
        P3_U2938) );
  AOI22_X1 U21108 ( .A1(n19326), .A2(n19048), .B1(n19307), .B2(n19047), .ZN(
        n19034) );
  AOI22_X1 U21109 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19309), .B1(
        n19320), .B2(n19049), .ZN(n19033) );
  OAI211_X1 U21110 ( .C1(n19300), .C2(n19052), .A(n19034), .B(n19033), .ZN(
        P3_U2930) );
  AOI22_X1 U21111 ( .A1(n19326), .A2(n19049), .B1(n19313), .B2(n19047), .ZN(
        n19036) );
  AOI22_X1 U21112 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19315), .B1(
        n19331), .B2(n19048), .ZN(n19035) );
  OAI211_X1 U21113 ( .C1(n19306), .C2(n19052), .A(n19036), .B(n19035), .ZN(
        P3_U2922) );
  AOI22_X1 U21114 ( .A1(n19331), .A2(n19049), .B1(n19319), .B2(n19047), .ZN(
        n19038) );
  AOI22_X1 U21115 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19321), .B1(
        n19337), .B2(n19048), .ZN(n19037) );
  OAI211_X1 U21116 ( .C1(n19312), .C2(n19052), .A(n19038), .B(n19037), .ZN(
        P3_U2914) );
  AOI22_X1 U21117 ( .A1(n19337), .A2(n19049), .B1(n19325), .B2(n19047), .ZN(
        n19040) );
  AOI22_X1 U21118 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19327), .B1(
        n19345), .B2(n19048), .ZN(n19039) );
  OAI211_X1 U21119 ( .C1(n19318), .C2(n19052), .A(n19040), .B(n19039), .ZN(
        P3_U2906) );
  AOI22_X1 U21120 ( .A1(n19330), .A2(n19047), .B1(n19355), .B2(n19048), .ZN(
        n19042) );
  AOI22_X1 U21121 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19332), .B1(
        n19345), .B2(n19049), .ZN(n19041) );
  OAI211_X1 U21122 ( .C1(n19240), .C2(n19052), .A(n19042), .B(n19041), .ZN(
        P3_U2898) );
  AOI22_X1 U21123 ( .A1(n19344), .A2(n19048), .B1(n19336), .B2(n19047), .ZN(
        n19044) );
  AOI22_X1 U21124 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19338), .B1(
        n19355), .B2(n19049), .ZN(n19043) );
  OAI211_X1 U21125 ( .C1(n19324), .C2(n19052), .A(n19044), .B(n19043), .ZN(
        P3_U2890) );
  AOI22_X1 U21126 ( .A1(n19344), .A2(n19049), .B1(n19342), .B2(n19047), .ZN(
        n19046) );
  AOI22_X1 U21127 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19346), .B1(
        n19268), .B2(n19048), .ZN(n19045) );
  OAI211_X1 U21128 ( .C1(n19335), .C2(n19052), .A(n19046), .B(n19045), .ZN(
        P3_U2882) );
  AOI22_X1 U21129 ( .A1(n19353), .A2(n19048), .B1(n19351), .B2(n19047), .ZN(
        n19051) );
  AOI22_X1 U21130 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19356), .B1(
        n19268), .B2(n19049), .ZN(n19050) );
  OAI211_X1 U21131 ( .C1(n19341), .C2(n19052), .A(n19051), .B(n19050), .ZN(
        P3_U2874) );
  INV_X1 U21132 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n19053) );
  INV_X1 U21133 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n20839) );
  AOI22_X1 U21134 ( .A1(n19095), .A2(n19053), .B1(n20839), .B2(U215), .ZN(U256) );
  NAND2_X1 U21135 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n19215), .ZN(n19083) );
  NOR2_X1 U21136 ( .A1(n20921), .A2(n19054), .ZN(n19080) );
  NOR2_X2 U21137 ( .A1(n20839), .A2(n19173), .ZN(n19088) );
  AOI22_X1 U21138 ( .A1(n19279), .A2(n19080), .B1(n19260), .B2(n19088), .ZN(
        n19057) );
  NOR2_X2 U21139 ( .A1(n19055), .A2(n19261), .ZN(n19090) );
  AOI22_X1 U21140 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19263), .B1(
        n19344), .B2(n19090), .ZN(n19056) );
  OAI211_X1 U21141 ( .C1(n19266), .C2(n19083), .A(n19057), .B(n19056), .ZN(
        P3_U2993) );
  AOI22_X1 U21142 ( .A1(n19285), .A2(n19080), .B1(n19267), .B2(n19088), .ZN(
        n19059) );
  AOI22_X1 U21143 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19269), .B1(
        n19268), .B2(n19090), .ZN(n19058) );
  OAI211_X1 U21144 ( .C1(n19219), .C2(n19083), .A(n19059), .B(n19058), .ZN(
        P3_U2985) );
  INV_X1 U21145 ( .A(n19080), .ZN(n19093) );
  INV_X1 U21146 ( .A(n19083), .ZN(n19089) );
  AOI22_X1 U21147 ( .A1(n19285), .A2(n19089), .B1(n19273), .B2(n19088), .ZN(
        n19061) );
  AOI22_X1 U21148 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19274), .B1(
        n19353), .B2(n19090), .ZN(n19060) );
  OAI211_X1 U21149 ( .C1(n19277), .C2(n19093), .A(n19061), .B(n19060), .ZN(
        P3_U2977) );
  AOI22_X1 U21150 ( .A1(n19290), .A2(n19089), .B1(n19278), .B2(n19088), .ZN(
        n19063) );
  AOI22_X1 U21151 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19280), .B1(
        n19279), .B2(n19090), .ZN(n19062) );
  OAI211_X1 U21152 ( .C1(n19283), .C2(n19093), .A(n19063), .B(n19062), .ZN(
        P3_U2969) );
  AOI22_X1 U21153 ( .A1(n19296), .A2(n19089), .B1(n19284), .B2(n19088), .ZN(
        n19065) );
  AOI22_X1 U21154 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19286), .B1(
        n19285), .B2(n19090), .ZN(n19064) );
  OAI211_X1 U21155 ( .C1(n19294), .C2(n19093), .A(n19065), .B(n19064), .ZN(
        P3_U2961) );
  AOI22_X1 U21156 ( .A1(n19302), .A2(n19089), .B1(n19289), .B2(n19088), .ZN(
        n19067) );
  AOI22_X1 U21157 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19291), .B1(
        n19290), .B2(n19090), .ZN(n19066) );
  OAI211_X1 U21158 ( .C1(n19300), .C2(n19093), .A(n19067), .B(n19066), .ZN(
        P3_U2953) );
  AOI22_X1 U21159 ( .A1(n19314), .A2(n19080), .B1(n19295), .B2(n19088), .ZN(
        n19069) );
  AOI22_X1 U21160 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19297), .B1(
        n19296), .B2(n19090), .ZN(n19068) );
  OAI211_X1 U21161 ( .C1(n19300), .C2(n19083), .A(n19069), .B(n19068), .ZN(
        P3_U2945) );
  AOI22_X1 U21162 ( .A1(n19314), .A2(n19089), .B1(n19301), .B2(n19088), .ZN(
        n19071) );
  AOI22_X1 U21163 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19303), .B1(
        n19302), .B2(n19090), .ZN(n19070) );
  OAI211_X1 U21164 ( .C1(n19312), .C2(n19093), .A(n19071), .B(n19070), .ZN(
        P3_U2937) );
  AOI22_X1 U21165 ( .A1(n19320), .A2(n19089), .B1(n19307), .B2(n19088), .ZN(
        n19073) );
  AOI22_X1 U21166 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19309), .B1(
        n19308), .B2(n19090), .ZN(n19072) );
  OAI211_X1 U21167 ( .C1(n19318), .C2(n19093), .A(n19073), .B(n19072), .ZN(
        P3_U2929) );
  AOI22_X1 U21168 ( .A1(n19331), .A2(n19080), .B1(n19313), .B2(n19088), .ZN(
        n19075) );
  AOI22_X1 U21169 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19315), .B1(
        n19314), .B2(n19090), .ZN(n19074) );
  OAI211_X1 U21170 ( .C1(n19318), .C2(n19083), .A(n19075), .B(n19074), .ZN(
        P3_U2921) );
  AOI22_X1 U21171 ( .A1(n19331), .A2(n19089), .B1(n19319), .B2(n19088), .ZN(
        n19077) );
  AOI22_X1 U21172 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19321), .B1(
        n19320), .B2(n19090), .ZN(n19076) );
  OAI211_X1 U21173 ( .C1(n19324), .C2(n19093), .A(n19077), .B(n19076), .ZN(
        P3_U2913) );
  AOI22_X1 U21174 ( .A1(n19337), .A2(n19089), .B1(n19325), .B2(n19088), .ZN(
        n19079) );
  AOI22_X1 U21175 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19327), .B1(
        n19326), .B2(n19090), .ZN(n19078) );
  OAI211_X1 U21176 ( .C1(n19335), .C2(n19093), .A(n19079), .B(n19078), .ZN(
        P3_U2905) );
  AOI22_X1 U21177 ( .A1(n19330), .A2(n19088), .B1(n19355), .B2(n19080), .ZN(
        n19082) );
  AOI22_X1 U21178 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19332), .B1(
        n19331), .B2(n19090), .ZN(n19081) );
  OAI211_X1 U21179 ( .C1(n19335), .C2(n19083), .A(n19082), .B(n19081), .ZN(
        P3_U2897) );
  AOI22_X1 U21180 ( .A1(n19355), .A2(n19089), .B1(n19336), .B2(n19088), .ZN(
        n19085) );
  AOI22_X1 U21181 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19338), .B1(
        n19337), .B2(n19090), .ZN(n19084) );
  OAI211_X1 U21182 ( .C1(n19203), .C2(n19093), .A(n19085), .B(n19084), .ZN(
        P3_U2889) );
  AOI22_X1 U21183 ( .A1(n19344), .A2(n19089), .B1(n19342), .B2(n19088), .ZN(
        n19087) );
  AOI22_X1 U21184 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19346), .B1(
        n19345), .B2(n19090), .ZN(n19086) );
  OAI211_X1 U21185 ( .C1(n19360), .C2(n19093), .A(n19087), .B(n19086), .ZN(
        P3_U2881) );
  AOI22_X1 U21186 ( .A1(n19268), .A2(n19089), .B1(n19351), .B2(n19088), .ZN(
        n19092) );
  AOI22_X1 U21187 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19356), .B1(
        n19355), .B2(n19090), .ZN(n19091) );
  OAI211_X1 U21188 ( .C1(n19266), .C2(n19093), .A(n19092), .B(n19091), .ZN(
        P3_U2873) );
  INV_X1 U21189 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n19094) );
  AOI22_X1 U21190 ( .A1(n19095), .A2(n19094), .B1(n20843), .B2(U215), .ZN(U255) );
  INV_X1 U21191 ( .A(n19131), .ZN(n19120) );
  AOI22_X1 U21192 ( .A1(n19120), .A2(n19279), .B1(n19126), .B2(n19260), .ZN(
        n19097) );
  AOI22_X1 U21193 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19263), .B1(
        n19128), .B2(n19344), .ZN(n19096) );
  OAI211_X1 U21194 ( .C1(n19123), .C2(n19266), .A(n19097), .B(n19096), .ZN(
        P3_U2992) );
  AOI22_X1 U21195 ( .A1(n19127), .A2(n19279), .B1(n19126), .B2(n19267), .ZN(
        n19099) );
  AOI22_X1 U21196 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19269), .B1(
        n19128), .B2(n19268), .ZN(n19098) );
  OAI211_X1 U21197 ( .C1(n19131), .C2(n19272), .A(n19099), .B(n19098), .ZN(
        P3_U2984) );
  AOI22_X1 U21198 ( .A1(n19127), .A2(n19285), .B1(n19126), .B2(n19273), .ZN(
        n19101) );
  AOI22_X1 U21199 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19274), .B1(
        n19128), .B2(n19353), .ZN(n19100) );
  OAI211_X1 U21200 ( .C1(n19131), .C2(n19277), .A(n19101), .B(n19100), .ZN(
        P3_U2976) );
  AOI22_X1 U21201 ( .A1(n19127), .A2(n19290), .B1(n19126), .B2(n19278), .ZN(
        n19103) );
  AOI22_X1 U21202 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19280), .B1(
        n19128), .B2(n19279), .ZN(n19102) );
  OAI211_X1 U21203 ( .C1(n19131), .C2(n19283), .A(n19103), .B(n19102), .ZN(
        P3_U2968) );
  AOI22_X1 U21204 ( .A1(n19120), .A2(n19302), .B1(n19126), .B2(n19284), .ZN(
        n19105) );
  AOI22_X1 U21205 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19286), .B1(
        n19128), .B2(n19285), .ZN(n19104) );
  OAI211_X1 U21206 ( .C1(n19283), .C2(n19123), .A(n19105), .B(n19104), .ZN(
        P3_U2960) );
  AOI22_X1 U21207 ( .A1(n19127), .A2(n19302), .B1(n19126), .B2(n19289), .ZN(
        n19107) );
  AOI22_X1 U21208 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19291), .B1(
        n19128), .B2(n19290), .ZN(n19106) );
  OAI211_X1 U21209 ( .C1(n19131), .C2(n19300), .A(n19107), .B(n19106), .ZN(
        P3_U2952) );
  AOI22_X1 U21210 ( .A1(n19120), .A2(n19320), .B1(n19126), .B2(n19301), .ZN(
        n19109) );
  AOI22_X1 U21211 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19303), .B1(
        n19128), .B2(n19302), .ZN(n19108) );
  OAI211_X1 U21212 ( .C1(n19306), .C2(n19123), .A(n19109), .B(n19108), .ZN(
        P3_U2936) );
  AOI22_X1 U21213 ( .A1(n19120), .A2(n19326), .B1(n19126), .B2(n19307), .ZN(
        n19111) );
  AOI22_X1 U21214 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19309), .B1(
        n19128), .B2(n19308), .ZN(n19110) );
  OAI211_X1 U21215 ( .C1(n19123), .C2(n19312), .A(n19111), .B(n19110), .ZN(
        P3_U2928) );
  AOI22_X1 U21216 ( .A1(n19120), .A2(n19331), .B1(n19126), .B2(n19313), .ZN(
        n19113) );
  AOI22_X1 U21217 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19315), .B1(
        n19314), .B2(n19128), .ZN(n19112) );
  OAI211_X1 U21218 ( .C1(n19123), .C2(n19318), .A(n19113), .B(n19112), .ZN(
        P3_U2920) );
  AOI22_X1 U21219 ( .A1(n19127), .A2(n19331), .B1(n19126), .B2(n19319), .ZN(
        n19115) );
  AOI22_X1 U21220 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19321), .B1(
        n19128), .B2(n19320), .ZN(n19114) );
  OAI211_X1 U21221 ( .C1(n19131), .C2(n19324), .A(n19115), .B(n19114), .ZN(
        P3_U2912) );
  AOI22_X1 U21222 ( .A1(n19127), .A2(n19337), .B1(n19126), .B2(n19325), .ZN(
        n19117) );
  AOI22_X1 U21223 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19327), .B1(
        n19128), .B2(n19326), .ZN(n19116) );
  OAI211_X1 U21224 ( .C1(n19131), .C2(n19335), .A(n19117), .B(n19116), .ZN(
        P3_U2904) );
  AOI22_X1 U21225 ( .A1(n19127), .A2(n19345), .B1(n19126), .B2(n19330), .ZN(
        n19119) );
  AOI22_X1 U21226 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19332), .B1(
        n19128), .B2(n19331), .ZN(n19118) );
  OAI211_X1 U21227 ( .C1(n19131), .C2(n19341), .A(n19119), .B(n19118), .ZN(
        P3_U2896) );
  AOI22_X1 U21228 ( .A1(n19120), .A2(n19344), .B1(n19126), .B2(n19336), .ZN(
        n19122) );
  AOI22_X1 U21229 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19338), .B1(
        n19128), .B2(n19337), .ZN(n19121) );
  OAI211_X1 U21230 ( .C1(n19123), .C2(n19341), .A(n19122), .B(n19121), .ZN(
        P3_U2888) );
  AOI22_X1 U21231 ( .A1(n19127), .A2(n19344), .B1(n19126), .B2(n19342), .ZN(
        n19125) );
  AOI22_X1 U21232 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19346), .B1(
        n19128), .B2(n19345), .ZN(n19124) );
  OAI211_X1 U21233 ( .C1(n19131), .C2(n19360), .A(n19125), .B(n19124), .ZN(
        P3_U2880) );
  AOI22_X1 U21234 ( .A1(n19127), .A2(n19268), .B1(n19126), .B2(n19351), .ZN(
        n19130) );
  AOI22_X1 U21235 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19356), .B1(
        n19128), .B2(n19355), .ZN(n19129) );
  OAI211_X1 U21236 ( .C1(n19131), .C2(n19266), .A(n19130), .B(n19129), .ZN(
        P3_U2872) );
  INV_X1 U21237 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n19132) );
  INV_X1 U21238 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n20848) );
  AOI22_X1 U21239 ( .A1(n19257), .A2(n19132), .B1(n20848), .B2(U215), .ZN(U254) );
  NAND2_X1 U21240 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19215), .ZN(n19155) );
  NAND2_X1 U21241 ( .A1(BUF2_REG_19__SCAN_IN), .A2(n19215), .ZN(n19171) );
  INV_X1 U21242 ( .A(n19171), .ZN(n19152) );
  NOR2_X2 U21243 ( .A1(n20848), .A2(n19173), .ZN(n19166) );
  AOI22_X1 U21244 ( .A1(n19353), .A2(n19152), .B1(n19260), .B2(n19166), .ZN(
        n19135) );
  NOR2_X2 U21245 ( .A1(n19133), .A2(n19261), .ZN(n19168) );
  AOI22_X1 U21246 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19263), .B1(
        n19344), .B2(n19168), .ZN(n19134) );
  OAI211_X1 U21247 ( .C1(n19219), .C2(n19155), .A(n19135), .B(n19134), .ZN(
        P3_U2991) );
  AOI22_X1 U21248 ( .A1(n19279), .A2(n19152), .B1(n19267), .B2(n19166), .ZN(
        n19137) );
  AOI22_X1 U21249 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19269), .B1(
        n19268), .B2(n19168), .ZN(n19136) );
  OAI211_X1 U21250 ( .C1(n19272), .C2(n19155), .A(n19137), .B(n19136), .ZN(
        P3_U2983) );
  AOI22_X1 U21251 ( .A1(n19285), .A2(n19152), .B1(n19273), .B2(n19166), .ZN(
        n19139) );
  AOI22_X1 U21252 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19274), .B1(
        n19353), .B2(n19168), .ZN(n19138) );
  OAI211_X1 U21253 ( .C1(n19277), .C2(n19155), .A(n19139), .B(n19138), .ZN(
        P3_U2975) );
  INV_X1 U21254 ( .A(n19155), .ZN(n19167) );
  AOI22_X1 U21255 ( .A1(n19296), .A2(n19167), .B1(n19278), .B2(n19166), .ZN(
        n19141) );
  AOI22_X1 U21256 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19280), .B1(
        n19279), .B2(n19168), .ZN(n19140) );
  OAI211_X1 U21257 ( .C1(n19277), .C2(n19171), .A(n19141), .B(n19140), .ZN(
        P3_U2967) );
  AOI22_X1 U21258 ( .A1(n19302), .A2(n19167), .B1(n19284), .B2(n19166), .ZN(
        n19143) );
  AOI22_X1 U21259 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19286), .B1(
        n19285), .B2(n19168), .ZN(n19142) );
  OAI211_X1 U21260 ( .C1(n19283), .C2(n19171), .A(n19143), .B(n19142), .ZN(
        P3_U2959) );
  AOI22_X1 U21261 ( .A1(n19308), .A2(n19167), .B1(n19289), .B2(n19166), .ZN(
        n19145) );
  AOI22_X1 U21262 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19291), .B1(
        n19290), .B2(n19168), .ZN(n19144) );
  OAI211_X1 U21263 ( .C1(n19294), .C2(n19171), .A(n19145), .B(n19144), .ZN(
        P3_U2951) );
  AOI22_X1 U21264 ( .A1(n19308), .A2(n19152), .B1(n19295), .B2(n19166), .ZN(
        n19147) );
  AOI22_X1 U21265 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19297), .B1(
        n19296), .B2(n19168), .ZN(n19146) );
  OAI211_X1 U21266 ( .C1(n19306), .C2(n19155), .A(n19147), .B(n19146), .ZN(
        P3_U2943) );
  AOI22_X1 U21267 ( .A1(n19314), .A2(n19152), .B1(n19301), .B2(n19166), .ZN(
        n19149) );
  AOI22_X1 U21268 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19303), .B1(
        n19302), .B2(n19168), .ZN(n19148) );
  OAI211_X1 U21269 ( .C1(n19312), .C2(n19155), .A(n19149), .B(n19148), .ZN(
        P3_U2935) );
  AOI22_X1 U21270 ( .A1(n19320), .A2(n19152), .B1(n19307), .B2(n19166), .ZN(
        n19151) );
  AOI22_X1 U21271 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19309), .B1(
        n19308), .B2(n19168), .ZN(n19150) );
  OAI211_X1 U21272 ( .C1(n19318), .C2(n19155), .A(n19151), .B(n19150), .ZN(
        P3_U2927) );
  AOI22_X1 U21273 ( .A1(n19326), .A2(n19152), .B1(n19313), .B2(n19166), .ZN(
        n19154) );
  AOI22_X1 U21274 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19315), .B1(
        n19314), .B2(n19168), .ZN(n19153) );
  OAI211_X1 U21275 ( .C1(n19240), .C2(n19155), .A(n19154), .B(n19153), .ZN(
        P3_U2919) );
  AOI22_X1 U21276 ( .A1(n19319), .A2(n19166), .B1(n19337), .B2(n19167), .ZN(
        n19157) );
  AOI22_X1 U21277 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19321), .B1(
        n19320), .B2(n19168), .ZN(n19156) );
  OAI211_X1 U21278 ( .C1(n19240), .C2(n19171), .A(n19157), .B(n19156), .ZN(
        P3_U2911) );
  AOI22_X1 U21279 ( .A1(n19345), .A2(n19167), .B1(n19325), .B2(n19166), .ZN(
        n19159) );
  AOI22_X1 U21280 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19327), .B1(
        n19326), .B2(n19168), .ZN(n19158) );
  OAI211_X1 U21281 ( .C1(n19324), .C2(n19171), .A(n19159), .B(n19158), .ZN(
        P3_U2903) );
  AOI22_X1 U21282 ( .A1(n19330), .A2(n19166), .B1(n19355), .B2(n19167), .ZN(
        n19161) );
  AOI22_X1 U21283 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19332), .B1(
        n19331), .B2(n19168), .ZN(n19160) );
  OAI211_X1 U21284 ( .C1(n19335), .C2(n19171), .A(n19161), .B(n19160), .ZN(
        P3_U2895) );
  AOI22_X1 U21285 ( .A1(n19344), .A2(n19167), .B1(n19336), .B2(n19166), .ZN(
        n19163) );
  AOI22_X1 U21286 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19338), .B1(
        n19337), .B2(n19168), .ZN(n19162) );
  OAI211_X1 U21287 ( .C1(n19341), .C2(n19171), .A(n19163), .B(n19162), .ZN(
        P3_U2887) );
  AOI22_X1 U21288 ( .A1(n19268), .A2(n19167), .B1(n19342), .B2(n19166), .ZN(
        n19165) );
  AOI22_X1 U21289 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19346), .B1(
        n19345), .B2(n19168), .ZN(n19164) );
  OAI211_X1 U21290 ( .C1(n19203), .C2(n19171), .A(n19165), .B(n19164), .ZN(
        P3_U2879) );
  AOI22_X1 U21291 ( .A1(n19353), .A2(n19167), .B1(n19351), .B2(n19166), .ZN(
        n19170) );
  AOI22_X1 U21292 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19356), .B1(
        n19355), .B2(n19168), .ZN(n19169) );
  OAI211_X1 U21293 ( .C1(n19360), .C2(n19171), .A(n19170), .B(n19169), .ZN(
        P3_U2871) );
  INV_X1 U21294 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n19172) );
  INV_X1 U21295 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n20854) );
  AOI22_X1 U21296 ( .A1(n19257), .A2(n19172), .B1(n20854), .B2(U215), .ZN(U253) );
  NAND2_X1 U21297 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19215), .ZN(n19207) );
  NAND2_X1 U21298 ( .A1(n19215), .A2(BUF2_REG_18__SCAN_IN), .ZN(n19213) );
  INV_X1 U21299 ( .A(n19213), .ZN(n19204) );
  NOR2_X2 U21300 ( .A1(n19173), .A2(n20854), .ZN(n19208) );
  AOI22_X1 U21301 ( .A1(n19353), .A2(n19204), .B1(n19260), .B2(n19208), .ZN(
        n19176) );
  NOR2_X2 U21302 ( .A1(n19174), .A2(n19261), .ZN(n19210) );
  AOI22_X1 U21303 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19263), .B1(
        n19344), .B2(n19210), .ZN(n19175) );
  OAI211_X1 U21304 ( .C1(n19219), .C2(n19207), .A(n19176), .B(n19175), .ZN(
        P3_U2990) );
  INV_X1 U21305 ( .A(n19207), .ZN(n19209) );
  AOI22_X1 U21306 ( .A1(n19285), .A2(n19209), .B1(n19267), .B2(n19208), .ZN(
        n19178) );
  AOI22_X1 U21307 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19269), .B1(
        n19268), .B2(n19210), .ZN(n19177) );
  OAI211_X1 U21308 ( .C1(n19219), .C2(n19213), .A(n19178), .B(n19177), .ZN(
        P3_U2982) );
  AOI22_X1 U21309 ( .A1(n19285), .A2(n19204), .B1(n19273), .B2(n19208), .ZN(
        n19180) );
  AOI22_X1 U21310 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19274), .B1(
        n19353), .B2(n19210), .ZN(n19179) );
  OAI211_X1 U21311 ( .C1(n19277), .C2(n19207), .A(n19180), .B(n19179), .ZN(
        P3_U2974) );
  AOI22_X1 U21312 ( .A1(n19290), .A2(n19204), .B1(n19278), .B2(n19208), .ZN(
        n19182) );
  AOI22_X1 U21313 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19280), .B1(
        n19279), .B2(n19210), .ZN(n19181) );
  OAI211_X1 U21314 ( .C1(n19283), .C2(n19207), .A(n19182), .B(n19181), .ZN(
        P3_U2966) );
  AOI22_X1 U21315 ( .A1(n19302), .A2(n19209), .B1(n19284), .B2(n19208), .ZN(
        n19184) );
  AOI22_X1 U21316 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19286), .B1(
        n19285), .B2(n19210), .ZN(n19183) );
  OAI211_X1 U21317 ( .C1(n19283), .C2(n19213), .A(n19184), .B(n19183), .ZN(
        P3_U2958) );
  AOI22_X1 U21318 ( .A1(n19308), .A2(n19209), .B1(n19289), .B2(n19208), .ZN(
        n19186) );
  AOI22_X1 U21319 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19291), .B1(
        n19290), .B2(n19210), .ZN(n19185) );
  OAI211_X1 U21320 ( .C1(n19294), .C2(n19213), .A(n19186), .B(n19185), .ZN(
        P3_U2950) );
  AOI22_X1 U21321 ( .A1(n19308), .A2(n19204), .B1(n19295), .B2(n19208), .ZN(
        n19188) );
  AOI22_X1 U21322 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19297), .B1(
        n19296), .B2(n19210), .ZN(n19187) );
  OAI211_X1 U21323 ( .C1(n19306), .C2(n19207), .A(n19188), .B(n19187), .ZN(
        P3_U2942) );
  AOI22_X1 U21324 ( .A1(n19320), .A2(n19209), .B1(n19301), .B2(n19208), .ZN(
        n19190) );
  AOI22_X1 U21325 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19303), .B1(
        n19302), .B2(n19210), .ZN(n19189) );
  OAI211_X1 U21326 ( .C1(n19306), .C2(n19213), .A(n19190), .B(n19189), .ZN(
        P3_U2934) );
  AOI22_X1 U21327 ( .A1(n19326), .A2(n19209), .B1(n19307), .B2(n19208), .ZN(
        n19192) );
  AOI22_X1 U21328 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19309), .B1(
        n19308), .B2(n19210), .ZN(n19191) );
  OAI211_X1 U21329 ( .C1(n19312), .C2(n19213), .A(n19192), .B(n19191), .ZN(
        P3_U2926) );
  AOI22_X1 U21330 ( .A1(n19326), .A2(n19204), .B1(n19313), .B2(n19208), .ZN(
        n19194) );
  AOI22_X1 U21331 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19315), .B1(
        n19314), .B2(n19210), .ZN(n19193) );
  OAI211_X1 U21332 ( .C1(n19240), .C2(n19207), .A(n19194), .B(n19193), .ZN(
        P3_U2918) );
  AOI22_X1 U21333 ( .A1(n19319), .A2(n19208), .B1(n19337), .B2(n19209), .ZN(
        n19196) );
  AOI22_X1 U21334 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19321), .B1(
        n19320), .B2(n19210), .ZN(n19195) );
  OAI211_X1 U21335 ( .C1(n19240), .C2(n19213), .A(n19196), .B(n19195), .ZN(
        P3_U2910) );
  AOI22_X1 U21336 ( .A1(n19337), .A2(n19204), .B1(n19325), .B2(n19208), .ZN(
        n19198) );
  AOI22_X1 U21337 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19327), .B1(
        n19326), .B2(n19210), .ZN(n19197) );
  OAI211_X1 U21338 ( .C1(n19335), .C2(n19207), .A(n19198), .B(n19197), .ZN(
        P3_U2902) );
  AOI22_X1 U21339 ( .A1(n19345), .A2(n19204), .B1(n19330), .B2(n19208), .ZN(
        n19200) );
  AOI22_X1 U21340 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19332), .B1(
        n19331), .B2(n19210), .ZN(n19199) );
  OAI211_X1 U21341 ( .C1(n19341), .C2(n19207), .A(n19200), .B(n19199), .ZN(
        P3_U2894) );
  AOI22_X1 U21342 ( .A1(n19355), .A2(n19204), .B1(n19336), .B2(n19208), .ZN(
        n19202) );
  AOI22_X1 U21343 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19338), .B1(
        n19337), .B2(n19210), .ZN(n19201) );
  OAI211_X1 U21344 ( .C1(n19203), .C2(n19207), .A(n19202), .B(n19201), .ZN(
        P3_U2886) );
  AOI22_X1 U21345 ( .A1(n19344), .A2(n19204), .B1(n19342), .B2(n19208), .ZN(
        n19206) );
  AOI22_X1 U21346 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19346), .B1(
        n19345), .B2(n19210), .ZN(n19205) );
  OAI211_X1 U21347 ( .C1(n19360), .C2(n19207), .A(n19206), .B(n19205), .ZN(
        P3_U2878) );
  AOI22_X1 U21348 ( .A1(n19353), .A2(n19209), .B1(n19351), .B2(n19208), .ZN(
        n19212) );
  AOI22_X1 U21349 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19356), .B1(
        n19355), .B2(n19210), .ZN(n19211) );
  OAI211_X1 U21350 ( .C1(n19360), .C2(n19213), .A(n19212), .B(n19211), .ZN(
        P3_U2870) );
  OAI22_X1 U21351 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19257), .ZN(n19214) );
  INV_X1 U21352 ( .A(n19214), .ZN(U252) );
  NAND2_X1 U21353 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19215), .ZN(n19256) );
  NAND2_X1 U21354 ( .A1(n19215), .A2(BUF2_REG_17__SCAN_IN), .ZN(n19248) );
  INV_X1 U21355 ( .A(n19248), .ZN(n19252) );
  AND2_X1 U21356 ( .A1(n19259), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19251) );
  AOI22_X1 U21357 ( .A1(n19353), .A2(n19252), .B1(n19260), .B2(n19251), .ZN(
        n19218) );
  NOR2_X2 U21358 ( .A1(n19216), .A2(n19261), .ZN(n19253) );
  AOI22_X1 U21359 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19263), .B1(
        n19344), .B2(n19253), .ZN(n19217) );
  OAI211_X1 U21360 ( .C1(n19219), .C2(n19256), .A(n19218), .B(n19217), .ZN(
        P3_U2989) );
  AOI22_X1 U21361 ( .A1(n19279), .A2(n19252), .B1(n19267), .B2(n19251), .ZN(
        n19221) );
  AOI22_X1 U21362 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19269), .B1(
        n19268), .B2(n19253), .ZN(n19220) );
  OAI211_X1 U21363 ( .C1(n19272), .C2(n19256), .A(n19221), .B(n19220), .ZN(
        P3_U2981) );
  AOI22_X1 U21364 ( .A1(n19285), .A2(n19252), .B1(n19273), .B2(n19251), .ZN(
        n19223) );
  AOI22_X1 U21365 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19274), .B1(
        n19353), .B2(n19253), .ZN(n19222) );
  OAI211_X1 U21366 ( .C1(n19277), .C2(n19256), .A(n19223), .B(n19222), .ZN(
        P3_U2973) );
  INV_X1 U21367 ( .A(n19256), .ZN(n19245) );
  AOI22_X1 U21368 ( .A1(n19296), .A2(n19245), .B1(n19278), .B2(n19251), .ZN(
        n19225) );
  AOI22_X1 U21369 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19280), .B1(
        n19279), .B2(n19253), .ZN(n19224) );
  OAI211_X1 U21370 ( .C1(n19277), .C2(n19248), .A(n19225), .B(n19224), .ZN(
        P3_U2965) );
  AOI22_X1 U21371 ( .A1(n19296), .A2(n19252), .B1(n19284), .B2(n19251), .ZN(
        n19227) );
  AOI22_X1 U21372 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19286), .B1(
        n19285), .B2(n19253), .ZN(n19226) );
  OAI211_X1 U21373 ( .C1(n19294), .C2(n19256), .A(n19227), .B(n19226), .ZN(
        P3_U2957) );
  AOI22_X1 U21374 ( .A1(n19302), .A2(n19252), .B1(n19289), .B2(n19251), .ZN(
        n19229) );
  AOI22_X1 U21375 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19291), .B1(
        n19290), .B2(n19253), .ZN(n19228) );
  OAI211_X1 U21376 ( .C1(n19300), .C2(n19256), .A(n19229), .B(n19228), .ZN(
        P3_U2949) );
  AOI22_X1 U21377 ( .A1(n19314), .A2(n19245), .B1(n19295), .B2(n19251), .ZN(
        n19231) );
  AOI22_X1 U21378 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19297), .B1(
        n19296), .B2(n19253), .ZN(n19230) );
  OAI211_X1 U21379 ( .C1(n19300), .C2(n19248), .A(n19231), .B(n19230), .ZN(
        P3_U2941) );
  AOI22_X1 U21380 ( .A1(n19320), .A2(n19245), .B1(n19301), .B2(n19251), .ZN(
        n19233) );
  AOI22_X1 U21381 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19303), .B1(
        n19302), .B2(n19253), .ZN(n19232) );
  OAI211_X1 U21382 ( .C1(n19306), .C2(n19248), .A(n19233), .B(n19232), .ZN(
        P3_U2933) );
  AOI22_X1 U21383 ( .A1(n19326), .A2(n19245), .B1(n19307), .B2(n19251), .ZN(
        n19235) );
  AOI22_X1 U21384 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19309), .B1(
        n19308), .B2(n19253), .ZN(n19234) );
  OAI211_X1 U21385 ( .C1(n19312), .C2(n19248), .A(n19235), .B(n19234), .ZN(
        P3_U2925) );
  AOI22_X1 U21386 ( .A1(n19331), .A2(n19245), .B1(n19313), .B2(n19251), .ZN(
        n19237) );
  AOI22_X1 U21387 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19315), .B1(
        n19314), .B2(n19253), .ZN(n19236) );
  OAI211_X1 U21388 ( .C1(n19318), .C2(n19248), .A(n19237), .B(n19236), .ZN(
        P3_U2917) );
  AOI22_X1 U21389 ( .A1(n19319), .A2(n19251), .B1(n19337), .B2(n19245), .ZN(
        n19239) );
  AOI22_X1 U21390 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19321), .B1(
        n19320), .B2(n19253), .ZN(n19238) );
  OAI211_X1 U21391 ( .C1(n19240), .C2(n19248), .A(n19239), .B(n19238), .ZN(
        P3_U2909) );
  AOI22_X1 U21392 ( .A1(n19345), .A2(n19245), .B1(n19325), .B2(n19251), .ZN(
        n19242) );
  AOI22_X1 U21393 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19327), .B1(
        n19326), .B2(n19253), .ZN(n19241) );
  OAI211_X1 U21394 ( .C1(n19324), .C2(n19248), .A(n19242), .B(n19241), .ZN(
        P3_U2901) );
  AOI22_X1 U21395 ( .A1(n19345), .A2(n19252), .B1(n19330), .B2(n19251), .ZN(
        n19244) );
  AOI22_X1 U21396 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19332), .B1(
        n19331), .B2(n19253), .ZN(n19243) );
  OAI211_X1 U21397 ( .C1(n19341), .C2(n19256), .A(n19244), .B(n19243), .ZN(
        P3_U2893) );
  AOI22_X1 U21398 ( .A1(n19344), .A2(n19245), .B1(n19336), .B2(n19251), .ZN(
        n19247) );
  AOI22_X1 U21399 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19338), .B1(
        n19337), .B2(n19253), .ZN(n19246) );
  OAI211_X1 U21400 ( .C1(n19341), .C2(n19248), .A(n19247), .B(n19246), .ZN(
        P3_U2885) );
  AOI22_X1 U21401 ( .A1(n19344), .A2(n19252), .B1(n19342), .B2(n19251), .ZN(
        n19250) );
  AOI22_X1 U21402 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19346), .B1(
        n19345), .B2(n19253), .ZN(n19249) );
  OAI211_X1 U21403 ( .C1(n19360), .C2(n19256), .A(n19250), .B(n19249), .ZN(
        P3_U2877) );
  AOI22_X1 U21404 ( .A1(n19268), .A2(n19252), .B1(n19351), .B2(n19251), .ZN(
        n19255) );
  AOI22_X1 U21405 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19356), .B1(
        n19355), .B2(n19253), .ZN(n19254) );
  OAI211_X1 U21406 ( .C1(n19266), .C2(n19256), .A(n19255), .B(n19254), .ZN(
        P3_U2869) );
  OAI22_X1 U21407 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19257), .ZN(n19258) );
  INV_X1 U21408 ( .A(n19258), .ZN(U251) );
  NAND2_X1 U21409 ( .A1(n19215), .A2(BUF2_REG_16__SCAN_IN), .ZN(n19359) );
  NAND2_X1 U21410 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19215), .ZN(n19349) );
  INV_X1 U21411 ( .A(n19349), .ZN(n19352) );
  AND2_X1 U21412 ( .A1(n19259), .A2(BUF2_REG_0__SCAN_IN), .ZN(n19350) );
  AOI22_X1 U21413 ( .A1(n19279), .A2(n19352), .B1(n19260), .B2(n19350), .ZN(
        n19265) );
  NOR2_X2 U21414 ( .A1(n19262), .A2(n19261), .ZN(n19354) );
  AOI22_X1 U21415 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19263), .B1(
        n19344), .B2(n19354), .ZN(n19264) );
  OAI211_X1 U21416 ( .C1(n19266), .C2(n19359), .A(n19265), .B(n19264), .ZN(
        P3_U2988) );
  INV_X1 U21417 ( .A(n19359), .ZN(n19343) );
  AOI22_X1 U21418 ( .A1(n19279), .A2(n19343), .B1(n19267), .B2(n19350), .ZN(
        n19271) );
  AOI22_X1 U21419 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19269), .B1(
        n19268), .B2(n19354), .ZN(n19270) );
  OAI211_X1 U21420 ( .C1(n19272), .C2(n19349), .A(n19271), .B(n19270), .ZN(
        P3_U2980) );
  AOI22_X1 U21421 ( .A1(n19285), .A2(n19343), .B1(n19273), .B2(n19350), .ZN(
        n19276) );
  AOI22_X1 U21422 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19274), .B1(
        n19353), .B2(n19354), .ZN(n19275) );
  OAI211_X1 U21423 ( .C1(n19277), .C2(n19349), .A(n19276), .B(n19275), .ZN(
        P3_U2972) );
  AOI22_X1 U21424 ( .A1(n19290), .A2(n19343), .B1(n19278), .B2(n19350), .ZN(
        n19282) );
  AOI22_X1 U21425 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19280), .B1(
        n19279), .B2(n19354), .ZN(n19281) );
  OAI211_X1 U21426 ( .C1(n19283), .C2(n19349), .A(n19282), .B(n19281), .ZN(
        P3_U2964) );
  AOI22_X1 U21427 ( .A1(n19296), .A2(n19343), .B1(n19284), .B2(n19350), .ZN(
        n19288) );
  AOI22_X1 U21428 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19286), .B1(
        n19285), .B2(n19354), .ZN(n19287) );
  OAI211_X1 U21429 ( .C1(n19294), .C2(n19349), .A(n19288), .B(n19287), .ZN(
        P3_U2956) );
  AOI22_X1 U21430 ( .A1(n19308), .A2(n19352), .B1(n19289), .B2(n19350), .ZN(
        n19293) );
  AOI22_X1 U21431 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19291), .B1(
        n19290), .B2(n19354), .ZN(n19292) );
  OAI211_X1 U21432 ( .C1(n19294), .C2(n19359), .A(n19293), .B(n19292), .ZN(
        P3_U2948) );
  AOI22_X1 U21433 ( .A1(n19314), .A2(n19352), .B1(n19295), .B2(n19350), .ZN(
        n19299) );
  AOI22_X1 U21434 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19297), .B1(
        n19296), .B2(n19354), .ZN(n19298) );
  OAI211_X1 U21435 ( .C1(n19300), .C2(n19359), .A(n19299), .B(n19298), .ZN(
        P3_U2940) );
  AOI22_X1 U21436 ( .A1(n19320), .A2(n19352), .B1(n19301), .B2(n19350), .ZN(
        n19305) );
  AOI22_X1 U21437 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19303), .B1(
        n19302), .B2(n19354), .ZN(n19304) );
  OAI211_X1 U21438 ( .C1(n19306), .C2(n19359), .A(n19305), .B(n19304), .ZN(
        P3_U2932) );
  AOI22_X1 U21439 ( .A1(n19326), .A2(n19352), .B1(n19307), .B2(n19350), .ZN(
        n19311) );
  AOI22_X1 U21440 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19309), .B1(
        n19308), .B2(n19354), .ZN(n19310) );
  OAI211_X1 U21441 ( .C1(n19312), .C2(n19359), .A(n19311), .B(n19310), .ZN(
        P3_U2924) );
  AOI22_X1 U21442 ( .A1(n19331), .A2(n19352), .B1(n19313), .B2(n19350), .ZN(
        n19317) );
  AOI22_X1 U21443 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19315), .B1(
        n19314), .B2(n19354), .ZN(n19316) );
  OAI211_X1 U21444 ( .C1(n19318), .C2(n19359), .A(n19317), .B(n19316), .ZN(
        P3_U2916) );
  AOI22_X1 U21445 ( .A1(n19331), .A2(n19343), .B1(n19319), .B2(n19350), .ZN(
        n19323) );
  AOI22_X1 U21446 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19321), .B1(
        n19320), .B2(n19354), .ZN(n19322) );
  OAI211_X1 U21447 ( .C1(n19324), .C2(n19349), .A(n19323), .B(n19322), .ZN(
        P3_U2908) );
  AOI22_X1 U21448 ( .A1(n19337), .A2(n19343), .B1(n19325), .B2(n19350), .ZN(
        n19329) );
  AOI22_X1 U21449 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19327), .B1(
        n19326), .B2(n19354), .ZN(n19328) );
  OAI211_X1 U21450 ( .C1(n19335), .C2(n19349), .A(n19329), .B(n19328), .ZN(
        P3_U2900) );
  AOI22_X1 U21451 ( .A1(n19330), .A2(n19350), .B1(n19355), .B2(n19352), .ZN(
        n19334) );
  AOI22_X1 U21452 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19332), .B1(
        n19331), .B2(n19354), .ZN(n19333) );
  OAI211_X1 U21453 ( .C1(n19335), .C2(n19359), .A(n19334), .B(n19333), .ZN(
        P3_U2892) );
  AOI22_X1 U21454 ( .A1(n19344), .A2(n19352), .B1(n19336), .B2(n19350), .ZN(
        n19340) );
  AOI22_X1 U21455 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19338), .B1(
        n19337), .B2(n19354), .ZN(n19339) );
  OAI211_X1 U21456 ( .C1(n19341), .C2(n19359), .A(n19340), .B(n19339), .ZN(
        P3_U2884) );
  AOI22_X1 U21457 ( .A1(n19344), .A2(n19343), .B1(n19342), .B2(n19350), .ZN(
        n19348) );
  AOI22_X1 U21458 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19346), .B1(
        n19345), .B2(n19354), .ZN(n19347) );
  OAI211_X1 U21459 ( .C1(n19360), .C2(n19349), .A(n19348), .B(n19347), .ZN(
        P3_U2876) );
  AOI22_X1 U21460 ( .A1(n19353), .A2(n19352), .B1(n19351), .B2(n19350), .ZN(
        n19358) );
  AOI22_X1 U21461 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19356), .B1(
        n19355), .B2(n19354), .ZN(n19357) );
  OAI211_X1 U21462 ( .C1(n19360), .C2(n19359), .A(n19358), .B(n19357), .ZN(
        P3_U2868) );
  AOI22_X1 U21463 ( .A1(n19369), .A2(n19361), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n19579), .ZN(n19362) );
  OAI21_X1 U21464 ( .B1(n19367), .B2(n19363), .A(n19362), .ZN(P2_U2905) );
  AOI22_X1 U21465 ( .A1(n19369), .A2(n19364), .B1(P2_EAX_REG_11__SCAN_IN), 
        .B2(n19579), .ZN(n19365) );
  OAI21_X1 U21466 ( .B1(n19367), .B2(n19366), .A(n19365), .ZN(P2_U2908) );
  INV_X1 U21467 ( .A(n19367), .ZN(n19371) );
  AOI22_X1 U21468 ( .A1(n19371), .A2(n19370), .B1(n19369), .B2(n19368), .ZN(
        n19372) );
  OAI21_X1 U21469 ( .B1(n19374), .B2(n19373), .A(n19372), .ZN(P2_U2910) );
  NOR3_X4 U21470 ( .A1(n21819), .A2(n19375), .A3(n19391), .ZN(n19843) );
  NOR3_X4 U21471 ( .A1(n19376), .A2(n21819), .A3(n19391), .ZN(n19842) );
  AOI22_X1 U21472 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19843), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19842), .ZN(n19578) );
  NAND3_X1 U21473 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19389) );
  INV_X1 U21474 ( .A(n19570), .ZN(n19840) );
  OAI21_X1 U21475 ( .B1(n19383), .B2(n19840), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19377) );
  OAI21_X1 U21476 ( .B1(n19389), .B2(n19549), .A(n19377), .ZN(n19841) );
  NOR2_X2 U21477 ( .A1(n19380), .A2(n19839), .ZN(n19562) );
  AOI22_X1 U21478 ( .A1(n19841), .A2(n19379), .B1(n19840), .B2(n19562), .ZN(
        n19388) );
  AOI22_X1 U21479 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19843), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19842), .ZN(n19533) );
  OAI21_X1 U21480 ( .B1(n19381), .B2(n21819), .A(n19389), .ZN(n19386) );
  NAND2_X1 U21481 ( .A1(n19459), .A2(n19382), .ZN(n19553) );
  INV_X1 U21482 ( .A(n19553), .ZN(n19568) );
  AOI211_X1 U21483 ( .C1(n19383), .C2(n19568), .A(n19840), .B(n19564), .ZN(
        n19384) );
  NOR2_X1 U21484 ( .A1(n19837), .A2(n19384), .ZN(n19385) );
  NAND2_X1 U21485 ( .A1(n19386), .A2(n19385), .ZN(n19844) );
  AOI22_X1 U21486 ( .A1(n19563), .A2(n19796), .B1(
        P2_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n19844), .ZN(n19387) );
  OAI211_X1 U21487 ( .C1(n19578), .C2(n19950), .A(n19388), .B(n19387), .ZN(
        P2_U3175) );
  INV_X1 U21488 ( .A(n19860), .ZN(n19849) );
  NOR2_X1 U21489 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19389), .ZN(
        n19848) );
  AOI22_X1 U21490 ( .A1(n19563), .A2(n19849), .B1(n19562), .B2(n19848), .ZN(
        n19399) );
  NAND3_X1 U21491 ( .A1(n19854), .A2(n19564), .A3(n19860), .ZN(n19390) );
  NAND2_X1 U21492 ( .A1(n19564), .A2(n21819), .ZN(n19565) );
  NAND2_X1 U21493 ( .A1(n19390), .A2(n19565), .ZN(n19394) );
  NAND3_X1 U21494 ( .A1(n19523), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19413) );
  NOR2_X1 U21495 ( .A1(n19424), .A2(n19413), .ZN(n19855) );
  INV_X1 U21496 ( .A(n19855), .ZN(n19403) );
  INV_X1 U21497 ( .A(n19391), .ZN(n19567) );
  AOI21_X1 U21498 ( .B1(n19395), .B2(n19568), .A(n19567), .ZN(n19392) );
  AOI21_X1 U21499 ( .B1(n19394), .B2(n19403), .A(n19392), .ZN(n19393) );
  OAI21_X1 U21500 ( .B1(n19848), .B2(n19855), .A(n19394), .ZN(n19397) );
  OAI21_X1 U21501 ( .B1(n19395), .B2(n19848), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19396) );
  NAND2_X1 U21502 ( .A1(n19397), .A2(n19396), .ZN(n19850) );
  AOI22_X1 U21503 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19851), .B1(
        n19379), .B2(n19850), .ZN(n19398) );
  OAI211_X1 U21504 ( .C1(n19578), .C2(n19854), .A(n19399), .B(n19398), .ZN(
        P2_U3167) );
  OAI21_X1 U21505 ( .B1(n19400), .B2(n19855), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19401) );
  OAI21_X1 U21506 ( .B1(n19413), .B2(n19549), .A(n19401), .ZN(n19856) );
  AOI22_X1 U21507 ( .A1(n19856), .A2(n19379), .B1(n19562), .B2(n19855), .ZN(
        n19407) );
  NOR2_X2 U21508 ( .A1(n19402), .A2(n19557), .ZN(n19863) );
  NAND2_X1 U21509 ( .A1(n19408), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19554) );
  OAI21_X1 U21510 ( .B1(n19402), .B2(n19554), .A(n19413), .ZN(n19405) );
  OAI211_X1 U21511 ( .C1(n11628), .C2(n19553), .A(n19403), .B(n19549), .ZN(
        n19404) );
  NAND3_X1 U21512 ( .A1(n19405), .A2(n19571), .A3(n19404), .ZN(n19857) );
  AOI22_X1 U21513 ( .A1(n19563), .A2(n19863), .B1(
        P2_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n19857), .ZN(n19406) );
  OAI211_X1 U21514 ( .C1(n19578), .C2(n19860), .A(n19407), .B(n19406), .ZN(
        P2_U3159) );
  NOR2_X1 U21515 ( .A1(n19408), .A2(n19455), .ZN(n19503) );
  INV_X1 U21516 ( .A(n19503), .ZN(n19409) );
  INV_X1 U21517 ( .A(n19410), .ZN(n19415) );
  INV_X1 U21518 ( .A(n19411), .ZN(n19412) );
  NAND2_X1 U21519 ( .A1(n19412), .A2(n19481), .ZN(n19506) );
  NOR2_X1 U21520 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19413), .ZN(
        n19861) );
  OAI21_X1 U21521 ( .B1(n19417), .B2(n19861), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19414) );
  OAI21_X1 U21522 ( .B1(n19415), .B2(n19506), .A(n19414), .ZN(n19862) );
  AOI22_X1 U21523 ( .A1(n19862), .A2(n19379), .B1(n19562), .B2(n19861), .ZN(
        n19422) );
  INV_X1 U21524 ( .A(n19873), .ZN(n19803) );
  OAI21_X1 U21525 ( .B1(n19803), .B2(n19863), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19416) );
  OAI21_X1 U21526 ( .B1(n19506), .B2(n14101), .A(n19416), .ZN(n19420) );
  AOI211_X1 U21527 ( .C1(n19417), .C2(n19568), .A(n19564), .B(n19861), .ZN(
        n19418) );
  NOR2_X1 U21528 ( .A1(n19837), .A2(n19418), .ZN(n19419) );
  NAND2_X1 U21529 ( .A1(n19420), .A2(n19419), .ZN(n19864) );
  INV_X1 U21530 ( .A(n19578), .ZN(n19520) );
  AOI22_X1 U21531 ( .A1(n19864), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n19520), .B2(n19863), .ZN(n19421) );
  OAI211_X1 U21532 ( .C1(n19533), .C2(n19873), .A(n19422), .B(n19421), .ZN(
        P2_U3151) );
  NAND2_X1 U21533 ( .A1(n19423), .A2(n19455), .ZN(n19517) );
  NAND3_X1 U21534 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n19518), .ZN(n19433) );
  NOR2_X1 U21535 ( .A1(n19424), .A2(n19433), .ZN(n19867) );
  OAI21_X1 U21536 ( .B1(n11508), .B2(n19867), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19425) );
  OAI21_X1 U21537 ( .B1(n19433), .B2(n19549), .A(n19425), .ZN(n19868) );
  AOI22_X1 U21538 ( .A1(n19868), .A2(n19379), .B1(n19562), .B2(n19867), .ZN(
        n19431) );
  OAI21_X1 U21539 ( .B1(n19426), .B2(n19522), .A(n19433), .ZN(n19429) );
  INV_X1 U21540 ( .A(n19867), .ZN(n19427) );
  OAI211_X1 U21541 ( .C1(n11624), .C2(n19553), .A(n19427), .B(n19549), .ZN(
        n19428) );
  NAND3_X1 U21542 ( .A1(n19429), .A2(n19571), .A3(n19428), .ZN(n19869) );
  AOI22_X1 U21543 ( .A1(n19520), .A2(n19803), .B1(
        P2_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n19869), .ZN(n19430) );
  OAI211_X1 U21544 ( .C1(n19533), .C2(n19879), .A(n19431), .B(n19430), .ZN(
        P2_U3143) );
  NOR2_X1 U21545 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19433), .ZN(
        n19874) );
  AOI22_X1 U21546 ( .A1(n19563), .A2(n19881), .B1(n19562), .B2(n19874), .ZN(
        n19444) );
  OAI21_X1 U21547 ( .B1(n19881), .B2(n19870), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19434) );
  NAND2_X1 U21548 ( .A1(n19434), .A2(n19564), .ZN(n19442) );
  NAND3_X1 U21549 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19518), .A3(
        n19523), .ZN(n19456) );
  INV_X1 U21550 ( .A(n19456), .ZN(n19449) );
  NAND2_X1 U21551 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19449), .ZN(
        n19446) );
  INV_X1 U21552 ( .A(n19874), .ZN(n19435) );
  NAND2_X1 U21553 ( .A1(n19446), .A2(n19435), .ZN(n19438) );
  NAND2_X1 U21554 ( .A1(n19439), .A2(n19459), .ZN(n19436) );
  AOI21_X1 U21555 ( .B1(n19436), .B2(n19435), .A(n19837), .ZN(n19437) );
  INV_X1 U21556 ( .A(n19438), .ZN(n19441) );
  OAI21_X1 U21557 ( .B1(n19439), .B2(n19874), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19440) );
  AOI22_X1 U21558 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19876), .B1(
        n19379), .B2(n19875), .ZN(n19443) );
  OAI211_X1 U21559 ( .C1(n19578), .C2(n19879), .A(n19444), .B(n19443), .ZN(
        P2_U3135) );
  INV_X1 U21560 ( .A(n19446), .ZN(n19880) );
  AOI22_X1 U21561 ( .A1(n19520), .A2(n19881), .B1(n19562), .B2(n19880), .ZN(
        n19454) );
  OAI21_X1 U21562 ( .B1(n19445), .B2(n19554), .A(n19564), .ZN(n19452) );
  OAI211_X1 U21563 ( .C1(n19447), .C2(n19553), .A(n19446), .B(n19549), .ZN(
        n19448) );
  OAI211_X1 U21564 ( .C1(n19452), .C2(n19449), .A(n19571), .B(n19448), .ZN(
        n19883) );
  OAI21_X1 U21565 ( .B1(n19450), .B2(n19880), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19451) );
  OAI21_X1 U21566 ( .B1(n19452), .B2(n19456), .A(n19451), .ZN(n19882) );
  AOI22_X1 U21567 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19883), .B1(
        n19379), .B2(n19882), .ZN(n19453) );
  OAI211_X1 U21568 ( .C1(n19533), .C2(n19886), .A(n19454), .B(n19453), .ZN(
        P2_U3127) );
  NOR2_X1 U21569 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19456), .ZN(
        n19887) );
  AOI22_X1 U21570 ( .A1(n19563), .A2(n19813), .B1(n19887), .B2(n19562), .ZN(
        n19466) );
  NAND3_X1 U21571 ( .A1(n19899), .A2(n19564), .A3(n19886), .ZN(n19457) );
  NAND2_X1 U21572 ( .A1(n19457), .A2(n19565), .ZN(n19462) );
  NOR2_X1 U21573 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19518), .ZN(
        n19492) );
  NAND2_X1 U21574 ( .A1(n19458), .A2(n19492), .ZN(n19471) );
  OAI21_X1 U21575 ( .B1(n11620), .B2(n19470), .A(n19459), .ZN(n19460) );
  AOI21_X1 U21576 ( .B1(n19462), .B2(n19471), .A(n19460), .ZN(n19461) );
  INV_X1 U21577 ( .A(n19471), .ZN(n19893) );
  OAI21_X1 U21578 ( .B1(n19893), .B2(n19887), .A(n19462), .ZN(n19464) );
  OAI21_X1 U21579 ( .B1(n11620), .B2(n19887), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19463) );
  NAND2_X1 U21580 ( .A1(n19464), .A2(n19463), .ZN(n19889) );
  AOI22_X1 U21581 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19890), .B1(
        n19889), .B2(n19379), .ZN(n19465) );
  OAI211_X1 U21582 ( .C1(n19578), .C2(n19886), .A(n19466), .B(n19465), .ZN(
        P2_U3119) );
  NOR2_X1 U21583 ( .A1(n19468), .A2(n19893), .ZN(n19472) );
  NAND2_X1 U21584 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19492), .ZN(
        n19469) );
  OAI22_X1 U21585 ( .A1(n19472), .A2(n19470), .B1(n19469), .B2(n19549), .ZN(
        n19894) );
  AOI22_X1 U21586 ( .A1(n19894), .A2(n19379), .B1(n19893), .B2(n19562), .ZN(
        n19477) );
  OAI22_X1 U21587 ( .A1(n19472), .A2(n19553), .B1(n19837), .B2(n19471), .ZN(
        n19475) );
  INV_X1 U21588 ( .A(n19492), .ZN(n19490) );
  OAI22_X1 U21589 ( .A1(n19523), .A2(n19490), .B1(n21819), .B2(n19473), .ZN(
        n19474) );
  OAI21_X1 U21590 ( .B1(n19567), .B2(n19475), .A(n19474), .ZN(n19896) );
  AOI22_X1 U21591 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19896), .B1(
        n19813), .B2(n19520), .ZN(n19476) );
  OAI211_X1 U21592 ( .C1(n19533), .C2(n19905), .A(n19477), .B(n19476), .ZN(
        P2_U3111) );
  NOR2_X1 U21593 ( .A1(n19534), .A2(n19490), .ZN(n19900) );
  OAI21_X1 U21594 ( .B1(n19478), .B2(n19900), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19479) );
  OAI21_X1 U21595 ( .B1(n19535), .B2(n19490), .A(n19479), .ZN(n19901) );
  AOI22_X1 U21596 ( .A1(n19901), .A2(n19379), .B1(n19562), .B2(n19900), .ZN(
        n19487) );
  INV_X1 U21597 ( .A(n19900), .ZN(n19480) );
  OAI211_X1 U21598 ( .C1(n11633), .C2(n19553), .A(n19480), .B(n19549), .ZN(
        n19485) );
  INV_X1 U21599 ( .A(n19481), .ZN(n19482) );
  NAND2_X1 U21600 ( .A1(n19492), .A2(n19482), .ZN(n19483) );
  OAI221_X1 U21601 ( .B1(n21819), .B2(n19818), .C1(n21819), .C2(n19905), .A(
        n19483), .ZN(n19484) );
  NAND3_X1 U21602 ( .A1(n19485), .A2(n19571), .A3(n19484), .ZN(n19902) );
  AOI22_X1 U21603 ( .A1(n19563), .A2(n19907), .B1(
        P2_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n19902), .ZN(n19486) );
  OAI211_X1 U21604 ( .C1(n19578), .C2(n19905), .A(n19487), .B(n19486), .ZN(
        P2_U3103) );
  INV_X1 U21605 ( .A(n19557), .ZN(n19488) );
  NOR2_X1 U21606 ( .A1(n19547), .A2(n19490), .ZN(n19906) );
  AOI22_X1 U21607 ( .A1(n19520), .A2(n19907), .B1(n19562), .B2(n19906), .ZN(
        n19501) );
  OAI21_X1 U21608 ( .B1(n19491), .B2(n19554), .A(n19564), .ZN(n19499) );
  NAND2_X1 U21609 ( .A1(n19492), .A2(n19523), .ZN(n19504) );
  INV_X1 U21610 ( .A(n19504), .ZN(n19496) );
  OAI21_X1 U21611 ( .B1(n19564), .B2(n19906), .A(n19571), .ZN(n19493) );
  OAI21_X1 U21612 ( .B1(n19494), .B2(n19553), .A(n19493), .ZN(n19495) );
  OAI21_X1 U21613 ( .B1(n19499), .B2(n19496), .A(n19495), .ZN(n19909) );
  OAI21_X1 U21614 ( .B1(n19497), .B2(n19906), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19498) );
  OAI21_X1 U21615 ( .B1(n19499), .B2(n19504), .A(n19498), .ZN(n19908) );
  AOI22_X1 U21616 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19909), .B1(
        n19379), .B2(n19908), .ZN(n19500) );
  OAI211_X1 U21617 ( .C1(n19533), .C2(n19912), .A(n19501), .B(n19500), .ZN(
        P2_U3095) );
  NOR2_X1 U21618 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19504), .ZN(
        n19913) );
  AOI22_X1 U21619 ( .A1(n19520), .A2(n19914), .B1(n19913), .B2(n19562), .ZN(
        n19516) );
  OAI21_X1 U21620 ( .B1(n19658), .B2(n19914), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19505) );
  NAND2_X1 U21621 ( .A1(n19505), .A2(n19564), .ZN(n19514) );
  NOR2_X1 U21622 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19506), .ZN(
        n19510) );
  INV_X1 U21623 ( .A(n19913), .ZN(n19508) );
  INV_X1 U21624 ( .A(n11632), .ZN(n19511) );
  NOR2_X1 U21625 ( .A1(n19913), .A2(n19511), .ZN(n19507) );
  AOI211_X1 U21626 ( .C1(n19553), .C2(n19508), .A(n19837), .B(n19507), .ZN(
        n19509) );
  INV_X1 U21627 ( .A(n19510), .ZN(n19513) );
  OAI21_X1 U21628 ( .B1(n19511), .B2(n19913), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19512) );
  AOI22_X1 U21629 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19916), .B1(
        n19379), .B2(n19915), .ZN(n19515) );
  OAI211_X1 U21630 ( .C1(n19533), .C2(n19925), .A(n19516), .B(n19515), .ZN(
        P2_U3087) );
  NAND2_X1 U21631 ( .A1(n14101), .A2(n19518), .ZN(n19546) );
  NOR2_X1 U21632 ( .A1(n19519), .A2(n19546), .ZN(n19919) );
  AOI22_X1 U21633 ( .A1(n19520), .A2(n19658), .B1(n19562), .B2(n19919), .ZN(
        n19532) );
  OAI21_X1 U21634 ( .B1(n19522), .B2(n19521), .A(n19564), .ZN(n19530) );
  NOR2_X1 U21635 ( .A1(n19523), .A2(n19546), .ZN(n19527) );
  OAI21_X1 U21636 ( .B1(n19564), .B2(n19919), .A(n19571), .ZN(n19524) );
  OAI21_X1 U21637 ( .B1(n19525), .B2(n19553), .A(n19524), .ZN(n19526) );
  OAI21_X1 U21638 ( .B1(n19530), .B2(n19527), .A(n19526), .ZN(n19922) );
  INV_X1 U21639 ( .A(n19527), .ZN(n19529) );
  OAI21_X1 U21640 ( .B1(n11619), .B2(n19919), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19528) );
  OAI21_X1 U21641 ( .B1(n19530), .B2(n19529), .A(n19528), .ZN(n19921) );
  AOI22_X1 U21642 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19922), .B1(
        n19379), .B2(n19921), .ZN(n19531) );
  OAI211_X1 U21643 ( .C1(n19533), .C2(n19782), .A(n19532), .B(n19531), .ZN(
        P2_U3079) );
  NOR2_X1 U21644 ( .A1(n19534), .A2(n19546), .ZN(n19927) );
  OAI21_X1 U21645 ( .B1(n11621), .B2(n19927), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19536) );
  OR2_X1 U21646 ( .A1(n19535), .A2(n19546), .ZN(n19540) );
  NAND2_X1 U21647 ( .A1(n19536), .A2(n19540), .ZN(n19928) );
  AOI22_X1 U21648 ( .A1(n19928), .A2(n19379), .B1(n19562), .B2(n19927), .ZN(
        n19545) );
  INV_X1 U21649 ( .A(n11621), .ZN(n19537) );
  AOI21_X1 U21650 ( .B1(n19537), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19543) );
  OAI21_X1 U21651 ( .B1(n19929), .B2(n19936), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19541) );
  NAND3_X1 U21652 ( .A1(n19541), .A2(n19564), .A3(n19540), .ZN(n19542) );
  OAI211_X1 U21653 ( .C1(n19927), .C2(n19543), .A(n19542), .B(n19571), .ZN(
        n19930) );
  AOI22_X1 U21654 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19930), .B1(
        n19936), .B2(n19563), .ZN(n19544) );
  OAI211_X1 U21655 ( .C1(n19578), .C2(n19782), .A(n19545), .B(n19544), .ZN(
        P2_U3071) );
  OR2_X1 U21656 ( .A1(n19546), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19561) );
  NOR2_X1 U21657 ( .A1(n19547), .A2(n19546), .ZN(n19934) );
  OAI21_X1 U21658 ( .B1(n19550), .B2(n19934), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19548) );
  OAI21_X1 U21659 ( .B1(n19561), .B2(n19549), .A(n19548), .ZN(n19935) );
  AOI22_X1 U21660 ( .A1(n19935), .A2(n19379), .B1(n19562), .B2(n19934), .ZN(
        n19560) );
  INV_X1 U21661 ( .A(n19934), .ZN(n19552) );
  NOR2_X1 U21662 ( .A1(n19934), .A2(n19550), .ZN(n19551) );
  AOI211_X1 U21663 ( .C1(n19553), .C2(n19552), .A(n19837), .B(n19551), .ZN(
        n19556) );
  OAI21_X1 U21664 ( .B1(n19558), .B2(n19554), .A(n19561), .ZN(n19555) );
  OAI21_X1 U21665 ( .B1(n19556), .B2(n19567), .A(n19555), .ZN(n19937) );
  AOI22_X1 U21666 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19937), .B1(
        n19943), .B2(n19563), .ZN(n19559) );
  OAI211_X1 U21667 ( .C1(n19578), .C2(n19933), .A(n19560), .B(n19559), .ZN(
        P2_U3063) );
  NOR2_X1 U21668 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19561), .ZN(
        n19942) );
  AOI22_X1 U21669 ( .A1(n19563), .A2(n19845), .B1(n19562), .B2(n19942), .ZN(
        n19577) );
  NAND3_X1 U21670 ( .A1(n19940), .A2(n19564), .A3(n19950), .ZN(n19566) );
  NAND2_X1 U21671 ( .A1(n19566), .A2(n19565), .ZN(n19573) );
  AOI21_X1 U21672 ( .B1(n11517), .B2(n19568), .A(n19567), .ZN(n19569) );
  AOI21_X1 U21673 ( .B1(n19573), .B2(n19570), .A(n19569), .ZN(n19572) );
  OAI21_X1 U21674 ( .B1(n19840), .B2(n19942), .A(n19573), .ZN(n19575) );
  OAI21_X1 U21675 ( .B1(n11517), .B2(n19942), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19574) );
  NAND2_X1 U21676 ( .A1(n19575), .A2(n19574), .ZN(n19946) );
  AOI22_X1 U21677 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19947), .B1(
        n19379), .B2(n19946), .ZN(n19576) );
  OAI211_X1 U21678 ( .C1(n19578), .C2(n19940), .A(n19577), .B(n19576), .ZN(
        P2_U3055) );
  AOI22_X1 U21679 ( .A1(n19581), .A2(n19580), .B1(n19579), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n19590) );
  AOI22_X1 U21680 ( .A1(n19583), .A2(BUF2_REG_22__SCAN_IN), .B1(n19582), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n19589) );
  AOI22_X1 U21681 ( .A1(n19587), .A2(n19586), .B1(n19585), .B2(n19584), .ZN(
        n19588) );
  NAND3_X1 U21682 ( .A1(n19590), .A2(n19589), .A3(n19588), .ZN(P2_U2897) );
  AOI22_X1 U21683 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19842), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n19843), .ZN(n19630) );
  NOR2_X2 U21684 ( .A1(n19591), .A2(n19837), .ZN(n19627) );
  NOR2_X2 U21685 ( .A1(n19592), .A2(n19839), .ZN(n19625) );
  AOI22_X1 U21686 ( .A1(n19841), .A2(n19627), .B1(n19840), .B2(n19625), .ZN(
        n19594) );
  AOI22_X1 U21687 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19843), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19842), .ZN(n19622) );
  AOI22_X1 U21688 ( .A1(n19626), .A2(n19845), .B1(
        P2_INSTQUEUE_REG_15__6__SCAN_IN), .B2(n19844), .ZN(n19593) );
  OAI211_X1 U21689 ( .C1(n19630), .C2(n19854), .A(n19594), .B(n19593), .ZN(
        P2_U3174) );
  AOI22_X1 U21690 ( .A1(n19626), .A2(n19796), .B1(n19625), .B2(n19848), .ZN(
        n19596) );
  AOI22_X1 U21691 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19851), .B1(
        n19627), .B2(n19850), .ZN(n19595) );
  OAI211_X1 U21692 ( .C1(n19630), .C2(n19860), .A(n19596), .B(n19595), .ZN(
        P2_U3166) );
  AOI22_X1 U21693 ( .A1(n19856), .A2(n19627), .B1(n19625), .B2(n19855), .ZN(
        n19598) );
  INV_X1 U21694 ( .A(n19630), .ZN(n19619) );
  AOI22_X1 U21695 ( .A1(n19619), .A2(n19863), .B1(
        P2_INSTQUEUE_REG_13__6__SCAN_IN), .B2(n19857), .ZN(n19597) );
  OAI211_X1 U21696 ( .C1(n19622), .C2(n19860), .A(n19598), .B(n19597), .ZN(
        P2_U3158) );
  AOI22_X1 U21697 ( .A1(n19862), .A2(n19627), .B1(n19625), .B2(n19861), .ZN(
        n19600) );
  AOI22_X1 U21698 ( .A1(n19864), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n19863), .B2(n19626), .ZN(n19599) );
  OAI211_X1 U21699 ( .C1(n19630), .C2(n19873), .A(n19600), .B(n19599), .ZN(
        P2_U3150) );
  AOI22_X1 U21700 ( .A1(n19868), .A2(n19627), .B1(n19625), .B2(n19867), .ZN(
        n19602) );
  AOI22_X1 U21701 ( .A1(n19626), .A2(n19803), .B1(
        P2_INSTQUEUE_REG_11__6__SCAN_IN), .B2(n19869), .ZN(n19601) );
  OAI211_X1 U21702 ( .C1(n19630), .C2(n19879), .A(n19602), .B(n19601), .ZN(
        P2_U3142) );
  AOI22_X1 U21703 ( .A1(n19619), .A2(n19881), .B1(n19625), .B2(n19874), .ZN(
        n19604) );
  AOI22_X1 U21704 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19876), .B1(
        n19627), .B2(n19875), .ZN(n19603) );
  OAI211_X1 U21705 ( .C1(n19622), .C2(n19879), .A(n19604), .B(n19603), .ZN(
        P2_U3134) );
  INV_X1 U21706 ( .A(n19886), .ZN(n19888) );
  AOI22_X1 U21707 ( .A1(n19619), .A2(n19888), .B1(n19625), .B2(n19880), .ZN(
        n19606) );
  AOI22_X1 U21708 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19883), .B1(
        n19627), .B2(n19882), .ZN(n19605) );
  OAI211_X1 U21709 ( .C1(n19622), .C2(n19808), .A(n19606), .B(n19605), .ZN(
        P2_U3126) );
  AOI22_X1 U21710 ( .A1(n19619), .A2(n19813), .B1(n19887), .B2(n19625), .ZN(
        n19608) );
  AOI22_X1 U21711 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19890), .B1(
        n19889), .B2(n19627), .ZN(n19607) );
  OAI211_X1 U21712 ( .C1(n19622), .C2(n19886), .A(n19608), .B(n19607), .ZN(
        P2_U3118) );
  AOI22_X1 U21713 ( .A1(n19894), .A2(n19627), .B1(n19893), .B2(n19625), .ZN(
        n19610) );
  INV_X1 U21714 ( .A(n19905), .ZN(n19895) );
  AOI22_X1 U21715 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19896), .B1(
        n19895), .B2(n19619), .ZN(n19609) );
  OAI211_X1 U21716 ( .C1(n19622), .C2(n19899), .A(n19610), .B(n19609), .ZN(
        P2_U3110) );
  AOI22_X1 U21717 ( .A1(n19901), .A2(n19627), .B1(n19625), .B2(n19900), .ZN(
        n19612) );
  AOI22_X1 U21718 ( .A1(n19619), .A2(n19907), .B1(
        P2_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n19902), .ZN(n19611) );
  OAI211_X1 U21719 ( .C1(n19622), .C2(n19905), .A(n19612), .B(n19611), .ZN(
        P2_U3102) );
  AOI22_X1 U21720 ( .A1(n19626), .A2(n19907), .B1(n19625), .B2(n19906), .ZN(
        n19614) );
  AOI22_X1 U21721 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19909), .B1(
        n19627), .B2(n19908), .ZN(n19613) );
  OAI211_X1 U21722 ( .C1(n19630), .C2(n19912), .A(n19614), .B(n19613), .ZN(
        P2_U3094) );
  AOI22_X1 U21723 ( .A1(n19626), .A2(n19914), .B1(n19913), .B2(n19625), .ZN(
        n19616) );
  AOI22_X1 U21724 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19916), .B1(
        n19627), .B2(n19915), .ZN(n19615) );
  OAI211_X1 U21725 ( .C1(n19630), .C2(n19925), .A(n19616), .B(n19615), .ZN(
        P2_U3086) );
  AOI22_X1 U21726 ( .A1(n19626), .A2(n19658), .B1(n19625), .B2(n19919), .ZN(
        n19618) );
  AOI22_X1 U21727 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19922), .B1(
        n19627), .B2(n19921), .ZN(n19617) );
  OAI211_X1 U21728 ( .C1(n19630), .C2(n19782), .A(n19618), .B(n19617), .ZN(
        P2_U3078) );
  AOI22_X1 U21729 ( .A1(n19928), .A2(n19627), .B1(n19625), .B2(n19927), .ZN(
        n19621) );
  AOI22_X1 U21730 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19930), .B1(
        n19936), .B2(n19619), .ZN(n19620) );
  OAI211_X1 U21731 ( .C1(n19622), .C2(n19782), .A(n19621), .B(n19620), .ZN(
        P2_U3070) );
  AOI22_X1 U21732 ( .A1(n19935), .A2(n19627), .B1(n19625), .B2(n19934), .ZN(
        n19624) );
  AOI22_X1 U21733 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19937), .B1(
        n19936), .B2(n19626), .ZN(n19623) );
  OAI211_X1 U21734 ( .C1(n19630), .C2(n19940), .A(n19624), .B(n19623), .ZN(
        P2_U3062) );
  AOI22_X1 U21735 ( .A1(n19626), .A2(n19943), .B1(n19625), .B2(n19942), .ZN(
        n19629) );
  AOI22_X1 U21736 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19947), .B1(
        n19946), .B2(n19627), .ZN(n19628) );
  OAI211_X1 U21737 ( .C1(n19630), .C2(n19950), .A(n19629), .B(n19628), .ZN(
        P2_U3054) );
  AOI22_X1 U21738 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19843), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19842), .ZN(n19671) );
  NOR2_X2 U21739 ( .A1(n19633), .A2(n19839), .ZN(n19667) );
  AOI22_X1 U21740 ( .A1(n19841), .A2(n19632), .B1(n19840), .B2(n19667), .ZN(
        n19635) );
  AOI22_X1 U21741 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19843), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19842), .ZN(n19666) );
  AOI22_X1 U21742 ( .A1(n19668), .A2(n19796), .B1(
        P2_INSTQUEUE_REG_15__5__SCAN_IN), .B2(n19844), .ZN(n19634) );
  OAI211_X1 U21743 ( .C1(n19671), .C2(n19950), .A(n19635), .B(n19634), .ZN(
        P2_U3173) );
  AOI22_X1 U21744 ( .A1(n19668), .A2(n19849), .B1(n19667), .B2(n19848), .ZN(
        n19637) );
  AOI22_X1 U21745 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19851), .B1(
        n19632), .B2(n19850), .ZN(n19636) );
  OAI211_X1 U21746 ( .C1(n19671), .C2(n19854), .A(n19637), .B(n19636), .ZN(
        P2_U3165) );
  AOI22_X1 U21747 ( .A1(n19856), .A2(n19632), .B1(n19667), .B2(n19855), .ZN(
        n19639) );
  AOI22_X1 U21748 ( .A1(n19668), .A2(n19863), .B1(
        P2_INSTQUEUE_REG_13__5__SCAN_IN), .B2(n19857), .ZN(n19638) );
  OAI211_X1 U21749 ( .C1(n19671), .C2(n19860), .A(n19639), .B(n19638), .ZN(
        P2_U3157) );
  AOI22_X1 U21750 ( .A1(n19862), .A2(n19632), .B1(n19667), .B2(n19861), .ZN(
        n19641) );
  INV_X1 U21751 ( .A(n19671), .ZN(n19663) );
  AOI22_X1 U21752 ( .A1(n19864), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n19863), .B2(n19663), .ZN(n19640) );
  OAI211_X1 U21753 ( .C1(n19666), .C2(n19873), .A(n19641), .B(n19640), .ZN(
        P2_U3149) );
  AOI22_X1 U21754 ( .A1(n19868), .A2(n19632), .B1(n19667), .B2(n19867), .ZN(
        n19643) );
  AOI22_X1 U21755 ( .A1(n19668), .A2(n19870), .B1(
        P2_INSTQUEUE_REG_11__5__SCAN_IN), .B2(n19869), .ZN(n19642) );
  OAI211_X1 U21756 ( .C1(n19671), .C2(n19873), .A(n19643), .B(n19642), .ZN(
        P2_U3141) );
  AOI22_X1 U21757 ( .A1(n19663), .A2(n19870), .B1(n19667), .B2(n19874), .ZN(
        n19645) );
  AOI22_X1 U21758 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19876), .B1(
        n19632), .B2(n19875), .ZN(n19644) );
  OAI211_X1 U21759 ( .C1(n19666), .C2(n19808), .A(n19645), .B(n19644), .ZN(
        P2_U3133) );
  AOI22_X1 U21760 ( .A1(n19663), .A2(n19881), .B1(n19667), .B2(n19880), .ZN(
        n19647) );
  AOI22_X1 U21761 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19883), .B1(
        n19632), .B2(n19882), .ZN(n19646) );
  OAI211_X1 U21762 ( .C1(n19666), .C2(n19886), .A(n19647), .B(n19646), .ZN(
        P2_U3125) );
  AOI22_X1 U21763 ( .A1(n19668), .A2(n19813), .B1(n19887), .B2(n19667), .ZN(
        n19649) );
  AOI22_X1 U21764 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19890), .B1(
        n19889), .B2(n19632), .ZN(n19648) );
  OAI211_X1 U21765 ( .C1(n19671), .C2(n19886), .A(n19649), .B(n19648), .ZN(
        P2_U3117) );
  AOI22_X1 U21766 ( .A1(n19894), .A2(n19632), .B1(n19893), .B2(n19667), .ZN(
        n19651) );
  AOI22_X1 U21767 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19896), .B1(
        n19813), .B2(n19663), .ZN(n19650) );
  OAI211_X1 U21768 ( .C1(n19666), .C2(n19905), .A(n19651), .B(n19650), .ZN(
        P2_U3109) );
  AOI22_X1 U21769 ( .A1(n19901), .A2(n19632), .B1(n19667), .B2(n19900), .ZN(
        n19653) );
  AOI22_X1 U21770 ( .A1(n19668), .A2(n19907), .B1(
        P2_INSTQUEUE_REG_6__5__SCAN_IN), .B2(n19902), .ZN(n19652) );
  OAI211_X1 U21771 ( .C1(n19671), .C2(n19905), .A(n19653), .B(n19652), .ZN(
        P2_U3101) );
  AOI22_X1 U21772 ( .A1(n19668), .A2(n19914), .B1(n19667), .B2(n19906), .ZN(
        n19655) );
  AOI22_X1 U21773 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19909), .B1(
        n19632), .B2(n19908), .ZN(n19654) );
  OAI211_X1 U21774 ( .C1(n19671), .C2(n19818), .A(n19655), .B(n19654), .ZN(
        P2_U3093) );
  AOI22_X1 U21775 ( .A1(n19663), .A2(n19914), .B1(n19913), .B2(n19667), .ZN(
        n19657) );
  AOI22_X1 U21776 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19916), .B1(
        n19632), .B2(n19915), .ZN(n19656) );
  OAI211_X1 U21777 ( .C1(n19666), .C2(n19925), .A(n19657), .B(n19656), .ZN(
        P2_U3085) );
  AOI22_X1 U21778 ( .A1(n19663), .A2(n19658), .B1(n19667), .B2(n19919), .ZN(
        n19660) );
  AOI22_X1 U21779 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19922), .B1(
        n19632), .B2(n19921), .ZN(n19659) );
  OAI211_X1 U21780 ( .C1(n19666), .C2(n19782), .A(n19660), .B(n19659), .ZN(
        P2_U3077) );
  AOI22_X1 U21781 ( .A1(n19928), .A2(n19632), .B1(n19667), .B2(n19927), .ZN(
        n19662) );
  AOI22_X1 U21782 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19930), .B1(
        n19936), .B2(n19668), .ZN(n19661) );
  OAI211_X1 U21783 ( .C1(n19671), .C2(n19782), .A(n19662), .B(n19661), .ZN(
        P2_U3069) );
  AOI22_X1 U21784 ( .A1(n19935), .A2(n19632), .B1(n19667), .B2(n19934), .ZN(
        n19665) );
  AOI22_X1 U21785 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19937), .B1(
        n19936), .B2(n19663), .ZN(n19664) );
  OAI211_X1 U21786 ( .C1(n19666), .C2(n19940), .A(n19665), .B(n19664), .ZN(
        P2_U3061) );
  AOI22_X1 U21787 ( .A1(n19668), .A2(n19845), .B1(n19667), .B2(n19942), .ZN(
        n19670) );
  AOI22_X1 U21788 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19947), .B1(
        n19946), .B2(n19632), .ZN(n19669) );
  OAI211_X1 U21789 ( .C1(n19671), .C2(n19940), .A(n19670), .B(n19669), .ZN(
        P2_U3053) );
  AOI22_X1 U21790 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19842), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19843), .ZN(n19706) );
  NOR2_X2 U21791 ( .A1(n19674), .A2(n19839), .ZN(n19707) );
  AOI22_X1 U21792 ( .A1(n19841), .A2(n19673), .B1(n19840), .B2(n19707), .ZN(
        n19676) );
  AOI22_X1 U21793 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19843), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19842), .ZN(n19711) );
  INV_X1 U21794 ( .A(n19711), .ZN(n19703) );
  AOI22_X1 U21795 ( .A1(n19703), .A2(n19845), .B1(
        P2_INSTQUEUE_REG_15__4__SCAN_IN), .B2(n19844), .ZN(n19675) );
  OAI211_X1 U21796 ( .C1(n19706), .C2(n19854), .A(n19676), .B(n19675), .ZN(
        P2_U3172) );
  AOI22_X1 U21797 ( .A1(n19703), .A2(n19796), .B1(n19848), .B2(n19707), .ZN(
        n19678) );
  AOI22_X1 U21798 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19851), .B1(
        n19673), .B2(n19850), .ZN(n19677) );
  OAI211_X1 U21799 ( .C1(n19706), .C2(n19860), .A(n19678), .B(n19677), .ZN(
        P2_U3164) );
  AOI22_X1 U21800 ( .A1(n19856), .A2(n19673), .B1(n19707), .B2(n19855), .ZN(
        n19680) );
  AOI22_X1 U21801 ( .A1(n19708), .A2(n19863), .B1(
        P2_INSTQUEUE_REG_13__4__SCAN_IN), .B2(n19857), .ZN(n19679) );
  OAI211_X1 U21802 ( .C1(n19711), .C2(n19860), .A(n19680), .B(n19679), .ZN(
        P2_U3156) );
  AOI22_X1 U21803 ( .A1(n19862), .A2(n19673), .B1(n19707), .B2(n19861), .ZN(
        n19682) );
  AOI22_X1 U21804 ( .A1(n19864), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n19863), .B2(n19703), .ZN(n19681) );
  OAI211_X1 U21805 ( .C1(n19706), .C2(n19873), .A(n19682), .B(n19681), .ZN(
        P2_U3148) );
  AOI22_X1 U21806 ( .A1(n19868), .A2(n19673), .B1(n19707), .B2(n19867), .ZN(
        n19684) );
  AOI22_X1 U21807 ( .A1(n19708), .A2(n19870), .B1(
        P2_INSTQUEUE_REG_11__4__SCAN_IN), .B2(n19869), .ZN(n19683) );
  OAI211_X1 U21808 ( .C1(n19711), .C2(n19873), .A(n19684), .B(n19683), .ZN(
        P2_U3140) );
  AOI22_X1 U21809 ( .A1(n19708), .A2(n19881), .B1(n19707), .B2(n19874), .ZN(
        n19686) );
  AOI22_X1 U21810 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19876), .B1(
        n19673), .B2(n19875), .ZN(n19685) );
  OAI211_X1 U21811 ( .C1(n19711), .C2(n19879), .A(n19686), .B(n19685), .ZN(
        P2_U3132) );
  AOI22_X1 U21812 ( .A1(n19708), .A2(n19888), .B1(n19707), .B2(n19880), .ZN(
        n19688) );
  AOI22_X1 U21813 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19883), .B1(
        n19673), .B2(n19882), .ZN(n19687) );
  OAI211_X1 U21814 ( .C1(n19711), .C2(n19808), .A(n19688), .B(n19687), .ZN(
        P2_U3124) );
  AOI22_X1 U21815 ( .A1(n19703), .A2(n19888), .B1(n19887), .B2(n19707), .ZN(
        n19690) );
  AOI22_X1 U21816 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19890), .B1(
        n19889), .B2(n19673), .ZN(n19689) );
  OAI211_X1 U21817 ( .C1(n19706), .C2(n19899), .A(n19690), .B(n19689), .ZN(
        P2_U3116) );
  AOI22_X1 U21818 ( .A1(n19894), .A2(n19673), .B1(n19893), .B2(n19707), .ZN(
        n19692) );
  AOI22_X1 U21819 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19896), .B1(
        n19813), .B2(n19703), .ZN(n19691) );
  OAI211_X1 U21820 ( .C1(n19706), .C2(n19905), .A(n19692), .B(n19691), .ZN(
        P2_U3108) );
  AOI22_X1 U21821 ( .A1(n19901), .A2(n19673), .B1(n19707), .B2(n19900), .ZN(
        n19694) );
  AOI22_X1 U21822 ( .A1(n19708), .A2(n19907), .B1(
        P2_INSTQUEUE_REG_6__4__SCAN_IN), .B2(n19902), .ZN(n19693) );
  OAI211_X1 U21823 ( .C1(n19711), .C2(n19905), .A(n19694), .B(n19693), .ZN(
        P2_U3100) );
  AOI22_X1 U21824 ( .A1(n19708), .A2(n19914), .B1(n19707), .B2(n19906), .ZN(
        n19696) );
  AOI22_X1 U21825 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19909), .B1(
        n19673), .B2(n19908), .ZN(n19695) );
  OAI211_X1 U21826 ( .C1(n19711), .C2(n19818), .A(n19696), .B(n19695), .ZN(
        P2_U3092) );
  AOI22_X1 U21827 ( .A1(n19703), .A2(n19914), .B1(n19913), .B2(n19707), .ZN(
        n19698) );
  AOI22_X1 U21828 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19916), .B1(
        n19673), .B2(n19915), .ZN(n19697) );
  OAI211_X1 U21829 ( .C1(n19706), .C2(n19925), .A(n19698), .B(n19697), .ZN(
        P2_U3084) );
  AOI22_X1 U21830 ( .A1(n19708), .A2(n19929), .B1(n19707), .B2(n19919), .ZN(
        n19700) );
  AOI22_X1 U21831 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19922), .B1(
        n19673), .B2(n19921), .ZN(n19699) );
  OAI211_X1 U21832 ( .C1(n19711), .C2(n19925), .A(n19700), .B(n19699), .ZN(
        P2_U3076) );
  AOI22_X1 U21833 ( .A1(n19928), .A2(n19673), .B1(n19707), .B2(n19927), .ZN(
        n19702) );
  AOI22_X1 U21834 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19930), .B1(
        n19936), .B2(n19708), .ZN(n19701) );
  OAI211_X1 U21835 ( .C1(n19711), .C2(n19782), .A(n19702), .B(n19701), .ZN(
        P2_U3068) );
  AOI22_X1 U21836 ( .A1(n19935), .A2(n19673), .B1(n19707), .B2(n19934), .ZN(
        n19705) );
  AOI22_X1 U21837 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19937), .B1(
        n19936), .B2(n19703), .ZN(n19704) );
  OAI211_X1 U21838 ( .C1(n19706), .C2(n19940), .A(n19705), .B(n19704), .ZN(
        P2_U3060) );
  AOI22_X1 U21839 ( .A1(n19708), .A2(n19845), .B1(n19942), .B2(n19707), .ZN(
        n19710) );
  AOI22_X1 U21840 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19947), .B1(
        n19946), .B2(n19673), .ZN(n19709) );
  OAI211_X1 U21841 ( .C1(n19711), .C2(n19940), .A(n19710), .B(n19709), .ZN(
        P2_U3052) );
  AOI22_X1 U21842 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19843), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19842), .ZN(n19750) );
  NOR2_X2 U21843 ( .A1(n11377), .A2(n19839), .ZN(n19746) );
  AOI22_X1 U21844 ( .A1(n19841), .A2(n19713), .B1(n19840), .B2(n19746), .ZN(
        n19715) );
  AOI22_X1 U21845 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19843), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19842), .ZN(n19745) );
  INV_X1 U21846 ( .A(n19745), .ZN(n19747) );
  AOI22_X1 U21847 ( .A1(n19747), .A2(n19845), .B1(
        P2_INSTQUEUE_REG_15__3__SCAN_IN), .B2(n19844), .ZN(n19714) );
  OAI211_X1 U21848 ( .C1(n19750), .C2(n19854), .A(n19715), .B(n19714), .ZN(
        P2_U3171) );
  AOI22_X1 U21849 ( .A1(n19747), .A2(n19796), .B1(n19746), .B2(n19848), .ZN(
        n19717) );
  AOI22_X1 U21850 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19851), .B1(
        n19713), .B2(n19850), .ZN(n19716) );
  OAI211_X1 U21851 ( .C1(n19750), .C2(n19860), .A(n19717), .B(n19716), .ZN(
        P2_U3163) );
  AOI22_X1 U21852 ( .A1(n19856), .A2(n19713), .B1(n19746), .B2(n19855), .ZN(
        n19719) );
  AOI22_X1 U21853 ( .A1(n19742), .A2(n19863), .B1(
        P2_INSTQUEUE_REG_13__3__SCAN_IN), .B2(n19857), .ZN(n19718) );
  OAI211_X1 U21854 ( .C1(n19745), .C2(n19860), .A(n19719), .B(n19718), .ZN(
        P2_U3155) );
  AOI22_X1 U21855 ( .A1(n19862), .A2(n19713), .B1(n19746), .B2(n19861), .ZN(
        n19721) );
  AOI22_X1 U21856 ( .A1(n19864), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n19863), .B2(n19747), .ZN(n19720) );
  OAI211_X1 U21857 ( .C1(n19750), .C2(n19873), .A(n19721), .B(n19720), .ZN(
        P2_U3147) );
  AOI22_X1 U21858 ( .A1(n19868), .A2(n19713), .B1(n19746), .B2(n19867), .ZN(
        n19723) );
  AOI22_X1 U21859 ( .A1(n19742), .A2(n19870), .B1(
        P2_INSTQUEUE_REG_11__3__SCAN_IN), .B2(n19869), .ZN(n19722) );
  OAI211_X1 U21860 ( .C1(n19745), .C2(n19873), .A(n19723), .B(n19722), .ZN(
        P2_U3139) );
  AOI22_X1 U21861 ( .A1(n19742), .A2(n19881), .B1(n19746), .B2(n19874), .ZN(
        n19725) );
  AOI22_X1 U21862 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19876), .B1(
        n19713), .B2(n19875), .ZN(n19724) );
  OAI211_X1 U21863 ( .C1(n19745), .C2(n19879), .A(n19725), .B(n19724), .ZN(
        P2_U3131) );
  AOI22_X1 U21864 ( .A1(n19747), .A2(n19881), .B1(n19746), .B2(n19880), .ZN(
        n19727) );
  AOI22_X1 U21865 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19883), .B1(
        n19713), .B2(n19882), .ZN(n19726) );
  OAI211_X1 U21866 ( .C1(n19750), .C2(n19886), .A(n19727), .B(n19726), .ZN(
        P2_U3123) );
  AOI22_X1 U21867 ( .A1(n19742), .A2(n19813), .B1(n19887), .B2(n19746), .ZN(
        n19729) );
  AOI22_X1 U21868 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19890), .B1(
        n19889), .B2(n19713), .ZN(n19728) );
  OAI211_X1 U21869 ( .C1(n19745), .C2(n19886), .A(n19729), .B(n19728), .ZN(
        P2_U3115) );
  AOI22_X1 U21870 ( .A1(n19894), .A2(n19713), .B1(n19893), .B2(n19746), .ZN(
        n19731) );
  AOI22_X1 U21871 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19896), .B1(
        n19895), .B2(n19742), .ZN(n19730) );
  OAI211_X1 U21872 ( .C1(n19745), .C2(n19899), .A(n19731), .B(n19730), .ZN(
        P2_U3107) );
  AOI22_X1 U21873 ( .A1(n19901), .A2(n19713), .B1(n19746), .B2(n19900), .ZN(
        n19733) );
  AOI22_X1 U21874 ( .A1(n19742), .A2(n19907), .B1(
        P2_INSTQUEUE_REG_6__3__SCAN_IN), .B2(n19902), .ZN(n19732) );
  OAI211_X1 U21875 ( .C1(n19745), .C2(n19905), .A(n19733), .B(n19732), .ZN(
        P2_U3099) );
  AOI22_X1 U21876 ( .A1(n19742), .A2(n19914), .B1(n19746), .B2(n19906), .ZN(
        n19735) );
  AOI22_X1 U21877 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19909), .B1(
        n19713), .B2(n19908), .ZN(n19734) );
  OAI211_X1 U21878 ( .C1(n19745), .C2(n19818), .A(n19735), .B(n19734), .ZN(
        P2_U3091) );
  AOI22_X1 U21879 ( .A1(n19747), .A2(n19914), .B1(n19913), .B2(n19746), .ZN(
        n19737) );
  AOI22_X1 U21880 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19916), .B1(
        n19713), .B2(n19915), .ZN(n19736) );
  OAI211_X1 U21881 ( .C1(n19750), .C2(n19925), .A(n19737), .B(n19736), .ZN(
        P2_U3083) );
  AOI22_X1 U21882 ( .A1(n19742), .A2(n19929), .B1(n19746), .B2(n19919), .ZN(
        n19739) );
  AOI22_X1 U21883 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19922), .B1(
        n19713), .B2(n19921), .ZN(n19738) );
  OAI211_X1 U21884 ( .C1(n19745), .C2(n19925), .A(n19739), .B(n19738), .ZN(
        P2_U3075) );
  AOI22_X1 U21885 ( .A1(n19928), .A2(n19713), .B1(n19746), .B2(n19927), .ZN(
        n19741) );
  AOI22_X1 U21886 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19930), .B1(
        n19936), .B2(n19742), .ZN(n19740) );
  OAI211_X1 U21887 ( .C1(n19745), .C2(n19782), .A(n19741), .B(n19740), .ZN(
        P2_U3067) );
  AOI22_X1 U21888 ( .A1(n19935), .A2(n19713), .B1(n19746), .B2(n19934), .ZN(
        n19744) );
  AOI22_X1 U21889 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19937), .B1(
        n19943), .B2(n19742), .ZN(n19743) );
  OAI211_X1 U21890 ( .C1(n19745), .C2(n19933), .A(n19744), .B(n19743), .ZN(
        P2_U3059) );
  AOI22_X1 U21891 ( .A1(n19747), .A2(n19943), .B1(n19746), .B2(n19942), .ZN(
        n19749) );
  AOI22_X1 U21892 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19947), .B1(
        n19946), .B2(n19713), .ZN(n19748) );
  OAI211_X1 U21893 ( .C1(n19750), .C2(n19950), .A(n19749), .B(n19748), .ZN(
        P2_U3051) );
  AOI22_X1 U21894 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19843), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19842), .ZN(n19786) );
  NOR2_X2 U21895 ( .A1(n19753), .A2(n19839), .ZN(n19787) );
  AOI22_X1 U21896 ( .A1(n19841), .A2(n19752), .B1(n19840), .B2(n19787), .ZN(
        n19755) );
  AOI22_X1 U21897 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19843), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19842), .ZN(n19791) );
  AOI22_X1 U21898 ( .A1(n19783), .A2(n19796), .B1(
        P2_INSTQUEUE_REG_15__2__SCAN_IN), .B2(n19844), .ZN(n19754) );
  OAI211_X1 U21899 ( .C1(n19786), .C2(n19950), .A(n19755), .B(n19754), .ZN(
        P2_U3170) );
  AOI22_X1 U21900 ( .A1(n19783), .A2(n19849), .B1(n19787), .B2(n19848), .ZN(
        n19757) );
  AOI22_X1 U21901 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19851), .B1(
        n19752), .B2(n19850), .ZN(n19756) );
  OAI211_X1 U21902 ( .C1(n19786), .C2(n19854), .A(n19757), .B(n19756), .ZN(
        P2_U3162) );
  AOI22_X1 U21903 ( .A1(n19856), .A2(n19752), .B1(n19787), .B2(n19855), .ZN(
        n19759) );
  AOI22_X1 U21904 ( .A1(n19783), .A2(n19863), .B1(
        P2_INSTQUEUE_REG_13__2__SCAN_IN), .B2(n19857), .ZN(n19758) );
  OAI211_X1 U21905 ( .C1(n19786), .C2(n19860), .A(n19759), .B(n19758), .ZN(
        P2_U3154) );
  AOI22_X1 U21906 ( .A1(n19862), .A2(n19752), .B1(n19787), .B2(n19861), .ZN(
        n19761) );
  INV_X1 U21907 ( .A(n19786), .ZN(n19788) );
  AOI22_X1 U21908 ( .A1(n19864), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n19863), .B2(n19788), .ZN(n19760) );
  OAI211_X1 U21909 ( .C1(n19791), .C2(n19873), .A(n19761), .B(n19760), .ZN(
        P2_U3146) );
  AOI22_X1 U21910 ( .A1(n19868), .A2(n19752), .B1(n19787), .B2(n19867), .ZN(
        n19763) );
  AOI22_X1 U21911 ( .A1(n19783), .A2(n19870), .B1(
        P2_INSTQUEUE_REG_11__2__SCAN_IN), .B2(n19869), .ZN(n19762) );
  OAI211_X1 U21912 ( .C1(n19786), .C2(n19873), .A(n19763), .B(n19762), .ZN(
        P2_U3138) );
  AOI22_X1 U21913 ( .A1(n19788), .A2(n19870), .B1(n19787), .B2(n19874), .ZN(
        n19765) );
  AOI22_X1 U21914 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19876), .B1(
        n19752), .B2(n19875), .ZN(n19764) );
  OAI211_X1 U21915 ( .C1(n19791), .C2(n19808), .A(n19765), .B(n19764), .ZN(
        P2_U3130) );
  AOI22_X1 U21916 ( .A1(n19788), .A2(n19881), .B1(n19787), .B2(n19880), .ZN(
        n19767) );
  AOI22_X1 U21917 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19883), .B1(
        n19752), .B2(n19882), .ZN(n19766) );
  OAI211_X1 U21918 ( .C1(n19791), .C2(n19886), .A(n19767), .B(n19766), .ZN(
        P2_U3122) );
  AOI22_X1 U21919 ( .A1(n19783), .A2(n19813), .B1(n19887), .B2(n19787), .ZN(
        n19769) );
  AOI22_X1 U21920 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19890), .B1(
        n19889), .B2(n19752), .ZN(n19768) );
  OAI211_X1 U21921 ( .C1(n19786), .C2(n19886), .A(n19769), .B(n19768), .ZN(
        P2_U3114) );
  AOI22_X1 U21922 ( .A1(n19894), .A2(n19752), .B1(n19893), .B2(n19787), .ZN(
        n19771) );
  AOI22_X1 U21923 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19896), .B1(
        n19813), .B2(n19788), .ZN(n19770) );
  OAI211_X1 U21924 ( .C1(n19791), .C2(n19905), .A(n19771), .B(n19770), .ZN(
        P2_U3106) );
  AOI22_X1 U21925 ( .A1(n19901), .A2(n19752), .B1(n19787), .B2(n19900), .ZN(
        n19773) );
  AOI22_X1 U21926 ( .A1(n19783), .A2(n19907), .B1(
        P2_INSTQUEUE_REG_6__2__SCAN_IN), .B2(n19902), .ZN(n19772) );
  OAI211_X1 U21927 ( .C1(n19786), .C2(n19905), .A(n19773), .B(n19772), .ZN(
        P2_U3098) );
  AOI22_X1 U21928 ( .A1(n19783), .A2(n19914), .B1(n19787), .B2(n19906), .ZN(
        n19775) );
  AOI22_X1 U21929 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19909), .B1(
        n19752), .B2(n19908), .ZN(n19774) );
  OAI211_X1 U21930 ( .C1(n19786), .C2(n19818), .A(n19775), .B(n19774), .ZN(
        P2_U3090) );
  AOI22_X1 U21931 ( .A1(n19788), .A2(n19914), .B1(n19913), .B2(n19787), .ZN(
        n19777) );
  AOI22_X1 U21932 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19916), .B1(
        n19752), .B2(n19915), .ZN(n19776) );
  OAI211_X1 U21933 ( .C1(n19791), .C2(n19925), .A(n19777), .B(n19776), .ZN(
        P2_U3082) );
  AOI22_X1 U21934 ( .A1(n19783), .A2(n19929), .B1(n19787), .B2(n19919), .ZN(
        n19779) );
  AOI22_X1 U21935 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19922), .B1(
        n19752), .B2(n19921), .ZN(n19778) );
  OAI211_X1 U21936 ( .C1(n19786), .C2(n19925), .A(n19779), .B(n19778), .ZN(
        P2_U3074) );
  AOI22_X1 U21937 ( .A1(n19928), .A2(n19752), .B1(n19787), .B2(n19927), .ZN(
        n19781) );
  AOI22_X1 U21938 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19930), .B1(
        n19936), .B2(n19783), .ZN(n19780) );
  OAI211_X1 U21939 ( .C1(n19786), .C2(n19782), .A(n19781), .B(n19780), .ZN(
        P2_U3066) );
  AOI22_X1 U21940 ( .A1(n19935), .A2(n19752), .B1(n19787), .B2(n19934), .ZN(
        n19785) );
  AOI22_X1 U21941 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19937), .B1(
        n19943), .B2(n19783), .ZN(n19784) );
  OAI211_X1 U21942 ( .C1(n19786), .C2(n19933), .A(n19785), .B(n19784), .ZN(
        P2_U3058) );
  AOI22_X1 U21943 ( .A1(n19788), .A2(n19943), .B1(n19787), .B2(n19942), .ZN(
        n19790) );
  AOI22_X1 U21944 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19947), .B1(
        n19946), .B2(n19752), .ZN(n19789) );
  OAI211_X1 U21945 ( .C1(n19791), .C2(n19950), .A(n19790), .B(n19789), .ZN(
        P2_U3050) );
  AOI22_X2 U21946 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19842), .B1(
        BUF1_REG_25__SCAN_IN), .B2(n19843), .ZN(n19836) );
  NOR2_X2 U21947 ( .A1(n19792), .A2(n19837), .ZN(n19833) );
  NOR2_X2 U21948 ( .A1(n10959), .A2(n19839), .ZN(n19831) );
  AOI22_X1 U21949 ( .A1(n19841), .A2(n19833), .B1(n19840), .B2(n19831), .ZN(
        n19795) );
  AOI22_X1 U21950 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19843), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19842), .ZN(n19826) );
  AOI22_X1 U21951 ( .A1(n19832), .A2(n19845), .B1(
        P2_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n19844), .ZN(n19794) );
  OAI211_X1 U21952 ( .C1(n19836), .C2(n19854), .A(n19795), .B(n19794), .ZN(
        P2_U3169) );
  AOI22_X1 U21953 ( .A1(n19832), .A2(n19796), .B1(n19848), .B2(n19831), .ZN(
        n19798) );
  AOI22_X1 U21954 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19851), .B1(
        n19833), .B2(n19850), .ZN(n19797) );
  OAI211_X1 U21955 ( .C1(n19836), .C2(n19860), .A(n19798), .B(n19797), .ZN(
        P2_U3161) );
  AOI22_X1 U21956 ( .A1(n19856), .A2(n19833), .B1(n19831), .B2(n19855), .ZN(
        n19800) );
  INV_X1 U21957 ( .A(n19836), .ZN(n19823) );
  AOI22_X1 U21958 ( .A1(n19823), .A2(n19863), .B1(
        P2_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n19857), .ZN(n19799) );
  OAI211_X1 U21959 ( .C1(n19826), .C2(n19860), .A(n19800), .B(n19799), .ZN(
        P2_U3153) );
  AOI22_X1 U21960 ( .A1(n19862), .A2(n19833), .B1(n19831), .B2(n19861), .ZN(
        n19802) );
  AOI22_X1 U21961 ( .A1(n19864), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n19863), .B2(n19832), .ZN(n19801) );
  OAI211_X1 U21962 ( .C1(n19836), .C2(n19873), .A(n19802), .B(n19801), .ZN(
        P2_U3145) );
  AOI22_X1 U21963 ( .A1(n19868), .A2(n19833), .B1(n19831), .B2(n19867), .ZN(
        n19805) );
  AOI22_X1 U21964 ( .A1(n19832), .A2(n19803), .B1(
        P2_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n19869), .ZN(n19804) );
  OAI211_X1 U21965 ( .C1(n19836), .C2(n19879), .A(n19805), .B(n19804), .ZN(
        P2_U3137) );
  AOI22_X1 U21966 ( .A1(n19832), .A2(n19870), .B1(n19831), .B2(n19874), .ZN(
        n19807) );
  AOI22_X1 U21967 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19876), .B1(
        n19833), .B2(n19875), .ZN(n19806) );
  OAI211_X1 U21968 ( .C1(n19836), .C2(n19808), .A(n19807), .B(n19806), .ZN(
        P2_U3129) );
  AOI22_X1 U21969 ( .A1(n19832), .A2(n19881), .B1(n19831), .B2(n19880), .ZN(
        n19810) );
  AOI22_X1 U21970 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19883), .B1(
        n19833), .B2(n19882), .ZN(n19809) );
  OAI211_X1 U21971 ( .C1(n19836), .C2(n19886), .A(n19810), .B(n19809), .ZN(
        P2_U3121) );
  AOI22_X1 U21972 ( .A1(n19832), .A2(n19888), .B1(n19887), .B2(n19831), .ZN(
        n19812) );
  AOI22_X1 U21973 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19890), .B1(
        n19889), .B2(n19833), .ZN(n19811) );
  OAI211_X1 U21974 ( .C1(n19836), .C2(n19899), .A(n19812), .B(n19811), .ZN(
        P2_U3113) );
  AOI22_X1 U21975 ( .A1(n19894), .A2(n19833), .B1(n19893), .B2(n19831), .ZN(
        n19815) );
  AOI22_X1 U21976 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19896), .B1(
        n19813), .B2(n19832), .ZN(n19814) );
  OAI211_X1 U21977 ( .C1(n19836), .C2(n19905), .A(n19815), .B(n19814), .ZN(
        P2_U3105) );
  AOI22_X1 U21978 ( .A1(n19901), .A2(n19833), .B1(n19831), .B2(n19900), .ZN(
        n19817) );
  AOI22_X1 U21979 ( .A1(n19832), .A2(n19895), .B1(
        P2_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n19902), .ZN(n19816) );
  OAI211_X1 U21980 ( .C1(n19836), .C2(n19818), .A(n19817), .B(n19816), .ZN(
        P2_U3097) );
  AOI22_X1 U21981 ( .A1(n19832), .A2(n19907), .B1(n19831), .B2(n19906), .ZN(
        n19820) );
  AOI22_X1 U21982 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19909), .B1(
        n19833), .B2(n19908), .ZN(n19819) );
  OAI211_X1 U21983 ( .C1(n19836), .C2(n19912), .A(n19820), .B(n19819), .ZN(
        P2_U3089) );
  AOI22_X1 U21984 ( .A1(n19832), .A2(n19914), .B1(n19913), .B2(n19831), .ZN(
        n19822) );
  AOI22_X1 U21985 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19916), .B1(
        n19833), .B2(n19915), .ZN(n19821) );
  OAI211_X1 U21986 ( .C1(n19836), .C2(n19925), .A(n19822), .B(n19821), .ZN(
        P2_U3081) );
  AOI22_X1 U21987 ( .A1(n19823), .A2(n19929), .B1(n19831), .B2(n19919), .ZN(
        n19825) );
  AOI22_X1 U21988 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19922), .B1(
        n19833), .B2(n19921), .ZN(n19824) );
  OAI211_X1 U21989 ( .C1(n19826), .C2(n19925), .A(n19825), .B(n19824), .ZN(
        P2_U3073) );
  AOI22_X1 U21990 ( .A1(n19928), .A2(n19833), .B1(n19831), .B2(n19927), .ZN(
        n19828) );
  AOI22_X1 U21991 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19930), .B1(
        n19929), .B2(n19832), .ZN(n19827) );
  OAI211_X1 U21992 ( .C1(n19836), .C2(n19933), .A(n19828), .B(n19827), .ZN(
        P2_U3065) );
  AOI22_X1 U21993 ( .A1(n19935), .A2(n19833), .B1(n19831), .B2(n19934), .ZN(
        n19830) );
  AOI22_X1 U21994 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19937), .B1(
        n19936), .B2(n19832), .ZN(n19829) );
  OAI211_X1 U21995 ( .C1(n19836), .C2(n19940), .A(n19830), .B(n19829), .ZN(
        P2_U3057) );
  AOI22_X1 U21996 ( .A1(n19832), .A2(n19943), .B1(n19942), .B2(n19831), .ZN(
        n19835) );
  AOI22_X1 U21997 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19947), .B1(
        n19946), .B2(n19833), .ZN(n19834) );
  OAI211_X1 U21998 ( .C1(n19836), .C2(n19950), .A(n19835), .B(n19834), .ZN(
        P2_U3049) );
  AOI22_X1 U21999 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19843), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19842), .ZN(n19951) );
  NOR2_X2 U22000 ( .A1(n19838), .A2(n19837), .ZN(n19945) );
  NOR2_X2 U22001 ( .A1(n11411), .A2(n19839), .ZN(n19941) );
  AOI22_X1 U22002 ( .A1(n19841), .A2(n19945), .B1(n19840), .B2(n19941), .ZN(
        n19847) );
  AOI22_X1 U22003 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19843), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19842), .ZN(n19926) );
  AOI22_X1 U22004 ( .A1(n19944), .A2(n19845), .B1(
        P2_INSTQUEUE_REG_15__0__SCAN_IN), .B2(n19844), .ZN(n19846) );
  OAI211_X1 U22005 ( .C1(n19951), .C2(n19854), .A(n19847), .B(n19846), .ZN(
        P2_U3168) );
  INV_X1 U22006 ( .A(n19951), .ZN(n19920) );
  AOI22_X1 U22007 ( .A1(n19920), .A2(n19849), .B1(n19848), .B2(n19941), .ZN(
        n19853) );
  AOI22_X1 U22008 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19851), .B1(
        n19945), .B2(n19850), .ZN(n19852) );
  OAI211_X1 U22009 ( .C1(n19926), .C2(n19854), .A(n19853), .B(n19852), .ZN(
        P2_U3160) );
  AOI22_X1 U22010 ( .A1(n19856), .A2(n19945), .B1(n19941), .B2(n19855), .ZN(
        n19859) );
  AOI22_X1 U22011 ( .A1(n19920), .A2(n19863), .B1(
        P2_INSTQUEUE_REG_13__0__SCAN_IN), .B2(n19857), .ZN(n19858) );
  OAI211_X1 U22012 ( .C1(n19926), .C2(n19860), .A(n19859), .B(n19858), .ZN(
        P2_U3152) );
  AOI22_X1 U22013 ( .A1(n19862), .A2(n19945), .B1(n19941), .B2(n19861), .ZN(
        n19866) );
  AOI22_X1 U22014 ( .A1(n19864), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n19863), .B2(n19944), .ZN(n19865) );
  OAI211_X1 U22015 ( .C1(n19951), .C2(n19873), .A(n19866), .B(n19865), .ZN(
        P2_U3144) );
  AOI22_X1 U22016 ( .A1(n19868), .A2(n19945), .B1(n19941), .B2(n19867), .ZN(
        n19872) );
  AOI22_X1 U22017 ( .A1(n19920), .A2(n19870), .B1(
        P2_INSTQUEUE_REG_11__0__SCAN_IN), .B2(n19869), .ZN(n19871) );
  OAI211_X1 U22018 ( .C1(n19926), .C2(n19873), .A(n19872), .B(n19871), .ZN(
        P2_U3136) );
  AOI22_X1 U22019 ( .A1(n19920), .A2(n19881), .B1(n19874), .B2(n19941), .ZN(
        n19878) );
  AOI22_X1 U22020 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19876), .B1(
        n19945), .B2(n19875), .ZN(n19877) );
  OAI211_X1 U22021 ( .C1(n19926), .C2(n19879), .A(n19878), .B(n19877), .ZN(
        P2_U3128) );
  AOI22_X1 U22022 ( .A1(n19944), .A2(n19881), .B1(n19880), .B2(n19941), .ZN(
        n19885) );
  AOI22_X1 U22023 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19883), .B1(
        n19945), .B2(n19882), .ZN(n19884) );
  OAI211_X1 U22024 ( .C1(n19951), .C2(n19886), .A(n19885), .B(n19884), .ZN(
        P2_U3120) );
  AOI22_X1 U22025 ( .A1(n19944), .A2(n19888), .B1(n19887), .B2(n19941), .ZN(
        n19892) );
  AOI22_X1 U22026 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19890), .B1(
        n19889), .B2(n19945), .ZN(n19891) );
  OAI211_X1 U22027 ( .C1(n19951), .C2(n19899), .A(n19892), .B(n19891), .ZN(
        P2_U3112) );
  AOI22_X1 U22028 ( .A1(n19894), .A2(n19945), .B1(n19893), .B2(n19941), .ZN(
        n19898) );
  AOI22_X1 U22029 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19896), .B1(
        n19895), .B2(n19920), .ZN(n19897) );
  OAI211_X1 U22030 ( .C1(n19926), .C2(n19899), .A(n19898), .B(n19897), .ZN(
        P2_U3104) );
  AOI22_X1 U22031 ( .A1(n19901), .A2(n19945), .B1(n19941), .B2(n19900), .ZN(
        n19904) );
  AOI22_X1 U22032 ( .A1(n19920), .A2(n19907), .B1(
        P2_INSTQUEUE_REG_6__0__SCAN_IN), .B2(n19902), .ZN(n19903) );
  OAI211_X1 U22033 ( .C1(n19926), .C2(n19905), .A(n19904), .B(n19903), .ZN(
        P2_U3096) );
  AOI22_X1 U22034 ( .A1(n19944), .A2(n19907), .B1(n19941), .B2(n19906), .ZN(
        n19911) );
  AOI22_X1 U22035 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19909), .B1(
        n19945), .B2(n19908), .ZN(n19910) );
  OAI211_X1 U22036 ( .C1(n19951), .C2(n19912), .A(n19911), .B(n19910), .ZN(
        P2_U3088) );
  AOI22_X1 U22037 ( .A1(n19944), .A2(n19914), .B1(n19913), .B2(n19941), .ZN(
        n19918) );
  AOI22_X1 U22038 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19916), .B1(
        n19945), .B2(n19915), .ZN(n19917) );
  OAI211_X1 U22039 ( .C1(n19951), .C2(n19925), .A(n19918), .B(n19917), .ZN(
        P2_U3080) );
  AOI22_X1 U22040 ( .A1(n19920), .A2(n19929), .B1(n19941), .B2(n19919), .ZN(
        n19924) );
  AOI22_X1 U22041 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19922), .B1(
        n19945), .B2(n19921), .ZN(n19923) );
  OAI211_X1 U22042 ( .C1(n19926), .C2(n19925), .A(n19924), .B(n19923), .ZN(
        P2_U3072) );
  AOI22_X1 U22043 ( .A1(n19928), .A2(n19945), .B1(n19941), .B2(n19927), .ZN(
        n19932) );
  AOI22_X1 U22044 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19930), .B1(
        n19929), .B2(n19944), .ZN(n19931) );
  OAI211_X1 U22045 ( .C1(n19951), .C2(n19933), .A(n19932), .B(n19931), .ZN(
        P2_U3064) );
  AOI22_X1 U22046 ( .A1(n19935), .A2(n19945), .B1(n19941), .B2(n19934), .ZN(
        n19939) );
  AOI22_X1 U22047 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19937), .B1(
        n19936), .B2(n19944), .ZN(n19938) );
  OAI211_X1 U22048 ( .C1(n19951), .C2(n19940), .A(n19939), .B(n19938), .ZN(
        P2_U3056) );
  AOI22_X1 U22049 ( .A1(n19944), .A2(n19943), .B1(n19942), .B2(n19941), .ZN(
        n19949) );
  AOI22_X1 U22050 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19947), .B1(
        n19946), .B2(n19945), .ZN(n19948) );
  OAI211_X1 U22051 ( .C1(n19951), .C2(n19950), .A(n19949), .B(n19948), .ZN(
        P2_U3048) );
  INV_X1 U22052 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n20269) );
  INV_X1 U22053 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n19952) );
  AOI222_X1 U22054 ( .A1(n20269), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n20272), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n19952), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n19953) );
  INV_X2 U22055 ( .A(n19953), .ZN(n20013) );
  INV_X1 U22056 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19955) );
  AOI22_X1 U22057 ( .A1(n20002), .A2(n19955), .B1(n19954), .B2(n20013), .ZN(
        U376) );
  INV_X1 U22058 ( .A(n20013), .ZN(n20016) );
  INV_X1 U22059 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19957) );
  AOI22_X1 U22060 ( .A1(n20016), .A2(n19957), .B1(n19956), .B2(n20013), .ZN(
        U365) );
  INV_X1 U22061 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19959) );
  AOI22_X1 U22062 ( .A1(n20002), .A2(n19959), .B1(n19958), .B2(n20013), .ZN(
        U354) );
  INV_X1 U22063 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19961) );
  AOI22_X1 U22064 ( .A1(n20002), .A2(n19961), .B1(n19960), .B2(n20013), .ZN(
        U353) );
  INV_X1 U22065 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19963) );
  AOI22_X1 U22066 ( .A1(n20002), .A2(n19963), .B1(n19962), .B2(n20013), .ZN(
        U352) );
  INV_X1 U22067 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19965) );
  AOI22_X1 U22068 ( .A1(n20002), .A2(n19965), .B1(n19964), .B2(n20013), .ZN(
        U351) );
  INV_X1 U22069 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19967) );
  AOI22_X1 U22070 ( .A1(n20016), .A2(n19967), .B1(n19966), .B2(n20013), .ZN(
        U350) );
  INV_X1 U22071 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19969) );
  AOI22_X1 U22072 ( .A1(n20002), .A2(n19969), .B1(n19968), .B2(n20013), .ZN(
        U349) );
  INV_X1 U22073 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19971) );
  AOI22_X1 U22074 ( .A1(n20002), .A2(n19971), .B1(n19970), .B2(n20013), .ZN(
        U348) );
  INV_X1 U22075 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19973) );
  AOI22_X1 U22076 ( .A1(n20002), .A2(n19973), .B1(n19972), .B2(n20013), .ZN(
        U347) );
  INV_X1 U22077 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19975) );
  AOI22_X1 U22078 ( .A1(n20002), .A2(n19975), .B1(n19974), .B2(n20013), .ZN(
        U375) );
  INV_X1 U22079 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19977) );
  AOI22_X1 U22080 ( .A1(n20002), .A2(n19977), .B1(n19976), .B2(n20013), .ZN(
        U374) );
  INV_X1 U22081 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19979) );
  AOI22_X1 U22082 ( .A1(n20002), .A2(n19979), .B1(n19978), .B2(n20013), .ZN(
        U373) );
  INV_X1 U22083 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19981) );
  AOI22_X1 U22084 ( .A1(n20002), .A2(n19981), .B1(n19980), .B2(n20013), .ZN(
        U372) );
  INV_X1 U22085 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19983) );
  AOI22_X1 U22086 ( .A1(n20002), .A2(n19983), .B1(n19982), .B2(n20013), .ZN(
        U371) );
  INV_X1 U22087 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19985) );
  AOI22_X1 U22088 ( .A1(n20002), .A2(n19985), .B1(n19984), .B2(n20013), .ZN(
        U370) );
  INV_X1 U22089 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19987) );
  AOI22_X1 U22090 ( .A1(n20002), .A2(n19987), .B1(n19986), .B2(n20013), .ZN(
        U369) );
  INV_X1 U22091 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19989) );
  AOI22_X1 U22092 ( .A1(n20002), .A2(n19989), .B1(n19988), .B2(n20013), .ZN(
        U368) );
  INV_X1 U22093 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19991) );
  AOI22_X1 U22094 ( .A1(n20002), .A2(n19991), .B1(n19990), .B2(n20013), .ZN(
        U367) );
  INV_X1 U22095 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19993) );
  AOI22_X1 U22096 ( .A1(n20002), .A2(n19993), .B1(n19992), .B2(n20013), .ZN(
        U366) );
  INV_X1 U22097 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19995) );
  AOI22_X1 U22098 ( .A1(n20002), .A2(n19995), .B1(n19994), .B2(n20013), .ZN(
        U364) );
  INV_X1 U22099 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19997) );
  AOI22_X1 U22100 ( .A1(n20002), .A2(n19997), .B1(n19996), .B2(n20013), .ZN(
        U363) );
  INV_X1 U22101 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19999) );
  AOI22_X1 U22102 ( .A1(n20002), .A2(n19999), .B1(n19998), .B2(n20013), .ZN(
        U362) );
  INV_X1 U22103 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n20001) );
  AOI22_X1 U22104 ( .A1(n20002), .A2(n20001), .B1(n20000), .B2(n20013), .ZN(
        U361) );
  INV_X1 U22105 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n20004) );
  AOI22_X1 U22106 ( .A1(n20016), .A2(n20004), .B1(n20003), .B2(n20013), .ZN(
        U360) );
  INV_X1 U22107 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n20006) );
  AOI22_X1 U22108 ( .A1(n20016), .A2(n20006), .B1(n20005), .B2(n20013), .ZN(
        U359) );
  INV_X1 U22109 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n20008) );
  AOI22_X1 U22110 ( .A1(n20016), .A2(n20008), .B1(n20007), .B2(n20013), .ZN(
        U358) );
  INV_X1 U22111 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n20010) );
  AOI22_X1 U22112 ( .A1(n20016), .A2(n20010), .B1(n20009), .B2(n20013), .ZN(
        U357) );
  INV_X1 U22113 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n20012) );
  AOI22_X1 U22114 ( .A1(n20016), .A2(n20012), .B1(n20011), .B2(n20013), .ZN(
        U356) );
  INV_X1 U22115 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n20015) );
  AOI22_X1 U22116 ( .A1(n20016), .A2(n20015), .B1(n20014), .B2(n20013), .ZN(
        U355) );
  AOI22_X1 U22117 ( .A1(n21515), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20018) );
  OAI21_X1 U22118 ( .B1(n20019), .B2(n20044), .A(n20018), .ZN(P1_U2936) );
  INV_X1 U22119 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20021) );
  AOI22_X1 U22120 ( .A1(n20031), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20020) );
  OAI21_X1 U22121 ( .B1(n20021), .B2(n20044), .A(n20020), .ZN(P1_U2935) );
  AOI22_X1 U22122 ( .A1(n20031), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20022) );
  OAI21_X1 U22123 ( .B1(n20023), .B2(n20044), .A(n20022), .ZN(P1_U2934) );
  AOI22_X1 U22124 ( .A1(n20031), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20024) );
  OAI21_X1 U22125 ( .B1(n20025), .B2(n20044), .A(n20024), .ZN(P1_U2933) );
  AOI22_X1 U22126 ( .A1(n20031), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20026) );
  OAI21_X1 U22127 ( .B1(n20027), .B2(n20044), .A(n20026), .ZN(P1_U2932) );
  AOI22_X1 U22128 ( .A1(n20031), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20028) );
  OAI21_X1 U22129 ( .B1(n13169), .B2(n20044), .A(n20028), .ZN(P1_U2931) );
  AOI22_X1 U22130 ( .A1(n20031), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20029) );
  OAI21_X1 U22131 ( .B1(n13176), .B2(n20044), .A(n20029), .ZN(P1_U2930) );
  AOI22_X1 U22132 ( .A1(n21515), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20030) );
  OAI21_X1 U22133 ( .B1(n13184), .B2(n20044), .A(n20030), .ZN(P1_U2929) );
  INV_X1 U22134 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n21891) );
  AOI22_X1 U22135 ( .A1(n20031), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20032) );
  OAI21_X1 U22136 ( .B1(n21891), .B2(n20044), .A(n20032), .ZN(P1_U2928) );
  AOI22_X1 U22137 ( .A1(n21515), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20033) );
  OAI21_X1 U22138 ( .B1(n21899), .B2(n20044), .A(n20033), .ZN(P1_U2927) );
  INV_X1 U22139 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20036) );
  AOI22_X1 U22140 ( .A1(n21515), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20035) );
  OAI21_X1 U22141 ( .B1(n20036), .B2(n20044), .A(n20035), .ZN(P1_U2926) );
  AOI22_X1 U22142 ( .A1(n21515), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20037) );
  OAI21_X1 U22143 ( .B1(n21919), .B2(n20044), .A(n20037), .ZN(P1_U2925) );
  AOI22_X1 U22144 ( .A1(n21515), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20038) );
  OAI21_X1 U22145 ( .B1(n21929), .B2(n20044), .A(n20038), .ZN(P1_U2924) );
  INV_X1 U22146 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20040) );
  AOI22_X1 U22147 ( .A1(n21515), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20039) );
  OAI21_X1 U22148 ( .B1(n20040), .B2(n20044), .A(n20039), .ZN(P1_U2923) );
  INV_X1 U22149 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20042) );
  AOI22_X1 U22150 ( .A1(n21515), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20041) );
  OAI21_X1 U22151 ( .B1(n20042), .B2(n20044), .A(n20041), .ZN(P1_U2922) );
  AOI22_X1 U22152 ( .A1(n21515), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n20034), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20043) );
  OAI21_X1 U22153 ( .B1(n20045), .B2(n20044), .A(n20043), .ZN(P1_U2921) );
  AND2_X1 U22154 ( .A1(n22401), .A2(n21840), .ZN(n20065) );
  INV_X2 U22155 ( .A(n20065), .ZN(n20090) );
  AND2_X1 U22156 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n22401), .ZN(n20068) );
  OAI222_X1 U22157 ( .A1(n20090), .A2(n20047), .B1(n20046), .B2(n22401), .C1(
        n14907), .C2(n10965), .ZN(P1_U3197) );
  INV_X1 U22158 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n20048) );
  OAI222_X1 U22159 ( .A1(n20090), .A2(n20049), .B1(n20048), .B2(n22401), .C1(
        n20047), .C2(n10965), .ZN(P1_U3198) );
  INV_X1 U22160 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20050) );
  OAI222_X1 U22161 ( .A1(n20090), .A2(n21621), .B1(n20050), .B2(n22401), .C1(
        n20049), .C2(n10965), .ZN(P1_U3199) );
  INV_X1 U22162 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20051) );
  OAI222_X1 U22163 ( .A1(n20090), .A2(n21627), .B1(n20051), .B2(n22401), .C1(
        n21621), .C2(n10965), .ZN(P1_U3200) );
  INV_X1 U22164 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n20052) );
  OAI222_X1 U22165 ( .A1(n20090), .A2(n20053), .B1(n20052), .B2(n22401), .C1(
        n21627), .C2(n10965), .ZN(P1_U3201) );
  INV_X1 U22166 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n20054) );
  OAI222_X1 U22167 ( .A1(n20090), .A2(n21655), .B1(n20054), .B2(n22401), .C1(
        n20053), .C2(n10965), .ZN(P1_U3202) );
  INV_X1 U22168 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n20055) );
  OAI222_X1 U22169 ( .A1(n10965), .A2(n21655), .B1(n20055), .B2(n22401), .C1(
        n21667), .C2(n20090), .ZN(P1_U3203) );
  AOI22_X1 U22170 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n20065), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n22398), .ZN(n20056) );
  OAI21_X1 U22171 ( .B1(n21667), .B2(n10965), .A(n20056), .ZN(P1_U3204) );
  INV_X1 U22172 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20058) );
  AOI22_X1 U22173 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n20065), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n22398), .ZN(n20057) );
  OAI21_X1 U22174 ( .B1(n20058), .B2(n10965), .A(n20057), .ZN(P1_U3205) );
  AOI22_X1 U22175 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n20068), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n22398), .ZN(n20059) );
  OAI21_X1 U22176 ( .B1(n21696), .B2(n20090), .A(n20059), .ZN(P1_U3206) );
  INV_X1 U22177 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n20060) );
  OAI222_X1 U22178 ( .A1(n10965), .A2(n21696), .B1(n20060), .B2(n22401), .C1(
        n21709), .C2(n20090), .ZN(P1_U3207) );
  INV_X1 U22179 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n20061) );
  OAI222_X1 U22180 ( .A1(n10965), .A2(n21709), .B1(n20061), .B2(n22401), .C1(
        n20063), .C2(n20090), .ZN(P1_U3208) );
  AOI22_X1 U22181 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n20065), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n22398), .ZN(n20062) );
  OAI21_X1 U22182 ( .B1(n20063), .B2(n10965), .A(n20062), .ZN(P1_U3209) );
  AOI22_X1 U22183 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n20068), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n22398), .ZN(n20064) );
  OAI21_X1 U22184 ( .B1(n20067), .B2(n20090), .A(n20064), .ZN(P1_U3210) );
  AOI22_X1 U22185 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n20065), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n22398), .ZN(n20066) );
  OAI21_X1 U22186 ( .B1(n20067), .B2(n10965), .A(n20066), .ZN(P1_U3211) );
  AOI22_X1 U22187 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n20068), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n22398), .ZN(n20069) );
  OAI21_X1 U22188 ( .B1(n20070), .B2(n20090), .A(n20069), .ZN(P1_U3212) );
  INV_X1 U22189 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n20071) );
  OAI222_X1 U22190 ( .A1(n20090), .A2(n21743), .B1(n20071), .B2(n22401), .C1(
        n20070), .C2(n10965), .ZN(P1_U3213) );
  INV_X1 U22191 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n20072) );
  INV_X1 U22192 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21744) );
  OAI222_X1 U22193 ( .A1(n10965), .A2(n21743), .B1(n20072), .B2(n22401), .C1(
        n21744), .C2(n20090), .ZN(P1_U3214) );
  INV_X1 U22194 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n20073) );
  OAI222_X1 U22195 ( .A1(n10965), .A2(n21744), .B1(n20073), .B2(n22401), .C1(
        n20074), .C2(n20090), .ZN(P1_U3215) );
  INV_X1 U22196 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n20075) );
  OAI222_X1 U22197 ( .A1(n20090), .A2(n20076), .B1(n20075), .B2(n22401), .C1(
        n20074), .C2(n10965), .ZN(P1_U3216) );
  INV_X1 U22198 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20077) );
  OAI222_X1 U22199 ( .A1(n20090), .A2(n20078), .B1(n20077), .B2(n22401), .C1(
        n20076), .C2(n10965), .ZN(P1_U3217) );
  INV_X1 U22200 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n20079) );
  OAI222_X1 U22201 ( .A1(n20090), .A2(n21599), .B1(n20079), .B2(n22401), .C1(
        n20078), .C2(n10965), .ZN(P1_U3218) );
  INV_X1 U22202 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n20080) );
  OAI222_X1 U22203 ( .A1(n20090), .A2(n16118), .B1(n20080), .B2(n22401), .C1(
        n21599), .C2(n10965), .ZN(P1_U3219) );
  INV_X1 U22204 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20081) );
  OAI222_X1 U22205 ( .A1(n10965), .A2(n16118), .B1(n20081), .B2(n22401), .C1(
        n20082), .C2(n20090), .ZN(P1_U3220) );
  INV_X1 U22206 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20083) );
  OAI222_X1 U22207 ( .A1(n20090), .A2(n20085), .B1(n20083), .B2(n22401), .C1(
        n20082), .C2(n10965), .ZN(P1_U3221) );
  INV_X1 U22208 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20084) );
  OAI222_X1 U22209 ( .A1(n10965), .A2(n20085), .B1(n20084), .B2(n22401), .C1(
        n21578), .C2(n20090), .ZN(P1_U3222) );
  INV_X1 U22210 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n20086) );
  OAI222_X1 U22211 ( .A1(n20090), .A2(n13652), .B1(n20086), .B2(n22401), .C1(
        n21578), .C2(n10965), .ZN(P1_U3223) );
  INV_X1 U22212 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n20087) );
  OAI222_X1 U22213 ( .A1(n10965), .A2(n13652), .B1(n20087), .B2(n22401), .C1(
        n20089), .C2(n20090), .ZN(P1_U3224) );
  INV_X1 U22214 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n20088) );
  OAI222_X1 U22215 ( .A1(n10965), .A2(n20089), .B1(n20088), .B2(n22401), .C1(
        n20093), .C2(n20090), .ZN(P1_U3225) );
  INV_X1 U22216 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20092) );
  OAI222_X1 U22217 ( .A1(n10965), .A2(n20093), .B1(n20092), .B2(n22401), .C1(
        n20091), .C2(n20090), .ZN(P1_U3226) );
  INV_X1 U22218 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20094) );
  AOI22_X1 U22219 ( .A1(n22401), .A2(n20095), .B1(n20094), .B2(n22398), .ZN(
        P1_U3458) );
  AOI221_X1 U22220 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(P1_REIP_REG_1__SCAN_IN), 
        .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(P1_REIP_REG_1__SCAN_IN), .A(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20106) );
  NOR4_X1 U22221 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20099) );
  NOR4_X1 U22222 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20098) );
  NOR4_X1 U22223 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n20097) );
  NOR4_X1 U22224 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n20096) );
  NAND4_X1 U22225 ( .A1(n20099), .A2(n20098), .A3(n20097), .A4(n20096), .ZN(
        n20105) );
  NOR4_X1 U22226 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n20103) );
  AOI211_X1 U22227 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_31__SCAN_IN), .B(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n20102) );
  NOR4_X1 U22228 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20101) );
  NOR4_X1 U22229 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20100) );
  NAND4_X1 U22230 ( .A1(n20103), .A2(n20102), .A3(n20101), .A4(n20100), .ZN(
        n20104) );
  NOR2_X1 U22231 ( .A1(n20105), .A2(n20104), .ZN(n20118) );
  MUX2_X1 U22232 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .B(n20106), .S(n20118), 
        .Z(P1_U2808) );
  INV_X1 U22233 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20107) );
  AOI22_X1 U22234 ( .A1(n22401), .A2(n20110), .B1(n20107), .B2(n22398), .ZN(
        P1_U3459) );
  AOI21_X1 U22235 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20108) );
  OAI221_X1 U22236 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20108), .C1(n14907), 
        .C2(P1_REIP_REG_0__SCAN_IN), .A(n20118), .ZN(n20109) );
  OAI21_X1 U22237 ( .B1(n20118), .B2(n20110), .A(n20109), .ZN(P1_U3481) );
  INV_X1 U22238 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20111) );
  AOI22_X1 U22239 ( .A1(n22401), .A2(n20114), .B1(n20111), .B2(n22398), .ZN(
        P1_U3460) );
  NOR3_X1 U22240 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20112) );
  OAI21_X1 U22241 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20112), .A(n20118), .ZN(
        n20113) );
  OAI21_X1 U22242 ( .B1(n20118), .B2(n20114), .A(n20113), .ZN(P1_U2807) );
  INV_X1 U22243 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20115) );
  AOI22_X1 U22244 ( .A1(n22401), .A2(n20117), .B1(n20115), .B2(n22398), .ZN(
        P1_U3461) );
  OAI21_X1 U22245 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20118), .ZN(n20116) );
  OAI21_X1 U22246 ( .B1(n20118), .B2(n20117), .A(n20116), .ZN(P1_U3482) );
  AOI22_X1 U22247 ( .A1(n20120), .A2(n13627), .B1(n13631), .B2(n20119), .ZN(
        n20121) );
  OAI21_X1 U22248 ( .B1(n20137), .B2(n20122), .A(n20121), .ZN(P1_U2869) );
  AOI22_X1 U22249 ( .A1(n20173), .A2(n13627), .B1(n20123), .B2(n13631), .ZN(
        n20124) );
  OAI21_X1 U22250 ( .B1(n20137), .B2(n20125), .A(n20124), .ZN(P1_U2855) );
  INV_X1 U22251 ( .A(n20126), .ZN(n21723) );
  AOI22_X1 U22252 ( .A1(n21725), .A2(n13627), .B1(n13631), .B2(n21723), .ZN(
        n20127) );
  OAI21_X1 U22253 ( .B1(n20137), .B2(n21719), .A(n20127), .ZN(P1_U2857) );
  AOI22_X1 U22254 ( .A1(n21679), .A2(n13627), .B1(n13631), .B2(n21673), .ZN(
        n20128) );
  OAI21_X1 U22255 ( .B1(n20137), .B2(n21676), .A(n20128), .ZN(P1_U2863) );
  AOI22_X1 U22256 ( .A1(n21665), .A2(n13627), .B1(n13631), .B2(n21662), .ZN(
        n20129) );
  OAI21_X1 U22257 ( .B1(n20137), .B2(n20130), .A(n20129), .ZN(P1_U2864) );
  AND2_X1 U22258 ( .A1(n20132), .A2(n20131), .ZN(n20133) );
  NOR2_X1 U22259 ( .A1(n20134), .A2(n20133), .ZN(n21625) );
  AOI22_X1 U22260 ( .A1(n21632), .A2(n13627), .B1(n13631), .B2(n21625), .ZN(
        n20135) );
  OAI21_X1 U22261 ( .B1(n20137), .B2(n20136), .A(n20135), .ZN(P1_U2867) );
  OR2_X1 U22262 ( .A1(n20192), .A2(n20138), .ZN(n20141) );
  INV_X1 U22263 ( .A(n20139), .ZN(n20140) );
  AOI22_X1 U22264 ( .A1(n20141), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B1(
        n20188), .B2(n20140), .ZN(n20143) );
  OAI211_X1 U22265 ( .C1(n20144), .C2(n20194), .A(n20143), .B(n20142), .ZN(
        P1_U2999) );
  INV_X1 U22266 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20149) );
  XOR2_X1 U22267 ( .A(n11005), .B(n20146), .Z(n21549) );
  INV_X1 U22268 ( .A(n21635), .ZN(n20147) );
  AOI222_X1 U22269 ( .A1(n21549), .A2(n20188), .B1(n20186), .B2(n21632), .C1(
        n20147), .C2(n20172), .ZN(n20148) );
  NAND2_X1 U22270 ( .A1(n21585), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n21545) );
  OAI211_X1 U22271 ( .C1(n20155), .C2(n20149), .A(n20148), .B(n21545), .ZN(
        P1_U2994) );
  INV_X1 U22272 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20154) );
  OAI22_X1 U22273 ( .A1(n21657), .A2(n20194), .B1(n21661), .B2(n20200), .ZN(
        n20150) );
  AOI21_X1 U22274 ( .B1(n20151), .B2(n20188), .A(n20150), .ZN(n20153) );
  OAI211_X1 U22275 ( .C1(n20155), .C2(n20154), .A(n20153), .B(n20152), .ZN(
        P1_U2992) );
  AOI22_X1 U22276 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n20192), .B1(
        n21585), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n20158) );
  INV_X1 U22277 ( .A(n20156), .ZN(n21688) );
  AOI22_X1 U22278 ( .A1(n21689), .A2(n20186), .B1(n20172), .B2(n21688), .ZN(
        n20157) );
  OAI211_X1 U22279 ( .C1(n21789), .C2(n20159), .A(n20158), .B(n20157), .ZN(
        P1_U2989) );
  OAI22_X1 U22280 ( .A1(n20160), .A2(n21789), .B1(n20200), .B2(n21701), .ZN(
        n20161) );
  OAI21_X1 U22281 ( .B1(n20194), .B2(n21698), .A(n20163), .ZN(P1_U2988) );
  AOI22_X1 U22282 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n20192), .B1(
        n21585), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n20166) );
  AOI22_X1 U22283 ( .A1(n20172), .A2(n21713), .B1(n20186), .B2(n20164), .ZN(
        n20165) );
  OAI211_X1 U22284 ( .C1(n20167), .C2(n21789), .A(n20166), .B(n20165), .ZN(
        P1_U2987) );
  AOI22_X1 U22285 ( .A1(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n20192), .B1(
        n21585), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n20169) );
  AOI22_X1 U22286 ( .A1(n21725), .A2(n20186), .B1(n21722), .B2(n20172), .ZN(
        n20168) );
  OAI211_X1 U22287 ( .C1(n20170), .C2(n21789), .A(n20169), .B(n20168), .ZN(
        P1_U2984) );
  AOI22_X1 U22288 ( .A1(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n20192), .B1(
        n21585), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n20175) );
  AOI22_X1 U22289 ( .A1(n20173), .A2(n20186), .B1(n20172), .B2(n20171), .ZN(
        n20174) );
  OAI211_X1 U22290 ( .C1(n20176), .C2(n21789), .A(n20175), .B(n20174), .ZN(
        P1_U2982) );
  AOI22_X1 U22291 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n20192), .B1(
        n21585), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n20179) );
  AOI22_X1 U22292 ( .A1(n21755), .A2(n20186), .B1(n20188), .B2(n20177), .ZN(
        n20178) );
  OAI211_X1 U22293 ( .C1(n20200), .C2(n21746), .A(n20179), .B(n20178), .ZN(
        P1_U2980) );
  AOI22_X1 U22294 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n20192), .B1(
        n21585), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n20190) );
  NAND2_X1 U22295 ( .A1(n20183), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n20180) );
  OAI211_X1 U22296 ( .C1(n20183), .C2(n20182), .A(n20181), .B(n20180), .ZN(
        n20184) );
  XNOR2_X1 U22297 ( .A(n20184), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n21568) );
  INV_X1 U22298 ( .A(n20185), .ZN(n20187) );
  AOI22_X1 U22299 ( .A1(n20188), .A2(n21568), .B1(n20187), .B2(n20186), .ZN(
        n20189) );
  OAI211_X1 U22300 ( .C1(n20200), .C2(n20191), .A(n20190), .B(n20189), .ZN(
        P1_U2978) );
  AOI22_X1 U22301 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n20192), .B1(
        n21585), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n20198) );
  XNOR2_X1 U22302 ( .A(n20182), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n20193) );
  XNOR2_X1 U22303 ( .A(n11000), .B(n20193), .ZN(n21593) );
  OAI22_X1 U22304 ( .A1(n20195), .A2(n20194), .B1(n21593), .B2(n21789), .ZN(
        n20196) );
  INV_X1 U22305 ( .A(n20196), .ZN(n20197) );
  OAI211_X1 U22306 ( .C1(n20200), .C2(n20199), .A(n20198), .B(n20197), .ZN(
        P1_U2976) );
  NOR2_X1 U22307 ( .A1(n20201), .A2(n21813), .ZN(n20203) );
  OAI22_X1 U22308 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20204), .B1(n20203), 
        .B2(n20202), .ZN(P1_U2803) );
  INV_X1 U22309 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n20205) );
  OAI222_X1 U22310 ( .A1(n22401), .A2(n20206), .B1(n22401), .B2(n20205), .C1(
        P1_CODEFETCH_REG_SCAN_IN), .C2(n22398), .ZN(P1_U2804) );
  AOI22_X1 U22311 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n10964), .ZN(n20208) );
  OAI21_X1 U22312 ( .B1(n20209), .B2(n20271), .A(n20208), .ZN(U247) );
  AOI22_X1 U22313 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n10964), .ZN(n20210) );
  OAI21_X1 U22314 ( .B1(n20211), .B2(n20271), .A(n20210), .ZN(U246) );
  AOI22_X1 U22315 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n10964), .ZN(n20212) );
  OAI21_X1 U22316 ( .B1(n20213), .B2(n20271), .A(n20212), .ZN(U245) );
  AOI22_X1 U22317 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n10964), .ZN(n20214) );
  OAI21_X1 U22318 ( .B1(n20215), .B2(n20271), .A(n20214), .ZN(U244) );
  AOI22_X1 U22319 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n10964), .ZN(n20216) );
  OAI21_X1 U22320 ( .B1(n20217), .B2(n20271), .A(n20216), .ZN(U243) );
  AOI22_X1 U22321 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n10964), .ZN(n20218) );
  OAI21_X1 U22322 ( .B1(n20219), .B2(n20271), .A(n20218), .ZN(U242) );
  AOI22_X1 U22323 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n10964), .ZN(n20220) );
  OAI21_X1 U22324 ( .B1(n20221), .B2(n20271), .A(n20220), .ZN(U241) );
  AOI22_X1 U22325 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n10964), .ZN(n20222) );
  OAI21_X1 U22326 ( .B1(n20223), .B2(n20271), .A(n20222), .ZN(U240) );
  INV_X1 U22327 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n20225) );
  AOI22_X1 U22328 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n10964), .ZN(n20224) );
  OAI21_X1 U22329 ( .B1(n20225), .B2(n20271), .A(n20224), .ZN(U239) );
  AOI22_X1 U22330 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n10964), .ZN(n20226) );
  OAI21_X1 U22331 ( .B1(n20227), .B2(n20271), .A(n20226), .ZN(U238) );
  AOI22_X1 U22332 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10964), .ZN(n20228) );
  OAI21_X1 U22333 ( .B1(n14671), .B2(n20271), .A(n20228), .ZN(U237) );
  AOI22_X1 U22334 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n10964), .ZN(n20229) );
  OAI21_X1 U22335 ( .B1(n20230), .B2(n20271), .A(n20229), .ZN(U236) );
  INV_X1 U22336 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n20232) );
  AOI22_X1 U22337 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n10964), .ZN(n20231) );
  OAI21_X1 U22338 ( .B1(n20232), .B2(n20271), .A(n20231), .ZN(U235) );
  AOI22_X1 U22339 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n10964), .ZN(n20233) );
  OAI21_X1 U22340 ( .B1(n20234), .B2(n20271), .A(n20233), .ZN(U234) );
  AOI22_X1 U22341 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n10964), .ZN(n20235) );
  OAI21_X1 U22342 ( .B1(n20236), .B2(n20271), .A(n20235), .ZN(U233) );
  AOI22_X1 U22343 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n10964), .ZN(n20237) );
  OAI21_X1 U22344 ( .B1(n14746), .B2(n20271), .A(n20237), .ZN(U232) );
  AOI22_X1 U22345 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n10964), .ZN(n20238) );
  OAI21_X1 U22346 ( .B1(n20239), .B2(n20271), .A(n20238), .ZN(U231) );
  AOI22_X1 U22347 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10964), .ZN(n20240) );
  OAI21_X1 U22348 ( .B1(n20241), .B2(n20271), .A(n20240), .ZN(U230) );
  AOI22_X1 U22349 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10964), .ZN(n20242) );
  OAI21_X1 U22350 ( .B1(n20243), .B2(n20271), .A(n20242), .ZN(U229) );
  AOI22_X1 U22351 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n10964), .ZN(n20244) );
  OAI21_X1 U22352 ( .B1(n20245), .B2(n20271), .A(n20244), .ZN(U228) );
  AOI22_X1 U22353 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n10964), .ZN(n20246) );
  OAI21_X1 U22354 ( .B1(n20247), .B2(n20271), .A(n20246), .ZN(U227) );
  AOI22_X1 U22355 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n10964), .ZN(n20248) );
  OAI21_X1 U22356 ( .B1(n20249), .B2(n20271), .A(n20248), .ZN(U226) );
  AOI22_X1 U22357 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n10964), .ZN(n20250) );
  OAI21_X1 U22358 ( .B1(n20251), .B2(n20271), .A(n20250), .ZN(U225) );
  AOI22_X1 U22359 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n10964), .ZN(n20252) );
  OAI21_X1 U22360 ( .B1(n20253), .B2(n20271), .A(n20252), .ZN(U224) );
  AOI22_X1 U22361 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n10964), .ZN(n20254) );
  OAI21_X1 U22362 ( .B1(n20255), .B2(n20271), .A(n20254), .ZN(U223) );
  AOI22_X1 U22363 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n10964), .ZN(n20256) );
  OAI21_X1 U22364 ( .B1(n20257), .B2(n20271), .A(n20256), .ZN(U222) );
  AOI22_X1 U22365 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n10964), .ZN(n20259) );
  OAI21_X1 U22366 ( .B1(n20260), .B2(n20271), .A(n20259), .ZN(U221) );
  AOI22_X1 U22367 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n10964), .ZN(n20261) );
  OAI21_X1 U22368 ( .B1(n20262), .B2(n20271), .A(n20261), .ZN(U220) );
  AOI22_X1 U22369 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n10964), .ZN(n20263) );
  OAI21_X1 U22370 ( .B1(n20264), .B2(n20271), .A(n20263), .ZN(U219) );
  AOI22_X1 U22371 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n10964), .ZN(n20265) );
  OAI21_X1 U22372 ( .B1(n20266), .B2(n20271), .A(n20265), .ZN(U218) );
  AOI22_X1 U22373 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n20258), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n10964), .ZN(n20267) );
  OAI21_X1 U22374 ( .B1(n20268), .B2(n20271), .A(n20267), .ZN(U217) );
  OAI222_X1 U22375 ( .A1(U212), .A2(n20272), .B1(n20271), .B2(n20270), .C1(
        U214), .C2(n20269), .ZN(U216) );
  AOI22_X1 U22376 ( .A1(n22401), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20273), 
        .B2(n22398), .ZN(P1_U3483) );
  OAI21_X1 U22377 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n20351), .A(n20348), 
        .ZN(n20274) );
  AOI211_X1 U22378 ( .C1(n20275), .C2(n20274), .A(n21876), .B(n21352), .ZN(
        n20277) );
  OAI21_X1 U22379 ( .B1(n20277), .B2(n20337), .A(n20276), .ZN(n20282) );
  AOI22_X1 U22380 ( .A1(n20279), .A2(n21478), .B1(n20278), .B2(n21500), .ZN(
        n20280) );
  NAND2_X1 U22381 ( .A1(n20280), .A2(n20339), .ZN(n20281) );
  MUX2_X1 U22382 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .B(n20282), .S(n20281), 
        .Z(P3_U3296) );
  NOR2_X1 U22383 ( .A1(n21476), .A2(n20283), .ZN(n20285) );
  NOR3_X1 U22384 ( .A1(n21876), .A2(n20284), .A3(n20283), .ZN(n20297) );
  AOI22_X1 U22385 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20333), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n20332), .ZN(n20286) );
  OAI21_X1 U22386 ( .B1(n20952), .B2(n20335), .A(n20286), .ZN(P3_U2768) );
  AOI22_X1 U22387 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20333), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n20332), .ZN(n20287) );
  OAI21_X1 U22388 ( .B1(n20890), .B2(n20335), .A(n20287), .ZN(P3_U2769) );
  AOI22_X1 U22389 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20333), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n20332), .ZN(n20288) );
  OAI21_X1 U22390 ( .B1(n20289), .B2(n20335), .A(n20288), .ZN(P3_U2770) );
  AOI22_X1 U22391 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20333), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n20332), .ZN(n20290) );
  OAI21_X1 U22392 ( .B1(n20291), .B2(n20335), .A(n20290), .ZN(P3_U2771) );
  AOI22_X1 U22393 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20333), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n20332), .ZN(n20292) );
  OAI21_X1 U22394 ( .B1(n20293), .B2(n20335), .A(n20292), .ZN(P3_U2772) );
  AOI22_X1 U22395 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20333), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n20332), .ZN(n20294) );
  OAI21_X1 U22396 ( .B1(n20860), .B2(n20335), .A(n20294), .ZN(P3_U2773) );
  AOI22_X1 U22397 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20333), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n20328), .ZN(n20295) );
  OAI21_X1 U22398 ( .B1(n20296), .B2(n20335), .A(n20295), .ZN(P3_U2774) );
  AOI22_X1 U22399 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20333), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n20328), .ZN(n20298) );
  OAI21_X1 U22400 ( .B1(n20943), .B2(n20335), .A(n20298), .ZN(P3_U2775) );
  AOI22_X1 U22401 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20333), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n20328), .ZN(n20299) );
  OAI21_X1 U22402 ( .B1(n20936), .B2(n20335), .A(n20299), .ZN(P3_U2776) );
  AOI22_X1 U22403 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20333), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n20328), .ZN(n20300) );
  OAI21_X1 U22404 ( .B1(n20896), .B2(n20335), .A(n20300), .ZN(P3_U2777) );
  AOI22_X1 U22405 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20333), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n20328), .ZN(n20301) );
  OAI21_X1 U22406 ( .B1(n20302), .B2(n20335), .A(n20301), .ZN(P3_U2778) );
  AOI22_X1 U22407 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20333), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n20328), .ZN(n20303) );
  OAI21_X1 U22408 ( .B1(n20929), .B2(n20335), .A(n20303), .ZN(P3_U2779) );
  AOI22_X1 U22409 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20333), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n20332), .ZN(n20304) );
  OAI21_X1 U22410 ( .B1(n20305), .B2(n20335), .A(n20304), .ZN(P3_U2780) );
  AOI22_X1 U22411 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20333), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n20332), .ZN(n20306) );
  OAI21_X1 U22412 ( .B1(n20307), .B2(n20335), .A(n20306), .ZN(P3_U2781) );
  AOI22_X1 U22413 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20333), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n20332), .ZN(n20308) );
  OAI21_X1 U22414 ( .B1(n20915), .B2(n20335), .A(n20308), .ZN(P3_U2782) );
  AOI22_X1 U22415 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20333), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n20332), .ZN(n20309) );
  OAI21_X1 U22416 ( .B1(n20979), .B2(n20335), .A(n20309), .ZN(P3_U2783) );
  AOI22_X1 U22417 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20333), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n20332), .ZN(n20310) );
  OAI21_X1 U22418 ( .B1(n20829), .B2(n20335), .A(n20310), .ZN(P3_U2784) );
  AOI22_X1 U22419 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20333), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n20332), .ZN(n20311) );
  OAI21_X1 U22420 ( .B1(n20312), .B2(n20335), .A(n20311), .ZN(P3_U2785) );
  AOI22_X1 U22421 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20333), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n20332), .ZN(n20313) );
  OAI21_X1 U22422 ( .B1(n20830), .B2(n20335), .A(n20313), .ZN(P3_U2786) );
  AOI22_X1 U22423 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20333), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n20332), .ZN(n20314) );
  OAI21_X1 U22424 ( .B1(n20315), .B2(n20335), .A(n20314), .ZN(P3_U2787) );
  AOI22_X1 U22425 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20333), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n20332), .ZN(n20316) );
  OAI21_X1 U22426 ( .B1(n20831), .B2(n20335), .A(n20316), .ZN(P3_U2788) );
  AOI22_X1 U22427 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20333), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n20332), .ZN(n20317) );
  OAI21_X1 U22428 ( .B1(n20318), .B2(n20335), .A(n20317), .ZN(P3_U2789) );
  AOI22_X1 U22429 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20333), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n20332), .ZN(n20319) );
  OAI21_X1 U22430 ( .B1(n20800), .B2(n20335), .A(n20319), .ZN(P3_U2790) );
  AOI22_X1 U22431 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20333), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n20332), .ZN(n20320) );
  OAI21_X1 U22432 ( .B1(n20975), .B2(n20335), .A(n20320), .ZN(P3_U2791) );
  AOI22_X1 U22433 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20333), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n20328), .ZN(n20321) );
  OAI21_X1 U22434 ( .B1(n20322), .B2(n20335), .A(n20321), .ZN(P3_U2792) );
  AOI22_X1 U22435 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20333), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n20328), .ZN(n20323) );
  OAI21_X1 U22436 ( .B1(n20324), .B2(n20335), .A(n20323), .ZN(P3_U2793) );
  AOI22_X1 U22437 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20333), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n20328), .ZN(n20325) );
  OAI21_X1 U22438 ( .B1(n20802), .B2(n20335), .A(n20325), .ZN(P3_U2794) );
  AOI22_X1 U22439 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20333), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n20328), .ZN(n20326) );
  OAI21_X1 U22440 ( .B1(n20327), .B2(n20335), .A(n20326), .ZN(P3_U2795) );
  AOI22_X1 U22441 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20333), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n20328), .ZN(n20329) );
  OAI21_X1 U22442 ( .B1(n20330), .B2(n20335), .A(n20329), .ZN(P3_U2796) );
  AOI22_X1 U22443 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20333), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n20332), .ZN(n20331) );
  OAI21_X1 U22444 ( .B1(n20960), .B2(n20335), .A(n20331), .ZN(P3_U2797) );
  AOI22_X1 U22445 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n20333), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n20332), .ZN(n20334) );
  OAI21_X1 U22446 ( .B1(n20336), .B2(n20335), .A(n20334), .ZN(P3_U2798) );
  AND4_X1 U22447 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n20337), .A3(n21352), 
        .A4(n21823), .ZN(n20606) );
  NAND2_X1 U22448 ( .A1(n21481), .A2(n20338), .ZN(n21497) );
  NAND4_X1 U22449 ( .A1(n21379), .A2(n20339), .A3(n21485), .A4(n21497), .ZN(
        n20612) );
  NAND2_X1 U22450 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n20351), .ZN(n20342) );
  AOI211_X4 U22451 ( .C1(n21478), .C2(n21823), .A(n20349), .B(n20342), .ZN(
        n20787) );
  INV_X1 U22452 ( .A(n20343), .ZN(n20345) );
  NOR2_X1 U22453 ( .A1(n20345), .A2(n20344), .ZN(n20998) );
  AOI22_X1 U22454 ( .A1(n20787), .A2(n20346), .B1(n20998), .B2(n20390), .ZN(
        n20356) );
  INV_X1 U22455 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n20783) );
  NOR2_X1 U22456 ( .A1(n20765), .A2(n20783), .ZN(n20347) );
  OR2_X1 U22457 ( .A1(n21485), .A2(n20347), .ZN(n20504) );
  AOI21_X1 U22458 ( .B1(n20606), .B2(n20347), .A(n20708), .ZN(n20353) );
  OAI211_X1 U22459 ( .C1(n20348), .C2(n20351), .A(n21478), .B(n21823), .ZN(
        n21477) );
  INV_X1 U22460 ( .A(n21477), .ZN(n20350) );
  AOI211_X4 U22461 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n20351), .A(n20350), .B(
        n20349), .ZN(n20788) );
  AOI22_X1 U22462 ( .A1(n20357), .A2(n20614), .B1(n20788), .B2(
        P3_EBX_REG_1__SCAN_IN), .ZN(n20352) );
  OAI221_X1 U22463 ( .B1(n20504), .B2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C1(
        n20353), .C2(n11129), .A(n20352), .ZN(n20354) );
  INV_X1 U22464 ( .A(n20354), .ZN(n20355) );
  OAI211_X1 U22465 ( .C1(n20357), .C2(n20612), .A(n20356), .B(n20355), .ZN(
        P3_U2670) );
  NAND2_X1 U22466 ( .A1(n20606), .A2(n20765), .ZN(n20506) );
  INV_X1 U22467 ( .A(n20358), .ZN(n20369) );
  INV_X1 U22468 ( .A(n20359), .ZN(n20360) );
  NOR3_X1 U22469 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .ZN(n20379) );
  AOI211_X1 U22470 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n20360), .A(n20379), .B(
        n20757), .ZN(n20365) );
  INV_X1 U22471 ( .A(n20612), .ZN(n20784) );
  OAI21_X1 U22472 ( .B1(n20344), .B2(n21006), .A(n21012), .ZN(n21010) );
  AOI22_X1 U22473 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n20784), .B1(n20390), 
        .B2(n21010), .ZN(n20362) );
  NAND2_X1 U22474 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .ZN(n20372) );
  OAI211_X1 U22475 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(P3_REIP_REG_1__SCAN_IN), 
        .A(n20614), .B(n20372), .ZN(n20361) );
  OAI211_X1 U22476 ( .C1(n20770), .C2(n20363), .A(n20362), .B(n20361), .ZN(
        n20364) );
  AOI211_X1 U22477 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n20788), .A(n20365), .B(
        n20364), .ZN(n20368) );
  NOR2_X1 U22478 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n11129), .ZN(
        n20591) );
  AOI21_X1 U22479 ( .B1(n20366), .B2(n20783), .A(n20765), .ZN(n20374) );
  OAI211_X1 U22480 ( .C1(n20591), .C2(n20369), .A(n20606), .B(n20374), .ZN(
        n20367) );
  OAI211_X1 U22481 ( .C1(n20506), .C2(n20369), .A(n20368), .B(n20367), .ZN(
        P3_U2669) );
  INV_X1 U22482 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20382) );
  INV_X1 U22483 ( .A(n21028), .ZN(n21030) );
  AOI21_X1 U22484 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21030), .A(
        n21461), .ZN(n21033) );
  NOR2_X1 U22485 ( .A1(n20370), .A2(n21033), .ZN(n21019) );
  NAND3_X1 U22486 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .A3(P3_REIP_REG_1__SCAN_IN), .ZN(n20398) );
  NAND2_X1 U22487 ( .A1(n20614), .A2(n20398), .ZN(n20371) );
  OAI22_X1 U22488 ( .A1(n21019), .A2(n20791), .B1(n20372), .B2(n20371), .ZN(
        n20377) );
  AOI21_X1 U22489 ( .B1(n20614), .B2(n20398), .A(n20784), .ZN(n20397) );
  XOR2_X1 U22490 ( .A(n20374), .B(n20373), .Z(n20375) );
  OAI22_X1 U22491 ( .A1(n20397), .A2(n21090), .B1(n21485), .B2(n20375), .ZN(
        n20376) );
  AOI211_X1 U22492 ( .C1(n20788), .C2(P3_EBX_REG_3__SCAN_IN), .A(n20377), .B(
        n20376), .ZN(n20381) );
  INV_X1 U22493 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n20378) );
  NAND2_X1 U22494 ( .A1(n20379), .A2(n20378), .ZN(n20389) );
  OAI211_X1 U22495 ( .C1(n20379), .C2(n20378), .A(n20787), .B(n20389), .ZN(
        n20380) );
  OAI211_X1 U22496 ( .C1(n20770), .C2(n20382), .A(n20381), .B(n20380), .ZN(
        P3_U2668) );
  INV_X1 U22497 ( .A(n20385), .ZN(n20384) );
  NAND2_X1 U22498 ( .A1(n20592), .A2(n20606), .ZN(n20383) );
  AOI211_X1 U22499 ( .C1(n18413), .C2(n20591), .A(n20384), .B(n20383), .ZN(
        n20388) );
  AOI211_X1 U22500 ( .C1(n20592), .C2(n20386), .A(n20385), .B(n20504), .ZN(
        n20387) );
  AOI211_X1 U22501 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n20788), .A(n20388), .B(
        n20387), .ZN(n20396) );
  NOR2_X1 U22502 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n20389), .ZN(n20407) );
  AOI211_X1 U22503 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n20389), .A(n20407), .B(
        n20757), .ZN(n20394) );
  NAND2_X1 U22504 ( .A1(n20614), .A2(n20399), .ZN(n20392) );
  OAI21_X1 U22505 ( .B1(n17998), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n20390), .ZN(n20391) );
  OAI211_X1 U22506 ( .C1(n20398), .C2(n20392), .A(n21379), .B(n20391), .ZN(
        n20393) );
  AOI211_X1 U22507 ( .C1(n20708), .C2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20394), .B(n20393), .ZN(n20395) );
  OAI211_X1 U22508 ( .C1(n20397), .C2(n20399), .A(n20396), .B(n20395), .ZN(
        P3_U2667) );
  NOR2_X1 U22509 ( .A1(n20399), .A2(n20398), .ZN(n20400) );
  NAND2_X1 U22510 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n20400), .ZN(n20429) );
  AOI21_X1 U22511 ( .B1(n20614), .B2(n20429), .A(n20784), .ZN(n20425) );
  AOI21_X1 U22512 ( .B1(n20614), .B2(n20400), .A(P3_REIP_REG_5__SCAN_IN), .ZN(
        n20404) );
  AOI21_X1 U22513 ( .B1(n18413), .B2(n20591), .A(n20765), .ZN(n20401) );
  XNOR2_X1 U22514 ( .A(n20402), .B(n20401), .ZN(n20403) );
  OAI22_X1 U22515 ( .A1(n20425), .A2(n20404), .B1(n21485), .B2(n20403), .ZN(
        n20405) );
  AOI211_X1 U22516 ( .C1(n20788), .C2(P3_EBX_REG_5__SCAN_IN), .A(n21401), .B(
        n20405), .ZN(n20409) );
  INV_X1 U22517 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n20406) );
  NAND2_X1 U22518 ( .A1(n20407), .A2(n20406), .ZN(n20411) );
  OAI211_X1 U22519 ( .C1(n20407), .C2(n20406), .A(n20787), .B(n20411), .ZN(
        n20408) );
  OAI211_X1 U22520 ( .C1(n20770), .C2(n20410), .A(n20409), .B(n20408), .ZN(
        P3_U2666) );
  INV_X1 U22521 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n20422) );
  AOI211_X1 U22522 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n20411), .A(n20432), .B(
        n20757), .ZN(n20420) );
  INV_X1 U22523 ( .A(n20412), .ZN(n20413) );
  AOI21_X1 U22524 ( .B1(n20592), .B2(n20413), .A(n20504), .ZN(n20417) );
  NAND2_X1 U22525 ( .A1(n20414), .A2(n20591), .ZN(n20491) );
  NAND2_X1 U22526 ( .A1(n20592), .A2(n20491), .ZN(n20479) );
  OAI21_X1 U22527 ( .B1(n21485), .B2(n20479), .A(n20416), .ZN(n20415) );
  OAI21_X1 U22528 ( .B1(n20417), .B2(n20416), .A(n20415), .ZN(n20418) );
  OAI211_X1 U22529 ( .C1(n20425), .C2(n20430), .A(n20418), .B(n21379), .ZN(
        n20419) );
  AOI211_X1 U22530 ( .C1(n20708), .C2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n20420), .B(n20419), .ZN(n20421) );
  OR3_X1 U22531 ( .A1(n20598), .A2(n20429), .A3(P3_REIP_REG_6__SCAN_IN), .ZN(
        n20424) );
  OAI211_X1 U22532 ( .C1(n20422), .C2(n20768), .A(n20421), .B(n20424), .ZN(
        P3_U2665) );
  XNOR2_X1 U22533 ( .A(n20423), .B(n20479), .ZN(n20428) );
  AOI21_X1 U22534 ( .B1(n20425), .B2(n20424), .A(n21128), .ZN(n20427) );
  OAI22_X1 U22535 ( .A1(n20436), .A2(n20770), .B1(n20768), .B2(n20431), .ZN(
        n20426) );
  AOI211_X1 U22536 ( .C1(n20606), .C2(n20428), .A(n20427), .B(n20426), .ZN(
        n20435) );
  NOR2_X1 U22537 ( .A1(n20430), .A2(n20429), .ZN(n20441) );
  NAND3_X1 U22538 ( .A1(n20614), .A2(n20441), .A3(n21128), .ZN(n20434) );
  NAND2_X1 U22539 ( .A1(n20432), .A2(n20431), .ZN(n20439) );
  OAI211_X1 U22540 ( .C1(n20432), .C2(n20431), .A(n20787), .B(n20439), .ZN(
        n20433) );
  NAND4_X1 U22541 ( .A1(n20435), .A2(n21379), .A3(n20434), .A4(n20433), .ZN(
        P3_U2664) );
  OAI21_X1 U22542 ( .B1(n20436), .B2(n20491), .A(n20592), .ZN(n20437) );
  XNOR2_X1 U22543 ( .A(n20438), .B(n20437), .ZN(n20449) );
  AOI211_X1 U22544 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n20439), .A(n20459), .B(
        n20757), .ZN(n20440) );
  AOI21_X1 U22545 ( .B1(n20708), .B2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n20440), .ZN(n20448) );
  NAND2_X1 U22546 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n20441), .ZN(n20445) );
  NOR2_X1 U22547 ( .A1(n20442), .A2(n20445), .ZN(n20463) );
  OAI21_X1 U22548 ( .B1(n20463), .B2(n20598), .A(n20612), .ZN(n20469) );
  INV_X1 U22549 ( .A(n20463), .ZN(n20452) );
  NAND2_X1 U22550 ( .A1(n20614), .A2(n20452), .ZN(n20444) );
  OAI22_X1 U22551 ( .A1(n20445), .A2(n20444), .B1(n20768), .B2(n20443), .ZN(
        n20446) );
  AOI211_X1 U22552 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n20469), .A(n21401), .B(
        n20446), .ZN(n20447) );
  OAI211_X1 U22553 ( .C1(n21485), .C2(n20449), .A(n20448), .B(n20447), .ZN(
        P3_U2663) );
  AOI211_X1 U22554 ( .C1(n20450), .C2(n20506), .A(n20453), .B(n20504), .ZN(
        n20458) );
  OAI21_X1 U22555 ( .B1(n20451), .B2(n20491), .A(n20592), .ZN(n20467) );
  NOR2_X1 U22556 ( .A1(n21485), .A2(n20467), .ZN(n20454) );
  NOR3_X1 U22557 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n20598), .A3(n20452), .ZN(
        n20470) );
  AOI21_X1 U22558 ( .B1(n20454), .B2(n20453), .A(n20470), .ZN(n20455) );
  OAI211_X1 U22559 ( .C1(n20456), .C2(n20770), .A(n20455), .B(n21379), .ZN(
        n20457) );
  AOI211_X1 U22560 ( .C1(P3_REIP_REG_9__SCAN_IN), .C2(n20469), .A(n20458), .B(
        n20457), .ZN(n20461) );
  NAND2_X1 U22561 ( .A1(n20459), .A2(n20462), .ZN(n20464) );
  OAI211_X1 U22562 ( .C1(n20459), .C2(n20462), .A(n20787), .B(n20464), .ZN(
        n20460) );
  OAI211_X1 U22563 ( .C1(n20462), .C2(n20768), .A(n20461), .B(n20460), .ZN(
        P3_U2662) );
  AOI22_X1 U22564 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n20708), .B1(
        n20788), .B2(P3_EBX_REG_10__SCAN_IN), .ZN(n20474) );
  NAND2_X1 U22565 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n20463), .ZN(n20475) );
  NOR2_X1 U22566 ( .A1(n20598), .A2(n20475), .ZN(n20478) );
  AOI211_X1 U22567 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n20464), .A(n20487), .B(
        n20757), .ZN(n20465) );
  AOI211_X1 U22568 ( .C1(n20478), .C2(n20477), .A(n21401), .B(n20465), .ZN(
        n20473) );
  AOI21_X1 U22569 ( .B1(n20468), .B2(n20467), .A(n21485), .ZN(n20466) );
  OAI21_X1 U22570 ( .B1(n20468), .B2(n20467), .A(n20466), .ZN(n20472) );
  OAI21_X1 U22571 ( .B1(n20470), .B2(n20469), .A(P3_REIP_REG_10__SCAN_IN), 
        .ZN(n20471) );
  NAND4_X1 U22572 ( .A1(n20474), .A2(n20473), .A3(n20472), .A4(n20471), .ZN(
        P3_U2661) );
  NOR3_X1 U22573 ( .A1(n20477), .A2(n20476), .A3(n20475), .ZN(n20568) );
  OAI21_X1 U22574 ( .B1(n20568), .B2(n20598), .A(n20612), .ZN(n20526) );
  INV_X1 U22575 ( .A(n20526), .ZN(n20501) );
  AOI21_X1 U22576 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n20478), .A(
        P3_REIP_REG_11__SCAN_IN), .ZN(n20484) );
  OAI21_X1 U22577 ( .B1(n20480), .B2(n20765), .A(n20479), .ZN(n20481) );
  XNOR2_X1 U22578 ( .A(n20482), .B(n20481), .ZN(n20483) );
  OAI22_X1 U22579 ( .A1(n20501), .A2(n20484), .B1(n21485), .B2(n20483), .ZN(
        n20485) );
  AOI211_X1 U22580 ( .C1(n20788), .C2(P3_EBX_REG_11__SCAN_IN), .A(n21401), .B(
        n20485), .ZN(n20489) );
  NAND2_X1 U22581 ( .A1(n20487), .A2(n20486), .ZN(n20496) );
  OAI211_X1 U22582 ( .C1(n20487), .C2(n20486), .A(n20787), .B(n20496), .ZN(
        n20488) );
  OAI211_X1 U22583 ( .C1(n20770), .C2(n20490), .A(n20489), .B(n20488), .ZN(
        P3_U2660) );
  NAND2_X1 U22584 ( .A1(n20614), .A2(n20568), .ZN(n20537) );
  NOR2_X1 U22585 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n20537), .ZN(n20513) );
  AOI211_X1 U22586 ( .C1(n20788), .C2(P3_EBX_REG_12__SCAN_IN), .A(n21401), .B(
        n20513), .ZN(n20500) );
  OAI21_X1 U22587 ( .B1(n20492), .B2(n20491), .A(n20592), .ZN(n20495) );
  OAI21_X1 U22588 ( .B1(n20495), .B2(n20494), .A(n20606), .ZN(n20493) );
  AOI21_X1 U22589 ( .B1(n20495), .B2(n20494), .A(n20493), .ZN(n20498) );
  AOI211_X1 U22590 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n20496), .A(n20508), .B(
        n20757), .ZN(n20497) );
  AOI211_X1 U22591 ( .C1(n20708), .C2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n20498), .B(n20497), .ZN(n20499) );
  OAI211_X1 U22592 ( .C1(n20501), .C2(n20524), .A(n20500), .B(n20499), .ZN(
        P3_U2659) );
  NOR2_X1 U22593 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n20537), .ZN(n20503) );
  NOR2_X1 U22594 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20502), .ZN(
        n20533) );
  NOR3_X1 U22595 ( .A1(n20533), .A2(n21485), .A3(n20765), .ZN(n20523) );
  AOI22_X1 U22596 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n20503), .B1(n20523), 
        .B2(n20505), .ZN(n20516) );
  AOI211_X1 U22597 ( .C1(n20507), .C2(n20506), .A(n20505), .B(n20504), .ZN(
        n20512) );
  NAND2_X1 U22598 ( .A1(n20508), .A2(n20510), .ZN(n20517) );
  OAI211_X1 U22599 ( .C1(n20508), .C2(n20510), .A(n20787), .B(n20517), .ZN(
        n20509) );
  OAI211_X1 U22600 ( .C1(n20768), .C2(n20510), .A(n21379), .B(n20509), .ZN(
        n20511) );
  AOI211_X1 U22601 ( .C1(n20708), .C2(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n20512), .B(n20511), .ZN(n20515) );
  OAI21_X1 U22602 ( .B1(n20513), .B2(n20526), .A(P3_REIP_REG_13__SCAN_IN), 
        .ZN(n20514) );
  NAND3_X1 U22603 ( .A1(n20516), .A2(n20515), .A3(n20514), .ZN(P3_U2658) );
  INV_X1 U22604 ( .A(n20529), .ZN(n20522) );
  AOI211_X1 U22605 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n20517), .A(n20541), .B(
        n20757), .ZN(n20521) );
  OAI22_X1 U22606 ( .A1(n20519), .A2(n20770), .B1(n20768), .B2(n20518), .ZN(
        n20520) );
  AOI211_X1 U22607 ( .C1(n20523), .C2(n20522), .A(n20521), .B(n20520), .ZN(
        n20532) );
  NOR2_X1 U22608 ( .A1(n20525), .A2(n20524), .ZN(n20528) );
  INV_X1 U22609 ( .A(n20537), .ZN(n20552) );
  NAND3_X1 U22610 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .A3(P3_REIP_REG_12__SCAN_IN), .ZN(n20549) );
  NOR2_X1 U22611 ( .A1(n20614), .A2(n20784), .ZN(n20738) );
  INV_X1 U22612 ( .A(n20738), .ZN(n20786) );
  AOI21_X1 U22613 ( .B1(n20549), .B2(n20786), .A(n20526), .ZN(n20527) );
  INV_X1 U22614 ( .A(n20527), .ZN(n20557) );
  OAI221_X1 U22615 ( .B1(P3_REIP_REG_14__SCAN_IN), .B2(n20528), .C1(
        P3_REIP_REG_14__SCAN_IN), .C2(n20552), .A(n20557), .ZN(n20531) );
  OAI211_X1 U22616 ( .C1(n20533), .C2(n20765), .A(n20606), .B(n20529), .ZN(
        n20530) );
  NAND4_X1 U22617 ( .A1(n20532), .A2(n21379), .A3(n20531), .A4(n20530), .ZN(
        P3_U2657) );
  NAND2_X1 U22618 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n20533), .ZN(
        n20563) );
  NAND2_X1 U22619 ( .A1(n20592), .A2(n20563), .ZN(n20535) );
  OAI21_X1 U22620 ( .B1(n20536), .B2(n20535), .A(n20606), .ZN(n20534) );
  AOI21_X1 U22621 ( .B1(n20536), .B2(n20535), .A(n20534), .ZN(n20540) );
  NOR3_X1 U22622 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n20549), .A3(n20537), 
        .ZN(n20558) );
  AOI211_X1 U22623 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n20708), .A(
        n21401), .B(n20558), .ZN(n20538) );
  INV_X1 U22624 ( .A(n20538), .ZN(n20539) );
  AOI211_X1 U22625 ( .C1(P3_REIP_REG_15__SCAN_IN), .C2(n20557), .A(n20540), 
        .B(n20539), .ZN(n20543) );
  NAND2_X1 U22626 ( .A1(n20541), .A2(n20544), .ZN(n20548) );
  OAI211_X1 U22627 ( .C1(n20541), .C2(n20544), .A(n20787), .B(n20548), .ZN(
        n20542) );
  OAI211_X1 U22628 ( .C1(n20544), .C2(n20768), .A(n20543), .B(n20542), .ZN(
        P3_U2656) );
  OAI21_X1 U22629 ( .B1(n20545), .B2(n20563), .A(n20592), .ZN(n20546) );
  XNOR2_X1 U22630 ( .A(n20547), .B(n20546), .ZN(n20561) );
  AOI211_X1 U22631 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n20548), .A(n20576), .B(
        n20757), .ZN(n20556) );
  NOR2_X1 U22632 ( .A1(n20550), .A2(n20549), .ZN(n20567) );
  NAND3_X1 U22633 ( .A1(n20567), .A2(n20552), .A3(n20551), .ZN(n20553) );
  OAI211_X1 U22634 ( .C1(n20554), .C2(n20770), .A(n21379), .B(n20553), .ZN(
        n20555) );
  AOI211_X1 U22635 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n20788), .A(n20556), .B(
        n20555), .ZN(n20560) );
  OAI21_X1 U22636 ( .B1(n20558), .B2(n20557), .A(P3_REIP_REG_16__SCAN_IN), 
        .ZN(n20559) );
  OAI211_X1 U22637 ( .C1(n21485), .C2(n20561), .A(n20560), .B(n20559), .ZN(
        P3_U2655) );
  INV_X1 U22638 ( .A(n20562), .ZN(n20564) );
  NOR2_X1 U22639 ( .A1(n20564), .A2(n20563), .ZN(n20616) );
  NOR2_X1 U22640 ( .A1(n20616), .A2(n20765), .ZN(n20566) );
  XOR2_X1 U22641 ( .A(n20566), .B(n20565), .Z(n20575) );
  NAND3_X1 U22642 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n20568), .A3(n20567), 
        .ZN(n20569) );
  NOR2_X1 U22643 ( .A1(n20573), .A2(n20569), .ZN(n20597) );
  NOR2_X1 U22644 ( .A1(n20597), .A2(n20598), .ZN(n20570) );
  NOR2_X1 U22645 ( .A1(n20784), .A2(n20570), .ZN(n20609) );
  INV_X1 U22646 ( .A(n20569), .ZN(n20571) );
  AOI22_X1 U22647 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n20708), .B1(
        n20571), .B2(n20570), .ZN(n20572) );
  OAI211_X1 U22648 ( .C1(n20609), .C2(n20573), .A(n20572), .B(n21379), .ZN(
        n20574) );
  AOI21_X1 U22649 ( .B1(n20575), .B2(n20606), .A(n20574), .ZN(n20578) );
  NAND2_X1 U22650 ( .A1(n20576), .A2(n20579), .ZN(n20580) );
  OAI211_X1 U22651 ( .C1(n20576), .C2(n20579), .A(n20787), .B(n20580), .ZN(
        n20577) );
  OAI211_X1 U22652 ( .C1(n20579), .C2(n20768), .A(n20578), .B(n20577), .ZN(
        P3_U2654) );
  AOI211_X1 U22653 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n20580), .A(n20600), .B(
        n20757), .ZN(n20583) );
  INV_X1 U22654 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n20581) );
  NAND3_X1 U22655 ( .A1(n20614), .A2(n20597), .A3(n21378), .ZN(n20608) );
  OAI211_X1 U22656 ( .C1(n20581), .C2(n20770), .A(n21379), .B(n20608), .ZN(
        n20582) );
  AOI211_X1 U22657 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n20788), .A(n20583), .B(
        n20582), .ZN(n20590) );
  INV_X1 U22658 ( .A(n20584), .ZN(n20585) );
  OAI21_X1 U22659 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20585), .A(
        n20592), .ZN(n20588) );
  AOI21_X1 U22660 ( .B1(n20588), .B2(n20587), .A(n21485), .ZN(n20586) );
  OAI21_X1 U22661 ( .B1(n20588), .B2(n20587), .A(n20586), .ZN(n20589) );
  OAI211_X1 U22662 ( .C1(n20609), .C2(n21378), .A(n20590), .B(n20589), .ZN(
        P3_U2653) );
  INV_X1 U22663 ( .A(n20591), .ZN(n20593) );
  OAI21_X1 U22664 ( .B1(n20594), .B2(n20593), .A(n20592), .ZN(n20595) );
  XOR2_X1 U22665 ( .A(n20596), .B(n20595), .Z(n20605) );
  INV_X1 U22666 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n20603) );
  NAND2_X1 U22667 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n20597), .ZN(n20610) );
  NOR3_X1 U22668 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n20598), .A3(n20610), 
        .ZN(n20599) );
  AOI211_X1 U22669 ( .C1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(n20708), .A(
        n21401), .B(n20599), .ZN(n20602) );
  NAND2_X1 U22670 ( .A1(n20600), .A2(n20603), .ZN(n20620) );
  OAI211_X1 U22671 ( .C1(n20600), .C2(n20603), .A(n20787), .B(n20620), .ZN(
        n20601) );
  OAI211_X1 U22672 ( .C1(n20603), .C2(n20768), .A(n20602), .B(n20601), .ZN(
        n20604) );
  AOI21_X1 U22673 ( .B1(n20606), .B2(n20605), .A(n20604), .ZN(n20607) );
  OAI221_X1 U22674 ( .B1(n20611), .B2(n20609), .C1(n20611), .C2(n20608), .A(
        n20607), .ZN(P3_U2652) );
  NOR2_X1 U22675 ( .A1(n20611), .A2(n20610), .ZN(n20613) );
  NAND3_X1 U22676 ( .A1(n20613), .A2(P3_REIP_REG_20__SCAN_IN), .A3(n20612), 
        .ZN(n20652) );
  NAND2_X1 U22677 ( .A1(n20786), .A2(n20652), .ZN(n20650) );
  AOI22_X1 U22678 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n20708), .B1(
        n20626), .B2(n20625), .ZN(n20624) );
  NOR2_X1 U22679 ( .A1(n20619), .A2(n20618), .ZN(n20627) );
  AOI211_X1 U22680 ( .C1(n20619), .C2(n20618), .A(n20627), .B(n21485), .ZN(
        n20622) );
  AOI211_X1 U22681 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n20620), .A(n20630), .B(
        n20757), .ZN(n20621) );
  AOI211_X1 U22682 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n20788), .A(n20622), .B(
        n20621), .ZN(n20623) );
  OAI211_X1 U22683 ( .C1(n20625), .C2(n20650), .A(n20624), .B(n20623), .ZN(
        P3_U2651) );
  NAND2_X1 U22684 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n20626), .ZN(n20646) );
  NOR2_X1 U22685 ( .A1(n20627), .A2(n20765), .ZN(n20628) );
  AOI211_X1 U22686 ( .C1(n20629), .C2(n20628), .A(n20637), .B(n21485), .ZN(
        n20634) );
  NAND2_X1 U22687 ( .A1(n20630), .A2(n20632), .ZN(n20640) );
  OAI211_X1 U22688 ( .C1(n20630), .C2(n20632), .A(n20787), .B(n20640), .ZN(
        n20631) );
  OAI21_X1 U22689 ( .B1(n20632), .B2(n20768), .A(n20631), .ZN(n20633) );
  AOI211_X1 U22690 ( .C1(n20708), .C2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n20634), .B(n20633), .ZN(n20635) );
  OAI221_X1 U22691 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n20646), .C1(n20636), 
        .C2(n20650), .A(n20635), .ZN(P3_U2650) );
  AOI211_X1 U22692 ( .C1(n20639), .C2(n20638), .A(n20654), .B(n21485), .ZN(
        n20645) );
  AOI211_X1 U22693 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n20640), .A(n20657), .B(
        n20757), .ZN(n20644) );
  OAI22_X1 U22694 ( .A1(n20642), .A2(n20770), .B1(n20768), .B2(n20641), .ZN(
        n20643) );
  NOR3_X1 U22695 ( .A1(n20645), .A2(n20644), .A3(n20643), .ZN(n20649) );
  NAND2_X1 U22696 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .ZN(n20647) );
  OAI211_X1 U22697 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(P3_REIP_REG_21__SCAN_IN), .A(n20665), .B(n20647), .ZN(n20648) );
  OAI211_X1 U22698 ( .C1(n20651), .C2(n20650), .A(n20649), .B(n20648), .ZN(
        P3_U2649) );
  NAND3_X1 U22699 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .A3(n20665), .ZN(n20664) );
  NAND3_X1 U22700 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(P3_REIP_REG_22__SCAN_IN), 
        .A3(P3_REIP_REG_21__SCAN_IN), .ZN(n20653) );
  NOR2_X1 U22701 ( .A1(n20653), .A2(n20652), .ZN(n20684) );
  OR2_X1 U22702 ( .A1(n20738), .A2(n20684), .ZN(n20676) );
  NOR2_X1 U22703 ( .A1(n20656), .A2(n20655), .ZN(n20666) );
  AOI211_X1 U22704 ( .C1(n20656), .C2(n20655), .A(n20666), .B(n21485), .ZN(
        n20661) );
  NAND2_X1 U22705 ( .A1(n20657), .A2(n20659), .ZN(n20669) );
  OAI211_X1 U22706 ( .C1(n20657), .C2(n20659), .A(n20787), .B(n20669), .ZN(
        n20658) );
  OAI21_X1 U22707 ( .B1(n20659), .B2(n20768), .A(n20658), .ZN(n20660) );
  AOI211_X1 U22708 ( .C1(n20708), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n20661), .B(n20660), .ZN(n20662) );
  OAI221_X1 U22709 ( .B1(P3_REIP_REG_23__SCAN_IN), .B2(n20664), .C1(n20663), 
        .C2(n20676), .A(n20662), .ZN(P3_U2648) );
  NAND4_X1 U22710 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(P3_REIP_REG_22__SCAN_IN), 
        .A3(P3_REIP_REG_21__SCAN_IN), .A4(n20665), .ZN(n20677) );
  AOI211_X1 U22711 ( .C1(n20668), .C2(n20667), .A(n20680), .B(n21485), .ZN(
        n20674) );
  NOR2_X1 U22712 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n20669), .ZN(n20686) );
  AOI211_X1 U22713 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n20669), .A(n20686), .B(
        n20757), .ZN(n20673) );
  INV_X1 U22714 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n20670) );
  OAI22_X1 U22715 ( .A1(n20671), .A2(n20770), .B1(n20768), .B2(n20670), .ZN(
        n20672) );
  NOR3_X1 U22716 ( .A1(n20674), .A2(n20673), .A3(n20672), .ZN(n20675) );
  OAI221_X1 U22717 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n20677), .C1(n20678), 
        .C2(n20676), .A(n20675), .ZN(P3_U2647) );
  AOI22_X1 U22718 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n20708), .B1(
        n20788), .B2(P3_EBX_REG_25__SCAN_IN), .ZN(n20690) );
  NOR2_X1 U22719 ( .A1(n20678), .A2(n20677), .ZN(n20691) );
  INV_X1 U22720 ( .A(n20679), .ZN(n20682) );
  AOI211_X1 U22721 ( .C1(n20682), .C2(n20681), .A(n20695), .B(n21485), .ZN(
        n20683) );
  AOI21_X1 U22722 ( .B1(n20691), .B2(n20693), .A(n20683), .ZN(n20689) );
  NAND2_X1 U22723 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n20684), .ZN(n20692) );
  NAND3_X1 U22724 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n20786), .A3(n20692), 
        .ZN(n20688) );
  NAND2_X1 U22725 ( .A1(n20686), .A2(n20685), .ZN(n20698) );
  OAI211_X1 U22726 ( .C1(n20686), .C2(n20685), .A(n20787), .B(n20698), .ZN(
        n20687) );
  NAND4_X1 U22727 ( .A1(n20690), .A2(n20689), .A3(n20688), .A4(n20687), .ZN(
        P3_U2646) );
  NAND2_X1 U22728 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n20691), .ZN(n20706) );
  NOR3_X1 U22729 ( .A1(n20693), .A2(n20707), .A3(n20692), .ZN(n20739) );
  NOR2_X1 U22730 ( .A1(n20738), .A2(n20739), .ZN(n20720) );
  INV_X1 U22731 ( .A(n20720), .ZN(n20705) );
  INV_X1 U22732 ( .A(n20694), .ZN(n20697) );
  NOR2_X1 U22733 ( .A1(n20695), .A2(n20765), .ZN(n20696) );
  NOR2_X1 U22734 ( .A1(n20697), .A2(n20696), .ZN(n20712) );
  AOI211_X1 U22735 ( .C1(n20697), .C2(n20696), .A(n20712), .B(n21485), .ZN(
        n20703) );
  NOR2_X1 U22736 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n20698), .ZN(n20709) );
  AOI211_X1 U22737 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n20698), .A(n20709), .B(
        n20757), .ZN(n20702) );
  INV_X1 U22738 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n20700) );
  OAI22_X1 U22739 ( .A1(n20700), .A2(n20770), .B1(n20768), .B2(n20699), .ZN(
        n20701) );
  NOR3_X1 U22740 ( .A1(n20703), .A2(n20702), .A3(n20701), .ZN(n20704) );
  OAI221_X1 U22741 ( .B1(P3_REIP_REG_26__SCAN_IN), .B2(n20706), .C1(n20707), 
        .C2(n20705), .A(n20704), .ZN(P3_U2645) );
  INV_X1 U22742 ( .A(n20752), .ZN(n20719) );
  AOI22_X1 U22743 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n20708), .B1(
        P3_REIP_REG_27__SCAN_IN), .B2(n20720), .ZN(n20718) );
  NAND2_X1 U22744 ( .A1(n20709), .A2(n20710), .ZN(n20722) );
  NOR2_X1 U22745 ( .A1(n20709), .A2(n20710), .ZN(n20711) );
  OAI22_X1 U22746 ( .A1(n20757), .A2(n20711), .B1(n20768), .B2(n20710), .ZN(
        n20716) );
  NOR2_X1 U22747 ( .A1(n20712), .A2(n20765), .ZN(n20713) );
  AOI211_X1 U22748 ( .C1(n20714), .C2(n20713), .A(n20724), .B(n21485), .ZN(
        n20715) );
  AOI21_X1 U22749 ( .B1(n20722), .B2(n20716), .A(n20715), .ZN(n20717) );
  OAI211_X1 U22750 ( .C1(P3_REIP_REG_27__SCAN_IN), .C2(n20719), .A(n20718), 
        .B(n20717), .ZN(P3_U2644) );
  AOI22_X1 U22751 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n20720), .B1(n20788), 
        .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n20731) );
  NOR2_X1 U22752 ( .A1(n21317), .A2(n20721), .ZN(n20751) );
  AOI21_X1 U22753 ( .B1(n21317), .B2(n20721), .A(n20751), .ZN(n20729) );
  NOR2_X1 U22754 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n20722), .ZN(n20733) );
  AOI211_X1 U22755 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n20722), .A(n20733), .B(
        n20757), .ZN(n20728) );
  INV_X1 U22756 ( .A(n20723), .ZN(n20726) );
  AOI211_X1 U22757 ( .C1(n20726), .C2(n20725), .A(n20734), .B(n21485), .ZN(
        n20727) );
  AOI211_X1 U22758 ( .C1(n20729), .C2(n20752), .A(n20728), .B(n20727), .ZN(
        n20730) );
  OAI211_X1 U22759 ( .C1(n20732), .C2(n20770), .A(n20731), .B(n20730), .ZN(
        P3_U2643) );
  NOR2_X1 U22760 ( .A1(n20733), .A2(n15067), .ZN(n20749) );
  NAND2_X1 U22761 ( .A1(n20733), .A2(n15067), .ZN(n20756) );
  NAND2_X1 U22762 ( .A1(n20787), .A2(n20756), .ZN(n20754) );
  AOI21_X1 U22763 ( .B1(n11037), .B2(n20735), .A(n21485), .ZN(n20745) );
  INV_X1 U22764 ( .A(n20750), .ZN(n20744) );
  OAI22_X1 U22765 ( .A1(n20736), .A2(n20770), .B1(n20768), .B2(n15067), .ZN(
        n20737) );
  INV_X1 U22766 ( .A(n20737), .ZN(n20742) );
  AND2_X1 U22767 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n20751), .ZN(n20740) );
  AOI21_X1 U22768 ( .B1(n20740), .B2(n20739), .A(n20738), .ZN(n20777) );
  NAND2_X1 U22769 ( .A1(n20777), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n20741) );
  NAND3_X1 U22770 ( .A1(n20752), .A2(n20751), .A3(n20746), .ZN(n20747) );
  OAI211_X1 U22771 ( .C1(n20749), .C2(n20754), .A(n20748), .B(n20747), .ZN(
        P3_U2642) );
  NOR2_X1 U22772 ( .A1(n20750), .A2(n20765), .ZN(n20762) );
  XNOR2_X1 U22773 ( .A(n20763), .B(n20762), .ZN(n20760) );
  NAND3_X1 U22774 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n20752), .A3(n20751), 
        .ZN(n20782) );
  NOR2_X1 U22775 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n20782), .ZN(n20778) );
  OAI22_X1 U22776 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n20754), .B1(n20753), 
        .B2(n20770), .ZN(n20755) );
  AOI211_X1 U22777 ( .C1(P3_REIP_REG_30__SCAN_IN), .C2(n20777), .A(n20778), 
        .B(n20755), .ZN(n20759) );
  NOR2_X1 U22778 ( .A1(n20757), .A2(n20756), .ZN(n20767) );
  OAI21_X1 U22779 ( .B1(n20788), .B2(n20767), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n20758) );
  OAI211_X1 U22780 ( .C1(n20760), .C2(n21485), .A(n20759), .B(n20758), .ZN(
        P3_U2641) );
  NAND2_X1 U22781 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n20761), .ZN(n20781) );
  OR2_X1 U22782 ( .A1(n20763), .A2(n21485), .ZN(n20764) );
  NOR2_X1 U22783 ( .A1(n20765), .A2(n20764), .ZN(n20775) );
  INV_X1 U22784 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n20766) );
  NAND2_X1 U22785 ( .A1(n20767), .A2(n20766), .ZN(n20773) );
  INV_X1 U22786 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n20769) );
  OAI22_X1 U22787 ( .A1(n11131), .A2(n20770), .B1(n20769), .B2(n20768), .ZN(
        n20771) );
  OAI21_X1 U22788 ( .B1(n20778), .B2(n20777), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n20779) );
  OAI211_X1 U22789 ( .C1(n20782), .C2(n20781), .A(n20780), .B(n20779), .ZN(
        P3_U2640) );
  NOR3_X1 U22790 ( .A1(n20784), .A2(n21036), .A3(n20783), .ZN(n20785) );
  AOI21_X1 U22791 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(n20786), .A(n20785), .ZN(
        n20790) );
  OAI21_X1 U22792 ( .B1(n20788), .B2(n20787), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n20789) );
  OAI211_X1 U22793 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n20791), .A(
        n20790), .B(n20789), .ZN(P3_U2671) );
  NAND4_X1 U22794 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_5__SCAN_IN), .A4(P3_EAX_REG_4__SCAN_IN), .ZN(n20799) );
  INV_X1 U22795 ( .A(n20970), .ZN(n20827) );
  NOR4_X1 U22796 ( .A1(n20801), .A2(n20827), .A3(n20800), .A4(n20975), .ZN(
        n20821) );
  AND2_X1 U22797 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n20821), .ZN(n20824) );
  NAND2_X1 U22798 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n20824), .ZN(n20817) );
  NAND2_X1 U22799 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n20815), .ZN(n20808) );
  NAND2_X1 U22800 ( .A1(n20808), .A2(P3_EAX_REG_13__SCAN_IN), .ZN(n20807) );
  NAND2_X1 U22801 ( .A1(n20803), .A2(n20828), .ZN(n20853) );
  AOI22_X1 U22802 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20986), .B1(n20978), .B2(
        n20805), .ZN(n20806) );
  OAI221_X1 U22803 ( .B1(n20808), .B2(P3_EAX_REG_13__SCAN_IN), .C1(n20807), 
        .C2(n20959), .A(n20806), .ZN(P3_U2722) );
  INV_X1 U22804 ( .A(n20808), .ZN(n20957) );
  AOI21_X1 U22805 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n20966), .A(n20815), .ZN(
        n20810) );
  OAI222_X1 U22806 ( .A1(n20853), .A2(n20811), .B1(n20957), .B2(n20810), .C1(
        n20990), .C2(n20809), .ZN(P3_U2723) );
  INV_X1 U22807 ( .A(n20817), .ZN(n20812) );
  AOI21_X1 U22808 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n20966), .A(n20812), .ZN(
        n20814) );
  OAI222_X1 U22809 ( .A1(n20853), .A2(n20816), .B1(n20815), .B2(n20814), .C1(
        n20990), .C2(n20813), .ZN(P3_U2724) );
  NAND2_X1 U22810 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20986), .ZN(n20819) );
  OAI211_X1 U22811 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n20824), .A(n20966), .B(
        n20817), .ZN(n20818) );
  OAI211_X1 U22812 ( .C1(n20820), .C2(n20990), .A(n20819), .B(n20818), .ZN(
        P3_U2725) );
  AOI21_X1 U22813 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n20966), .A(n20821), .ZN(
        n20823) );
  OAI222_X1 U22814 ( .A1(n20853), .A2(n20900), .B1(n20824), .B2(n20823), .C1(
        n20990), .C2(n20822), .ZN(P3_U2726) );
  NAND2_X1 U22815 ( .A1(n20966), .A2(n20859), .ZN(n20974) );
  NOR2_X1 U22816 ( .A1(n20970), .A2(P3_EAX_REG_7__SCAN_IN), .ZN(n20825) );
  OAI222_X1 U22817 ( .A1(n20853), .A2(n20826), .B1(n20990), .B2(n21297), .C1(
        n20974), .C2(n20825), .ZN(P3_U2728) );
  INV_X1 U22818 ( .A(n20827), .ZN(n20834) );
  NAND2_X1 U22819 ( .A1(n20971), .A2(n20828), .ZN(n20980) );
  NOR3_X1 U22820 ( .A1(n20829), .A2(n20979), .A3(n20980), .ZN(n20849) );
  NAND2_X1 U22821 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n20849), .ZN(n20844) );
  NOR2_X1 U22822 ( .A1(n20830), .A2(n20844), .ZN(n20847) );
  NAND2_X1 U22823 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n20847), .ZN(n20835) );
  NOR2_X1 U22824 ( .A1(n20831), .A2(n20835), .ZN(n20838) );
  AOI21_X1 U22825 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n20966), .A(n20838), .ZN(
        n20833) );
  OAI222_X1 U22826 ( .A1(n20878), .A2(n20853), .B1(n20834), .B2(n20833), .C1(
        n20990), .C2(n20832), .ZN(P3_U2729) );
  INV_X1 U22827 ( .A(n20835), .ZN(n20842) );
  AOI21_X1 U22828 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n20966), .A(n20842), .ZN(
        n20837) );
  OAI222_X1 U22829 ( .A1(n20839), .A2(n20853), .B1(n20838), .B2(n20837), .C1(
        n20990), .C2(n20836), .ZN(P3_U2730) );
  AOI21_X1 U22830 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n20966), .A(n20847), .ZN(
        n20841) );
  OAI222_X1 U22831 ( .A1(n20843), .A2(n20853), .B1(n20842), .B2(n20841), .C1(
        n20990), .C2(n20840), .ZN(P3_U2731) );
  INV_X1 U22832 ( .A(n20844), .ZN(n20852) );
  AOI21_X1 U22833 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n20966), .A(n20852), .ZN(
        n20846) );
  OAI222_X1 U22834 ( .A1(n20848), .A2(n20853), .B1(n20847), .B2(n20846), .C1(
        n20990), .C2(n20845), .ZN(P3_U2732) );
  AOI21_X1 U22835 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n20966), .A(n20849), .ZN(
        n20851) );
  OAI222_X1 U22836 ( .A1(n20854), .A2(n20853), .B1(n20852), .B2(n20851), .C1(
        n20990), .C2(n20850), .ZN(P3_U2733) );
  NOR2_X2 U22837 ( .A1(n20855), .A2(n20966), .ZN(n20950) );
  NAND2_X1 U22838 ( .A1(n20959), .A2(n20856), .ZN(n20934) );
  AOI22_X1 U22839 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20950), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n20949), .ZN(n20866) );
  NAND2_X1 U22840 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .ZN(n20862) );
  NAND2_X1 U22841 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .ZN(n20861) );
  NAND3_X1 U22842 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .ZN(n20858) );
  NAND4_X1 U22843 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_14__SCAN_IN), 
        .A3(P3_EAX_REG_9__SCAN_IN), .A4(P3_EAX_REG_13__SCAN_IN), .ZN(n20857)
         );
  NAND2_X1 U22844 ( .A1(n20971), .A2(n20951), .ZN(n20889) );
  INV_X1 U22845 ( .A(n20880), .ZN(n20884) );
  NOR2_X1 U22846 ( .A1(n20862), .A2(n20884), .ZN(n20869) );
  NOR3_X1 U22847 ( .A1(n20862), .A2(n20861), .A3(n20860), .ZN(n20874) );
  INV_X1 U22848 ( .A(n20874), .ZN(n20863) );
  NOR2_X1 U22849 ( .A1(n20863), .A2(n20889), .ZN(n20875) );
  INV_X1 U22850 ( .A(n20875), .ZN(n20864) );
  OAI211_X1 U22851 ( .C1(n20869), .C2(P3_EAX_REG_21__SCAN_IN), .A(n20966), .B(
        n20864), .ZN(n20865) );
  OAI211_X1 U22852 ( .C1(n20867), .C2(n20990), .A(n20866), .B(n20865), .ZN(
        P3_U2714) );
  AOI22_X1 U22853 ( .A1(n20880), .A2(P3_EAX_REG_19__SCAN_IN), .B1(
        P3_EAX_REG_20__SCAN_IN), .B2(n20966), .ZN(n20868) );
  OAI22_X1 U22854 ( .A1(n20869), .A2(n20868), .B1(n15956), .B2(n20934), .ZN(
        n20870) );
  AOI21_X1 U22855 ( .B1(BUF2_REG_4__SCAN_IN), .B2(n20950), .A(n20870), .ZN(
        n20871) );
  OAI21_X1 U22856 ( .B1(n20872), .B2(n20990), .A(n20871), .ZN(P3_U2715) );
  INV_X1 U22857 ( .A(n20950), .ZN(n20901) );
  AOI22_X1 U22858 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n20949), .B1(n20978), .B2(
        n20873), .ZN(n20877) );
  NAND3_X1 U22859 ( .A1(n20951), .A2(n20874), .A3(P3_EAX_REG_22__SCAN_IN), 
        .ZN(n20944) );
  OAI211_X1 U22860 ( .C1(n20875), .C2(P3_EAX_REG_22__SCAN_IN), .A(n20966), .B(
        n20944), .ZN(n20876) );
  OAI211_X1 U22861 ( .C1(n20901), .C2(n20878), .A(n20877), .B(n20876), .ZN(
        P3_U2713) );
  AOI22_X1 U22862 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20950), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n20949), .ZN(n20882) );
  NAND2_X1 U22863 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n20880), .ZN(n20879) );
  OAI211_X1 U22864 ( .C1(n20880), .C2(P3_EAX_REG_19__SCAN_IN), .A(n20966), .B(
        n20879), .ZN(n20881) );
  OAI211_X1 U22865 ( .C1(n20883), .C2(n20990), .A(n20882), .B(n20881), .ZN(
        P3_U2716) );
  AOI22_X1 U22866 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20950), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n20949), .ZN(n20886) );
  NOR2_X1 U22867 ( .A1(n20890), .A2(n20889), .ZN(n20888) );
  OAI211_X1 U22868 ( .C1(n20888), .C2(P3_EAX_REG_18__SCAN_IN), .A(n20966), .B(
        n20884), .ZN(n20885) );
  OAI211_X1 U22869 ( .C1(n20887), .C2(n20990), .A(n20886), .B(n20885), .ZN(
        P3_U2717) );
  AOI22_X1 U22870 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20950), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n20949), .ZN(n20893) );
  AOI211_X1 U22871 ( .C1(n20890), .C2(n20889), .A(n20888), .B(n20959), .ZN(
        n20891) );
  INV_X1 U22872 ( .A(n20891), .ZN(n20892) );
  OAI211_X1 U22873 ( .C1(n20894), .C2(n20990), .A(n20893), .B(n20892), .ZN(
        P3_U2718) );
  AOI22_X1 U22874 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n20949), .B1(n20978), .B2(
        n20895), .ZN(n20899) );
  NAND2_X1 U22875 ( .A1(n20942), .A2(n20971), .ZN(n20935) );
  AOI211_X1 U22876 ( .C1(n20896), .C2(n20937), .A(n20902), .B(n20959), .ZN(
        n20897) );
  INV_X1 U22877 ( .A(n20897), .ZN(n20898) );
  OAI211_X1 U22878 ( .C1(n20901), .C2(n20900), .A(n20899), .B(n20898), .ZN(
        P3_U2710) );
  AOI22_X1 U22879 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20950), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n20949), .ZN(n20904) );
  OAI211_X1 U22880 ( .C1(n20902), .C2(P3_EAX_REG_26__SCAN_IN), .A(n20966), .B(
        n20928), .ZN(n20903) );
  OAI211_X1 U22881 ( .C1(n20905), .C2(n20990), .A(n20904), .B(n20903), .ZN(
        P3_U2709) );
  NAND2_X1 U22882 ( .A1(n20927), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n20922) );
  NOR2_X1 U22883 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n20917), .ZN(n20907) );
  NAND2_X1 U22884 ( .A1(n20966), .A2(n20917), .ZN(n20914) );
  OAI21_X1 U22885 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n20980), .A(n20914), .ZN(
        n20906) );
  AOI22_X1 U22886 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n20907), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n20906), .ZN(n20908) );
  OAI21_X1 U22887 ( .B1(n20909), .B2(n20934), .A(n20908), .ZN(P3_U2704) );
  OAI22_X1 U22888 ( .A1(n20911), .A2(n20990), .B1(n20910), .B2(n20934), .ZN(
        n20912) );
  AOI21_X1 U22889 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n20950), .A(n20912), .ZN(
        n20913) );
  OAI221_X1 U22890 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n20917), .C1(n20915), 
        .C2(n20914), .A(n20913), .ZN(P3_U2705) );
  AOI22_X1 U22891 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20950), .B1(n20978), .B2(
        n20916), .ZN(n20920) );
  OAI211_X1 U22892 ( .C1(n20918), .C2(P3_EAX_REG_29__SCAN_IN), .A(n20966), .B(
        n20917), .ZN(n20919) );
  OAI211_X1 U22893 ( .C1(n20934), .C2(n20921), .A(n20920), .B(n20919), .ZN(
        P3_U2706) );
  AOI22_X1 U22894 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20950), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n20949), .ZN(n20924) );
  OAI211_X1 U22895 ( .C1(n20927), .C2(P3_EAX_REG_28__SCAN_IN), .A(n20966), .B(
        n20922), .ZN(n20923) );
  OAI211_X1 U22896 ( .C1(n20925), .C2(n20990), .A(n20924), .B(n20923), .ZN(
        P3_U2707) );
  AOI22_X1 U22897 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20950), .B1(n20978), .B2(
        n20926), .ZN(n20932) );
  AOI211_X1 U22898 ( .C1(n20929), .C2(n20928), .A(n20927), .B(n20959), .ZN(
        n20930) );
  INV_X1 U22899 ( .A(n20930), .ZN(n20931) );
  OAI211_X1 U22900 ( .C1(n20934), .C2(n20933), .A(n20932), .B(n20931), .ZN(
        P3_U2708) );
  AOI22_X1 U22901 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20950), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n20949), .ZN(n20940) );
  OAI21_X1 U22902 ( .B1(n20936), .B2(n20959), .A(n20935), .ZN(n20938) );
  NAND2_X1 U22903 ( .A1(n20938), .A2(n20937), .ZN(n20939) );
  OAI211_X1 U22904 ( .C1(n20941), .C2(n20990), .A(n20940), .B(n20939), .ZN(
        P3_U2711) );
  AOI22_X1 U22905 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20950), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n20949), .ZN(n20948) );
  AOI211_X1 U22906 ( .C1(n20944), .C2(n20943), .A(n20959), .B(n20942), .ZN(
        n20945) );
  AOI21_X1 U22907 ( .B1(n20946), .B2(n20978), .A(n20945), .ZN(n20947) );
  NAND2_X1 U22908 ( .A1(n20948), .A2(n20947), .ZN(P3_U2712) );
  AOI22_X1 U22909 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20950), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n20949), .ZN(n20955) );
  AOI211_X1 U22910 ( .C1(n20965), .C2(n20952), .A(n20959), .B(n20951), .ZN(
        n20953) );
  INV_X1 U22911 ( .A(n20953), .ZN(n20954) );
  OAI211_X1 U22912 ( .C1(n20956), .C2(n20990), .A(n20955), .B(n20954), .ZN(
        P3_U2719) );
  NAND2_X1 U22913 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n20957), .ZN(n20963) );
  AOI22_X1 U22914 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20986), .B1(n20978), .B2(
        n20958), .ZN(n20962) );
  OR3_X1 U22915 ( .A1(n20960), .A2(n20959), .A3(n20967), .ZN(n20961) );
  OAI211_X1 U22916 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n20963), .A(n20962), .B(
        n20961), .ZN(P3_U2721) );
  AOI22_X1 U22917 ( .A1(n20978), .A2(n20964), .B1(BUF2_REG_15__SCAN_IN), .B2(
        n20986), .ZN(n20969) );
  OAI211_X1 U22918 ( .C1(n20967), .C2(P3_EAX_REG_15__SCAN_IN), .A(n20966), .B(
        n20965), .ZN(n20968) );
  NAND2_X1 U22919 ( .A1(n20969), .A2(n20968), .ZN(P3_U2720) );
  NAND3_X1 U22920 ( .A1(n20971), .A2(n20970), .A3(P3_EAX_REG_7__SCAN_IN), .ZN(
        n20976) );
  AOI22_X1 U22921 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20986), .B1(n20978), .B2(
        n20972), .ZN(n20973) );
  OAI221_X1 U22922 ( .B1(P3_EAX_REG_8__SCAN_IN), .B2(n20976), .C1(n20975), 
        .C2(n20974), .A(n20973), .ZN(P3_U2727) );
  AOI22_X1 U22923 ( .A1(n20986), .A2(BUF2_REG_1__SCAN_IN), .B1(n20978), .B2(
        n20977), .ZN(n20984) );
  NOR2_X1 U22924 ( .A1(n20979), .A2(n20980), .ZN(n20982) );
  NOR2_X1 U22925 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n20980), .ZN(n20987) );
  OAI22_X1 U22926 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n20982), .B1(n20987), .B2(
        n20981), .ZN(n20983) );
  NAND2_X1 U22927 ( .A1(n20984), .A2(n20983), .ZN(P3_U2734) );
  AOI22_X1 U22928 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20986), .B1(
        P3_EAX_REG_0__SCAN_IN), .B2(n20985), .ZN(n20989) );
  INV_X1 U22929 ( .A(n20987), .ZN(n20988) );
  OAI211_X1 U22930 ( .C1(n20991), .C2(n20990), .A(n20989), .B(n20988), .ZN(
        P3_U2735) );
  NAND2_X1 U22931 ( .A1(n21217), .A2(n20992), .ZN(n20994) );
  AOI22_X1 U22932 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21231), .B1(
        n20994), .B2(n21020), .ZN(n21451) );
  INV_X1 U22933 ( .A(n21451), .ZN(n21448) );
  AOI222_X1 U22934 ( .A1(n21071), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n21448), 
        .B2(n21036), .C1(n21020), .C2(n21490), .ZN(n20993) );
  AOI22_X1 U22935 ( .A1(n21040), .A2(n21020), .B1(n20993), .B2(n21038), .ZN(
        P3_U3290) );
  INV_X1 U22936 ( .A(n21231), .ZN(n21427) );
  AOI21_X1 U22937 ( .B1(n21427), .B2(n21020), .A(n21372), .ZN(n21026) );
  AOI22_X1 U22938 ( .A1(n20998), .A2(n20994), .B1(n21026), .B2(n21001), .ZN(
        n21453) );
  INV_X1 U22939 ( .A(n21453), .ZN(n20999) );
  INV_X1 U22940 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n20996) );
  AOI22_X1 U22941 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20996), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n20995), .ZN(n21011) );
  NOR2_X1 U22942 ( .A1(n20997), .A2(n21071), .ZN(n21014) );
  AOI222_X1 U22943 ( .A1(n20999), .A2(n21036), .B1(n20998), .B2(n21490), .C1(
        n21011), .C2(n21014), .ZN(n21000) );
  AOI22_X1 U22944 ( .A1(n21040), .A2(n21001), .B1(n21000), .B2(n21038), .ZN(
        P3_U3289) );
  OAI211_X1 U22945 ( .C1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n21026), .B(n21028), .ZN(
        n21009) );
  OAI22_X1 U22946 ( .A1(n21005), .A2(n21004), .B1(n21003), .B2(n21002), .ZN(
        n21034) );
  NOR2_X1 U22947 ( .A1(n20344), .A2(n21006), .ZN(n21016) );
  OAI21_X1 U22948 ( .B1(n21007), .B2(n21034), .A(n21016), .ZN(n21008) );
  OAI211_X1 U22949 ( .C1(n21438), .C2(n21010), .A(n21009), .B(n21008), .ZN(
        n21456) );
  INV_X1 U22950 ( .A(n21011), .ZN(n21015) );
  INV_X1 U22951 ( .A(n21012), .ZN(n21013) );
  AOI222_X1 U22952 ( .A1(n21456), .A2(n21036), .B1(n21015), .B2(n21014), .C1(
        n21013), .C2(n21490), .ZN(n21018) );
  AOI22_X1 U22953 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n21040), .B1(
        n21490), .B2(n21016), .ZN(n21017) );
  OAI21_X1 U22954 ( .B1(n21040), .B2(n21018), .A(n21017), .ZN(P3_U3288) );
  INV_X1 U22955 ( .A(n21019), .ZN(n21037) );
  NAND2_X1 U22956 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21020), .ZN(
        n21024) );
  OAI211_X1 U22957 ( .C1(n20344), .C2(n21022), .A(n21368), .B(n21021), .ZN(
        n21023) );
  OAI22_X1 U22958 ( .A1(n21025), .A2(n21024), .B1(n10956), .B2(n21023), .ZN(
        n21032) );
  INV_X1 U22959 ( .A(n21026), .ZN(n21027) );
  OAI33_X1 U22960 ( .A1(n21030), .A2(n21029), .A3(n21461), .B1(n21028), .B2(
        n21027), .B3(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n21031) );
  AOI211_X1 U22961 ( .C1(n21034), .C2(n21033), .A(n21032), .B(n21031), .ZN(
        n21460) );
  INV_X1 U22962 ( .A(n21460), .ZN(n21035) );
  AOI22_X1 U22963 ( .A1(n21490), .A2(n21037), .B1(n21036), .B2(n21035), .ZN(
        n21039) );
  AOI22_X1 U22964 ( .A1(n21040), .A2(n21461), .B1(n21039), .B2(n21038), .ZN(
        P3_U3285) );
  AOI22_X1 U22965 ( .A1(n21345), .A2(n21362), .B1(n21343), .B2(n21041), .ZN(
        n21153) );
  OAI21_X1 U22966 ( .B1(n21153), .B2(n21043), .A(n21042), .ZN(n21221) );
  NAND2_X1 U22967 ( .A1(n21403), .A2(n21221), .ZN(n21358) );
  AOI21_X1 U22968 ( .B1(n21050), .B2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n21427), .ZN(n21044) );
  AOI21_X1 U22969 ( .B1(n21368), .B2(n21045), .A(n21044), .ZN(n21339) );
  AOI22_X1 U22970 ( .A1(n21345), .A2(n21047), .B1(n21343), .B2(n21046), .ZN(
        n21048) );
  OAI211_X1 U22971 ( .C1(n21215), .C2(n21049), .A(n21339), .B(n21048), .ZN(
        n21219) );
  NAND2_X1 U22972 ( .A1(n21422), .A2(n21071), .ZN(n21365) );
  OAI211_X1 U22973 ( .C1(n21217), .C2(n21050), .A(n21403), .B(n21365), .ZN(
        n21340) );
  AOI211_X1 U22974 ( .C1(n21422), .C2(n21051), .A(n21219), .B(n21340), .ZN(
        n21052) );
  NOR3_X1 U22975 ( .A1(n21401), .A2(n21052), .A3(n21220), .ZN(n21053) );
  AOI21_X1 U22976 ( .B1(n21432), .B2(n21054), .A(n21053), .ZN(n21056) );
  OAI211_X1 U22977 ( .C1(n21057), .C2(n21358), .A(n21056), .B(n21055), .ZN(
        P3_U2841) );
  NOR2_X1 U22978 ( .A1(n21368), .A2(n21422), .ZN(n21353) );
  AOI221_X1 U22979 ( .B1(n21353), .B2(n21071), .C1(n21427), .C2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n21430), .ZN(n21058) );
  AOI221_X1 U22980 ( .B1(n21271), .B2(n21060), .C1(n21131), .C2(n21059), .A(
        n21058), .ZN(n21062) );
  NAND2_X1 U22981 ( .A1(n21401), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n21061) );
  OAI211_X1 U22982 ( .C1(n21383), .C2(n21071), .A(n21062), .B(n21061), .ZN(
        P3_U2862) );
  AOI22_X1 U22983 ( .A1(n21401), .A2(P3_REIP_REG_1__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n21410), .ZN(n21069) );
  NOR2_X1 U22984 ( .A1(n21392), .A2(n21063), .ZN(n21065) );
  NOR2_X1 U22985 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21353), .ZN(
        n21064) );
  MUX2_X1 U22986 ( .A(n21065), .B(n21064), .S(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n21067) );
  AOI22_X1 U22987 ( .A1(n21403), .A2(n21067), .B1(n21131), .B2(n21066), .ZN(
        n21068) );
  OAI211_X1 U22988 ( .C1(n21070), .C2(n21239), .A(n21069), .B(n21068), .ZN(
        P3_U2861) );
  NOR2_X1 U22989 ( .A1(n21071), .A2(n21089), .ZN(n21087) );
  NOR2_X1 U22990 ( .A1(n21438), .A2(n21086), .ZN(n21073) );
  AOI211_X1 U22991 ( .C1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n21365), .A(
        n21372), .B(n21083), .ZN(n21072) );
  AOI211_X1 U22992 ( .C1(n21368), .C2(n21087), .A(n21073), .B(n21072), .ZN(
        n21075) );
  NAND3_X1 U22993 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21085), .A3(
        n21083), .ZN(n21074) );
  OAI211_X1 U22994 ( .C1(n21076), .C2(n21437), .A(n21075), .B(n21074), .ZN(
        n21080) );
  AOI21_X1 U22995 ( .B1(n21078), .B2(n21077), .A(n18447), .ZN(n21079) );
  AOI22_X1 U22996 ( .A1(n21403), .A2(n21080), .B1(n21131), .B2(n21079), .ZN(
        n21082) );
  OAI211_X1 U22997 ( .C1(n21383), .C2(n21083), .A(n21082), .B(n21081), .ZN(
        P3_U2860) );
  INV_X1 U22998 ( .A(n21089), .ZN(n21084) );
  AOI22_X1 U22999 ( .A1(n21368), .A2(n21086), .B1(n21085), .B2(n21084), .ZN(
        n21134) );
  OAI22_X1 U23000 ( .A1(n21217), .A2(n21087), .B1(n21438), .B2(n21086), .ZN(
        n21088) );
  AOI211_X1 U23001 ( .C1(n21231), .C2(n21089), .A(n21097), .B(n21088), .ZN(
        n21101) );
  AOI211_X1 U23002 ( .C1(n21134), .C2(n21097), .A(n21101), .B(n21430), .ZN(
        n21092) );
  OAI22_X1 U23003 ( .A1(n21379), .A2(n21090), .B1(n21097), .B2(n21383), .ZN(
        n21091) );
  AOI211_X1 U23004 ( .C1(n21093), .C2(n21131), .A(n21092), .B(n21091), .ZN(
        n21094) );
  OAI21_X1 U23005 ( .B1(n21239), .B2(n21095), .A(n21094), .ZN(P3_U2859) );
  INV_X1 U23006 ( .A(n21096), .ZN(n21107) );
  NOR3_X1 U23007 ( .A1(n21134), .A2(n21097), .A3(n21430), .ZN(n21099) );
  AOI221_X1 U23008 ( .B1(n21410), .B2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(
        n21099), .C2(n21100), .A(n21098), .ZN(n21106) );
  NOR3_X1 U23009 ( .A1(n21392), .A2(n21101), .A3(n21100), .ZN(n21104) );
  INV_X1 U23010 ( .A(n21102), .ZN(n21442) );
  OAI221_X1 U23011 ( .B1(n21104), .B2(n21103), .C1(n21104), .C2(n21442), .A(
        n21403), .ZN(n21105) );
  OAI211_X1 U23012 ( .C1(n21107), .C2(n21239), .A(n21106), .B(n21105), .ZN(
        P3_U2858) );
  OR2_X1 U23013 ( .A1(n21430), .A2(n21134), .ZN(n21120) );
  NOR2_X1 U23014 ( .A1(n21108), .A2(n21120), .ZN(n21114) );
  NAND2_X1 U23015 ( .A1(n21368), .A2(n21109), .ZN(n21110) );
  OAI211_X1 U23016 ( .C1(n21372), .C2(n21111), .A(n21110), .B(n21365), .ZN(
        n21112) );
  AOI21_X1 U23017 ( .B1(n21403), .B2(n21112), .A(n21410), .ZN(n21113) );
  INV_X1 U23018 ( .A(n21113), .ZN(n21121) );
  MUX2_X1 U23019 ( .A(n21114), .B(n21121), .S(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(n21115) );
  AOI21_X1 U23020 ( .B1(n21131), .B2(n21116), .A(n21115), .ZN(n21118) );
  NAND2_X1 U23021 ( .A1(n21401), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n21117) );
  OAI211_X1 U23022 ( .C1(n21119), .C2(n21239), .A(n21118), .B(n21117), .ZN(
        P3_U2857) );
  NOR2_X1 U23023 ( .A1(n21133), .A2(n21120), .ZN(n21122) );
  MUX2_X1 U23024 ( .A(n21122), .B(n21121), .S(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .Z(n21123) );
  AOI21_X1 U23025 ( .B1(n21131), .B2(n21124), .A(n21123), .ZN(n21126) );
  NAND2_X1 U23026 ( .A1(n21401), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n21125) );
  OAI211_X1 U23027 ( .C1(n21127), .C2(n21239), .A(n21126), .B(n21125), .ZN(
        P3_U2856) );
  OAI22_X1 U23028 ( .A1(n21428), .A2(n21128), .B1(n21135), .B2(n21383), .ZN(
        n21129) );
  AOI21_X1 U23029 ( .B1(n21131), .B2(n21130), .A(n21129), .ZN(n21140) );
  NOR3_X1 U23030 ( .A1(n21134), .A2(n21133), .A3(n21132), .ZN(n21152) );
  INV_X1 U23031 ( .A(n21372), .ZN(n21421) );
  AOI21_X1 U23032 ( .B1(n21421), .B2(n21136), .A(n21135), .ZN(n21137) );
  OAI211_X1 U23033 ( .C1(n21138), .C2(n21438), .A(n21137), .B(n21365), .ZN(
        n21142) );
  OAI211_X1 U23034 ( .C1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n21152), .A(
        n21403), .B(n21142), .ZN(n21139) );
  OAI211_X1 U23035 ( .C1(n21141), .C2(n21239), .A(n21140), .B(n21139), .ZN(
        P3_U2855) );
  NAND3_X1 U23036 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21334), .A3(
        n21142), .ZN(n21144) );
  NAND3_X1 U23037 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n21152), .A3(
        n21423), .ZN(n21143) );
  OAI211_X1 U23038 ( .C1(n21145), .C2(n21437), .A(n21144), .B(n21143), .ZN(
        n21146) );
  AOI21_X1 U23039 ( .B1(n21345), .B2(n21147), .A(n21146), .ZN(n21151) );
  AOI22_X1 U23040 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21410), .B1(
        n21432), .B2(n21148), .ZN(n21150) );
  OAI211_X1 U23041 ( .C1(n21151), .C2(n21430), .A(n21150), .B(n21149), .ZN(
        P3_U2854) );
  NAND3_X1 U23042 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n21152), .ZN(n21206) );
  NAND2_X1 U23043 ( .A1(n21153), .A2(n21206), .ZN(n21174) );
  NAND2_X1 U23044 ( .A1(n21403), .A2(n21174), .ZN(n21436) );
  NAND2_X1 U23045 ( .A1(n21361), .A2(n21437), .ZN(n21371) );
  INV_X1 U23046 ( .A(n21371), .ZN(n21157) );
  NOR2_X1 U23047 ( .A1(n21362), .A2(n21361), .ZN(n21154) );
  AND2_X1 U23048 ( .A1(n21194), .A2(n21368), .ZN(n21165) );
  AOI211_X1 U23049 ( .C1(n21155), .C2(n21343), .A(n21154), .B(n21165), .ZN(
        n21425) );
  INV_X1 U23050 ( .A(n21195), .ZN(n21413) );
  NAND2_X1 U23051 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21413), .ZN(
        n21420) );
  OAI21_X1 U23052 ( .B1(n21435), .B2(n21420), .A(n21422), .ZN(n21156) );
  OAI211_X1 U23053 ( .C1(n21158), .C2(n21157), .A(n21425), .B(n21156), .ZN(
        n21409) );
  OR2_X1 U23054 ( .A1(n21438), .A2(n21175), .ZN(n21182) );
  OAI221_X1 U23055 ( .B1(n21427), .B2(n21158), .C1(n21427), .C2(n21413), .A(
        n21182), .ZN(n21167) );
  AOI211_X1 U23056 ( .C1(n21422), .C2(n21412), .A(n21409), .B(n21167), .ZN(
        n21159) );
  OAI21_X1 U23057 ( .B1(n21159), .B2(n21430), .A(n21383), .ZN(n21161) );
  AOI22_X1 U23058 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n21161), .B1(
        n21432), .B2(n21160), .ZN(n21163) );
  OAI211_X1 U23059 ( .C1(n21164), .C2(n21436), .A(n21163), .B(n21162), .ZN(
        P3_U2851) );
  AOI221_X1 U23060 ( .B1(n21166), .B2(n21422), .C1(n21420), .C2(n21422), .A(
        n21165), .ZN(n21181) );
  AOI21_X1 U23061 ( .B1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n21427), .ZN(n21172) );
  AOI21_X1 U23062 ( .B1(n21343), .B2(n21168), .A(n21167), .ZN(n21169) );
  OAI21_X1 U23063 ( .B1(n21170), .B2(n21361), .A(n21169), .ZN(n21171) );
  NOR2_X1 U23064 ( .A1(n21172), .A2(n21171), .ZN(n21402) );
  NAND3_X1 U23065 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n21181), .A3(
        n21402), .ZN(n21173) );
  OAI221_X1 U23066 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n21175), 
        .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n21174), .A(n21173), .ZN(
        n21179) );
  AOI22_X1 U23067 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n21410), .B1(
        n21432), .B2(n21176), .ZN(n21178) );
  OAI211_X1 U23068 ( .C1(n21430), .C2(n21179), .A(n21178), .B(n21177), .ZN(
        P3_U2850) );
  NOR3_X1 U23069 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n21196), .A3(
        n21206), .ZN(n21188) );
  NAND2_X1 U23070 ( .A1(n21180), .A2(n21413), .ZN(n21184) );
  OAI21_X1 U23071 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n21438), .A(
        n21181), .ZN(n21405) );
  OAI21_X1 U23072 ( .B1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n21353), .A(
        n21182), .ZN(n21183) );
  AOI211_X1 U23073 ( .C1(n21231), .C2(n21184), .A(n21405), .B(n21183), .ZN(
        n21186) );
  OAI22_X1 U23074 ( .A1(n21186), .A2(n13871), .B1(n21437), .B2(n21185), .ZN(
        n21187) );
  AOI211_X1 U23075 ( .C1(n21189), .C2(n21345), .A(n21188), .B(n21187), .ZN(
        n21193) );
  AOI22_X1 U23076 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n21410), .B1(
        n21432), .B2(n21190), .ZN(n21192) );
  OAI211_X1 U23077 ( .C1(n21193), .C2(n21430), .A(n21192), .B(n21191), .ZN(
        P3_U2848) );
  NOR2_X1 U23078 ( .A1(n21374), .A2(n21194), .ZN(n21363) );
  NOR3_X1 U23079 ( .A1(n13871), .A2(n21196), .A3(n21195), .ZN(n21197) );
  OAI21_X1 U23080 ( .B1(n21217), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n21197), .ZN(n21198) );
  OAI21_X1 U23081 ( .B1(n21231), .B2(n21422), .A(n21198), .ZN(n21199) );
  OAI211_X1 U23082 ( .C1(n21363), .C2(n21438), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n21199), .ZN(n21204) );
  OAI22_X1 U23083 ( .A1(n21207), .A2(n21361), .B1(n21360), .B2(n21437), .ZN(
        n21394) );
  AOI221_X1 U23084 ( .B1(n21204), .B2(n21403), .C1(n21394), .C2(n21403), .A(
        n21410), .ZN(n21214) );
  NOR3_X1 U23085 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21200), .A3(
        n21239), .ZN(n21201) );
  AOI211_X1 U23086 ( .C1(n21432), .C2(n21203), .A(n21202), .B(n21201), .ZN(
        n21212) );
  INV_X1 U23087 ( .A(n21204), .ZN(n21391) );
  NOR3_X1 U23088 ( .A1(n21391), .A2(n21206), .A3(n21205), .ZN(n21210) );
  NOR2_X1 U23089 ( .A1(n21207), .A2(n21361), .ZN(n21209) );
  OAI221_X1 U23090 ( .B1(n21210), .B2(n21209), .C1(n21210), .C2(n21208), .A(
        n21403), .ZN(n21211) );
  OAI211_X1 U23091 ( .C1(n21214), .C2(n21213), .A(n21212), .B(n21211), .ZN(
        P3_U2847) );
  INV_X1 U23092 ( .A(n21215), .ZN(n21411) );
  NAND2_X1 U23093 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n21216), .ZN(
        n21230) );
  INV_X1 U23094 ( .A(n21230), .ZN(n21218) );
  AOI21_X1 U23095 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21218), .A(
        n21217), .ZN(n21229) );
  AOI211_X1 U23096 ( .C1(n21411), .C2(n21220), .A(n21229), .B(n21219), .ZN(
        n21223) );
  NAND2_X1 U23097 ( .A1(n21222), .A2(n21221), .ZN(n21330) );
  AOI221_X1 U23098 ( .B1(n21223), .B2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), 
        .C1(n21330), .C2(n21257), .A(n21430), .ZN(n21224) );
  AOI21_X1 U23099 ( .B1(n21225), .B2(n21432), .A(n21224), .ZN(n21227) );
  OAI211_X1 U23100 ( .C1(n21383), .C2(n21257), .A(n21227), .B(n21226), .ZN(
        P3_U2840) );
  NAND2_X1 U23101 ( .A1(n21228), .A2(n21247), .ZN(n21234) );
  AOI21_X1 U23102 ( .B1(n21231), .B2(n21230), .A(n21229), .ZN(n21322) );
  INV_X1 U23103 ( .A(n21322), .ZN(n21232) );
  AOI211_X1 U23104 ( .C1(n21334), .C2(n21233), .A(n21323), .B(n21232), .ZN(
        n21250) );
  OAI22_X1 U23105 ( .A1(n21235), .A2(n21234), .B1(n21250), .B2(n21247), .ZN(
        n21236) );
  AOI21_X1 U23106 ( .B1(n21345), .B2(n21237), .A(n21236), .ZN(n21240) );
  OAI22_X1 U23107 ( .A1(n21240), .A2(n21430), .B1(n21239), .B2(n21238), .ZN(
        n21241) );
  AOI21_X1 U23108 ( .B1(n21432), .B2(n21242), .A(n21241), .ZN(n21244) );
  OAI211_X1 U23109 ( .C1(n21383), .C2(n21247), .A(n21244), .B(n21243), .ZN(
        P3_U2837) );
  AOI22_X1 U23110 ( .A1(n21401), .A2(P3_REIP_REG_26__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n21410), .ZN(n21255) );
  INV_X1 U23111 ( .A(n21330), .ZN(n21253) );
  NOR2_X1 U23112 ( .A1(n21245), .A2(n21361), .ZN(n21261) );
  AOI211_X1 U23113 ( .C1(n21334), .C2(n21247), .A(n21261), .B(n21246), .ZN(
        n21249) );
  NAND2_X1 U23114 ( .A1(n21271), .A2(n21248), .ZN(n21262) );
  OAI221_X1 U23115 ( .B1(n21430), .B2(n21250), .C1(n21430), .C2(n21249), .A(
        n21262), .ZN(n21251) );
  OAI221_X1 U23116 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n21253), 
        .C1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n21252), .A(n21251), .ZN(
        n21254) );
  OAI211_X1 U23117 ( .C1(n21256), .C2(n21337), .A(n21255), .B(n21254), .ZN(
        P3_U2836) );
  NOR2_X1 U23118 ( .A1(n21330), .A2(n21257), .ZN(n21325) );
  NAND2_X1 U23119 ( .A1(n21325), .A2(n21259), .ZN(n21307) );
  AND2_X1 U23120 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n21258), .ZN(
        n21273) );
  OAI211_X1 U23121 ( .C1(n21372), .C2(n21259), .A(n21273), .B(n21322), .ZN(
        n21260) );
  OAI21_X1 U23122 ( .B1(n21261), .B2(n21260), .A(n21403), .ZN(n21263) );
  AOI22_X1 U23123 ( .A1(n21307), .A2(n21306), .B1(n21263), .B2(n21262), .ZN(
        n21264) );
  AOI211_X1 U23124 ( .C1(n21432), .C2(n21266), .A(n21265), .B(n21264), .ZN(
        n21267) );
  OAI21_X1 U23125 ( .B1(n21306), .B2(n21383), .A(n21267), .ZN(P3_U2835) );
  AOI221_X1 U23126 ( .B1(n21361), .B2(n21270), .C1(n21269), .C2(n21270), .A(
        n21268), .ZN(n21272) );
  AOI22_X1 U23127 ( .A1(n21403), .A2(n21272), .B1(n11245), .B2(n21271), .ZN(
        n21289) );
  OAI22_X1 U23128 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n21353), .B1(
        n21273), .B2(n21438), .ZN(n21281) );
  NAND2_X1 U23129 ( .A1(n21275), .A2(n21274), .ZN(n21276) );
  AOI22_X1 U23130 ( .A1(n21345), .A2(n21277), .B1(n21343), .B2(n21276), .ZN(
        n21285) );
  OAI211_X1 U23131 ( .C1(n21427), .C2(n21279), .A(n21278), .B(n21285), .ZN(
        n21280) );
  AOI221_X1 U23132 ( .B1(n21281), .B2(n21403), .C1(n21280), .C2(n21403), .A(
        n21410), .ZN(n21284) );
  AOI22_X1 U23133 ( .A1(n21401), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n21432), 
        .B2(n21282), .ZN(n21283) );
  OAI221_X1 U23134 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n21289), 
        .C1(n21288), .C2(n21284), .A(n21283), .ZN(P3_U2833) );
  NAND2_X1 U23135 ( .A1(n21286), .A2(n21285), .ZN(n21290) );
  INV_X1 U23136 ( .A(n21290), .ZN(n21287) );
  OAI21_X1 U23137 ( .B1(n21287), .B2(n21430), .A(n21383), .ZN(n21292) );
  NOR2_X1 U23138 ( .A1(n21289), .A2(n21288), .ZN(n21291) );
  AOI22_X1 U23139 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n21292), .B1(
        n21291), .B2(n21290), .ZN(n21294) );
  OAI211_X1 U23140 ( .C1(n21295), .C2(n21337), .A(n21294), .B(n21293), .ZN(
        P3_U2832) );
  NOR2_X1 U23141 ( .A1(n11245), .A2(n21437), .ZN(n21298) );
  AOI21_X1 U23142 ( .B1(n21300), .B2(n21299), .A(n21298), .ZN(n21305) );
  AOI211_X1 U23143 ( .C1(n21411), .C2(n21306), .A(n21410), .B(n21302), .ZN(
        n21303) );
  NAND3_X1 U23144 ( .A1(n21305), .A2(n21304), .A3(n21303), .ZN(n21313) );
  NAND2_X1 U23145 ( .A1(n21309), .A2(n21403), .ZN(n21311) );
  INV_X1 U23146 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n21310) );
  NAND2_X1 U23147 ( .A1(n21311), .A2(n21310), .ZN(n21312) );
  NAND2_X1 U23148 ( .A1(n21313), .A2(n21312), .ZN(n21318) );
  OR3_X1 U23149 ( .A1(n21315), .A2(n21337), .A3(n21314), .ZN(n21316) );
  OAI221_X1 U23150 ( .B1(n21401), .B2(n21318), .C1(n21379), .C2(n21317), .A(
        n21316), .ZN(P3_U2834) );
  AOI22_X1 U23151 ( .A1(n21345), .A2(n21320), .B1(n21343), .B2(n21319), .ZN(
        n21321) );
  NAND3_X1 U23152 ( .A1(n21322), .A2(n21321), .A3(n21383), .ZN(n21333) );
  NOR2_X1 U23153 ( .A1(n21333), .A2(n21323), .ZN(n21324) );
  AOI21_X1 U23154 ( .B1(n21324), .B2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n21401), .ZN(n21332) );
  OAI221_X1 U23155 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n21325), 
        .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n21383), .A(n21332), .ZN(
        n21326) );
  OAI211_X1 U23156 ( .C1(n21328), .C2(n21337), .A(n21327), .B(n21326), .ZN(
        P3_U2839) );
  NOR4_X1 U23157 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n21330), .A3(
        n21430), .A4(n21329), .ZN(n21331) );
  AOI21_X1 U23158 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n21401), .A(n21331), 
        .ZN(n21336) );
  OAI211_X1 U23159 ( .C1(n21334), .C2(n21333), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n21332), .ZN(n21335) );
  OAI211_X1 U23160 ( .C1(n21338), .C2(n21337), .A(n21336), .B(n21335), .ZN(
        P3_U2838) );
  INV_X1 U23161 ( .A(n21339), .ZN(n21341) );
  AOI211_X1 U23162 ( .C1(n21343), .C2(n21342), .A(n21341), .B(n21340), .ZN(
        n21347) );
  NAND2_X1 U23163 ( .A1(n21345), .A2(n21344), .ZN(n21346) );
  AOI21_X1 U23164 ( .B1(n21347), .B2(n21346), .A(n21401), .ZN(n21355) );
  AOI22_X1 U23165 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n21355), .B1(
        n21432), .B2(n21348), .ZN(n21350) );
  OAI211_X1 U23166 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n21358), .A(
        n21350), .B(n21349), .ZN(P3_U2843) );
  AOI22_X1 U23167 ( .A1(n21401), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n21432), 
        .B2(n21351), .ZN(n21357) );
  NOR3_X1 U23168 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n21353), .A3(
        n21352), .ZN(n21354) );
  OAI21_X1 U23169 ( .B1(n21355), .B2(n21354), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n21356) );
  OAI211_X1 U23170 ( .C1(n21359), .C2(n21358), .A(n21357), .B(n21356), .ZN(
        P3_U2842) );
  OAI211_X1 U23171 ( .C1(n21362), .C2(n21361), .A(n21364), .B(n21360), .ZN(
        n21370) );
  NAND2_X1 U23172 ( .A1(n21364), .A2(n21363), .ZN(n21369) );
  NAND4_X1 U23173 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n21366), .A3(
        n21413), .A4(n21365), .ZN(n21367) );
  AOI222_X1 U23174 ( .A1(n21371), .A2(n21370), .B1(n21369), .B2(n21368), .C1(
        n21367), .C2(n21421), .ZN(n21384) );
  OAI211_X1 U23175 ( .C1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n21372), .A(
        n21403), .B(n21384), .ZN(n21373) );
  NAND2_X1 U23176 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n21373), .ZN(
        n21380) );
  NOR2_X1 U23177 ( .A1(n21374), .A2(n21436), .ZN(n21382) );
  AOI22_X1 U23178 ( .A1(n21432), .A2(n21376), .B1(n21375), .B2(n21382), .ZN(
        n21377) );
  OAI221_X1 U23179 ( .B1(n21401), .B2(n21380), .C1(n21379), .C2(n21378), .A(
        n21377), .ZN(P3_U2844) );
  INV_X1 U23180 ( .A(n21381), .ZN(n21390) );
  INV_X1 U23181 ( .A(n21382), .ZN(n21399) );
  OAI21_X1 U23182 ( .B1(n21384), .B2(n21430), .A(n21383), .ZN(n21386) );
  AOI22_X1 U23183 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n21386), .B1(
        n21432), .B2(n21385), .ZN(n21389) );
  INV_X1 U23184 ( .A(n21387), .ZN(n21388) );
  OAI211_X1 U23185 ( .C1(n21390), .C2(n21399), .A(n21389), .B(n21388), .ZN(
        P3_U2845) );
  OAI21_X1 U23186 ( .B1(n21392), .B2(n21391), .A(n21403), .ZN(n21393) );
  OAI21_X1 U23187 ( .B1(n21394), .B2(n21393), .A(n21428), .ZN(n21397) );
  AOI22_X1 U23188 ( .A1(n21401), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n21432), 
        .B2(n21395), .ZN(n21396) );
  OAI221_X1 U23189 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n21399), 
        .C1(n21398), .C2(n21397), .A(n21396), .ZN(P3_U2846) );
  AOI22_X1 U23190 ( .A1(n21401), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n21432), 
        .B2(n21400), .ZN(n21407) );
  NAND2_X1 U23191 ( .A1(n21403), .A2(n21402), .ZN(n21404) );
  OAI211_X1 U23192 ( .C1(n21405), .C2(n21404), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n21428), .ZN(n21406) );
  OAI211_X1 U23193 ( .C1(n21436), .C2(n21408), .A(n21407), .B(n21406), .ZN(
        P3_U2849) );
  NAND2_X1 U23194 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n21412), .ZN(
        n21419) );
  AOI211_X1 U23195 ( .C1(n21411), .C2(n21435), .A(n21410), .B(n21409), .ZN(
        n21414) );
  AOI221_X1 U23196 ( .B1(n21427), .B2(n21414), .C1(n21413), .C2(n21414), .A(
        n21412), .ZN(n21415) );
  AOI22_X1 U23197 ( .A1(n21416), .A2(n21432), .B1(n21415), .B2(n21428), .ZN(
        n21418) );
  OAI211_X1 U23198 ( .C1(n21436), .C2(n21419), .A(n21418), .B(n21417), .ZN(
        P3_U2852) );
  OAI211_X1 U23199 ( .C1(n21423), .C2(n21422), .A(n21421), .B(n21420), .ZN(
        n21424) );
  OAI211_X1 U23200 ( .C1(n21427), .C2(n21426), .A(n21425), .B(n21424), .ZN(
        n21429) );
  OAI21_X1 U23201 ( .B1(n21430), .B2(n21429), .A(n21428), .ZN(n21434) );
  AOI22_X1 U23202 ( .A1(n21401), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n21432), 
        .B2(n21431), .ZN(n21433) );
  OAI221_X1 U23203 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21436), .C1(
        n21435), .C2(n21434), .A(n21433), .ZN(P3_U2853) );
  NAND2_X1 U23204 ( .A1(n21876), .A2(n21489), .ZN(n21484) );
  NAND2_X1 U23205 ( .A1(n21438), .A2(n21437), .ZN(n21444) );
  OR2_X1 U23206 ( .A1(n21440), .A2(n21439), .ZN(n21441) );
  AOI222_X1 U23207 ( .A1(n21445), .A2(n21444), .B1(n21443), .B2(n21442), .C1(
        n21441), .C2(n21471), .ZN(n21503) );
  AOI211_X1 U23208 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n11085), .A(
        n21447), .B(n21446), .ZN(n21474) );
  INV_X1 U23209 ( .A(n11085), .ZN(n21459) );
  NOR3_X1 U23210 ( .A1(n21450), .A2(n21449), .A3(n21448), .ZN(n21452) );
  OAI22_X1 U23211 ( .A1(n21453), .A2(n21452), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n21451), .ZN(n21455) );
  AOI21_X1 U23212 ( .B1(n21459), .B2(n21455), .A(n21454), .ZN(n21458) );
  AOI22_X1 U23213 ( .A1(n11085), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n21456), .B2(n21459), .ZN(n21463) );
  OR2_X1 U23214 ( .A1(n21463), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n21457) );
  AOI221_X1 U23215 ( .B1(n21458), .B2(n21457), .C1(n21463), .C2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21467) );
  AOI22_X1 U23216 ( .A1(n11085), .A2(n21461), .B1(n21460), .B2(n21459), .ZN(
        n21466) );
  OAI21_X1 U23217 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n21463), .ZN(n21464) );
  AOI222_X1 U23218 ( .A1(n21467), .A2(n21466), .B1(n21467), .B2(n21465), .C1(
        n21466), .C2(n21464), .ZN(n21473) );
  INV_X1 U23219 ( .A(n21468), .ZN(n21470) );
  NOR3_X1 U23220 ( .A1(n21471), .A2(n21470), .A3(n21469), .ZN(n21501) );
  OAI21_X1 U23221 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(P3_MORE_REG_SCAN_IN), .A(
        n21501), .ZN(n21472) );
  OAI211_X1 U23222 ( .C1(n21477), .C2(n21476), .A(n21475), .B(n21499), .ZN(
        n21487) );
  OAI21_X1 U23223 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n21478), .A(n21487), 
        .ZN(n21493) );
  INV_X1 U23224 ( .A(n21493), .ZN(n21480) );
  NAND3_X1 U23225 ( .A1(n21481), .A2(n21480), .A3(n21479), .ZN(n21482) );
  NAND4_X1 U23226 ( .A1(n21485), .A2(n21484), .A3(n21483), .A4(n21482), .ZN(
        P3_U2997) );
  OAI221_X1 U23227 ( .B1(n21488), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n21488), 
        .C2(n21487), .A(n21486), .ZN(P3_U3282) );
  AOI22_X1 U23228 ( .A1(n21491), .A2(n21490), .B1(n21876), .B2(n21489), .ZN(
        n21492) );
  INV_X1 U23229 ( .A(n21492), .ZN(n21496) );
  NOR2_X1 U23230 ( .A1(n21494), .A2(n21493), .ZN(n21495) );
  MUX2_X1 U23231 ( .A(n21496), .B(n21495), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n21498) );
  OAI211_X1 U23232 ( .C1(n21499), .C2(n21500), .A(n21498), .B(n21497), .ZN(
        P3_U2996) );
  NOR2_X1 U23233 ( .A1(n21501), .A2(n21500), .ZN(n21507) );
  INV_X1 U23234 ( .A(n21507), .ZN(n21504) );
  NAND2_X1 U23235 ( .A1(n21504), .A2(P3_MORE_REG_SCAN_IN), .ZN(n21502) );
  OAI21_X1 U23236 ( .B1(n21504), .B2(n21503), .A(n21502), .ZN(P3_U3295) );
  OAI21_X1 U23237 ( .B1(n21507), .B2(n21506), .A(n21505), .ZN(P3_U2637) );
  INV_X1 U23238 ( .A(n21508), .ZN(n21509) );
  AOI211_X1 U23239 ( .C1(n21510), .C2(n15084), .A(n22106), .B(n21509), .ZN(
        n21512) );
  OAI21_X1 U23240 ( .B1(n21512), .B2(n21804), .A(n21511), .ZN(n21517) );
  AOI211_X1 U23241 ( .C1(n21515), .C2(n21834), .A(n21514), .B(n21513), .ZN(
        n21516) );
  MUX2_X1 U23242 ( .A(n21517), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n21516), 
        .Z(P1_U3485) );
  AOI22_X1 U23243 ( .A1(n21519), .A2(n21596), .B1(n21595), .B2(n21518), .ZN(
        n21528) );
  NAND2_X1 U23244 ( .A1(n21585), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n21527) );
  OR3_X1 U23245 ( .A1(n21521), .A2(n21520), .A3(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21526) );
  NOR2_X1 U23246 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n21522), .ZN(
        n21524) );
  OAI21_X1 U23247 ( .B1(n21524), .B2(n21523), .A(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21525) );
  NAND4_X1 U23248 ( .A1(n21528), .A2(n21527), .A3(n21526), .A4(n21525), .ZN(
        P1_U3017) );
  INV_X1 U23249 ( .A(n21529), .ZN(n21534) );
  OAI21_X1 U23250 ( .B1(n21531), .B2(n21534), .A(n21530), .ZN(n21532) );
  AOI21_X1 U23251 ( .B1(n21544), .B2(n21542), .A(n21532), .ZN(n21553) );
  NAND3_X1 U23252 ( .A1(n21534), .A2(n21533), .A3(n21552), .ZN(n21550) );
  NAND2_X1 U23253 ( .A1(n21595), .A2(n21637), .ZN(n21536) );
  OAI211_X1 U23254 ( .C1(n21537), .C2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n21536), .B(n21535), .ZN(n21538) );
  AOI21_X1 U23255 ( .B1(n21539), .B2(n21596), .A(n21538), .ZN(n21540) );
  OAI221_X1 U23256 ( .B1(n21541), .B2(n21553), .C1(n21541), .C2(n21550), .A(
        n21540), .ZN(P1_U3025) );
  INV_X1 U23257 ( .A(n21625), .ZN(n21547) );
  NAND3_X1 U23258 ( .A1(n21544), .A2(n21543), .A3(n21542), .ZN(n21546) );
  OAI211_X1 U23259 ( .C1(n21560), .C2(n21547), .A(n21546), .B(n21545), .ZN(
        n21548) );
  AOI21_X1 U23260 ( .B1(n21549), .B2(n21596), .A(n21548), .ZN(n21551) );
  OAI211_X1 U23261 ( .C1(n21553), .C2(n21552), .A(n21551), .B(n21550), .ZN(
        P1_U3026) );
  INV_X1 U23262 ( .A(n21554), .ZN(n21562) );
  INV_X1 U23263 ( .A(n21555), .ZN(n21557) );
  NAND3_X1 U23264 ( .A1(n21558), .A2(n21557), .A3(n21556), .ZN(n21559) );
  OAI21_X1 U23265 ( .B1(n21560), .B2(n21742), .A(n21559), .ZN(n21561) );
  AOI21_X1 U23266 ( .B1(n21562), .B2(n21596), .A(n21561), .ZN(n21564) );
  NAND2_X1 U23267 ( .A1(n21585), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n21563) );
  OAI211_X1 U23268 ( .C1(n21566), .C2(n21565), .A(n21564), .B(n21563), .ZN(
        P1_U3015) );
  AOI22_X1 U23269 ( .A1(n21568), .A2(n21596), .B1(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n21567), .ZN(n21573) );
  NAND2_X1 U23270 ( .A1(n21585), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n21572) );
  NAND2_X1 U23271 ( .A1(n21569), .A2(n21595), .ZN(n21571) );
  NAND4_X1 U23272 ( .A1(n21573), .A2(n21572), .A3(n21571), .A4(n21570), .ZN(
        P1_U3010) );
  INV_X1 U23273 ( .A(n21574), .ZN(n21577) );
  INV_X1 U23274 ( .A(n21575), .ZN(n21576) );
  NOR2_X1 U23275 ( .A1(n21600), .A2(n21578), .ZN(n21579) );
  AOI221_X1 U23276 ( .B1(n21582), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), 
        .C1(n21581), .C2(n21580), .A(n21579), .ZN(n21583) );
  NAND2_X1 U23277 ( .A1(n21584), .A2(n21583), .ZN(P1_U3004) );
  AOI22_X1 U23278 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n21586), .B1(
        n21585), .B2(P1_REIP_REG_25__SCAN_IN), .ZN(n21591) );
  INV_X1 U23279 ( .A(n21587), .ZN(n21589) );
  AOI22_X1 U23280 ( .A1(n21589), .A2(n21596), .B1(n21595), .B2(n21588), .ZN(
        n21590) );
  OAI211_X1 U23281 ( .C1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n21592), .A(
        n21591), .B(n21590), .ZN(P1_U3006) );
  INV_X1 U23282 ( .A(n21593), .ZN(n21597) );
  AOI22_X1 U23283 ( .A1(n21597), .A2(n21596), .B1(n21595), .B2(n21594), .ZN(
        n21606) );
  INV_X1 U23284 ( .A(n21598), .ZN(n21604) );
  NOR2_X1 U23285 ( .A1(n21600), .A2(n21599), .ZN(n21601) );
  AOI221_X1 U23286 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n21604), 
        .C1(n21603), .C2(n21602), .A(n21601), .ZN(n21605) );
  NAND2_X1 U23287 ( .A1(n21606), .A2(n21605), .ZN(P1_U3008) );
  OAI21_X1 U23288 ( .B1(n21622), .B2(n21623), .A(n21738), .ZN(n21628) );
  INV_X1 U23289 ( .A(n21607), .ZN(n21618) );
  NAND2_X1 U23290 ( .A1(n21782), .A2(n21608), .ZN(n21615) );
  AOI22_X1 U23291 ( .A1(n21724), .A2(n21611), .B1(n21610), .B2(n21609), .ZN(
        n21612) );
  NAND2_X1 U23292 ( .A1(n21729), .A2(n21612), .ZN(n21613) );
  AOI21_X1 U23293 ( .B1(n21773), .B2(P1_EBX_REG_4__SCAN_IN), .A(n21613), .ZN(
        n21614) );
  OAI211_X1 U23294 ( .C1(n21776), .C2(n21616), .A(n21615), .B(n21614), .ZN(
        n21617) );
  AOI21_X1 U23295 ( .B1(n21618), .B2(n21631), .A(n21617), .ZN(n21619) );
  OAI221_X1 U23296 ( .B1(n21628), .B2(n21621), .C1(n21628), .C2(n21620), .A(
        n21619), .ZN(P1_U2836) );
  NOR2_X1 U23297 ( .A1(n21623), .A2(n21622), .ZN(n21624) );
  AOI22_X1 U23298 ( .A1(n21724), .A2(n21625), .B1(n21624), .B2(n21627), .ZN(
        n21634) );
  AOI21_X1 U23299 ( .B1(n21773), .B2(P1_EBX_REG_5__SCAN_IN), .A(n21745), .ZN(
        n21626) );
  OAI21_X1 U23300 ( .B1(n21776), .B2(n20149), .A(n21626), .ZN(n21630) );
  NOR2_X1 U23301 ( .A1(n21628), .A2(n21627), .ZN(n21629) );
  AOI211_X1 U23302 ( .C1(n21632), .C2(n21631), .A(n21630), .B(n21629), .ZN(
        n21633) );
  OAI211_X1 U23303 ( .C1(n21635), .C2(n21702), .A(n21634), .B(n21633), .ZN(
        P1_U2835) );
  AND2_X1 U23304 ( .A1(n21738), .A2(n21636), .ZN(n21654) );
  AOI22_X1 U23305 ( .A1(n21724), .A2(n21637), .B1(P1_REIP_REG_6__SCAN_IN), 
        .B2(n21654), .ZN(n21648) );
  NOR2_X1 U23306 ( .A1(n21638), .A2(P1_REIP_REG_6__SCAN_IN), .ZN(n21641) );
  INV_X1 U23307 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n21639) );
  OAI21_X1 U23308 ( .B1(n21761), .B2(n21639), .A(n21729), .ZN(n21640) );
  NOR2_X1 U23309 ( .A1(n21641), .A2(n21640), .ZN(n21642) );
  OAI21_X1 U23310 ( .B1(n21776), .B2(n21643), .A(n21642), .ZN(n21644) );
  INV_X1 U23311 ( .A(n21644), .ZN(n21647) );
  OR2_X1 U23312 ( .A1(n21645), .A2(n21777), .ZN(n21646) );
  AND3_X1 U23313 ( .A1(n21648), .A2(n21647), .A3(n21646), .ZN(n21649) );
  OAI21_X1 U23314 ( .B1(n21650), .B2(n21702), .A(n21649), .ZN(P1_U2834) );
  AOI22_X1 U23315 ( .A1(n21748), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n21773), .B2(P1_EBX_REG_7__SCAN_IN), .ZN(n21651) );
  OAI211_X1 U23316 ( .C1(n21788), .C2(n21652), .A(n21651), .B(n21729), .ZN(
        n21653) );
  AOI221_X1 U23317 ( .B1(n21656), .B2(n21655), .C1(n21654), .C2(
        P1_REIP_REG_7__SCAN_IN), .A(n21653), .ZN(n21660) );
  INV_X1 U23318 ( .A(n21657), .ZN(n21658) );
  NAND2_X1 U23319 ( .A1(n21658), .A2(n21754), .ZN(n21659) );
  OAI211_X1 U23320 ( .C1(n21702), .C2(n21661), .A(n21660), .B(n21659), .ZN(
        P1_U2833) );
  AOI22_X1 U23321 ( .A1(n21662), .A2(n21724), .B1(n21773), .B2(
        P1_EBX_REG_8__SCAN_IN), .ZN(n21672) );
  AOI21_X1 U23322 ( .B1(n21748), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n21745), .ZN(n21671) );
  INV_X1 U23323 ( .A(n21663), .ZN(n21664) );
  AOI22_X1 U23324 ( .A1(n21665), .A2(n21754), .B1(n21664), .B2(n21782), .ZN(
        n21670) );
  INV_X1 U23325 ( .A(n21666), .ZN(n21668) );
  NOR2_X1 U23326 ( .A1(n21667), .A2(n21666), .ZN(n21683) );
  NOR2_X1 U23327 ( .A1(n21683), .A2(n21710), .ZN(n21678) );
  OAI21_X1 U23328 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(n21668), .A(n21678), .ZN(
        n21669) );
  NAND4_X1 U23329 ( .A1(n21672), .A2(n21671), .A3(n21670), .A4(n21669), .ZN(
        P1_U2832) );
  INV_X1 U23330 ( .A(n21683), .ZN(n21682) );
  INV_X1 U23331 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n21676) );
  AOI22_X1 U23332 ( .A1(n21674), .A2(n21782), .B1(n21724), .B2(n21673), .ZN(
        n21675) );
  OAI211_X1 U23333 ( .C1(n21761), .C2(n21676), .A(n21729), .B(n21675), .ZN(
        n21677) );
  AOI21_X1 U23334 ( .B1(n21748), .B2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n21677), .ZN(n21681) );
  AOI22_X1 U23335 ( .A1(n21679), .A2(n21754), .B1(P1_REIP_REG_9__SCAN_IN), 
        .B2(n21678), .ZN(n21680) );
  OAI211_X1 U23336 ( .C1(P1_REIP_REG_9__SCAN_IN), .C2(n21682), .A(n21681), .B(
        n21680), .ZN(P1_U2831) );
  NAND2_X1 U23337 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n21683), .ZN(n21692) );
  NOR2_X1 U23338 ( .A1(n21710), .A2(n21684), .ZN(n21697) );
  AOI22_X1 U23339 ( .A1(n21685), .A2(n21724), .B1(n21773), .B2(
        P1_EBX_REG_10__SCAN_IN), .ZN(n21686) );
  OAI211_X1 U23340 ( .C1(n21776), .C2(n13219), .A(n21686), .B(n21729), .ZN(
        n21687) );
  AOI21_X1 U23341 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(n21697), .A(n21687), 
        .ZN(n21691) );
  AOI22_X1 U23342 ( .A1(n21689), .A2(n21754), .B1(n21782), .B2(n21688), .ZN(
        n21690) );
  OAI211_X1 U23343 ( .C1(P1_REIP_REG_10__SCAN_IN), .C2(n21692), .A(n21691), 
        .B(n21690), .ZN(P1_U2830) );
  AOI22_X1 U23344 ( .A1(n21693), .A2(n21724), .B1(n21773), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n21694) );
  OAI211_X1 U23345 ( .C1(n21776), .C2(n13283), .A(n21694), .B(n21729), .ZN(
        n21695) );
  AOI221_X1 U23346 ( .B1(n21697), .B2(P1_REIP_REG_11__SCAN_IN), .C1(n21707), 
        .C2(n21696), .A(n21695), .ZN(n21700) );
  OR2_X1 U23347 ( .A1(n21777), .A2(n21698), .ZN(n21699) );
  OAI211_X1 U23348 ( .C1(n21702), .C2(n21701), .A(n21700), .B(n21699), .ZN(
        P1_U2829) );
  INV_X1 U23349 ( .A(n21703), .ZN(n21705) );
  AOI21_X1 U23350 ( .B1(n21773), .B2(P1_EBX_REG_12__SCAN_IN), .A(n21745), .ZN(
        n21704) );
  OAI21_X1 U23351 ( .B1(n21705), .B2(n21788), .A(n21704), .ZN(n21706) );
  AOI21_X1 U23352 ( .B1(n21748), .B2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n21706), .ZN(n21715) );
  NAND2_X1 U23353 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n21707), .ZN(n21708) );
  OAI21_X1 U23354 ( .B1(n21710), .B2(n21709), .A(n21708), .ZN(n21711) );
  AOI22_X1 U23355 ( .A1(n21713), .A2(n21782), .B1(n21712), .B2(n21711), .ZN(
        n21714) );
  OAI211_X1 U23356 ( .C1(n21777), .C2(n21716), .A(n21715), .B(n21714), .ZN(
        P1_U2828) );
  INV_X1 U23357 ( .A(n21717), .ZN(n21718) );
  AOI21_X1 U23358 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n21738), .A(n21718), 
        .ZN(n21728) );
  OAI22_X1 U23359 ( .A1(n21776), .A2(n21720), .B1(n21719), .B2(n21761), .ZN(
        n21721) );
  AOI211_X1 U23360 ( .C1(n21782), .C2(n21722), .A(n21745), .B(n21721), .ZN(
        n21727) );
  AOI22_X1 U23361 ( .A1(n21725), .A2(n21754), .B1(n21724), .B2(n21723), .ZN(
        n21726) );
  OAI211_X1 U23362 ( .C1(n21739), .C2(n21728), .A(n21727), .B(n21726), .ZN(
        P1_U2825) );
  OAI21_X1 U23363 ( .B1(n21761), .B2(n21730), .A(n21729), .ZN(n21731) );
  AOI21_X1 U23364 ( .B1(n21748), .B2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n21731), .ZN(n21734) );
  NAND2_X1 U23365 ( .A1(n21782), .A2(n21732), .ZN(n21733) );
  OAI211_X1 U23366 ( .C1(n21735), .C2(n21777), .A(n21734), .B(n21733), .ZN(
        n21736) );
  INV_X1 U23367 ( .A(n21736), .ZN(n21741) );
  OAI211_X1 U23368 ( .C1(n21739), .C2(P1_REIP_REG_16__SCAN_IN), .A(n21738), 
        .B(n21737), .ZN(n21740) );
  OAI211_X1 U23369 ( .C1(n21742), .C2(n21788), .A(n21741), .B(n21740), .ZN(
        P1_U2824) );
  NOR2_X1 U23370 ( .A1(n21744), .A2(n21743), .ZN(n21760) );
  OAI21_X1 U23371 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(P1_REIP_REG_18__SCAN_IN), 
        .A(n21759), .ZN(n21758) );
  AOI21_X1 U23372 ( .B1(n21773), .B2(P1_EBX_REG_19__SCAN_IN), .A(n21745), .ZN(
        n21750) );
  INV_X1 U23373 ( .A(n21746), .ZN(n21747) );
  AOI22_X1 U23374 ( .A1(n21748), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n21782), .B2(n21747), .ZN(n21749) );
  OAI211_X1 U23375 ( .C1(n21751), .C2(n21788), .A(n21750), .B(n21749), .ZN(
        n21752) );
  INV_X1 U23376 ( .A(n21752), .ZN(n21757) );
  AOI22_X1 U23377 ( .A1(n21755), .A2(n21754), .B1(P1_REIP_REG_19__SCAN_IN), 
        .B2(n21753), .ZN(n21756) );
  OAI211_X1 U23378 ( .C1(n21760), .C2(n21758), .A(n21757), .B(n21756), .ZN(
        P1_U2821) );
  AOI21_X1 U23379 ( .B1(n21760), .B2(n21759), .A(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n21771) );
  OAI22_X1 U23380 ( .A1(n21776), .A2(n21763), .B1(n21762), .B2(n21761), .ZN(
        n21767) );
  OAI22_X1 U23381 ( .A1(n21765), .A2(n21777), .B1(n21764), .B2(n21788), .ZN(
        n21766) );
  AOI211_X1 U23382 ( .C1(n21768), .C2(n21782), .A(n21767), .B(n21766), .ZN(
        n21769) );
  OAI21_X1 U23383 ( .B1(n21771), .B2(n21770), .A(n21769), .ZN(P1_U2820) );
  AOI22_X1 U23384 ( .A1(n21773), .A2(P1_EBX_REG_24__SCAN_IN), .B1(
        P1_REIP_REG_24__SCAN_IN), .B2(n21772), .ZN(n21774) );
  OAI21_X1 U23385 ( .B1(n21776), .B2(n21775), .A(n21774), .ZN(n21780) );
  NOR2_X1 U23386 ( .A1(n21778), .A2(n21777), .ZN(n21779) );
  AOI211_X1 U23387 ( .C1(n21782), .C2(n21781), .A(n21780), .B(n21779), .ZN(
        n21783) );
  INV_X1 U23388 ( .A(n21783), .ZN(n21784) );
  AOI21_X1 U23389 ( .B1(n21785), .B2(n16118), .A(n21784), .ZN(n21786) );
  OAI21_X1 U23390 ( .B1(n21788), .B2(n21787), .A(n21786), .ZN(P1_U2816) );
  OAI21_X1 U23391 ( .B1(n21791), .B2(n21790), .A(n21789), .ZN(P1_U2806) );
  OAI22_X1 U23392 ( .A1(n21795), .A2(n21794), .B1(n21793), .B2(n21792), .ZN(
        n21797) );
  MUX2_X1 U23393 ( .A(n21797), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n21796), .Z(P1_U3469) );
  NOR4_X1 U23394 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21841), .A3(n21798), 
        .A4(n21804), .ZN(n21799) );
  NOR2_X1 U23395 ( .A1(n21800), .A2(n21799), .ZN(n21802) );
  OAI211_X1 U23396 ( .C1(n21805), .C2(n22106), .A(n21802), .B(n21801), .ZN(
        P1_U3163) );
  OAI22_X1 U23397 ( .A1(n21805), .A2(n22072), .B1(n21804), .B2(n21803), .ZN(
        P1_U3466) );
  AOI21_X1 U23398 ( .B1(n21808), .B2(n21807), .A(n21806), .ZN(n21809) );
  OAI22_X1 U23399 ( .A1(n21811), .A2(n21810), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n21809), .ZN(n21812) );
  OAI21_X1 U23400 ( .B1(n21814), .B2(n21813), .A(n21812), .ZN(P1_U3161) );
  AOI21_X1 U23401 ( .B1(n17343), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21816), 
        .ZN(n21815) );
  INV_X1 U23402 ( .A(n21815), .ZN(P1_U2805) );
  AOI21_X1 U23403 ( .B1(n17343), .B2(P1_DATAWIDTH_REG_1__SCAN_IN), .A(n21816), 
        .ZN(n21817) );
  INV_X1 U23404 ( .A(n21817), .ZN(P1_U3465) );
  INV_X1 U23405 ( .A(n21818), .ZN(n21820) );
  OAI21_X1 U23406 ( .B1(n21822), .B2(n21819), .A(n21820), .ZN(P2_U2818) );
  OAI21_X1 U23407 ( .B1(n21822), .B2(n21821), .A(n21820), .ZN(P2_U3592) );
  OAI21_X1 U23408 ( .B1(n21826), .B2(n21823), .A(n21824), .ZN(P3_U2636) );
  OAI21_X1 U23409 ( .B1(n21826), .B2(n21825), .A(n21824), .ZN(P3_U3281) );
  INV_X1 U23410 ( .A(HOLD), .ZN(n21869) );
  OAI21_X1 U23411 ( .B1(n21869), .B2(n21827), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21828) );
  INV_X1 U23412 ( .A(n21828), .ZN(n21830) );
  AOI21_X1 U23413 ( .B1(n21876), .B2(P3_STATE_REG_1__SCAN_IN), .A(n21881), 
        .ZN(n21883) );
  OAI21_X1 U23414 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n21833), .A(
        P3_STATE_REG_2__SCAN_IN), .ZN(n21882) );
  INV_X1 U23415 ( .A(n21882), .ZN(n21829) );
  OAI22_X1 U23416 ( .A1(n21831), .A2(n21830), .B1(n21883), .B2(n21829), .ZN(
        P3_U3029) );
  AOI21_X1 U23417 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21841), .A(n21847), 
        .ZN(n21849) );
  INV_X1 U23418 ( .A(n21849), .ZN(n21832) );
  OAI211_X1 U23419 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n21833), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n21832), .ZN(n21839) );
  NOR3_X1 U23420 ( .A1(NA), .A2(n21847), .A3(n21834), .ZN(n21836) );
  OAI21_X1 U23421 ( .B1(n21840), .B2(n21869), .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21845) );
  OAI211_X1 U23422 ( .C1(n21836), .C2(n21835), .A(HOLD), .B(n21845), .ZN(
        n21838) );
  NAND3_X1 U23423 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(
        P1_REQUESTPENDING_REG_SCAN_IN), .A3(n21836), .ZN(n21837) );
  NAND3_X1 U23424 ( .A1(n21839), .A2(n21838), .A3(n21837), .ZN(P1_U3196) );
  OAI221_X1 U23425 ( .B1(n21841), .B2(HOLD), .C1(n21841), .C2(n21840), .A(
        P1_STATE_REG_1__SCAN_IN), .ZN(n21843) );
  OAI211_X1 U23426 ( .C1(n21847), .C2(n21845), .A(n21843), .B(n21842), .ZN(
        P1_U3195) );
  INV_X1 U23427 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n21844) );
  NOR2_X1 U23428 ( .A1(n21844), .A2(n21869), .ZN(n21846) );
  AOI211_X1 U23429 ( .C1(NA), .C2(n21847), .A(n21846), .B(n21845), .ZN(n21848)
         );
  OAI22_X1 U23430 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21849), .B1(n22401), 
        .B2(n21848), .ZN(P1_U3194) );
  OAI21_X1 U23431 ( .B1(P2_STATE_REG_2__SCAN_IN), .B2(P2_STATE_REG_1__SCAN_IN), 
        .A(HOLD), .ZN(n21854) );
  NAND2_X1 U23432 ( .A1(n21850), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n21861) );
  NAND2_X1 U23433 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n21861), .ZN(n21865) );
  INV_X1 U23434 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n21856) );
  AOI22_X1 U23435 ( .A1(n21851), .A2(n21865), .B1(n21856), .B2(n17762), .ZN(
        n21853) );
  NAND2_X1 U23436 ( .A1(n21852), .A2(NA), .ZN(n21864) );
  OAI211_X1 U23437 ( .C1(n21855), .C2(n21854), .A(n21853), .B(n21864), .ZN(
        P2_U3209) );
  NAND2_X1 U23438 ( .A1(n21869), .A2(n21856), .ZN(n21863) );
  AOI211_X1 U23439 ( .C1(P2_STATE_REG_2__SCAN_IN), .C2(HOLD), .A(n21867), .B(
        n21856), .ZN(n21858) );
  AOI211_X1 U23440 ( .C1(n21859), .C2(n21863), .A(n21858), .B(n21857), .ZN(
        n21860) );
  NAND2_X1 U23441 ( .A1(n21860), .A2(n21861), .ZN(P2_U3210) );
  OAI22_X1 U23442 ( .A1(NA), .A2(n21861), .B1(P2_STATE_REG_1__SCAN_IN), .B2(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n21862) );
  AOI22_X1 U23443 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(HOLD), .B1(n21863), .B2(
        n21862), .ZN(n21868) );
  NAND3_X1 U23444 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n21865), .A3(n21864), 
        .ZN(n21866) );
  OAI21_X1 U23445 ( .B1(n21868), .B2(n21867), .A(n21866), .ZN(P2_U3211) );
  NOR2_X1 U23446 ( .A1(n21871), .A2(n21869), .ZN(n21879) );
  NOR2_X1 U23447 ( .A1(HOLD), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21875)
         );
  INV_X1 U23448 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21872) );
  OAI211_X1 U23449 ( .C1(n21881), .C2(n21872), .A(n21871), .B(n21870), .ZN(
        n21873) );
  OAI21_X1 U23450 ( .B1(n21876), .B2(n18553), .A(n21873), .ZN(n21874) );
  AOI221_X1 U23451 ( .B1(n21879), .B2(n21883), .C1(n21875), .C2(n21883), .A(
        n21874), .ZN(P3_U3030) );
  NAND2_X1 U23452 ( .A1(n21876), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n21877) );
  OAI22_X1 U23453 ( .A1(NA), .A2(n21877), .B1(P3_STATE_REG_1__SCAN_IN), .B2(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21878) );
  OAI22_X1 U23454 ( .A1(n21879), .A2(n21878), .B1(HOLD), .B2(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21880) );
  OAI22_X1 U23455 ( .A1(n21883), .A2(n21882), .B1(n21881), .B2(n21880), .ZN(
        P3_U3031) );
  INV_X1 U23456 ( .A(n21884), .ZN(n21885) );
  NOR2_X1 U23457 ( .A1(n21886), .A2(n21885), .ZN(n21889) );
  AOI21_X1 U23458 ( .B1(P1_UWORD_REG_8__SCAN_IN), .B2(n21945), .A(n21889), 
        .ZN(n21887) );
  OAI21_X1 U23459 ( .B1(n21888), .B2(n21951), .A(n21887), .ZN(P1_U2945) );
  AOI21_X1 U23460 ( .B1(P1_LWORD_REG_8__SCAN_IN), .B2(n21945), .A(n21889), 
        .ZN(n21890) );
  OAI21_X1 U23461 ( .B1(n21891), .B2(n21951), .A(n21890), .ZN(P1_U2960) );
  INV_X1 U23462 ( .A(n21892), .ZN(n21893) );
  NAND2_X1 U23463 ( .A1(n21943), .A2(n21893), .ZN(n21901) );
  INV_X1 U23464 ( .A(n21901), .ZN(n21894) );
  AOI21_X1 U23465 ( .B1(P1_UWORD_REG_9__SCAN_IN), .B2(n21945), .A(n21894), 
        .ZN(n21895) );
  OAI21_X1 U23466 ( .B1(n21896), .B2(n21951), .A(n21895), .ZN(P1_U2946) );
  INV_X1 U23467 ( .A(P1_LWORD_REG_9__SCAN_IN), .ZN(n21897) );
  OR2_X1 U23468 ( .A1(n21949), .A2(n21897), .ZN(n21898) );
  OAI21_X1 U23469 ( .B1(n21951), .B2(n21899), .A(n21898), .ZN(n21900) );
  INV_X1 U23470 ( .A(n21900), .ZN(n21902) );
  NAND2_X1 U23471 ( .A1(n21902), .A2(n21901), .ZN(P1_U2961) );
  NAND2_X1 U23472 ( .A1(n21943), .A2(n21903), .ZN(n21910) );
  INV_X1 U23473 ( .A(n21910), .ZN(n21904) );
  AOI21_X1 U23474 ( .B1(P1_UWORD_REG_10__SCAN_IN), .B2(n21945), .A(n21904), 
        .ZN(n21905) );
  OAI21_X1 U23475 ( .B1(n21906), .B2(n21951), .A(n21905), .ZN(P1_U2947) );
  INV_X1 U23476 ( .A(P1_LWORD_REG_10__SCAN_IN), .ZN(n21907) );
  OR2_X1 U23477 ( .A1(n21949), .A2(n21907), .ZN(n21908) );
  OAI21_X1 U23478 ( .B1(n21951), .B2(n20036), .A(n21908), .ZN(n21909) );
  INV_X1 U23479 ( .A(n21909), .ZN(n21911) );
  NAND2_X1 U23480 ( .A1(n21911), .A2(n21910), .ZN(P1_U2962) );
  INV_X1 U23481 ( .A(n21912), .ZN(n21913) );
  NAND2_X1 U23482 ( .A1(n21943), .A2(n21913), .ZN(n21921) );
  INV_X1 U23483 ( .A(n21921), .ZN(n21914) );
  AOI21_X1 U23484 ( .B1(P1_UWORD_REG_11__SCAN_IN), .B2(n21945), .A(n21914), 
        .ZN(n21915) );
  OAI21_X1 U23485 ( .B1(n21916), .B2(n21951), .A(n21915), .ZN(P1_U2948) );
  INV_X1 U23486 ( .A(P1_LWORD_REG_11__SCAN_IN), .ZN(n21917) );
  OR2_X1 U23487 ( .A1(n21949), .A2(n21917), .ZN(n21918) );
  OAI21_X1 U23488 ( .B1(n21951), .B2(n21919), .A(n21918), .ZN(n21920) );
  INV_X1 U23489 ( .A(n21920), .ZN(n21922) );
  NAND2_X1 U23490 ( .A1(n21922), .A2(n21921), .ZN(P1_U2963) );
  NAND2_X1 U23491 ( .A1(n21943), .A2(n21923), .ZN(n21931) );
  INV_X1 U23492 ( .A(n21931), .ZN(n21924) );
  AOI21_X1 U23493 ( .B1(P1_UWORD_REG_12__SCAN_IN), .B2(n21945), .A(n21924), 
        .ZN(n21925) );
  OAI21_X1 U23494 ( .B1(n21926), .B2(n21951), .A(n21925), .ZN(P1_U2949) );
  INV_X1 U23495 ( .A(P1_LWORD_REG_12__SCAN_IN), .ZN(n21927) );
  OR2_X1 U23496 ( .A1(n21949), .A2(n21927), .ZN(n21928) );
  OAI21_X1 U23497 ( .B1(n21951), .B2(n21929), .A(n21928), .ZN(n21930) );
  INV_X1 U23498 ( .A(n21930), .ZN(n21932) );
  NAND2_X1 U23499 ( .A1(n21932), .A2(n21931), .ZN(P1_U2964) );
  NAND2_X1 U23500 ( .A1(n21943), .A2(n21933), .ZN(n21940) );
  INV_X1 U23501 ( .A(n21940), .ZN(n21934) );
  AOI21_X1 U23502 ( .B1(P1_UWORD_REG_13__SCAN_IN), .B2(n21945), .A(n21934), 
        .ZN(n21935) );
  OAI21_X1 U23503 ( .B1(n21936), .B2(n21951), .A(n21935), .ZN(P1_U2950) );
  INV_X1 U23504 ( .A(P1_LWORD_REG_13__SCAN_IN), .ZN(n21937) );
  OR2_X1 U23505 ( .A1(n21949), .A2(n21937), .ZN(n21938) );
  OAI21_X1 U23506 ( .B1(n21951), .B2(n20040), .A(n21938), .ZN(n21939) );
  INV_X1 U23507 ( .A(n21939), .ZN(n21941) );
  NAND2_X1 U23508 ( .A1(n21941), .A2(n21940), .ZN(P1_U2965) );
  NAND2_X1 U23509 ( .A1(n21943), .A2(n21942), .ZN(n21953) );
  INV_X1 U23510 ( .A(n21953), .ZN(n21944) );
  AOI21_X1 U23511 ( .B1(P1_UWORD_REG_14__SCAN_IN), .B2(n21945), .A(n21944), 
        .ZN(n21946) );
  OAI21_X1 U23512 ( .B1(n21947), .B2(n21951), .A(n21946), .ZN(P1_U2951) );
  INV_X1 U23513 ( .A(P1_LWORD_REG_14__SCAN_IN), .ZN(n21948) );
  OR2_X1 U23514 ( .A1(n21949), .A2(n21948), .ZN(n21950) );
  OAI21_X1 U23515 ( .B1(n21951), .B2(n20042), .A(n21950), .ZN(n21952) );
  INV_X1 U23516 ( .A(n21952), .ZN(n21954) );
  NAND2_X1 U23517 ( .A1(n21954), .A2(n21953), .ZN(P1_U2966) );
  INV_X1 U23518 ( .A(n22393), .ZN(n21957) );
  NAND2_X1 U23519 ( .A1(n21957), .A2(n22117), .ZN(n21958) );
  NOR2_X1 U23520 ( .A1(n22115), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n22000) );
  INV_X1 U23521 ( .A(n22000), .ZN(n22060) );
  OAI21_X1 U23522 ( .B1(n21958), .B2(n22317), .A(n22060), .ZN(n21965) );
  INV_X1 U23523 ( .A(n22063), .ZN(n21959) );
  OR2_X1 U23524 ( .A1(n22015), .A2(n21959), .ZN(n21987) );
  INV_X1 U23525 ( .A(n11019), .ZN(n22086) );
  NOR2_X1 U23526 ( .A1(n21987), .A2(n22086), .ZN(n21962) );
  INV_X1 U23527 ( .A(n21960), .ZN(n21967) );
  NAND3_X1 U23528 ( .A1(n22105), .A2(n22039), .A3(n22066), .ZN(n21971) );
  NOR2_X1 U23529 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21971), .ZN(
        n22310) );
  AOI22_X1 U23530 ( .A1(n22109), .A2(n22310), .B1(n22393), .B2(n11070), .ZN(
        n21969) );
  INV_X1 U23531 ( .A(n21962), .ZN(n21964) );
  INV_X1 U23532 ( .A(n22310), .ZN(n21963) );
  AOI22_X1 U23533 ( .A1(n21965), .A2(n21964), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n21963), .ZN(n21966) );
  AOI22_X1 U23534 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n22311), .B1(
        n22317), .B2(n11072), .ZN(n21968) );
  OAI211_X1 U23535 ( .C1(n22314), .C2(n22075), .A(n21969), .B(n21968), .ZN(
        P1_U3033) );
  NOR2_X1 U23536 ( .A1(n22076), .A2(n21971), .ZN(n22316) );
  INV_X1 U23537 ( .A(n21987), .ZN(n21970) );
  AOI21_X1 U23538 ( .B1(n21970), .B2(n22077), .A(n22316), .ZN(n21972) );
  OAI22_X1 U23539 ( .A1(n21972), .A2(n22115), .B1(n21971), .B2(n22106), .ZN(
        n22315) );
  AOI22_X1 U23540 ( .A1(n22109), .A2(n22316), .B1(n22108), .B2(n22315), .ZN(
        n21976) );
  INV_X1 U23541 ( .A(n21971), .ZN(n21974) );
  OAI211_X1 U23542 ( .C1(n21988), .C2(n15084), .A(n22059), .B(n21972), .ZN(
        n21973) );
  OAI211_X1 U23543 ( .C1(n22059), .C2(n21974), .A(n22113), .B(n21973), .ZN(
        n22318) );
  AOI22_X1 U23544 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n22318), .B1(
        n22317), .B2(n11070), .ZN(n21975) );
  OAI211_X1 U23545 ( .C1(n11071), .C2(n22321), .A(n21976), .B(n21975), .ZN(
        P1_U3041) );
  NOR3_X1 U23546 ( .A1(n22330), .A2(n22323), .A3(n22115), .ZN(n21977) );
  NOR2_X1 U23547 ( .A1(n21977), .A2(n22000), .ZN(n21983) );
  INV_X1 U23548 ( .A(n21983), .ZN(n21979) );
  NOR2_X1 U23549 ( .A1(n21987), .A2(n11019), .ZN(n21982) );
  NOR2_X1 U23550 ( .A1(n21978), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n22003) );
  NAND3_X1 U23551 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n22105), .A3(
        n22039), .ZN(n21993) );
  NOR2_X1 U23552 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21993), .ZN(
        n22322) );
  AOI22_X1 U23553 ( .A1(n22323), .A2(n11070), .B1(n22109), .B2(n22322), .ZN(
        n21985) );
  INV_X1 U23554 ( .A(n22322), .ZN(n21980) );
  NOR2_X1 U23555 ( .A1(n22003), .A2(n22106), .ZN(n22005) );
  AOI21_X1 U23556 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21980), .A(n22005), 
        .ZN(n21981) );
  AOI22_X1 U23557 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n22324), .B1(
        n22330), .B2(n11072), .ZN(n21984) );
  OAI211_X1 U23558 ( .C1(n22327), .C2(n22075), .A(n21985), .B(n21984), .ZN(
        P1_U3049) );
  INV_X1 U23559 ( .A(n21993), .ZN(n21990) );
  NOR2_X1 U23560 ( .A1(n22076), .A2(n21993), .ZN(n22328) );
  INV_X1 U23561 ( .A(n22328), .ZN(n21986) );
  OAI21_X1 U23562 ( .B1(n21987), .B2(n22100), .A(n21986), .ZN(n21995) );
  OR2_X1 U23563 ( .A1(n21988), .A2(n22111), .ZN(n21989) );
  AND2_X1 U23564 ( .A1(n21989), .A2(n22059), .ZN(n21991) );
  AOI22_X1 U23565 ( .A1(n22329), .A2(n11072), .B1(n22109), .B2(n22328), .ZN(
        n21998) );
  INV_X1 U23566 ( .A(n21991), .ZN(n21996) );
  AOI21_X1 U23567 ( .B1(n22115), .B2(n21993), .A(n21992), .ZN(n21994) );
  OAI21_X1 U23568 ( .B1(n21996), .B2(n21995), .A(n21994), .ZN(n22331) );
  AOI22_X1 U23569 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n22331), .B1(
        n22330), .B2(n11070), .ZN(n21997) );
  OAI211_X1 U23570 ( .C1(n22334), .C2(n22075), .A(n21998), .B(n21997), .ZN(
        P1_U3057) );
  NOR2_X1 U23571 ( .A1(n22337), .A2(n22115), .ZN(n22001) );
  AOI21_X1 U23572 ( .B1(n22001), .B2(n22010), .A(n22000), .ZN(n22009) );
  INV_X1 U23573 ( .A(n22009), .ZN(n22004) );
  NOR2_X1 U23574 ( .A1(n22002), .A2(n11019), .ZN(n22008) );
  NOR3_X2 U23575 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n22104), .ZN(n22336) );
  AOI22_X1 U23576 ( .A1(n22109), .A2(n22336), .B1(n22337), .B2(n11072), .ZN(
        n22012) );
  INV_X1 U23577 ( .A(n22336), .ZN(n22006) );
  AOI21_X1 U23578 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22006), .A(n22005), 
        .ZN(n22007) );
  OAI211_X1 U23579 ( .C1(n22009), .C2(n22008), .A(n22094), .B(n22007), .ZN(
        n22338) );
  AOI22_X1 U23580 ( .A1(n22338), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11070), .B2(n22335), .ZN(n22011) );
  OAI211_X1 U23581 ( .C1(n22341), .C2(n22075), .A(n22012), .B(n22011), .ZN(
        P1_U3081) );
  INV_X1 U23582 ( .A(n22058), .ZN(n22014) );
  NAND3_X1 U23583 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n22039), .A3(
        n22066), .ZN(n22025) );
  NOR2_X1 U23584 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22025), .ZN(
        n22343) );
  AND2_X1 U23585 ( .A1(n22015), .A2(n22063), .ZN(n22049) );
  AOI21_X1 U23586 ( .B1(n22049), .B2(n11019), .A(n22343), .ZN(n22020) );
  INV_X1 U23587 ( .A(n22037), .ZN(n22018) );
  INV_X1 U23588 ( .A(n22016), .ZN(n22017) );
  NOR2_X1 U23589 ( .A1(n22017), .A2(n22036), .ZN(n22065) );
  INV_X1 U23590 ( .A(n22065), .ZN(n22068) );
  OAI22_X1 U23591 ( .A1(n22020), .A2(n22115), .B1(n22018), .B2(n22068), .ZN(
        n22342) );
  AOI22_X1 U23592 ( .A1(n22109), .A2(n22343), .B1(n22108), .B2(n22342), .ZN(
        n22024) );
  INV_X1 U23593 ( .A(n22353), .ZN(n22019) );
  OAI21_X1 U23594 ( .B1(n22019), .B2(n22344), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n22021) );
  NAND2_X1 U23595 ( .A1(n22021), .A2(n22020), .ZN(n22022) );
  AOI22_X1 U23596 ( .A1(n22345), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11070), .B2(n22344), .ZN(n22023) );
  OAI211_X1 U23597 ( .C1(n11071), .C2(n22353), .A(n22024), .B(n22023), .ZN(
        P1_U3097) );
  NOR2_X1 U23598 ( .A1(n22076), .A2(n22025), .ZN(n22349) );
  AOI21_X1 U23599 ( .B1(n22049), .B2(n22077), .A(n22349), .ZN(n22026) );
  OAI22_X1 U23600 ( .A1(n22026), .A2(n22115), .B1(n22025), .B2(n22106), .ZN(
        n22348) );
  AOI22_X1 U23601 ( .A1(n22109), .A2(n22349), .B1(n22108), .B2(n22348), .ZN(
        n22031) );
  INV_X1 U23602 ( .A(n22025), .ZN(n22028) );
  OAI211_X1 U23603 ( .C1(n22055), .C2(n15084), .A(n22117), .B(n22026), .ZN(
        n22027) );
  OAI211_X1 U23604 ( .C1(n22059), .C2(n22028), .A(n22113), .B(n22027), .ZN(
        n22350) );
  INV_X1 U23605 ( .A(n22082), .ZN(n22029) );
  AOI22_X1 U23606 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n22350), .B1(
        n22354), .B2(n11072), .ZN(n22030) );
  OAI211_X1 U23607 ( .C1(n11069), .C2(n22353), .A(n22031), .B(n22030), .ZN(
        P1_U3105) );
  INV_X1 U23608 ( .A(n22354), .ZN(n22034) );
  INV_X1 U23609 ( .A(n22085), .ZN(n22032) );
  NAND3_X1 U23610 ( .A1(n22034), .A2(n22117), .A3(n22366), .ZN(n22035) );
  NAND2_X1 U23611 ( .A1(n22035), .A2(n22060), .ZN(n22043) );
  AND2_X1 U23612 ( .A1(n22049), .A2(n22086), .ZN(n22040) );
  NAND2_X1 U23613 ( .A1(n22036), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n22089) );
  INV_X1 U23614 ( .A(n22089), .ZN(n22038) );
  NAND3_X1 U23615 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n22039), .ZN(n22050) );
  NOR2_X1 U23616 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22050), .ZN(
        n22355) );
  AOI22_X1 U23617 ( .A1(n22109), .A2(n22355), .B1(n22354), .B2(n11070), .ZN(
        n22047) );
  INV_X1 U23618 ( .A(n22040), .ZN(n22042) );
  INV_X1 U23619 ( .A(n22355), .ZN(n22041) );
  AOI22_X1 U23620 ( .A1(n22043), .A2(n22042), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n22041), .ZN(n22044) );
  NAND2_X1 U23621 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n22089), .ZN(n22093) );
  NAND3_X1 U23622 ( .A1(n22045), .A2(n22044), .A3(n22093), .ZN(n22357) );
  AOI22_X1 U23623 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n22357), .B1(
        n22356), .B2(n11072), .ZN(n22046) );
  OAI211_X1 U23624 ( .C1(n22360), .C2(n22075), .A(n22047), .B(n22046), .ZN(
        P1_U3113) );
  NOR2_X1 U23625 ( .A1(n22076), .A2(n22050), .ZN(n22362) );
  INV_X1 U23626 ( .A(n22100), .ZN(n22048) );
  AOI21_X1 U23627 ( .B1(n22049), .B2(n22048), .A(n22362), .ZN(n22051) );
  OAI22_X1 U23628 ( .A1(n22051), .A2(n22115), .B1(n22050), .B2(n22106), .ZN(
        n22361) );
  AOI22_X1 U23629 ( .A1(n22109), .A2(n22362), .B1(n22108), .B2(n22361), .ZN(
        n22057) );
  INV_X1 U23630 ( .A(n22050), .ZN(n22053) );
  OAI211_X1 U23631 ( .C1(n22055), .C2(n22111), .A(n22059), .B(n22051), .ZN(
        n22052) );
  OAI211_X1 U23632 ( .C1(n22059), .C2(n22053), .A(n22113), .B(n22052), .ZN(
        n22363) );
  AOI22_X1 U23633 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n22363), .B1(
        n22369), .B2(n11072), .ZN(n22056) );
  OAI211_X1 U23634 ( .C1(n11069), .C2(n22366), .A(n22057), .B(n22056), .ZN(
        P1_U3121) );
  NAND2_X1 U23635 ( .A1(n22380), .A2(n22059), .ZN(n22061) );
  OAI21_X1 U23636 ( .B1(n22369), .B2(n22061), .A(n22060), .ZN(n22070) );
  OR2_X1 U23637 ( .A1(n22063), .A2(n22062), .ZN(n22101) );
  NOR2_X1 U23638 ( .A1(n22101), .A2(n22086), .ZN(n22067) );
  NAND3_X1 U23639 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n22066), .ZN(n22078) );
  NOR2_X1 U23640 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22078), .ZN(
        n22368) );
  AOI22_X1 U23641 ( .A1(n22109), .A2(n22368), .B1(n22367), .B2(n11072), .ZN(
        n22074) );
  INV_X1 U23642 ( .A(n22067), .ZN(n22069) );
  AOI22_X1 U23643 ( .A1(n22070), .A2(n22069), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n22068), .ZN(n22071) );
  AOI22_X1 U23644 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n22370), .B1(
        n22369), .B2(n11070), .ZN(n22073) );
  OAI211_X1 U23645 ( .C1(n22374), .C2(n22075), .A(n22074), .B(n22073), .ZN(
        P1_U3129) );
  NOR2_X1 U23646 ( .A1(n22076), .A2(n22078), .ZN(n22376) );
  INV_X1 U23647 ( .A(n22101), .ZN(n22087) );
  AOI21_X1 U23648 ( .B1(n22087), .B2(n22077), .A(n22376), .ZN(n22079) );
  OAI22_X1 U23649 ( .A1(n22079), .A2(n22115), .B1(n22078), .B2(n22106), .ZN(
        n22375) );
  AOI22_X1 U23650 ( .A1(n22109), .A2(n22376), .B1(n22108), .B2(n22375), .ZN(
        n22084) );
  INV_X1 U23651 ( .A(n22078), .ZN(n22081) );
  OAI21_X1 U23652 ( .B1(n22112), .B2(n15084), .A(n22079), .ZN(n22080) );
  OAI221_X1 U23653 ( .B1(n22117), .B2(n22081), .C1(n22115), .C2(n22080), .A(
        n22113), .ZN(n22377) );
  AOI22_X1 U23654 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n22377), .B1(
        n22384), .B2(n11072), .ZN(n22083) );
  OAI211_X1 U23655 ( .C1(n11069), .C2(n22380), .A(n22084), .B(n22083), .ZN(
        P1_U3137) );
  NOR3_X2 U23656 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22105), .A3(
        n22104), .ZN(n22382) );
  NAND2_X1 U23657 ( .A1(n22087), .A2(n22086), .ZN(n22091) );
  OAI22_X1 U23658 ( .A1(n22091), .A2(n22115), .B1(n22089), .B2(n22088), .ZN(
        n22381) );
  AOI22_X1 U23659 ( .A1(n22109), .A2(n22382), .B1(n22108), .B2(n22381), .ZN(
        n22098) );
  INV_X1 U23660 ( .A(n22397), .ZN(n22090) );
  OAI21_X1 U23661 ( .B1(n22384), .B2(n22090), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n22092) );
  AOI21_X1 U23662 ( .B1(n22092), .B2(n22091), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n22095) );
  AOI22_X1 U23663 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n22385), .B1(
        n22384), .B2(n11070), .ZN(n22097) );
  OAI211_X1 U23664 ( .C1(n11071), .C2(n22397), .A(n22098), .B(n22097), .ZN(
        P1_U3145) );
  NAND2_X1 U23665 ( .A1(n22099), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n22102) );
  INV_X1 U23666 ( .A(n22102), .ZN(n22390) );
  OR2_X1 U23667 ( .A1(n22101), .A2(n22100), .ZN(n22103) );
  AND2_X1 U23668 ( .A1(n22103), .A2(n22102), .ZN(n22110) );
  NOR2_X1 U23669 ( .A1(n22105), .A2(n22104), .ZN(n22116) );
  INV_X1 U23670 ( .A(n22116), .ZN(n22107) );
  OAI22_X1 U23671 ( .A1(n22110), .A2(n22115), .B1(n22107), .B2(n22106), .ZN(
        n22388) );
  AOI22_X1 U23672 ( .A1(n22109), .A2(n22390), .B1(n22108), .B2(n22388), .ZN(
        n22120) );
  OAI21_X1 U23673 ( .B1(n22112), .B2(n22111), .A(n22110), .ZN(n22114) );
  OAI221_X1 U23674 ( .B1(n22117), .B2(n22116), .C1(n22115), .C2(n22114), .A(
        n22113), .ZN(n22394) );
  AOI22_X1 U23675 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n22394), .B1(
        n22393), .B2(n11072), .ZN(n22119) );
  OAI211_X1 U23676 ( .C1(n11069), .C2(n22397), .A(n22120), .B(n22119), .ZN(
        P1_U3153) );
  AOI22_X1 U23677 ( .A1(n22148), .A2(n22310), .B1(n22393), .B2(n11062), .ZN(
        n22122) );
  AOI22_X1 U23678 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n22311), .B1(
        n22317), .B2(n11080), .ZN(n22121) );
  OAI211_X1 U23679 ( .C1(n22314), .C2(n22141), .A(n22122), .B(n22121), .ZN(
        P1_U3034) );
  AOI22_X1 U23680 ( .A1(n22148), .A2(n22316), .B1(n22147), .B2(n22315), .ZN(
        n22124) );
  AOI22_X1 U23681 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n22318), .B1(
        n22317), .B2(n11062), .ZN(n22123) );
  OAI211_X1 U23682 ( .C1(n11079), .C2(n22321), .A(n22124), .B(n22123), .ZN(
        P1_U3042) );
  AOI22_X1 U23683 ( .A1(n22323), .A2(n11062), .B1(n22148), .B2(n22322), .ZN(
        n22126) );
  AOI22_X1 U23684 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n22324), .B1(
        n22330), .B2(n11080), .ZN(n22125) );
  OAI211_X1 U23685 ( .C1(n22327), .C2(n22141), .A(n22126), .B(n22125), .ZN(
        P1_U3050) );
  AOI22_X1 U23686 ( .A1(n22329), .A2(n11080), .B1(n22148), .B2(n22328), .ZN(
        n22128) );
  AOI22_X1 U23687 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n22331), .B1(
        n22330), .B2(n11062), .ZN(n22127) );
  OAI211_X1 U23688 ( .C1(n22334), .C2(n22141), .A(n22128), .B(n22127), .ZN(
        P1_U3058) );
  AOI22_X1 U23689 ( .A1(n22148), .A2(n22336), .B1(n22337), .B2(n11080), .ZN(
        n22130) );
  AOI22_X1 U23690 ( .A1(n22338), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11062), .B2(n22335), .ZN(n22129) );
  OAI211_X1 U23691 ( .C1(n22341), .C2(n22141), .A(n22130), .B(n22129), .ZN(
        P1_U3082) );
  AOI22_X1 U23692 ( .A1(n22148), .A2(n22343), .B1(n22147), .B2(n22342), .ZN(
        n22132) );
  AOI22_X1 U23693 ( .A1(n22345), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n22344), .B2(n11062), .ZN(n22131) );
  OAI211_X1 U23694 ( .C1(n11079), .C2(n22353), .A(n22132), .B(n22131), .ZN(
        P1_U3098) );
  AOI22_X1 U23695 ( .A1(n22148), .A2(n22349), .B1(n22147), .B2(n22348), .ZN(
        n22134) );
  AOI22_X1 U23696 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n22350), .B1(
        n22354), .B2(n11080), .ZN(n22133) );
  OAI211_X1 U23697 ( .C1(n11061), .C2(n22353), .A(n22134), .B(n22133), .ZN(
        P1_U3106) );
  AOI22_X1 U23698 ( .A1(n22148), .A2(n22355), .B1(n22354), .B2(n11062), .ZN(
        n22136) );
  AOI22_X1 U23699 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n22357), .B1(
        n22356), .B2(n11080), .ZN(n22135) );
  OAI211_X1 U23700 ( .C1(n22360), .C2(n22141), .A(n22136), .B(n22135), .ZN(
        P1_U3114) );
  AOI22_X1 U23701 ( .A1(n22148), .A2(n22362), .B1(n22147), .B2(n22361), .ZN(
        n22138) );
  AOI22_X1 U23702 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n22363), .B1(
        n22369), .B2(n11080), .ZN(n22137) );
  OAI211_X1 U23703 ( .C1(n11061), .C2(n22366), .A(n22138), .B(n22137), .ZN(
        P1_U3122) );
  AOI22_X1 U23704 ( .A1(n22148), .A2(n22368), .B1(n22367), .B2(n11080), .ZN(
        n22140) );
  AOI22_X1 U23705 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n22370), .B1(
        n22369), .B2(n11062), .ZN(n22139) );
  OAI211_X1 U23706 ( .C1(n22374), .C2(n22141), .A(n22140), .B(n22139), .ZN(
        P1_U3130) );
  AOI22_X1 U23707 ( .A1(n22148), .A2(n22376), .B1(n22147), .B2(n22375), .ZN(
        n22143) );
  AOI22_X1 U23708 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n22377), .B1(
        n22384), .B2(n11080), .ZN(n22142) );
  OAI211_X1 U23709 ( .C1(n11061), .C2(n22380), .A(n22143), .B(n22142), .ZN(
        P1_U3138) );
  AOI22_X1 U23710 ( .A1(n22148), .A2(n22382), .B1(n22147), .B2(n22381), .ZN(
        n22146) );
  AOI22_X1 U23711 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n22385), .B1(
        n22384), .B2(n11062), .ZN(n22145) );
  OAI211_X1 U23712 ( .C1(n11079), .C2(n22397), .A(n22146), .B(n22145), .ZN(
        P1_U3146) );
  AOI22_X1 U23713 ( .A1(n22148), .A2(n22390), .B1(n22147), .B2(n22388), .ZN(
        n22151) );
  AOI22_X1 U23714 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n22394), .B1(
        n22393), .B2(n11080), .ZN(n22150) );
  OAI211_X1 U23715 ( .C1(n11061), .C2(n22397), .A(n22151), .B(n22150), .ZN(
        P1_U3154) );
  AOI22_X1 U23716 ( .A1(n22180), .A2(n22310), .B1(n22393), .B2(n22175), .ZN(
        n22153) );
  AOI22_X1 U23717 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n22311), .B1(
        n22317), .B2(n22181), .ZN(n22152) );
  OAI211_X1 U23718 ( .C1(n22314), .C2(n22172), .A(n22153), .B(n22152), .ZN(
        P1_U3035) );
  AOI22_X1 U23719 ( .A1(n22180), .A2(n22316), .B1(n22179), .B2(n22315), .ZN(
        n22155) );
  AOI22_X1 U23720 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n22318), .B1(
        n22317), .B2(n22175), .ZN(n22154) );
  OAI211_X1 U23721 ( .C1(n22178), .C2(n22321), .A(n22155), .B(n22154), .ZN(
        P1_U3043) );
  AOI22_X1 U23722 ( .A1(n22330), .A2(n22181), .B1(n22180), .B2(n22322), .ZN(
        n22157) );
  AOI22_X1 U23723 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n22324), .B1(
        n22323), .B2(n22175), .ZN(n22156) );
  OAI211_X1 U23724 ( .C1(n22327), .C2(n22172), .A(n22157), .B(n22156), .ZN(
        P1_U3051) );
  AOI22_X1 U23725 ( .A1(n22329), .A2(n22181), .B1(n22180), .B2(n22328), .ZN(
        n22159) );
  AOI22_X1 U23726 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n22331), .B1(
        n22330), .B2(n22175), .ZN(n22158) );
  OAI211_X1 U23727 ( .C1(n22334), .C2(n22172), .A(n22159), .B(n22158), .ZN(
        P1_U3059) );
  AOI22_X1 U23728 ( .A1(n22180), .A2(n22336), .B1(n22175), .B2(n22335), .ZN(
        n22161) );
  AOI22_X1 U23729 ( .A1(n22338), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n22337), .B2(n22181), .ZN(n22160) );
  OAI211_X1 U23730 ( .C1(n22341), .C2(n22172), .A(n22161), .B(n22160), .ZN(
        P1_U3083) );
  AOI22_X1 U23731 ( .A1(n22180), .A2(n22343), .B1(n22179), .B2(n22342), .ZN(
        n22163) );
  AOI22_X1 U23732 ( .A1(n22345), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n22344), .B2(n22175), .ZN(n22162) );
  OAI211_X1 U23733 ( .C1(n22178), .C2(n22353), .A(n22163), .B(n22162), .ZN(
        P1_U3099) );
  AOI22_X1 U23734 ( .A1(n22180), .A2(n22349), .B1(n22179), .B2(n22348), .ZN(
        n22165) );
  AOI22_X1 U23735 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n22350), .B1(
        n22354), .B2(n22181), .ZN(n22164) );
  OAI211_X1 U23736 ( .C1(n22184), .C2(n22353), .A(n22165), .B(n22164), .ZN(
        P1_U3107) );
  AOI22_X1 U23737 ( .A1(n22180), .A2(n22355), .B1(n22354), .B2(n22175), .ZN(
        n22167) );
  AOI22_X1 U23738 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n22357), .B1(
        n22356), .B2(n22181), .ZN(n22166) );
  OAI211_X1 U23739 ( .C1(n22360), .C2(n22172), .A(n22167), .B(n22166), .ZN(
        P1_U3115) );
  AOI22_X1 U23740 ( .A1(n22180), .A2(n22362), .B1(n22179), .B2(n22361), .ZN(
        n22169) );
  AOI22_X1 U23741 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n22363), .B1(
        n22369), .B2(n22181), .ZN(n22168) );
  OAI211_X1 U23742 ( .C1(n22184), .C2(n22366), .A(n22169), .B(n22168), .ZN(
        P1_U3123) );
  AOI22_X1 U23743 ( .A1(n22180), .A2(n22368), .B1(n22367), .B2(n22181), .ZN(
        n22171) );
  AOI22_X1 U23744 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n22370), .B1(
        n22369), .B2(n22175), .ZN(n22170) );
  OAI211_X1 U23745 ( .C1(n22374), .C2(n22172), .A(n22171), .B(n22170), .ZN(
        P1_U3131) );
  AOI22_X1 U23746 ( .A1(n22180), .A2(n22376), .B1(n22179), .B2(n22375), .ZN(
        n22174) );
  AOI22_X1 U23747 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n22377), .B1(
        n22384), .B2(n22181), .ZN(n22173) );
  OAI211_X1 U23748 ( .C1(n22184), .C2(n22380), .A(n22174), .B(n22173), .ZN(
        P1_U3139) );
  AOI22_X1 U23749 ( .A1(n22180), .A2(n22382), .B1(n22179), .B2(n22381), .ZN(
        n22177) );
  AOI22_X1 U23750 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n22385), .B1(
        n22384), .B2(n22175), .ZN(n22176) );
  OAI211_X1 U23751 ( .C1(n22178), .C2(n22397), .A(n22177), .B(n22176), .ZN(
        P1_U3147) );
  AOI22_X1 U23752 ( .A1(n22180), .A2(n22390), .B1(n22179), .B2(n22388), .ZN(
        n22183) );
  AOI22_X1 U23753 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n22394), .B1(
        n22393), .B2(n22181), .ZN(n22182) );
  OAI211_X1 U23754 ( .C1(n22184), .C2(n22397), .A(n22183), .B(n22182), .ZN(
        P1_U3155) );
  AOI22_X1 U23755 ( .A1(n22212), .A2(n22310), .B1(n22393), .B2(n11068), .ZN(
        n22186) );
  AOI22_X1 U23756 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n22311), .B1(
        n22317), .B2(n11074), .ZN(n22185) );
  OAI211_X1 U23757 ( .C1(n22314), .C2(n22205), .A(n22186), .B(n22185), .ZN(
        P1_U3036) );
  AOI22_X1 U23758 ( .A1(n22212), .A2(n22316), .B1(n22211), .B2(n22315), .ZN(
        n22188) );
  AOI22_X1 U23759 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n22318), .B1(
        n22317), .B2(n11068), .ZN(n22187) );
  OAI211_X1 U23760 ( .C1(n11073), .C2(n22321), .A(n22188), .B(n22187), .ZN(
        P1_U3044) );
  AOI22_X1 U23761 ( .A1(n22323), .A2(n11068), .B1(n22212), .B2(n22322), .ZN(
        n22190) );
  AOI22_X1 U23762 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n22324), .B1(
        n22330), .B2(n11074), .ZN(n22189) );
  OAI211_X1 U23763 ( .C1(n22327), .C2(n22205), .A(n22190), .B(n22189), .ZN(
        P1_U3052) );
  AOI22_X1 U23764 ( .A1(n22330), .A2(n11068), .B1(n22212), .B2(n22328), .ZN(
        n22192) );
  AOI22_X1 U23765 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n22331), .B1(
        n22329), .B2(n11074), .ZN(n22191) );
  OAI211_X1 U23766 ( .C1(n22334), .C2(n22205), .A(n22192), .B(n22191), .ZN(
        P1_U3060) );
  AOI22_X1 U23767 ( .A1(n22212), .A2(n22336), .B1(n11068), .B2(n22335), .ZN(
        n22194) );
  AOI22_X1 U23768 ( .A1(n22338), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n22337), .B2(n11074), .ZN(n22193) );
  OAI211_X1 U23769 ( .C1(n22341), .C2(n22205), .A(n22194), .B(n22193), .ZN(
        P1_U3084) );
  AOI22_X1 U23770 ( .A1(n22212), .A2(n22343), .B1(n22211), .B2(n22342), .ZN(
        n22196) );
  AOI22_X1 U23771 ( .A1(n22345), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n22344), .B2(n11068), .ZN(n22195) );
  OAI211_X1 U23772 ( .C1(n11073), .C2(n22353), .A(n22196), .B(n22195), .ZN(
        P1_U3100) );
  AOI22_X1 U23773 ( .A1(n22212), .A2(n22349), .B1(n22211), .B2(n22348), .ZN(
        n22198) );
  AOI22_X1 U23774 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n22350), .B1(
        n22354), .B2(n11074), .ZN(n22197) );
  OAI211_X1 U23775 ( .C1(n11067), .C2(n22353), .A(n22198), .B(n22197), .ZN(
        P1_U3108) );
  AOI22_X1 U23776 ( .A1(n22212), .A2(n22355), .B1(n22354), .B2(n11068), .ZN(
        n22200) );
  AOI22_X1 U23777 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n22357), .B1(
        n22356), .B2(n11074), .ZN(n22199) );
  OAI211_X1 U23778 ( .C1(n22360), .C2(n22205), .A(n22200), .B(n22199), .ZN(
        P1_U3116) );
  AOI22_X1 U23779 ( .A1(n22212), .A2(n22362), .B1(n22211), .B2(n22361), .ZN(
        n22202) );
  AOI22_X1 U23780 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n22363), .B1(
        n22369), .B2(n11074), .ZN(n22201) );
  OAI211_X1 U23781 ( .C1(n11067), .C2(n22366), .A(n22202), .B(n22201), .ZN(
        P1_U3124) );
  AOI22_X1 U23782 ( .A1(n22212), .A2(n22368), .B1(n22367), .B2(n11074), .ZN(
        n22204) );
  AOI22_X1 U23783 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n22370), .B1(
        n22369), .B2(n11068), .ZN(n22203) );
  OAI211_X1 U23784 ( .C1(n22374), .C2(n22205), .A(n22204), .B(n22203), .ZN(
        P1_U3132) );
  AOI22_X1 U23785 ( .A1(n22212), .A2(n22376), .B1(n22211), .B2(n22375), .ZN(
        n22207) );
  AOI22_X1 U23786 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n22377), .B1(
        n22384), .B2(n11074), .ZN(n22206) );
  OAI211_X1 U23787 ( .C1(n11067), .C2(n22380), .A(n22207), .B(n22206), .ZN(
        P1_U3140) );
  AOI22_X1 U23788 ( .A1(n22212), .A2(n22382), .B1(n22211), .B2(n22381), .ZN(
        n22210) );
  AOI22_X1 U23789 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n22385), .B1(
        n22384), .B2(n11068), .ZN(n22209) );
  OAI211_X1 U23790 ( .C1(n11073), .C2(n22397), .A(n22210), .B(n22209), .ZN(
        P1_U3148) );
  AOI22_X1 U23791 ( .A1(n22212), .A2(n22390), .B1(n22211), .B2(n22388), .ZN(
        n22215) );
  AOI22_X1 U23792 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n22394), .B1(
        n22393), .B2(n11074), .ZN(n22214) );
  OAI211_X1 U23793 ( .C1(n11067), .C2(n22397), .A(n22215), .B(n22214), .ZN(
        P1_U3156) );
  AOI22_X1 U23794 ( .A1(n22243), .A2(n22310), .B1(n22393), .B2(n11066), .ZN(
        n22217) );
  AOI22_X1 U23795 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n22311), .B1(
        n22317), .B2(n11084), .ZN(n22216) );
  OAI211_X1 U23796 ( .C1(n22314), .C2(n22236), .A(n22217), .B(n22216), .ZN(
        P1_U3037) );
  AOI22_X1 U23797 ( .A1(n22243), .A2(n22316), .B1(n22242), .B2(n22315), .ZN(
        n22219) );
  AOI22_X1 U23798 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n22318), .B1(
        n22317), .B2(n11066), .ZN(n22218) );
  OAI211_X1 U23799 ( .C1(n11083), .C2(n22321), .A(n22219), .B(n22218), .ZN(
        P1_U3045) );
  AOI22_X1 U23800 ( .A1(n22323), .A2(n11066), .B1(n22243), .B2(n22322), .ZN(
        n22221) );
  AOI22_X1 U23801 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n22324), .B1(
        n22330), .B2(n11084), .ZN(n22220) );
  OAI211_X1 U23802 ( .C1(n22327), .C2(n22236), .A(n22221), .B(n22220), .ZN(
        P1_U3053) );
  AOI22_X1 U23803 ( .A1(n22329), .A2(n11084), .B1(n22243), .B2(n22328), .ZN(
        n22223) );
  AOI22_X1 U23804 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n22331), .B1(
        n22330), .B2(n11066), .ZN(n22222) );
  OAI211_X1 U23805 ( .C1(n22334), .C2(n22236), .A(n22223), .B(n22222), .ZN(
        P1_U3061) );
  AOI22_X1 U23806 ( .A1(n22243), .A2(n22336), .B1(n11066), .B2(n22335), .ZN(
        n22225) );
  AOI22_X1 U23807 ( .A1(n22338), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n22337), .B2(n11084), .ZN(n22224) );
  OAI211_X1 U23808 ( .C1(n22341), .C2(n22236), .A(n22225), .B(n22224), .ZN(
        P1_U3085) );
  AOI22_X1 U23809 ( .A1(n22243), .A2(n22343), .B1(n22242), .B2(n22342), .ZN(
        n22227) );
  AOI22_X1 U23810 ( .A1(n22345), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n22344), .B2(n11066), .ZN(n22226) );
  OAI211_X1 U23811 ( .C1(n11083), .C2(n22353), .A(n22227), .B(n22226), .ZN(
        P1_U3101) );
  AOI22_X1 U23812 ( .A1(n22243), .A2(n22349), .B1(n22242), .B2(n22348), .ZN(
        n22229) );
  AOI22_X1 U23813 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n22350), .B1(
        n22354), .B2(n11084), .ZN(n22228) );
  OAI211_X1 U23814 ( .C1(n11065), .C2(n22353), .A(n22229), .B(n22228), .ZN(
        P1_U3109) );
  AOI22_X1 U23815 ( .A1(n22243), .A2(n22355), .B1(n22354), .B2(n11066), .ZN(
        n22231) );
  AOI22_X1 U23816 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n22357), .B1(
        n22356), .B2(n11084), .ZN(n22230) );
  OAI211_X1 U23817 ( .C1(n22360), .C2(n22236), .A(n22231), .B(n22230), .ZN(
        P1_U3117) );
  AOI22_X1 U23818 ( .A1(n22243), .A2(n22362), .B1(n22242), .B2(n22361), .ZN(
        n22233) );
  AOI22_X1 U23819 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n22363), .B1(
        n22369), .B2(n11084), .ZN(n22232) );
  OAI211_X1 U23820 ( .C1(n11065), .C2(n22366), .A(n22233), .B(n22232), .ZN(
        P1_U3125) );
  AOI22_X1 U23821 ( .A1(n22243), .A2(n22368), .B1(n22367), .B2(n11084), .ZN(
        n22235) );
  AOI22_X1 U23822 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n22370), .B1(
        n22369), .B2(n11066), .ZN(n22234) );
  OAI211_X1 U23823 ( .C1(n22374), .C2(n22236), .A(n22235), .B(n22234), .ZN(
        P1_U3133) );
  AOI22_X1 U23824 ( .A1(n22243), .A2(n22376), .B1(n22242), .B2(n22375), .ZN(
        n22238) );
  AOI22_X1 U23825 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n22377), .B1(
        n22384), .B2(n11084), .ZN(n22237) );
  OAI211_X1 U23826 ( .C1(n11065), .C2(n22380), .A(n22238), .B(n22237), .ZN(
        P1_U3141) );
  AOI22_X1 U23827 ( .A1(n22243), .A2(n22382), .B1(n22242), .B2(n22381), .ZN(
        n22241) );
  AOI22_X1 U23828 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n22385), .B1(
        n22384), .B2(n11066), .ZN(n22240) );
  OAI211_X1 U23829 ( .C1(n11083), .C2(n22397), .A(n22241), .B(n22240), .ZN(
        P1_U3149) );
  AOI22_X1 U23830 ( .A1(n22243), .A2(n22390), .B1(n22242), .B2(n22388), .ZN(
        n22246) );
  AOI22_X1 U23831 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n22394), .B1(
        n22393), .B2(n11084), .ZN(n22245) );
  OAI211_X1 U23832 ( .C1(n11065), .C2(n22397), .A(n22246), .B(n22245), .ZN(
        P1_U3157) );
  AOI22_X1 U23833 ( .A1(n22274), .A2(n22310), .B1(n22393), .B2(n22270), .ZN(
        n22248) );
  AOI22_X1 U23834 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n22311), .B1(
        n22317), .B2(n11076), .ZN(n22247) );
  OAI211_X1 U23835 ( .C1(n22314), .C2(n22267), .A(n22248), .B(n22247), .ZN(
        P1_U3038) );
  AOI22_X1 U23836 ( .A1(n22274), .A2(n22316), .B1(n22273), .B2(n22315), .ZN(
        n22250) );
  AOI22_X1 U23837 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n22318), .B1(
        n22317), .B2(n22270), .ZN(n22249) );
  OAI211_X1 U23838 ( .C1(n11075), .C2(n22321), .A(n22250), .B(n22249), .ZN(
        P1_U3046) );
  AOI22_X1 U23839 ( .A1(n22323), .A2(n22270), .B1(n22274), .B2(n22322), .ZN(
        n22252) );
  AOI22_X1 U23840 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n22324), .B1(
        n22330), .B2(n11076), .ZN(n22251) );
  OAI211_X1 U23841 ( .C1(n22327), .C2(n22267), .A(n22252), .B(n22251), .ZN(
        P1_U3054) );
  AOI22_X1 U23842 ( .A1(n22330), .A2(n22270), .B1(n22274), .B2(n22328), .ZN(
        n22254) );
  AOI22_X1 U23843 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n22331), .B1(
        n22329), .B2(n11076), .ZN(n22253) );
  OAI211_X1 U23844 ( .C1(n22334), .C2(n22267), .A(n22254), .B(n22253), .ZN(
        P1_U3062) );
  AOI22_X1 U23845 ( .A1(n22274), .A2(n22336), .B1(n22337), .B2(n11076), .ZN(
        n22256) );
  AOI22_X1 U23846 ( .A1(n22338), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n22270), .B2(n22335), .ZN(n22255) );
  OAI211_X1 U23847 ( .C1(n22341), .C2(n22267), .A(n22256), .B(n22255), .ZN(
        P1_U3086) );
  AOI22_X1 U23848 ( .A1(n22274), .A2(n22343), .B1(n22273), .B2(n22342), .ZN(
        n22258) );
  AOI22_X1 U23849 ( .A1(n22345), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n22344), .B2(n22270), .ZN(n22257) );
  OAI211_X1 U23850 ( .C1(n11075), .C2(n22353), .A(n22258), .B(n22257), .ZN(
        P1_U3102) );
  AOI22_X1 U23851 ( .A1(n22274), .A2(n22349), .B1(n22273), .B2(n22348), .ZN(
        n22260) );
  AOI22_X1 U23852 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n22350), .B1(
        n22354), .B2(n11076), .ZN(n22259) );
  OAI211_X1 U23853 ( .C1(n22278), .C2(n22353), .A(n22260), .B(n22259), .ZN(
        P1_U3110) );
  AOI22_X1 U23854 ( .A1(n22274), .A2(n22355), .B1(n22354), .B2(n22270), .ZN(
        n22262) );
  AOI22_X1 U23855 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n22357), .B1(
        n22356), .B2(n11076), .ZN(n22261) );
  OAI211_X1 U23856 ( .C1(n22360), .C2(n22267), .A(n22262), .B(n22261), .ZN(
        P1_U3118) );
  AOI22_X1 U23857 ( .A1(n22274), .A2(n22362), .B1(n22273), .B2(n22361), .ZN(
        n22264) );
  AOI22_X1 U23858 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n22363), .B1(
        n22369), .B2(n11076), .ZN(n22263) );
  OAI211_X1 U23859 ( .C1(n22278), .C2(n22366), .A(n22264), .B(n22263), .ZN(
        P1_U3126) );
  AOI22_X1 U23860 ( .A1(n22274), .A2(n22368), .B1(n22367), .B2(n11076), .ZN(
        n22266) );
  AOI22_X1 U23861 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n22370), .B1(
        n22369), .B2(n22270), .ZN(n22265) );
  OAI211_X1 U23862 ( .C1(n22374), .C2(n22267), .A(n22266), .B(n22265), .ZN(
        P1_U3134) );
  AOI22_X1 U23863 ( .A1(n22274), .A2(n22376), .B1(n22273), .B2(n22375), .ZN(
        n22269) );
  AOI22_X1 U23864 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n22377), .B1(
        n22384), .B2(n11076), .ZN(n22268) );
  OAI211_X1 U23865 ( .C1(n22278), .C2(n22380), .A(n22269), .B(n22268), .ZN(
        P1_U3142) );
  AOI22_X1 U23866 ( .A1(n22274), .A2(n22382), .B1(n22273), .B2(n22381), .ZN(
        n22272) );
  AOI22_X1 U23867 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n22385), .B1(
        n22384), .B2(n22270), .ZN(n22271) );
  OAI211_X1 U23868 ( .C1(n11075), .C2(n22397), .A(n22272), .B(n22271), .ZN(
        P1_U3150) );
  AOI22_X1 U23869 ( .A1(n22274), .A2(n22390), .B1(n22273), .B2(n22388), .ZN(
        n22277) );
  AOI22_X1 U23870 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n22394), .B1(
        n22393), .B2(n11076), .ZN(n22276) );
  OAI211_X1 U23871 ( .C1(n22278), .C2(n22397), .A(n22277), .B(n22276), .ZN(
        P1_U3158) );
  AOI22_X1 U23872 ( .A1(n22306), .A2(n22310), .B1(n22393), .B2(n11064), .ZN(
        n22280) );
  AOI22_X1 U23873 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n22311), .B1(
        n22317), .B2(n11082), .ZN(n22279) );
  OAI211_X1 U23874 ( .C1(n22314), .C2(n22299), .A(n22280), .B(n22279), .ZN(
        P1_U3039) );
  AOI22_X1 U23875 ( .A1(n22306), .A2(n22316), .B1(n22305), .B2(n22315), .ZN(
        n22282) );
  AOI22_X1 U23876 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n22318), .B1(
        n22317), .B2(n11064), .ZN(n22281) );
  OAI211_X1 U23877 ( .C1(n11081), .C2(n22321), .A(n22282), .B(n22281), .ZN(
        P1_U3047) );
  AOI22_X1 U23878 ( .A1(n22330), .A2(n11082), .B1(n22306), .B2(n22322), .ZN(
        n22284) );
  AOI22_X1 U23879 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n22324), .B1(
        n22323), .B2(n11064), .ZN(n22283) );
  OAI211_X1 U23880 ( .C1(n22327), .C2(n22299), .A(n22284), .B(n22283), .ZN(
        P1_U3055) );
  AOI22_X1 U23881 ( .A1(n22330), .A2(n11064), .B1(n22306), .B2(n22328), .ZN(
        n22286) );
  AOI22_X1 U23882 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n22331), .B1(
        n22329), .B2(n11082), .ZN(n22285) );
  OAI211_X1 U23883 ( .C1(n22334), .C2(n22299), .A(n22286), .B(n22285), .ZN(
        P1_U3063) );
  AOI22_X1 U23884 ( .A1(n22306), .A2(n22336), .B1(n11064), .B2(n22335), .ZN(
        n22288) );
  AOI22_X1 U23885 ( .A1(n22338), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n22337), .B2(n11082), .ZN(n22287) );
  OAI211_X1 U23886 ( .C1(n22341), .C2(n22299), .A(n22288), .B(n22287), .ZN(
        P1_U3087) );
  AOI22_X1 U23887 ( .A1(n22306), .A2(n22343), .B1(n22305), .B2(n22342), .ZN(
        n22290) );
  AOI22_X1 U23888 ( .A1(n22345), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n22344), .B2(n11064), .ZN(n22289) );
  OAI211_X1 U23889 ( .C1(n11081), .C2(n22353), .A(n22290), .B(n22289), .ZN(
        P1_U3103) );
  AOI22_X1 U23890 ( .A1(n22306), .A2(n22349), .B1(n22305), .B2(n22348), .ZN(
        n22292) );
  AOI22_X1 U23891 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n22350), .B1(
        n22354), .B2(n11082), .ZN(n22291) );
  OAI211_X1 U23892 ( .C1(n11063), .C2(n22353), .A(n22292), .B(n22291), .ZN(
        P1_U3111) );
  AOI22_X1 U23893 ( .A1(n22306), .A2(n22355), .B1(n22354), .B2(n11064), .ZN(
        n22294) );
  AOI22_X1 U23894 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n22357), .B1(
        n22356), .B2(n11082), .ZN(n22293) );
  OAI211_X1 U23895 ( .C1(n22360), .C2(n22299), .A(n22294), .B(n22293), .ZN(
        P1_U3119) );
  AOI22_X1 U23896 ( .A1(n22306), .A2(n22362), .B1(n22305), .B2(n22361), .ZN(
        n22296) );
  AOI22_X1 U23897 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n22363), .B1(
        n22369), .B2(n11082), .ZN(n22295) );
  OAI211_X1 U23898 ( .C1(n11063), .C2(n22366), .A(n22296), .B(n22295), .ZN(
        P1_U3127) );
  AOI22_X1 U23899 ( .A1(n22306), .A2(n22368), .B1(n22367), .B2(n11082), .ZN(
        n22298) );
  AOI22_X1 U23900 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n22370), .B1(
        n22369), .B2(n11064), .ZN(n22297) );
  OAI211_X1 U23901 ( .C1(n22374), .C2(n22299), .A(n22298), .B(n22297), .ZN(
        P1_U3135) );
  AOI22_X1 U23902 ( .A1(n22306), .A2(n22376), .B1(n22305), .B2(n22375), .ZN(
        n22301) );
  AOI22_X1 U23903 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n22377), .B1(
        n22384), .B2(n11082), .ZN(n22300) );
  OAI211_X1 U23904 ( .C1(n11063), .C2(n22380), .A(n22301), .B(n22300), .ZN(
        P1_U3143) );
  AOI22_X1 U23905 ( .A1(n22306), .A2(n22382), .B1(n22305), .B2(n22381), .ZN(
        n22304) );
  AOI22_X1 U23906 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n22385), .B1(
        n22384), .B2(n11064), .ZN(n22303) );
  OAI211_X1 U23907 ( .C1(n11081), .C2(n22397), .A(n22304), .B(n22303), .ZN(
        P1_U3151) );
  AOI22_X1 U23908 ( .A1(n22306), .A2(n22390), .B1(n22305), .B2(n22388), .ZN(
        n22309) );
  AOI22_X1 U23909 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n22394), .B1(
        n22393), .B2(n11082), .ZN(n22308) );
  OAI211_X1 U23910 ( .C1(n11063), .C2(n22397), .A(n22309), .B(n22308), .ZN(
        P1_U3159) );
  AOI22_X1 U23911 ( .A1(n22391), .A2(n22310), .B1(n22393), .B2(n11060), .ZN(
        n22313) );
  AOI22_X1 U23912 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n22311), .B1(
        n22317), .B2(n11078), .ZN(n22312) );
  OAI211_X1 U23913 ( .C1(n22314), .C2(n22373), .A(n22313), .B(n22312), .ZN(
        P1_U3040) );
  AOI22_X1 U23914 ( .A1(n22391), .A2(n22316), .B1(n22389), .B2(n22315), .ZN(
        n22320) );
  AOI22_X1 U23915 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n22318), .B1(
        n22317), .B2(n11060), .ZN(n22319) );
  OAI211_X1 U23916 ( .C1(n11077), .C2(n22321), .A(n22320), .B(n22319), .ZN(
        P1_U3048) );
  AOI22_X1 U23917 ( .A1(n22323), .A2(n11060), .B1(n22391), .B2(n22322), .ZN(
        n22326) );
  AOI22_X1 U23918 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n22324), .B1(
        n22330), .B2(n11078), .ZN(n22325) );
  OAI211_X1 U23919 ( .C1(n22327), .C2(n22373), .A(n22326), .B(n22325), .ZN(
        P1_U3056) );
  AOI22_X1 U23920 ( .A1(n22329), .A2(n11078), .B1(n22391), .B2(n22328), .ZN(
        n22333) );
  AOI22_X1 U23921 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n22331), .B1(
        n22330), .B2(n11060), .ZN(n22332) );
  OAI211_X1 U23922 ( .C1(n22334), .C2(n22373), .A(n22333), .B(n22332), .ZN(
        P1_U3064) );
  AOI22_X1 U23923 ( .A1(n22391), .A2(n22336), .B1(n11060), .B2(n22335), .ZN(
        n22340) );
  AOI22_X1 U23924 ( .A1(n22338), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n22337), .B2(n11078), .ZN(n22339) );
  OAI211_X1 U23925 ( .C1(n22341), .C2(n22373), .A(n22340), .B(n22339), .ZN(
        P1_U3088) );
  AOI22_X1 U23926 ( .A1(n22391), .A2(n22343), .B1(n22389), .B2(n22342), .ZN(
        n22347) );
  AOI22_X1 U23927 ( .A1(n22345), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n22344), .B2(n11060), .ZN(n22346) );
  OAI211_X1 U23928 ( .C1(n11077), .C2(n22353), .A(n22347), .B(n22346), .ZN(
        P1_U3104) );
  AOI22_X1 U23929 ( .A1(n22391), .A2(n22349), .B1(n22389), .B2(n22348), .ZN(
        n22352) );
  AOI22_X1 U23930 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n22350), .B1(
        n22354), .B2(n11078), .ZN(n22351) );
  OAI211_X1 U23931 ( .C1(n11059), .C2(n22353), .A(n22352), .B(n22351), .ZN(
        P1_U3112) );
  AOI22_X1 U23932 ( .A1(n22391), .A2(n22355), .B1(n22354), .B2(n11060), .ZN(
        n22359) );
  AOI22_X1 U23933 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n22357), .B1(
        n22356), .B2(n11078), .ZN(n22358) );
  OAI211_X1 U23934 ( .C1(n22360), .C2(n22373), .A(n22359), .B(n22358), .ZN(
        P1_U3120) );
  AOI22_X1 U23935 ( .A1(n22391), .A2(n22362), .B1(n22389), .B2(n22361), .ZN(
        n22365) );
  AOI22_X1 U23936 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n22363), .B1(
        n22369), .B2(n11078), .ZN(n22364) );
  OAI211_X1 U23937 ( .C1(n11059), .C2(n22366), .A(n22365), .B(n22364), .ZN(
        P1_U3128) );
  AOI22_X1 U23938 ( .A1(n22391), .A2(n22368), .B1(n22367), .B2(n11078), .ZN(
        n22372) );
  AOI22_X1 U23939 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n22370), .B1(
        n22369), .B2(n11060), .ZN(n22371) );
  OAI211_X1 U23940 ( .C1(n22374), .C2(n22373), .A(n22372), .B(n22371), .ZN(
        P1_U3136) );
  AOI22_X1 U23941 ( .A1(n22391), .A2(n22376), .B1(n22389), .B2(n22375), .ZN(
        n22379) );
  AOI22_X1 U23942 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n22377), .B1(
        n22384), .B2(n11078), .ZN(n22378) );
  OAI211_X1 U23943 ( .C1(n11059), .C2(n22380), .A(n22379), .B(n22378), .ZN(
        P1_U3144) );
  AOI22_X1 U23944 ( .A1(n22391), .A2(n22382), .B1(n22389), .B2(n22381), .ZN(
        n22387) );
  AOI22_X1 U23945 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n22385), .B1(
        n22384), .B2(n11060), .ZN(n22386) );
  OAI211_X1 U23946 ( .C1(n11077), .C2(n22397), .A(n22387), .B(n22386), .ZN(
        P1_U3152) );
  AOI22_X1 U23947 ( .A1(n22391), .A2(n22390), .B1(n22389), .B2(n22388), .ZN(
        n22396) );
  AOI22_X1 U23948 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n22394), .B1(
        n22393), .B2(n11078), .ZN(n22395) );
  OAI211_X1 U23949 ( .C1(n11059), .C2(n22397), .A(n22396), .B(n22395), .ZN(
        P1_U3160) );
  INV_X1 U23950 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n22400) );
  AOI22_X1 U23951 ( .A1(n22401), .A2(n22400), .B1(n22399), .B2(n22398), .ZN(
        P1_U3486) );
  AND2_X1 U11188 ( .A1(n12446), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11091) );
  AND2_X1 U11458 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15212) );
  OR2_X1 U13079 ( .A1(n11496), .A2(n11495), .ZN(n11512) );
  AND2_X1 U12465 ( .A1(n14464), .A2(n14462), .ZN(n16633) );
  CLKBUF_X1 U11108 ( .A(n19793), .Z(n10958) );
  CLKBUF_X1 U11130 ( .A(n12808), .Z(n13526) );
  CLKBUF_X3 U11135 ( .A(n11370), .Z(n14483) );
  NOR2_X1 U11145 ( .A1(n11526), .A2(n11525), .ZN(n11578) );
  AND2_X1 U11146 ( .A1(n16728), .A2(n16729), .ZN(n14511) );
  NAND2_X1 U11168 ( .A1(n11321), .A2(n11322), .ZN(n11379) );
  AOI21_X2 U11171 ( .B1(n10994), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n11437), .ZN(n11451) );
  CLKBUF_X1 U11173 ( .A(n13790), .Z(n20370) );
  CLKBUF_X1 U11179 ( .A(n13126), .Z(n22013) );
  AND4_X2 U11180 ( .A1(n12535), .A2(n12534), .A3(n12533), .A4(n12532), .ZN(
        n12966) );
  OR2_X1 U11416 ( .A1(n14461), .A2(n14460), .ZN(n14464) );
  XNOR2_X1 U11477 ( .A(n14396), .B(n11228), .ZN(n16660) );
  CLKBUF_X1 U11482 ( .A(n11973), .Z(n11008) );
  CLKBUF_X1 U11509 ( .A(n12601), .Z(n14745) );
  CLKBUF_X1 U11510 ( .A(n15382), .Z(n11019) );
  CLKBUF_X1 U11528 ( .A(n16784), .Z(n16785) );
  CLKBUF_X1 U11578 ( .A(n18525), .Z(n18532) );
  CLKBUF_X1 U11776 ( .A(n20328), .Z(n20332) );
  CLKBUF_X1 U12235 ( .A(n19095), .Z(n19257) );
  AND2_X2 U12236 ( .A1(n11969), .A2(n19459), .ZN(n11983) );
  CLKBUF_X1 U12238 ( .A(n21489), .Z(n20279) );
endmodule

