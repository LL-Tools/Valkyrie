

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944;

  OAI21_X1 U2387 ( .B1(n3368), .B2(n3367), .A(n3366), .ZN(n3387) );
  INV_X2 U2388 ( .A(n3016), .ZN(n3674) );
  OAI22_X2 U2389 ( .A1(n3565), .A2(n2341), .B1(n2343), .B2(n2187), .ZN(n3740)
         );
  INV_X2 U2390 ( .A(n3675), .ZN(n3639) );
  CLKBUF_X2 U2391 ( .A(n2463), .Z(n2152) );
  AND4_X1 U2392 ( .A1(n2451), .A2(n2452), .A3(n2449), .A4(n2450), .ZN(n3029)
         );
  NAND2_X1 U2393 ( .A1(n3621), .A2(n3752), .ZN(n3724) );
  INV_X1 U2394 ( .A(IR_REG_31__SCAN_IN), .ZN(n2846) );
  BUF_X4 U2395 ( .A(n2468), .Z(n2145) );
  NAND2_X1 U2396 ( .A1(n2431), .A2(n2844), .ZN(n2468) );
  AOI22_X2 U2397 ( .A1(n3387), .A2(n3386), .B1(n3385), .B2(n3384), .ZN(n3393)
         );
  XNOR2_X2 U2398 ( .A(n2424), .B(IR_REG_30__SCAN_IN), .ZN(n2848) );
  OAI21_X2 U2399 ( .B1(n3646), .B2(n3647), .A(n3648), .ZN(n3565) );
  NAND2_X2 U2400 ( .A1(n2222), .A2(n2354), .ZN(n3646) );
  CLKBUF_X3 U2401 ( .A(n3631), .Z(n2146) );
  AND2_X1 U2402 ( .A1(n3052), .A2(n3012), .ZN(n3631) );
  NAND2_X1 U2403 ( .A1(n2466), .A2(n2397), .ZN(n3529) );
  NAND4_X1 U2404 ( .A1(n2462), .A2(n2461), .A3(n2460), .A4(n2459), .ZN(n3998)
         );
  BUF_X2 U2405 ( .A(n2463), .Z(n2151) );
  MUX2_X1 U2406 ( .A(n4915), .B(n3543), .S(n4657), .Z(n3544) );
  AND2_X1 U2407 ( .A1(n2296), .A2(n2195), .ZN(n4124) );
  OR2_X1 U2408 ( .A1(n4153), .A2(n3882), .ZN(n4136) );
  NAND2_X1 U2409 ( .A1(n4371), .A2(n2402), .ZN(n4168) );
  OAI21_X1 U2410 ( .B1(n4227), .B2(n3838), .A(n3842), .ZN(n4208) );
  OR2_X1 U2411 ( .A1(n4251), .A2(n2736), .ZN(n4227) );
  NAND2_X1 U2412 ( .A1(n2306), .A2(n2164), .ZN(n4251) );
  NAND2_X1 U2413 ( .A1(n2375), .A2(n2374), .ZN(n4210) );
  AND2_X1 U2414 ( .A1(n2359), .A2(n3710), .ZN(n2221) );
  AND2_X1 U2415 ( .A1(n2229), .A2(n2228), .ZN(n3294) );
  AND2_X2 U2416 ( .A1(n2824), .A2(n4603), .ZN(n4625) );
  NAND2_X1 U2417 ( .A1(n2482), .A2(n2170), .ZN(n3225) );
  BUF_X2 U2418 ( .A(n2479), .Z(n2148) );
  INV_X2 U2419 ( .A(n2447), .ZN(n2458) );
  AND2_X1 U2420 ( .A1(n3081), .A2(n3117), .ZN(n3537) );
  NAND2_X1 U2421 ( .A1(n2791), .A2(n4501), .ZN(n3012) );
  BUF_X4 U2422 ( .A(n2469), .Z(n2149) );
  INV_X1 U2423 ( .A(n3043), .ZN(n3117) );
  CLKBUF_X1 U2424 ( .A(n2791), .Z(n3978) );
  XNOR2_X1 U2425 ( .A(n2364), .B(IR_REG_20__SCAN_IN), .ZN(n2791) );
  NAND2_X1 U2426 ( .A1(n2774), .A2(n4498), .ZN(n3052) );
  XNOR2_X1 U2427 ( .A(n2717), .B(n2716), .ZN(n4065) );
  NAND2_X1 U2428 ( .A1(n2658), .A2(IR_REG_31__SCAN_IN), .ZN(n2717) );
  AND2_X1 U2429 ( .A1(n2772), .A2(n2771), .ZN(n4498) );
  XNOR2_X1 U2430 ( .A(n2765), .B(n2764), .ZN(n2840) );
  NAND2_X1 U2431 ( .A1(n2425), .A2(IR_REG_31__SCAN_IN), .ZN(n2424) );
  OR2_X1 U2432 ( .A1(n2426), .A2(n2846), .ZN(n2427) );
  OR2_X1 U2433 ( .A1(n2755), .A2(n2400), .ZN(n2440) );
  NAND2_X1 U2434 ( .A1(n2763), .A2(IR_REG_31__SCAN_IN), .ZN(n2765) );
  MUX2_X1 U2435 ( .A(IR_REG_31__SCAN_IN), .B(n2770), .S(IR_REG_26__SCAN_IN), 
        .Z(n2772) );
  NAND2_X1 U2436 ( .A1(n2771), .A2(IR_REG_31__SCAN_IN), .ZN(n2755) );
  AND2_X1 U2437 ( .A1(n2388), .A2(n2300), .ZN(n2299) );
  AND2_X1 U2438 ( .A1(n2388), .A2(n2421), .ZN(n2298) );
  XNOR2_X1 U2439 ( .A(n2448), .B(IR_REG_2__SCAN_IN), .ZN(n4509) );
  AND2_X1 U2440 ( .A1(n2159), .A2(n2389), .ZN(n2388) );
  INV_X2 U2441 ( .A(n2497), .ZN(n2147) );
  NAND2_X1 U2442 ( .A1(n2249), .A2(n2252), .ZN(n4510) );
  AND2_X1 U2443 ( .A1(n2420), .A2(n2421), .ZN(n2232) );
  AND4_X1 U2444 ( .A1(n2419), .A2(n2418), .A3(n2417), .A4(n4878), .ZN(n2420)
         );
  AND2_X1 U2445 ( .A1(n2416), .A2(n2386), .ZN(n2160) );
  AND3_X1 U2446 ( .A1(n2392), .A2(n2422), .A3(n2391), .ZN(n2159) );
  NAND2_X1 U2447 ( .A1(n4893), .A2(n2753), .ZN(n2438) );
  NAND4_X1 U2448 ( .A1(n2414), .A2(n2413), .A3(n2412), .A4(n2411), .ZN(n2415)
         );
  NOR2_X1 U2449 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2422)
         );
  NOR2_X1 U2450 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2413)
         );
  NOR2_X1 U2451 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2412)
         );
  NOR2_X1 U2452 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2411)
         );
  NOR2_X1 U2453 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2417)
         );
  NOR2_X1 U2454 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2419)
         );
  NOR2_X1 U2455 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2418)
         );
  NOR2_X2 U2456 ( .A1(n3417), .A2(n3552), .ZN(n3441) );
  AND2_X4 U2457 ( .A1(n2945), .A2(n3052), .ZN(n3016) );
  NAND2_X1 U2458 ( .A1(n2844), .A2(n2848), .ZN(n2479) );
  NOR2_X2 U2459 ( .A1(n4265), .A2(n4230), .ZN(n4239) );
  OR2_X2 U2460 ( .A1(n4283), .A2(n4263), .ZN(n4265) );
  INV_X2 U2461 ( .A(n2447), .ZN(n2150) );
  OR2_X1 U2462 ( .A1(n2844), .A2(n2848), .ZN(n2447) );
  NAND2_X2 U2463 ( .A1(n4212), .A2(n4198), .ZN(n4200) );
  AND2_X2 U2464 ( .A1(n4239), .A2(n4219), .ZN(n4212) );
  NOR2_X2 U2465 ( .A1(n4398), .A2(n4297), .ZN(n4298) );
  INV_X2 U2466 ( .A(n3101), .ZN(n3023) );
  NAND4_X1 U2467 ( .A1(n3101), .A2(n2456), .A3(n2301), .A4(n2457), .ZN(n3915)
         );
  AND2_X2 U2468 ( .A1(n4155), .A2(n4145), .ZN(n4143) );
  NOR3_X4 U2469 ( .A1(n4200), .A2(n4356), .A3(n2790), .ZN(n4155) );
  AND2_X1 U2470 ( .A1(n4013), .A2(n4014), .ZN(n2261) );
  NAND2_X1 U2471 ( .A1(n2690), .A2(n2384), .ZN(n2296) );
  NAND2_X1 U2472 ( .A1(n4362), .A2(n4145), .ZN(n2384) );
  NAND2_X1 U2473 ( .A1(n3243), .A2(n2290), .ZN(n2289) );
  AND2_X1 U2474 ( .A1(n2371), .A2(n2288), .ZN(n2287) );
  NAND2_X1 U2475 ( .A1(n2290), .A2(n2291), .ZN(n2288) );
  INV_X1 U2476 ( .A(IR_REG_26__SCAN_IN), .ZN(n2392) );
  INV_X1 U2477 ( .A(IR_REG_21__SCAN_IN), .ZN(n2386) );
  INV_X1 U2478 ( .A(n2632), .ZN(n2634) );
  AOI21_X1 U2479 ( .B1(n3322), .B2(n2348), .A(n2176), .ZN(n2347) );
  NAND2_X1 U2480 ( .A1(n3322), .A2(n2350), .ZN(n2349) );
  NAND2_X1 U2481 ( .A1(n3122), .A2(n2396), .ZN(n3123) );
  NAND2_X1 U2482 ( .A1(n3996), .A2(n3016), .ZN(n3122) );
  NAND2_X1 U2483 ( .A1(n2755), .A2(n2438), .ZN(n2439) );
  AND2_X1 U2484 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2400)
         );
  NAND2_X1 U2485 ( .A1(n3591), .A2(n3590), .ZN(n3592) );
  OAI21_X1 U2486 ( .B1(n4509), .B2(REG2_REG_2__SCAN_IN), .A(n2259), .ZN(n4015)
         );
  NAND2_X1 U2487 ( .A1(n4509), .A2(REG2_REG_2__SCAN_IN), .ZN(n2259) );
  AOI22_X1 U2488 ( .A1(n2897), .A2(REG2_REG_3__SCAN_IN), .B1(n4508), .B2(n2896), .ZN(n2898) );
  NAND2_X1 U2489 ( .A1(n2263), .A2(n2262), .ZN(n4556) );
  OR2_X1 U2490 ( .A1(n4043), .A2(n2266), .ZN(n2262) );
  OR2_X1 U2491 ( .A1(n4139), .A2(n4157), .ZN(n2689) );
  INV_X1 U2492 ( .A(n2279), .ZN(n2278) );
  OAI21_X1 U2493 ( .B1(n2162), .B2(n2281), .A(n2623), .ZN(n2279) );
  NAND2_X1 U2494 ( .A1(n3225), .A2(n3536), .ZN(n3924) );
  INV_X1 U2495 ( .A(n2724), .ZN(n3872) );
  AND2_X1 U2496 ( .A1(n2760), .A2(n2759), .ZN(n2977) );
  AND2_X1 U2497 ( .A1(n2708), .A2(n2707), .ZN(n4338) );
  OR2_X1 U2498 ( .A1(n4617), .A2(n4500), .ZN(n3446) );
  INV_X1 U2499 ( .A(IR_REG_29__SCAN_IN), .ZN(n2423) );
  INV_X1 U2500 ( .A(n3225), .ZN(n3132) );
  NAND2_X1 U2501 ( .A1(n2358), .A2(n2356), .ZN(n2355) );
  NAND2_X1 U2502 ( .A1(n3774), .A2(n3555), .ZN(n2356) );
  INV_X1 U2503 ( .A(n2276), .ZN(n2272) );
  INV_X1 U2504 ( .A(n3897), .ZN(n2603) );
  INV_X1 U2505 ( .A(n2372), .ZN(n2371) );
  OAI21_X1 U2506 ( .B1(n2569), .B2(n2373), .A(n2582), .ZN(n2372) );
  NAND2_X1 U2507 ( .A1(n3991), .A2(n3552), .ZN(n2582) );
  INV_X1 U2508 ( .A(n2571), .ZN(n2373) );
  NAND2_X1 U2509 ( .A1(n2178), .A2(n2558), .ZN(n2290) );
  INV_X1 U2510 ( .A(n3936), .ZN(n2319) );
  INV_X1 U2511 ( .A(n3924), .ZN(n2314) );
  INV_X1 U2512 ( .A(n3939), .ZN(n2312) );
  AND2_X1 U2513 ( .A1(n2454), .A2(n2455), .ZN(n2301) );
  AND2_X1 U2514 ( .A1(n2152), .A2(DATAI_20_), .ZN(n4230) );
  AND2_X1 U2515 ( .A1(n4500), .A2(n4501), .ZN(n2979) );
  AND2_X1 U2516 ( .A1(n2160), .A2(n2422), .ZN(n2230) );
  NOR2_X1 U2517 ( .A1(n2415), .A2(IR_REG_13__SCAN_IN), .ZN(n2387) );
  INV_X1 U2518 ( .A(IR_REG_6__SCAN_IN), .ZN(n2521) );
  NOR2_X1 U2519 ( .A1(n3292), .A2(n3291), .ZN(n2351) );
  NOR2_X1 U2520 ( .A1(n3295), .A2(n3293), .ZN(n2348) );
  NOR2_X1 U2521 ( .A1(n2165), .A2(n2191), .ZN(n2225) );
  INV_X1 U2522 ( .A(n2362), .ZN(n2226) );
  INV_X1 U2523 ( .A(n2182), .ZN(n2227) );
  INV_X1 U2524 ( .A(n3806), .ZN(n2340) );
  AOI21_X1 U2525 ( .B1(n3636), .B2(n3998), .A(n2949), .ZN(n2953) );
  AOI21_X1 U2526 ( .B1(n2993), .B2(n3016), .A(n2947), .ZN(n2948) );
  NAND2_X1 U2527 ( .A1(n3467), .A2(n3469), .ZN(n3470) );
  AND2_X1 U2528 ( .A1(n2344), .A2(n3733), .ZN(n2343) );
  OR2_X1 U2529 ( .A1(n2345), .A2(n2187), .ZN(n2341) );
  NAND2_X1 U2530 ( .A1(n3567), .A2(n3818), .ZN(n2344) );
  NAND2_X1 U2531 ( .A1(n3248), .A2(n3247), .ZN(n2228) );
  NAND2_X1 U2532 ( .A1(n3052), .A2(n2857), .ZN(n2989) );
  OR2_X1 U2533 ( .A1(n2682), .A2(n3755), .ZN(n2684) );
  NOR2_X1 U2534 ( .A1(n2595), .A2(n2594), .ZN(n2605) );
  NAND2_X1 U2535 ( .A1(n4018), .A2(n2876), .ZN(n2901) );
  NOR2_X1 U2536 ( .A1(n4012), .A2(n2260), .ZN(n2895) );
  NAND2_X1 U2537 ( .A1(n2961), .A2(REG1_REG_4__SCAN_IN), .ZN(n2960) );
  NOR2_X1 U2538 ( .A1(n2936), .A2(n2255), .ZN(n2254) );
  NOR2_X1 U2539 ( .A1(n2936), .A2(n2965), .ZN(n2253) );
  AND2_X1 U2540 ( .A1(n2257), .A2(n2256), .ZN(n2924) );
  NAND2_X1 U2541 ( .A1(n4506), .A2(REG2_REG_5__SCAN_IN), .ZN(n2256) );
  OR2_X1 U2542 ( .A1(n3173), .A2(n4605), .ZN(n2276) );
  AND2_X1 U2543 ( .A1(n4518), .A2(n2186), .ZN(n2274) );
  NAND2_X1 U2544 ( .A1(n4529), .A2(n3178), .ZN(n4534) );
  NAND2_X1 U2545 ( .A1(n4534), .A2(n4535), .ZN(n4533) );
  NAND2_X1 U2546 ( .A1(n2410), .A2(n2399), .ZN(n2497) );
  INV_X1 U2547 ( .A(IR_REG_4__SCAN_IN), .ZN(n2409) );
  OR2_X1 U2548 ( .A1(n4503), .A2(REG2_REG_13__SCAN_IN), .ZN(n2270) );
  NOR2_X1 U2549 ( .A1(n4556), .A2(n4557), .ZN(n4555) );
  NOR2_X1 U2550 ( .A1(n2242), .A2(n2198), .ZN(n2240) );
  OR2_X1 U2551 ( .A1(n2243), .A2(n2198), .ZN(n2238) );
  AOI21_X1 U2552 ( .B1(n2155), .B2(n3966), .A(n3848), .ZN(n2330) );
  NAND2_X1 U2553 ( .A1(n2304), .A2(n3866), .ZN(n4153) );
  OAI21_X1 U2554 ( .B1(n4208), .B2(n3843), .A(n2744), .ZN(n2304) );
  AOI21_X1 U2555 ( .B1(n4168), .B2(n2681), .A(n2395), .ZN(n4151) );
  INV_X1 U2556 ( .A(n2378), .ZN(n2377) );
  OAI21_X1 U2557 ( .B1(n2650), .B2(n2154), .A(n2659), .ZN(n2378) );
  OR2_X1 U2558 ( .A1(n3511), .A2(n2622), .ZN(n2306) );
  AOI21_X1 U2559 ( .B1(n4322), .B2(n2309), .A(n2308), .ZN(n2307) );
  INV_X1 U2560 ( .A(n3834), .ZN(n2309) );
  NAND2_X1 U2561 ( .A1(n2380), .A2(n2613), .ZN(n2379) );
  INV_X1 U2562 ( .A(n2604), .ZN(n2380) );
  OR2_X1 U2563 ( .A1(n3510), .A2(n3867), .ZN(n3511) );
  NAND2_X1 U2564 ( .A1(n2294), .A2(n3376), .ZN(n2293) );
  NAND2_X1 U2565 ( .A1(n2322), .A2(n2183), .ZN(n2321) );
  INV_X1 U2566 ( .A(n2325), .ZN(n2322) );
  INV_X1 U2567 ( .A(n3930), .ZN(n2326) );
  AND2_X1 U2568 ( .A1(n3931), .A2(n3936), .ZN(n3870) );
  NAND2_X1 U2569 ( .A1(n2502), .A2(n2285), .ZN(n2284) );
  INV_X1 U2570 ( .A(n3527), .ZN(n2316) );
  AND2_X1 U2571 ( .A1(n3923), .A2(n3939), .ZN(n3893) );
  AND2_X1 U2572 ( .A1(n4606), .A2(n4427), .ZN(n4161) );
  INV_X1 U2573 ( .A(n4345), .ZN(n3906) );
  INV_X1 U2574 ( .A(n4162), .ZN(n4362) );
  INV_X1 U2575 ( .A(n4417), .ZN(n3825) );
  INV_X1 U2576 ( .A(n4428), .ZN(n3652) );
  INV_X1 U2577 ( .A(n3066), .ZN(n3140) );
  AND2_X1 U2578 ( .A1(n2791), .A2(n2977), .ZN(n4412) );
  AND2_X1 U2579 ( .A1(n2997), .A2(n2979), .ZN(n4429) );
  AND2_X1 U2580 ( .A1(n2773), .A2(n4498), .ZN(n2850) );
  INV_X1 U2581 ( .A(n2438), .ZN(n2389) );
  NAND2_X1 U2582 ( .A1(n2423), .A2(IR_REG_31__SCAN_IN), .ZN(n2428) );
  AND2_X1 U2583 ( .A1(n2422), .A2(n2391), .ZN(n2390) );
  INV_X1 U2584 ( .A(IR_REG_23__SCAN_IN), .ZN(n2775) );
  INV_X1 U2585 ( .A(IR_REG_19__SCAN_IN), .ZN(n2716) );
  INV_X1 U2586 ( .A(IR_REG_17__SCAN_IN), .ZN(n2352) );
  AND2_X1 U2587 ( .A1(n2250), .A2(n2251), .ZN(n2249) );
  NAND2_X1 U2588 ( .A1(IR_REG_1__SCAN_IN), .A2(n2846), .ZN(n2251) );
  INV_X1 U2589 ( .A(n4399), .ZN(n3745) );
  INV_X1 U2590 ( .A(n3529), .ZN(n3141) );
  INV_X1 U2591 ( .A(n3990), .ZN(n4421) );
  NAND2_X1 U2592 ( .A1(n3166), .A2(n4544), .ZN(n4043) );
  NOR2_X1 U2593 ( .A1(n4084), .A2(n2206), .ZN(n2205) );
  NOR2_X1 U2594 ( .A1(n4082), .A2(n4603), .ZN(n2206) );
  NAND2_X1 U2595 ( .A1(n3872), .A2(n2303), .ZN(n2813) );
  INV_X1 U2596 ( .A(n2812), .ZN(n2303) );
  INV_X2 U2597 ( .A(n4655), .ZN(n4657) );
  NAND2_X1 U2598 ( .A1(n4331), .A2(n2207), .ZN(n4083) );
  OR2_X1 U2599 ( .A1(n2807), .A2(n4077), .ZN(n2207) );
  OR2_X1 U2600 ( .A1(n4084), .A2(n2761), .ZN(n2762) );
  INV_X1 U2601 ( .A(n2351), .ZN(n2350) );
  AOI21_X1 U2602 ( .B1(n2216), .B2(n2219), .A(n2214), .ZN(n2213) );
  INV_X1 U2603 ( .A(n3668), .ZN(n2214) );
  NOR2_X1 U2604 ( .A1(n3605), .A2(n2363), .ZN(n2362) );
  NOR2_X1 U2605 ( .A1(n3567), .A2(n3818), .ZN(n2345) );
  AND2_X1 U2606 ( .A1(n2252), .A2(REG1_REG_1__SCAN_IN), .ZN(n2246) );
  AND2_X1 U2607 ( .A1(n2270), .A2(n4632), .ZN(n2267) );
  OR2_X1 U2608 ( .A1(n4632), .A2(n2270), .ZN(n2268) );
  NAND2_X1 U2609 ( .A1(n2267), .A2(n4042), .ZN(n2265) );
  OR2_X1 U2610 ( .A1(n4042), .A2(n4632), .ZN(n2266) );
  INV_X1 U2611 ( .A(n4060), .ZN(n2241) );
  NAND2_X1 U2612 ( .A1(n2292), .A2(n2558), .ZN(n2291) );
  INV_X1 U2613 ( .A(n2548), .ZN(n2292) );
  INV_X1 U2614 ( .A(n3896), .ZN(n2569) );
  AND2_X1 U2615 ( .A1(n2476), .A2(REG3_REG_5__SCAN_IN), .ZN(n2488) );
  INV_X1 U2616 ( .A(n2487), .ZN(n2285) );
  AND2_X1 U2617 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2476) );
  AND2_X1 U2618 ( .A1(n2978), .A2(n2979), .ZN(n2983) );
  OAI21_X1 U2619 ( .B1(n2330), .B2(n2329), .A(n2709), .ZN(n2328) );
  INV_X1 U2620 ( .A(n3853), .ZN(n2329) );
  NAND2_X1 U2621 ( .A1(n2212), .A2(n4320), .ZN(n4297) );
  NOR2_X1 U2622 ( .A1(n3514), .A2(n4417), .ZN(n2212) );
  INV_X1 U2623 ( .A(n3344), .ZN(n3324) );
  INV_X1 U2624 ( .A(IR_REG_28__SCAN_IN), .ZN(n4893) );
  INV_X1 U2625 ( .A(IR_REG_27__SCAN_IN), .ZN(n2753) );
  INV_X1 U2626 ( .A(IR_REG_25__SCAN_IN), .ZN(n2391) );
  AOI21_X1 U2627 ( .B1(n2717), .B2(n2716), .A(n2846), .ZN(n2364) );
  NOR2_X1 U2628 ( .A1(IR_REG_15__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2633)
         );
  INV_X1 U2629 ( .A(IR_REG_14__SCAN_IN), .ZN(n2611) );
  OR3_X1 U2630 ( .A1(n2546), .A2(IR_REG_7__SCAN_IN), .A3(IR_REG_8__SCAN_IN), 
        .ZN(n2556) );
  CLKBUF_X1 U2631 ( .A(n2497), .Z(n2498) );
  INV_X1 U2632 ( .A(IR_REG_2__SCAN_IN), .ZN(n2408) );
  INV_X1 U2633 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2594) );
  NAND2_X1 U2634 ( .A1(n2357), .A2(n3774), .ZN(n2354) );
  NAND2_X1 U2635 ( .A1(n3556), .A2(n2355), .ZN(n2222) );
  AOI21_X1 U2636 ( .B1(n2185), .B2(n2218), .A(n2217), .ZN(n2216) );
  INV_X1 U2637 ( .A(n3579), .ZN(n2218) );
  INV_X1 U2638 ( .A(n3795), .ZN(n2217) );
  INV_X1 U2639 ( .A(n2185), .ZN(n2219) );
  INV_X1 U2640 ( .A(n2337), .ZN(n2336) );
  OAI21_X1 U2641 ( .B1(n3806), .B2(n2338), .A(n3804), .ZN(n2337) );
  NAND2_X1 U2642 ( .A1(n3723), .A2(n2339), .ZN(n2338) );
  INV_X1 U2643 ( .A(n3722), .ZN(n2339) );
  NAND2_X1 U2644 ( .A1(n2146), .A2(n2993), .ZN(n3014) );
  NAND2_X1 U2645 ( .A1(n3660), .A2(n3617), .ZN(n3751) );
  AOI21_X1 U2646 ( .B1(n2225), .B2(n2227), .A(n2192), .ZN(n2224) );
  NAND2_X1 U2647 ( .A1(n3761), .A2(n2225), .ZN(n2223) );
  INV_X1 U2648 ( .A(n2146), .ZN(n3677) );
  NAND2_X1 U2649 ( .A1(n3761), .A2(n2362), .ZN(n2361) );
  XNOR2_X1 U2650 ( .A(n3020), .B(n3639), .ZN(n3032) );
  OR2_X1 U2651 ( .A1(n2684), .A2(n2406), .ZN(n2692) );
  NAND2_X1 U2652 ( .A1(n2342), .A2(n3567), .ZN(n3817) );
  INV_X1 U2653 ( .A(n3565), .ZN(n2342) );
  NAND2_X1 U2654 ( .A1(n2685), .A2(REG1_REG_4__SCAN_IN), .ZN(n2297) );
  NAND2_X1 U2655 ( .A1(n2302), .A2(REG3_REG_2__SCAN_IN), .ZN(n2449) );
  NAND2_X1 U2656 ( .A1(n2302), .A2(REG3_REG_1__SCAN_IN), .ZN(n2455) );
  OAI211_X1 U2657 ( .C1(n2249), .C2(REG1_REG_1__SCAN_IN), .A(n2245), .B(n2247), 
        .ZN(n4001) );
  NAND2_X1 U2658 ( .A1(n2248), .A2(n3107), .ZN(n2247) );
  NAND2_X1 U2659 ( .A1(n2246), .A2(n2249), .ZN(n2245) );
  INV_X1 U2660 ( .A(n2252), .ZN(n2248) );
  NAND2_X1 U2661 ( .A1(n4001), .A2(n4000), .ZN(n3999) );
  NAND2_X1 U2662 ( .A1(n2940), .A2(n2244), .ZN(n2920) );
  OR2_X1 U2663 ( .A1(n2906), .A2(n3158), .ZN(n2244) );
  AOI22_X1 U2664 ( .A1(n2926), .A2(REG2_REG_6__SCAN_IN), .B1(n4505), .B2(n2925), .ZN(n2928) );
  NAND2_X1 U2665 ( .A1(n4514), .A2(n3175), .ZN(n3177) );
  AOI21_X1 U2666 ( .B1(n2274), .B2(n2272), .A(n2188), .ZN(n2271) );
  INV_X1 U2667 ( .A(n2274), .ZN(n2273) );
  NAND2_X1 U2668 ( .A1(n4533), .A2(n3179), .ZN(n3180) );
  NOR2_X1 U2669 ( .A1(REG1_REG_16__SCAN_IN), .A2(n4578), .ZN(n4577) );
  INV_X1 U2670 ( .A(n4596), .ZN(n2242) );
  NAND2_X1 U2671 ( .A1(n4124), .A2(n2383), .ZN(n2382) );
  NAND2_X1 U2672 ( .A1(n4336), .A2(n4344), .ZN(n2383) );
  NAND2_X1 U2673 ( .A1(n2677), .A2(REG3_REG_23__SCAN_IN), .ZN(n2682) );
  AND2_X1 U2674 ( .A1(n2673), .A2(REG3_REG_22__SCAN_IN), .ZN(n2677) );
  AOI21_X1 U2675 ( .B1(n2163), .B2(n2154), .A(n2189), .ZN(n2374) );
  NAND2_X1 U2676 ( .A1(n4280), .A2(n2163), .ZN(n2375) );
  INV_X1 U2677 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3767) );
  OR2_X1 U2678 ( .A1(n2626), .A2(n2405), .ZN(n2642) );
  AND2_X1 U2679 ( .A1(n3832), .A2(n3833), .ZN(n3897) );
  OR2_X1 U2680 ( .A1(n2574), .A2(n2404), .ZN(n2583) );
  INV_X1 U2681 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3185) );
  OR2_X1 U2682 ( .A1(n2583), .A2(n3185), .ZN(n2595) );
  AOI21_X1 U2683 ( .B1(n2371), .B2(n2373), .A(n2174), .ZN(n2369) );
  NAND2_X1 U2684 ( .A1(n2289), .A2(n2287), .ZN(n2370) );
  NAND2_X1 U2685 ( .A1(n2286), .A2(n2290), .ZN(n2570) );
  OR2_X1 U2686 ( .A1(n3243), .A2(n2291), .ZN(n2286) );
  NAND2_X1 U2687 ( .A1(n2570), .A2(n2569), .ZN(n3400) );
  AND2_X1 U2688 ( .A1(n3911), .A2(n3947), .ZN(n3896) );
  AOI21_X1 U2689 ( .B1(n2321), .B2(n2324), .A(n2319), .ZN(n2318) );
  INV_X1 U2690 ( .A(n2321), .ZN(n2320) );
  AND2_X1 U2691 ( .A1(n2488), .A2(REG3_REG_6__SCAN_IN), .ZN(n2516) );
  NAND2_X1 U2692 ( .A1(n2310), .A2(n2311), .ZN(n3192) );
  AOI21_X1 U2693 ( .B1(n2313), .B2(n2727), .A(n2312), .ZN(n2311) );
  AND2_X1 U2694 ( .A1(n3920), .A2(n3917), .ZN(n3871) );
  NOR2_X1 U2695 ( .A1(n2725), .A2(n2453), .ZN(n2464) );
  AND2_X1 U2696 ( .A1(n4606), .A2(n4429), .ZN(n4313) );
  NOR2_X1 U2697 ( .A1(n2989), .A2(n2983), .ZN(n2821) );
  NOR2_X1 U2698 ( .A1(n4331), .A2(n4333), .ZN(n4330) );
  AND2_X1 U2699 ( .A1(n2152), .A2(DATAI_30_), .ZN(n4333) );
  AND2_X1 U2700 ( .A1(n2151), .A2(DATAI_28_), .ZN(n4092) );
  NOR2_X1 U2701 ( .A1(n4106), .A2(n4092), .ZN(n2807) );
  OR2_X1 U2702 ( .A1(n4125), .A2(n4335), .ZN(n4106) );
  AND2_X1 U2703 ( .A1(n2152), .A2(DATAI_27_), .ZN(n4335) );
  NAND2_X1 U2704 ( .A1(n4143), .A2(n4129), .ZN(n4125) );
  NAND2_X1 U2705 ( .A1(n2151), .A2(DATAI_24_), .ZN(n4157) );
  INV_X1 U2706 ( .A(n4157), .ZN(n4356) );
  NAND2_X1 U2707 ( .A1(n2151), .A2(DATAI_22_), .ZN(n4198) );
  NAND2_X1 U2708 ( .A1(n4298), .A2(n4284), .ZN(n4283) );
  INV_X1 U2709 ( .A(n2212), .ZN(n4312) );
  AND2_X1 U2710 ( .A1(n3441), .A2(n3780), .ZN(n3459) );
  OR2_X1 U2711 ( .A1(n3409), .A2(n3403), .ZN(n3417) );
  INV_X1 U2712 ( .A(n3391), .ZN(n3394) );
  NOR2_X1 U2713 ( .A1(n2209), .A2(n3369), .ZN(n3282) );
  NAND2_X1 U2714 ( .A1(n3196), .A2(n2208), .ZN(n3339) );
  AND2_X1 U2715 ( .A1(n3254), .A2(n3303), .ZN(n2208) );
  NAND2_X1 U2716 ( .A1(n3196), .A2(n3254), .ZN(n3214) );
  INV_X1 U2717 ( .A(n3200), .ZN(n3254) );
  INV_X1 U2718 ( .A(n4432), .ZN(n4357) );
  INV_X1 U2719 ( .A(n3230), .ZN(n3154) );
  NAND2_X1 U2720 ( .A1(n3537), .A2(n3536), .ZN(n3535) );
  NOR2_X2 U2721 ( .A1(n3535), .A2(n3154), .ZN(n3196) );
  NAND2_X1 U2722 ( .A1(n4502), .A2(n2977), .ZN(n4258) );
  NAND2_X1 U2723 ( .A1(n4237), .A2(n3446), .ZN(n4423) );
  INV_X1 U2724 ( .A(n4429), .ZN(n4361) );
  INV_X1 U2725 ( .A(n4258), .ZN(n4427) );
  INV_X1 U2726 ( .A(n2820), .ZN(n2975) );
  INV_X1 U2727 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4862) );
  XNOR2_X1 U2728 ( .A(n2756), .B(IR_REG_28__SCAN_IN), .ZN(n2997) );
  NAND2_X1 U2729 ( .A1(n2169), .A2(n2159), .ZN(n2771) );
  NAND2_X1 U2730 ( .A1(n2172), .A2(n2768), .ZN(n2853) );
  NAND2_X1 U2731 ( .A1(n2634), .A2(n2633), .ZN(n2353) );
  INV_X1 U2732 ( .A(IR_REG_3__SCAN_IN), .ZN(n2483) );
  OAI21_X1 U2733 ( .B1(n3294), .B2(n2351), .A(n2346), .ZN(n3323) );
  INV_X1 U2734 ( .A(n2348), .ZN(n2346) );
  INV_X1 U2735 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4672) );
  NAND2_X1 U2736 ( .A1(n2151), .A2(DATAI_23_), .ZN(n4181) );
  OAI21_X1 U2737 ( .B1(n3761), .B2(n2227), .A(n2225), .ZN(n3660) );
  NAND2_X1 U2738 ( .A1(n3393), .A2(n3392), .ZN(n3471) );
  NAND2_X1 U2739 ( .A1(n3050), .A2(n3049), .ZN(n3089) );
  NAND2_X1 U2740 ( .A1(n2335), .A2(n2333), .ZN(n3698) );
  AND2_X1 U2741 ( .A1(n2336), .A2(n2334), .ZN(n2333) );
  INV_X1 U2742 ( .A(n3682), .ZN(n2334) );
  NAND2_X1 U2743 ( .A1(n3761), .A2(n3764), .ZN(n3703) );
  INV_X1 U2744 ( .A(n3483), .ZN(n3715) );
  NAND2_X1 U2745 ( .A1(n2152), .A2(DATAI_25_), .ZN(n4145) );
  INV_X1 U2746 ( .A(n3224), .ZN(n3301) );
  NAND2_X1 U2747 ( .A1(n3129), .A2(n3128), .ZN(n3130) );
  NAND2_X1 U2748 ( .A1(n3125), .A2(n3127), .ZN(n3128) );
  NAND2_X1 U2749 ( .A1(n2361), .A2(n3604), .ZN(n3786) );
  NOR2_X1 U2750 ( .A1(n3034), .A2(n3033), .ZN(n3035) );
  AND2_X1 U2751 ( .A1(n3032), .A2(n3031), .ZN(n3033) );
  INV_X1 U2752 ( .A(n4275), .ZN(n4233) );
  NAND2_X1 U2753 ( .A1(n3740), .A2(n3579), .ZN(n2220) );
  INV_X1 U2754 ( .A(n3995), .ZN(n3345) );
  NAND2_X1 U2755 ( .A1(n2233), .A2(n3723), .ZN(n3808) );
  NAND2_X1 U2756 ( .A1(n3724), .A2(n3722), .ZN(n2233) );
  INV_X1 U2757 ( .A(n3815), .ZN(n3820) );
  INV_X1 U2758 ( .A(n3813), .ZN(n3831) );
  AND3_X1 U2759 ( .A1(n2752), .A2(n2751), .A3(n2750), .ZN(n3861) );
  NAND2_X1 U2760 ( .A1(n2698), .A2(n2697), .ZN(n4345) );
  OR2_X1 U2761 ( .A1(n3641), .A2(n2148), .ZN(n2698) );
  NAND2_X1 U2762 ( .A1(n2445), .A2(n2444), .ZN(n4162) );
  NAND2_X1 U2763 ( .A1(n2496), .A2(n2167), .ZN(n3996) );
  AND3_X1 U2764 ( .A1(n2472), .A2(n2471), .A3(n2470), .ZN(n2397) );
  OR2_X1 U2765 ( .A1(n2148), .A2(n3000), .ZN(n2460) );
  CLKBUF_X2 U2766 ( .A(U4043), .Z(n3997) );
  OAI211_X1 U2767 ( .C1(n4510), .C2(REG2_REG_1__SCAN_IN), .A(n2258), .B(n2168), 
        .ZN(n4014) );
  XNOR2_X1 U2768 ( .A(n2895), .B(n4508), .ZN(n2897) );
  NAND2_X1 U2769 ( .A1(n2960), .A2(n2173), .ZN(n2941) );
  NAND2_X1 U2770 ( .A1(n2941), .A2(n2942), .ZN(n2940) );
  AOI21_X1 U2771 ( .B1(n2959), .B2(REG2_REG_4__SCAN_IN), .A(n2200), .ZN(n2937)
         );
  XNOR2_X1 U2772 ( .A(n2924), .B(n4505), .ZN(n2926) );
  XNOR2_X1 U2773 ( .A(n3160), .B(n3173), .ZN(n3161) );
  NAND2_X1 U2774 ( .A1(n4515), .A2(n4516), .ZN(n4514) );
  NAND2_X1 U2775 ( .A1(n2237), .A2(n2235), .ZN(n4515) );
  NAND2_X1 U2776 ( .A1(n3172), .A2(n2236), .ZN(n2235) );
  NAND2_X1 U2777 ( .A1(n3171), .A2(REG1_REG_8__SCAN_IN), .ZN(n2237) );
  INV_X1 U2778 ( .A(n3173), .ZN(n2236) );
  NAND2_X1 U2779 ( .A1(n2275), .A2(n2274), .ZN(n4517) );
  NAND2_X1 U2780 ( .A1(n3160), .A2(n2276), .ZN(n2275) );
  XNOR2_X1 U2781 ( .A(n3180), .B(n4553), .ZN(n4550) );
  NOR2_X1 U2782 ( .A1(n4555), .A2(n4045), .ZN(n4566) );
  OR2_X1 U2783 ( .A1(n4043), .A2(n4042), .ZN(n2264) );
  AND2_X1 U2784 ( .A1(n2872), .A2(n3984), .ZN(n4584) );
  NAND2_X1 U2785 ( .A1(n2872), .A2(n2997), .ZN(n4602) );
  AND2_X1 U2786 ( .A1(n2861), .A2(n2865), .ZN(n4594) );
  AND2_X1 U2787 ( .A1(n2238), .A2(n2239), .ZN(n4061) );
  NOR2_X1 U2788 ( .A1(n2240), .A2(n2199), .ZN(n2239) );
  INV_X1 U2789 ( .A(n4584), .ZN(n4588) );
  OAI21_X1 U2790 ( .B1(n4086), .B2(n4327), .A(n4085), .ZN(n2202) );
  NAND2_X1 U2791 ( .A1(n2327), .A2(n2330), .ZN(n2802) );
  NAND2_X1 U2792 ( .A1(n4136), .A2(n2155), .ZN(n2327) );
  INV_X1 U2793 ( .A(n4335), .ZN(n4112) );
  NAND2_X1 U2794 ( .A1(n2331), .A2(n2155), .ZN(n4105) );
  NAND2_X1 U2795 ( .A1(n2331), .A2(n2746), .ZN(n4103) );
  INV_X1 U2796 ( .A(n2690), .ZN(n4134) );
  NAND2_X1 U2797 ( .A1(n2152), .A2(DATAI_21_), .ZN(n4219) );
  NAND2_X1 U2798 ( .A1(n2376), .A2(n2377), .ZN(n4224) );
  OR2_X1 U2799 ( .A1(n4280), .A2(n2154), .ZN(n2376) );
  NAND2_X1 U2800 ( .A1(n4280), .A2(n2650), .ZN(n4249) );
  NAND2_X1 U2801 ( .A1(n2306), .A2(n2307), .ZN(n4292) );
  NAND2_X1 U2802 ( .A1(n4323), .A2(n4322), .ZN(n4321) );
  NAND2_X1 U2803 ( .A1(n3511), .A2(n3834), .ZN(n4323) );
  AND2_X1 U2804 ( .A1(n2282), .A2(n2161), .ZN(n4310) );
  NAND2_X1 U2805 ( .A1(n2282), .A2(n2280), .ZN(n4309) );
  NAND2_X1 U2806 ( .A1(n2381), .A2(n2162), .ZN(n2282) );
  NAND2_X1 U2807 ( .A1(n3456), .A2(n2604), .ZN(n3513) );
  INV_X1 U2808 ( .A(n3484), .ZN(n4433) );
  NAND2_X1 U2809 ( .A1(n2295), .A2(n2293), .ZN(n3281) );
  OR2_X1 U2810 ( .A1(n3243), .A2(n2548), .ZN(n2295) );
  NAND2_X1 U2811 ( .A1(n2317), .A2(n2321), .ZN(n3235) );
  NAND2_X1 U2812 ( .A1(n3209), .A2(n2323), .ZN(n2317) );
  AND2_X1 U2813 ( .A1(n4238), .A2(n4065), .ZN(n4285) );
  INV_X1 U2814 ( .A(n3996), .ZN(n3252) );
  INV_X1 U2815 ( .A(n4327), .ZN(n4296) );
  NAND2_X1 U2816 ( .A1(n2315), .A2(n3924), .ZN(n3150) );
  NAND2_X1 U2817 ( .A1(n2316), .A2(n3921), .ZN(n2315) );
  INV_X1 U2818 ( .A(n2822), .ZN(n2823) );
  INV_X1 U2819 ( .A(n4161), .ZN(n4319) );
  NAND2_X1 U2820 ( .A1(n4285), .A2(n4412), .ZN(n4266) );
  NAND2_X1 U2821 ( .A1(n2970), .A2(n2724), .ZN(n2814) );
  AND2_X1 U2822 ( .A1(n2210), .A2(n3082), .ZN(n3272) );
  INV_X1 U2823 ( .A(n3537), .ZN(n2210) );
  INV_X1 U2824 ( .A(n4627), .ZN(n2857) );
  NAND2_X1 U2825 ( .A1(n2852), .A2(n2851), .ZN(n4942) );
  AND2_X1 U2826 ( .A1(n2423), .A2(n2421), .ZN(n2300) );
  INV_X1 U2827 ( .A(n2997), .ZN(n4497) );
  INV_X1 U2828 ( .A(IR_REG_24__SCAN_IN), .ZN(n2764) );
  XNOR2_X1 U2829 ( .A(n2722), .B(IR_REG_22__SCAN_IN), .ZN(n4500) );
  AND2_X1 U2830 ( .A1(n2721), .A2(n2231), .ZN(n4501) );
  XNOR2_X1 U2831 ( .A(n2649), .B(IR_REG_18__SCAN_IN), .ZN(n4059) );
  AND2_X1 U2832 ( .A1(n2532), .A2(n2525), .ZN(n4504) );
  NAND2_X1 U2833 ( .A1(n2367), .A2(n2366), .ZN(n2365) );
  CLKBUF_X1 U2834 ( .A(IR_REG_0__SCAN_IN), .Z(n4877) );
  INV_X2 U2835 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND2_X1 U2836 ( .A1(n2203), .A2(n2201), .ZN(U3354) );
  NAND2_X1 U2837 ( .A1(n2204), .A2(n4238), .ZN(n2203) );
  INV_X1 U2838 ( .A(n2202), .ZN(n2201) );
  OAI21_X1 U2839 ( .B1(n4083), .B2(n4266), .A(n2205), .ZN(n2204) );
  OR2_X1 U2840 ( .A1(n4083), .A2(n4441), .ZN(n2792) );
  OR2_X1 U2841 ( .A1(n4083), .A2(n4495), .ZN(n2797) );
  OR2_X1 U2842 ( .A1(n4096), .A2(n4495), .ZN(n2810) );
  NAND2_X1 U2843 ( .A1(n3224), .A2(n3200), .ZN(n2153) );
  AND2_X1 U2844 ( .A1(n4275), .A2(n4263), .ZN(n2154) );
  INV_X1 U2845 ( .A(n2145), .ZN(n2685) );
  AND2_X1 U2846 ( .A1(n2746), .A2(n3879), .ZN(n2155) );
  INV_X1 U2847 ( .A(n3993), .ZN(n2294) );
  AND2_X1 U2848 ( .A1(n2361), .A2(n2182), .ZN(n2156) );
  AND2_X1 U2849 ( .A1(n3301), .A2(n3254), .ZN(n2157) );
  AND2_X1 U2850 ( .A1(n2220), .A2(n2184), .ZN(n2158) );
  AND2_X1 U2851 ( .A1(n2177), .A2(n2379), .ZN(n2161) );
  NAND2_X1 U2852 ( .A1(n2175), .A2(n2147), .ZN(n2718) );
  NAND2_X1 U2853 ( .A1(n2367), .A2(IR_REG_1__SCAN_IN), .ZN(n2252) );
  AND2_X1 U2854 ( .A1(n2603), .A2(n2613), .ZN(n2162) );
  AND2_X1 U2855 ( .A1(n2377), .A2(n2190), .ZN(n2163) );
  AND2_X1 U2856 ( .A1(n2307), .A2(n2305), .ZN(n2164) );
  OR2_X1 U2857 ( .A1(n3658), .A2(n3659), .ZN(n2165) );
  NAND2_X1 U2858 ( .A1(n3132), .A2(n3528), .ZN(n3921) );
  AND2_X1 U2859 ( .A1(n2726), .A2(n3918), .ZN(n2725) );
  OR2_X1 U2860 ( .A1(n3992), .A2(n3391), .ZN(n2166) );
  AND3_X1 U2861 ( .A1(n2495), .A2(n2494), .A3(n2493), .ZN(n2167) );
  NAND2_X1 U2862 ( .A1(n2622), .A2(n2161), .ZN(n2281) );
  AND2_X1 U2863 ( .A1(n4877), .A2(REG2_REG_0__SCAN_IN), .ZN(n2168) );
  AND4_X1 U2864 ( .A1(n2232), .A2(n2147), .A3(n2385), .A4(n2160), .ZN(n2169)
         );
  AND2_X1 U2865 ( .A1(n2481), .A2(n2297), .ZN(n2170) );
  OAI21_X1 U2866 ( .B1(n3740), .B2(n2219), .A(n2216), .ZN(n3667) );
  NOR2_X1 U2867 ( .A1(n4598), .A2(n4034), .ZN(n2171) );
  NAND2_X1 U2868 ( .A1(n2169), .A2(n2390), .ZN(n2172) );
  INV_X1 U2869 ( .A(n3879), .ZN(n4102) );
  INV_X1 U2870 ( .A(n2231), .ZN(n2720) );
  NAND2_X1 U2871 ( .A1(n2425), .A2(n2430), .ZN(n2432) );
  INV_X1 U2872 ( .A(n2432), .ZN(n2844) );
  INV_X1 U2873 ( .A(n2324), .ZN(n2323) );
  NAND2_X1 U2874 ( .A1(n2183), .A2(n3937), .ZN(n2324) );
  OR2_X1 U2875 ( .A1(n2905), .A2(n2965), .ZN(n2173) );
  AND2_X1 U2876 ( .A1(n3777), .A2(n3716), .ZN(n2174) );
  OR2_X1 U2877 ( .A1(n4577), .A2(n4033), .ZN(n2243) );
  AND2_X1 U2878 ( .A1(n2387), .A2(n2420), .ZN(n2175) );
  AND2_X1 U2879 ( .A1(n3321), .A2(n3320), .ZN(n2176) );
  NAND2_X1 U2880 ( .A1(n4410), .A2(n3825), .ZN(n2177) );
  INV_X1 U2881 ( .A(IR_REG_13__SCAN_IN), .ZN(n2416) );
  NAND2_X1 U2882 ( .A1(n2293), .A2(n2166), .ZN(n2178) );
  AND2_X1 U2883 ( .A1(n2633), .A2(n2352), .ZN(n2179) );
  NOR2_X1 U2884 ( .A1(n2148), .A2(n3538), .ZN(n2180) );
  AND2_X1 U2885 ( .A1(n2155), .A2(n3853), .ZN(n2181) );
  NOR2_X1 U2886 ( .A1(n3149), .A2(n2314), .ZN(n2313) );
  INV_X1 U2887 ( .A(n2281), .ZN(n2280) );
  AND2_X1 U2888 ( .A1(n3607), .A2(n3604), .ZN(n2182) );
  NAND2_X1 U2889 ( .A1(n3994), .A2(n3344), .ZN(n2183) );
  NAND2_X1 U2890 ( .A1(n3565), .A2(n3566), .ZN(n3731) );
  OR2_X1 U2891 ( .A1(n3742), .A2(n3741), .ZN(n2184) );
  AND2_X1 U2892 ( .A1(n3796), .A2(n2184), .ZN(n2185) );
  NAND2_X1 U2893 ( .A1(n3173), .A2(n4605), .ZN(n2186) );
  NAND2_X1 U2894 ( .A1(n3400), .A2(n2571), .ZN(n3415) );
  AND2_X1 U2895 ( .A1(n3574), .A2(n3573), .ZN(n2187) );
  NAND2_X1 U2896 ( .A1(n3471), .A2(n3470), .ZN(n3547) );
  AND2_X1 U2897 ( .A1(n3556), .A2(n3555), .ZN(n3772) );
  AND2_X1 U2898 ( .A1(n3170), .A2(REG2_REG_9__SCAN_IN), .ZN(n2188) );
  AND2_X1 U2899 ( .A1(n2147), .A2(n2387), .ZN(n2612) );
  AND2_X1 U2900 ( .A1(n4214), .A2(n4230), .ZN(n2189) );
  OR2_X1 U2901 ( .A1(n4214), .A2(n4230), .ZN(n2190) );
  INV_X1 U2902 ( .A(n2149), .ZN(n2492) );
  INV_X1 U2903 ( .A(n2211), .ZN(n4180) );
  NOR2_X1 U2904 ( .A1(n4200), .A2(n2790), .ZN(n2211) );
  NAND2_X1 U2905 ( .A1(n2381), .A2(n2603), .ZN(n3456) );
  AND2_X1 U2906 ( .A1(n2182), .A2(n2226), .ZN(n2191) );
  NOR2_X1 U2907 ( .A1(n3614), .A2(n3613), .ZN(n2192) );
  AND2_X1 U2908 ( .A1(n2634), .A2(n2179), .ZN(n2657) );
  INV_X1 U2909 ( .A(n2358), .ZN(n2357) );
  OAI21_X1 U2910 ( .B1(n3555), .B2(n3774), .A(n3773), .ZN(n2358) );
  AND2_X1 U2911 ( .A1(n2360), .A2(n2359), .ZN(n2193) );
  AND2_X1 U2912 ( .A1(n2340), .A2(n3723), .ZN(n2194) );
  NAND2_X1 U2913 ( .A1(n4162), .A2(n3622), .ZN(n2195) );
  INV_X1 U2914 ( .A(n3837), .ZN(n2308) );
  OAI22_X1 U2915 ( .A1(n3440), .A2(n2593), .B1(n4433), .B2(n3780), .ZN(n3458)
         );
  INV_X1 U2916 ( .A(n3458), .ZN(n2381) );
  INV_X1 U2917 ( .A(n4632), .ZN(n2269) );
  INV_X1 U2918 ( .A(n3764), .ZN(n2363) );
  NAND2_X1 U2919 ( .A1(n2368), .A2(n2475), .ZN(n3524) );
  OR2_X1 U2920 ( .A1(n3339), .A2(n3324), .ZN(n2209) );
  NAND2_X1 U2921 ( .A1(n3130), .A2(n3131), .ZN(n2229) );
  INV_X1 U2922 ( .A(n3887), .ZN(n2305) );
  NAND2_X1 U2923 ( .A1(n2265), .A2(n2268), .ZN(n2196) );
  AND2_X1 U2924 ( .A1(n2275), .A2(n2186), .ZN(n2197) );
  OR2_X1 U2925 ( .A1(n2241), .A2(n4034), .ZN(n2198) );
  NAND2_X1 U2926 ( .A1(n3523), .A2(n2487), .ZN(n3148) );
  AND2_X1 U2927 ( .A1(n4059), .A2(REG1_REG_18__SCAN_IN), .ZN(n2199) );
  AND2_X1 U2928 ( .A1(n2899), .A2(n4507), .ZN(n2200) );
  NAND2_X1 U2929 ( .A1(n2151), .A2(DATAI_26_), .ZN(n4129) );
  INV_X1 U2930 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2255) );
  NAND4_X1 U2931 ( .A1(n2457), .A2(n2455), .A3(n2454), .A4(n2456), .ZN(n3017)
         );
  INV_X1 U2932 ( .A(IR_REG_1__SCAN_IN), .ZN(n2366) );
  INV_X1 U2933 ( .A(IR_REG_0__SCAN_IN), .ZN(n2367) );
  INV_X1 U2934 ( .A(n2209), .ZN(n3340) );
  NAND2_X1 U2935 ( .A1(n3740), .A2(n2216), .ZN(n2215) );
  NAND2_X1 U2936 ( .A1(n2215), .A2(n2213), .ZN(n3593) );
  NAND2_X1 U2937 ( .A1(n2221), .A2(n2360), .ZN(n3556) );
  NAND2_X1 U2938 ( .A1(n2223), .A2(n2224), .ZN(n3620) );
  OAI21_X2 U2939 ( .B1(n3294), .B2(n2349), .A(n2347), .ZN(n3368) );
  NAND4_X1 U2940 ( .A1(n2232), .A2(n2147), .A3(n2385), .A4(n2230), .ZN(n2766)
         );
  NAND4_X1 U2941 ( .A1(n2147), .A2(n2385), .A3(n2160), .A4(n2420), .ZN(n2231)
         );
  NAND2_X1 U2942 ( .A1(n3014), .A2(n2234), .ZN(n2951) );
  OR2_X1 U2943 ( .A1(n3052), .A2(n2950), .ZN(n2234) );
  AND2_X1 U2944 ( .A1(n2243), .A2(n2242), .ZN(n4598) );
  INV_X1 U2945 ( .A(n2243), .ZN(n4597) );
  NAND3_X1 U2946 ( .A1(n2366), .A2(IR_REG_31__SCAN_IN), .A3(n4877), .ZN(n2250)
         );
  AOI22_X1 U2947 ( .A1(n2959), .A2(n2254), .B1(n2899), .B2(n2253), .ZN(n2257)
         );
  INV_X1 U2948 ( .A(n2257), .ZN(n2935) );
  NAND2_X1 U2949 ( .A1(n4510), .A2(REG2_REG_1__SCAN_IN), .ZN(n2258) );
  AND2_X1 U2950 ( .A1(n4509), .A2(REG2_REG_2__SCAN_IN), .ZN(n2260) );
  NOR2_X1 U2951 ( .A1(n4015), .A2(n2261), .ZN(n4012) );
  AOI21_X1 U2952 ( .B1(n4043), .B2(n2267), .A(n2196), .ZN(n2263) );
  NAND2_X1 U2953 ( .A1(n2264), .A2(n2270), .ZN(n4044) );
  OAI21_X1 U2954 ( .B1(n3160), .B2(n2273), .A(n2271), .ZN(n3162) );
  NAND2_X1 U2955 ( .A1(n3458), .A2(n2280), .ZN(n2277) );
  NAND2_X1 U2956 ( .A1(n2277), .A2(n2278), .ZN(n4295) );
  NAND3_X1 U2957 ( .A1(n2284), .A2(n2503), .A3(n2283), .ZN(n3191) );
  NAND4_X1 U2958 ( .A1(n3525), .A2(n2368), .A3(n2502), .A4(n2475), .ZN(n2283)
         );
  NAND3_X1 U2959 ( .A1(n3525), .A2(n2368), .A3(n2475), .ZN(n3523) );
  INV_X1 U2960 ( .A(n2570), .ZN(n3402) );
  AND2_X1 U2961 ( .A1(n2720), .A2(n2298), .ZN(n2426) );
  NAND2_X1 U2962 ( .A1(n2720), .A2(n2299), .ZN(n2425) );
  NAND2_X1 U2963 ( .A1(n3217), .A2(n3874), .ZN(n4651) );
  AOI21_X1 U2964 ( .B1(n4295), .B2(n2640), .A(n2639), .ZN(n4282) );
  NAND2_X1 U2965 ( .A1(n4195), .A2(n4189), .ZN(n4371) );
  AOI22_X1 U2966 ( .A1(n2800), .A2(n2801), .B1(n4092), .B2(n4108), .ZN(n2715)
         );
  INV_X1 U2967 ( .A(n3191), .ZN(n2514) );
  AOI21_X2 U2968 ( .B1(n2514), .B2(n2153), .A(n2157), .ZN(n3217) );
  OAI22_X2 U2969 ( .A1(n4101), .A2(n2699), .B1(n3906), .B2(n4112), .ZN(n2800)
         );
  NAND2_X1 U2970 ( .A1(n3075), .A2(n2474), .ZN(n2368) );
  AOI21_X1 U2971 ( .B1(n4151), .B2(n2689), .A(n2688), .ZN(n2690) );
  NAND2_X1 U2972 ( .A1(n2382), .A2(n2691), .ZN(n4101) );
  XNOR2_X1 U2973 ( .A(n2715), .B(n3904), .ZN(n4076) );
  AOI21_X1 U2974 ( .B1(n2672), .B2(n2394), .A(n2401), .ZN(n4195) );
  NAND2_X1 U2975 ( .A1(n2464), .A2(n3062), .ZN(n3063) );
  NAND2_X2 U2976 ( .A1(n4282), .A2(n4281), .ZN(n4280) );
  NAND2_X1 U2977 ( .A1(n3912), .A2(n3915), .ZN(n2724) );
  INV_X1 U2978 ( .A(n2479), .ZN(n2302) );
  NAND2_X1 U2979 ( .A1(n2429), .A2(n2428), .ZN(n2430) );
  NAND2_X1 U2980 ( .A1(n2370), .A2(n2369), .ZN(n3440) );
  NAND2_X1 U2981 ( .A1(n2150), .A2(REG0_REG_1__SCAN_IN), .ZN(n2457) );
  OR2_X1 U2982 ( .A1(n2145), .A2(n3107), .ZN(n2454) );
  NAND2_X1 U2983 ( .A1(n2313), .A2(n3527), .ZN(n2310) );
  OAI21_X1 U2984 ( .B1(n3209), .B2(n2320), .A(n2318), .ZN(n2731) );
  OAI21_X1 U2985 ( .B1(n3209), .B2(n2730), .A(n3937), .ZN(n3343) );
  AOI21_X1 U2986 ( .B1(n2730), .B2(n3937), .A(n2326), .ZN(n2325) );
  OR2_X1 U2987 ( .A1(n4136), .A2(n3966), .ZN(n2331) );
  AOI21_X1 U2988 ( .B1(n4136), .B2(n2181), .A(n2328), .ZN(n2747) );
  INV_X1 U2989 ( .A(n3724), .ZN(n2332) );
  NAND2_X1 U2990 ( .A1(n2332), .A2(n2194), .ZN(n2335) );
  NAND2_X1 U2991 ( .A1(n2335), .A2(n2336), .ZN(n3683) );
  NAND2_X1 U2992 ( .A1(n2353), .A2(IR_REG_31__SCAN_IN), .ZN(n2635) );
  NAND2_X1 U2993 ( .A1(n3547), .A2(n3546), .ZN(n2359) );
  OAI21_X1 U2994 ( .B1(n3547), .B2(n3546), .A(n3548), .ZN(n2360) );
  NAND3_X1 U2995 ( .A1(n2366), .A2(n2367), .A3(n2408), .ZN(n2473) );
  NAND2_X1 U2996 ( .A1(IR_REG_31__SCAN_IN), .A2(n2365), .ZN(n2448) );
  NAND2_X1 U2997 ( .A1(n3924), .A2(n3921), .ZN(n3525) );
  INV_X1 U2998 ( .A(n2415), .ZN(n2385) );
  NOR2_X1 U2999 ( .A1(n2497), .A2(n2415), .ZN(n2589) );
  INV_X1 U3000 ( .A(n3017), .ZN(n3015) );
  NAND2_X1 U3001 ( .A1(n2437), .A2(n2436), .ZN(n4336) );
  NAND2_X1 U3002 ( .A1(n4475), .A2(n4412), .ZN(n4495) );
  AND2_X1 U3003 ( .A1(n3687), .A2(n3820), .ZN(n2393) );
  NAND2_X1 U3004 ( .A1(n4231), .A2(n4377), .ZN(n2394) );
  AND2_X1 U3005 ( .A1(n4358), .A2(n2790), .ZN(n2395) );
  OR2_X1 U3006 ( .A1(n3230), .A2(n3677), .ZN(n2396) );
  AND2_X1 U3007 ( .A1(n2149), .A2(REG2_REG_4__SCAN_IN), .ZN(n2398) );
  AND2_X1 U3008 ( .A1(n2409), .A2(n2483), .ZN(n2399) );
  NAND2_X1 U3009 ( .A1(n4657), .A2(n4412), .ZN(n4441) );
  OAI22_X1 U3010 ( .A1(n3301), .A2(n3042), .B1(n3674), .B2(n3254), .ZN(n3291)
         );
  NAND2_X1 U3011 ( .A1(n3063), .A2(n2465), .ZN(n3075) );
  INV_X1 U3012 ( .A(n3619), .ZN(n3616) );
  AND2_X1 U3013 ( .A1(n3955), .A2(n3837), .ZN(n4322) );
  AND2_X1 U3014 ( .A1(n3788), .A2(n4219), .ZN(n2401) );
  OR2_X1 U3015 ( .A1(n4175), .A2(n4198), .ZN(n2402) );
  INV_X1 U3016 ( .A(n4625), .ZN(n4238) );
  NOR2_X1 U3017 ( .A1(n4177), .A2(n4356), .ZN(n2688) );
  INV_X1 U3018 ( .A(n3468), .ZN(n3469) );
  INV_X1 U3019 ( .A(n3711), .ZN(n3555) );
  AND2_X1 U3020 ( .A1(n2946), .A2(n4877), .ZN(n2947) );
  OR4_X1 U3021 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_29__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2780) );
  NAND2_X1 U3022 ( .A1(n3529), .A2(n3016), .ZN(n3045) );
  AND2_X1 U3023 ( .A1(n4338), .A2(n4092), .ZN(n3849) );
  INV_X1 U3024 ( .A(IR_REG_18__SCAN_IN), .ZN(n4878) );
  INV_X1 U3025 ( .A(n3292), .ZN(n3295) );
  INV_X1 U3026 ( .A(n3126), .ZN(n3127) );
  NOR2_X1 U3027 ( .A1(n2192), .A2(n3616), .ZN(n3617) );
  INV_X1 U3028 ( .A(n3787), .ZN(n3607) );
  NAND2_X1 U3029 ( .A1(n3726), .A2(n4129), .ZN(n2691) );
  INV_X1 U3030 ( .A(n4304), .ZN(n4398) );
  INV_X1 U3031 ( .A(IR_REG_11__SCAN_IN), .ZN(n2566) );
  INV_X1 U3032 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3705) );
  INV_X1 U3033 ( .A(n4430), .ZN(n4410) );
  INV_X1 U3034 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3755) );
  OR2_X1 U3035 ( .A1(n4090), .A2(n2148), .ZN(n2708) );
  AOI21_X1 U3036 ( .B1(n3998), .B2(n3016), .A(n2951), .ZN(n2952) );
  AND2_X1 U3037 ( .A1(n2151), .A2(n2860), .ZN(n2866) );
  AND3_X1 U3038 ( .A1(n2885), .A2(n2884), .A3(n2883), .ZN(n4072) );
  INV_X1 U3039 ( .A(n2801), .ZN(n2799) );
  AND2_X1 U3040 ( .A1(n3889), .A2(n3888), .ZN(n4255) );
  INV_X1 U3041 ( .A(n4322), .ZN(n2622) );
  INV_X1 U3042 ( .A(n4065), .ZN(n3539) );
  OR2_X1 U3043 ( .A1(n3446), .A2(n4501), .ZN(n2822) );
  INV_X1 U3044 ( .A(n4181), .ZN(n2790) );
  INV_X1 U3045 ( .A(n4274), .ZN(n4284) );
  INV_X1 U3046 ( .A(n2592), .ZN(n3780) );
  INV_X1 U3047 ( .A(n3369), .ZN(n3376) );
  AND2_X1 U3048 ( .A1(n3862), .A2(n2748), .ZN(n4261) );
  NAND2_X1 U3049 ( .A1(n4497), .A2(n2979), .ZN(n4432) );
  INV_X1 U3050 ( .A(n4498), .ZN(n2787) );
  NOR2_X1 U3051 ( .A1(n2840), .A2(n2853), .ZN(n2774) );
  AND2_X1 U3052 ( .A1(n3688), .A2(n2393), .ZN(n3686) );
  NOR2_X1 U3053 ( .A1(n2666), .A2(n3705), .ZN(n2673) );
  AOI22_X1 U3054 ( .A1(n3089), .A2(n3088), .B1(n3087), .B2(n3086), .ZN(n3094)
         );
  OR2_X1 U3055 ( .A1(n2660), .A2(n3767), .ZN(n2666) );
  NOR2_X1 U3056 ( .A1(n2642), .A2(n4862), .ZN(n2651) );
  AND2_X1 U3057 ( .A1(n2692), .A2(n2407), .ZN(n4126) );
  XNOR2_X1 U3058 ( .A(n2776), .B(n2775), .ZN(n3051) );
  OAI211_X1 U3059 ( .C1(n2492), .C2(n4158), .A(n2687), .B(n2686), .ZN(n4177)
         );
  AND2_X1 U3060 ( .A1(n2866), .A2(n2865), .ZN(n2872) );
  AND2_X1 U3061 ( .A1(n2872), .A2(n2954), .ZN(n4595) );
  INV_X1 U3062 ( .A(n4079), .ZN(n4314) );
  INV_X1 U3063 ( .A(n4261), .ZN(n4437) );
  AND2_X1 U3064 ( .A1(n3926), .A2(n3938), .ZN(n3875) );
  INV_X1 U3065 ( .A(n4266), .ZN(n4611) );
  NAND2_X1 U3066 ( .A1(n2823), .A2(n2851), .ZN(n4603) );
  NAND2_X1 U3067 ( .A1(n2788), .A2(n2856), .ZN(n2820) );
  AOI21_X1 U3068 ( .B1(n4087), .B2(n4423), .A(n2805), .ZN(n3543) );
  INV_X1 U3069 ( .A(n3403), .ZN(n3477) );
  INV_X1 U3070 ( .A(n2989), .ZN(n2851) );
  INV_X1 U3071 ( .A(n2850), .ZN(n2852) );
  AND2_X1 U3072 ( .A1(n2580), .A2(n2568), .ZN(n3169) );
  NAND2_X1 U3073 ( .A1(n3051), .A2(STATE_REG_SCAN_IN), .ZN(n4627) );
  NAND2_X1 U3074 ( .A1(n2991), .A2(n2988), .ZN(n3815) );
  INV_X1 U3075 ( .A(n4338), .ZN(n4108) );
  OAI211_X1 U3076 ( .C1(n4183), .C2(n2148), .A(n2680), .B(n2679), .ZN(n4358)
         );
  INV_X1 U3077 ( .A(n4594), .ZN(n4587) );
  NAND2_X1 U3078 ( .A1(n4606), .A2(n3111), .ZN(n4327) );
  OR2_X1 U3079 ( .A1(n2794), .A2(n2820), .ZN(n4655) );
  OR2_X1 U3080 ( .A1(n3459), .A2(n3442), .ZN(n3509) );
  OR2_X1 U3081 ( .A1(n3282), .A2(n3237), .ZN(n3319) );
  INV_X1 U3082 ( .A(n4475), .ZN(n4653) );
  INV_X1 U3083 ( .A(n4942), .ZN(n4626) );
  INV_X1 U3084 ( .A(D_REG_0__SCAN_IN), .ZN(n2859) );
  INV_X1 U3085 ( .A(n3169), .ZN(n4637) );
  NOR2_X1 U3086 ( .A1(n3052), .A2(n4627), .ZN(U4043) );
  INV_X1 U3087 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2789) );
  NAND2_X1 U3088 ( .A1(n2516), .A2(REG3_REG_7__SCAN_IN), .ZN(n2539) );
  NAND2_X1 U3089 ( .A1(REG3_REG_8__SCAN_IN), .A2(REG3_REG_9__SCAN_IN), .ZN(
        n2403) );
  NOR2_X1 U3090 ( .A1(n2539), .A2(n2403), .ZN(n2550) );
  NAND2_X1 U3091 ( .A1(n2550), .A2(REG3_REG_10__SCAN_IN), .ZN(n2574) );
  NAND2_X1 U3092 ( .A1(REG3_REG_12__SCAN_IN), .A2(REG3_REG_11__SCAN_IN), .ZN(
        n2404) );
  NAND2_X1 U3093 ( .A1(n2605), .A2(REG3_REG_15__SCAN_IN), .ZN(n2626) );
  NAND2_X1 U3094 ( .A1(REG3_REG_16__SCAN_IN), .A2(REG3_REG_17__SCAN_IN), .ZN(
        n2405) );
  NAND2_X1 U3095 ( .A1(n2651), .A2(REG3_REG_19__SCAN_IN), .ZN(n2660) );
  NAND2_X1 U3096 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2406) );
  INV_X1 U3097 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4680) );
  INV_X1 U3098 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3809) );
  OAI21_X1 U3099 ( .B1(n2684), .B2(n4680), .A(n3809), .ZN(n2407) );
  INV_X1 U3100 ( .A(n2473), .ZN(n2410) );
  NOR2_X1 U3101 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2414)
         );
  INV_X1 U3102 ( .A(IR_REG_22__SCAN_IN), .ZN(n2421) );
  NAND2_X1 U3103 ( .A1(n2427), .A2(IR_REG_29__SCAN_IN), .ZN(n2429) );
  NAND2_X1 U3104 ( .A1(n4126), .A2(n2302), .ZN(n2437) );
  INV_X1 U3105 ( .A(n2848), .ZN(n2431) );
  INV_X1 U3106 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4350) );
  AND2_X2 U3107 ( .A1(n2848), .A2(n2432), .ZN(n2469) );
  NAND2_X1 U3108 ( .A1(n2149), .A2(REG2_REG_26__SCAN_IN), .ZN(n2434) );
  NAND2_X1 U3109 ( .A1(n2458), .A2(REG0_REG_26__SCAN_IN), .ZN(n2433) );
  OAI211_X1 U3110 ( .C1(n2145), .C2(n4350), .A(n2434), .B(n2433), .ZN(n2435)
         );
  INV_X1 U3111 ( .A(n2435), .ZN(n2436) );
  INV_X1 U3112 ( .A(n4336), .ZN(n3726) );
  NAND2_X2 U3113 ( .A1(n2440), .A2(n2439), .ZN(n2463) );
  INV_X1 U3114 ( .A(n4145), .ZN(n3622) );
  XNOR2_X1 U3115 ( .A(n2684), .B(REG3_REG_25__SCAN_IN), .ZN(n4146) );
  NAND2_X1 U3116 ( .A1(n4146), .A2(n2302), .ZN(n2445) );
  INV_X1 U3117 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4354) );
  NAND2_X1 U3118 ( .A1(n2150), .A2(REG0_REG_25__SCAN_IN), .ZN(n2442) );
  NAND2_X1 U3119 ( .A1(n2149), .A2(REG2_REG_25__SCAN_IN), .ZN(n2441) );
  OAI211_X1 U3120 ( .C1(n2145), .C2(n4354), .A(n2442), .B(n2441), .ZN(n2443)
         );
  INV_X1 U3121 ( .A(n2443), .ZN(n2444) );
  INV_X1 U3122 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2446) );
  OR2_X1 U3123 ( .A1(n2447), .A2(n2446), .ZN(n2451) );
  INV_X1 U3124 ( .A(REG1_REG_2__SCAN_IN), .ZN(n4885) );
  OR2_X2 U3125 ( .A1(n2145), .A2(n4885), .ZN(n2452) );
  NAND2_X1 U3126 ( .A1(n2149), .A2(REG2_REG_2__SCAN_IN), .ZN(n2450) );
  MUX2_X1 U3127 ( .A(n4509), .B(DATAI_2_), .S(n2463), .Z(n3066) );
  NAND2_X1 U3128 ( .A1(n3029), .A2(n3066), .ZN(n2726) );
  NAND4_X1 U3129 ( .A1(n2452), .A2(n2451), .A3(n2450), .A4(n2449), .ZN(n2828)
         );
  NAND2_X1 U3130 ( .A1(n2828), .A2(n3140), .ZN(n3918) );
  INV_X1 U3131 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3025) );
  INV_X1 U3132 ( .A(REG1_REG_1__SCAN_IN), .ZN(n3107) );
  NAND2_X1 U3133 ( .A1(n2149), .A2(REG2_REG_1__SCAN_IN), .ZN(n2456) );
  MUX2_X1 U3134 ( .A(n4510), .B(DATAI_1_), .S(n2463), .Z(n3101) );
  NAND2_X1 U3135 ( .A1(n3017), .A2(n3101), .ZN(n3061) );
  INV_X1 U3136 ( .A(n3061), .ZN(n2453) );
  NAND2_X1 U3137 ( .A1(n3017), .A2(n3023), .ZN(n3912) );
  INV_X1 U3138 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2950) );
  OR2_X1 U3139 ( .A1(n2145), .A2(n2950), .ZN(n2462) );
  NAND2_X1 U3140 ( .A1(n2458), .A2(REG0_REG_0__SCAN_IN), .ZN(n2461) );
  INV_X1 U3141 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3000) );
  NAND2_X1 U3142 ( .A1(n2149), .A2(REG2_REG_0__SCAN_IN), .ZN(n2459) );
  MUX2_X1 U3143 ( .A(n4877), .B(DATAI_0_), .S(n2463), .Z(n2993) );
  AND2_X1 U3144 ( .A1(n3998), .A2(n2993), .ZN(n2812) );
  NAND2_X1 U3145 ( .A1(n2724), .A2(n2812), .ZN(n3062) );
  NAND2_X1 U3146 ( .A1(n3029), .A2(n3140), .ZN(n2465) );
  OR2_X1 U3147 ( .A1(n2148), .A2(REG3_REG_3__SCAN_IN), .ZN(n2466) );
  INV_X1 U31480 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2467) );
  OR2_X1 U31490 ( .A1(n2145), .A2(n2467), .ZN(n2472) );
  NAND2_X1 U3150 ( .A1(n2458), .A2(REG0_REG_3__SCAN_IN), .ZN(n2471) );
  NAND2_X1 U3151 ( .A1(n2149), .A2(REG2_REG_3__SCAN_IN), .ZN(n2470) );
  NAND2_X1 U3152 ( .A1(n2473), .A2(IR_REG_31__SCAN_IN), .ZN(n2484) );
  XNOR2_X1 U3153 ( .A(n2484), .B(IR_REG_3__SCAN_IN), .ZN(n4508) );
  MUX2_X1 U3154 ( .A(n4508), .B(DATAI_3_), .S(n2463), .Z(n3043) );
  NAND2_X1 U3155 ( .A1(n3529), .A2(n3043), .ZN(n2474) );
  NAND2_X1 U3156 ( .A1(n3141), .A2(n3117), .ZN(n2475) );
  INV_X1 U3157 ( .A(n2476), .ZN(n2490) );
  INV_X1 U3158 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2477) );
  INV_X1 U3159 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4894) );
  NAND2_X1 U3160 ( .A1(n2477), .A2(n4894), .ZN(n2478) );
  NAND2_X1 U3161 ( .A1(n2490), .A2(n2478), .ZN(n3538) );
  NOR2_X1 U3162 ( .A1(n2398), .A2(n2180), .ZN(n2482) );
  INV_X1 U3163 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2480) );
  NAND2_X1 U3164 ( .A1(n2458), .A2(REG0_REG_4__SCAN_IN), .ZN(n2481) );
  NAND2_X1 U3165 ( .A1(n2484), .A2(n2483), .ZN(n2485) );
  NAND2_X1 U3166 ( .A1(n2485), .A2(IR_REG_31__SCAN_IN), .ZN(n2486) );
  XNOR2_X1 U3167 ( .A(n2486), .B(IR_REG_4__SCAN_IN), .ZN(n4507) );
  MUX2_X1 U3168 ( .A(n4507), .B(DATAI_4_), .S(n2152), .Z(n3528) );
  INV_X1 U3169 ( .A(n3528), .ZN(n3536) );
  NAND2_X1 U3170 ( .A1(n3225), .A2(n3528), .ZN(n2487) );
  NAND2_X1 U3171 ( .A1(n2458), .A2(REG0_REG_5__SCAN_IN), .ZN(n2496) );
  INV_X1 U3172 ( .A(n2488), .ZN(n2506) );
  INV_X1 U3173 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2489) );
  NAND2_X1 U3174 ( .A1(n2490), .A2(n2489), .ZN(n2491) );
  NAND2_X1 U3175 ( .A1(n2506), .A2(n2491), .ZN(n3226) );
  OR2_X1 U3176 ( .A1(n2148), .A2(n3226), .ZN(n2495) );
  INV_X1 U3177 ( .A(REG1_REG_5__SCAN_IN), .ZN(n3158) );
  OR2_X1 U3178 ( .A1(n2145), .A2(n3158), .ZN(n2494) );
  NAND2_X1 U3179 ( .A1(n2149), .A2(REG2_REG_5__SCAN_IN), .ZN(n2493) );
  NAND2_X1 U3180 ( .A1(n2498), .A2(IR_REG_31__SCAN_IN), .ZN(n2499) );
  MUX2_X1 U3181 ( .A(IR_REG_31__SCAN_IN), .B(n2499), .S(IR_REG_5__SCAN_IN), 
        .Z(n2501) );
  NOR2_X1 U3182 ( .A1(n2498), .A2(IR_REG_5__SCAN_IN), .ZN(n2522) );
  INV_X1 U3183 ( .A(n2522), .ZN(n2500) );
  NAND2_X1 U3184 ( .A1(n2501), .A2(n2500), .ZN(n2906) );
  INV_X1 U3185 ( .A(DATAI_5_), .ZN(n4869) );
  MUX2_X1 U3186 ( .A(n2906), .B(n4869), .S(n2151), .Z(n3230) );
  NAND2_X1 U3187 ( .A1(n3252), .A2(n3230), .ZN(n2502) );
  NAND2_X1 U3188 ( .A1(n3996), .A2(n3154), .ZN(n2503) );
  NAND2_X1 U3189 ( .A1(n2149), .A2(REG2_REG_6__SCAN_IN), .ZN(n2512) );
  NAND2_X1 U3190 ( .A1(n2458), .A2(REG0_REG_6__SCAN_IN), .ZN(n2511) );
  INV_X1 U3191 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2504) );
  OR2_X1 U3192 ( .A1(n2145), .A2(n2504), .ZN(n2510) );
  INV_X1 U3193 ( .A(n2516), .ZN(n2508) );
  INV_X1 U3194 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2505) );
  NAND2_X1 U3195 ( .A1(n2506), .A2(n2505), .ZN(n2507) );
  NAND2_X1 U3196 ( .A1(n2508), .A2(n2507), .ZN(n3259) );
  OR2_X1 U3197 ( .A1(n2148), .A2(n3259), .ZN(n2509) );
  NAND4_X1 U3198 ( .A1(n2512), .A2(n2511), .A3(n2510), .A4(n2509), .ZN(n3224)
         );
  OR2_X1 U3199 ( .A1(n2522), .A2(n2846), .ZN(n2513) );
  XNOR2_X1 U3200 ( .A(n2513), .B(IR_REG_6__SCAN_IN), .ZN(n4505) );
  MUX2_X1 U3201 ( .A(n4505), .B(DATAI_6_), .S(n2152), .Z(n3200) );
  NAND2_X1 U3202 ( .A1(n2149), .A2(REG2_REG_7__SCAN_IN), .ZN(n2520) );
  NAND2_X1 U3203 ( .A1(n2458), .A2(REG0_REG_7__SCAN_IN), .ZN(n2519) );
  INV_X1 U3204 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2515) );
  OR2_X1 U3205 ( .A1(n2145), .A2(n2515), .ZN(n2518) );
  OAI21_X1 U3206 ( .B1(n2516), .B2(REG3_REG_7__SCAN_IN), .A(n2539), .ZN(n3308)
         );
  OR2_X1 U3207 ( .A1(n2148), .A2(n3308), .ZN(n2517) );
  NAND4_X1 U3208 ( .A1(n2520), .A2(n2519), .A3(n2518), .A4(n2517), .ZN(n3995)
         );
  NAND2_X1 U3209 ( .A1(n2522), .A2(n2521), .ZN(n2546) );
  NAND2_X1 U32100 ( .A1(n2546), .A2(IR_REG_31__SCAN_IN), .ZN(n2524) );
  INV_X1 U32110 ( .A(IR_REG_7__SCAN_IN), .ZN(n2523) );
  NAND2_X1 U32120 ( .A1(n2524), .A2(n2523), .ZN(n2532) );
  OR2_X1 U32130 ( .A1(n2524), .A2(n2523), .ZN(n2525) );
  MUX2_X1 U32140 ( .A(n4504), .B(DATAI_7_), .S(n2151), .Z(n3296) );
  NAND2_X1 U32150 ( .A1(n3345), .A2(n3296), .ZN(n2729) );
  INV_X1 U32160 ( .A(n3296), .ZN(n3303) );
  NAND2_X1 U32170 ( .A1(n3995), .A2(n3303), .ZN(n3937) );
  NAND2_X1 U32180 ( .A1(n2729), .A2(n3937), .ZN(n3874) );
  NAND2_X1 U32190 ( .A1(n3995), .A2(n3296), .ZN(n2526) );
  NAND2_X1 U32200 ( .A1(n4651), .A2(n2526), .ZN(n3342) );
  NAND2_X1 U32210 ( .A1(n2149), .A2(REG2_REG_8__SCAN_IN), .ZN(n2531) );
  NAND2_X1 U32220 ( .A1(n2458), .A2(REG0_REG_8__SCAN_IN), .ZN(n2530) );
  INV_X1 U32230 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3174) );
  OR2_X1 U32240 ( .A1(n2145), .A2(n3174), .ZN(n2529) );
  INV_X1 U32250 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2527) );
  XNOR2_X1 U32260 ( .A(n2539), .B(n2527), .ZN(n4604) );
  OR2_X1 U32270 ( .A1(n2148), .A2(n4604), .ZN(n2528) );
  NAND4_X1 U32280 ( .A1(n2531), .A2(n2530), .A3(n2529), .A4(n2528), .ZN(n3994)
         );
  INV_X1 U32290 ( .A(n3994), .ZN(n3374) );
  NAND2_X1 U32300 ( .A1(n2532), .A2(IR_REG_31__SCAN_IN), .ZN(n2534) );
  INV_X1 U32310 ( .A(IR_REG_8__SCAN_IN), .ZN(n2533) );
  XNOR2_X1 U32320 ( .A(n2534), .B(n2533), .ZN(n3173) );
  INV_X1 U32330 ( .A(DATAI_8_), .ZN(n2834) );
  MUX2_X1 U32340 ( .A(n3173), .B(n2834), .S(n2152), .Z(n3344) );
  NAND2_X1 U32350 ( .A1(n3374), .A2(n3344), .ZN(n2535) );
  NAND2_X1 U32360 ( .A1(n3342), .A2(n2535), .ZN(n2537) );
  NAND2_X1 U32370 ( .A1(n3994), .A2(n3324), .ZN(n2536) );
  NAND2_X1 U32380 ( .A1(n2537), .A2(n2536), .ZN(n3243) );
  NAND2_X1 U32390 ( .A1(n2150), .A2(REG0_REG_9__SCAN_IN), .ZN(n2545) );
  NAND2_X1 U32400 ( .A1(n2149), .A2(REG2_REG_9__SCAN_IN), .ZN(n2544) );
  INV_X1 U32410 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2538) );
  OR2_X1 U32420 ( .A1(n2145), .A2(n2538), .ZN(n2543) );
  INV_X1 U32430 ( .A(n2539), .ZN(n2540) );
  AOI21_X1 U32440 ( .B1(n2540), .B2(REG3_REG_8__SCAN_IN), .A(
        REG3_REG_9__SCAN_IN), .ZN(n2541) );
  OR2_X1 U32450 ( .A1(n2541), .A2(n2550), .ZN(n3381) );
  OR2_X1 U32460 ( .A1(n2148), .A2(n3381), .ZN(n2542) );
  NAND4_X1 U32470 ( .A1(n2545), .A2(n2544), .A3(n2543), .A4(n2542), .ZN(n3993)
         );
  NAND2_X1 U32480 ( .A1(n2556), .A2(IR_REG_31__SCAN_IN), .ZN(n2547) );
  XNOR2_X1 U32490 ( .A(n2547), .B(IR_REG_9__SCAN_IN), .ZN(n3170) );
  MUX2_X1 U32500 ( .A(n3170), .B(DATAI_9_), .S(n2151), .Z(n3369) );
  AND2_X1 U32510 ( .A1(n3993), .A2(n3369), .ZN(n2548) );
  NAND2_X1 U32520 ( .A1(n2149), .A2(REG2_REG_10__SCAN_IN), .ZN(n2555) );
  NAND2_X1 U32530 ( .A1(n2458), .A2(REG0_REG_10__SCAN_IN), .ZN(n2554) );
  INV_X1 U32540 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2549) );
  OR2_X1 U32550 ( .A1(n2145), .A2(n2549), .ZN(n2553) );
  OR2_X1 U32560 ( .A1(n2550), .A2(REG3_REG_10__SCAN_IN), .ZN(n2551) );
  NAND2_X1 U32570 ( .A1(n2574), .A2(n2551), .ZN(n3399) );
  OR2_X1 U32580 ( .A1(n2148), .A2(n3399), .ZN(n2552) );
  NAND4_X1 U32590 ( .A1(n2555), .A2(n2554), .A3(n2553), .A4(n2552), .ZN(n3992)
         );
  NOR2_X1 U32600 ( .A1(n2556), .A2(IR_REG_9__SCAN_IN), .ZN(n2564) );
  OR2_X1 U32610 ( .A1(n2564), .A2(n2846), .ZN(n2557) );
  XNOR2_X1 U32620 ( .A(n2557), .B(IR_REG_10__SCAN_IN), .ZN(n3176) );
  MUX2_X1 U32630 ( .A(n3176), .B(DATAI_10_), .S(n2152), .Z(n3391) );
  NAND2_X1 U32640 ( .A1(n3992), .A2(n3391), .ZN(n2558) );
  NAND2_X1 U32650 ( .A1(n2149), .A2(REG2_REG_11__SCAN_IN), .ZN(n2562) );
  NAND2_X1 U32660 ( .A1(n2150), .A2(REG0_REG_11__SCAN_IN), .ZN(n2561) );
  INV_X1 U32670 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3450) );
  OR2_X1 U32680 ( .A1(n2145), .A2(n3450), .ZN(n2560) );
  INV_X1 U32690 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2573) );
  XNOR2_X1 U32700 ( .A(n2574), .B(n2573), .ZN(n3482) );
  OR2_X1 U32710 ( .A1(n2148), .A2(n3482), .ZN(n2559) );
  NAND4_X1 U32720 ( .A1(n2562), .A2(n2561), .A3(n2560), .A4(n2559), .ZN(n3483)
         );
  INV_X1 U32730 ( .A(IR_REG_10__SCAN_IN), .ZN(n2563) );
  NAND2_X1 U32740 ( .A1(n2564), .A2(n2563), .ZN(n2565) );
  NAND2_X1 U32750 ( .A1(n2565), .A2(IR_REG_31__SCAN_IN), .ZN(n2567) );
  NAND2_X1 U32760 ( .A1(n2567), .A2(n2566), .ZN(n2580) );
  OR2_X1 U32770 ( .A1(n2567), .A2(n2566), .ZN(n2568) );
  MUX2_X1 U32780 ( .A(n3169), .B(DATAI_11_), .S(n2151), .Z(n3403) );
  NAND2_X1 U32790 ( .A1(n3715), .A2(n3403), .ZN(n3911) );
  NAND2_X1 U32800 ( .A1(n3483), .A2(n3477), .ZN(n3947) );
  NAND2_X1 U32810 ( .A1(n3715), .A2(n3477), .ZN(n2571) );
  NAND2_X1 U32820 ( .A1(n2149), .A2(REG2_REG_12__SCAN_IN), .ZN(n2579) );
  NAND2_X1 U32830 ( .A1(n2150), .A2(REG0_REG_12__SCAN_IN), .ZN(n2578) );
  INV_X1 U32840 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4762) );
  OR2_X1 U32850 ( .A1(n2145), .A2(n4762), .ZN(n2577) );
  INV_X1 U32860 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2572) );
  OAI21_X1 U32870 ( .B1(n2574), .B2(n2573), .A(n2572), .ZN(n2575) );
  NAND2_X1 U32880 ( .A1(n2575), .A2(n2583), .ZN(n3721) );
  OR2_X1 U32890 ( .A1(n2148), .A2(n3721), .ZN(n2576) );
  NAND4_X1 U32900 ( .A1(n2579), .A2(n2578), .A3(n2577), .A4(n2576), .ZN(n3991)
         );
  NAND2_X1 U32910 ( .A1(n2580), .A2(IR_REG_31__SCAN_IN), .ZN(n2581) );
  XNOR2_X1 U32920 ( .A(n2581), .B(IR_REG_12__SCAN_IN), .ZN(n4634) );
  MUX2_X1 U32930 ( .A(n4634), .B(DATAI_12_), .S(n2151), .Z(n3552) );
  INV_X1 U32940 ( .A(n3991), .ZN(n3777) );
  INV_X1 U32950 ( .A(n3552), .ZN(n3716) );
  NAND2_X1 U32960 ( .A1(n2150), .A2(REG0_REG_13__SCAN_IN), .ZN(n2588) );
  NAND2_X1 U32970 ( .A1(n2149), .A2(REG2_REG_13__SCAN_IN), .ZN(n2587) );
  INV_X1 U32980 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3182) );
  OR2_X1 U32990 ( .A1(n2145), .A2(n3182), .ZN(n2586) );
  NAND2_X1 U33000 ( .A1(n2583), .A2(n3185), .ZN(n2584) );
  NAND2_X1 U33010 ( .A1(n2595), .A2(n2584), .ZN(n3785) );
  OR2_X1 U33020 ( .A1(n2148), .A2(n3785), .ZN(n2585) );
  NAND4_X1 U33030 ( .A1(n2588), .A2(n2587), .A3(n2586), .A4(n2585), .ZN(n3484)
         );
  NOR2_X1 U33040 ( .A1(n2589), .A2(n2846), .ZN(n2590) );
  MUX2_X1 U33050 ( .A(n2846), .B(n2590), .S(IR_REG_13__SCAN_IN), .Z(n2591) );
  OR2_X1 U33060 ( .A1(n2591), .A2(n2612), .ZN(n3188) );
  INV_X1 U33070 ( .A(n3188), .ZN(n4503) );
  MUX2_X1 U33080 ( .A(n4503), .B(DATAI_13_), .S(n2151), .Z(n2592) );
  NOR2_X1 U33090 ( .A1(n3484), .A2(n2592), .ZN(n2593) );
  NAND2_X1 U33100 ( .A1(n2149), .A2(REG2_REG_14__SCAN_IN), .ZN(n2601) );
  NAND2_X1 U33110 ( .A1(n2458), .A2(REG0_REG_14__SCAN_IN), .ZN(n2600) );
  INV_X1 U33120 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4439) );
  OR2_X1 U33130 ( .A1(n2145), .A2(n4439), .ZN(n2599) );
  INV_X1 U33140 ( .A(n2605), .ZN(n2597) );
  NAND2_X1 U33150 ( .A1(n2595), .A2(n2594), .ZN(n2596) );
  NAND2_X1 U33160 ( .A1(n2597), .A2(n2596), .ZN(n3657) );
  OR2_X1 U33170 ( .A1(n2148), .A2(n3657), .ZN(n2598) );
  NAND4_X1 U33180 ( .A1(n2601), .A2(n2600), .A3(n2599), .A4(n2598), .ZN(n3990)
         );
  OR2_X1 U33190 ( .A1(n2612), .A2(n2846), .ZN(n2602) );
  XNOR2_X1 U33200 ( .A(n2602), .B(IR_REG_14__SCAN_IN), .ZN(n4632) );
  MUX2_X1 U33210 ( .A(n4632), .B(DATAI_14_), .S(n2152), .Z(n4428) );
  NAND2_X1 U33220 ( .A1(n4421), .A2(n4428), .ZN(n3832) );
  NAND2_X1 U33230 ( .A1(n3990), .A2(n3652), .ZN(n3833) );
  NAND2_X1 U33240 ( .A1(n4421), .A2(n3652), .ZN(n2604) );
  NAND2_X1 U33250 ( .A1(n2149), .A2(REG2_REG_15__SCAN_IN), .ZN(n2610) );
  NAND2_X1 U33260 ( .A1(n2458), .A2(REG0_REG_15__SCAN_IN), .ZN(n2609) );
  INV_X1 U33270 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4425) );
  OR2_X1 U33280 ( .A1(n2145), .A2(n4425), .ZN(n2608) );
  OR2_X1 U33290 ( .A1(n2605), .A2(REG3_REG_15__SCAN_IN), .ZN(n2606) );
  NAND2_X1 U33300 ( .A1(n2626), .A2(n2606), .ZN(n3830) );
  OR2_X1 U33310 ( .A1(n2148), .A2(n3830), .ZN(n2607) );
  NAND4_X1 U33320 ( .A1(n2610), .A2(n2609), .A3(n2608), .A4(n2607), .ZN(n4430)
         );
  NAND2_X1 U33330 ( .A1(n2612), .A2(n2611), .ZN(n2632) );
  NAND2_X1 U33340 ( .A1(n2632), .A2(IR_REG_31__SCAN_IN), .ZN(n2619) );
  XNOR2_X1 U33350 ( .A(n2619), .B(IR_REG_15__SCAN_IN), .ZN(n4047) );
  MUX2_X1 U33360 ( .A(n4047), .B(DATAI_15_), .S(n2152), .Z(n4417) );
  NAND2_X1 U33370 ( .A1(n4430), .A2(n4417), .ZN(n2613) );
  NAND2_X1 U33380 ( .A1(n2149), .A2(REG2_REG_16__SCAN_IN), .ZN(n2617) );
  NAND2_X1 U33390 ( .A1(n2458), .A2(REG0_REG_16__SCAN_IN), .ZN(n2616) );
  INV_X1 U33400 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4774) );
  OR2_X1 U33410 ( .A1(n2145), .A2(n4774), .ZN(n2615) );
  INV_X1 U33420 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2625) );
  XNOR2_X1 U33430 ( .A(n2626), .B(n2625), .ZN(n4315) );
  OR2_X1 U33440 ( .A1(n2148), .A2(n4315), .ZN(n2614) );
  NAND4_X1 U33450 ( .A1(n2617), .A2(n2616), .A3(n2615), .A4(n2614), .ZN(n4418)
         );
  INV_X1 U33460 ( .A(n4418), .ZN(n4402) );
  INV_X1 U33470 ( .A(IR_REG_15__SCAN_IN), .ZN(n2618) );
  NAND2_X1 U33480 ( .A1(n2619), .A2(n2618), .ZN(n2620) );
  NAND2_X1 U33490 ( .A1(n2620), .A2(IR_REG_31__SCAN_IN), .ZN(n2621) );
  XNOR2_X1 U33500 ( .A(n2621), .B(IR_REG_16__SCAN_IN), .ZN(n4049) );
  MUX2_X1 U33510 ( .A(n4049), .B(DATAI_16_), .S(n2152), .Z(n4407) );
  NAND2_X1 U33520 ( .A1(n4402), .A2(n4407), .ZN(n3955) );
  INV_X1 U3353 ( .A(n4407), .ZN(n4320) );
  NAND2_X1 U33540 ( .A1(n4418), .A2(n4320), .ZN(n3837) );
  NAND2_X1 U3355 ( .A1(n4418), .A2(n4407), .ZN(n2623) );
  NAND2_X1 U3356 ( .A1(n2149), .A2(REG2_REG_17__SCAN_IN), .ZN(n2631) );
  NAND2_X1 U3357 ( .A1(n2150), .A2(REG0_REG_17__SCAN_IN), .ZN(n2630) );
  INV_X1 U3358 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4405) );
  OR2_X1 U3359 ( .A1(n2145), .A2(n4405), .ZN(n2629) );
  INV_X1 U3360 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2624) );
  OAI21_X1 U3361 ( .B1(n2626), .B2(n2625), .A(n2624), .ZN(n2627) );
  NAND2_X1 U3362 ( .A1(n2627), .A2(n2642), .ZN(n4300) );
  OR2_X1 U3363 ( .A1(n2148), .A2(n4300), .ZN(n2628) );
  NAND4_X1 U3364 ( .A1(n2631), .A2(n2630), .A3(n2629), .A4(n2628), .ZN(n4408)
         );
  INV_X1 U3365 ( .A(n4408), .ZN(n4277) );
  MUX2_X1 U3366 ( .A(IR_REG_31__SCAN_IN), .B(n2635), .S(IR_REG_17__SCAN_IN), 
        .Z(n2636) );
  INV_X1 U3367 ( .A(n2636), .ZN(n2637) );
  NOR2_X1 U3368 ( .A1(n2637), .A2(n2657), .ZN(n4629) );
  INV_X1 U3369 ( .A(n4629), .ZN(n4601) );
  INV_X1 U3370 ( .A(DATAI_17_), .ZN(n2638) );
  MUX2_X1 U3371 ( .A(n4601), .B(n2638), .S(n2152), .Z(n4304) );
  NAND2_X1 U3372 ( .A1(n4277), .A2(n4304), .ZN(n2640) );
  AND2_X1 U3373 ( .A1(n4408), .A2(n4398), .ZN(n2639) );
  NAND2_X1 U3374 ( .A1(n2149), .A2(REG2_REG_18__SCAN_IN), .ZN(n2647) );
  NAND2_X1 U3375 ( .A1(n2150), .A2(REG0_REG_18__SCAN_IN), .ZN(n2646) );
  INV_X1 U3376 ( .A(REG1_REG_18__SCAN_IN), .ZN(n2641) );
  OR2_X1 U3377 ( .A1(n2145), .A2(n2641), .ZN(n2645) );
  AND2_X1 U3378 ( .A1(n2642), .A2(n4862), .ZN(n2643) );
  OR2_X1 U3379 ( .A1(n2643), .A2(n2651), .ZN(n4287) );
  OR2_X1 U3380 ( .A1(n2148), .A2(n4287), .ZN(n2644) );
  NAND4_X1 U3381 ( .A1(n2647), .A2(n2646), .A3(n2645), .A4(n2644), .ZN(n4399)
         );
  INV_X1 U3382 ( .A(n2657), .ZN(n2648) );
  NAND2_X1 U3383 ( .A1(n2648), .A2(IR_REG_31__SCAN_IN), .ZN(n2649) );
  MUX2_X1 U3384 ( .A(n4059), .B(DATAI_18_), .S(n2151), .Z(n4274) );
  NAND2_X1 U3385 ( .A1(n3745), .A2(n4274), .ZN(n4252) );
  NAND2_X1 U3386 ( .A1(n4399), .A2(n4284), .ZN(n4253) );
  NAND2_X1 U3387 ( .A1(n4252), .A2(n4253), .ZN(n4281) );
  NAND2_X1 U3388 ( .A1(n3745), .A2(n4284), .ZN(n2650) );
  NAND2_X1 U3389 ( .A1(n2149), .A2(REG2_REG_19__SCAN_IN), .ZN(n2656) );
  NAND2_X1 U3390 ( .A1(n2458), .A2(REG0_REG_19__SCAN_IN), .ZN(n2655) );
  INV_X1 U3391 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4392) );
  OR2_X1 U3392 ( .A1(n2145), .A2(n4392), .ZN(n2654) );
  OR2_X1 U3393 ( .A1(n2651), .A2(REG3_REG_19__SCAN_IN), .ZN(n2652) );
  NAND2_X1 U3394 ( .A1(n2660), .A2(n2652), .ZN(n4267) );
  OR2_X1 U3395 ( .A1(n2148), .A2(n4267), .ZN(n2653) );
  NAND4_X1 U3396 ( .A1(n2656), .A2(n2655), .A3(n2654), .A4(n2653), .ZN(n4275)
         );
  NAND2_X1 U3397 ( .A1(n2657), .A2(n4878), .ZN(n2658) );
  MUX2_X1 U3398 ( .A(n3539), .B(DATAI_19_), .S(n2152), .Z(n4263) );
  INV_X1 U3399 ( .A(n4263), .ZN(n4257) );
  NAND2_X1 U3400 ( .A1(n4233), .A2(n4257), .ZN(n2659) );
  NAND2_X1 U3401 ( .A1(n2149), .A2(REG2_REG_20__SCAN_IN), .ZN(n2665) );
  NAND2_X1 U3402 ( .A1(n2458), .A2(REG0_REG_20__SCAN_IN), .ZN(n2664) );
  INV_X1 U3403 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4776) );
  OR2_X1 U3404 ( .A1(n2145), .A2(n4776), .ZN(n2663) );
  NAND2_X1 U3405 ( .A1(n2660), .A2(n3767), .ZN(n2661) );
  NAND2_X1 U3406 ( .A1(n2666), .A2(n2661), .ZN(n4243) );
  OR2_X1 U3407 ( .A1(n2148), .A2(n4243), .ZN(n2662) );
  NAND4_X1 U3408 ( .A1(n2665), .A2(n2664), .A3(n2663), .A4(n2662), .ZN(n4214)
         );
  INV_X1 U3409 ( .A(n4210), .ZN(n2672) );
  AND2_X1 U3410 ( .A1(n2666), .A2(n3705), .ZN(n2667) );
  OR2_X1 U3411 ( .A1(n2667), .A2(n2673), .ZN(n4215) );
  NAND2_X1 U3412 ( .A1(n2149), .A2(REG2_REG_21__SCAN_IN), .ZN(n2669) );
  INV_X1 U3413 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4384) );
  OR2_X1 U3414 ( .A1(n2145), .A2(n4384), .ZN(n2668) );
  AND2_X1 U3415 ( .A1(n2669), .A2(n2668), .ZN(n2671) );
  NAND2_X1 U3416 ( .A1(n2150), .A2(REG0_REG_21__SCAN_IN), .ZN(n2670) );
  OAI211_X1 U3417 ( .C1(n2148), .C2(n4215), .A(n2671), .B(n2670), .ZN(n4231)
         );
  INV_X1 U3418 ( .A(n4219), .ZN(n4377) );
  INV_X1 U3419 ( .A(n4231), .ZN(n3788) );
  NOR2_X1 U3420 ( .A1(n2673), .A2(REG3_REG_22__SCAN_IN), .ZN(n2674) );
  OR2_X1 U3421 ( .A1(n2677), .A2(n2674), .ZN(n4201) );
  AOI22_X1 U3422 ( .A1(n2685), .A2(REG1_REG_22__SCAN_IN), .B1(n2149), .B2(
        REG2_REG_22__SCAN_IN), .ZN(n2676) );
  NAND2_X1 U3423 ( .A1(n2150), .A2(REG0_REG_22__SCAN_IN), .ZN(n2675) );
  OAI211_X1 U3424 ( .C1(n4201), .C2(n2148), .A(n2676), .B(n2675), .ZN(n4378)
         );
  OR2_X1 U3425 ( .A1(n4378), .A2(n4198), .ZN(n4172) );
  NAND2_X1 U3426 ( .A1(n4378), .A2(n4198), .ZN(n2742) );
  NAND2_X1 U3427 ( .A1(n4172), .A2(n2742), .ZN(n4189) );
  INV_X1 U3428 ( .A(n4378), .ZN(n4175) );
  OR2_X1 U3429 ( .A1(n2677), .A2(REG3_REG_23__SCAN_IN), .ZN(n2678) );
  NAND2_X1 U3430 ( .A1(n2682), .A2(n2678), .ZN(n4183) );
  AOI22_X1 U3431 ( .A1(n2685), .A2(REG1_REG_23__SCAN_IN), .B1(n2458), .B2(
        REG0_REG_23__SCAN_IN), .ZN(n2680) );
  NAND2_X1 U3432 ( .A1(n2149), .A2(REG2_REG_23__SCAN_IN), .ZN(n2679) );
  INV_X1 U3433 ( .A(n4358), .ZN(n3789) );
  NAND2_X1 U3434 ( .A1(n3789), .A2(n4181), .ZN(n2681) );
  INV_X1 U3435 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4158) );
  NAND2_X1 U3436 ( .A1(n2682), .A2(n3755), .ZN(n2683) );
  NAND2_X1 U3437 ( .A1(n2684), .A2(n2683), .ZN(n4159) );
  OR2_X1 U3438 ( .A1(n4159), .A2(n2148), .ZN(n2687) );
  AOI22_X1 U3439 ( .A1(n2685), .A2(REG1_REG_24__SCAN_IN), .B1(n2150), .B2(
        REG0_REG_24__SCAN_IN), .ZN(n2686) );
  INV_X1 U3440 ( .A(n4177), .ZN(n4139) );
  INV_X1 U3441 ( .A(n4129), .ZN(n4344) );
  NOR2_X1 U3442 ( .A1(n2692), .A2(n4672), .ZN(n2700) );
  INV_X1 U3443 ( .A(n2700), .ZN(n2702) );
  NAND2_X1 U3444 ( .A1(n2692), .A2(n4672), .ZN(n2693) );
  NAND2_X1 U3445 ( .A1(n2702), .A2(n2693), .ZN(n3641) );
  INV_X1 U3446 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4342) );
  NAND2_X1 U3447 ( .A1(n2149), .A2(REG2_REG_27__SCAN_IN), .ZN(n2695) );
  NAND2_X1 U3448 ( .A1(n2458), .A2(REG0_REG_27__SCAN_IN), .ZN(n2694) );
  OAI211_X1 U3449 ( .C1(n2145), .C2(n4342), .A(n2695), .B(n2694), .ZN(n2696)
         );
  INV_X1 U3450 ( .A(n2696), .ZN(n2697) );
  NOR2_X1 U3451 ( .A1(n4345), .A2(n4335), .ZN(n2699) );
  NAND2_X1 U3452 ( .A1(n2700), .A2(REG3_REG_28__SCAN_IN), .ZN(n4082) );
  INV_X1 U3453 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2701) );
  NAND2_X1 U3454 ( .A1(n2702), .A2(n2701), .ZN(n2703) );
  NAND2_X1 U3455 ( .A1(n4082), .A2(n2703), .ZN(n4090) );
  INV_X1 U3456 ( .A(REG1_REG_28__SCAN_IN), .ZN(n4915) );
  NAND2_X1 U3457 ( .A1(n2149), .A2(REG2_REG_28__SCAN_IN), .ZN(n2705) );
  NAND2_X1 U34580 ( .A1(n2150), .A2(REG0_REG_28__SCAN_IN), .ZN(n2704) );
  OAI211_X1 U34590 ( .C1(n2145), .C2(n4915), .A(n2705), .B(n2704), .ZN(n2706)
         );
  INV_X1 U3460 ( .A(n2706), .ZN(n2707) );
  INV_X1 U3461 ( .A(n3849), .ZN(n2709) );
  INV_X1 U3462 ( .A(n4092), .ZN(n3678) );
  NAND2_X1 U3463 ( .A1(n4108), .A2(n3678), .ZN(n3853) );
  NAND2_X1 U3464 ( .A1(n2709), .A2(n3853), .ZN(n2801) );
  OR2_X1 U3465 ( .A1(n4082), .A2(n2148), .ZN(n2714) );
  NAND2_X1 U3466 ( .A1(n2149), .A2(REG2_REG_29__SCAN_IN), .ZN(n2711) );
  NAND2_X1 U34670 ( .A1(n2458), .A2(REG0_REG_29__SCAN_IN), .ZN(n2710) );
  OAI211_X1 U3468 ( .C1(n2789), .C2(n2145), .A(n2711), .B(n2710), .ZN(n2712)
         );
  INV_X1 U34690 ( .A(n2712), .ZN(n2713) );
  NAND2_X1 U3470 ( .A1(n2714), .A2(n2713), .ZN(n4093) );
  NAND2_X1 U34710 ( .A1(n2152), .A2(DATAI_29_), .ZN(n4077) );
  XNOR2_X1 U3472 ( .A(n4093), .B(n4077), .ZN(n3904) );
  NAND2_X1 U34730 ( .A1(n2718), .A2(IR_REG_31__SCAN_IN), .ZN(n2719) );
  MUX2_X1 U3474 ( .A(IR_REG_31__SCAN_IN), .B(n2719), .S(IR_REG_21__SCAN_IN), 
        .Z(n2721) );
  NAND2_X1 U34750 ( .A1(n2231), .A2(IR_REG_31__SCAN_IN), .ZN(n2722) );
  XNOR2_X1 U3476 ( .A(n3012), .B(n4500), .ZN(n2723) );
  NAND2_X1 U34770 ( .A1(n2723), .A2(n4065), .ZN(n4237) );
  NAND2_X1 U3478 ( .A1(n3978), .A2(n3539), .ZN(n4617) );
  INV_X1 U34790 ( .A(n2993), .ZN(n2969) );
  NOR2_X1 U3480 ( .A1(n3998), .A2(n2969), .ZN(n3914) );
  NAND2_X1 U34810 ( .A1(n3872), .A2(n3914), .ZN(n2815) );
  NAND2_X1 U3482 ( .A1(n2815), .A2(n3915), .ZN(n3069) );
  NAND2_X1 U34830 ( .A1(n3069), .A2(n2725), .ZN(n3068) );
  NAND2_X1 U3484 ( .A1(n3068), .A2(n2726), .ZN(n3077) );
  NAND2_X1 U34850 ( .A1(n3141), .A2(n3043), .ZN(n3920) );
  NAND2_X1 U3486 ( .A1(n3529), .A2(n3117), .ZN(n3917) );
  NAND2_X1 U34870 ( .A1(n3077), .A2(n3871), .ZN(n3076) );
  NAND2_X1 U3488 ( .A1(n3076), .A2(n3920), .ZN(n3527) );
  INV_X1 U34890 ( .A(n3921), .ZN(n2727) );
  AND2_X1 U3490 ( .A1(n3996), .A2(n3230), .ZN(n3149) );
  NAND2_X1 U34910 ( .A1(n3252), .A2(n3154), .ZN(n3939) );
  NAND2_X1 U3492 ( .A1(n3224), .A2(n3254), .ZN(n3938) );
  NAND2_X1 U34930 ( .A1(n3192), .A2(n3938), .ZN(n2728) );
  NAND2_X1 U3494 ( .A1(n3301), .A2(n3200), .ZN(n3926) );
  NAND2_X1 U34950 ( .A1(n2728), .A2(n3926), .ZN(n3209) );
  INV_X1 U3496 ( .A(n2729), .ZN(n2730) );
  NAND2_X1 U34970 ( .A1(n3374), .A2(n3324), .ZN(n3930) );
  NAND2_X1 U3498 ( .A1(n3993), .A2(n3376), .ZN(n3936) );
  NAND2_X1 U34990 ( .A1(n2294), .A2(n3369), .ZN(n3931) );
  NAND2_X1 U3500 ( .A1(n2731), .A2(n3931), .ZN(n3280) );
  NAND2_X1 U35010 ( .A1(n3992), .A2(n3394), .ZN(n3946) );
  NAND2_X1 U3502 ( .A1(n3280), .A2(n3946), .ZN(n2732) );
  INV_X1 U35030 ( .A(n3992), .ZN(n3475) );
  NAND2_X1 U3504 ( .A1(n3475), .A2(n3391), .ZN(n3943) );
  NAND2_X1 U35050 ( .A1(n2732), .A2(n3943), .ZN(n3404) );
  NAND2_X1 U35060 ( .A1(n3404), .A2(n3947), .ZN(n2733) );
  NAND2_X1 U35070 ( .A1(n2733), .A2(n3911), .ZN(n3431) );
  NAND2_X1 U35080 ( .A1(n3991), .A2(n3716), .ZN(n3429) );
  NAND2_X1 U35090 ( .A1(n3484), .A2(n3780), .ZN(n3432) );
  AND2_X1 U35100 ( .A1(n3429), .A2(n3432), .ZN(n3948) );
  NAND2_X1 U35110 ( .A1(n3431), .A2(n3948), .ZN(n2734) );
  NOR2_X1 U35120 ( .A1(n3991), .A2(n3716), .ZN(n3430) );
  NOR2_X1 U35130 ( .A1(n3484), .A2(n3780), .ZN(n3433) );
  AOI21_X1 U35140 ( .B1(n3948), .B2(n3430), .A(n3433), .ZN(n3909) );
  NAND2_X1 U35150 ( .A1(n2734), .A2(n3909), .ZN(n3836) );
  NAND2_X1 U35160 ( .A1(n3836), .A2(n3897), .ZN(n2735) );
  NAND2_X1 U35170 ( .A1(n2735), .A2(n3832), .ZN(n3510) );
  NAND2_X1 U35180 ( .A1(n4410), .A2(n4417), .ZN(n3835) );
  NAND2_X1 U35190 ( .A1(n4430), .A2(n3825), .ZN(n3834) );
  NAND2_X1 U35200 ( .A1(n3835), .A2(n3834), .ZN(n3867) );
  AND2_X1 U35210 ( .A1(n4408), .A2(n4304), .ZN(n3887) );
  NAND2_X1 U35220 ( .A1(n4275), .A2(n4257), .ZN(n3888) );
  NAND2_X1 U35230 ( .A1(n4253), .A2(n3888), .ZN(n2736) );
  INV_X1 U35240 ( .A(n4230), .ZN(n4241) );
  AND2_X1 U35250 ( .A1(n4214), .A2(n4241), .ZN(n3838) );
  NAND2_X1 U35260 ( .A1(n4277), .A2(n4398), .ZN(n4250) );
  NAND2_X1 U35270 ( .A1(n4252), .A2(n4250), .ZN(n2737) );
  INV_X1 U35280 ( .A(n2736), .ZN(n3839) );
  NAND2_X1 U35290 ( .A1(n2737), .A2(n3839), .ZN(n2738) );
  NAND2_X1 U35300 ( .A1(n4233), .A2(n4263), .ZN(n3889) );
  NAND2_X1 U35310 ( .A1(n2738), .A2(n3889), .ZN(n4225) );
  NOR2_X1 U35320 ( .A1(n4214), .A2(n4241), .ZN(n2739) );
  OR2_X1 U35330 ( .A1(n4225), .A2(n2739), .ZN(n2741) );
  INV_X1 U35340 ( .A(n3838), .ZN(n2740) );
  NAND2_X1 U35350 ( .A1(n2741), .A2(n2740), .ZN(n3842) );
  OR2_X1 U35360 ( .A1(n4231), .A2(n4219), .ZN(n4169) );
  AND2_X1 U35370 ( .A1(n4172), .A2(n4169), .ZN(n3961) );
  INV_X1 U35380 ( .A(n3961), .ZN(n3843) );
  NAND2_X1 U35390 ( .A1(n4358), .A2(n4181), .ZN(n3865) );
  AND2_X1 U35400 ( .A1(n3865), .A2(n2742), .ZN(n3968) );
  AND2_X1 U35410 ( .A1(n4231), .A2(n4219), .ZN(n3963) );
  NAND2_X1 U35420 ( .A1(n4172), .A2(n3963), .ZN(n2743) );
  NAND2_X1 U35430 ( .A1(n3968), .A2(n2743), .ZN(n3846) );
  INV_X1 U35440 ( .A(n3846), .ZN(n2744) );
  OR2_X1 U35450 ( .A1(n4358), .A2(n4181), .ZN(n3866) );
  NOR2_X1 U35460 ( .A1(n4177), .A2(n4157), .ZN(n3882) );
  OR2_X1 U35470 ( .A1(n4162), .A2(n4145), .ZN(n4118) );
  OAI21_X1 U35480 ( .B1(n4336), .B2(n4129), .A(n4118), .ZN(n3966) );
  NAND2_X1 U35490 ( .A1(n4162), .A2(n4145), .ZN(n3869) );
  NAND2_X1 U35500 ( .A1(n4177), .A2(n4157), .ZN(n4135) );
  AND2_X1 U35510 ( .A1(n3869), .A2(n4135), .ZN(n4117) );
  OR2_X1 U35520 ( .A1(n4117), .A2(n3966), .ZN(n2745) );
  NAND2_X1 U35530 ( .A1(n4336), .A2(n4129), .ZN(n3854) );
  NAND2_X1 U35540 ( .A1(n2745), .A2(n3854), .ZN(n3971) );
  INV_X1 U35550 ( .A(n3971), .ZN(n2746) );
  XNOR2_X1 U35560 ( .A(n4345), .B(n4335), .ZN(n3879) );
  NOR2_X1 U35570 ( .A1(n4345), .A2(n4112), .ZN(n3848) );
  XOR2_X1 U35580 ( .A(n2747), .B(n3904), .Z(n2758) );
  INV_X1 U35590 ( .A(n3978), .ZN(n4502) );
  NAND2_X1 U35600 ( .A1(n4502), .A2(n4501), .ZN(n3862) );
  NAND2_X1 U35610 ( .A1(n3539), .A2(n4500), .ZN(n2748) );
  NAND2_X1 U35620 ( .A1(n2149), .A2(REG2_REG_30__SCAN_IN), .ZN(n2752) );
  NAND2_X1 U35630 ( .A1(n2458), .A2(REG0_REG_30__SCAN_IN), .ZN(n2751) );
  INV_X1 U35640 ( .A(REG1_REG_30__SCAN_IN), .ZN(n2749) );
  OR2_X1 U35650 ( .A1(n2145), .A2(n2749), .ZN(n2750) );
  XNOR2_X1 U35660 ( .A(n2755), .B(n2753), .ZN(n2954) );
  INV_X1 U35670 ( .A(B_REG_SCAN_IN), .ZN(n2757) );
  NAND2_X1 U35680 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(
        n2754) );
  NAND2_X1 U35690 ( .A1(n2755), .A2(n2754), .ZN(n2756) );
  OAI21_X1 U35700 ( .B1(n2954), .B2(n2757), .A(n4429), .ZN(n4071) );
  OAI22_X1 U35710 ( .A1(n2758), .A2(n4261), .B1(n3861), .B2(n4071), .ZN(n4084)
         );
  INV_X1 U35720 ( .A(n4500), .ZN(n2760) );
  INV_X1 U35730 ( .A(n4501), .ZN(n2759) );
  OAI22_X1 U35740 ( .A1(n4338), .A2(n4432), .B1(n4077), .B2(n4258), .ZN(n2761)
         );
  AOI21_X1 U35750 ( .B1(n4076), .B2(n4423), .A(n2762), .ZN(n2795) );
  OR2_X1 U35760 ( .A1(n2169), .A2(n2846), .ZN(n2776) );
  NAND2_X1 U35770 ( .A1(n2776), .A2(n2775), .ZN(n2763) );
  NAND2_X1 U35780 ( .A1(n2766), .A2(IR_REG_31__SCAN_IN), .ZN(n2767) );
  MUX2_X1 U35790 ( .A(IR_REG_31__SCAN_IN), .B(n2767), .S(IR_REG_25__SCAN_IN), 
        .Z(n2768) );
  NAND2_X1 U35800 ( .A1(n2840), .A2(n2853), .ZN(n2769) );
  MUX2_X1 U35810 ( .A(n2840), .B(n2769), .S(B_REG_SCAN_IN), .Z(n2773) );
  NAND2_X1 U3582 ( .A1(n2172), .A2(IR_REG_31__SCAN_IN), .ZN(n2770) );
  INV_X1 U3583 ( .A(D_REG_1__SCAN_IN), .ZN(n2855) );
  NAND2_X1 U3584 ( .A1(n2850), .A2(n2855), .ZN(n2973) );
  NAND2_X1 U3585 ( .A1(n2787), .A2(n2853), .ZN(n2818) );
  NAND2_X1 U3586 ( .A1(n2973), .A2(n2818), .ZN(n2786) );
  NAND2_X1 U3587 ( .A1(n3978), .A2(n4065), .ZN(n2978) );
  NOR3_X1 U3588 ( .A1(D_REG_12__SCAN_IN), .A2(D_REG_2__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .ZN(n2779) );
  NOR4_X1 U3589 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_19__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2778) );
  NOR4_X1 U3590 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_26__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2777) );
  NAND3_X1 U3591 ( .A1(n2779), .A2(n2778), .A3(n2777), .ZN(n4932) );
  NOR4_X1 U3592 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_28__SCAN_IN), .ZN(n2784) );
  NOR4_X1 U3593 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(n2780), .ZN(n2783) );
  NOR4_X1 U3594 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_13__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2782) );
  NOR4_X1 U3595 ( .A1(D_REG_3__SCAN_IN), .A2(D_REG_4__SCAN_IN), .A3(
        D_REG_7__SCAN_IN), .A4(D_REG_10__SCAN_IN), .ZN(n2781) );
  NAND4_X1 U3596 ( .A1(n2784), .A2(n2783), .A3(n2782), .A4(n2781), .ZN(n2785)
         );
  OAI21_X1 U3597 ( .B1(n4932), .B2(n2785), .A(n2850), .ZN(n2819) );
  NAND4_X1 U3598 ( .A1(n2786), .A2(n2821), .A3(n2819), .A4(n2822), .ZN(n2794)
         );
  NAND2_X1 U3599 ( .A1(n2850), .A2(n2859), .ZN(n2788) );
  NAND2_X1 U3600 ( .A1(n2787), .A2(n2840), .ZN(n2856) );
  MUX2_X1 U3601 ( .A(n2789), .B(n2795), .S(n4657), .Z(n2793) );
  NAND2_X1 U3602 ( .A1(n3023), .A2(n2969), .ZN(n3073) );
  NOR2_X1 U3603 ( .A1(n3073), .A2(n3066), .ZN(n3081) );
  NAND2_X1 U3604 ( .A1(n3282), .A2(n3394), .ZN(n3409) );
  NAND2_X1 U3605 ( .A1(n3459), .A2(n3652), .ZN(n3514) );
  NAND2_X1 U3606 ( .A1(n2807), .A2(n4077), .ZN(n4331) );
  NAND2_X1 U3607 ( .A1(n2793), .A2(n2792), .ZN(U3547) );
  INV_X1 U3608 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2796) );
  NOR2_X4 U3609 ( .A1(n2794), .A2(n2975), .ZN(n4475) );
  MUX2_X1 U3610 ( .A(n2796), .B(n2795), .S(n4475), .Z(n2798) );
  NAND2_X1 U3611 ( .A1(n2798), .A2(n2797), .ZN(U3515) );
  INV_X1 U3612 ( .A(REG0_REG_28__SCAN_IN), .ZN(n2806) );
  XNOR2_X1 U3613 ( .A(n2800), .B(n2799), .ZN(n4087) );
  XNOR2_X1 U3614 ( .A(n2802), .B(n2799), .ZN(n2803) );
  NAND2_X1 U3615 ( .A1(n2803), .A2(n4437), .ZN(n4088) );
  AOI22_X1 U3616 ( .A1(n4093), .A2(n4429), .B1(n4427), .B2(n4092), .ZN(n2804)
         );
  OAI211_X1 U3617 ( .C1(n3906), .C2(n4432), .A(n4088), .B(n2804), .ZN(n2805)
         );
  MUX2_X1 U3618 ( .A(n2806), .B(n3543), .S(n4475), .Z(n2811) );
  INV_X1 U3619 ( .A(n4106), .ZN(n2809) );
  INV_X1 U3620 ( .A(n2807), .ZN(n2808) );
  OAI21_X1 U3621 ( .B1(n2809), .B2(n3678), .A(n2808), .ZN(n4096) );
  NAND2_X1 U3622 ( .A1(n2811), .A2(n2810), .ZN(U3514) );
  NAND2_X1 U3623 ( .A1(n3062), .A2(n2813), .ZN(n3100) );
  INV_X1 U3624 ( .A(n3914), .ZN(n2970) );
  NAND2_X1 U3625 ( .A1(n2815), .A2(n2814), .ZN(n2816) );
  NAND2_X1 U3626 ( .A1(n2816), .A2(n4437), .ZN(n2817) );
  OAI21_X1 U3627 ( .B1(n3100), .B2(n4237), .A(n2817), .ZN(n3104) );
  AND2_X1 U3628 ( .A1(n2819), .A2(n2818), .ZN(n2974) );
  NAND4_X1 U3629 ( .A1(n2974), .A2(n2821), .A3(n2820), .A4(n2973), .ZN(n2824)
         );
  MUX2_X1 U3630 ( .A(REG2_REG_1__SCAN_IN), .B(n3104), .S(n4606), .Z(n2833) );
  OR2_X1 U3631 ( .A1(n3012), .A2(n4065), .ZN(n3110) );
  INV_X1 U3632 ( .A(n3110), .ZN(n2825) );
  NAND2_X1 U3633 ( .A1(n4606), .A2(n2825), .ZN(n4608) );
  INV_X1 U3634 ( .A(n4603), .ZN(n4619) );
  AOI22_X1 U3635 ( .A1(n4161), .A2(n3101), .B1(REG3_REG_1__SCAN_IN), .B2(n4619), .ZN(n2826) );
  OAI21_X1 U3636 ( .B1(n3100), .B2(n4608), .A(n2826), .ZN(n2832) );
  NAND2_X1 U3637 ( .A1(n3101), .A2(n2993), .ZN(n2827) );
  NAND2_X1 U3638 ( .A1(n3073), .A2(n2827), .ZN(n3276) );
  NAND2_X1 U3639 ( .A1(n4313), .A2(n2828), .ZN(n2830) );
  NAND2_X1 U3640 ( .A1(n4238), .A2(n4357), .ZN(n4079) );
  NAND2_X1 U3641 ( .A1(n4314), .A2(n3998), .ZN(n2829) );
  OAI211_X1 U3642 ( .C1(n4266), .C2(n3276), .A(n2830), .B(n2829), .ZN(n2831)
         );
  OR3_X1 U3643 ( .A1(n2833), .A2(n2832), .A3(n2831), .ZN(U3289) );
  MUX2_X1 U3644 ( .A(n2834), .B(n3173), .S(STATE_REG_SCAN_IN), .Z(n2835) );
  INV_X1 U3645 ( .A(n2835), .ZN(U3344) );
  INV_X1 U3646 ( .A(DATAI_16_), .ZN(n2837) );
  NAND2_X1 U3647 ( .A1(n4049), .A2(STATE_REG_SCAN_IN), .ZN(n2836) );
  OAI21_X1 U3648 ( .B1(STATE_REG_SCAN_IN), .B2(n2837), .A(n2836), .ZN(U3336)
         );
  INV_X1 U3649 ( .A(DATAI_18_), .ZN(n2839) );
  NAND2_X1 U3650 ( .A1(n4059), .A2(STATE_REG_SCAN_IN), .ZN(n2838) );
  OAI21_X1 U3651 ( .B1(STATE_REG_SCAN_IN), .B2(n2839), .A(n2838), .ZN(U3334)
         );
  INV_X1 U3652 ( .A(DATAI_24_), .ZN(n4872) );
  MUX2_X1 U3653 ( .A(n2840), .B(n4872), .S(U3149), .Z(n2841) );
  INV_X1 U3654 ( .A(n2841), .ZN(U3328) );
  INV_X1 U3655 ( .A(DATAI_19_), .ZN(n4664) );
  MUX2_X1 U3656 ( .A(n4664), .B(n4065), .S(STATE_REG_SCAN_IN), .Z(n2842) );
  INV_X1 U3657 ( .A(n2842), .ZN(U3333) );
  INV_X1 U3658 ( .A(DATAI_27_), .ZN(n4660) );
  INV_X1 U3659 ( .A(n2954), .ZN(n2862) );
  NAND2_X1 U3660 ( .A1(n2862), .A2(STATE_REG_SCAN_IN), .ZN(n2843) );
  OAI21_X1 U3661 ( .B1(STATE_REG_SCAN_IN), .B2(n4660), .A(n2843), .ZN(U3325)
         );
  INV_X1 U3662 ( .A(DATAI_29_), .ZN(n4866) );
  NAND2_X1 U3663 ( .A1(n2844), .A2(STATE_REG_SCAN_IN), .ZN(n2845) );
  OAI21_X1 U3664 ( .B1(STATE_REG_SCAN_IN), .B2(n4866), .A(n2845), .ZN(U3323)
         );
  INV_X1 U3665 ( .A(DATAI_31_), .ZN(n4864) );
  OR4_X1 U3666 ( .A1(n2425), .A2(IR_REG_30__SCAN_IN), .A3(n2846), .A4(U3149), 
        .ZN(n2847) );
  OAI21_X1 U3667 ( .B1(STATE_REG_SCAN_IN), .B2(n4864), .A(n2847), .ZN(U3321)
         );
  INV_X1 U3668 ( .A(DATAI_30_), .ZN(n4865) );
  NAND2_X1 U3669 ( .A1(n2848), .A2(STATE_REG_SCAN_IN), .ZN(n2849) );
  OAI21_X1 U3670 ( .B1(STATE_REG_SCAN_IN), .B2(n4865), .A(n2849), .ZN(U3322)
         );
  INV_X1 U3671 ( .A(n2853), .ZN(n4499) );
  NOR3_X1 U3672 ( .A1(n4498), .A2(n4499), .A3(n4627), .ZN(n2854) );
  AOI21_X1 U3673 ( .B1(n4942), .B2(n2855), .A(n2854), .ZN(U3459) );
  INV_X1 U3674 ( .A(n2856), .ZN(n2858) );
  AOI22_X1 U3675 ( .A1(n4942), .A2(n2859), .B1(n2858), .B2(n2857), .ZN(U3458)
         );
  NAND2_X1 U3676 ( .A1(n3051), .A2(n2979), .ZN(n2860) );
  INV_X1 U3677 ( .A(n2866), .ZN(n2861) );
  OR2_X1 U3678 ( .A1(n3051), .A2(U3149), .ZN(n3988) );
  NAND2_X1 U3679 ( .A1(n2989), .A2(n3988), .ZN(n2865) );
  INV_X1 U3680 ( .A(ADDR_REG_0__SCAN_IN), .ZN(n2870) );
  INV_X1 U3681 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4623) );
  AOI21_X1 U3682 ( .B1(n2862), .B2(n4623), .A(n2997), .ZN(n2956) );
  OAI21_X1 U3683 ( .B1(n2862), .B2(REG1_REG_0__SCAN_IN), .A(n2367), .ZN(n2864)
         );
  NOR2_X1 U3684 ( .A1(n2956), .A2(n4877), .ZN(n2863) );
  AOI21_X1 U3685 ( .B1(n2956), .B2(n2864), .A(n2863), .ZN(n2867) );
  AOI22_X1 U3686 ( .A1(n2867), .A2(n2872), .B1(REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n2869) );
  NAND3_X1 U3687 ( .A1(n4595), .A2(n4877), .A3(n2950), .ZN(n2868) );
  OAI211_X1 U3688 ( .C1(n4587), .C2(n2870), .A(n2869), .B(n2868), .ZN(U3240)
         );
  NOR2_X1 U3689 ( .A1(n4594), .A2(n3997), .ZN(U3148) );
  INV_X1 U3690 ( .A(REG2_REG_1__SCAN_IN), .ZN(n4002) );
  NAND2_X1 U3691 ( .A1(n4510), .A2(REG2_REG_1__SCAN_IN), .ZN(n4013) );
  INV_X1 U3692 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2871) );
  XNOR2_X1 U3693 ( .A(n2897), .B(REG2_REG_3__SCAN_IN), .ZN(n2881) );
  NOR2_X1 U3694 ( .A1(n2997), .A2(n2954), .ZN(n3984) );
  INV_X1 U3695 ( .A(n4602), .ZN(n4036) );
  INV_X1 U3696 ( .A(ADDR_REG_3__SCAN_IN), .ZN(n2873) );
  OAI22_X1 U3697 ( .A1(n4587), .A2(n2873), .B1(STATE_REG_SCAN_IN), .B2(n4894), 
        .ZN(n2874) );
  AOI21_X1 U3698 ( .B1(n4508), .B2(n4036), .A(n2874), .ZN(n2880) );
  XNOR2_X1 U3699 ( .A(n4509), .B(n4885), .ZN(n4020) );
  AND2_X1 U3700 ( .A1(n4877), .A2(REG1_REG_0__SCAN_IN), .ZN(n4000) );
  NAND2_X1 U3701 ( .A1(n4510), .A2(REG1_REG_1__SCAN_IN), .ZN(n2875) );
  NAND2_X1 U3702 ( .A1(n3999), .A2(n2875), .ZN(n4019) );
  NAND2_X1 U3703 ( .A1(n4020), .A2(n4019), .ZN(n4018) );
  NAND2_X1 U3704 ( .A1(n4509), .A2(REG1_REG_2__SCAN_IN), .ZN(n2876) );
  INV_X1 U3705 ( .A(n4508), .ZN(n2877) );
  XNOR2_X1 U3706 ( .A(n2901), .B(n2877), .ZN(n2878) );
  NAND2_X1 U3707 ( .A1(n2878), .A2(REG1_REG_3__SCAN_IN), .ZN(n2903) );
  OAI211_X1 U3708 ( .C1(REG1_REG_3__SCAN_IN), .C2(n2878), .A(n4595), .B(n2903), 
        .ZN(n2879) );
  OAI211_X1 U3709 ( .C1(n2881), .C2(n4588), .A(n2880), .B(n2879), .ZN(U3243)
         );
  INV_X1 U3710 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n4820) );
  NAND2_X1 U3711 ( .A1(n3225), .A2(U4043), .ZN(n2882) );
  OAI21_X1 U3712 ( .B1(n3997), .B2(n4820), .A(n2882), .ZN(U3554) );
  INV_X1 U3713 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n4842) );
  NAND2_X1 U3714 ( .A1(n2149), .A2(REG2_REG_31__SCAN_IN), .ZN(n2885) );
  NAND2_X1 U3715 ( .A1(n2150), .A2(REG0_REG_31__SCAN_IN), .ZN(n2884) );
  INV_X1 U3716 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4328) );
  OR2_X1 U3717 ( .A1(n2145), .A2(n4328), .ZN(n2883) );
  INV_X1 U3718 ( .A(n4072), .ZN(n3883) );
  NAND2_X1 U3719 ( .A1(n3883), .A2(U4043), .ZN(n2886) );
  OAI21_X1 U3720 ( .B1(n3997), .B2(n4842), .A(n2886), .ZN(U3581) );
  INV_X1 U3721 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n4836) );
  INV_X1 U3722 ( .A(n3861), .ZN(n2887) );
  NAND2_X1 U3723 ( .A1(n2887), .A2(U4043), .ZN(n2888) );
  OAI21_X1 U3724 ( .B1(U4043), .B2(n4836), .A(n2888), .ZN(U3580) );
  INV_X1 U3725 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n4923) );
  NAND2_X1 U3726 ( .A1(n3224), .A2(U4043), .ZN(n2889) );
  OAI21_X1 U3727 ( .B1(U4043), .B2(n4923), .A(n2889), .ZN(U3556) );
  INV_X1 U3728 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n4921) );
  NAND2_X1 U3729 ( .A1(n4214), .A2(n3997), .ZN(n2890) );
  OAI21_X1 U3730 ( .B1(n3997), .B2(n4921), .A(n2890), .ZN(U3570) );
  INV_X1 U3731 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n4920) );
  NAND2_X1 U3732 ( .A1(n3529), .A2(U4043), .ZN(n2891) );
  OAI21_X1 U3733 ( .B1(U4043), .B2(n4920), .A(n2891), .ZN(U3553) );
  INV_X1 U3734 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n4834) );
  NAND2_X1 U3735 ( .A1(n4162), .A2(n3997), .ZN(n2892) );
  OAI21_X1 U3736 ( .B1(n3997), .B2(n4834), .A(n2892), .ZN(U3575) );
  INV_X1 U3737 ( .A(DATAO_REG_15__SCAN_IN), .ZN(n4825) );
  NAND2_X1 U3738 ( .A1(n4430), .A2(n3997), .ZN(n2893) );
  OAI21_X1 U3739 ( .B1(n3997), .B2(n4825), .A(n2893), .ZN(U3565) );
  INV_X1 U3740 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n4919) );
  NAND2_X1 U3741 ( .A1(n2828), .A2(n3997), .ZN(n2894) );
  OAI21_X1 U3742 ( .B1(n3997), .B2(n4919), .A(n2894), .ZN(U3552) );
  INV_X1 U3743 ( .A(n2906), .ZN(n4506) );
  INV_X1 U3744 ( .A(n2895), .ZN(n2896) );
  XNOR2_X1 U3745 ( .A(n2898), .B(n4507), .ZN(n2959) );
  INV_X1 U3746 ( .A(n2898), .ZN(n2899) );
  INV_X1 U3747 ( .A(REG2_REG_5__SCAN_IN), .ZN(n4900) );
  MUX2_X1 U3748 ( .A(REG2_REG_5__SCAN_IN), .B(n4900), .S(n2906), .Z(n2936) );
  XNOR2_X1 U3749 ( .A(n2926), .B(REG2_REG_6__SCAN_IN), .ZN(n2911) );
  NAND2_X1 U3750 ( .A1(n4594), .A2(ADDR_REG_6__SCAN_IN), .ZN(n2900) );
  NAND2_X1 U3751 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3253) );
  NAND2_X1 U3752 ( .A1(n2900), .A2(n3253), .ZN(n2909) );
  NAND2_X1 U3753 ( .A1(n2901), .A2(n4508), .ZN(n2902) );
  NAND2_X1 U3754 ( .A1(n2903), .A2(n2902), .ZN(n2904) );
  INV_X1 U3755 ( .A(n2904), .ZN(n2905) );
  INV_X1 U3756 ( .A(n4507), .ZN(n2965) );
  XNOR2_X1 U3757 ( .A(n2904), .B(n2965), .ZN(n2961) );
  XNOR2_X1 U3758 ( .A(n2906), .B(REG1_REG_5__SCAN_IN), .ZN(n2942) );
  XNOR2_X1 U3759 ( .A(n2920), .B(n4505), .ZN(n2907) );
  NOR2_X1 U3760 ( .A1(n2907), .A2(n2504), .ZN(n2919) );
  INV_X1 U3761 ( .A(n4595), .ZN(n4580) );
  AOI211_X1 U3762 ( .C1(n2907), .C2(n2504), .A(n2919), .B(n4580), .ZN(n2908)
         );
  AOI211_X1 U3763 ( .C1(n4036), .C2(n4505), .A(n2909), .B(n2908), .ZN(n2910)
         );
  OAI21_X1 U3764 ( .B1(n2911), .B2(n4588), .A(n2910), .ZN(U3246) );
  INV_X1 U3765 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n4924) );
  NAND2_X1 U3766 ( .A1(n3483), .A2(n3997), .ZN(n2912) );
  OAI21_X1 U3767 ( .B1(n3997), .B2(n4924), .A(n2912), .ZN(U3561) );
  INV_X1 U3768 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n4832) );
  NAND2_X1 U3769 ( .A1(n4378), .A2(n3997), .ZN(n2913) );
  OAI21_X1 U3770 ( .B1(n3997), .B2(n4832), .A(n2913), .ZN(U3572) );
  INV_X1 U3771 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n4824) );
  NAND2_X1 U3772 ( .A1(n4399), .A2(n3997), .ZN(n2914) );
  OAI21_X1 U3773 ( .B1(n3997), .B2(n4824), .A(n2914), .ZN(U3568) );
  INV_X1 U3774 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n4922) );
  NAND2_X1 U3775 ( .A1(n4275), .A2(n3997), .ZN(n2915) );
  OAI21_X1 U3776 ( .B1(U4043), .B2(n4922), .A(n2915), .ZN(U3569) );
  INV_X1 U3777 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n4822) );
  NAND2_X1 U3778 ( .A1(n3484), .A2(n3997), .ZN(n2916) );
  OAI21_X1 U3779 ( .B1(n3997), .B2(n4822), .A(n2916), .ZN(U3563) );
  INV_X1 U3780 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n4917) );
  NAND2_X1 U3781 ( .A1(n4336), .A2(n3997), .ZN(n2917) );
  OAI21_X1 U3782 ( .B1(n3997), .B2(n4917), .A(n2917), .ZN(U3576) );
  INV_X1 U3783 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n4916) );
  NAND2_X1 U3784 ( .A1(n4177), .A2(n3997), .ZN(n2918) );
  OAI21_X1 U3785 ( .B1(n3997), .B2(n4916), .A(n2918), .ZN(U3574) );
  AOI21_X1 U3786 ( .B1(n4505), .B2(n2920), .A(n2919), .ZN(n3003) );
  MUX2_X1 U3787 ( .A(REG1_REG_7__SCAN_IN), .B(n2515), .S(n4504), .Z(n2921) );
  XNOR2_X1 U3788 ( .A(n3003), .B(n2921), .ZN(n2931) );
  INV_X1 U3789 ( .A(n4504), .ZN(n3001) );
  INV_X1 U3790 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2922) );
  OR2_X1 U3791 ( .A1(STATE_REG_SCAN_IN), .A2(n2922), .ZN(n3302) );
  NAND2_X1 U3792 ( .A1(n4594), .A2(ADDR_REG_7__SCAN_IN), .ZN(n2923) );
  OAI211_X1 U3793 ( .C1(n4602), .C2(n3001), .A(n3302), .B(n2923), .ZN(n2930)
         );
  INV_X1 U3794 ( .A(n2924), .ZN(n2925) );
  INV_X1 U3795 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3216) );
  MUX2_X1 U3796 ( .A(n3216), .B(REG2_REG_7__SCAN_IN), .S(n4504), .Z(n2927) );
  NOR2_X1 U3797 ( .A1(n2928), .A2(n2927), .ZN(n3004) );
  AOI211_X1 U3798 ( .C1(n2928), .C2(n2927), .A(n4588), .B(n3004), .ZN(n2929)
         );
  AOI211_X1 U3799 ( .C1(n4595), .C2(n2931), .A(n2930), .B(n2929), .ZN(n2932)
         );
  INV_X1 U3800 ( .A(n2932), .ZN(U3247) );
  INV_X1 U3801 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n4918) );
  NAND2_X1 U3802 ( .A1(n4345), .A2(n3997), .ZN(n2933) );
  OAI21_X1 U3803 ( .B1(n3997), .B2(n4918), .A(n2933), .ZN(U3577) );
  INV_X1 U3804 ( .A(ADDR_REG_5__SCAN_IN), .ZN(n2934) );
  OR2_X1 U3805 ( .A1(STATE_REG_SCAN_IN), .A2(n2489), .ZN(n3133) );
  OAI21_X1 U3806 ( .B1(n4587), .B2(n2934), .A(n3133), .ZN(n2939) );
  AOI211_X1 U3807 ( .C1(n2937), .C2(n2936), .A(n4588), .B(n2935), .ZN(n2938)
         );
  AOI211_X1 U3808 ( .C1(n4036), .C2(n4506), .A(n2939), .B(n2938), .ZN(n2944)
         );
  OAI211_X1 U3809 ( .C1(n2942), .C2(n2941), .A(n4595), .B(n2940), .ZN(n2943)
         );
  NAND2_X1 U3810 ( .A1(n2944), .A2(n2943), .ZN(U3245) );
  INV_X1 U3811 ( .A(n4412), .ZN(n3213) );
  AND2_X4 U3812 ( .A1(n3631), .A2(n3213), .ZN(n3636) );
  INV_X1 U3813 ( .A(n3012), .ZN(n2945) );
  INV_X1 U3814 ( .A(n3052), .ZN(n2946) );
  INV_X1 U3815 ( .A(n2948), .ZN(n2949) );
  NOR2_X1 U3816 ( .A1(n2952), .A2(n2953), .ZN(n3013) );
  AOI21_X1 U3817 ( .B1(n2953), .B2(n2952), .A(n3013), .ZN(n2994) );
  NAND2_X1 U3818 ( .A1(n4497), .A2(n2954), .ZN(n2958) );
  NAND2_X1 U3819 ( .A1(n3984), .A2(REG2_REG_0__SCAN_IN), .ZN(n2955) );
  MUX2_X1 U3820 ( .A(n2956), .B(n2955), .S(n4877), .Z(n2957) );
  OAI211_X1 U3821 ( .C1(n2994), .C2(n2958), .A(n3997), .B(n2957), .ZN(n4024)
         );
  XOR2_X1 U3822 ( .A(REG2_REG_4__SCAN_IN), .B(n2959), .Z(n2967) );
  OAI211_X1 U3823 ( .C1(REG1_REG_4__SCAN_IN), .C2(n2961), .A(n4595), .B(n2960), 
        .ZN(n2964) );
  NAND2_X1 U3824 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3095) );
  INV_X1 U3825 ( .A(n3095), .ZN(n2962) );
  AOI21_X1 U3826 ( .B1(n4594), .B2(ADDR_REG_4__SCAN_IN), .A(n2962), .ZN(n2963)
         );
  OAI211_X1 U3827 ( .C1(n4602), .C2(n2965), .A(n2964), .B(n2963), .ZN(n2966)
         );
  AOI21_X1 U3828 ( .B1(n4584), .B2(n2967), .A(n2966), .ZN(n2968) );
  NAND2_X1 U3829 ( .A1(n4024), .A2(n2968), .ZN(U3244) );
  INV_X1 U3830 ( .A(n3446), .ZN(n4645) );
  NAND2_X1 U3831 ( .A1(n3998), .A2(n2969), .ZN(n3913) );
  NAND2_X1 U3832 ( .A1(n2970), .A2(n3913), .ZN(n4621) );
  AND2_X1 U3833 ( .A1(n2993), .A2(n2977), .ZN(n4618) );
  INV_X1 U3834 ( .A(n4237), .ZN(n3350) );
  OAI21_X1 U3835 ( .B1(n3350), .B2(n4437), .A(n4621), .ZN(n2971) );
  OAI21_X1 U3836 ( .B1(n3015), .B2(n4361), .A(n2971), .ZN(n4616) );
  AOI211_X1 U3837 ( .C1(n4645), .C2(n4621), .A(n4618), .B(n4616), .ZN(n4640)
         );
  NAND2_X1 U3838 ( .A1(n4655), .A2(REG1_REG_0__SCAN_IN), .ZN(n2972) );
  OAI21_X1 U3839 ( .B1(n4640), .B2(n4655), .A(n2972), .ZN(U3518) );
  NAND3_X1 U3840 ( .A1(n2975), .A2(n2974), .A3(n2973), .ZN(n2996) );
  NAND2_X1 U3841 ( .A1(n4065), .A2(n4500), .ZN(n3011) );
  NOR2_X1 U3842 ( .A1(n3011), .A2(n4627), .ZN(n2976) );
  NAND2_X1 U3843 ( .A1(n3016), .A2(n2976), .ZN(n2995) );
  INV_X1 U3844 ( .A(n2995), .ZN(n3985) );
  NAND2_X1 U3845 ( .A1(n2996), .A2(n3985), .ZN(n3055) );
  INV_X1 U3846 ( .A(n3055), .ZN(n2986) );
  NAND2_X1 U3847 ( .A1(n2978), .A2(n2977), .ZN(n2981) );
  INV_X1 U3848 ( .A(n2979), .ZN(n2980) );
  NAND2_X1 U3849 ( .A1(n2981), .A2(n2980), .ZN(n2987) );
  NAND2_X1 U3850 ( .A1(n2987), .A2(n4258), .ZN(n2982) );
  NAND2_X1 U3851 ( .A1(n2996), .A2(n2982), .ZN(n2985) );
  INV_X1 U3852 ( .A(n2983), .ZN(n2984) );
  NAND2_X1 U3853 ( .A1(n2985), .A2(n2984), .ZN(n3054) );
  NOR3_X1 U3854 ( .A1(n2986), .A2(n3054), .A3(n2989), .ZN(n3037) );
  INV_X1 U3855 ( .A(n2996), .ZN(n2991) );
  NOR2_X1 U3856 ( .A1(n2989), .A2(n2987), .ZN(n2988) );
  NOR2_X1 U3857 ( .A1(n2989), .A2(n4258), .ZN(n2990) );
  NAND2_X1 U3858 ( .A1(n2991), .A2(n2990), .ZN(n2992) );
  AND2_X2 U3859 ( .A1(n2992), .A2(n4603), .ZN(n3810) );
  INV_X1 U3860 ( .A(n3810), .ZN(n3691) );
  AOI22_X1 U3861 ( .A1(n2994), .A2(n3820), .B1(n2993), .B2(n3691), .ZN(n2999)
         );
  NOR2_X1 U3862 ( .A1(n2996), .A2(n2995), .ZN(n3024) );
  NAND2_X2 U3863 ( .A1(n3024), .A2(n2997), .ZN(n3822) );
  INV_X1 U3864 ( .A(n3822), .ZN(n3689) );
  NAND2_X1 U3865 ( .A1(n3689), .A2(n3017), .ZN(n2998) );
  OAI211_X1 U3866 ( .C1(n3037), .C2(n3000), .A(n2999), .B(n2998), .ZN(U3229)
         );
  NOR2_X1 U3867 ( .A1(n4504), .A2(REG1_REG_7__SCAN_IN), .ZN(n3002) );
  OAI22_X1 U3868 ( .A1(n3003), .A2(n3002), .B1(n2515), .B2(n3001), .ZN(n3172)
         );
  XNOR2_X1 U3869 ( .A(n3172), .B(n3173), .ZN(n3171) );
  XNOR2_X1 U3870 ( .A(n3171), .B(REG1_REG_8__SCAN_IN), .ZN(n3010) );
  AOI21_X1 U3871 ( .B1(n4504), .B2(REG2_REG_7__SCAN_IN), .A(n3004), .ZN(n3160)
         );
  XNOR2_X1 U3872 ( .A(REG2_REG_8__SCAN_IN), .B(n3161), .ZN(n3005) );
  NAND2_X1 U3873 ( .A1(n4584), .A2(n3005), .ZN(n3006) );
  NAND2_X1 U3874 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3334) );
  NAND2_X1 U3875 ( .A1(n3006), .A2(n3334), .ZN(n3008) );
  NOR2_X1 U3876 ( .A1(n4602), .A2(n3173), .ZN(n3007) );
  AOI211_X1 U3877 ( .C1(n4594), .C2(ADDR_REG_8__SCAN_IN), .A(n3008), .B(n3007), 
        .ZN(n3009) );
  OAI21_X1 U3878 ( .B1(n3010), .B2(n4580), .A(n3009), .ZN(U3248) );
  AND2_X2 U3879 ( .A1(n3012), .A2(n3011), .ZN(n3675) );
  AOI21_X1 U3880 ( .B1(n3675), .B2(n3014), .A(n3013), .ZN(n3022) );
  INV_X2 U3881 ( .A(n3636), .ZN(n3042) );
  OAI22_X1 U3882 ( .A1(n3042), .A2(n3015), .B1(n3023), .B2(n3674), .ZN(n3031)
         );
  NAND2_X1 U3883 ( .A1(n3017), .A2(n3016), .ZN(n3019) );
  NAND2_X1 U3884 ( .A1(n3101), .A2(n2146), .ZN(n3018) );
  NAND2_X1 U3885 ( .A1(n3019), .A2(n3018), .ZN(n3020) );
  XNOR2_X1 U3886 ( .A(n3031), .B(n3032), .ZN(n3021) );
  NOR2_X1 U3887 ( .A1(n3022), .A2(n3021), .ZN(n3034) );
  AOI211_X1 U3888 ( .C1(n3022), .C2(n3021), .A(n3815), .B(n3034), .ZN(n3028)
         );
  OAI22_X1 U3889 ( .A1(n3029), .A2(n3822), .B1(n3810), .B2(n3023), .ZN(n3027)
         );
  INV_X1 U3890 ( .A(n3998), .ZN(n3103) );
  NAND2_X2 U3891 ( .A1(n3024), .A2(n4497), .ZN(n3823) );
  OAI22_X1 U3892 ( .A1(n3037), .A2(n3025), .B1(n3103), .B2(n3823), .ZN(n3026)
         );
  OR3_X1 U3893 ( .A1(n3028), .A2(n3027), .A3(n3026), .ZN(U3219) );
  OAI22_X1 U3894 ( .A1(n3029), .A2(n3042), .B1(n3140), .B2(n3674), .ZN(n3047)
         );
  OAI22_X1 U3895 ( .A1(n3029), .A2(n3674), .B1(n3140), .B2(n3677), .ZN(n3030)
         );
  XNOR2_X1 U3896 ( .A(n3030), .B(n3639), .ZN(n3048) );
  XOR2_X1 U3897 ( .A(n3047), .B(n3048), .Z(n3036) );
  NAND2_X1 U3898 ( .A1(n3035), .A2(n3036), .ZN(n3050) );
  OAI21_X1 U3899 ( .B1(n3036), .B2(n3035), .A(n3050), .ZN(n3040) );
  OAI22_X1 U3900 ( .A1(n3141), .A2(n3822), .B1(n3810), .B2(n3140), .ZN(n3039)
         );
  INV_X1 U3901 ( .A(REG3_REG_2__SCAN_IN), .ZN(n4009) );
  OAI22_X1 U3902 ( .A1(n3037), .A2(n4009), .B1(n3015), .B2(n3823), .ZN(n3038)
         );
  AOI211_X1 U3903 ( .C1(n3040), .C2(n3820), .A(n3039), .B(n3038), .ZN(n3041)
         );
  INV_X1 U3904 ( .A(n3041), .ZN(U3234) );
  OAI22_X1 U3905 ( .A1(n3141), .A2(n3042), .B1(n3674), .B2(n3117), .ZN(n3085)
         );
  NAND2_X1 U3906 ( .A1(n3043), .A2(n2146), .ZN(n3044) );
  NAND2_X1 U3907 ( .A1(n3045), .A2(n3044), .ZN(n3046) );
  XNOR2_X1 U3908 ( .A(n3046), .B(n3639), .ZN(n3084) );
  XOR2_X1 U3909 ( .A(n3085), .B(n3084), .Z(n3088) );
  OR2_X1 U3910 ( .A1(n3048), .A2(n3047), .ZN(n3049) );
  XOR2_X1 U3911 ( .A(n3088), .B(n3089), .Z(n3060) );
  INV_X1 U3912 ( .A(n3823), .ZN(n3690) );
  OAI22_X1 U3913 ( .A1(n3132), .A2(n3822), .B1(n3810), .B2(n3117), .ZN(n3058)
         );
  NAND2_X1 U3914 ( .A1(n3052), .A2(n3051), .ZN(n3053) );
  OAI21_X1 U3915 ( .B1(n3054), .B2(n3053), .A(STATE_REG_SCAN_IN), .ZN(n3056)
         );
  NAND2_X1 U3916 ( .A1(n3056), .A2(n3055), .ZN(n3813) );
  MUX2_X1 U3917 ( .A(n3813), .B(U3149), .S(REG3_REG_3__SCAN_IN), .Z(n3057) );
  AOI211_X1 U3918 ( .C1(n3690), .C2(n2828), .A(n3058), .B(n3057), .ZN(n3059)
         );
  OAI21_X1 U3919 ( .B1(n3060), .B2(n3815), .A(n3059), .ZN(U3215) );
  AND2_X1 U3920 ( .A1(n3062), .A2(n3061), .ZN(n3065) );
  INV_X1 U3921 ( .A(n2725), .ZN(n3064) );
  OAI21_X1 U3922 ( .B1(n3065), .B2(n3064), .A(n3063), .ZN(n3138) );
  AOI22_X1 U3923 ( .A1(n3529), .A2(n4429), .B1(n3066), .B2(n4427), .ZN(n3067)
         );
  OAI21_X1 U3924 ( .B1(n3015), .B2(n4432), .A(n3067), .ZN(n3072) );
  OAI21_X1 U3925 ( .B1(n2725), .B2(n3069), .A(n3068), .ZN(n3070) );
  AOI22_X1 U3926 ( .A1(n3138), .A2(n3350), .B1(n3070), .B2(n4437), .ZN(n3139)
         );
  INV_X1 U3927 ( .A(n3139), .ZN(n3071) );
  AOI211_X1 U3928 ( .C1(n4645), .C2(n3138), .A(n3072), .B(n3071), .ZN(n3267)
         );
  INV_X1 U3929 ( .A(n4441), .ZN(n3494) );
  XNOR2_X1 U3930 ( .A(n3073), .B(n3140), .ZN(n3265) );
  AOI22_X1 U3931 ( .A1(n3494), .A2(n3265), .B1(REG1_REG_2__SCAN_IN), .B2(n4655), .ZN(n3074) );
  OAI21_X1 U3932 ( .B1(n3267), .B2(n4655), .A(n3074), .ZN(U3520) );
  XOR2_X1 U3933 ( .A(n3075), .B(n3871), .Z(n3112) );
  OAI22_X1 U3934 ( .A1(n3132), .A2(n4361), .B1(n4258), .B2(n3117), .ZN(n3080)
         );
  OAI21_X1 U3935 ( .B1(n3871), .B2(n3077), .A(n3076), .ZN(n3078) );
  AOI22_X1 U3936 ( .A1(n3078), .A2(n4437), .B1(n4357), .B2(n2828), .ZN(n3079)
         );
  INV_X1 U3937 ( .A(n3079), .ZN(n3119) );
  AOI211_X1 U3938 ( .C1(n4423), .C2(n3112), .A(n3080), .B(n3119), .ZN(n3274)
         );
  OR2_X1 U3939 ( .A1(n3081), .A2(n3117), .ZN(n3082) );
  AOI22_X1 U3940 ( .A1(n3272), .A2(n3494), .B1(REG1_REG_3__SCAN_IN), .B2(n4655), .ZN(n3083) );
  OAI21_X1 U3941 ( .B1(n3274), .B2(n4655), .A(n3083), .ZN(U3521) );
  INV_X1 U3942 ( .A(n3084), .ZN(n3087) );
  INV_X1 U3943 ( .A(n3085), .ZN(n3086) );
  NAND2_X1 U3944 ( .A1(n3225), .A2(n3016), .ZN(n3091) );
  NAND2_X1 U3945 ( .A1(n3528), .A2(n3631), .ZN(n3090) );
  NAND2_X1 U3946 ( .A1(n3091), .A2(n3090), .ZN(n3092) );
  XNOR2_X1 U3947 ( .A(n3092), .B(n3639), .ZN(n3125) );
  AOI22_X1 U3948 ( .A1(n3225), .A2(n3636), .B1(n3016), .B2(n3528), .ZN(n3126)
         );
  XNOR2_X1 U3949 ( .A(n3125), .B(n3126), .ZN(n3093) );
  NAND2_X1 U3950 ( .A1(n3094), .A2(n3093), .ZN(n3129) );
  OAI211_X1 U3951 ( .C1(n3094), .C2(n3093), .A(n3129), .B(n3820), .ZN(n3099)
         );
  OAI22_X1 U3952 ( .A1(n3252), .A2(n3822), .B1(n3823), .B2(n3141), .ZN(n3097)
         );
  OAI21_X1 U3953 ( .B1(n3810), .B2(n3536), .A(n3095), .ZN(n3096) );
  NOR2_X1 U3954 ( .A1(n3097), .A2(n3096), .ZN(n3098) );
  OAI211_X1 U3955 ( .C1(n3831), .C2(n3538), .A(n3099), .B(n3098), .ZN(U3227)
         );
  INV_X1 U3956 ( .A(n3100), .ZN(n3106) );
  AOI22_X1 U3957 ( .A1(n2828), .A2(n4429), .B1(n4427), .B2(n3101), .ZN(n3102)
         );
  OAI21_X1 U3958 ( .B1(n3103), .B2(n4432), .A(n3102), .ZN(n3105) );
  AOI211_X1 U3959 ( .C1(n4645), .C2(n3106), .A(n3105), .B(n3104), .ZN(n3279)
         );
  OAI22_X1 U3960 ( .A1(n4441), .A2(n3276), .B1(n4657), .B2(n3107), .ZN(n3108)
         );
  INV_X1 U3961 ( .A(n3108), .ZN(n3109) );
  OAI21_X1 U3962 ( .B1(n3279), .B2(n4655), .A(n3109), .ZN(U3519) );
  NAND2_X1 U3963 ( .A1(n4237), .A2(n3110), .ZN(n3111) );
  INV_X1 U3964 ( .A(n3112), .ZN(n3121) );
  NAND2_X1 U3965 ( .A1(n4611), .A2(n3272), .ZN(n3116) );
  INV_X1 U3966 ( .A(n4625), .ZN(n4606) );
  INV_X1 U3967 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3113) );
  OAI22_X1 U3968 ( .A1(n4606), .A2(n3113), .B1(REG3_REG_3__SCAN_IN), .B2(n4603), .ZN(n3114) );
  AOI21_X1 U3969 ( .B1(n4313), .B2(n3225), .A(n3114), .ZN(n3115) );
  OAI211_X1 U3970 ( .C1(n4319), .C2(n3117), .A(n3116), .B(n3115), .ZN(n3118)
         );
  AOI21_X1 U3971 ( .B1(n3119), .B2(n4238), .A(n3118), .ZN(n3120) );
  OAI21_X1 U3972 ( .B1(n4327), .B2(n3121), .A(n3120), .ZN(U3287) );
  XNOR2_X1 U3973 ( .A(n3123), .B(n3639), .ZN(n3247) );
  NOR2_X1 U3974 ( .A1(n3230), .A2(n3674), .ZN(n3124) );
  AOI21_X1 U3975 ( .B1(n3996), .B2(n3636), .A(n3124), .ZN(n3246) );
  XNOR2_X1 U3976 ( .A(n3247), .B(n3246), .ZN(n3131) );
  OAI211_X1 U3977 ( .C1(n3131), .C2(n3130), .A(n2229), .B(n3820), .ZN(n3137)
         );
  OAI22_X1 U3978 ( .A1(n3132), .A2(n3823), .B1(n3822), .B2(n3301), .ZN(n3135)
         );
  OAI21_X1 U3979 ( .B1(n3810), .B2(n3230), .A(n3133), .ZN(n3134) );
  NOR2_X1 U3980 ( .A1(n3135), .A2(n3134), .ZN(n3136) );
  OAI211_X1 U3981 ( .C1(n3831), .C2(n3226), .A(n3137), .B(n3136), .ZN(U3224)
         );
  INV_X1 U3982 ( .A(n3138), .ZN(n3147) );
  MUX2_X1 U3983 ( .A(n2871), .B(n3139), .S(n4606), .Z(n3146) );
  OAI22_X1 U3984 ( .A1(n4319), .A2(n3140), .B1(n4009), .B2(n4603), .ZN(n3144)
         );
  INV_X1 U3985 ( .A(n4313), .ZN(n3142) );
  OAI22_X1 U3986 ( .A1(n3142), .A2(n3141), .B1(n3015), .B2(n4079), .ZN(n3143)
         );
  AOI211_X1 U3987 ( .C1(n4611), .C2(n3265), .A(n3144), .B(n3143), .ZN(n3145)
         );
  OAI211_X1 U3988 ( .C1(n3147), .C2(n4608), .A(n3146), .B(n3145), .ZN(U3288)
         );
  INV_X1 U3989 ( .A(n4423), .ZN(n4647) );
  INV_X1 U3990 ( .A(n3149), .ZN(n3923) );
  XOR2_X1 U3991 ( .A(n3148), .B(n3893), .Z(n3234) );
  OAI22_X1 U3992 ( .A1(n3301), .A2(n4361), .B1(n4258), .B2(n3230), .ZN(n3152)
         );
  XNOR2_X1 U3993 ( .A(n3150), .B(n3893), .ZN(n3151) );
  NOR2_X1 U3994 ( .A1(n3151), .A2(n4261), .ZN(n3223) );
  AOI211_X1 U3995 ( .C1(n4357), .C2(n3225), .A(n3152), .B(n3223), .ZN(n3153)
         );
  OAI21_X1 U3996 ( .B1(n4647), .B2(n3234), .A(n3153), .ZN(n3268) );
  NAND2_X1 U3997 ( .A1(n3268), .A2(n4657), .ZN(n3157) );
  AND2_X1 U3998 ( .A1(n3535), .A2(n3154), .ZN(n3155) );
  NOR2_X1 U3999 ( .A1(n3196), .A2(n3155), .ZN(n3269) );
  NAND2_X1 U4000 ( .A1(n3269), .A2(n3494), .ZN(n3156) );
  OAI211_X1 U4001 ( .C1(n4657), .C2(n3158), .A(n3157), .B(n3156), .ZN(U3523)
         );
  INV_X1 U4002 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3159) );
  NOR2_X1 U4003 ( .A1(n3188), .A2(n3159), .ZN(n4042) );
  AOI21_X1 U4004 ( .B1(n3159), .B2(n3188), .A(n4042), .ZN(n3168) );
  NAND2_X1 U4005 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3169), .ZN(n3164) );
  INV_X1 U4006 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3408) );
  AOI22_X1 U4007 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3169), .B1(n4637), .B2(
        n3408), .ZN(n4538) );
  INV_X1 U4008 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3238) );
  INV_X1 U4009 ( .A(n3170), .ZN(n4639) );
  AOI22_X1 U4010 ( .A1(n3170), .A2(REG2_REG_9__SCAN_IN), .B1(n3238), .B2(n4639), .ZN(n4518) );
  INV_X1 U4011 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4605) );
  NAND2_X1 U4012 ( .A1(n3176), .A2(n3162), .ZN(n3163) );
  INV_X1 U4013 ( .A(n3176), .ZN(n4638) );
  XNOR2_X1 U4014 ( .A(n3162), .B(n4638), .ZN(n4525) );
  NAND2_X1 U4015 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4525), .ZN(n4524) );
  NAND2_X1 U4016 ( .A1(n3163), .A2(n4524), .ZN(n4537) );
  NAND2_X1 U4017 ( .A1(n4538), .A2(n4537), .ZN(n4536) );
  NAND2_X1 U4018 ( .A1(n3164), .A2(n4536), .ZN(n3165) );
  NAND2_X1 U4019 ( .A1(n4634), .A2(n3165), .ZN(n3166) );
  INV_X1 U4020 ( .A(n4634), .ZN(n4553) );
  XNOR2_X1 U4021 ( .A(n3165), .B(n4553), .ZN(n4545) );
  NAND2_X1 U4022 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4545), .ZN(n4544) );
  OAI21_X1 U4023 ( .B1(n3168), .B2(n4043), .A(n4584), .ZN(n3167) );
  AOI21_X1 U4024 ( .B1(n3168), .B2(n4043), .A(n3167), .ZN(n3190) );
  NAND2_X1 U4025 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3169), .ZN(n3179) );
  AOI22_X1 U4026 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3169), .B1(n4637), .B2(
        n3450), .ZN(n4535) );
  NAND2_X1 U4027 ( .A1(n3170), .A2(REG1_REG_9__SCAN_IN), .ZN(n3175) );
  AOI22_X1 U4028 ( .A1(n3170), .A2(REG1_REG_9__SCAN_IN), .B1(n2538), .B2(n4639), .ZN(n4516) );
  NAND2_X1 U4029 ( .A1(n3176), .A2(n3177), .ZN(n3178) );
  XNOR2_X1 U4030 ( .A(n3177), .B(n4638), .ZN(n4530) );
  NAND2_X1 U4031 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4530), .ZN(n4529) );
  NAND2_X1 U4032 ( .A1(n4634), .A2(n3180), .ZN(n3181) );
  NAND2_X1 U4033 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4550), .ZN(n4549) );
  NAND2_X1 U4034 ( .A1(n3181), .A2(n4549), .ZN(n3184) );
  NOR2_X1 U4035 ( .A1(n3188), .A2(n3182), .ZN(n4025) );
  AOI21_X1 U4036 ( .B1(n3182), .B2(n3188), .A(n4025), .ZN(n3183) );
  NAND2_X1 U4037 ( .A1(n3183), .A2(n3184), .ZN(n4026) );
  OAI211_X1 U4038 ( .C1(n3184), .C2(n3183), .A(n4595), .B(n4026), .ZN(n3187)
         );
  NOR2_X1 U4039 ( .A1(STATE_REG_SCAN_IN), .A2(n3185), .ZN(n3778) );
  AOI21_X1 U4040 ( .B1(n4594), .B2(ADDR_REG_13__SCAN_IN), .A(n3778), .ZN(n3186) );
  OAI211_X1 U4041 ( .C1(n4602), .C2(n3188), .A(n3187), .B(n3186), .ZN(n3189)
         );
  OR2_X1 U4042 ( .A1(n3190), .A2(n3189), .ZN(U3253) );
  XNOR2_X1 U40430 ( .A(n3191), .B(n3875), .ZN(n3205) );
  XOR2_X1 U4044 ( .A(n3875), .B(n3192), .Z(n3208) );
  OAI22_X1 U4045 ( .A1(n3345), .A2(n4361), .B1(n4258), .B2(n3254), .ZN(n3193)
         );
  AOI21_X1 U4046 ( .B1(n4357), .B2(n3996), .A(n3193), .ZN(n3194) );
  OAI21_X1 U4047 ( .B1(n3208), .B2(n4261), .A(n3194), .ZN(n3195) );
  AOI21_X1 U4048 ( .B1(n3205), .B2(n4423), .A(n3195), .ZN(n3264) );
  INV_X1 U4049 ( .A(n3196), .ZN(n3198) );
  INV_X1 U4050 ( .A(n3214), .ZN(n3197) );
  AOI21_X1 U4051 ( .B1(n3200), .B2(n3198), .A(n3197), .ZN(n3262) );
  AOI22_X1 U4052 ( .A1(n3262), .A2(n3494), .B1(n4655), .B2(REG1_REG_6__SCAN_IN), .ZN(n3199) );
  OAI21_X1 U4053 ( .B1(n3264), .B2(n4655), .A(n3199), .ZN(U3524) );
  NOR2_X1 U4054 ( .A1(n4625), .A2(n4261), .ZN(n3465) );
  INV_X1 U4055 ( .A(n3465), .ZN(n3290) );
  AOI22_X1 U4056 ( .A1(n4161), .A2(n3200), .B1(n4313), .B2(n3995), .ZN(n3203)
         );
  INV_X1 U4057 ( .A(n3259), .ZN(n3201) );
  AOI22_X1 U4058 ( .A1(n4625), .A2(REG2_REG_6__SCAN_IN), .B1(n3201), .B2(n4619), .ZN(n3202) );
  OAI211_X1 U4059 ( .C1(n3252), .C2(n4079), .A(n3203), .B(n3202), .ZN(n3204)
         );
  AOI21_X1 U4060 ( .B1(n3262), .B2(n4611), .A(n3204), .ZN(n3207) );
  NAND2_X1 U4061 ( .A1(n3205), .A2(n4296), .ZN(n3206) );
  OAI211_X1 U4062 ( .C1(n3208), .C2(n3290), .A(n3207), .B(n3206), .ZN(U3284)
         );
  XNOR2_X1 U4063 ( .A(n3209), .B(n3874), .ZN(n3212) );
  OAI22_X1 U4064 ( .A1(n3374), .A2(n4361), .B1(n3303), .B2(n4258), .ZN(n3210)
         );
  AOI21_X1 U4065 ( .B1(n4357), .B2(n3224), .A(n3210), .ZN(n3211) );
  OAI21_X1 U4066 ( .B1(n3212), .B2(n4261), .A(n3211), .ZN(n4649) );
  INV_X1 U4067 ( .A(n4649), .ZN(n3222) );
  AOI21_X1 U4068 ( .B1(n3214), .B2(n3296), .A(n3213), .ZN(n3215) );
  AND2_X1 U4069 ( .A1(n3215), .A2(n3339), .ZN(n4650) );
  OAI22_X1 U4070 ( .A1(n4606), .A2(n3216), .B1(n3308), .B2(n4603), .ZN(n3220)
         );
  NOR2_X1 U4071 ( .A1(n3217), .A2(n3874), .ZN(n4648) );
  INV_X1 U4072 ( .A(n4651), .ZN(n3218) );
  NOR3_X1 U4073 ( .A1(n4648), .A2(n3218), .A3(n4327), .ZN(n3219) );
  AOI211_X1 U4074 ( .C1(n4285), .C2(n4650), .A(n3220), .B(n3219), .ZN(n3221)
         );
  OAI21_X1 U4075 ( .B1(n4625), .B2(n3222), .A(n3221), .ZN(U3283) );
  NAND2_X1 U4076 ( .A1(n3223), .A2(n4238), .ZN(n3233) );
  AOI22_X1 U4077 ( .A1(n4314), .A2(n3225), .B1(n4313), .B2(n3224), .ZN(n3229)
         );
  INV_X1 U4078 ( .A(n3226), .ZN(n3227) );
  AOI22_X1 U4079 ( .A1(n4625), .A2(REG2_REG_5__SCAN_IN), .B1(n3227), .B2(n4619), .ZN(n3228) );
  OAI211_X1 U4080 ( .C1(n3230), .C2(n4319), .A(n3229), .B(n3228), .ZN(n3231)
         );
  AOI21_X1 U4081 ( .B1(n3269), .B2(n4611), .A(n3231), .ZN(n3232) );
  OAI211_X1 U4082 ( .C1(n3234), .C2(n4327), .A(n3233), .B(n3232), .ZN(U3285)
         );
  XNOR2_X1 U4083 ( .A(n3235), .B(n3870), .ZN(n3236) );
  NAND2_X1 U4084 ( .A1(n3236), .A2(n4437), .ZN(n3313) );
  NOR2_X1 U4085 ( .A1(n3340), .A2(n3376), .ZN(n3237) );
  INV_X1 U4086 ( .A(n3319), .ZN(n3242) );
  OAI22_X1 U4087 ( .A1(n3381), .A2(n4603), .B1(n3238), .B2(n4606), .ZN(n3241)
         );
  AOI22_X1 U4088 ( .A1(n4161), .A2(n3369), .B1(n4313), .B2(n3992), .ZN(n3239)
         );
  OAI21_X1 U4089 ( .B1(n3374), .B2(n4079), .A(n3239), .ZN(n3240) );
  AOI211_X1 U4090 ( .C1(n3242), .C2(n4611), .A(n3241), .B(n3240), .ZN(n3245)
         );
  XNOR2_X1 U4091 ( .A(n3243), .B(n3870), .ZN(n3309) );
  NAND2_X1 U4092 ( .A1(n3309), .A2(n4296), .ZN(n3244) );
  OAI211_X1 U4093 ( .C1(n3313), .C2(n4625), .A(n3245), .B(n3244), .ZN(U3281)
         );
  INV_X1 U4094 ( .A(n3246), .ZN(n3248) );
  OAI22_X1 U4095 ( .A1(n3301), .A2(n3674), .B1(n3677), .B2(n3254), .ZN(n3249)
         );
  XNOR2_X1 U4096 ( .A(n3249), .B(n3639), .ZN(n3292) );
  INV_X1 U4097 ( .A(n3291), .ZN(n3293) );
  XNOR2_X1 U4098 ( .A(n3292), .B(n3293), .ZN(n3250) );
  XNOR2_X1 U4099 ( .A(n3294), .B(n3250), .ZN(n3251) );
  NAND2_X1 U4100 ( .A1(n3251), .A2(n3820), .ZN(n3258) );
  OAI22_X1 U4101 ( .A1(n3252), .A2(n3823), .B1(n3822), .B2(n3345), .ZN(n3256)
         );
  OAI21_X1 U4102 ( .B1(n3810), .B2(n3254), .A(n3253), .ZN(n3255) );
  NOR2_X1 U4103 ( .A1(n3256), .A2(n3255), .ZN(n3257) );
  OAI211_X1 U4104 ( .C1(n3831), .C2(n3259), .A(n3258), .B(n3257), .ZN(U3236)
         );
  INV_X1 U4105 ( .A(n4495), .ZN(n3498) );
  INV_X1 U4106 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3260) );
  NOR2_X1 U4107 ( .A1(n4475), .A2(n3260), .ZN(n3261) );
  AOI21_X1 U4108 ( .B1(n3262), .B2(n3498), .A(n3261), .ZN(n3263) );
  OAI21_X1 U4109 ( .B1(n3264), .B2(n4653), .A(n3263), .ZN(U3479) );
  AOI22_X1 U4110 ( .A1(n3498), .A2(n3265), .B1(REG0_REG_2__SCAN_IN), .B2(n4653), .ZN(n3266) );
  OAI21_X1 U4111 ( .B1(n3267), .B2(n4653), .A(n3266), .ZN(U3471) );
  INV_X1 U4112 ( .A(n3268), .ZN(n3271) );
  AOI22_X1 U4113 ( .A1(n3269), .A2(n3498), .B1(REG0_REG_5__SCAN_IN), .B2(n4653), .ZN(n3270) );
  OAI21_X1 U4114 ( .B1(n3271), .B2(n4653), .A(n3270), .ZN(U3477) );
  AOI22_X1 U4115 ( .A1(n3272), .A2(n3498), .B1(REG0_REG_3__SCAN_IN), .B2(n4653), .ZN(n3273) );
  OAI21_X1 U4116 ( .B1(n3274), .B2(n4653), .A(n3273), .ZN(U3473) );
  INV_X1 U4117 ( .A(REG0_REG_1__SCAN_IN), .ZN(n3275) );
  OAI22_X1 U4118 ( .A1(n4495), .A2(n3276), .B1(n4475), .B2(n3275), .ZN(n3277)
         );
  INV_X1 U4119 ( .A(n3277), .ZN(n3278) );
  OAI21_X1 U4120 ( .B1(n3279), .B2(n4653), .A(n3278), .ZN(U3469) );
  AND2_X1 U4121 ( .A1(n3943), .A2(n3946), .ZN(n3892) );
  XOR2_X1 U4122 ( .A(n3892), .B(n3280), .Z(n3358) );
  XOR2_X1 U4123 ( .A(n3892), .B(n3281), .Z(n3360) );
  NAND2_X1 U4124 ( .A1(n3360), .A2(n4296), .ZN(n3289) );
  OAI21_X1 U4125 ( .B1(n3282), .B2(n3394), .A(n3409), .ZN(n3365) );
  INV_X1 U4126 ( .A(n3365), .ZN(n3287) );
  AOI22_X1 U4127 ( .A1(n4161), .A2(n3391), .B1(n4313), .B2(n3483), .ZN(n3285)
         );
  INV_X1 U4128 ( .A(n3399), .ZN(n3283) );
  AOI22_X1 U4129 ( .A1(n4625), .A2(REG2_REG_10__SCAN_IN), .B1(n3283), .B2(
        n4619), .ZN(n3284) );
  OAI211_X1 U4130 ( .C1(n2294), .C2(n4079), .A(n3285), .B(n3284), .ZN(n3286)
         );
  AOI21_X1 U4131 ( .B1(n3287), .B2(n4611), .A(n3286), .ZN(n3288) );
  OAI211_X1 U4132 ( .C1(n3358), .C2(n3290), .A(n3289), .B(n3288), .ZN(U3280)
         );
  NAND2_X1 U4133 ( .A1(n3995), .A2(n3016), .ZN(n3298) );
  NAND2_X1 U4134 ( .A1(n3296), .A2(n2146), .ZN(n3297) );
  NAND2_X1 U4135 ( .A1(n3298), .A2(n3297), .ZN(n3299) );
  XNOR2_X1 U4136 ( .A(n3299), .B(n3639), .ZN(n3321) );
  OAI22_X1 U4137 ( .A1(n3345), .A2(n3042), .B1(n3674), .B2(n3303), .ZN(n3320)
         );
  XOR2_X1 U4138 ( .A(n3321), .B(n3320), .Z(n3322) );
  XOR2_X1 U4139 ( .A(n3323), .B(n3322), .Z(n3300) );
  NAND2_X1 U4140 ( .A1(n3300), .A2(n3820), .ZN(n3307) );
  OAI22_X1 U4141 ( .A1(n3374), .A2(n3822), .B1(n3823), .B2(n3301), .ZN(n3305)
         );
  OAI21_X1 U4142 ( .B1(n3810), .B2(n3303), .A(n3302), .ZN(n3304) );
  NOR2_X1 U4143 ( .A1(n3305), .A2(n3304), .ZN(n3306) );
  OAI211_X1 U4144 ( .C1(n3831), .C2(n3308), .A(n3307), .B(n3306), .ZN(U3210)
         );
  NAND2_X1 U4145 ( .A1(n3309), .A2(n4423), .ZN(n3312) );
  AOI22_X1 U4146 ( .A1(n3992), .A2(n4429), .B1(n4427), .B2(n3369), .ZN(n3311)
         );
  NAND2_X1 U4147 ( .A1(n3994), .A2(n4357), .ZN(n3310) );
  NAND4_X1 U4148 ( .A1(n3313), .A2(n3312), .A3(n3311), .A4(n3310), .ZN(n3316)
         );
  MUX2_X1 U4149 ( .A(REG1_REG_9__SCAN_IN), .B(n3316), .S(n4657), .Z(n3314) );
  INV_X1 U4150 ( .A(n3314), .ZN(n3315) );
  OAI21_X1 U4151 ( .B1(n4441), .B2(n3319), .A(n3315), .ZN(U3527) );
  MUX2_X1 U4152 ( .A(REG0_REG_9__SCAN_IN), .B(n3316), .S(n4475), .Z(n3317) );
  INV_X1 U4153 ( .A(n3317), .ZN(n3318) );
  OAI21_X1 U4154 ( .B1(n3319), .B2(n4495), .A(n3318), .ZN(U3485) );
  NAND2_X1 U4155 ( .A1(n3994), .A2(n3016), .ZN(n3326) );
  NAND2_X1 U4156 ( .A1(n3324), .A2(n2146), .ZN(n3325) );
  NAND2_X1 U4157 ( .A1(n3326), .A2(n3325), .ZN(n3327) );
  XNOR2_X1 U4158 ( .A(n3327), .B(n3675), .ZN(n3330) );
  NOR2_X1 U4159 ( .A1(n3344), .A2(n3674), .ZN(n3328) );
  AOI21_X1 U4160 ( .B1(n3994), .B2(n3636), .A(n3328), .ZN(n3329) );
  NOR2_X1 U4161 ( .A1(n3330), .A2(n3329), .ZN(n3367) );
  INV_X1 U4162 ( .A(n3367), .ZN(n3331) );
  NAND2_X1 U4163 ( .A1(n3330), .A2(n3329), .ZN(n3366) );
  NAND2_X1 U4164 ( .A1(n3331), .A2(n3366), .ZN(n3332) );
  XNOR2_X1 U4165 ( .A(n3368), .B(n3332), .ZN(n3333) );
  NAND2_X1 U4166 ( .A1(n3333), .A2(n3820), .ZN(n3338) );
  OAI22_X1 U4167 ( .A1(n3345), .A2(n3823), .B1(n3822), .B2(n2294), .ZN(n3336)
         );
  OAI21_X1 U4168 ( .B1(n3810), .B2(n3344), .A(n3334), .ZN(n3335) );
  NOR2_X1 U4169 ( .A1(n3336), .A2(n3335), .ZN(n3337) );
  OAI211_X1 U4170 ( .C1(n3831), .C2(n4604), .A(n3338), .B(n3337), .ZN(U3218)
         );
  INV_X1 U4171 ( .A(n3339), .ZN(n3341) );
  OAI21_X1 U4172 ( .B1(n3341), .B2(n3344), .A(n2209), .ZN(n4609) );
  AND2_X1 U4173 ( .A1(n2183), .A2(n3930), .ZN(n3873) );
  XNOR2_X1 U4174 ( .A(n3342), .B(n3873), .ZN(n4612) );
  XNOR2_X1 U4175 ( .A(n3343), .B(n3873), .ZN(n3348) );
  OAI22_X1 U4176 ( .A1(n3345), .A2(n4432), .B1(n4258), .B2(n3344), .ZN(n3346)
         );
  AOI21_X1 U4177 ( .B1(n4429), .B2(n3993), .A(n3346), .ZN(n3347) );
  OAI21_X1 U4178 ( .B1(n3348), .B2(n4261), .A(n3347), .ZN(n3349) );
  AOI21_X1 U4179 ( .B1(n3350), .B2(n4612), .A(n3349), .ZN(n4615) );
  INV_X1 U4180 ( .A(n4615), .ZN(n3351) );
  AOI21_X1 U4181 ( .B1(n4645), .B2(n4612), .A(n3351), .ZN(n3353) );
  MUX2_X1 U4182 ( .A(n3174), .B(n3353), .S(n4657), .Z(n3352) );
  OAI21_X1 U4183 ( .B1(n4609), .B2(n4441), .A(n3352), .ZN(U3526) );
  INV_X1 U4184 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3354) );
  MUX2_X1 U4185 ( .A(n3354), .B(n3353), .S(n4475), .Z(n3355) );
  OAI21_X1 U4186 ( .B1(n4609), .B2(n4495), .A(n3355), .ZN(U3483) );
  OAI22_X1 U4187 ( .A1(n3715), .A2(n4361), .B1(n4258), .B2(n3394), .ZN(n3356)
         );
  AOI21_X1 U4188 ( .B1(n4357), .B2(n3993), .A(n3356), .ZN(n3357) );
  OAI21_X1 U4189 ( .B1(n3358), .B2(n4261), .A(n3357), .ZN(n3359) );
  AOI21_X1 U4190 ( .B1(n4423), .B2(n3360), .A(n3359), .ZN(n3362) );
  MUX2_X1 U4191 ( .A(n2549), .B(n3362), .S(n4657), .Z(n3361) );
  OAI21_X1 U4192 ( .B1(n3365), .B2(n4441), .A(n3361), .ZN(U3528) );
  INV_X1 U4193 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3363) );
  MUX2_X1 U4194 ( .A(n3363), .B(n3362), .S(n4475), .Z(n3364) );
  OAI21_X1 U4195 ( .B1(n3365), .B2(n4495), .A(n3364), .ZN(U3487) );
  NAND2_X1 U4196 ( .A1(n3993), .A2(n3016), .ZN(n3371) );
  NAND2_X1 U4197 ( .A1(n3369), .A2(n3631), .ZN(n3370) );
  NAND2_X1 U4198 ( .A1(n3371), .A2(n3370), .ZN(n3372) );
  XNOR2_X1 U4199 ( .A(n3372), .B(n3639), .ZN(n3382) );
  OAI22_X1 U4200 ( .A1(n2294), .A2(n3042), .B1(n3674), .B2(n3376), .ZN(n3383)
         );
  XOR2_X1 U4201 ( .A(n3382), .B(n3383), .Z(n3386) );
  XNOR2_X1 U4202 ( .A(n3387), .B(n3386), .ZN(n3373) );
  NAND2_X1 U4203 ( .A1(n3373), .A2(n3820), .ZN(n3380) );
  OAI22_X1 U4204 ( .A1(n3374), .A2(n3823), .B1(n3822), .B2(n3475), .ZN(n3378)
         );
  AND2_X1 U4205 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4522) );
  INV_X1 U4206 ( .A(n4522), .ZN(n3375) );
  OAI21_X1 U4207 ( .B1(n3810), .B2(n3376), .A(n3375), .ZN(n3377) );
  NOR2_X1 U4208 ( .A1(n3378), .A2(n3377), .ZN(n3379) );
  OAI211_X1 U4209 ( .C1(n3831), .C2(n3381), .A(n3380), .B(n3379), .ZN(U3228)
         );
  INV_X1 U4210 ( .A(n3382), .ZN(n3385) );
  INV_X1 U4211 ( .A(n3383), .ZN(n3384) );
  NAND2_X1 U4212 ( .A1(n3992), .A2(n3016), .ZN(n3389) );
  NAND2_X1 U4213 ( .A1(n3391), .A2(n3631), .ZN(n3388) );
  NAND2_X1 U4214 ( .A1(n3389), .A2(n3388), .ZN(n3390) );
  XNOR2_X1 U4215 ( .A(n3390), .B(n3639), .ZN(n3467) );
  AOI22_X1 U4216 ( .A1(n3992), .A2(n3636), .B1(n3016), .B2(n3391), .ZN(n3468)
         );
  XNOR2_X1 U4217 ( .A(n3467), .B(n3468), .ZN(n3392) );
  OAI211_X1 U4218 ( .C1(n3393), .C2(n3392), .A(n3471), .B(n3820), .ZN(n3398)
         );
  OAI22_X1 U4219 ( .A1(n2294), .A2(n3823), .B1(n3822), .B2(n3715), .ZN(n3396)
         );
  NAND2_X1 U4220 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4526) );
  OAI21_X1 U4221 ( .B1(n3810), .B2(n3394), .A(n4526), .ZN(n3395) );
  NOR2_X1 U4222 ( .A1(n3396), .A2(n3395), .ZN(n3397) );
  OAI211_X1 U4223 ( .C1(n3831), .C2(n3399), .A(n3398), .B(n3397), .ZN(U3214)
         );
  INV_X1 U4224 ( .A(n3400), .ZN(n3401) );
  AOI21_X1 U4225 ( .B1(n3896), .B2(n3402), .A(n3401), .ZN(n3447) );
  AOI22_X1 U4226 ( .A1(n3991), .A2(n4429), .B1(n3403), .B2(n4427), .ZN(n3407)
         );
  XNOR2_X1 U4227 ( .A(n3404), .B(n3896), .ZN(n3405) );
  NAND2_X1 U4228 ( .A1(n3405), .A2(n4437), .ZN(n3406) );
  OAI211_X1 U4229 ( .C1(n3447), .C2(n4237), .A(n3407), .B(n3406), .ZN(n3449)
         );
  NAND2_X1 U4230 ( .A1(n3449), .A2(n4238), .ZN(n3414) );
  OAI22_X1 U4231 ( .A1(n4606), .A2(n3408), .B1(n3482), .B2(n4603), .ZN(n3412)
         );
  INV_X1 U4232 ( .A(n3409), .ZN(n3410) );
  OAI21_X1 U4233 ( .B1(n3410), .B2(n3477), .A(n3417), .ZN(n3455) );
  NOR2_X1 U4234 ( .A1(n3455), .A2(n4266), .ZN(n3411) );
  AOI211_X1 U4235 ( .C1(n4314), .C2(n3992), .A(n3412), .B(n3411), .ZN(n3413)
         );
  OAI211_X1 U4236 ( .C1(n3447), .C2(n4608), .A(n3414), .B(n3413), .ZN(U3279)
         );
  INV_X1 U4237 ( .A(n3429), .ZN(n3416) );
  OR2_X1 U4238 ( .A1(n3416), .A2(n3430), .ZN(n3424) );
  XNOR2_X1 U4239 ( .A(n3415), .B(n3424), .ZN(n3490) );
  AND2_X1 U4240 ( .A1(n3417), .A2(n3552), .ZN(n3418) );
  NOR2_X1 U4241 ( .A1(n3441), .A2(n3418), .ZN(n3499) );
  NAND2_X1 U4242 ( .A1(n3499), .A2(n4611), .ZN(n3423) );
  INV_X1 U4243 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3419) );
  OAI22_X1 U4244 ( .A1(n4606), .A2(n3419), .B1(n3721), .B2(n4603), .ZN(n3420)
         );
  AOI21_X1 U4245 ( .B1(n3552), .B2(n4161), .A(n3420), .ZN(n3422) );
  AOI22_X1 U4246 ( .A1(n4314), .A2(n3483), .B1(n4313), .B2(n3484), .ZN(n3421)
         );
  NAND3_X1 U4247 ( .A1(n3423), .A2(n3422), .A3(n3421), .ZN(n3427) );
  INV_X1 U4248 ( .A(n3424), .ZN(n3894) );
  XNOR2_X1 U4249 ( .A(n3431), .B(n3894), .ZN(n3425) );
  NAND2_X1 U4250 ( .A1(n3425), .A2(n4437), .ZN(n3489) );
  NOR2_X1 U4251 ( .A1(n3489), .A2(n4625), .ZN(n3426) );
  AOI211_X1 U4252 ( .C1(n4296), .C2(n3490), .A(n3427), .B(n3426), .ZN(n3428)
         );
  INV_X1 U4253 ( .A(n3428), .ZN(U3278) );
  OAI21_X1 U4254 ( .B1(n3431), .B2(n3430), .A(n3429), .ZN(n3435) );
  INV_X1 U4255 ( .A(n3432), .ZN(n3434) );
  OR2_X1 U4256 ( .A1(n3434), .A2(n3433), .ZN(n3886) );
  XNOR2_X1 U4257 ( .A(n3435), .B(n3886), .ZN(n3439) );
  NAND2_X1 U4258 ( .A1(n3991), .A2(n4357), .ZN(n3437) );
  NAND2_X1 U4259 ( .A1(n3990), .A2(n4429), .ZN(n3436) );
  OAI211_X1 U4260 ( .C1(n4258), .C2(n3780), .A(n3437), .B(n3436), .ZN(n3438)
         );
  AOI21_X1 U4261 ( .B1(n3439), .B2(n4437), .A(n3438), .ZN(n3503) );
  XNOR2_X1 U4262 ( .A(n3440), .B(n3886), .ZN(n3501) );
  NOR2_X1 U4263 ( .A1(n3441), .A2(n3780), .ZN(n3442) );
  NOR2_X1 U4264 ( .A1(n3509), .A2(n4266), .ZN(n3444) );
  OAI22_X1 U4265 ( .A1(n4606), .A2(n3159), .B1(n3785), .B2(n4603), .ZN(n3443)
         );
  AOI211_X1 U4266 ( .C1(n3501), .C2(n4296), .A(n3444), .B(n3443), .ZN(n3445)
         );
  OAI21_X1 U4267 ( .B1(n4625), .B2(n3503), .A(n3445), .ZN(U3277) );
  OAI22_X1 U4268 ( .A1(n3447), .A2(n3446), .B1(n3475), .B2(n4432), .ZN(n3448)
         );
  NOR2_X1 U4269 ( .A1(n3449), .A2(n3448), .ZN(n3452) );
  MUX2_X1 U4270 ( .A(n3450), .B(n3452), .S(n4657), .Z(n3451) );
  OAI21_X1 U4271 ( .B1(n4441), .B2(n3455), .A(n3451), .ZN(U3529) );
  INV_X1 U4272 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3453) );
  MUX2_X1 U4273 ( .A(n3453), .B(n3452), .S(n4475), .Z(n3454) );
  OAI21_X1 U4274 ( .B1(n3455), .B2(n4495), .A(n3454), .ZN(U3489) );
  INV_X1 U4275 ( .A(n3456), .ZN(n3457) );
  AOI21_X1 U4276 ( .B1(n3897), .B2(n3458), .A(n3457), .ZN(n4434) );
  XNOR2_X1 U4277 ( .A(n3836), .B(n3897), .ZN(n4438) );
  OAI21_X1 U4278 ( .B1(n3459), .B2(n3652), .A(n3514), .ZN(n4496) );
  NOR2_X1 U4279 ( .A1(n4496), .A2(n4266), .ZN(n3464) );
  AOI22_X1 U4280 ( .A1(n4428), .A2(n4161), .B1(n4313), .B2(n4430), .ZN(n3462)
         );
  INV_X1 U4281 ( .A(n3657), .ZN(n3460) );
  AOI22_X1 U4282 ( .A1(n4625), .A2(REG2_REG_14__SCAN_IN), .B1(n3460), .B2(
        n4619), .ZN(n3461) );
  OAI211_X1 U4283 ( .C1(n4433), .C2(n4079), .A(n3462), .B(n3461), .ZN(n3463)
         );
  AOI211_X1 U4284 ( .C1(n4438), .C2(n3465), .A(n3464), .B(n3463), .ZN(n3466)
         );
  OAI21_X1 U4285 ( .B1(n4434), .B2(n4327), .A(n3466), .ZN(U3276) );
  OAI22_X1 U4286 ( .A1(n3715), .A2(n3674), .B1(n3677), .B2(n3477), .ZN(n3472)
         );
  XNOR2_X1 U4287 ( .A(n3472), .B(n3639), .ZN(n3548) );
  OAI22_X1 U4288 ( .A1(n3715), .A2(n3042), .B1(n3674), .B2(n3477), .ZN(n3546)
         );
  XNOR2_X1 U4289 ( .A(n3548), .B(n3546), .ZN(n3473) );
  XNOR2_X1 U4290 ( .A(n3547), .B(n3473), .ZN(n3474) );
  NAND2_X1 U4291 ( .A1(n3474), .A2(n3820), .ZN(n3481) );
  OAI22_X1 U4292 ( .A1(n3777), .A2(n3822), .B1(n3823), .B2(n3475), .ZN(n3479)
         );
  AND2_X1 U4293 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4542) );
  INV_X1 U4294 ( .A(n4542), .ZN(n3476) );
  OAI21_X1 U4295 ( .B1(n3810), .B2(n3477), .A(n3476), .ZN(n3478) );
  NOR2_X1 U4296 ( .A1(n3479), .A2(n3478), .ZN(n3480) );
  OAI211_X1 U4297 ( .C1(n3831), .C2(n3482), .A(n3481), .B(n3480), .ZN(U3233)
         );
  NAND2_X1 U4298 ( .A1(n3483), .A2(n4357), .ZN(n3486) );
  NAND2_X1 U4299 ( .A1(n3484), .A2(n4429), .ZN(n3485) );
  OAI211_X1 U4300 ( .C1(n4258), .C2(n3716), .A(n3486), .B(n3485), .ZN(n3487)
         );
  INV_X1 U4301 ( .A(n3487), .ZN(n3488) );
  AND2_X1 U4302 ( .A1(n3489), .A2(n3488), .ZN(n3492) );
  NAND2_X1 U4303 ( .A1(n3490), .A2(n4423), .ZN(n3491) );
  NAND2_X1 U4304 ( .A1(n3492), .A2(n3491), .ZN(n3496) );
  MUX2_X1 U4305 ( .A(REG1_REG_12__SCAN_IN), .B(n3496), .S(n4657), .Z(n3493) );
  AOI21_X1 U4306 ( .B1(n3494), .B2(n3499), .A(n3493), .ZN(n3495) );
  INV_X1 U4307 ( .A(n3495), .ZN(U3530) );
  MUX2_X1 U4308 ( .A(REG0_REG_12__SCAN_IN), .B(n3496), .S(n4475), .Z(n3497) );
  AOI21_X1 U4309 ( .B1(n3499), .B2(n3498), .A(n3497), .ZN(n3500) );
  INV_X1 U4310 ( .A(n3500), .ZN(U3491) );
  NAND2_X1 U4311 ( .A1(n3501), .A2(n4423), .ZN(n3502) );
  NAND2_X1 U4312 ( .A1(n3503), .A2(n3502), .ZN(n3506) );
  MUX2_X1 U4313 ( .A(REG1_REG_13__SCAN_IN), .B(n3506), .S(n4657), .Z(n3504) );
  INV_X1 U4314 ( .A(n3504), .ZN(n3505) );
  OAI21_X1 U4315 ( .B1(n4441), .B2(n3509), .A(n3505), .ZN(U3531) );
  MUX2_X1 U4316 ( .A(REG0_REG_13__SCAN_IN), .B(n3506), .S(n4475), .Z(n3507) );
  INV_X1 U4317 ( .A(n3507), .ZN(n3508) );
  OAI21_X1 U4318 ( .B1(n3509), .B2(n4495), .A(n3508), .ZN(U3493) );
  AOI21_X1 U4319 ( .B1(n3510), .B2(n3867), .A(n4261), .ZN(n3512) );
  NAND2_X1 U4320 ( .A1(n3512), .A2(n3511), .ZN(n4420) );
  XNOR2_X1 U4321 ( .A(n3513), .B(n3867), .ZN(n4424) );
  NAND2_X1 U4322 ( .A1(n4424), .A2(n4296), .ZN(n3522) );
  INV_X1 U4323 ( .A(n3514), .ZN(n3515) );
  OAI21_X1 U4324 ( .B1(n3515), .B2(n3825), .A(n4312), .ZN(n4492) );
  INV_X1 U4325 ( .A(n4492), .ZN(n3520) );
  AOI22_X1 U4326 ( .A1(n4314), .A2(n3990), .B1(n4313), .B2(n4418), .ZN(n3518)
         );
  INV_X1 U4327 ( .A(n3830), .ZN(n3516) );
  AOI22_X1 U4328 ( .A1(n4625), .A2(REG2_REG_15__SCAN_IN), .B1(n3516), .B2(
        n4619), .ZN(n3517) );
  OAI211_X1 U4329 ( .C1(n3825), .C2(n4319), .A(n3518), .B(n3517), .ZN(n3519)
         );
  AOI21_X1 U4330 ( .B1(n3520), .B2(n4611), .A(n3519), .ZN(n3521) );
  OAI211_X1 U4331 ( .C1(n4625), .C2(n4420), .A(n3522), .B(n3521), .ZN(U3275)
         );
  INV_X1 U4332 ( .A(n3525), .ZN(n3895) );
  NAND2_X1 U4333 ( .A1(n3524), .A2(n3895), .ZN(n3526) );
  NAND2_X1 U4334 ( .A1(n3523), .A2(n3526), .ZN(n4641) );
  XNOR2_X1 U4335 ( .A(n3895), .B(n3527), .ZN(n3533) );
  AOI22_X1 U4336 ( .A1(n3529), .A2(n4357), .B1(n3528), .B2(n4427), .ZN(n3531)
         );
  NAND2_X1 U4337 ( .A1(n3996), .A2(n4429), .ZN(n3530) );
  OAI211_X1 U4338 ( .C1(n4641), .C2(n4237), .A(n3531), .B(n3530), .ZN(n3532)
         );
  AOI21_X1 U4339 ( .B1(n3533), .B2(n4437), .A(n3532), .ZN(n3534) );
  INV_X1 U4340 ( .A(n3534), .ZN(n4643) );
  OAI211_X1 U4341 ( .C1(n3537), .C2(n3536), .A(n4412), .B(n3535), .ZN(n4642)
         );
  OAI22_X1 U4342 ( .A1(n4642), .A2(n3539), .B1(n4603), .B2(n3538), .ZN(n3540)
         );
  OAI21_X1 U4343 ( .B1(n4643), .B2(n3540), .A(n4606), .ZN(n3542) );
  NAND2_X1 U4344 ( .A1(n4625), .A2(REG2_REG_4__SCAN_IN), .ZN(n3541) );
  OAI211_X1 U4345 ( .C1(n4641), .C2(n4608), .A(n3542), .B(n3541), .ZN(U3286)
         );
  OAI21_X1 U4346 ( .B1(n4441), .B2(n4096), .A(n3544), .ZN(U3546) );
  OAI22_X1 U4347 ( .A1(n4433), .A2(n3674), .B1(n3677), .B2(n3780), .ZN(n3545)
         );
  XNOR2_X1 U4348 ( .A(n3545), .B(n3639), .ZN(n3774) );
  NAND2_X1 U4349 ( .A1(n3991), .A2(n3016), .ZN(n3550) );
  NAND2_X1 U4350 ( .A1(n3552), .A2(n2146), .ZN(n3549) );
  NAND2_X1 U4351 ( .A1(n3550), .A2(n3549), .ZN(n3551) );
  XNOR2_X1 U4352 ( .A(n3551), .B(n3675), .ZN(n3554) );
  AOI22_X1 U4353 ( .A1(n3991), .A2(n3636), .B1(n3016), .B2(n3552), .ZN(n3553)
         );
  OR2_X1 U4354 ( .A1(n3554), .A2(n3553), .ZN(n3710) );
  AND2_X1 U4355 ( .A1(n3554), .A2(n3553), .ZN(n3711) );
  OAI22_X1 U4356 ( .A1(n4433), .A2(n3042), .B1(n3674), .B2(n3780), .ZN(n3773)
         );
  NAND2_X1 U4357 ( .A1(n3990), .A2(n3016), .ZN(n3558) );
  NAND2_X1 U4358 ( .A1(n4428), .A2(n2146), .ZN(n3557) );
  NAND2_X1 U4359 ( .A1(n3558), .A2(n3557), .ZN(n3559) );
  XNOR2_X1 U4360 ( .A(n3559), .B(n3675), .ZN(n3561) );
  AOI22_X1 U4361 ( .A1(n3990), .A2(n3636), .B1(n3016), .B2(n4428), .ZN(n3560)
         );
  NOR2_X1 U4362 ( .A1(n3561), .A2(n3560), .ZN(n3647) );
  NAND2_X1 U4363 ( .A1(n3561), .A2(n3560), .ZN(n3648) );
  OAI22_X1 U4364 ( .A1(n4410), .A2(n3674), .B1(n3825), .B2(n3677), .ZN(n3562)
         );
  XOR2_X1 U4365 ( .A(n3639), .B(n3562), .Z(n3566) );
  NAND2_X1 U4366 ( .A1(n4430), .A2(n3636), .ZN(n3564) );
  NAND2_X1 U4367 ( .A1(n4417), .A2(n3016), .ZN(n3563) );
  NAND2_X1 U4368 ( .A1(n3564), .A2(n3563), .ZN(n3818) );
  INV_X1 U4369 ( .A(n3566), .ZN(n3567) );
  OAI22_X1 U4370 ( .A1(n4402), .A2(n3042), .B1(n4320), .B2(n3674), .ZN(n3572)
         );
  NAND2_X1 U4371 ( .A1(n4418), .A2(n3016), .ZN(n3569) );
  NAND2_X1 U4372 ( .A1(n4407), .A2(n2146), .ZN(n3568) );
  NAND2_X1 U4373 ( .A1(n3569), .A2(n3568), .ZN(n3570) );
  XNOR2_X1 U4374 ( .A(n3570), .B(n3639), .ZN(n3571) );
  XOR2_X1 U4375 ( .A(n3572), .B(n3571), .Z(n3733) );
  INV_X1 U4376 ( .A(n3571), .ZN(n3574) );
  INV_X1 U4377 ( .A(n3572), .ZN(n3573) );
  NAND2_X1 U4378 ( .A1(n4408), .A2(n3016), .ZN(n3576) );
  NAND2_X1 U4379 ( .A1(n4398), .A2(n3631), .ZN(n3575) );
  NAND2_X1 U4380 ( .A1(n3576), .A2(n3575), .ZN(n3577) );
  XNOR2_X1 U4381 ( .A(n3577), .B(n3675), .ZN(n3742) );
  NOR2_X1 U4382 ( .A1(n4304), .A2(n3674), .ZN(n3578) );
  AOI21_X1 U4383 ( .B1(n4408), .B2(n3636), .A(n3578), .ZN(n3741) );
  NAND2_X1 U4384 ( .A1(n3742), .A2(n3741), .ZN(n3579) );
  NAND2_X1 U4385 ( .A1(n4399), .A2(n3016), .ZN(n3581) );
  NAND2_X1 U4386 ( .A1(n4274), .A2(n3631), .ZN(n3580) );
  NAND2_X1 U4387 ( .A1(n3581), .A2(n3580), .ZN(n3582) );
  XNOR2_X1 U4388 ( .A(n3582), .B(n3675), .ZN(n3584) );
  AOI22_X1 U4389 ( .A1(n4399), .A2(n3636), .B1(n3016), .B2(n4274), .ZN(n3583)
         );
  OR2_X1 U4390 ( .A1(n3584), .A2(n3583), .ZN(n3796) );
  NAND2_X1 U4391 ( .A1(n3584), .A2(n3583), .ZN(n3795) );
  OAI22_X1 U4392 ( .A1(n4233), .A2(n3042), .B1(n3674), .B2(n4257), .ZN(n3589)
         );
  NAND2_X1 U4393 ( .A1(n4275), .A2(n3016), .ZN(n3586) );
  NAND2_X1 U4394 ( .A1(n4263), .A2(n3631), .ZN(n3585) );
  NAND2_X1 U4395 ( .A1(n3586), .A2(n3585), .ZN(n3587) );
  XNOR2_X1 U4396 ( .A(n3587), .B(n3639), .ZN(n3588) );
  XOR2_X1 U4397 ( .A(n3589), .B(n3588), .Z(n3668) );
  INV_X1 U4398 ( .A(n3588), .ZN(n3591) );
  INV_X1 U4399 ( .A(n3589), .ZN(n3590) );
  NAND2_X1 U4400 ( .A1(n3593), .A2(n3592), .ZN(n3762) );
  NAND2_X1 U4401 ( .A1(n4214), .A2(n3016), .ZN(n3595) );
  NAND2_X1 U4402 ( .A1(n4230), .A2(n2146), .ZN(n3594) );
  NAND2_X1 U4403 ( .A1(n3595), .A2(n3594), .ZN(n3596) );
  XNOR2_X1 U4404 ( .A(n3596), .B(n3675), .ZN(n3598) );
  AOI22_X1 U4405 ( .A1(n4214), .A2(n3636), .B1(n3016), .B2(n4230), .ZN(n3597)
         );
  OR2_X1 U4406 ( .A1(n3598), .A2(n3597), .ZN(n3763) );
  NAND2_X1 U4407 ( .A1(n3762), .A2(n3763), .ZN(n3761) );
  NAND2_X1 U4408 ( .A1(n3598), .A2(n3597), .ZN(n3764) );
  NAND2_X1 U4409 ( .A1(n4231), .A2(n3016), .ZN(n3600) );
  NAND2_X1 U4410 ( .A1(n4377), .A2(n3631), .ZN(n3599) );
  NAND2_X1 U4411 ( .A1(n3600), .A2(n3599), .ZN(n3601) );
  XNOR2_X1 U4412 ( .A(n3601), .B(n3639), .ZN(n3700) );
  NAND2_X1 U4413 ( .A1(n4231), .A2(n3636), .ZN(n3603) );
  NAND2_X1 U4414 ( .A1(n4377), .A2(n3016), .ZN(n3602) );
  NAND2_X1 U4415 ( .A1(n3603), .A2(n3602), .ZN(n3701) );
  NOR2_X1 U4416 ( .A1(n3700), .A2(n3701), .ZN(n3605) );
  NAND2_X1 U4417 ( .A1(n3700), .A2(n3701), .ZN(n3604) );
  OAI22_X1 U4418 ( .A1(n4175), .A2(n3674), .B1(n4198), .B2(n3677), .ZN(n3606)
         );
  XNOR2_X1 U4419 ( .A(n3606), .B(n3639), .ZN(n3611) );
  OAI22_X1 U4420 ( .A1(n4175), .A2(n3042), .B1(n4198), .B2(n3674), .ZN(n3610)
         );
  XNOR2_X1 U4421 ( .A(n3611), .B(n3610), .ZN(n3787) );
  NOR2_X1 U4422 ( .A1(n4181), .A2(n3674), .ZN(n3608) );
  AOI21_X1 U4423 ( .B1(n4358), .B2(n3636), .A(n3608), .ZN(n3613) );
  OAI22_X1 U4424 ( .A1(n3789), .A2(n3674), .B1(n3677), .B2(n4181), .ZN(n3609)
         );
  XNOR2_X1 U4425 ( .A(n3609), .B(n3639), .ZN(n3612) );
  XOR2_X1 U4426 ( .A(n3613), .B(n3612), .Z(n3658) );
  NOR2_X1 U4427 ( .A1(n3611), .A2(n3610), .ZN(n3659) );
  INV_X1 U4428 ( .A(n3612), .ZN(n3614) );
  NOR2_X1 U4429 ( .A1(n4157), .A2(n3674), .ZN(n3615) );
  AOI21_X1 U4430 ( .B1(n4177), .B2(n3636), .A(n3615), .ZN(n3619) );
  OAI22_X1 U4431 ( .A1(n4139), .A2(n3674), .B1(n3677), .B2(n4157), .ZN(n3618)
         );
  XNOR2_X1 U4432 ( .A(n3618), .B(n3639), .ZN(n3754) );
  NAND2_X1 U4433 ( .A1(n3751), .A2(n3754), .ZN(n3621) );
  NAND2_X1 U4434 ( .A1(n3620), .A2(n3616), .ZN(n3752) );
  NAND2_X1 U4435 ( .A1(n4162), .A2(n3016), .ZN(n3624) );
  NAND2_X1 U4436 ( .A1(n3622), .A2(n2146), .ZN(n3623) );
  NAND2_X1 U4437 ( .A1(n3624), .A2(n3623), .ZN(n3625) );
  XNOR2_X1 U4438 ( .A(n3625), .B(n3675), .ZN(n3627) );
  NOR2_X1 U4439 ( .A1(n4145), .A2(n3674), .ZN(n3626) );
  AOI21_X1 U4440 ( .B1(n4162), .B2(n3636), .A(n3626), .ZN(n3628) );
  NAND2_X1 U4441 ( .A1(n3627), .A2(n3628), .ZN(n3722) );
  INV_X1 U4442 ( .A(n3627), .ZN(n3630) );
  INV_X1 U4443 ( .A(n3628), .ZN(n3629) );
  NAND2_X1 U4444 ( .A1(n3630), .A2(n3629), .ZN(n3723) );
  NAND2_X1 U4445 ( .A1(n4336), .A2(n3016), .ZN(n3633) );
  NAND2_X1 U4446 ( .A1(n4344), .A2(n3631), .ZN(n3632) );
  NAND2_X1 U4447 ( .A1(n3633), .A2(n3632), .ZN(n3634) );
  XNOR2_X1 U4448 ( .A(n3634), .B(n3675), .ZN(n3638) );
  NOR2_X1 U4449 ( .A1(n4129), .A2(n3674), .ZN(n3635) );
  AOI21_X1 U4450 ( .B1(n4336), .B2(n3636), .A(n3635), .ZN(n3637) );
  NOR2_X1 U4451 ( .A1(n3638), .A2(n3637), .ZN(n3806) );
  NAND2_X1 U4452 ( .A1(n3638), .A2(n3637), .ZN(n3804) );
  OAI22_X1 U4453 ( .A1(n3906), .A2(n3674), .B1(n3677), .B2(n4112), .ZN(n3640)
         );
  XNOR2_X1 U4454 ( .A(n3640), .B(n3639), .ZN(n3685) );
  OAI22_X1 U4455 ( .A1(n3906), .A2(n3042), .B1(n3674), .B2(n4112), .ZN(n3684)
         );
  XNOR2_X1 U4456 ( .A(n3685), .B(n3684), .ZN(n3682) );
  XNOR2_X1 U4457 ( .A(n3683), .B(n3682), .ZN(n3645) );
  INV_X1 U4458 ( .A(n3641), .ZN(n4109) );
  OAI22_X1 U4459 ( .A1(n3810), .A2(n4112), .B1(STATE_REG_SCAN_IN), .B2(n4672), 
        .ZN(n3643) );
  OAI22_X1 U4460 ( .A1(n4338), .A2(n3822), .B1(n3726), .B2(n3823), .ZN(n3642)
         );
  AOI211_X1 U4461 ( .C1(n4109), .C2(n3813), .A(n3643), .B(n3642), .ZN(n3644)
         );
  OAI21_X1 U4462 ( .B1(n3645), .B2(n3815), .A(n3644), .ZN(U3211) );
  INV_X1 U4463 ( .A(n3647), .ZN(n3649) );
  NAND2_X1 U4464 ( .A1(n3649), .A2(n3648), .ZN(n3650) );
  XNOR2_X1 U4465 ( .A(n3646), .B(n3650), .ZN(n3651) );
  NAND2_X1 U4466 ( .A1(n3651), .A2(n3820), .ZN(n3656) );
  OAI22_X1 U4467 ( .A1(n4410), .A2(n3822), .B1(n3823), .B2(n4433), .ZN(n3654)
         );
  NAND2_X1 U4468 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4554) );
  OAI21_X1 U4469 ( .B1(n3810), .B2(n3652), .A(n4554), .ZN(n3653) );
  NOR2_X1 U4470 ( .A1(n3654), .A2(n3653), .ZN(n3655) );
  OAI211_X1 U4471 ( .C1(n3831), .C2(n3657), .A(n3656), .B(n3655), .ZN(U3212)
         );
  OAI21_X1 U4472 ( .B1(n2156), .B2(n3659), .A(n3658), .ZN(n3661) );
  NAND3_X1 U4473 ( .A1(n3661), .A2(n3820), .A3(n3660), .ZN(n3666) );
  NAND2_X1 U4474 ( .A1(n3689), .A2(n4177), .ZN(n3662) );
  OAI21_X1 U4475 ( .B1(n4175), .B2(n3823), .A(n3662), .ZN(n3664) );
  INV_X1 U4476 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4890) );
  OAI22_X1 U4477 ( .A1(n3810), .A2(n4181), .B1(STATE_REG_SCAN_IN), .B2(n4890), 
        .ZN(n3663) );
  NOR2_X1 U4478 ( .A1(n3664), .A2(n3663), .ZN(n3665) );
  OAI211_X1 U4479 ( .C1(n3831), .C2(n4183), .A(n3666), .B(n3665), .ZN(U3213)
         );
  XNOR2_X1 U4480 ( .A(n3667), .B(n3668), .ZN(n3669) );
  NAND2_X1 U4481 ( .A1(n3669), .A2(n3820), .ZN(n3673) );
  INV_X1 U4482 ( .A(n4214), .ZN(n4381) );
  OAI22_X1 U4483 ( .A1(n3745), .A2(n3823), .B1(n3822), .B2(n4381), .ZN(n3671)
         );
  NAND2_X1 U4484 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4064) );
  OAI21_X1 U4485 ( .B1(n3810), .B2(n4257), .A(n4064), .ZN(n3670) );
  NOR2_X1 U4486 ( .A1(n3671), .A2(n3670), .ZN(n3672) );
  OAI211_X1 U4487 ( .C1(n3831), .C2(n4267), .A(n3673), .B(n3672), .ZN(U3216)
         );
  OAI22_X1 U4488 ( .A1(n4338), .A2(n3042), .B1(n3678), .B2(n3674), .ZN(n3676)
         );
  XNOR2_X1 U4489 ( .A(n3676), .B(n3675), .ZN(n3680) );
  OAI22_X1 U4490 ( .A1(n4338), .A2(n3674), .B1(n3678), .B2(n3677), .ZN(n3679)
         );
  XNOR2_X1 U4491 ( .A(n3680), .B(n3679), .ZN(n3688) );
  INV_X1 U4492 ( .A(n3688), .ZN(n3681) );
  NAND2_X1 U4493 ( .A1(n3681), .A2(n3820), .ZN(n3699) );
  NAND2_X1 U4494 ( .A1(n3685), .A2(n3684), .ZN(n3687) );
  NAND2_X1 U4495 ( .A1(n3698), .A2(n3686), .ZN(n3697) );
  NOR3_X1 U4496 ( .A1(n3688), .A2(n3687), .A3(n3815), .ZN(n3695) );
  AOI22_X1 U4497 ( .A1(n4345), .A2(n3690), .B1(n3689), .B2(n4093), .ZN(n3693)
         );
  AOI22_X1 U4498 ( .A1(n3691), .A2(n4092), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3692) );
  OAI211_X1 U4499 ( .C1(n3831), .C2(n4090), .A(n3693), .B(n3692), .ZN(n3694)
         );
  NOR2_X1 U4500 ( .A1(n3695), .A2(n3694), .ZN(n3696) );
  OAI211_X1 U4501 ( .C1(n3699), .C2(n3698), .A(n3697), .B(n3696), .ZN(U3217)
         );
  XOR2_X1 U4502 ( .A(n3701), .B(n3700), .Z(n3702) );
  XNOR2_X1 U4503 ( .A(n3703), .B(n3702), .ZN(n3704) );
  NAND2_X1 U4504 ( .A1(n3704), .A2(n3820), .ZN(n3709) );
  OAI22_X1 U4505 ( .A1(n4175), .A2(n3822), .B1(n3823), .B2(n4381), .ZN(n3707)
         );
  OAI22_X1 U4506 ( .A1(n3810), .A2(n4219), .B1(STATE_REG_SCAN_IN), .B2(n3705), 
        .ZN(n3706) );
  NOR2_X1 U4507 ( .A1(n3707), .A2(n3706), .ZN(n3708) );
  OAI211_X1 U4508 ( .C1(n3831), .C2(n4215), .A(n3709), .B(n3708), .ZN(U3220)
         );
  INV_X1 U4509 ( .A(n3710), .ZN(n3712) );
  NOR2_X1 U4510 ( .A1(n3712), .A2(n3711), .ZN(n3713) );
  XNOR2_X1 U4511 ( .A(n2193), .B(n3713), .ZN(n3714) );
  NAND2_X1 U4512 ( .A1(n3714), .A2(n3820), .ZN(n3720) );
  OAI22_X1 U4513 ( .A1(n3715), .A2(n3823), .B1(n3822), .B2(n4433), .ZN(n3718)
         );
  NAND2_X1 U4514 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4546) );
  OAI21_X1 U4515 ( .B1(n3810), .B2(n3716), .A(n4546), .ZN(n3717) );
  NOR2_X1 U4516 ( .A1(n3718), .A2(n3717), .ZN(n3719) );
  OAI211_X1 U4517 ( .C1(n3831), .C2(n3721), .A(n3720), .B(n3719), .ZN(U3221)
         );
  NAND2_X1 U4518 ( .A1(n3723), .A2(n3722), .ZN(n3725) );
  XOR2_X1 U4519 ( .A(n3725), .B(n3724), .Z(n3730) );
  OAI22_X1 U4520 ( .A1(n3810), .A2(n4145), .B1(STATE_REG_SCAN_IN), .B2(n4680), 
        .ZN(n3728) );
  OAI22_X1 U4521 ( .A1(n3726), .A2(n3822), .B1(n4139), .B2(n3823), .ZN(n3727)
         );
  AOI211_X1 U4522 ( .C1(n4146), .C2(n3813), .A(n3728), .B(n3727), .ZN(n3729)
         );
  OAI21_X1 U4523 ( .B1(n3730), .B2(n3815), .A(n3729), .ZN(U3222) );
  INV_X1 U4524 ( .A(n3817), .ZN(n3732) );
  OAI21_X1 U4525 ( .B1(n3732), .B2(n3818), .A(n3731), .ZN(n3734) );
  XNOR2_X1 U4526 ( .A(n3734), .B(n3733), .ZN(n3735) );
  NAND2_X1 U4527 ( .A1(n3735), .A2(n3820), .ZN(n3739) );
  OAI22_X1 U4528 ( .A1(n4277), .A2(n3822), .B1(n3823), .B2(n4410), .ZN(n3737)
         );
  NAND2_X1 U4529 ( .A1(REG3_REG_16__SCAN_IN), .A2(U3149), .ZN(n4585) );
  OAI21_X1 U4530 ( .B1(n3810), .B2(n4320), .A(n4585), .ZN(n3736) );
  NOR2_X1 U4531 ( .A1(n3737), .A2(n3736), .ZN(n3738) );
  OAI211_X1 U4532 ( .C1(n3831), .C2(n4315), .A(n3739), .B(n3738), .ZN(U3223)
         );
  XNOR2_X1 U4533 ( .A(n3742), .B(n3741), .ZN(n3743) );
  XNOR2_X1 U4534 ( .A(n3740), .B(n3743), .ZN(n3744) );
  NAND2_X1 U4535 ( .A1(n3744), .A2(n3820), .ZN(n3750) );
  OAI22_X1 U4536 ( .A1(n4402), .A2(n3823), .B1(n3822), .B2(n3745), .ZN(n3748)
         );
  AND2_X1 U4537 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4593) );
  INV_X1 U4538 ( .A(n4593), .ZN(n3746) );
  OAI21_X1 U4539 ( .B1(n3810), .B2(n4304), .A(n3746), .ZN(n3747) );
  NOR2_X1 U4540 ( .A1(n3748), .A2(n3747), .ZN(n3749) );
  OAI211_X1 U4541 ( .C1(n3831), .C2(n4300), .A(n3750), .B(n3749), .ZN(U3225)
         );
  NAND2_X1 U4542 ( .A1(n3752), .A2(n3751), .ZN(n3753) );
  XOR2_X1 U4543 ( .A(n3754), .B(n3753), .Z(n3760) );
  INV_X1 U4544 ( .A(n4159), .ZN(n3758) );
  OAI22_X1 U4545 ( .A1(n3810), .A2(n4157), .B1(STATE_REG_SCAN_IN), .B2(n3755), 
        .ZN(n3757) );
  OAI22_X1 U4546 ( .A1(n4362), .A2(n3822), .B1(n3789), .B2(n3823), .ZN(n3756)
         );
  AOI211_X1 U4547 ( .C1(n3758), .C2(n3813), .A(n3757), .B(n3756), .ZN(n3759)
         );
  OAI21_X1 U4548 ( .B1(n3760), .B2(n3815), .A(n3759), .ZN(U3226) );
  NOR2_X1 U4549 ( .A1(n3761), .A2(n2363), .ZN(n3766) );
  AOI21_X1 U4550 ( .B1(n3764), .B2(n3763), .A(n3762), .ZN(n3765) );
  OAI21_X1 U4551 ( .B1(n3766), .B2(n3765), .A(n3820), .ZN(n3771) );
  OAI22_X1 U4552 ( .A1(n4233), .A2(n3823), .B1(n3822), .B2(n3788), .ZN(n3769)
         );
  OAI22_X1 U4553 ( .A1(n3810), .A2(n4241), .B1(STATE_REG_SCAN_IN), .B2(n3767), 
        .ZN(n3768) );
  NOR2_X1 U4554 ( .A1(n3769), .A2(n3768), .ZN(n3770) );
  OAI211_X1 U4555 ( .C1(n3831), .C2(n4243), .A(n3771), .B(n3770), .ZN(U3230)
         );
  XNOR2_X1 U4556 ( .A(n3774), .B(n3773), .ZN(n3775) );
  XNOR2_X1 U4557 ( .A(n3772), .B(n3775), .ZN(n3776) );
  NAND2_X1 U4558 ( .A1(n3776), .A2(n3820), .ZN(n3784) );
  OAI22_X1 U4559 ( .A1(n3777), .A2(n3823), .B1(n3822), .B2(n4421), .ZN(n3782)
         );
  INV_X1 U4560 ( .A(n3778), .ZN(n3779) );
  OAI21_X1 U4561 ( .B1(n3810), .B2(n3780), .A(n3779), .ZN(n3781) );
  NOR2_X1 U4562 ( .A1(n3782), .A2(n3781), .ZN(n3783) );
  OAI211_X1 U4563 ( .C1(n3831), .C2(n3785), .A(n3784), .B(n3783), .ZN(U3231)
         );
  AOI21_X1 U4564 ( .B1(n3787), .B2(n3786), .A(n2156), .ZN(n3794) );
  INV_X1 U4565 ( .A(n4201), .ZN(n3792) );
  INV_X1 U4566 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4863) );
  OAI22_X1 U4567 ( .A1(n3810), .A2(n4198), .B1(STATE_REG_SCAN_IN), .B2(n4863), 
        .ZN(n3791) );
  OAI22_X1 U4568 ( .A1(n3789), .A2(n3822), .B1(n3823), .B2(n3788), .ZN(n3790)
         );
  AOI211_X1 U4569 ( .C1(n3792), .C2(n3813), .A(n3791), .B(n3790), .ZN(n3793)
         );
  OAI21_X1 U4570 ( .B1(n3794), .B2(n3815), .A(n3793), .ZN(U3232) );
  NAND2_X1 U4571 ( .A1(n3796), .A2(n3795), .ZN(n3797) );
  XOR2_X1 U4572 ( .A(n3797), .B(n2158), .Z(n3798) );
  NAND2_X1 U4573 ( .A1(n3798), .A2(n3820), .ZN(n3803) );
  OAI22_X1 U4574 ( .A1(n4233), .A2(n3822), .B1(n3823), .B2(n4277), .ZN(n3801)
         );
  NOR2_X1 U4575 ( .A1(STATE_REG_SCAN_IN), .A2(n4862), .ZN(n4035) );
  INV_X1 U4576 ( .A(n4035), .ZN(n3799) );
  OAI21_X1 U4577 ( .B1(n3810), .B2(n4284), .A(n3799), .ZN(n3800) );
  NOR2_X1 U4578 ( .A1(n3801), .A2(n3800), .ZN(n3802) );
  OAI211_X1 U4579 ( .C1(n3831), .C2(n4287), .A(n3803), .B(n3802), .ZN(U3235)
         );
  INV_X1 U4580 ( .A(n3804), .ZN(n3805) );
  NOR2_X1 U4581 ( .A1(n3806), .A2(n3805), .ZN(n3807) );
  XNOR2_X1 U4582 ( .A(n3808), .B(n3807), .ZN(n3816) );
  OAI22_X1 U4583 ( .A1(n3810), .A2(n4129), .B1(STATE_REG_SCAN_IN), .B2(n3809), 
        .ZN(n3812) );
  OAI22_X1 U4584 ( .A1(n3906), .A2(n3822), .B1(n4362), .B2(n3823), .ZN(n3811)
         );
  AOI211_X1 U4585 ( .C1(n4126), .C2(n3813), .A(n3812), .B(n3811), .ZN(n3814)
         );
  OAI21_X1 U4586 ( .B1(n3816), .B2(n3815), .A(n3814), .ZN(U3237) );
  NAND2_X1 U4587 ( .A1(n3817), .A2(n3731), .ZN(n3819) );
  XNOR2_X1 U4588 ( .A(n3819), .B(n3818), .ZN(n3821) );
  NAND2_X1 U4589 ( .A1(n3821), .A2(n3820), .ZN(n3829) );
  OAI22_X1 U4590 ( .A1(n4421), .A2(n3823), .B1(n3822), .B2(n4402), .ZN(n3827)
         );
  INV_X1 U4591 ( .A(REG3_REG_15__SCAN_IN), .ZN(n4843) );
  NOR2_X1 U4592 ( .A1(STATE_REG_SCAN_IN), .A2(n4843), .ZN(n4568) );
  INV_X1 U4593 ( .A(n4568), .ZN(n3824) );
  OAI21_X1 U4594 ( .B1(n3810), .B2(n3825), .A(n3824), .ZN(n3826) );
  NOR2_X1 U4595 ( .A1(n3827), .A2(n3826), .ZN(n3828) );
  OAI211_X1 U4596 ( .C1(n3831), .C2(n3830), .A(n3829), .B(n3828), .ZN(U3238)
         );
  NAND2_X1 U4597 ( .A1(n3832), .A2(n3835), .ZN(n3907) );
  NAND2_X1 U4598 ( .A1(n3834), .A2(n3833), .ZN(n3933) );
  NAND2_X1 U4599 ( .A1(n3933), .A2(n3835), .ZN(n3954) );
  OAI21_X1 U4600 ( .B1(n3836), .B2(n3907), .A(n3954), .ZN(n3841) );
  NOR2_X1 U4601 ( .A1(n3838), .A2(n3887), .ZN(n3840) );
  NAND2_X1 U4602 ( .A1(n3840), .A2(n3839), .ZN(n3957) );
  AOI211_X1 U4603 ( .C1(n3841), .C2(n3955), .A(n2308), .B(n3957), .ZN(n3844)
         );
  INV_X1 U4604 ( .A(n3842), .ZN(n3958) );
  NOR3_X1 U4605 ( .A1(n3844), .A2(n3958), .A3(n3843), .ZN(n3847) );
  INV_X1 U4606 ( .A(n3866), .ZN(n3845) );
  NOR2_X1 U4607 ( .A1(n3882), .A2(n3845), .ZN(n3964) );
  OAI21_X1 U4608 ( .B1(n3847), .B2(n3846), .A(n3964), .ZN(n3851) );
  OR2_X1 U4609 ( .A1(n3849), .A2(n3848), .ZN(n3856) );
  NAND2_X1 U4610 ( .A1(n3861), .A2(n4333), .ZN(n3850) );
  NAND2_X1 U4611 ( .A1(n2151), .A2(DATAI_31_), .ZN(n4070) );
  NAND2_X1 U4612 ( .A1(n3883), .A2(n4070), .ZN(n3974) );
  AND2_X1 U4613 ( .A1(n3850), .A2(n3974), .ZN(n3890) );
  OAI21_X1 U4614 ( .B1(n4093), .B2(n4077), .A(n3890), .ZN(n3855) );
  AOI211_X1 U4615 ( .C1(n4117), .C2(n3851), .A(n3856), .B(n3855), .ZN(n3859)
         );
  INV_X1 U4616 ( .A(n3966), .ZN(n3858) );
  NAND2_X1 U4617 ( .A1(n4093), .A2(n4077), .ZN(n3852) );
  AND2_X1 U4618 ( .A1(n3853), .A2(n3852), .ZN(n3969) );
  NAND3_X1 U4619 ( .A1(n3879), .A2(n3969), .A3(n3854), .ZN(n3857) );
  AOI21_X1 U4620 ( .B1(n3969), .B2(n3856), .A(n3855), .ZN(n3976) );
  AOI22_X1 U4621 ( .A1(n3859), .A2(n3858), .B1(n3857), .B2(n3976), .ZN(n3860)
         );
  AOI21_X1 U4622 ( .B1(n4072), .B2(n4333), .A(n3860), .ZN(n3864) );
  OR2_X1 U4623 ( .A1(n3861), .A2(n4333), .ZN(n3885) );
  AOI21_X1 U4624 ( .B1(n3885), .B2(n3883), .A(n4070), .ZN(n3863) );
  NOR3_X1 U4625 ( .A1(n3864), .A2(n3863), .A3(n3862), .ZN(n3982) );
  XNOR2_X1 U4626 ( .A(n4214), .B(n4230), .ZN(n4228) );
  NAND2_X1 U4627 ( .A1(n3866), .A2(n3865), .ZN(n4173) );
  INV_X1 U4628 ( .A(n3963), .ZN(n4171) );
  NAND2_X1 U4629 ( .A1(n4171), .A2(n4169), .ZN(n4211) );
  NOR4_X1 U4630 ( .A1(n4173), .A2(n4211), .A3(n4621), .A4(n3867), .ZN(n3868)
         );
  NAND3_X1 U4631 ( .A1(n2799), .A2(n4228), .A3(n3868), .ZN(n3878) );
  NAND2_X1 U4632 ( .A1(n4118), .A2(n3869), .ZN(n4138) );
  NAND4_X1 U4633 ( .A1(n3873), .A2(n3872), .A3(n3871), .A4(n3870), .ZN(n3877)
         );
  INV_X1 U4634 ( .A(n4189), .ZN(n4196) );
  INV_X1 U4635 ( .A(n3874), .ZN(n3927) );
  NAND4_X1 U4636 ( .A1(n4196), .A2(n4322), .A3(n3927), .A4(n3875), .ZN(n3876)
         );
  NOR4_X1 U4637 ( .A1(n3878), .A2(n4138), .A3(n3877), .A4(n3876), .ZN(n3880)
         );
  NAND2_X1 U4638 ( .A1(n3880), .A2(n3879), .ZN(n3905) );
  XNOR2_X1 U4639 ( .A(n4336), .B(n4129), .ZN(n4123) );
  INV_X1 U4640 ( .A(n4135), .ZN(n3881) );
  NOR2_X1 U4641 ( .A1(n3882), .A2(n3881), .ZN(n4152) );
  OR2_X1 U4642 ( .A1(n3883), .A2(n4070), .ZN(n3884) );
  NAND2_X1 U4643 ( .A1(n3885), .A2(n3884), .ZN(n3975) );
  NOR2_X1 U4644 ( .A1(n3975), .A2(n4501), .ZN(n3902) );
  INV_X1 U4645 ( .A(n3886), .ZN(n3891) );
  AND2_X1 U4646 ( .A1(n2305), .A2(n4250), .ZN(n4294) );
  AND4_X1 U4647 ( .A1(n3891), .A2(n4294), .A3(n4255), .A4(n3890), .ZN(n3901)
         );
  INV_X1 U4648 ( .A(n4281), .ZN(n4272) );
  NAND4_X1 U4649 ( .A1(n3894), .A2(n4272), .A3(n3893), .A4(n3892), .ZN(n3899)
         );
  NAND4_X1 U4650 ( .A1(n3897), .A2(n3896), .A3(n3895), .A4(n2725), .ZN(n3898)
         );
  NOR2_X1 U4651 ( .A1(n3899), .A2(n3898), .ZN(n3900) );
  NAND4_X1 U4652 ( .A1(n4152), .A2(n3902), .A3(n3901), .A4(n3900), .ZN(n3903)
         );
  NOR4_X1 U4653 ( .A1(n3905), .A2(n3904), .A3(n4123), .A4(n3903), .ZN(n3980)
         );
  NOR2_X1 U4654 ( .A1(n3906), .A2(n4335), .ZN(n3973) );
  INV_X1 U4655 ( .A(n3948), .ZN(n3910) );
  INV_X1 U4656 ( .A(n3907), .ZN(n3908) );
  OAI211_X1 U4657 ( .C1(n3911), .C2(n3910), .A(n3909), .B(n3908), .ZN(n3953)
         );
  OAI211_X1 U4658 ( .C1(n3914), .C2(n4501), .A(n3913), .B(n3912), .ZN(n3916)
         );
  NAND3_X1 U4659 ( .A1(n3916), .A2(n2726), .A3(n3915), .ZN(n3919) );
  NAND3_X1 U4660 ( .A1(n3919), .A2(n3918), .A3(n3917), .ZN(n3922) );
  NAND3_X1 U4661 ( .A1(n3922), .A2(n3921), .A3(n3920), .ZN(n3925) );
  NAND4_X1 U4662 ( .A1(n3925), .A2(n3924), .A3(n3923), .A4(n3938), .ZN(n3928)
         );
  NAND3_X1 U4663 ( .A1(n3928), .A2(n3927), .A3(n3926), .ZN(n3929) );
  NAND3_X1 U4664 ( .A1(n3929), .A2(n3937), .A3(n2183), .ZN(n3932) );
  NAND3_X1 U4665 ( .A1(n3932), .A2(n3931), .A3(n3930), .ZN(n3935) );
  INV_X1 U4666 ( .A(n3933), .ZN(n3934) );
  NAND3_X1 U4667 ( .A1(n3935), .A2(n3934), .A3(n3936), .ZN(n3951) );
  NAND2_X1 U4668 ( .A1(n2183), .A2(n3936), .ZN(n3942) );
  INV_X1 U4669 ( .A(n3937), .ZN(n3941) );
  INV_X1 U4670 ( .A(n3938), .ZN(n3940) );
  NOR4_X1 U4671 ( .A1(n3942), .A2(n3941), .A3(n3940), .A4(n3939), .ZN(n3945)
         );
  INV_X1 U4672 ( .A(n3943), .ZN(n3944) );
  OAI21_X1 U4673 ( .B1(n3945), .B2(n3944), .A(n3954), .ZN(n3950) );
  NAND3_X1 U4674 ( .A1(n3948), .A2(n3947), .A3(n3946), .ZN(n3949) );
  AOI21_X1 U4675 ( .B1(n3951), .B2(n3950), .A(n3949), .ZN(n3952) );
  AOI21_X1 U4676 ( .B1(n3954), .B2(n3953), .A(n3952), .ZN(n3956) );
  OAI21_X1 U4677 ( .B1(n3956), .B2(n2308), .A(n3955), .ZN(n3960) );
  INV_X1 U4678 ( .A(n3957), .ZN(n3959) );
  AOI21_X1 U4679 ( .B1(n3960), .B2(n3959), .A(n3958), .ZN(n3962) );
  OAI21_X1 U4680 ( .B1(n3963), .B2(n3962), .A(n3961), .ZN(n3967) );
  INV_X1 U4681 ( .A(n3964), .ZN(n3965) );
  AOI211_X1 U4682 ( .C1(n3968), .C2(n3967), .A(n3966), .B(n3965), .ZN(n3972)
         );
  INV_X1 U4683 ( .A(n3969), .ZN(n3970) );
  OR4_X1 U4684 ( .A1(n3973), .A2(n3972), .A3(n3971), .A4(n3970), .ZN(n3977) );
  AOI22_X1 U4685 ( .A1(n3977), .A2(n3976), .B1(n3975), .B2(n3974), .ZN(n3979)
         );
  MUX2_X1 U4686 ( .A(n3980), .B(n3979), .S(n3978), .Z(n3981) );
  NOR2_X1 U4687 ( .A1(n3982), .A2(n3981), .ZN(n3983) );
  XNOR2_X1 U4688 ( .A(n3983), .B(n4065), .ZN(n3989) );
  NAND2_X1 U4689 ( .A1(n3985), .A2(n3984), .ZN(n3986) );
  OAI211_X1 U4690 ( .C1(n4500), .C2(n3988), .A(n3986), .B(B_REG_SCAN_IN), .ZN(
        n3987) );
  OAI21_X1 U4691 ( .B1(n3989), .B2(n3988), .A(n3987), .ZN(U3239) );
  MUX2_X1 U4692 ( .A(DATAO_REG_29__SCAN_IN), .B(n4093), .S(n3997), .Z(U3579)
         );
  MUX2_X1 U4693 ( .A(DATAO_REG_28__SCAN_IN), .B(n4108), .S(n3997), .Z(U3578)
         );
  MUX2_X1 U4694 ( .A(DATAO_REG_23__SCAN_IN), .B(n4358), .S(n3997), .Z(U3573)
         );
  MUX2_X1 U4695 ( .A(DATAO_REG_21__SCAN_IN), .B(n4231), .S(n3997), .Z(U3571)
         );
  MUX2_X1 U4696 ( .A(DATAO_REG_17__SCAN_IN), .B(n4408), .S(n3997), .Z(U3567)
         );
  MUX2_X1 U4697 ( .A(DATAO_REG_16__SCAN_IN), .B(n4418), .S(n3997), .Z(U3566)
         );
  MUX2_X1 U4698 ( .A(DATAO_REG_14__SCAN_IN), .B(n3990), .S(n3997), .Z(U3564)
         );
  MUX2_X1 U4699 ( .A(DATAO_REG_12__SCAN_IN), .B(n3991), .S(n3997), .Z(U3562)
         );
  MUX2_X1 U4700 ( .A(DATAO_REG_10__SCAN_IN), .B(n3992), .S(n3997), .Z(U3560)
         );
  MUX2_X1 U4701 ( .A(DATAO_REG_9__SCAN_IN), .B(n3993), .S(n3997), .Z(U3559) );
  MUX2_X1 U4702 ( .A(DATAO_REG_8__SCAN_IN), .B(n3994), .S(n3997), .Z(U3558) );
  MUX2_X1 U4703 ( .A(DATAO_REG_7__SCAN_IN), .B(n3995), .S(n3997), .Z(U3557) );
  MUX2_X1 U4704 ( .A(DATAO_REG_5__SCAN_IN), .B(n3996), .S(n3997), .Z(U3555) );
  MUX2_X1 U4705 ( .A(DATAO_REG_1__SCAN_IN), .B(n3017), .S(n3997), .Z(U3551) );
  MUX2_X1 U4706 ( .A(DATAO_REG_0__SCAN_IN), .B(n3998), .S(n3997), .Z(U3550) );
  OAI211_X1 U4707 ( .C1(n4001), .C2(n4000), .A(n4595), .B(n3999), .ZN(n4008)
         );
  MUX2_X1 U4708 ( .A(n4002), .B(REG2_REG_1__SCAN_IN), .S(n4510), .Z(n4003) );
  OAI21_X1 U4709 ( .B1(n4623), .B2(n2367), .A(n4003), .ZN(n4004) );
  NAND3_X1 U4710 ( .A1(n4584), .A2(n4014), .A3(n4004), .ZN(n4007) );
  NAND2_X1 U4711 ( .A1(n4036), .A2(n4510), .ZN(n4006) );
  AOI22_X1 U4712 ( .A1(n4594), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4005) );
  NAND4_X1 U4713 ( .A1(n4008), .A2(n4007), .A3(n4006), .A4(n4005), .ZN(U3241)
         );
  INV_X1 U4714 ( .A(ADDR_REG_2__SCAN_IN), .ZN(n4010) );
  OAI22_X1 U4715 ( .A1(n4587), .A2(n4010), .B1(STATE_REG_SCAN_IN), .B2(n4009), 
        .ZN(n4011) );
  AOI21_X1 U4716 ( .B1(n4509), .B2(n4036), .A(n4011), .ZN(n4023) );
  INV_X1 U4717 ( .A(n4012), .ZN(n4017) );
  NAND3_X1 U4718 ( .A1(n4015), .A2(n4014), .A3(n4013), .ZN(n4016) );
  NAND3_X1 U4719 ( .A1(n4584), .A2(n4017), .A3(n4016), .ZN(n4022) );
  OAI211_X1 U4720 ( .C1(n4020), .C2(n4019), .A(n4595), .B(n4018), .ZN(n4021)
         );
  NAND4_X1 U4721 ( .A1(n4024), .A2(n4023), .A3(n4022), .A4(n4021), .ZN(U3242)
         );
  NOR2_X1 U4722 ( .A1(n4629), .A2(REG1_REG_17__SCAN_IN), .ZN(n4034) );
  NAND2_X1 U4723 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4047), .ZN(n4030) );
  INV_X1 U4724 ( .A(n4047), .ZN(n4631) );
  AOI22_X1 U4725 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4047), .B1(n4631), .B2(
        n4425), .ZN(n4571) );
  INV_X1 U4726 ( .A(n4025), .ZN(n4027) );
  NAND2_X1 U4727 ( .A1(n4027), .A2(n4026), .ZN(n4028) );
  NAND2_X1 U4728 ( .A1(n4632), .A2(n4028), .ZN(n4029) );
  XNOR2_X1 U4729 ( .A(n4028), .B(n2269), .ZN(n4561) );
  NAND2_X1 U4730 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4561), .ZN(n4560) );
  NAND2_X1 U4731 ( .A1(n4029), .A2(n4560), .ZN(n4570) );
  NAND2_X1 U4732 ( .A1(n4571), .A2(n4570), .ZN(n4569) );
  NAND2_X1 U4733 ( .A1(n4030), .A2(n4569), .ZN(n4031) );
  NOR2_X1 U4734 ( .A1(n4031), .A2(n4049), .ZN(n4033) );
  AOI21_X1 U4735 ( .B1(n4031), .B2(n4049), .A(n4033), .ZN(n4032) );
  INV_X1 U4736 ( .A(n4032), .ZN(n4578) );
  AOI22_X1 U4737 ( .A1(n4629), .A2(n4405), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4601), .ZN(n4596) );
  XOR2_X1 U4738 ( .A(REG1_REG_18__SCAN_IN), .B(n4059), .Z(n4060) );
  XNOR2_X1 U4739 ( .A(n2171), .B(n4060), .ZN(n4039) );
  AOI21_X1 U4740 ( .B1(n4594), .B2(ADDR_REG_18__SCAN_IN), .A(n4035), .ZN(n4038) );
  NAND2_X1 U4741 ( .A1(n4036), .A2(n4059), .ZN(n4037) );
  OAI211_X1 U4742 ( .C1(n4039), .C2(n4580), .A(n4038), .B(n4037), .ZN(n4055)
         );
  INV_X1 U4743 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4901) );
  NOR2_X1 U4744 ( .A1(n4059), .A2(n4901), .ZN(n4040) );
  AOI21_X1 U4745 ( .B1(n4059), .B2(n4901), .A(n4040), .ZN(n4053) );
  NOR2_X1 U4746 ( .A1(n4629), .A2(REG2_REG_17__SCAN_IN), .ZN(n4041) );
  AOI21_X1 U4747 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4629), .A(n4041), .ZN(n4591) );
  NOR2_X1 U4748 ( .A1(n2269), .A2(n4044), .ZN(n4045) );
  INV_X1 U4749 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4557) );
  NAND2_X1 U4750 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4047), .ZN(n4046) );
  OAI21_X1 U4751 ( .B1(REG2_REG_15__SCAN_IN), .B2(n4047), .A(n4046), .ZN(n4565) );
  NOR2_X1 U4752 ( .A1(n4566), .A2(n4565), .ZN(n4564) );
  AND2_X1 U4753 ( .A1(n4047), .A2(REG2_REG_15__SCAN_IN), .ZN(n4048) );
  NOR2_X1 U4754 ( .A1(n4564), .A2(n4048), .ZN(n4050) );
  INV_X1 U4755 ( .A(n4049), .ZN(n4579) );
  NAND2_X1 U4756 ( .A1(n4050), .A2(n4579), .ZN(n4051) );
  XNOR2_X1 U4757 ( .A(n4050), .B(n4049), .ZN(n4576) );
  INV_X1 U4758 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4575) );
  NAND2_X1 U4759 ( .A1(n4576), .A2(n4575), .ZN(n4574) );
  NAND2_X1 U4760 ( .A1(n4051), .A2(n4574), .ZN(n4589) );
  NAND2_X1 U4761 ( .A1(n4591), .A2(n4589), .ZN(n4590) );
  OAI21_X1 U4762 ( .B1(n4629), .B2(REG2_REG_17__SCAN_IN), .A(n4590), .ZN(n4052) );
  NOR2_X1 U4763 ( .A1(n4052), .A2(n4053), .ZN(n4056) );
  AOI211_X1 U4764 ( .C1(n4053), .C2(n4052), .A(n4056), .B(n4588), .ZN(n4054)
         );
  OR2_X1 U4765 ( .A1(n4055), .A2(n4054), .ZN(U3258) );
  INV_X1 U4766 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4910) );
  MUX2_X1 U4767 ( .A(n4910), .B(REG2_REG_19__SCAN_IN), .S(n4065), .Z(n4058) );
  AOI21_X1 U4768 ( .B1(n4059), .B2(REG2_REG_18__SCAN_IN), .A(n4056), .ZN(n4057) );
  XOR2_X1 U4769 ( .A(n4058), .B(n4057), .Z(n4069) );
  MUX2_X1 U4770 ( .A(REG1_REG_19__SCAN_IN), .B(n4392), .S(n4065), .Z(n4062) );
  XOR2_X1 U4771 ( .A(n4062), .B(n4061), .Z(n4067) );
  NAND2_X1 U4772 ( .A1(n4594), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4063) );
  OAI211_X1 U4773 ( .C1(n4602), .C2(n4065), .A(n4064), .B(n4063), .ZN(n4066)
         );
  AOI21_X1 U4774 ( .B1(n4067), .B2(n4595), .A(n4066), .ZN(n4068) );
  OAI21_X1 U4775 ( .B1(n4069), .B2(n4588), .A(n4068), .ZN(U3259) );
  XNOR2_X1 U4776 ( .A(n4330), .B(n4070), .ZN(n4445) );
  INV_X1 U4777 ( .A(n4070), .ZN(n4073) );
  NOR2_X1 U4778 ( .A1(n4072), .A2(n4071), .ZN(n4332) );
  AOI21_X1 U4779 ( .B1(n4073), .B2(n4427), .A(n4332), .ZN(n4442) );
  NOR2_X1 U4780 ( .A1(n4442), .A2(n4625), .ZN(n4074) );
  AOI21_X1 U4781 ( .B1(REG2_REG_31__SCAN_IN), .B2(n4625), .A(n4074), .ZN(n4075) );
  OAI21_X1 U4782 ( .B1(n4445), .B2(n4266), .A(n4075), .ZN(U3260) );
  INV_X1 U4783 ( .A(n4076), .ZN(n4086) );
  INV_X1 U4784 ( .A(n4077), .ZN(n4081) );
  INV_X1 U4785 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4078) );
  OAI22_X1 U4786 ( .A1(n4338), .A2(n4079), .B1(n4078), .B2(n4238), .ZN(n4080)
         );
  AOI21_X1 U4787 ( .B1(n4081), .B2(n4161), .A(n4080), .ZN(n4085) );
  INV_X1 U4788 ( .A(n4087), .ZN(n4100) );
  INV_X1 U4789 ( .A(n4088), .ZN(n4098) );
  INV_X1 U4790 ( .A(REG2_REG_28__SCAN_IN), .ZN(n4089) );
  OAI22_X1 U4791 ( .A1(n4090), .A2(n4603), .B1(n4089), .B2(n4238), .ZN(n4091)
         );
  AOI21_X1 U4792 ( .B1(n4092), .B2(n4161), .A(n4091), .ZN(n4095) );
  AOI22_X1 U4793 ( .A1(n4345), .A2(n4314), .B1(n4313), .B2(n4093), .ZN(n4094)
         );
  OAI211_X1 U4794 ( .C1(n4096), .C2(n4266), .A(n4095), .B(n4094), .ZN(n4097)
         );
  AOI21_X1 U4795 ( .B1(n4098), .B2(n4238), .A(n4097), .ZN(n4099) );
  OAI21_X1 U4796 ( .B1(n4100), .B2(n4327), .A(n4099), .ZN(U3262) );
  XNOR2_X1 U4797 ( .A(n4101), .B(n4102), .ZN(n4341) );
  INV_X1 U4798 ( .A(n4341), .ZN(n4116) );
  NAND2_X1 U4799 ( .A1(n4103), .A2(n4102), .ZN(n4104) );
  AOI21_X1 U4800 ( .B1(n4105), .B2(n4104), .A(n4261), .ZN(n4340) );
  INV_X1 U4801 ( .A(n4125), .ZN(n4107) );
  OAI21_X1 U4802 ( .B1(n4107), .B2(n4112), .A(n4106), .ZN(n4452) );
  NOR2_X1 U4803 ( .A1(n4452), .A2(n4266), .ZN(n4114) );
  AOI22_X1 U4804 ( .A1(n4108), .A2(n4313), .B1(n4314), .B2(n4336), .ZN(n4111)
         );
  AOI22_X1 U4805 ( .A1(n4109), .A2(n4619), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4625), .ZN(n4110) );
  OAI211_X1 U4806 ( .C1(n4112), .C2(n4319), .A(n4111), .B(n4110), .ZN(n4113)
         );
  AOI211_X1 U4807 ( .C1(n4340), .C2(n4606), .A(n4114), .B(n4113), .ZN(n4115)
         );
  OAI21_X1 U4808 ( .B1(n4116), .B2(n4327), .A(n4115), .ZN(U3263) );
  NAND2_X1 U4809 ( .A1(n4136), .A2(n4117), .ZN(n4119) );
  NAND2_X1 U4810 ( .A1(n4119), .A2(n4118), .ZN(n4121) );
  INV_X1 U4811 ( .A(n4123), .ZN(n4120) );
  XNOR2_X1 U4812 ( .A(n4121), .B(n4120), .ZN(n4122) );
  NAND2_X1 U4813 ( .A1(n4122), .A2(n4437), .ZN(n4347) );
  XNOR2_X1 U4814 ( .A(n4124), .B(n4123), .ZN(n4349) );
  NAND2_X1 U4815 ( .A1(n4349), .A2(n4296), .ZN(n4133) );
  OAI21_X1 U4816 ( .B1(n4143), .B2(n4129), .A(n4125), .ZN(n4455) );
  INV_X1 U4817 ( .A(n4455), .ZN(n4131) );
  AOI22_X1 U4818 ( .A1(n4345), .A2(n4313), .B1(n4314), .B2(n4162), .ZN(n4128)
         );
  AOI22_X1 U4819 ( .A1(n4126), .A2(n4619), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4625), .ZN(n4127) );
  OAI211_X1 U4820 ( .C1(n4129), .C2(n4319), .A(n4128), .B(n4127), .ZN(n4130)
         );
  AOI21_X1 U4821 ( .B1(n4131), .B2(n4611), .A(n4130), .ZN(n4132) );
  OAI211_X1 U4822 ( .C1(n4625), .C2(n4347), .A(n4133), .B(n4132), .ZN(U3264)
         );
  XNOR2_X1 U4823 ( .A(n4134), .B(n4138), .ZN(n4353) );
  INV_X1 U4824 ( .A(n4353), .ZN(n4150) );
  NAND2_X1 U4825 ( .A1(n4136), .A2(n4135), .ZN(n4137) );
  XOR2_X1 U4826 ( .A(n4138), .B(n4137), .Z(n4142) );
  OAI22_X1 U4827 ( .A1(n4139), .A2(n4432), .B1(n4145), .B2(n4258), .ZN(n4140)
         );
  AOI21_X1 U4828 ( .B1(n4429), .B2(n4336), .A(n4140), .ZN(n4141) );
  OAI21_X1 U4829 ( .B1(n4142), .B2(n4261), .A(n4141), .ZN(n4352) );
  INV_X1 U4830 ( .A(n4143), .ZN(n4144) );
  OAI21_X1 U4831 ( .B1(n4155), .B2(n4145), .A(n4144), .ZN(n4459) );
  AOI22_X1 U4832 ( .A1(n4146), .A2(n4619), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4625), .ZN(n4147) );
  OAI21_X1 U4833 ( .B1(n4459), .B2(n4266), .A(n4147), .ZN(n4148) );
  AOI21_X1 U4834 ( .B1(n4352), .B2(n4238), .A(n4148), .ZN(n4149) );
  OAI21_X1 U4835 ( .B1(n4150), .B2(n4327), .A(n4149), .ZN(U3265) );
  XOR2_X1 U4836 ( .A(n4152), .B(n4151), .Z(n4364) );
  XNOR2_X1 U4837 ( .A(n4153), .B(n4152), .ZN(n4154) );
  NAND2_X1 U4838 ( .A1(n4154), .A2(n4437), .ZN(n4360) );
  NOR2_X1 U4839 ( .A1(n4360), .A2(n4625), .ZN(n4166) );
  INV_X1 U4840 ( .A(n4155), .ZN(n4156) );
  OAI21_X1 U4841 ( .B1(n2211), .B2(n4157), .A(n4156), .ZN(n4462) );
  OAI22_X1 U4842 ( .A1(n4159), .A2(n4603), .B1(n4158), .B2(n4238), .ZN(n4160)
         );
  AOI21_X1 U4843 ( .B1(n4356), .B2(n4161), .A(n4160), .ZN(n4164) );
  AOI22_X1 U4844 ( .A1(n4162), .A2(n4313), .B1(n4314), .B2(n4358), .ZN(n4163)
         );
  OAI211_X1 U4845 ( .C1(n4462), .C2(n4266), .A(n4164), .B(n4163), .ZN(n4165)
         );
  AOI211_X1 U4846 ( .C1(n4364), .C2(n4296), .A(n4166), .B(n4165), .ZN(n4167)
         );
  INV_X1 U4847 ( .A(n4167), .ZN(U3266) );
  XOR2_X1 U4848 ( .A(n4173), .B(n4168), .Z(n4368) );
  INV_X1 U4849 ( .A(n4368), .ZN(n4188) );
  INV_X1 U4850 ( .A(n4169), .ZN(n4170) );
  AOI21_X1 U4851 ( .B1(n4208), .B2(n4171), .A(n4170), .ZN(n4190) );
  OAI21_X1 U4852 ( .B1(n4190), .B2(n4189), .A(n4172), .ZN(n4174) );
  XNOR2_X1 U4853 ( .A(n4174), .B(n4173), .ZN(n4179) );
  OAI22_X1 U4854 ( .A1(n4175), .A2(n4432), .B1(n4258), .B2(n4181), .ZN(n4176)
         );
  AOI21_X1 U4855 ( .B1(n4429), .B2(n4177), .A(n4176), .ZN(n4178) );
  OAI21_X1 U4856 ( .B1(n4179), .B2(n4261), .A(n4178), .ZN(n4367) );
  INV_X1 U4857 ( .A(n4200), .ZN(n4182) );
  OAI21_X1 U4858 ( .B1(n4182), .B2(n4181), .A(n4180), .ZN(n4466) );
  NOR2_X1 U4859 ( .A1(n4466), .A2(n4266), .ZN(n4186) );
  INV_X1 U4860 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4184) );
  OAI22_X1 U4861 ( .A1(n4184), .A2(n4238), .B1(n4183), .B2(n4603), .ZN(n4185)
         );
  AOI211_X1 U4862 ( .C1(n4367), .C2(n4606), .A(n4186), .B(n4185), .ZN(n4187)
         );
  OAI21_X1 U4863 ( .B1(n4188), .B2(n4327), .A(n4187), .ZN(U3267) );
  XNOR2_X1 U4864 ( .A(n4190), .B(n4189), .ZN(n4194) );
  NAND2_X1 U4865 ( .A1(n4358), .A2(n4429), .ZN(n4192) );
  NAND2_X1 U4866 ( .A1(n4231), .A2(n4357), .ZN(n4191) );
  OAI211_X1 U4867 ( .C1(n4258), .C2(n4198), .A(n4192), .B(n4191), .ZN(n4193)
         );
  AOI21_X1 U4868 ( .B1(n4194), .B2(n4437), .A(n4193), .ZN(n4373) );
  INV_X1 U4869 ( .A(n4195), .ZN(n4197) );
  NAND2_X1 U4870 ( .A1(n4197), .A2(n4196), .ZN(n4372) );
  NAND3_X1 U4871 ( .A1(n4372), .A2(n4296), .A3(n4371), .ZN(n4206) );
  OR2_X1 U4872 ( .A1(n4212), .A2(n4198), .ZN(n4199) );
  NAND2_X1 U4873 ( .A1(n4200), .A2(n4199), .ZN(n4470) );
  INV_X1 U4874 ( .A(n4470), .ZN(n4204) );
  INV_X1 U4875 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4202) );
  OAI22_X1 U4876 ( .A1(n4606), .A2(n4202), .B1(n4201), .B2(n4603), .ZN(n4203)
         );
  AOI21_X1 U4877 ( .B1(n4204), .B2(n4611), .A(n4203), .ZN(n4205) );
  OAI211_X1 U4878 ( .C1(n4625), .C2(n4373), .A(n4206), .B(n4205), .ZN(U3268)
         );
  INV_X1 U4879 ( .A(n4211), .ZN(n4207) );
  XNOR2_X1 U4880 ( .A(n4208), .B(n4207), .ZN(n4209) );
  NAND2_X1 U4881 ( .A1(n4209), .A2(n4437), .ZN(n4380) );
  XOR2_X1 U4882 ( .A(n4211), .B(n4210), .Z(n4383) );
  NAND2_X1 U4883 ( .A1(n4383), .A2(n4296), .ZN(n4223) );
  INV_X1 U4884 ( .A(n4212), .ZN(n4213) );
  OAI21_X1 U4885 ( .B1(n4239), .B2(n4219), .A(n4213), .ZN(n4474) );
  INV_X1 U4886 ( .A(n4474), .ZN(n4221) );
  AOI22_X1 U4887 ( .A1(n4314), .A2(n4214), .B1(n4378), .B2(n4313), .ZN(n4218)
         );
  INV_X1 U4888 ( .A(n4215), .ZN(n4216) );
  AOI22_X1 U4889 ( .A1(n4625), .A2(REG2_REG_21__SCAN_IN), .B1(n4216), .B2(
        n4619), .ZN(n4217) );
  OAI211_X1 U4890 ( .C1(n4219), .C2(n4319), .A(n4218), .B(n4217), .ZN(n4220)
         );
  AOI21_X1 U4891 ( .B1(n4221), .B2(n4611), .A(n4220), .ZN(n4222) );
  OAI211_X1 U4892 ( .C1(n4625), .C2(n4380), .A(n4223), .B(n4222), .ZN(U3269)
         );
  XNOR2_X1 U4893 ( .A(n4224), .B(n4228), .ZN(n4386) );
  INV_X1 U4894 ( .A(n4225), .ZN(n4226) );
  NAND2_X1 U4895 ( .A1(n4227), .A2(n4226), .ZN(n4229) );
  XNOR2_X1 U4896 ( .A(n4229), .B(n4228), .ZN(n4235) );
  AOI22_X1 U4897 ( .A1(n4231), .A2(n4429), .B1(n4427), .B2(n4230), .ZN(n4232)
         );
  OAI21_X1 U4898 ( .B1(n4233), .B2(n4432), .A(n4232), .ZN(n4234) );
  AOI21_X1 U4899 ( .B1(n4235), .B2(n4437), .A(n4234), .ZN(n4236) );
  OAI21_X1 U4900 ( .B1(n4386), .B2(n4237), .A(n4236), .ZN(n4387) );
  NAND2_X1 U4901 ( .A1(n4387), .A2(n4238), .ZN(n4248) );
  INV_X1 U4902 ( .A(n4265), .ZN(n4242) );
  INV_X1 U4903 ( .A(n4239), .ZN(n4240) );
  OAI21_X1 U4904 ( .B1(n4242), .B2(n4241), .A(n4240), .ZN(n4478) );
  INV_X1 U4905 ( .A(n4478), .ZN(n4246) );
  INV_X1 U4906 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4244) );
  OAI22_X1 U4907 ( .A1(n4606), .A2(n4244), .B1(n4243), .B2(n4603), .ZN(n4245)
         );
  AOI21_X1 U4908 ( .B1(n4246), .B2(n4611), .A(n4245), .ZN(n4247) );
  OAI211_X1 U4909 ( .C1(n4386), .C2(n4608), .A(n4248), .B(n4247), .ZN(U3270)
         );
  XOR2_X1 U4910 ( .A(n4255), .B(n4249), .Z(n4391) );
  INV_X1 U4911 ( .A(n4391), .ZN(n4271) );
  NAND2_X1 U4912 ( .A1(n4251), .A2(n4250), .ZN(n4273) );
  INV_X1 U4913 ( .A(n4252), .ZN(n4254) );
  OAI21_X1 U4914 ( .B1(n4273), .B2(n4254), .A(n4253), .ZN(n4256) );
  XNOR2_X1 U4915 ( .A(n4256), .B(n4255), .ZN(n4262) );
  OAI22_X1 U4916 ( .A1(n4381), .A2(n4361), .B1(n4258), .B2(n4257), .ZN(n4259)
         );
  AOI21_X1 U4917 ( .B1(n4357), .B2(n4399), .A(n4259), .ZN(n4260) );
  OAI21_X1 U4918 ( .B1(n4262), .B2(n4261), .A(n4260), .ZN(n4390) );
  NAND2_X1 U4919 ( .A1(n4283), .A2(n4263), .ZN(n4264) );
  NAND2_X1 U4920 ( .A1(n4265), .A2(n4264), .ZN(n4482) );
  NOR2_X1 U4921 ( .A1(n4482), .A2(n4266), .ZN(n4269) );
  OAI22_X1 U4922 ( .A1(n4606), .A2(n4910), .B1(n4267), .B2(n4603), .ZN(n4268)
         );
  AOI211_X1 U4923 ( .C1(n4390), .C2(n4606), .A(n4269), .B(n4268), .ZN(n4270)
         );
  OAI21_X1 U4924 ( .B1(n4271), .B2(n4327), .A(n4270), .ZN(U3271) );
  XNOR2_X1 U4925 ( .A(n4273), .B(n4272), .ZN(n4279) );
  AOI22_X1 U4926 ( .A1(n4275), .A2(n4429), .B1(n4274), .B2(n4427), .ZN(n4276)
         );
  OAI21_X1 U4927 ( .B1(n4277), .B2(n4432), .A(n4276), .ZN(n4278) );
  AOI21_X1 U4928 ( .B1(n4279), .B2(n4437), .A(n4278), .ZN(n4396) );
  OAI21_X1 U4929 ( .B1(n4282), .B2(n4281), .A(n4280), .ZN(n4394) );
  OAI211_X1 U4930 ( .C1(n4298), .C2(n4284), .A(n4283), .B(n4412), .ZN(n4395)
         );
  INV_X1 U4931 ( .A(n4285), .ZN(n4286) );
  NOR2_X1 U4932 ( .A1(n4395), .A2(n4286), .ZN(n4289) );
  OAI22_X1 U4933 ( .A1(n4606), .A2(n4901), .B1(n4287), .B2(n4603), .ZN(n4288)
         );
  AOI211_X1 U4934 ( .C1(n4394), .C2(n4296), .A(n4289), .B(n4288), .ZN(n4290)
         );
  OAI21_X1 U4935 ( .B1(n4625), .B2(n4396), .A(n4290), .ZN(U3272) );
  INV_X1 U4936 ( .A(n4294), .ZN(n4291) );
  XNOR2_X1 U4937 ( .A(n4292), .B(n4291), .ZN(n4293) );
  NAND2_X1 U4938 ( .A1(n4293), .A2(n4437), .ZN(n4401) );
  XNOR2_X1 U4939 ( .A(n4295), .B(n4294), .ZN(n4404) );
  NAND2_X1 U4940 ( .A1(n4404), .A2(n4296), .ZN(n4308) );
  INV_X1 U4941 ( .A(n4297), .ZN(n4311) );
  INV_X1 U4942 ( .A(n4298), .ZN(n4299) );
  OAI21_X1 U4943 ( .B1(n4311), .B2(n4304), .A(n4299), .ZN(n4487) );
  INV_X1 U4944 ( .A(n4487), .ZN(n4306) );
  AOI22_X1 U4945 ( .A1(n4314), .A2(n4418), .B1(n4313), .B2(n4399), .ZN(n4303)
         );
  INV_X1 U4946 ( .A(n4300), .ZN(n4301) );
  AOI22_X1 U4947 ( .A1(n4625), .A2(REG2_REG_17__SCAN_IN), .B1(n4301), .B2(
        n4619), .ZN(n4302) );
  OAI211_X1 U4948 ( .C1(n4304), .C2(n4319), .A(n4303), .B(n4302), .ZN(n4305)
         );
  AOI21_X1 U4949 ( .B1(n4306), .B2(n4611), .A(n4305), .ZN(n4307) );
  OAI211_X1 U4950 ( .C1(n4625), .C2(n4401), .A(n4308), .B(n4307), .ZN(U3273)
         );
  OAI21_X1 U4951 ( .B1(n4310), .B2(n2622), .A(n4309), .ZN(n4416) );
  AOI21_X1 U4952 ( .B1(n4407), .B2(n4312), .A(n4311), .ZN(n4413) );
  AOI22_X1 U4953 ( .A1(n4314), .A2(n4430), .B1(n4313), .B2(n4408), .ZN(n4318)
         );
  INV_X1 U4954 ( .A(n4315), .ZN(n4316) );
  AOI22_X1 U4955 ( .A1(n4625), .A2(REG2_REG_16__SCAN_IN), .B1(n4316), .B2(
        n4619), .ZN(n4317) );
  OAI211_X1 U4956 ( .C1(n4320), .C2(n4319), .A(n4318), .B(n4317), .ZN(n4325)
         );
  OAI211_X1 U4957 ( .C1(n4323), .C2(n4322), .A(n4321), .B(n4437), .ZN(n4414)
         );
  NOR2_X1 U4958 ( .A1(n4414), .A2(n4625), .ZN(n4324) );
  AOI211_X1 U4959 ( .C1(n4413), .C2(n4611), .A(n4325), .B(n4324), .ZN(n4326)
         );
  OAI21_X1 U4960 ( .B1(n4327), .B2(n4416), .A(n4326), .ZN(U3274) );
  MUX2_X1 U4961 ( .A(n4328), .B(n4442), .S(n4657), .Z(n4329) );
  OAI21_X1 U4962 ( .B1(n4445), .B2(n4441), .A(n4329), .ZN(U3549) );
  AOI21_X1 U4963 ( .B1(n4333), .B2(n4331), .A(n4330), .ZN(n4511) );
  INV_X1 U4964 ( .A(n4511), .ZN(n4448) );
  AOI21_X1 U4965 ( .B1(n4333), .B2(n4427), .A(n4332), .ZN(n4513) );
  MUX2_X1 U4966 ( .A(n2749), .B(n4513), .S(n4657), .Z(n4334) );
  OAI21_X1 U4967 ( .B1(n4448), .B2(n4441), .A(n4334), .ZN(U3548) );
  AOI22_X1 U4968 ( .A1(n4336), .A2(n4357), .B1(n4335), .B2(n4427), .ZN(n4337)
         );
  OAI21_X1 U4969 ( .B1(n4338), .B2(n4361), .A(n4337), .ZN(n4339) );
  AOI211_X1 U4970 ( .C1(n4341), .C2(n4423), .A(n4340), .B(n4339), .ZN(n4449)
         );
  MUX2_X1 U4971 ( .A(n4342), .B(n4449), .S(n4657), .Z(n4343) );
  OAI21_X1 U4972 ( .B1(n4441), .B2(n4452), .A(n4343), .ZN(U3545) );
  AOI22_X1 U4973 ( .A1(n4345), .A2(n4429), .B1(n4427), .B2(n4344), .ZN(n4346)
         );
  OAI211_X1 U4974 ( .C1(n4362), .C2(n4432), .A(n4347), .B(n4346), .ZN(n4348)
         );
  AOI21_X1 U4975 ( .B1(n4349), .B2(n4423), .A(n4348), .ZN(n4453) );
  MUX2_X1 U4976 ( .A(n4350), .B(n4453), .S(n4657), .Z(n4351) );
  OAI21_X1 U4977 ( .B1(n4441), .B2(n4455), .A(n4351), .ZN(U3544) );
  AOI21_X1 U4978 ( .B1(n4353), .B2(n4423), .A(n4352), .ZN(n4456) );
  MUX2_X1 U4979 ( .A(n4354), .B(n4456), .S(n4657), .Z(n4355) );
  OAI21_X1 U4980 ( .B1(n4441), .B2(n4459), .A(n4355), .ZN(U3543) );
  INV_X1 U4981 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4365) );
  AOI22_X1 U4982 ( .A1(n4358), .A2(n4357), .B1(n4356), .B2(n4427), .ZN(n4359)
         );
  OAI211_X1 U4983 ( .C1(n4362), .C2(n4361), .A(n4360), .B(n4359), .ZN(n4363)
         );
  AOI21_X1 U4984 ( .B1(n4364), .B2(n4423), .A(n4363), .ZN(n4460) );
  MUX2_X1 U4985 ( .A(n4365), .B(n4460), .S(n4657), .Z(n4366) );
  OAI21_X1 U4986 ( .B1(n4441), .B2(n4462), .A(n4366), .ZN(U3542) );
  INV_X1 U4987 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4369) );
  AOI21_X1 U4988 ( .B1(n4368), .B2(n4423), .A(n4367), .ZN(n4463) );
  MUX2_X1 U4989 ( .A(n4369), .B(n4463), .S(n4657), .Z(n4370) );
  OAI21_X1 U4990 ( .B1(n4441), .B2(n4466), .A(n4370), .ZN(U3541) );
  NAND3_X1 U4991 ( .A1(n4372), .A2(n4423), .A3(n4371), .ZN(n4374) );
  NAND2_X1 U4992 ( .A1(n4374), .A2(n4373), .ZN(n4467) );
  MUX2_X1 U4993 ( .A(REG1_REG_22__SCAN_IN), .B(n4467), .S(n4657), .Z(n4375) );
  INV_X1 U4994 ( .A(n4375), .ZN(n4376) );
  OAI21_X1 U4995 ( .B1(n4441), .B2(n4470), .A(n4376), .ZN(U3540) );
  AOI22_X1 U4996 ( .A1(n4378), .A2(n4429), .B1(n4427), .B2(n4377), .ZN(n4379)
         );
  OAI211_X1 U4997 ( .C1(n4381), .C2(n4432), .A(n4380), .B(n4379), .ZN(n4382)
         );
  AOI21_X1 U4998 ( .B1(n4383), .B2(n4423), .A(n4382), .ZN(n4471) );
  MUX2_X1 U4999 ( .A(n4384), .B(n4471), .S(n4657), .Z(n4385) );
  OAI21_X1 U5000 ( .B1(n4441), .B2(n4474), .A(n4385), .ZN(U3539) );
  INV_X1 U5001 ( .A(n4386), .ZN(n4388) );
  AOI21_X1 U5002 ( .B1(n4645), .B2(n4388), .A(n4387), .ZN(n4476) );
  MUX2_X1 U5003 ( .A(n4776), .B(n4476), .S(n4657), .Z(n4389) );
  OAI21_X1 U5004 ( .B1(n4441), .B2(n4478), .A(n4389), .ZN(U3538) );
  AOI21_X1 U5005 ( .B1(n4391), .B2(n4423), .A(n4390), .ZN(n4479) );
  MUX2_X1 U5006 ( .A(n4392), .B(n4479), .S(n4657), .Z(n4393) );
  OAI21_X1 U5007 ( .B1(n4441), .B2(n4482), .A(n4393), .ZN(U3537) );
  INV_X1 U5008 ( .A(n4394), .ZN(n4397) );
  OAI211_X1 U5009 ( .C1(n4397), .C2(n4647), .A(n4396), .B(n4395), .ZN(n4483)
         );
  MUX2_X1 U5010 ( .A(REG1_REG_18__SCAN_IN), .B(n4483), .S(n4657), .Z(U3536) );
  AOI22_X1 U5011 ( .A1(n4399), .A2(n4429), .B1(n4427), .B2(n4398), .ZN(n4400)
         );
  OAI211_X1 U5012 ( .C1(n4402), .C2(n4432), .A(n4401), .B(n4400), .ZN(n4403)
         );
  AOI21_X1 U5013 ( .B1(n4404), .B2(n4423), .A(n4403), .ZN(n4485) );
  MUX2_X1 U5014 ( .A(n4485), .B(n4405), .S(n4655), .Z(n4406) );
  OAI21_X1 U5015 ( .B1(n4441), .B2(n4487), .A(n4406), .ZN(U3535) );
  AOI22_X1 U5016 ( .A1(n4408), .A2(n4429), .B1(n4407), .B2(n4427), .ZN(n4409)
         );
  OAI21_X1 U5017 ( .B1(n4410), .B2(n4432), .A(n4409), .ZN(n4411) );
  AOI21_X1 U5018 ( .B1(n4413), .B2(n4412), .A(n4411), .ZN(n4415) );
  OAI211_X1 U5019 ( .C1(n4416), .C2(n4647), .A(n4415), .B(n4414), .ZN(n4488)
         );
  MUX2_X1 U5020 ( .A(REG1_REG_16__SCAN_IN), .B(n4488), .S(n4657), .Z(U3534) );
  AOI22_X1 U5021 ( .A1(n4418), .A2(n4429), .B1(n4427), .B2(n4417), .ZN(n4419)
         );
  OAI211_X1 U5022 ( .C1(n4421), .C2(n4432), .A(n4420), .B(n4419), .ZN(n4422)
         );
  AOI21_X1 U5023 ( .B1(n4424), .B2(n4423), .A(n4422), .ZN(n4489) );
  MUX2_X1 U5024 ( .A(n4425), .B(n4489), .S(n4657), .Z(n4426) );
  OAI21_X1 U5025 ( .B1(n4441), .B2(n4492), .A(n4426), .ZN(U3533) );
  AOI22_X1 U5026 ( .A1(n4430), .A2(n4429), .B1(n4428), .B2(n4427), .ZN(n4431)
         );
  OAI21_X1 U5027 ( .B1(n4433), .B2(n4432), .A(n4431), .ZN(n4436) );
  NOR2_X1 U5028 ( .A1(n4434), .A2(n4647), .ZN(n4435) );
  AOI211_X1 U5029 ( .C1(n4438), .C2(n4437), .A(n4436), .B(n4435), .ZN(n4493)
         );
  MUX2_X1 U5030 ( .A(n4439), .B(n4493), .S(n4657), .Z(n4440) );
  OAI21_X1 U5031 ( .B1(n4441), .B2(n4496), .A(n4440), .ZN(U3532) );
  NOR2_X1 U5032 ( .A1(n4442), .A2(n4653), .ZN(n4443) );
  AOI21_X1 U5033 ( .B1(REG0_REG_31__SCAN_IN), .B2(n4653), .A(n4443), .ZN(n4444) );
  OAI21_X1 U5034 ( .B1(n4445), .B2(n4495), .A(n4444), .ZN(U3517) );
  INV_X1 U5035 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4446) );
  MUX2_X1 U5036 ( .A(n4446), .B(n4513), .S(n4475), .Z(n4447) );
  OAI21_X1 U5037 ( .B1(n4448), .B2(n4495), .A(n4447), .ZN(U3516) );
  INV_X1 U5038 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4450) );
  MUX2_X1 U5039 ( .A(n4450), .B(n4449), .S(n4475), .Z(n4451) );
  OAI21_X1 U5040 ( .B1(n4452), .B2(n4495), .A(n4451), .ZN(U3513) );
  INV_X1 U5041 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4764) );
  MUX2_X1 U5042 ( .A(n4764), .B(n4453), .S(n4475), .Z(n4454) );
  OAI21_X1 U5043 ( .B1(n4455), .B2(n4495), .A(n4454), .ZN(U3512) );
  INV_X1 U5044 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4457) );
  MUX2_X1 U5045 ( .A(n4457), .B(n4456), .S(n4475), .Z(n4458) );
  OAI21_X1 U5046 ( .B1(n4459), .B2(n4495), .A(n4458), .ZN(U3511) );
  INV_X1 U5047 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4765) );
  MUX2_X1 U5048 ( .A(n4765), .B(n4460), .S(n4475), .Z(n4461) );
  OAI21_X1 U5049 ( .B1(n4462), .B2(n4495), .A(n4461), .ZN(U3510) );
  INV_X1 U5050 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4464) );
  MUX2_X1 U5051 ( .A(n4464), .B(n4463), .S(n4475), .Z(n4465) );
  OAI21_X1 U5052 ( .B1(n4466), .B2(n4495), .A(n4465), .ZN(U3509) );
  MUX2_X1 U5053 ( .A(REG0_REG_22__SCAN_IN), .B(n4467), .S(n4475), .Z(n4468) );
  INV_X1 U5054 ( .A(n4468), .ZN(n4469) );
  OAI21_X1 U5055 ( .B1(n4470), .B2(n4495), .A(n4469), .ZN(U3508) );
  INV_X1 U5056 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4472) );
  MUX2_X1 U5057 ( .A(n4472), .B(n4471), .S(n4475), .Z(n4473) );
  OAI21_X1 U5058 ( .B1(n4474), .B2(n4495), .A(n4473), .ZN(U3507) );
  INV_X1 U5059 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4750) );
  MUX2_X1 U5060 ( .A(n4750), .B(n4476), .S(n4475), .Z(n4477) );
  OAI21_X1 U5061 ( .B1(n4478), .B2(n4495), .A(n4477), .ZN(U3506) );
  INV_X1 U5062 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4480) );
  MUX2_X1 U5063 ( .A(n4480), .B(n4479), .S(n4475), .Z(n4481) );
  OAI21_X1 U5064 ( .B1(n4482), .B2(n4495), .A(n4481), .ZN(U3505) );
  MUX2_X1 U5065 ( .A(REG0_REG_18__SCAN_IN), .B(n4483), .S(n4475), .Z(U3503) );
  INV_X1 U5066 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4484) );
  MUX2_X1 U5067 ( .A(n4485), .B(n4484), .S(n4653), .Z(n4486) );
  OAI21_X1 U5068 ( .B1(n4487), .B2(n4495), .A(n4486), .ZN(U3501) );
  MUX2_X1 U5069 ( .A(REG0_REG_16__SCAN_IN), .B(n4488), .S(n4475), .Z(U3499) );
  INV_X1 U5070 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4490) );
  MUX2_X1 U5071 ( .A(n4490), .B(n4489), .S(n4475), .Z(n4491) );
  OAI21_X1 U5072 ( .B1(n4492), .B2(n4495), .A(n4491), .ZN(U3497) );
  INV_X1 U5073 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4748) );
  MUX2_X1 U5074 ( .A(n4748), .B(n4493), .S(n4475), .Z(n4494) );
  OAI21_X1 U5075 ( .B1(n4496), .B2(n4495), .A(n4494), .ZN(U3495) );
  MUX2_X1 U5076 ( .A(DATAI_28_), .B(n4497), .S(STATE_REG_SCAN_IN), .Z(U3324)
         );
  MUX2_X1 U5077 ( .A(n4498), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5078 ( .A(DATAI_25_), .B(n4499), .S(STATE_REG_SCAN_IN), .Z(U3327)
         );
  MUX2_X1 U5079 ( .A(n4500), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U5080 ( .A(n4501), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U5081 ( .A(DATAI_20_), .B(n4502), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5082 ( .A(n4503), .B(DATAI_13_), .S(U3149), .Z(U3339) );
  MUX2_X1 U5083 ( .A(n4504), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U5084 ( .A(n4505), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5085 ( .A(n4506), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5086 ( .A(DATAI_4_), .B(n4507), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5087 ( .A(DATAI_3_), .B(n4508), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U5088 ( .A(n4509), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5089 ( .A(n4510), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  MUX2_X1 U5090 ( .A(DATAI_0_), .B(n4877), .S(STATE_REG_SCAN_IN), .Z(U3352) );
  AOI22_X1 U5091 ( .A1(n4511), .A2(n4611), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4625), .ZN(n4512) );
  OAI21_X1 U5092 ( .B1(n4625), .B2(n4513), .A(n4512), .ZN(U3261) );
  OAI211_X1 U5093 ( .C1(n4516), .C2(n4515), .A(n4595), .B(n4514), .ZN(n4520)
         );
  OAI211_X1 U5094 ( .C1(n4518), .C2(n2197), .A(n4584), .B(n4517), .ZN(n4519)
         );
  OAI211_X1 U5095 ( .C1(n4602), .C2(n4639), .A(n4520), .B(n4519), .ZN(n4521)
         );
  AOI211_X1 U5096 ( .C1(n4594), .C2(ADDR_REG_9__SCAN_IN), .A(n4522), .B(n4521), 
        .ZN(n4523) );
  INV_X1 U5097 ( .A(n4523), .ZN(U3249) );
  OAI211_X1 U5098 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4525), .A(n4584), .B(n4524), .ZN(n4527) );
  NAND2_X1 U5099 ( .A1(n4527), .A2(n4526), .ZN(n4528) );
  AOI21_X1 U5100 ( .B1(n4594), .B2(ADDR_REG_10__SCAN_IN), .A(n4528), .ZN(n4532) );
  OAI211_X1 U5101 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4530), .A(n4595), .B(n4529), .ZN(n4531) );
  OAI211_X1 U5102 ( .C1(n4602), .C2(n4638), .A(n4532), .B(n4531), .ZN(U3250)
         );
  OAI211_X1 U5103 ( .C1(n4535), .C2(n4534), .A(n4595), .B(n4533), .ZN(n4540)
         );
  OAI211_X1 U5104 ( .C1(n4538), .C2(n4537), .A(n4584), .B(n4536), .ZN(n4539)
         );
  OAI211_X1 U5105 ( .C1(n4602), .C2(n4637), .A(n4540), .B(n4539), .ZN(n4541)
         );
  AOI211_X1 U5106 ( .C1(n4594), .C2(ADDR_REG_11__SCAN_IN), .A(n4542), .B(n4541), .ZN(n4543) );
  INV_X1 U5107 ( .A(n4543), .ZN(U3251) );
  OAI211_X1 U5108 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4545), .A(n4584), .B(n4544), .ZN(n4547) );
  NAND2_X1 U5109 ( .A1(n4547), .A2(n4546), .ZN(n4548) );
  AOI21_X1 U5110 ( .B1(n4594), .B2(ADDR_REG_12__SCAN_IN), .A(n4548), .ZN(n4552) );
  OAI211_X1 U5111 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4550), .A(n4595), .B(n4549), .ZN(n4551) );
  OAI211_X1 U5112 ( .C1(n4602), .C2(n4553), .A(n4552), .B(n4551), .ZN(U3252)
         );
  INV_X1 U5113 ( .A(n4554), .ZN(n4559) );
  AOI211_X1 U5114 ( .C1(n4557), .C2(n4556), .A(n4555), .B(n4588), .ZN(n4558)
         );
  AOI211_X1 U5115 ( .C1(n4594), .C2(ADDR_REG_14__SCAN_IN), .A(n4559), .B(n4558), .ZN(n4563) );
  OAI211_X1 U5116 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4561), .A(n4595), .B(n4560), .ZN(n4562) );
  OAI211_X1 U5117 ( .C1(n4602), .C2(n2269), .A(n4563), .B(n4562), .ZN(U3254)
         );
  AOI211_X1 U5118 ( .C1(n4566), .C2(n4565), .A(n4564), .B(n4588), .ZN(n4567)
         );
  AOI211_X1 U5119 ( .C1(n4594), .C2(ADDR_REG_15__SCAN_IN), .A(n4568), .B(n4567), .ZN(n4573) );
  OAI211_X1 U5120 ( .C1(n4571), .C2(n4570), .A(n4595), .B(n4569), .ZN(n4572)
         );
  OAI211_X1 U5121 ( .C1(n4602), .C2(n4631), .A(n4573), .B(n4572), .ZN(U3255)
         );
  INV_X1 U5122 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n4797) );
  OAI21_X1 U5123 ( .B1(n4576), .B2(n4575), .A(n4574), .ZN(n4583) );
  AOI21_X1 U5124 ( .B1(n4578), .B2(REG1_REG_16__SCAN_IN), .A(n4577), .ZN(n4581) );
  OAI22_X1 U5125 ( .A1(n4581), .A2(n4580), .B1(n4579), .B2(n4602), .ZN(n4582)
         );
  AOI21_X1 U5126 ( .B1(n4584), .B2(n4583), .A(n4582), .ZN(n4586) );
  OAI211_X1 U5127 ( .C1(n4587), .C2(n4797), .A(n4586), .B(n4585), .ZN(U3256)
         );
  AOI221_X1 U5128 ( .B1(n4591), .B2(n4590), .C1(n4589), .C2(n4590), .A(n4588), 
        .ZN(n4592) );
  AOI211_X1 U5129 ( .C1(n4594), .C2(ADDR_REG_17__SCAN_IN), .A(n4593), .B(n4592), .ZN(n4600) );
  OAI221_X1 U5130 ( .B1(n4598), .B2(n4597), .C1(n4598), .C2(n4596), .A(n4595), 
        .ZN(n4599) );
  OAI211_X1 U5131 ( .C1(n4602), .C2(n4601), .A(n4600), .B(n4599), .ZN(U3257)
         );
  OAI22_X1 U5132 ( .A1(n4606), .A2(n4605), .B1(n4604), .B2(n4603), .ZN(n4607)
         );
  INV_X1 U5133 ( .A(n4607), .ZN(n4614) );
  INV_X1 U5134 ( .A(n4608), .ZN(n4620) );
  INV_X1 U5135 ( .A(n4609), .ZN(n4610) );
  AOI22_X1 U5136 ( .A1(n4612), .A2(n4620), .B1(n4611), .B2(n4610), .ZN(n4613)
         );
  OAI211_X1 U5137 ( .C1(n4625), .C2(n4615), .A(n4614), .B(n4613), .ZN(U3282)
         );
  AOI21_X1 U5138 ( .B1(n4618), .B2(n4617), .A(n4616), .ZN(n4624) );
  AOI22_X1 U5139 ( .A1(n4621), .A2(n4620), .B1(REG3_REG_0__SCAN_IN), .B2(n4619), .ZN(n4622) );
  OAI221_X1 U5140 ( .B1(n4625), .B2(n4624), .C1(n4606), .C2(n4623), .A(n4622), 
        .ZN(U3290) );
  AND2_X1 U5141 ( .A1(D_REG_31__SCAN_IN), .A2(n4942), .ZN(U3291) );
  INV_X1 U5142 ( .A(D_REG_30__SCAN_IN), .ZN(n4737) );
  NOR2_X1 U5143 ( .A1(n4626), .A2(n4737), .ZN(U3292) );
  INV_X1 U5144 ( .A(D_REG_29__SCAN_IN), .ZN(n4736) );
  NOR2_X1 U5145 ( .A1(n4626), .A2(n4736), .ZN(U3293) );
  AND2_X1 U5146 ( .A1(D_REG_28__SCAN_IN), .A2(n4942), .ZN(U3294) );
  INV_X1 U5147 ( .A(D_REG_27__SCAN_IN), .ZN(n4734) );
  NOR2_X1 U5148 ( .A1(n4626), .A2(n4734), .ZN(U3295) );
  INV_X1 U5149 ( .A(D_REG_26__SCAN_IN), .ZN(n4733) );
  NOR2_X1 U5150 ( .A1(n4626), .A2(n4733), .ZN(U3296) );
  INV_X1 U5151 ( .A(D_REG_25__SCAN_IN), .ZN(n4730) );
  NOR2_X1 U5152 ( .A1(n4626), .A2(n4730), .ZN(U3297) );
  AND2_X1 U5153 ( .A1(D_REG_24__SCAN_IN), .A2(n4942), .ZN(U3298) );
  AND2_X1 U5154 ( .A1(D_REG_23__SCAN_IN), .A2(n4942), .ZN(U3299) );
  INV_X1 U5155 ( .A(D_REG_22__SCAN_IN), .ZN(n4731) );
  NOR2_X1 U5156 ( .A1(n4626), .A2(n4731), .ZN(U3300) );
  INV_X1 U5157 ( .A(D_REG_21__SCAN_IN), .ZN(n4724) );
  NOR2_X1 U5158 ( .A1(n4626), .A2(n4724), .ZN(U3301) );
  INV_X1 U5159 ( .A(D_REG_20__SCAN_IN), .ZN(n4723) );
  NOR2_X1 U5160 ( .A1(n4626), .A2(n4723), .ZN(U3302) );
  INV_X1 U5161 ( .A(D_REG_19__SCAN_IN), .ZN(n4720) );
  NOR2_X1 U5162 ( .A1(n4626), .A2(n4720), .ZN(U3303) );
  AND2_X1 U5163 ( .A1(D_REG_18__SCAN_IN), .A2(n4942), .ZN(U3304) );
  AND2_X1 U5164 ( .A1(D_REG_17__SCAN_IN), .A2(n4942), .ZN(U3305) );
  AND2_X1 U5165 ( .A1(D_REG_16__SCAN_IN), .A2(n4942), .ZN(U3306) );
  AND2_X1 U5166 ( .A1(D_REG_15__SCAN_IN), .A2(n4942), .ZN(U3307) );
  INV_X1 U5167 ( .A(D_REG_14__SCAN_IN), .ZN(n4721) );
  NOR2_X1 U5168 ( .A1(n4626), .A2(n4721), .ZN(U3308) );
  AND2_X1 U5169 ( .A1(D_REG_13__SCAN_IN), .A2(n4942), .ZN(U3309) );
  INV_X1 U5170 ( .A(D_REG_11__SCAN_IN), .ZN(n4717) );
  NOR2_X1 U5171 ( .A1(n4626), .A2(n4717), .ZN(U3311) );
  AND2_X1 U5172 ( .A1(D_REG_10__SCAN_IN), .A2(n4942), .ZN(U3312) );
  INV_X1 U5173 ( .A(D_REG_9__SCAN_IN), .ZN(n4848) );
  NOR2_X1 U5174 ( .A1(n4626), .A2(n4848), .ZN(U3313) );
  INV_X1 U5175 ( .A(D_REG_8__SCAN_IN), .ZN(n4846) );
  NOR2_X1 U5176 ( .A1(n4626), .A2(n4846), .ZN(U3314) );
  AND2_X1 U5177 ( .A1(D_REG_7__SCAN_IN), .A2(n4942), .ZN(U3315) );
  INV_X1 U5178 ( .A(D_REG_6__SCAN_IN), .ZN(n4714) );
  NOR2_X1 U5179 ( .A1(n4626), .A2(n4714), .ZN(U3316) );
  AND2_X1 U5180 ( .A1(D_REG_5__SCAN_IN), .A2(n4942), .ZN(U3317) );
  AND2_X1 U5181 ( .A1(D_REG_4__SCAN_IN), .A2(n4942), .ZN(U3318) );
  AND2_X1 U5182 ( .A1(D_REG_3__SCAN_IN), .A2(n4942), .ZN(U3319) );
  INV_X1 U5183 ( .A(D_REG_2__SCAN_IN), .ZN(n4715) );
  NOR2_X1 U5184 ( .A1(n4626), .A2(n4715), .ZN(U3320) );
  OAI21_X1 U5185 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4627), .ZN(
        n4628) );
  INV_X1 U5186 ( .A(n4628), .ZN(U3329) );
  OAI22_X1 U5187 ( .A1(U3149), .A2(n4629), .B1(DATAI_17_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4630) );
  INV_X1 U5188 ( .A(n4630), .ZN(U3335) );
  INV_X1 U5189 ( .A(DATAI_15_), .ZN(n4873) );
  AOI22_X1 U5190 ( .A1(STATE_REG_SCAN_IN), .A2(n4631), .B1(n4873), .B2(U3149), 
        .ZN(U3337) );
  OAI22_X1 U5191 ( .A1(U3149), .A2(n4632), .B1(DATAI_14_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4633) );
  INV_X1 U5192 ( .A(n4633), .ZN(U3338) );
  OAI22_X1 U5193 ( .A1(U3149), .A2(n4634), .B1(DATAI_12_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4635) );
  INV_X1 U5194 ( .A(n4635), .ZN(U3340) );
  INV_X1 U5195 ( .A(DATAI_11_), .ZN(n4636) );
  AOI22_X1 U5196 ( .A1(STATE_REG_SCAN_IN), .A2(n4637), .B1(n4636), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5197 ( .A(DATAI_10_), .ZN(n4871) );
  AOI22_X1 U5198 ( .A1(STATE_REG_SCAN_IN), .A2(n4638), .B1(n4871), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5199 ( .A(DATAI_9_), .ZN(n4870) );
  AOI22_X1 U5200 ( .A1(STATE_REG_SCAN_IN), .A2(n4639), .B1(n4870), .B2(U3149), 
        .ZN(U3343) );
  INV_X1 U5201 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4740) );
  AOI22_X1 U5202 ( .A1(n4475), .A2(n4640), .B1(n4740), .B2(n4653), .ZN(U3467)
         );
  INV_X1 U5203 ( .A(n4641), .ZN(n4646) );
  INV_X1 U5204 ( .A(n4642), .ZN(n4644) );
  AOI211_X1 U5205 ( .C1(n4646), .C2(n4645), .A(n4644), .B(n4643), .ZN(n4654)
         );
  INV_X1 U5206 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4739) );
  AOI22_X1 U5207 ( .A1(n4475), .A2(n4654), .B1(n4739), .B2(n4653), .ZN(U3475)
         );
  NOR2_X1 U5208 ( .A1(n4648), .A2(n4647), .ZN(n4652) );
  AOI211_X1 U5209 ( .C1(n4652), .C2(n4651), .A(n4650), .B(n4649), .ZN(n4656)
         );
  INV_X1 U5210 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4883) );
  AOI22_X1 U5211 ( .A1(n4475), .A2(n4656), .B1(n4883), .B2(n4653), .ZN(U3481)
         );
  AOI22_X1 U5212 ( .A1(n4657), .A2(n4654), .B1(n2480), .B2(n4655), .ZN(U3522)
         );
  AOI22_X1 U5213 ( .A1(n4657), .A2(n4656), .B1(n2515), .B2(n4655), .ZN(U3525)
         );
  AOI22_X1 U5214 ( .A1(n4864), .A2(keyinput65), .B1(n4865), .B2(keyinput2), 
        .ZN(n4658) );
  OAI221_X1 U5215 ( .B1(n4864), .B2(keyinput65), .C1(n4865), .C2(keyinput2), 
        .A(n4658), .ZN(n4668) );
  AOI22_X1 U5216 ( .A1(n4660), .A2(keyinput78), .B1(n4866), .B2(keyinput123), 
        .ZN(n4659) );
  OAI221_X1 U5217 ( .B1(n4660), .B2(keyinput78), .C1(n4866), .C2(keyinput123), 
        .A(n4659), .ZN(n4667) );
  INV_X1 U5218 ( .A(DATAI_21_), .ZN(n4662) );
  AOI22_X1 U5219 ( .A1(n4872), .A2(keyinput70), .B1(n4662), .B2(keyinput122), 
        .ZN(n4661) );
  OAI221_X1 U5220 ( .B1(n4872), .B2(keyinput70), .C1(n4662), .C2(keyinput122), 
        .A(n4661), .ZN(n4666) );
  AOI22_X1 U5221 ( .A1(n4664), .A2(keyinput35), .B1(keyinput74), .B2(n4873), 
        .ZN(n4663) );
  OAI221_X1 U5222 ( .B1(n4664), .B2(keyinput35), .C1(n4873), .C2(keyinput74), 
        .A(n4663), .ZN(n4665) );
  NOR4_X1 U5223 ( .A1(n4668), .A2(n4667), .A3(n4666), .A4(n4665), .ZN(n4702)
         );
  INV_X1 U5224 ( .A(DATAI_4_), .ZN(n4868) );
  AOI22_X1 U5225 ( .A1(n4868), .A2(keyinput100), .B1(n4869), .B2(keyinput8), 
        .ZN(n4669) );
  OAI221_X1 U5226 ( .B1(n4868), .B2(keyinput100), .C1(n4869), .C2(keyinput8), 
        .A(n4669), .ZN(n4678) );
  AOI22_X1 U5227 ( .A1(n4871), .A2(keyinput47), .B1(keyinput57), .B2(n4870), 
        .ZN(n4670) );
  OAI221_X1 U5228 ( .B1(n4871), .B2(keyinput47), .C1(n4870), .C2(keyinput57), 
        .A(n4670), .ZN(n4677) );
  AOI22_X1 U5229 ( .A1(n4890), .A2(keyinput60), .B1(n4672), .B2(keyinput112), 
        .ZN(n4671) );
  OAI221_X1 U5230 ( .B1(n4890), .B2(keyinput60), .C1(n4672), .C2(keyinput112), 
        .A(n4671), .ZN(n4676) );
  XNOR2_X1 U5231 ( .A(DATAI_0_), .B(keyinput6), .ZN(n4674) );
  XNOR2_X1 U5232 ( .A(DATAI_3_), .B(keyinput84), .ZN(n4673) );
  NAND2_X1 U5233 ( .A1(n4674), .A2(n4673), .ZN(n4675) );
  NOR4_X1 U5234 ( .A1(n4678), .A2(n4677), .A3(n4676), .A4(n4675), .ZN(n4701)
         );
  AOI22_X1 U5235 ( .A1(n4680), .A2(keyinput114), .B1(keyinput97), .B2(n2489), 
        .ZN(n4679) );
  OAI221_X1 U5236 ( .B1(n4680), .B2(keyinput114), .C1(n2489), .C2(keyinput97), 
        .A(n4679), .ZN(n4688) );
  AOI22_X1 U5237 ( .A1(n2701), .A2(keyinput125), .B1(keyinput72), .B2(n3705), 
        .ZN(n4681) );
  OAI221_X1 U5238 ( .B1(n2701), .B2(keyinput125), .C1(n3705), .C2(keyinput72), 
        .A(n4681), .ZN(n4687) );
  XNOR2_X1 U5239 ( .A(REG3_REG_10__SCAN_IN), .B(keyinput83), .ZN(n4685) );
  XNOR2_X1 U5240 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput44), .ZN(n4684) );
  XNOR2_X1 U5241 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput48), .ZN(n4683) );
  XNOR2_X1 U5242 ( .A(REG3_REG_24__SCAN_IN), .B(keyinput31), .ZN(n4682) );
  NAND4_X1 U5243 ( .A1(n4685), .A2(n4684), .A3(n4683), .A4(n4682), .ZN(n4686)
         );
  NOR3_X1 U5244 ( .A1(n4688), .A2(n4687), .A3(n4686), .ZN(n4700) );
  XNOR2_X1 U5245 ( .A(IR_REG_1__SCAN_IN), .B(keyinput23), .ZN(n4692) );
  XNOR2_X1 U5246 ( .A(n4877), .B(keyinput61), .ZN(n4691) );
  XNOR2_X1 U5247 ( .A(IR_REG_6__SCAN_IN), .B(keyinput28), .ZN(n4690) );
  XNOR2_X1 U5248 ( .A(IR_REG_4__SCAN_IN), .B(keyinput118), .ZN(n4689) );
  NAND4_X1 U5249 ( .A1(n4692), .A2(n4691), .A3(n4690), .A4(n4689), .ZN(n4698)
         );
  XNOR2_X1 U5250 ( .A(IR_REG_12__SCAN_IN), .B(keyinput116), .ZN(n4696) );
  XNOR2_X1 U5251 ( .A(IR_REG_7__SCAN_IN), .B(keyinput81), .ZN(n4695) );
  XNOR2_X1 U5252 ( .A(IR_REG_16__SCAN_IN), .B(keyinput14), .ZN(n4694) );
  XNOR2_X1 U5253 ( .A(IR_REG_13__SCAN_IN), .B(keyinput29), .ZN(n4693) );
  NAND4_X1 U5254 ( .A1(n4696), .A2(n4695), .A3(n4694), .A4(n4693), .ZN(n4697)
         );
  NOR2_X1 U5255 ( .A1(n4698), .A2(n4697), .ZN(n4699) );
  NAND4_X1 U5256 ( .A1(n4702), .A2(n4701), .A3(n4700), .A4(n4699), .ZN(n4861)
         );
  XNOR2_X1 U5257 ( .A(IR_REG_21__SCAN_IN), .B(keyinput76), .ZN(n4706) );
  XNOR2_X1 U5258 ( .A(IR_REG_18__SCAN_IN), .B(keyinput106), .ZN(n4705) );
  XNOR2_X1 U5259 ( .A(IR_REG_25__SCAN_IN), .B(keyinput24), .ZN(n4704) );
  XNOR2_X1 U5260 ( .A(IR_REG_24__SCAN_IN), .B(keyinput18), .ZN(n4703) );
  NAND4_X1 U5261 ( .A1(n4706), .A2(n4705), .A3(n4704), .A4(n4703), .ZN(n4712)
         );
  XNOR2_X1 U5262 ( .A(IR_REG_28__SCAN_IN), .B(keyinput33), .ZN(n4710) );
  XNOR2_X1 U5263 ( .A(IR_REG_26__SCAN_IN), .B(keyinput30), .ZN(n4709) );
  XNOR2_X1 U5264 ( .A(D_REG_0__SCAN_IN), .B(keyinput87), .ZN(n4708) );
  XNOR2_X1 U5265 ( .A(IR_REG_31__SCAN_IN), .B(keyinput16), .ZN(n4707) );
  NAND4_X1 U5266 ( .A1(n4710), .A2(n4709), .A3(n4708), .A4(n4707), .ZN(n4711)
         );
  NOR2_X1 U5267 ( .A1(n4712), .A2(n4711), .ZN(n4759) );
  AOI22_X1 U5268 ( .A1(n4715), .A2(keyinput56), .B1(keyinput38), .B2(n4714), 
        .ZN(n4713) );
  OAI221_X1 U5269 ( .B1(n4715), .B2(keyinput56), .C1(n4714), .C2(keyinput38), 
        .A(n4713), .ZN(n4728) );
  INV_X1 U5270 ( .A(D_REG_12__SCAN_IN), .ZN(n4718) );
  AOI22_X1 U5271 ( .A1(n4718), .A2(keyinput121), .B1(keyinput21), .B2(n4717), 
        .ZN(n4716) );
  OAI221_X1 U5272 ( .B1(n4718), .B2(keyinput121), .C1(n4717), .C2(keyinput21), 
        .A(n4716), .ZN(n4727) );
  AOI22_X1 U5273 ( .A1(n4721), .A2(keyinput85), .B1(n4720), .B2(keyinput103), 
        .ZN(n4719) );
  OAI221_X1 U5274 ( .B1(n4721), .B2(keyinput85), .C1(n4720), .C2(keyinput103), 
        .A(n4719), .ZN(n4726) );
  AOI22_X1 U5275 ( .A1(n4724), .A2(keyinput117), .B1(n4723), .B2(keyinput80), 
        .ZN(n4722) );
  OAI221_X1 U5276 ( .B1(n4724), .B2(keyinput117), .C1(n4723), .C2(keyinput80), 
        .A(n4722), .ZN(n4725) );
  NOR4_X1 U5277 ( .A1(n4728), .A2(n4727), .A3(n4726), .A4(n4725), .ZN(n4758)
         );
  AOI22_X1 U5278 ( .A1(n4731), .A2(keyinput49), .B1(keyinput68), .B2(n4730), 
        .ZN(n4729) );
  OAI221_X1 U5279 ( .B1(n4731), .B2(keyinput49), .C1(n4730), .C2(keyinput68), 
        .A(n4729), .ZN(n4744) );
  AOI22_X1 U5280 ( .A1(n4734), .A2(keyinput88), .B1(keyinput10), .B2(n4733), 
        .ZN(n4732) );
  OAI221_X1 U5281 ( .B1(n4734), .B2(keyinput88), .C1(n4733), .C2(keyinput10), 
        .A(n4732), .ZN(n4743) );
  AOI22_X1 U5282 ( .A1(n4737), .A2(keyinput94), .B1(keyinput34), .B2(n4736), 
        .ZN(n4735) );
  OAI221_X1 U5283 ( .B1(n4737), .B2(keyinput94), .C1(n4736), .C2(keyinput34), 
        .A(n4735), .ZN(n4742) );
  AOI22_X1 U5284 ( .A1(n4740), .A2(keyinput13), .B1(n4739), .B2(keyinput109), 
        .ZN(n4738) );
  OAI221_X1 U5285 ( .B1(n4740), .B2(keyinput13), .C1(n4739), .C2(keyinput109), 
        .A(n4738), .ZN(n4741) );
  NOR4_X1 U5286 ( .A1(n4744), .A2(n4743), .A3(n4742), .A4(n4741), .ZN(n4757)
         );
  INV_X1 U5287 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4746) );
  AOI22_X1 U5288 ( .A1(n4883), .A2(keyinput58), .B1(n4746), .B2(keyinput32), 
        .ZN(n4745) );
  OAI221_X1 U5289 ( .B1(n4883), .B2(keyinput58), .C1(n4746), .C2(keyinput32), 
        .A(n4745), .ZN(n4755) );
  AOI22_X1 U5290 ( .A1(n4748), .A2(keyinput46), .B1(keyinput67), .B2(n3453), 
        .ZN(n4747) );
  OAI221_X1 U5291 ( .B1(n4748), .B2(keyinput46), .C1(n3453), .C2(keyinput67), 
        .A(n4747), .ZN(n4754) );
  INV_X1 U5292 ( .A(REG0_REG_18__SCAN_IN), .ZN(n4884) );
  AOI22_X1 U5293 ( .A1(n4884), .A2(keyinput15), .B1(n4750), .B2(keyinput9), 
        .ZN(n4749) );
  OAI221_X1 U5294 ( .B1(n4884), .B2(keyinput15), .C1(n4750), .C2(keyinput9), 
        .A(n4749), .ZN(n4753) );
  AOI22_X1 U5295 ( .A1(n4472), .A2(keyinput7), .B1(n4464), .B2(keyinput51), 
        .ZN(n4751) );
  OAI221_X1 U5296 ( .B1(n4472), .B2(keyinput7), .C1(n4464), .C2(keyinput51), 
        .A(n4751), .ZN(n4752) );
  NOR4_X1 U5297 ( .A1(n4755), .A2(n4754), .A3(n4753), .A4(n4752), .ZN(n4756)
         );
  NAND4_X1 U5298 ( .A1(n4759), .A2(n4758), .A3(n4757), .A4(n4756), .ZN(n4860)
         );
  AOI22_X1 U5299 ( .A1(n2467), .A2(keyinput62), .B1(n2480), .B2(keyinput36), 
        .ZN(n4760) );
  OAI221_X1 U5300 ( .B1(n2467), .B2(keyinput62), .C1(n2480), .C2(keyinput36), 
        .A(n4760), .ZN(n4772) );
  AOI22_X1 U5301 ( .A1(n2504), .A2(keyinput41), .B1(n4762), .B2(keyinput91), 
        .ZN(n4761) );
  OAI221_X1 U5302 ( .B1(n2504), .B2(keyinput41), .C1(n4762), .C2(keyinput91), 
        .A(n4761), .ZN(n4771) );
  AOI22_X1 U5303 ( .A1(n4765), .A2(keyinput120), .B1(n4764), .B2(keyinput104), 
        .ZN(n4763) );
  OAI221_X1 U5304 ( .B1(n4765), .B2(keyinput120), .C1(n4764), .C2(keyinput104), 
        .A(n4763), .ZN(n4770) );
  INV_X1 U5305 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4766) );
  XOR2_X1 U5306 ( .A(n4766), .B(keyinput113), .Z(n4768) );
  XNOR2_X1 U5307 ( .A(REG1_REG_2__SCAN_IN), .B(keyinput4), .ZN(n4767) );
  NAND2_X1 U5308 ( .A1(n4768), .A2(n4767), .ZN(n4769) );
  NOR4_X1 U5309 ( .A1(n4772), .A2(n4771), .A3(n4770), .A4(n4769), .ZN(n4807)
         );
  AOI22_X1 U5310 ( .A1(n4425), .A2(keyinput25), .B1(n4774), .B2(keyinput111), 
        .ZN(n4773) );
  OAI221_X1 U5311 ( .B1(n4425), .B2(keyinput25), .C1(n4774), .C2(keyinput111), 
        .A(n4773), .ZN(n4782) );
  AOI22_X1 U5312 ( .A1(n4776), .A2(keyinput99), .B1(n4354), .B2(keyinput0), 
        .ZN(n4775) );
  OAI221_X1 U5313 ( .B1(n4776), .B2(keyinput99), .C1(n4354), .C2(keyinput0), 
        .A(n4775), .ZN(n4781) );
  AOI22_X1 U5314 ( .A1(n4342), .A2(keyinput79), .B1(n4915), .B2(keyinput102), 
        .ZN(n4777) );
  OAI221_X1 U5315 ( .B1(n4342), .B2(keyinput79), .C1(n4915), .C2(keyinput102), 
        .A(n4777), .ZN(n4780) );
  AOI22_X1 U5316 ( .A1(n2789), .A2(keyinput54), .B1(keyinput64), .B2(n4328), 
        .ZN(n4778) );
  OAI221_X1 U5317 ( .B1(n2789), .B2(keyinput54), .C1(n4328), .C2(keyinput64), 
        .A(n4778), .ZN(n4779) );
  NOR4_X1 U5318 ( .A1(n4782), .A2(n4781), .A3(n4780), .A4(n4779), .ZN(n4806)
         );
  AOI22_X1 U5319 ( .A1(n3113), .A2(keyinput73), .B1(n2255), .B2(keyinput40), 
        .ZN(n4783) );
  OAI221_X1 U5320 ( .B1(n3113), .B2(keyinput73), .C1(n2255), .C2(keyinput40), 
        .A(n4783), .ZN(n4791) );
  INV_X1 U5321 ( .A(REG2_REG_6__SCAN_IN), .ZN(n4785) );
  AOI22_X1 U5322 ( .A1(n4785), .A2(keyinput89), .B1(keyinput37), .B2(n4900), 
        .ZN(n4784) );
  OAI221_X1 U5323 ( .B1(n4785), .B2(keyinput89), .C1(n4900), .C2(keyinput37), 
        .A(n4784), .ZN(n4790) );
  AOI22_X1 U5324 ( .A1(n4605), .A2(keyinput53), .B1(n3419), .B2(keyinput93), 
        .ZN(n4786) );
  OAI221_X1 U5325 ( .B1(n4605), .B2(keyinput53), .C1(n3419), .C2(keyinput93), 
        .A(n4786), .ZN(n4789) );
  AOI22_X1 U5326 ( .A1(n4910), .A2(keyinput39), .B1(keyinput127), .B2(n4901), 
        .ZN(n4787) );
  OAI221_X1 U5327 ( .B1(n4910), .B2(keyinput39), .C1(n4901), .C2(keyinput127), 
        .A(n4787), .ZN(n4788) );
  NOR4_X1 U5328 ( .A1(n4791), .A2(n4790), .A3(n4789), .A4(n4788), .ZN(n4805)
         );
  INV_X1 U5329 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4793) );
  AOI22_X1 U5330 ( .A1(n4158), .A2(keyinput75), .B1(n4793), .B2(keyinput59), 
        .ZN(n4792) );
  OAI221_X1 U5331 ( .B1(n4158), .B2(keyinput75), .C1(n4793), .C2(keyinput59), 
        .A(n4792), .ZN(n4803) );
  INV_X1 U5332 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4795) );
  AOI22_X1 U5333 ( .A1(n4089), .A2(keyinput98), .B1(keyinput107), .B2(n4795), 
        .ZN(n4794) );
  OAI221_X1 U5334 ( .B1(n4089), .B2(keyinput98), .C1(n4795), .C2(keyinput107), 
        .A(n4794), .ZN(n4802) );
  AOI22_X1 U5335 ( .A1(n4078), .A2(keyinput66), .B1(keyinput17), .B2(n4797), 
        .ZN(n4796) );
  OAI221_X1 U5336 ( .B1(n4078), .B2(keyinput66), .C1(n4797), .C2(keyinput17), 
        .A(n4796), .ZN(n4801) );
  INV_X1 U5337 ( .A(ADDR_REG_12__SCAN_IN), .ZN(n4799) );
  INV_X1 U5338 ( .A(ADDR_REG_15__SCAN_IN), .ZN(n4905) );
  AOI22_X1 U5339 ( .A1(n4799), .A2(keyinput90), .B1(n4905), .B2(keyinput27), 
        .ZN(n4798) );
  OAI221_X1 U5340 ( .B1(n4799), .B2(keyinput90), .C1(n4905), .C2(keyinput27), 
        .A(n4798), .ZN(n4800) );
  NOR4_X1 U5341 ( .A1(n4803), .A2(n4802), .A3(n4801), .A4(n4800), .ZN(n4804)
         );
  NAND4_X1 U5342 ( .A1(n4807), .A2(n4806), .A3(n4805), .A4(n4804), .ZN(n4859)
         );
  INV_X1 U5343 ( .A(ADDR_REG_9__SCAN_IN), .ZN(n4809) );
  INV_X1 U5344 ( .A(ADDR_REG_10__SCAN_IN), .ZN(n4904) );
  AOI22_X1 U5345 ( .A1(n4809), .A2(keyinput5), .B1(n4904), .B2(keyinput86), 
        .ZN(n4808) );
  OAI221_X1 U5346 ( .B1(n4809), .B2(keyinput5), .C1(n4904), .C2(keyinput86), 
        .A(n4808), .ZN(n4817) );
  INV_X1 U5347 ( .A(ADDR_REG_4__SCAN_IN), .ZN(n4903) );
  AOI22_X1 U5348 ( .A1(n4903), .A2(keyinput124), .B1(keyinput20), .B2(n2934), 
        .ZN(n4810) );
  OAI221_X1 U5349 ( .B1(n4903), .B2(keyinput124), .C1(n2934), .C2(keyinput20), 
        .A(n4810), .ZN(n4816) );
  AOI22_X1 U5350 ( .A1(n2873), .A2(keyinput26), .B1(n4010), .B2(keyinput96), 
        .ZN(n4811) );
  OAI221_X1 U5351 ( .B1(n2873), .B2(keyinput26), .C1(n4010), .C2(keyinput96), 
        .A(n4811), .ZN(n4815) );
  INV_X1 U5352 ( .A(ADDR_REG_1__SCAN_IN), .ZN(n4813) );
  AOI22_X1 U5353 ( .A1(n2870), .A2(keyinput52), .B1(keyinput11), .B2(n4813), 
        .ZN(n4812) );
  OAI221_X1 U5354 ( .B1(n2870), .B2(keyinput52), .C1(n4813), .C2(keyinput11), 
        .A(n4812), .ZN(n4814) );
  NOR4_X1 U5355 ( .A1(n4817), .A2(n4816), .A3(n4815), .A4(n4814), .ZN(n4857)
         );
  AOI22_X1 U5356 ( .A1(n4919), .A2(keyinput105), .B1(n4920), .B2(keyinput82), 
        .ZN(n4818) );
  OAI221_X1 U5357 ( .B1(n4919), .B2(keyinput105), .C1(n4920), .C2(keyinput82), 
        .A(n4818), .ZN(n4829) );
  AOI22_X1 U5358 ( .A1(n4820), .A2(keyinput12), .B1(keyinput126), .B2(n4923), 
        .ZN(n4819) );
  OAI221_X1 U5359 ( .B1(n4820), .B2(keyinput12), .C1(n4923), .C2(keyinput126), 
        .A(n4819), .ZN(n4828) );
  AOI22_X1 U5360 ( .A1(n4924), .A2(keyinput1), .B1(keyinput77), .B2(n4822), 
        .ZN(n4821) );
  OAI221_X1 U5361 ( .B1(n4924), .B2(keyinput1), .C1(n4822), .C2(keyinput77), 
        .A(n4821), .ZN(n4827) );
  AOI22_X1 U5362 ( .A1(n4825), .A2(keyinput108), .B1(keyinput22), .B2(n4824), 
        .ZN(n4823) );
  OAI221_X1 U5363 ( .B1(n4825), .B2(keyinput108), .C1(n4824), .C2(keyinput22), 
        .A(n4823), .ZN(n4826) );
  NOR4_X1 U5364 ( .A1(n4829), .A2(n4828), .A3(n4827), .A4(n4826), .ZN(n4856)
         );
  AOI22_X1 U5365 ( .A1(n4922), .A2(keyinput19), .B1(keyinput119), .B2(n4921), 
        .ZN(n4830) );
  OAI221_X1 U5366 ( .B1(n4922), .B2(keyinput19), .C1(n4921), .C2(keyinput119), 
        .A(n4830), .ZN(n4840) );
  AOI22_X1 U5367 ( .A1(n4832), .A2(keyinput42), .B1(keyinput50), .B2(n4916), 
        .ZN(n4831) );
  OAI221_X1 U5368 ( .B1(n4832), .B2(keyinput42), .C1(n4916), .C2(keyinput50), 
        .A(n4831), .ZN(n4839) );
  AOI22_X1 U5369 ( .A1(n4834), .A2(keyinput45), .B1(n4917), .B2(keyinput3), 
        .ZN(n4833) );
  OAI221_X1 U5370 ( .B1(n4834), .B2(keyinput45), .C1(n4917), .C2(keyinput3), 
        .A(n4833), .ZN(n4838) );
  AOI22_X1 U5371 ( .A1(n4918), .A2(keyinput43), .B1(keyinput101), .B2(n4836), 
        .ZN(n4835) );
  OAI221_X1 U5372 ( .B1(n4918), .B2(keyinput43), .C1(n4836), .C2(keyinput101), 
        .A(n4835), .ZN(n4837) );
  NOR4_X1 U5373 ( .A1(n4840), .A2(n4839), .A3(n4838), .A4(n4837), .ZN(n4855)
         );
  AOI22_X1 U5374 ( .A1(n4843), .A2(keyinput115), .B1(keyinput95), .B2(n4842), 
        .ZN(n4841) );
  OAI221_X1 U5375 ( .B1(n4843), .B2(keyinput115), .C1(n4842), .C2(keyinput95), 
        .A(n4841), .ZN(n4853) );
  AOI22_X1 U5376 ( .A1(n4009), .A2(keyinput55), .B1(n4862), .B2(keyinput63), 
        .ZN(n4844) );
  OAI221_X1 U5377 ( .B1(n4009), .B2(keyinput55), .C1(n4862), .C2(keyinput63), 
        .A(n4844), .ZN(n4852) );
  AOI22_X1 U5378 ( .A1(n4863), .A2(keyinput69), .B1(n4846), .B2(keyinput92), 
        .ZN(n4845) );
  OAI221_X1 U5379 ( .B1(n4863), .B2(keyinput69), .C1(n4846), .C2(keyinput92), 
        .A(n4845), .ZN(n4851) );
  INV_X1 U5380 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4849) );
  AOI22_X1 U5381 ( .A1(n4849), .A2(keyinput71), .B1(n4848), .B2(keyinput110), 
        .ZN(n4847) );
  OAI221_X1 U5382 ( .B1(n4849), .B2(keyinput71), .C1(n4848), .C2(keyinput110), 
        .A(n4847), .ZN(n4850) );
  NOR4_X1 U5383 ( .A1(n4853), .A2(n4852), .A3(n4851), .A4(n4850), .ZN(n4854)
         );
  NAND4_X1 U5384 ( .A1(n4857), .A2(n4856), .A3(n4855), .A4(n4854), .ZN(n4858)
         );
  NOR4_X1 U5385 ( .A1(n4861), .A2(n4860), .A3(n4859), .A4(n4858), .ZN(n4941)
         );
  NAND4_X1 U5386 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_25__SCAN_IN), .A3(n4863), .A4(n4862), .ZN(n4939) );
  NAND4_X1 U5387 ( .A1(DATAI_27_), .A2(n4866), .A3(n4865), .A4(n4864), .ZN(
        n4867) );
  NOR3_X1 U5388 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .A3(n4867), 
        .ZN(n4882) );
  NAND4_X1 U5389 ( .A1(n4871), .A2(n4870), .A3(n4869), .A4(n4868), .ZN(n4880)
         );
  NAND4_X1 U5390 ( .A1(DATAI_19_), .A2(DATAI_21_), .A3(n4873), .A4(n4872), 
        .ZN(n4876) );
  INV_X1 U5391 ( .A(IR_REG_12__SCAN_IN), .ZN(n4874) );
  NAND4_X1 U5392 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .A3(
        IR_REG_7__SCAN_IN), .A4(n4874), .ZN(n4875) );
  OR4_X1 U5393 ( .A1(n4878), .A2(n4877), .A3(n4876), .A4(n4875), .ZN(n4879) );
  NOR4_X1 U5394 ( .A1(n4880), .A2(n4879), .A3(IR_REG_13__SCAN_IN), .A4(n2366), 
        .ZN(n4881) );
  NAND4_X1 U5395 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_26__SCAN_IN), .A3(n4882), .A4(n4881), .ZN(n4938) );
  NAND4_X1 U5396 ( .A1(REG0_REG_5__SCAN_IN), .A2(REG0_REG_14__SCAN_IN), .A3(
        REG0_REG_4__SCAN_IN), .A4(n4883), .ZN(n4889) );
  NAND4_X1 U5397 ( .A1(n4464), .A2(n4472), .A3(REG0_REG_20__SCAN_IN), .A4(
        REG0_REG_24__SCAN_IN), .ZN(n4888) );
  NAND4_X1 U5398 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_29__SCAN_IN), .A4(REG0_REG_0__SCAN_IN), .ZN(n4887) );
  NAND4_X1 U5399 ( .A1(n4885), .A2(n4884), .A3(REG0_REG_26__SCAN_IN), .A4(
        REG0_REG_11__SCAN_IN), .ZN(n4886) );
  NOR4_X1 U5400 ( .A1(n4889), .A2(n4888), .A3(n4887), .A4(n4886), .ZN(n4936)
         );
  NAND4_X1 U5401 ( .A1(REG3_REG_24__SCAN_IN), .A2(REG3_REG_25__SCAN_IN), .A3(
        REG3_REG_4__SCAN_IN), .A4(n2489), .ZN(n4898) );
  NAND4_X1 U5402 ( .A1(REG3_REG_27__SCAN_IN), .A2(DATAI_3_), .A3(DATAI_0_), 
        .A4(n4890), .ZN(n4891) );
  NOR2_X1 U5403 ( .A1(REG3_REG_21__SCAN_IN), .A2(n4891), .ZN(n4892) );
  NAND4_X1 U5404 ( .A1(n4893), .A2(D_REG_14__SCAN_IN), .A3(n2701), .A4(n4892), 
        .ZN(n4897) );
  INV_X1 U5405 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4895) );
  NAND4_X1 U5406 ( .A1(n4895), .A2(n4894), .A3(D_REG_0__SCAN_IN), .A4(
        D_REG_21__SCAN_IN), .ZN(n4896) );
  NOR3_X1 U5407 ( .A1(n4898), .A2(n4897), .A3(n4896), .ZN(n4935) );
  NOR4_X1 U5408 ( .A1(REG1_REG_27__SCAN_IN), .A2(REG1_REG_25__SCAN_IN), .A3(
        REG2_REG_6__SCAN_IN), .A4(n2255), .ZN(n4899) );
  NAND3_X1 U5409 ( .A1(REG2_REG_3__SCAN_IN), .A2(REG1_REG_31__SCAN_IN), .A3(
        n4899), .ZN(n4914) );
  NAND4_X1 U5410 ( .A1(REG2_REG_8__SCAN_IN), .A2(REG2_REG_24__SCAN_IN), .A3(
        n4901), .A4(n4900), .ZN(n4902) );
  NOR3_X1 U5411 ( .A1(REG2_REG_28__SCAN_IN), .A2(REG2_REG_21__SCAN_IN), .A3(
        n4902), .ZN(n4912) );
  NAND4_X1 U5412 ( .A1(REG1_REG_16__SCAN_IN), .A2(REG1_REG_20__SCAN_IN), .A3(
        REG1_REG_12__SCAN_IN), .A4(n4425), .ZN(n4909) );
  NAND4_X1 U5413 ( .A1(REG1_REG_6__SCAN_IN), .A2(REG1_REG_4__SCAN_IN), .A3(
        REG1_REG_3__SCAN_IN), .A4(REG0_REG_31__SCAN_IN), .ZN(n4908) );
  NAND4_X1 U5414 ( .A1(ADDR_REG_9__SCAN_IN), .A2(n4905), .A3(n4904), .A4(n4903), .ZN(n4907) );
  NAND4_X1 U5415 ( .A1(REG2_REG_27__SCAN_IN), .A2(ADDR_REG_16__SCAN_IN), .A3(
        ADDR_REG_12__SCAN_IN), .A4(n4078), .ZN(n4906) );
  NOR4_X1 U5416 ( .A1(n4909), .A2(n4908), .A3(n4907), .A4(n4906), .ZN(n4911)
         );
  NAND4_X1 U5417 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4912), .A3(n4911), .A4(
        n4910), .ZN(n4913) );
  NOR4_X1 U5418 ( .A1(REG1_REG_29__SCAN_IN), .A2(n4915), .A3(n4914), .A4(n4913), .ZN(n4934) );
  NAND4_X1 U5419 ( .A1(REG3_REG_15__SCAN_IN), .A2(REG3_REG_2__SCAN_IN), .A3(
        DATAO_REG_30__SCAN_IN), .A4(DATAO_REG_31__SCAN_IN), .ZN(n4931) );
  NAND4_X1 U5420 ( .A1(DATAO_REG_25__SCAN_IN), .A2(n4918), .A3(n4917), .A4(
        n4916), .ZN(n4930) );
  NOR4_X1 U5421 ( .A1(DATAO_REG_4__SCAN_IN), .A2(ADDR_REG_1__SCAN_IN), .A3(
        n4920), .A4(n4919), .ZN(n4928) );
  NOR4_X1 U5422 ( .A1(ADDR_REG_2__SCAN_IN), .A2(ADDR_REG_0__SCAN_IN), .A3(
        ADDR_REG_3__SCAN_IN), .A4(n2934), .ZN(n4927) );
  NOR4_X1 U5423 ( .A1(DATAO_REG_18__SCAN_IN), .A2(DATAO_REG_22__SCAN_IN), .A3(
        n4922), .A4(n4921), .ZN(n4926) );
  NOR4_X1 U5424 ( .A1(DATAO_REG_13__SCAN_IN), .A2(DATAO_REG_15__SCAN_IN), .A3(
        n4924), .A4(n4923), .ZN(n4925) );
  NAND4_X1 U5425 ( .A1(n4928), .A2(n4927), .A3(n4926), .A4(n4925), .ZN(n4929)
         );
  NOR4_X1 U5426 ( .A1(n4932), .A2(n4931), .A3(n4930), .A4(n4929), .ZN(n4933)
         );
  NAND4_X1 U5427 ( .A1(n4936), .A2(n4935), .A3(n4934), .A4(n4933), .ZN(n4937)
         );
  NOR4_X1 U5428 ( .A1(REG2_REG_26__SCAN_IN), .A2(n4939), .A3(n4938), .A4(n4937), .ZN(n4940) );
  XOR2_X1 U5429 ( .A(n4941), .B(n4940), .Z(n4944) );
  NAND2_X1 U5430 ( .A1(D_REG_12__SCAN_IN), .A2(n4942), .ZN(n4943) );
  XNOR2_X1 U5431 ( .A(n4944), .B(n4943), .ZN(U3310) );
endmodule

