

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput0, keyinput1, keyinput2, 
        keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, 
        keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, 
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, 
        keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, 
        keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, 
        keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, 
        keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, 
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, 
        keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, 
        keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, 
        keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, 
        keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, 
        keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, 
        keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, 
        keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, 
        keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, 
        keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, 
        keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, 
        keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, 
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, 
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, 
        keyinput124, keyinput125, keyinput126, keyinput127 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127;

  NOR2_X1 U3532 ( .A1(n5692), .A2(n5691), .ZN(n5693) );
  NAND2_X1 U3533 ( .A1(n3162), .A2(n3161), .ZN(n4884) );
  NAND2_X1 U3534 ( .A1(n3431), .A2(n3430), .ZN(n4324) );
  CLKBUF_X2 U3535 ( .A(n3487), .Z(n3086) );
  CLKBUF_X2 U3536 ( .A(n4075), .Z(n5124) );
  CLKBUF_X2 U3537 ( .A(n3497), .Z(n5115) );
  AND2_X1 U3539 ( .A1(n4492), .A2(n4315), .ZN(n3497) );
  AND2_X1 U3540 ( .A1(n3395), .A2(n3748), .ZN(n3148) );
  NAND2_X1 U3541 ( .A1(n3208), .A2(n3123), .ZN(n3653) );
  NAND2_X1 U3542 ( .A1(n4406), .A2(n5200), .ZN(n3771) );
  INV_X2 U3543 ( .A(n3290), .ZN(n4168) );
  INV_X1 U3544 ( .A(n3153), .ZN(n3851) );
  AND2_X2 U3545 ( .A1(n3299), .A2(n4315), .ZN(n3487) );
  OR2_X1 U3546 ( .A1(n5048), .A2(n5389), .ZN(n3251) );
  INV_X2 U3547 ( .A(n5813), .ZN(n5815) );
  INV_X1 U3548 ( .A(n3764), .ZN(n4991) );
  INV_X1 U3549 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6673) );
  INV_X1 U3551 ( .A(n6422), .ZN(n6435) );
  INV_X1 U3552 ( .A(n6451), .ZN(n6440) );
  AND4_X1 U3553 ( .A1(n3382), .A2(n3381), .A3(n3380), .A4(n3379), .ZN(n3084)
         );
  NAND2_X2 U3555 ( .A1(n3653), .A2(n3652), .ZN(n3659) );
  INV_X2 U3556 ( .A(n3912), .ZN(n6071) );
  NAND2_X2 U3557 ( .A1(n3314), .A2(n3099), .ZN(n3384) );
  NAND2_X2 U3559 ( .A1(n3150), .A2(n3199), .ZN(n5747) );
  OAI21_X4 U3560 ( .B1(n3729), .B2(n3735), .A(n3219), .ZN(n4376) );
  NOR2_X1 U3561 ( .A1(n4884), .A2(n3233), .ZN(n5377) );
  AOI21_X2 U3562 ( .B1(n5674), .B2(n5864), .A(n5236), .ZN(n5225) );
  AND2_X1 U3563 ( .A1(n5711), .A2(n5223), .ZN(n5699) );
  AOI21_X1 U3564 ( .B1(n5049), .B2(n5278), .A(n5056), .ZN(n4995) );
  INV_X4 U3565 ( .A(n5813), .ZN(n5824) );
  NOR3_X2 U3566 ( .A1(n5286), .A2(n4992), .A3(n3289), .ZN(n5048) );
  AND2_X1 U3567 ( .A1(n5303), .A2(n5304), .ZN(n5306) );
  INV_X1 U3568 ( .A(n3749), .ZN(n3386) );
  NOR2_X1 U3569 ( .A1(n4719), .A2(n3894), .ZN(n3839) );
  NOR2_X2 U3570 ( .A1(n3764), .A2(n5050), .ZN(n3763) );
  OR2_X1 U3571 ( .A1(n3405), .A2(n4531), .ZN(n3529) );
  OR2_X2 U3572 ( .A1(n3344), .A2(n3343), .ZN(n3400) );
  AND2_X1 U3573 ( .A1(n3157), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4319)
         );
  AND2_X1 U3574 ( .A1(n5879), .A2(n6653), .ZN(n3191) );
  NOR2_X1 U3575 ( .A1(n5764), .A2(n3137), .ZN(n5768) );
  NOR2_X1 U3576 ( .A1(n5032), .A2(n3277), .ZN(n3276) );
  AOI21_X1 U3577 ( .B1(n5267), .B2(n5839), .A(n5252), .ZN(n5253) );
  OAI21_X1 U3578 ( .B1(n5490), .B2(n5489), .A(n5488), .ZN(n5802) );
  AND2_X1 U3579 ( .A1(n5810), .A2(n5842), .ZN(n5834) );
  NOR2_X1 U3580 ( .A1(n5486), .A2(n5453), .ZN(n5487) );
  XNOR2_X1 U3581 ( .A(n5657), .B(n5454), .ZN(n5486) );
  AOI21_X1 U3582 ( .B1(n3184), .B2(n3183), .A(n3182), .ZN(n3181) );
  NOR2_X1 U3583 ( .A1(n6462), .A2(n5677), .ZN(n3227) );
  AND2_X1 U3584 ( .A1(n5452), .A2(n5451), .ZN(n5657) );
  INV_X2 U3585 ( .A(n6427), .ZN(n6462) );
  AND2_X1 U3586 ( .A1(n5377), .A2(n5594), .ZN(n5452) );
  AND2_X1 U3587 ( .A1(n5842), .A2(n3665), .ZN(n3666) );
  NOR2_X1 U3588 ( .A1(n3270), .A2(n3102), .ZN(n3268) );
  AND2_X1 U3589 ( .A1(n5809), .A2(n3661), .ZN(n3662) );
  AND2_X1 U3590 ( .A1(n5814), .A2(n3664), .ZN(n3665) );
  AND2_X1 U3591 ( .A1(n3113), .A2(n3667), .ZN(n3271) );
  AND2_X1 U3592 ( .A1(n4768), .A2(n4771), .ZN(n3161) );
  INV_X1 U3593 ( .A(n4769), .ZN(n3162) );
  AND2_X1 U3594 ( .A1(n5903), .A2(n5232), .ZN(n5871) );
  AND2_X1 U3595 ( .A1(n5881), .A2(n5228), .ZN(n5861) );
  NOR2_X1 U3596 ( .A1(n5278), .A2(n5277), .ZN(n5863) );
  NAND2_X1 U3597 ( .A1(n3647), .A2(n3646), .ZN(n3650) );
  NAND2_X1 U3598 ( .A1(n3938), .A2(n3937), .ZN(n4768) );
  NAND2_X1 U3599 ( .A1(n4462), .A2(n3931), .ZN(n4769) );
  INV_X1 U3600 ( .A(n4885), .ZN(n3235) );
  AND2_X1 U3601 ( .A1(n4533), .A2(n4883), .ZN(n3931) );
  AND2_X1 U3602 ( .A1(n5899), .A2(n5226), .ZN(n5881) );
  XNOR2_X1 U3603 ( .A(n3653), .B(n3118), .ZN(n3946) );
  OAI211_X1 U3604 ( .C1(n6582), .C2(INSTADDRPOINTER_REG_3__SCAN_IN), .A(n4588), 
        .B(n3571), .ZN(n3572) );
  NAND2_X1 U3605 ( .A1(n5306), .A2(n4986), .ZN(n5286) );
  NOR2_X1 U3606 ( .A1(n6203), .A2(n6056), .ZN(n4853) );
  XNOR2_X1 U3607 ( .A(n3615), .B(n3617), .ZN(n3890) );
  CLKBUF_X1 U3608 ( .A(n4542), .Z(n4583) );
  OR2_X1 U3609 ( .A1(n6026), .A2(n3876), .ZN(n5959) );
  AND2_X1 U3610 ( .A1(n5380), .A2(n3832), .ZN(n5373) );
  AND2_X1 U3611 ( .A1(n6203), .A2(n6071), .ZN(n6246) );
  NOR2_X1 U3612 ( .A1(n5394), .A2(n5428), .ZN(n5380) );
  OR2_X1 U3613 ( .A1(n4342), .A2(n4341), .ZN(n4344) );
  NAND2_X1 U3614 ( .A1(n6041), .A2(n6038), .ZN(n5967) );
  AND2_X1 U3615 ( .A1(n6004), .A2(n4352), .ZN(n6041) );
  AND2_X1 U3616 ( .A1(n3870), .A2(n3845), .ZN(n6636) );
  XNOR2_X1 U3617 ( .A(n4324), .B(n4780), .ZN(n4491) );
  OAI21_X1 U3618 ( .B1(n3915), .B2(STATE2_REG_0__SCAN_IN), .A(n3509), .ZN(
        n3197) );
  NOR2_X1 U3619 ( .A1(n3259), .A2(n3258), .ZN(n3257) );
  AOI21_X1 U3620 ( .B1(n4281), .B2(n3393), .A(n3839), .ZN(n3388) );
  NAND2_X1 U3621 ( .A1(n3770), .A2(n3769), .ZN(n3774) );
  AND2_X1 U3622 ( .A1(n3397), .A2(n3859), .ZN(n3417) );
  AND2_X2 U3623 ( .A1(n3386), .A2(n3385), .ZN(n3739) );
  NAND2_X1 U3624 ( .A1(n3407), .A2(n4531), .ZN(n3158) );
  NAND2_X1 U3625 ( .A1(n3288), .A2(n4279), .ZN(n4719) );
  AND2_X2 U3626 ( .A1(n3405), .A2(n3406), .ZN(n3713) );
  AND2_X2 U3627 ( .A1(n4413), .A2(n5200), .ZN(n5197) );
  AND2_X1 U3628 ( .A1(n4373), .A2(n3400), .ZN(n3391) );
  NAND2_X2 U3629 ( .A1(n3396), .A2(n5200), .ZN(n3764) );
  AND3_X2 U3630 ( .A1(n3210), .A2(n3212), .A3(n3211), .ZN(n3153) );
  INV_X2 U3631 ( .A(n5200), .ZN(n3410) );
  OR2_X2 U3632 ( .A1(n3305), .A2(n3304), .ZN(n3398) );
  AND3_X1 U3633 ( .A1(n3349), .A2(n3352), .A3(n3350), .ZN(n3210) );
  AND4_X1 U3634 ( .A1(n3378), .A2(n3377), .A3(n3376), .A4(n3375), .ZN(n3383)
         );
  AND2_X1 U3635 ( .A1(n3156), .A2(n3154), .ZN(n3349) );
  AND3_X1 U3636 ( .A1(n3348), .A2(n3351), .A3(n3347), .ZN(n3212) );
  AND4_X1 U3637 ( .A1(n3318), .A2(n3317), .A3(n3316), .A4(n3315), .ZN(n3334)
         );
  AND2_X1 U3638 ( .A1(n3346), .A2(n3353), .ZN(n3211) );
  AND4_X1 U3639 ( .A1(n3309), .A2(n3308), .A3(n3307), .A4(n3306), .ZN(n3314)
         );
  AND4_X1 U3640 ( .A1(n3326), .A2(n3325), .A3(n3324), .A4(n3323), .ZN(n3332)
         );
  BUF_X2 U3641 ( .A(n3495), .Z(n3496) );
  BUF_X2 U3642 ( .A(n3484), .Z(n5122) );
  BUF_X2 U3643 ( .A(n3460), .Z(n5107) );
  AND2_X2 U3644 ( .A1(n3298), .A2(n4315), .ZN(n4075) );
  AND2_X2 U3645 ( .A1(n3298), .A2(n3297), .ZN(n5116) );
  AND2_X2 U3646 ( .A1(n3297), .A2(n4492), .ZN(n3467) );
  BUF_X2 U3647 ( .A(n5007), .Z(n3088) );
  AND2_X2 U3648 ( .A1(n4319), .A2(n3299), .ZN(n3484) );
  AND2_X2 U3649 ( .A1(n4319), .A2(n4492), .ZN(n3485) );
  BUF_X2 U3650 ( .A(n3535), .Z(n5114) );
  BUF_X4 U3651 ( .A(n5007), .Z(n3087) );
  AND2_X2 U3652 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4315) );
  NOR2_X2 U3653 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4314) );
  NOR2_X4 U3654 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4492) );
  INV_X1 U3655 ( .A(n3907), .ZN(n6056) );
  OAI211_X1 U3656 ( .C1(n5613), .C2(n6435), .A(n3228), .B(n3224), .ZN(n3223)
         );
  NAND2_X2 U3657 ( .A1(n3930), .A2(n3929), .ZN(n4462) );
  NAND2_X1 U3658 ( .A1(n4717), .A2(n3400), .ZN(n3401) );
  NAND2_X1 U3659 ( .A1(n4717), .A2(n3745), .ZN(n3759) );
  NOR2_X4 U3660 ( .A1(n3387), .A2(n3398), .ZN(n3404) );
  NOR2_X4 U3661 ( .A1(n3869), .A2(n3374), .ZN(n3752) );
  NAND3_X2 U3662 ( .A1(n3386), .A2(n3411), .A3(n3851), .ZN(n3869) );
  AND4_X2 U3663 ( .A1(n3145), .A2(n3144), .A3(INSTQUEUERD_ADDR_REG_1__SCAN_IN), 
        .A4(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5007) );
  AND2_X1 U3664 ( .A1(n5251), .A2(n5188), .ZN(n3090) );
  NOR2_X2 U3665 ( .A1(n6263), .A2(n6262), .ZN(n6292) );
  AOI21_X4 U3666 ( .B1(n3907), .B2(n3710), .A(n3521), .ZN(n6578) );
  NOR2_X4 U3667 ( .A1(n5148), .A2(n5147), .ZN(n5323) );
  AND2_X2 U3668 ( .A1(n4314), .A2(n4492), .ZN(n3489) );
  AND2_X2 U3669 ( .A1(n4314), .A2(n3165), .ZN(n3535) );
  NAND2_X4 U3670 ( .A1(n3519), .A2(n3396), .ZN(n5050) );
  NAND2_X4 U3671 ( .A1(n3383), .A2(n3084), .ZN(n3396) );
  AND2_X1 U3672 ( .A1(n3115), .A2(n3672), .ZN(n3213) );
  INV_X1 U3673 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3155) );
  AND2_X1 U3674 ( .A1(n3630), .A2(n3629), .ZN(n3631) );
  NAND2_X1 U3675 ( .A1(n4581), .A2(n3209), .ZN(n3615) );
  NOR2_X1 U3676 ( .A1(n5447), .A2(n5208), .ZN(n5399) );
  NAND2_X1 U3677 ( .A1(n3235), .A2(n3231), .ZN(n3230) );
  AND2_X1 U3678 ( .A1(n3234), .A2(n3232), .ZN(n3231) );
  OR2_X1 U3679 ( .A1(n3400), .A2(n6673), .ZN(n3290) );
  INV_X1 U3680 ( .A(n5286), .ZN(n5051) );
  OAI21_X1 U3681 ( .B1(n3185), .B2(n5800), .A(n3181), .ZN(n3673) );
  INV_X1 U3682 ( .A(n5801), .ZN(n3183) );
  NAND2_X1 U3683 ( .A1(n3946), .A2(n3710), .ZN(n3647) );
  AND2_X1 U3684 ( .A1(n3151), .A2(n3387), .ZN(n3288) );
  OR2_X1 U3685 ( .A1(n5312), .A2(n3111), .ZN(n5195) );
  NAND2_X1 U3686 ( .A1(n5863), .A2(n6451), .ZN(n3226) );
  OR3_X1 U3687 ( .A1(n6808), .A2(n6577), .A3(n5044), .ZN(n6423) );
  AND2_X1 U3688 ( .A1(n6423), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5517) );
  INV_X1 U3689 ( .A(n5180), .ZN(n5060) );
  NAND2_X1 U3690 ( .A1(n3173), .A2(n3105), .ZN(n4715) );
  NAND2_X1 U3691 ( .A1(n3729), .A2(n3219), .ZN(n3173) );
  NAND2_X1 U3692 ( .A1(n3219), .A2(n3735), .ZN(n3218) );
  NOR2_X1 U3693 ( .A1(n5747), .A2(n3204), .ZN(n5236) );
  NAND2_X1 U3694 ( .A1(n3207), .A2(n3130), .ZN(n3204) );
  INV_X1 U3695 ( .A(n5224), .ZN(n3207) );
  NAND2_X1 U3696 ( .A1(n3282), .A2(n3281), .ZN(n3180) );
  INV_X1 U3697 ( .A(n5750), .ZN(n3281) );
  NAND2_X1 U3698 ( .A1(n5824), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3137) );
  AND4_X1 U3699 ( .A1(n3322), .A2(n3321), .A3(n3320), .A4(n3319), .ZN(n3333)
         );
  AND4_X1 U3700 ( .A1(n3330), .A2(n3329), .A3(n3328), .A4(n3327), .ZN(n3331)
         );
  NAND2_X1 U3701 ( .A1(n3479), .A2(n3480), .ZN(n3483) );
  AND2_X2 U3702 ( .A1(n3139), .A2(n3574), .ZN(n3907) );
  INV_X1 U3703 ( .A(n3141), .ZN(n3140) );
  INV_X1 U3704 ( .A(n3143), .ZN(n3142) );
  AND2_X1 U3705 ( .A1(n4673), .A2(n4604), .ZN(n6212) );
  INV_X2 U3706 ( .A(n3405), .ZN(n4717) );
  INV_X1 U3707 ( .A(n6651), .ZN(n6640) );
  INV_X1 U3708 ( .A(n3201), .ZN(n3182) );
  INV_X1 U3709 ( .A(n3631), .ZN(n3196) );
  OR2_X1 U3710 ( .A1(n3584), .A2(n3583), .ZN(n3634) );
  NAND2_X1 U3711 ( .A1(n3771), .A2(EBX_REG_1__SCAN_IN), .ZN(n3240) );
  NAND2_X2 U3712 ( .A1(n3530), .A2(n3529), .ZN(n3730) );
  AND2_X1 U3713 ( .A1(n5282), .A2(n3239), .ZN(n3238) );
  AND2_X1 U3714 ( .A1(n5296), .A2(n5309), .ZN(n3239) );
  AND2_X1 U3715 ( .A1(n4174), .A2(n5600), .ZN(n3234) );
  AND2_X1 U3716 ( .A1(n5378), .A2(n4173), .ZN(n4174) );
  NAND2_X1 U3717 ( .A1(n3975), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3992)
         );
  NAND2_X1 U3718 ( .A1(n3755), .A2(n3410), .ZN(n3747) );
  NOR2_X1 U3719 ( .A1(n3836), .A2(n3263), .ZN(n3262) );
  INV_X1 U3720 ( .A(n5372), .ZN(n3263) );
  INV_X1 U3721 ( .A(n5849), .ZN(n3134) );
  INV_X1 U3722 ( .A(n6565), .ZN(n3135) );
  NAND2_X1 U3723 ( .A1(n3244), .A2(n5587), .ZN(n3243) );
  INV_X1 U3724 ( .A(n3245), .ZN(n3244) );
  OR2_X1 U3725 ( .A1(n5602), .A2(n5596), .ZN(n3245) );
  INV_X1 U3726 ( .A(n3098), .ZN(n4987) );
  NAND2_X1 U3727 ( .A1(n3786), .A2(n3256), .ZN(n3259) );
  INV_X1 U3728 ( .A(n4667), .ZN(n3256) );
  OR2_X1 U3729 ( .A1(n3541), .A2(n3540), .ZN(n3587) );
  XNOR2_X1 U3730 ( .A(n3445), .B(n3444), .ZN(n3141) );
  AND2_X1 U3731 ( .A1(n3151), .A2(n3410), .ZN(n3860) );
  INV_X1 U3732 ( .A(n3220), .ZN(n3219) );
  NAND2_X1 U3733 ( .A1(n3737), .A2(n3736), .ZN(n3738) );
  NAND2_X1 U3734 ( .A1(n3498), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3156)
         );
  NAND2_X1 U3735 ( .A1(n3460), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3154) );
  INV_X1 U3736 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4839) );
  OR2_X2 U3737 ( .A1(n3363), .A2(n3362), .ZN(n3519) );
  NAND2_X1 U3738 ( .A1(n5341), .A2(n5193), .ZN(n5312) );
  NAND2_X1 U3739 ( .A1(n6459), .A2(n3128), .ZN(n5448) );
  NAND2_X1 U3740 ( .A1(n5491), .A2(n3129), .ZN(n5447) );
  AND2_X1 U3741 ( .A1(n6459), .A2(n5206), .ZN(n6389) );
  INV_X1 U3742 ( .A(n5325), .ZN(n5147) );
  INV_X1 U3743 ( .A(n5184), .ZN(n5274) );
  NAND2_X1 U3744 ( .A1(n5323), .A2(n5309), .ZN(n5308) );
  AND2_X1 U3745 ( .A1(n5323), .A2(n3239), .ZN(n5294) );
  NAND2_X1 U3746 ( .A1(n5142), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5159)
         );
  NAND2_X1 U3747 ( .A1(n5353), .A2(n4236), .ZN(n5021) );
  NAND2_X1 U3748 ( .A1(n4154), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4189)
         );
  INV_X1 U3749 ( .A(n4155), .ZN(n4154) );
  NAND2_X1 U3750 ( .A1(n3235), .A2(n5600), .ZN(n3233) );
  NAND2_X1 U3751 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n3949), .ZN(n3971)
         );
  AND2_X1 U3752 ( .A1(n3920), .A2(n3919), .ZN(n4341) );
  AND2_X1 U3753 ( .A1(n5051), .A2(n5275), .ZN(n5278) );
  NAND2_X1 U3754 ( .A1(n3215), .A2(n3107), .ZN(n5683) );
  NOR2_X1 U3755 ( .A1(n3200), .A2(n3674), .ZN(n3280) );
  AND2_X1 U3756 ( .A1(n5824), .A2(n5935), .ZN(n3674) );
  AOI21_X1 U3757 ( .B1(n3201), .B2(n3203), .A(n3200), .ZN(n3199) );
  NAND2_X1 U3758 ( .A1(n3814), .A2(n3252), .ZN(n5428) );
  NOR2_X1 U3759 ( .A1(n3253), .A2(n3122), .ZN(n3252) );
  INV_X1 U3760 ( .A(n3254), .ZN(n3253) );
  NAND2_X1 U3761 ( .A1(n3668), .A2(n3271), .ZN(n3269) );
  NAND2_X1 U3762 ( .A1(n5800), .A2(n5801), .ZN(n3668) );
  OR2_X1 U3763 ( .A1(n4304), .A2(n3844), .ZN(n4473) );
  NAND2_X1 U3764 ( .A1(n3166), .A2(n3408), .ZN(n3479) );
  NAND2_X1 U3765 ( .A1(n3197), .A2(n3556), .ZN(n3560) );
  OAI21_X1 U3766 ( .B1(n3507), .B2(n4531), .A(n3557), .ZN(n3508) );
  INV_X1 U3767 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4495) );
  NOR2_X1 U3768 ( .A1(n6203), .A2(n3907), .ZN(n4669) );
  AND2_X1 U3769 ( .A1(n4394), .A2(n4531), .ZN(n4673) );
  NAND2_X1 U3770 ( .A1(n6061), .A2(n4393), .ZN(n4394) );
  INV_X1 U3771 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6304) );
  INV_X1 U3772 ( .A(n3519), .ZN(n4406) );
  NAND2_X1 U3773 ( .A1(n3172), .A2(n4281), .ZN(n5040) );
  INV_X1 U3774 ( .A(n4715), .ZN(n3172) );
  INV_X1 U3775 ( .A(n5195), .ZN(n5288) );
  NOR2_X1 U3776 ( .A1(n3227), .A2(n3225), .ZN(n3224) );
  NAND2_X1 U3777 ( .A1(n3226), .A2(n5280), .ZN(n3225) );
  INV_X1 U3778 ( .A(n5211), .ZN(n3216) );
  AND2_X1 U3779 ( .A1(n6459), .A2(n3127), .ZN(n5476) );
  NAND2_X1 U3780 ( .A1(n6459), .A2(n3126), .ZN(n6384) );
  NOR2_X2 U3781 ( .A1(n5251), .A2(n5187), .ZN(n6422) );
  INV_X1 U3782 ( .A(n5243), .ZN(n5265) );
  AND2_X1 U3783 ( .A1(n5664), .A2(n4728), .ZN(n5645) );
  AND2_X1 U3784 ( .A1(n5664), .A2(n4729), .ZN(n5646) );
  NAND2_X1 U3785 ( .A1(n6362), .A2(n4239), .ZN(n5853) );
  INV_X1 U3786 ( .A(n6599), .ZN(n5855) );
  INV_X1 U3787 ( .A(n5853), .ZN(n6591) );
  NAND2_X1 U3788 ( .A1(n5055), .A2(n3249), .ZN(n5270) );
  INV_X1 U3789 ( .A(n5052), .ZN(n5053) );
  AOI21_X1 U3790 ( .B1(n5237), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5229), 
        .ZN(n3248) );
  OAI211_X1 U3791 ( .C1(n5681), .C2(n5875), .A(n3193), .B(n3192), .ZN(n5879)
         );
  NAND2_X1 U3792 ( .A1(n5681), .A2(n5682), .ZN(n3192) );
  INV_X1 U3793 ( .A(n3194), .ZN(n3193) );
  OAI21_X1 U3794 ( .B1(n5692), .B2(n3195), .A(n5683), .ZN(n3194) );
  NAND2_X1 U3795 ( .A1(n3274), .A2(n3272), .ZN(n3889) );
  NAND2_X1 U3796 ( .A1(n3276), .A2(n3273), .ZN(n3272) );
  AND2_X1 U3797 ( .A1(n3093), .A2(n5032), .ZN(n3275) );
  AOI21_X1 U3798 ( .B1(n3169), .B2(n3095), .A(n3125), .ZN(n3170) );
  AND2_X1 U3799 ( .A1(n3870), .A2(n3841), .ZN(n6651) );
  AND2_X1 U3800 ( .A1(n3870), .A2(n3762), .ZN(n6653) );
  CLKBUF_X1 U3801 ( .A(n4491), .Z(n6206) );
  INV_X1 U3802 ( .A(n6804), .ZN(n6663) );
  OR2_X1 U3803 ( .A1(n3604), .A2(n3603), .ZN(n3633) );
  INV_X1 U3804 ( .A(n3518), .ZN(n3543) );
  CLKBUF_X2 U3805 ( .A(n3489), .Z(n3461) );
  NAND2_X1 U3806 ( .A1(n5200), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3701) );
  OAI21_X1 U3807 ( .B1(n3177), .B2(n3176), .A(n3716), .ZN(n3175) );
  INV_X1 U3808 ( .A(n3713), .ZN(n3727) );
  INV_X1 U3809 ( .A(n3734), .ZN(n3737) );
  AND2_X1 U3810 ( .A1(n5410), .A2(n4153), .ZN(n5395) );
  AND2_X1 U3811 ( .A1(n5425), .A2(n5423), .ZN(n5410) );
  NAND2_X1 U3812 ( .A1(n3208), .A2(n3618), .ZN(n3632) );
  AOI21_X1 U3813 ( .B1(n3907), .B2(n4116), .A(n5245), .ZN(n3926) );
  INV_X1 U3814 ( .A(n3268), .ZN(n3202) );
  OR2_X1 U3815 ( .A1(n5776), .A2(n3138), .ZN(n5764) );
  NOR2_X1 U3816 ( .A1(n5813), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3138)
         );
  NAND2_X1 U3817 ( .A1(n3269), .A2(n3268), .ZN(n5756) );
  NOR2_X1 U3818 ( .A1(n3109), .A2(n5492), .ZN(n3254) );
  INV_X1 U3819 ( .A(n6041), .ZN(n4593) );
  NAND2_X1 U3820 ( .A1(n3410), .A2(n3519), .ZN(n3561) );
  OAI21_X1 U3821 ( .B1(n3763), .B2(EBX_REG_1__SCAN_IN), .A(n3240), .ZN(n3770)
         );
  AND2_X1 U3822 ( .A1(n3745), .A2(n3396), .ZN(n3710) );
  OR2_X1 U3823 ( .A1(n3504), .A2(n3503), .ZN(n3562) );
  OR2_X1 U3824 ( .A1(n3475), .A2(n3474), .ZN(n3654) );
  NAND2_X1 U3825 ( .A1(n4310), .A2(n4531), .ZN(n3131) );
  OR2_X1 U3826 ( .A1(n4376), .A2(n3844), .ZN(n4307) );
  NAND2_X1 U3827 ( .A1(n4491), .A2(n4531), .ZN(n3186) );
  OR2_X1 U3828 ( .A1(n5192), .A2(n5556), .ZN(n5341) );
  NOR2_X1 U3829 ( .A1(n5420), .A2(n5209), .ZN(n5384) );
  INV_X1 U3830 ( .A(n5498), .ZN(n3221) );
  NOR2_X1 U3831 ( .A1(n6386), .A2(n5191), .ZN(n5491) );
  OR2_X1 U3832 ( .A1(n6458), .A2(n5205), .ZN(n6386) );
  INV_X1 U3833 ( .A(n3404), .ZN(n4726) );
  NOR2_X1 U3834 ( .A1(n5274), .A2(n3237), .ZN(n3236) );
  INV_X1 U3835 ( .A(n3238), .ZN(n3237) );
  NAND2_X1 U3836 ( .A1(n5059), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5180)
         );
  NAND2_X1 U3837 ( .A1(n5323), .A2(n3238), .ZN(n5281) );
  OR3_X1 U3838 ( .A1(n5159), .A2(n5701), .A3(n5158), .ZN(n5171) );
  AND2_X1 U3839 ( .A1(n5058), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5142)
         );
  INV_X1 U3840 ( .A(n5057), .ZN(n5058) );
  NAND2_X1 U3841 ( .A1(n4231), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5057)
         );
  NAND2_X1 U3842 ( .A1(n4188), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4229)
         );
  NAND2_X1 U3843 ( .A1(n3235), .A2(n3234), .ZN(n3229) );
  OR2_X1 U3844 ( .A1(n4137), .A2(n3977), .ZN(n4155) );
  NAND2_X1 U3845 ( .A1(n4036), .A2(n3974), .ZN(n4122) );
  AND2_X1 U3846 ( .A1(n4100), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4074)
         );
  NAND2_X1 U3847 ( .A1(n3972), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4107)
         );
  NOR2_X1 U3848 ( .A1(n3948), .A2(n3947), .ZN(n3949) );
  INV_X1 U3849 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3947) );
  AOI21_X1 U3850 ( .B1(n3946), .B2(n4116), .A(n3955), .ZN(n4885) );
  NOR2_X1 U3851 ( .A1(n3900), .A2(n3891), .ZN(n3933) );
  INV_X1 U3852 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3891) );
  INV_X1 U3853 ( .A(n3922), .ZN(n3901) );
  NAND2_X1 U3854 ( .A1(n3901), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3900)
         );
  NAND2_X1 U3855 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3922) );
  OR2_X1 U3856 ( .A1(n5048), .A2(n5286), .ZN(n3250) );
  NAND2_X1 U3857 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n5869), .ZN(n3195) );
  AND2_X1 U3858 ( .A1(n3092), .A2(n3261), .ZN(n3260) );
  INV_X1 U3859 ( .A(n5319), .ZN(n3261) );
  NAND2_X1 U3860 ( .A1(n5373), .A2(n3092), .ZN(n5320) );
  NAND2_X1 U3861 ( .A1(n5373), .A2(n3262), .ZN(n5349) );
  INV_X1 U3862 ( .A(n3675), .ZN(n3277) );
  NOR2_X1 U3863 ( .A1(n3675), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3278)
         );
  AND2_X1 U3864 ( .A1(n5373), .A2(n5372), .ZN(n5370) );
  NAND2_X1 U3865 ( .A1(n5731), .A2(n5730), .ZN(n5729) );
  AND2_X1 U3866 ( .A1(n3766), .A2(n3765), .ZN(n5394) );
  NOR2_X1 U3867 ( .A1(n5815), .A2(n5935), .ZN(n5750) );
  INV_X1 U3868 ( .A(n5764), .ZN(n3169) );
  NAND2_X1 U3869 ( .A1(n5756), .A2(n3670), .ZN(n5776) );
  NAND2_X1 U3870 ( .A1(n3814), .A2(n3254), .ZN(n5461) );
  NAND2_X1 U3871 ( .A1(n3662), .A2(n3134), .ZN(n3133) );
  NAND2_X1 U3872 ( .A1(n3662), .A2(n3651), .ZN(n3136) );
  AND2_X1 U3873 ( .A1(n6636), .A2(n3883), .ZN(n5983) );
  NAND2_X1 U3874 ( .A1(n3241), .A2(n3108), .ZN(n6016) );
  INV_X1 U3875 ( .A(n3243), .ZN(n3242) );
  NOR2_X1 U3876 ( .A1(n5603), .A2(n3243), .ZN(n5589) );
  NOR2_X1 U3877 ( .A1(n5603), .A2(n3245), .ZN(n5595) );
  AND2_X1 U3878 ( .A1(n3800), .A2(n3799), .ZN(n5602) );
  NAND2_X1 U3879 ( .A1(n6565), .A2(n3651), .ZN(n5850) );
  INV_X1 U3880 ( .A(n6636), .ZN(n6038) );
  INV_X1 U3881 ( .A(n4775), .ZN(n3258) );
  NAND2_X1 U3882 ( .A1(n3178), .A2(n3614), .ZN(n3266) );
  NAND2_X1 U3883 ( .A1(n3787), .A2(n3287), .ZN(n4667) );
  NOR2_X1 U3884 ( .A1(n5536), .A2(n3259), .ZN(n4776) );
  NAND2_X1 U3885 ( .A1(n3523), .A2(n6582), .ZN(n3146) );
  OR2_X1 U3886 ( .A1(n5536), .A2(n4537), .ZN(n4666) );
  NAND2_X1 U3887 ( .A1(n4960), .A2(n4593), .ZN(n6628) );
  NAND2_X1 U3888 ( .A1(n4382), .A2(n4991), .ZN(n4381) );
  NAND2_X1 U3889 ( .A1(n3164), .A2(n3429), .ZN(n3163) );
  CLKBUF_X1 U3890 ( .A(n4315), .Z(n4943) );
  AND2_X2 U3891 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3165) );
  AND2_X1 U3892 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4496) );
  NAND2_X1 U3893 ( .A1(n3867), .A2(n3410), .ZN(n3374) );
  INV_X1 U3894 ( .A(n3398), .ZN(n4402) );
  NAND2_X1 U3895 ( .A1(n4673), .A2(STATE2_REG_3__SCAN_IN), .ZN(n4424) );
  NAND2_X1 U3896 ( .A1(n5040), .A2(n5039), .ZN(n6808) );
  NAND2_X1 U3897 ( .A1(n5384), .A2(REIP_REG_20__SCAN_IN), .ZN(n5369) );
  OR2_X1 U3898 ( .A1(n5448), .A2(n5208), .ZN(n5420) );
  AND2_X1 U3899 ( .A1(n5517), .A2(n5046), .ZN(n6451) );
  AND2_X1 U3900 ( .A1(n6423), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6452) );
  AND2_X1 U3901 ( .A1(n5517), .A2(n5190), .ZN(n6459) );
  AND2_X1 U3902 ( .A1(n5517), .A2(n5203), .ZN(n6441) );
  INV_X1 U3903 ( .A(n6441), .ZN(n6467) );
  AND2_X1 U3904 ( .A1(n5251), .A2(n5188), .ZN(n6427) );
  INV_X1 U3905 ( .A(n6452), .ZN(n6444) );
  AND2_X2 U3906 ( .A1(n4377), .A2(n4737), .ZN(n6480) );
  INV_X1 U3907 ( .A(n3400), .ZN(n5266) );
  OR2_X1 U3908 ( .A1(n5645), .A2(n5646), .ZN(n5659) );
  INV_X1 U3909 ( .A(n4826), .ZN(n6434) );
  AND2_X1 U3910 ( .A1(n4724), .A2(n4723), .ZN(n4725) );
  INV_X1 U3911 ( .A(n5659), .ZN(n5665) );
  INV_X1 U3912 ( .A(n6481), .ZN(n6490) );
  AND2_X1 U3913 ( .A1(n4363), .A2(n4472), .ZN(n6814) );
  OR2_X2 U3914 ( .A1(n5040), .A2(n4334), .ZN(n6556) );
  XNOR2_X1 U3915 ( .A(n5186), .B(n5258), .ZN(n5251) );
  OR2_X1 U3916 ( .A1(n5185), .A2(n5669), .ZN(n5186) );
  INV_X1 U3917 ( .A(n5308), .ZN(n5307) );
  OR2_X1 U3918 ( .A1(n5657), .A2(n5656), .ZN(n6472) );
  INV_X1 U3919 ( .A(n6639), .ZN(n6577) );
  XNOR2_X1 U3920 ( .A(n4995), .B(n4994), .ZN(n5243) );
  INV_X1 U3921 ( .A(n3251), .ZN(n5056) );
  XNOR2_X1 U3922 ( .A(n3205), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5254)
         );
  NAND2_X1 U3923 ( .A1(n3100), .A2(n3206), .ZN(n3205) );
  NAND2_X1 U3924 ( .A1(n5236), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3206) );
  NOR2_X1 U3925 ( .A1(n5231), .A2(n5230), .ZN(n5903) );
  OR2_X1 U3926 ( .A1(n5923), .A2(n5911), .ZN(n5231) );
  INV_X1 U3927 ( .A(n3180), .ZN(n5740) );
  NOR2_X1 U3928 ( .A1(n5962), .A2(n3886), .ZN(n5936) );
  AND2_X1 U3929 ( .A1(n3269), .A2(n3669), .ZN(n5786) );
  NAND2_X1 U3930 ( .A1(n3482), .A2(n3481), .ZN(n3198) );
  INV_X1 U3931 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3157) );
  INV_X1 U3932 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4952) );
  NAND2_X1 U3933 ( .A1(n4376), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6061) );
  OAI211_X1 U3934 ( .C1(n6112), .C2(n6116), .A(n6212), .B(n6300), .ZN(n6138)
         );
  OR2_X1 U3935 ( .A1(n4544), .A2(n4583), .ZN(n6107) );
  AND2_X1 U3936 ( .A1(n4543), .A2(n4670), .ZN(n4779) );
  AND2_X1 U3937 ( .A1(n4789), .A2(n4788), .ZN(n4813) );
  AND4_X1 U3938 ( .A1(n4607), .A2(n6212), .A3(n4606), .A4(n6315), .ZN(n4742)
         );
  OAI21_X1 U3939 ( .B1(n6215), .B2(n6668), .A(n6214), .ZN(n6238) );
  INV_X1 U3940 ( .A(n4846), .ZN(n4880) );
  INV_X1 U3941 ( .A(n6676), .ZN(n6306) );
  INV_X1 U3942 ( .A(n6683), .ZN(n6320) );
  INV_X1 U3943 ( .A(n6690), .ZN(n6325) );
  INV_X1 U3944 ( .A(n6697), .ZN(n6330) );
  INV_X1 U3945 ( .A(n6711), .ZN(n6340) );
  INV_X1 U3946 ( .A(n6718), .ZN(n6345) );
  INV_X1 U3947 ( .A(n6728), .ZN(n6351) );
  OAI21_X1 U3948 ( .B1(n5279), .B2(REIP_REG_29__SCAN_IN), .A(n3222), .ZN(U2798) );
  INV_X1 U3949 ( .A(n3223), .ZN(n3222) );
  OR2_X1 U3950 ( .A1(n5288), .A2(n6952), .ZN(n3228) );
  NAND2_X1 U3951 ( .A1(n3160), .A2(n6592), .ZN(n3159) );
  INV_X1 U3952 ( .A(n5897), .ZN(n3160) );
  NAND2_X1 U3953 ( .A1(n3889), .A2(n6592), .ZN(n4248) );
  OAI21_X1 U3954 ( .B1(n5628), .B2(n5858), .A(n4245), .ZN(n4246) );
  INV_X1 U3955 ( .A(n3168), .ZN(n3167) );
  OAI21_X1 U3956 ( .B1(n5774), .B2(n5858), .A(n5772), .ZN(n3168) );
  INV_X1 U3957 ( .A(n3247), .ZN(n5234) );
  OAI21_X1 U3958 ( .B1(n5270), .B2(n6640), .A(n3248), .ZN(n3247) );
  OR2_X1 U3959 ( .A1(n5878), .A2(n5877), .ZN(n3190) );
  NAND2_X1 U3960 ( .A1(n5955), .A2(n6653), .ZN(n5961) );
  AND2_X1 U3961 ( .A1(n6203), .A2(n3120), .ZN(n3091) );
  AND2_X1 U3962 ( .A1(n3262), .A2(n3121), .ZN(n3092) );
  AND2_X1 U3963 ( .A1(n5730), .A2(n3279), .ZN(n3093) );
  NAND2_X1 U3964 ( .A1(n4659), .A2(n4661), .ZN(n4660) );
  AND2_X1 U3965 ( .A1(n3124), .A2(n3614), .ZN(n3094) );
  NAND2_X1 U3966 ( .A1(n5813), .A2(n5930), .ZN(n3095) );
  NAND2_X1 U3967 ( .A1(n5824), .A2(n5738), .ZN(n3096) );
  AND2_X1 U3968 ( .A1(n5221), .A2(n3214), .ZN(n3097) );
  BUF_X1 U3969 ( .A(n5116), .Z(n4192) );
  INV_X1 U3970 ( .A(n3763), .ZN(n4980) );
  NOR2_X1 U3971 ( .A1(n5369), .A2(n5210), .ZN(n3217) );
  AND2_X1 U3972 ( .A1(n4991), .A2(n5050), .ZN(n3098) );
  AND2_X1 U3973 ( .A1(n5373), .A2(n3260), .ZN(n5303) );
  AND4_X1 U3974 ( .A1(n3313), .A2(n3312), .A3(n3311), .A4(n3310), .ZN(n3099)
         );
  AOI21_X1 U3975 ( .B1(n3423), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3428), 
        .ZN(n3429) );
  NOR2_X1 U3976 ( .A1(n6016), .A2(n6014), .ZN(n3814) );
  INV_X1 U3977 ( .A(n4581), .ZN(n4851) );
  NAND2_X1 U3978 ( .A1(n3186), .A2(n3542), .ZN(n4581) );
  OR3_X1 U3979 ( .A1(n5683), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3100) );
  AND2_X1 U3980 ( .A1(n3217), .A2(n3216), .ZN(n3101) );
  NAND2_X1 U3981 ( .A1(n3668), .A2(n3667), .ZN(n5793) );
  OAI21_X1 U3982 ( .B1(n7058), .B2(n3886), .A(n5815), .ZN(n3672) );
  INV_X1 U3983 ( .A(n3672), .ZN(n3200) );
  AND2_X1 U3984 ( .A1(n5813), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3102)
         );
  AND2_X1 U3985 ( .A1(n5813), .A2(n3671), .ZN(n3103) );
  AND2_X1 U3986 ( .A1(n5841), .A2(n5843), .ZN(n5809) );
  NOR2_X1 U3987 ( .A1(n4884), .A2(n4885), .ZN(n3104) );
  AND2_X1 U3988 ( .A1(n3218), .A2(n4737), .ZN(n3105) );
  OR2_X1 U3989 ( .A1(n5824), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5697)
         );
  INV_X1 U3990 ( .A(n5697), .ZN(n3214) );
  AND3_X1 U3991 ( .A1(n3414), .A2(n3413), .A3(n3854), .ZN(n3106) );
  INV_X1 U3992 ( .A(n3670), .ZN(n3203) );
  AND2_X1 U3993 ( .A1(n3097), .A2(n5235), .ZN(n3107) );
  AND2_X1 U3994 ( .A1(n3242), .A2(n5506), .ZN(n3108) );
  NAND2_X1 U3996 ( .A1(n5459), .A2(n5478), .ZN(n3109) );
  NOR2_X1 U3997 ( .A1(n5824), .A2(n5738), .ZN(n3110) );
  INV_X1 U3998 ( .A(n3185), .ZN(n3184) );
  NAND2_X1 U3999 ( .A1(n3271), .A2(n3670), .ZN(n3185) );
  AND2_X1 U4000 ( .A1(n6459), .A2(n5194), .ZN(n3111) );
  OR2_X1 U4001 ( .A1(n3418), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3112)
         );
  NAND2_X1 U4002 ( .A1(n5824), .A2(n5994), .ZN(n3113) );
  OR2_X1 U4003 ( .A1(n3543), .A2(n3529), .ZN(n3114) );
  NAND2_X1 U4004 ( .A1(n5824), .A2(n5710), .ZN(n3115) );
  INV_X1 U4005 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3144) );
  OR2_X1 U4006 ( .A1(n3191), .A2(n3190), .ZN(U2990) );
  INV_X1 U4007 ( .A(n3171), .ZN(n6660) );
  NOR2_X1 U4008 ( .A1(n4424), .A2(n3410), .ZN(n3171) );
  INV_X1 U4009 ( .A(n3152), .ZN(n6687) );
  NOR2_X1 U4010 ( .A1(n5493), .A2(n5492), .ZN(n5458) );
  NAND2_X1 U4011 ( .A1(n3188), .A2(n5389), .ZN(n3859) );
  NOR2_X1 U4012 ( .A1(n4884), .A2(n3229), .ZN(n3117) );
  NAND2_X1 U4013 ( .A1(n3641), .A2(n3640), .ZN(n3118) );
  AND2_X1 U4014 ( .A1(n3907), .A2(n4851), .ZN(n3119) );
  OR2_X1 U4015 ( .A1(n5603), .A2(n5602), .ZN(n3246) );
  INV_X1 U4016 ( .A(n5364), .ZN(n3232) );
  OR2_X1 U4017 ( .A1(n5824), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5720)
         );
  INV_X1 U4018 ( .A(n5720), .ZN(n3279) );
  AND2_X1 U4019 ( .A1(n3907), .A2(n4581), .ZN(n3120) );
  AND2_X1 U4020 ( .A1(n4973), .A2(n5026), .ZN(n3121) );
  OR2_X1 U4021 ( .A1(n5427), .A2(n5442), .ZN(n3122) );
  AND2_X1 U4022 ( .A1(n3618), .A2(n3196), .ZN(n3123) );
  AND2_X1 U4023 ( .A1(n3785), .A2(n3784), .ZN(n4537) );
  NAND2_X1 U4024 ( .A1(n4820), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3124)
         );
  AND2_X1 U4025 ( .A1(n3739), .A2(n5200), .ZN(n4281) );
  INV_X1 U4026 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n4531) );
  AND2_X1 U4027 ( .A1(n5765), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3125)
         );
  INV_X1 U4028 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3145) );
  INV_X1 U4029 ( .A(n3669), .ZN(n3270) );
  OR2_X1 U4030 ( .A1(n4715), .A2(n4516), .ZN(n6362) );
  INV_X1 U4031 ( .A(n6362), .ZN(n6592) );
  AND2_X1 U4032 ( .A1(n5206), .A2(n5207), .ZN(n3126) );
  NOR2_X1 U4033 ( .A1(n4467), .A2(n4466), .ZN(n4468) );
  AND2_X1 U4034 ( .A1(n3126), .A2(n3221), .ZN(n3127) );
  AND2_X1 U4035 ( .A1(n3127), .A2(REIP_REG_14__SCAN_IN), .ZN(n3128) );
  AND3_X1 U4036 ( .A1(REIP_REG_14__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .A3(
        REIP_REG_13__SCAN_IN), .ZN(n3129) );
  AND2_X1 U4037 ( .A1(n5682), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3130)
         );
  AND2_X4 U4038 ( .A1(n4315), .A2(n3165), .ZN(n3490) );
  NAND2_X2 U4039 ( .A1(n3131), .A2(n3459), .ZN(n3549) );
  XNOR2_X2 U4040 ( .A(n3132), .B(n3448), .ZN(n4310) );
  NAND2_X1 U4041 ( .A1(n3446), .A2(n3447), .ZN(n3132) );
  OAI211_X2 U4042 ( .C1(n3136), .C2(n3135), .A(n3666), .B(n3133), .ZN(n5800)
         );
  NAND2_X1 U4043 ( .A1(n5850), .A2(n5849), .ZN(n5808) );
  NAND2_X1 U4044 ( .A1(n3143), .A2(n3141), .ZN(n3574) );
  NAND2_X1 U4045 ( .A1(n3142), .A2(n3140), .ZN(n3139) );
  NAND2_X1 U4046 ( .A1(n3517), .A2(n3516), .ZN(n3143) );
  NAND3_X1 U4047 ( .A1(n3572), .A2(n3573), .A3(n3146), .ZN(n4659) );
  NAND4_X1 U4048 ( .A1(n3148), .A2(n3417), .A3(n3147), .A4(n3407), .ZN(n3149)
         );
  NAND2_X1 U4049 ( .A1(n4726), .A2(n3713), .ZN(n3407) );
  NAND2_X1 U4050 ( .A1(n3409), .A2(n3410), .ZN(n3147) );
  AND2_X2 U4051 ( .A1(n3149), .A2(n3158), .ZN(n3423) );
  OR2_X2 U4052 ( .A1(n5747), .A2(n5224), .ZN(n5681) );
  NAND2_X1 U4053 ( .A1(n3269), .A2(n3201), .ZN(n3150) );
  NAND2_X1 U4054 ( .A1(n3519), .A2(n3153), .ZN(n3848) );
  NAND4_X1 U4055 ( .A1(n4406), .A2(n3153), .A3(n5266), .A4(n4717), .ZN(n4375)
         );
  AND2_X1 U4056 ( .A1(n4406), .A2(n3153), .ZN(n3151) );
  MUX2_X1 U4057 ( .A(n3744), .B(n3743), .S(n3153), .Z(n3756) );
  NOR2_X1 U4058 ( .A1(n4424), .A2(n3153), .ZN(n3152) );
  AND2_X2 U4059 ( .A1(n4314), .A2(n3298), .ZN(n3460) );
  AND2_X2 U4060 ( .A1(n3155), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3298)
         );
  AND2_X2 U4061 ( .A1(n4319), .A2(n3165), .ZN(n3498) );
  NAND2_X1 U4062 ( .A1(n5706), .A2(n3159), .ZN(U2960) );
  AND2_X2 U4063 ( .A1(n5352), .A2(n5351), .ZN(n5353) );
  NOR2_X2 U4064 ( .A1(n3230), .A2(n4884), .ZN(n5352) );
  NAND2_X1 U4065 ( .A1(n3163), .A2(n4324), .ZN(n6455) );
  NAND3_X1 U4066 ( .A1(n3163), .A2(n4324), .A3(n4531), .ZN(n3189) );
  INV_X1 U4067 ( .A(n3431), .ZN(n3164) );
  NAND2_X1 U4068 ( .A1(n3165), .A2(n4525), .ZN(n4526) );
  AND2_X2 U4069 ( .A1(n3297), .A2(n3165), .ZN(n3486) );
  NOR2_X1 U4070 ( .A1(n4493), .A2(n3165), .ZN(n4502) );
  AND2_X2 U4071 ( .A1(n3422), .A2(n3447), .ZN(n3431) );
  NAND2_X1 U4072 ( .A1(n3423), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3166) );
  NAND2_X1 U4073 ( .A1(n5773), .A2(n3167), .ZN(U2969) );
  OAI21_X1 U4074 ( .B1(n5768), .B2(n3170), .A(n5767), .ZN(n5955) );
  NAND2_X2 U4075 ( .A1(n3410), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3530) );
  NAND2_X1 U4076 ( .A1(n3174), .A2(n3722), .ZN(n3725) );
  NAND2_X1 U4077 ( .A1(n3175), .A2(n3720), .ZN(n3174) );
  AOI21_X1 U4078 ( .B1(n3712), .B2(n3711), .A(n3734), .ZN(n3176) );
  OAI22_X1 U4079 ( .A1(n3712), .A2(n3709), .B1(n3708), .B2(n3707), .ZN(n3177)
         );
  NAND2_X2 U4080 ( .A1(n3345), .A2(n4373), .ZN(n3749) );
  NAND2_X1 U4081 ( .A1(n3179), .A2(n3094), .ZN(n3265) );
  NAND2_X1 U4082 ( .A1(n6571), .A2(n6570), .ZN(n3179) );
  CLKBUF_X1 U4083 ( .A(n3179), .Z(n3178) );
  OAI21_X1 U4084 ( .B1(n6571), .B2(n6570), .A(n3178), .ZN(n6572) );
  AOI21_X2 U4085 ( .B1(n3180), .B2(n3096), .A(n3110), .ZN(n5731) );
  CLKBUF_X1 U4086 ( .A(n5050), .Z(n3187) );
  NAND2_X1 U4087 ( .A1(n3187), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3793)
         );
  NAND2_X1 U4088 ( .A1(n3187), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4977) );
  INV_X2 U4089 ( .A(n5050), .ZN(n5389) );
  INV_X1 U4090 ( .A(n3759), .ZN(n3188) );
  NAND2_X1 U4091 ( .A1(n3771), .A2(n5050), .ZN(n4993) );
  NAND3_X1 U4092 ( .A1(n3776), .A2(n3775), .A3(n3187), .ZN(n3777) );
  NAND3_X1 U4093 ( .A1(n3811), .A2(n3810), .A3(n3187), .ZN(n3812) );
  NAND3_X1 U4094 ( .A1(n3790), .A2(n3789), .A3(n3187), .ZN(n3791) );
  NAND3_X1 U4095 ( .A1(n3798), .A2(n3797), .A3(n3187), .ZN(n3799) );
  NAND3_X1 U4096 ( .A1(n3804), .A2(n3803), .A3(n3187), .ZN(n3805) );
  NAND3_X1 U4097 ( .A1(n3819), .A2(n3818), .A3(n3187), .ZN(n3820) );
  OAI211_X1 U4098 ( .C1(n3764), .C2(EBX_REG_16__SCAN_IN), .A(n3824), .B(n3187), 
        .ZN(n3825) );
  MUX2_X1 U4099 ( .A(n4987), .B(n3187), .S(EBX_REG_5__SCAN_IN), .Z(n3787) );
  MUX2_X1 U4100 ( .A(n4987), .B(n3187), .S(EBX_REG_11__SCAN_IN), .Z(n3807) );
  MUX2_X1 U4101 ( .A(n4987), .B(n3187), .S(EBX_REG_15__SCAN_IN), .Z(n3816) );
  MUX2_X1 U4102 ( .A(n4987), .B(n3187), .S(EBX_REG_13__SCAN_IN), .Z(n3815) );
  MUX2_X1 U4103 ( .A(n4987), .B(n3187), .S(EBX_REG_17__SCAN_IN), .Z(n3822) );
  MUX2_X1 U4104 ( .A(n4987), .B(n3187), .S(EBX_REG_24__SCAN_IN), .Z(n4972) );
  MUX2_X1 U4105 ( .A(n3187), .B(n5391), .S(n5380), .Z(n5382) );
  NAND2_X1 U4106 ( .A1(n3189), .A2(n3114), .ZN(n3445) );
  NAND2_X2 U4107 ( .A1(n3198), .A2(n3483), .ZN(n3915) );
  AOI21_X2 U4108 ( .B1(n3202), .B2(n3670), .A(n3103), .ZN(n3201) );
  INV_X1 U4109 ( .A(n3615), .ZN(n3208) );
  INV_X1 U4110 ( .A(n3574), .ZN(n3209) );
  NAND2_X1 U4111 ( .A1(n3673), .A2(n3213), .ZN(n3215) );
  AND2_X1 U4112 ( .A1(n3215), .A2(n3097), .ZN(n5692) );
  NAND2_X1 U4113 ( .A1(n3215), .A2(n5221), .ZN(n5711) );
  INV_X2 U4114 ( .A(n3659), .ZN(n5813) );
  OAI21_X1 U4115 ( .B1(n3735), .B2(n3728), .A(n3738), .ZN(n3220) );
  AND2_X2 U4116 ( .A1(n5323), .A2(n3236), .ZN(n5273) );
  INV_X1 U4117 ( .A(n5603), .ZN(n3241) );
  NAND3_X1 U4118 ( .A1(n3251), .A2(n5047), .A3(n3250), .ZN(n3249) );
  INV_X1 U4119 ( .A(n5536), .ZN(n3255) );
  NAND2_X1 U4120 ( .A1(n3255), .A2(n3257), .ZN(n4887) );
  NAND2_X1 U4121 ( .A1(n3392), .A2(n3391), .ZN(n3850) );
  AND3_X2 U4122 ( .A1(n3392), .A2(n3391), .A3(n3264), .ZN(n3748) );
  INV_X1 U4123 ( .A(n3848), .ZN(n3264) );
  NAND2_X1 U4124 ( .A1(n3649), .A2(n3265), .ZN(n6565) );
  OAI21_X1 U4125 ( .B1(n4821), .B2(n3266), .A(n6563), .ZN(n4836) );
  NAND2_X1 U4126 ( .A1(n4821), .A2(n3266), .ZN(n6563) );
  INV_X1 U4127 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3267) );
  AND2_X2 U4128 ( .A1(n3267), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3297)
         );
  AND2_X1 U4129 ( .A1(n3145), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3699)
         );
  NAND2_X1 U4130 ( .A1(n4328), .A2(n3145), .ZN(n4329) );
  NAND2_X1 U4131 ( .A1(n5731), .A2(n3093), .ZN(n3273) );
  AOI21_X1 U4132 ( .B1(n5731), .B2(n3275), .A(n3278), .ZN(n3274) );
  NAND2_X1 U4133 ( .A1(n3673), .A2(n3280), .ZN(n3282) );
  INV_X1 U4134 ( .A(n3282), .ZN(n5746) );
  AND2_X2 U4135 ( .A1(n3144), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3299)
         );
  NAND2_X1 U4136 ( .A1(n3796), .A2(n3795), .ZN(n5603) );
  INV_X2 U4137 ( .A(n3396), .ZN(n4413) );
  XNOR2_X1 U4138 ( .A(n3574), .B(n4581), .ZN(n4542) );
  INV_X1 U4139 ( .A(n4887), .ZN(n3796) );
  OR2_X1 U4140 ( .A1(n5231), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3283)
         );
  AND2_X1 U4141 ( .A1(n3887), .A2(n3283), .ZN(n3284) );
  NAND2_X1 U4142 ( .A1(n6480), .A2(n5266), .ZN(n5605) );
  AND3_X1 U4143 ( .A1(n4054), .A2(n4053), .A3(n4052), .ZN(n3285) );
  OR2_X1 U4144 ( .A1(n4993), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3286)
         );
  OR2_X1 U4145 ( .A1(n4993), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3287)
         );
  AND2_X1 U4146 ( .A1(n4991), .A2(n4990), .ZN(n3289) );
  AND2_X1 U4147 ( .A1(n3545), .A2(n5197), .ZN(n3291) );
  OR2_X1 U4148 ( .A1(n4717), .A2(n3398), .ZN(n3292) );
  AND2_X1 U4149 ( .A1(n3394), .A2(n3842), .ZN(n3395) );
  AND2_X1 U4150 ( .A1(n6304), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3700)
         );
  AND2_X1 U4151 ( .A1(n3617), .A2(n3616), .ZN(n3618) );
  OR2_X1 U4152 ( .A1(n3442), .A2(n3441), .ZN(n3518) );
  OR3_X1 U4153 ( .A1(n3694), .A2(n6659), .A3(INSTQUEUERD_ADDR_REG_4__SCAN_IN), 
        .ZN(n3733) );
  INV_X1 U4154 ( .A(n3701), .ZN(n3406) );
  OR2_X1 U4155 ( .A1(n3628), .A2(n3627), .ZN(n3643) );
  OR2_X1 U4156 ( .A1(n3458), .A2(n3457), .ZN(n3553) );
  INV_X1 U4157 ( .A(n3508), .ZN(n3509) );
  NAND2_X1 U4158 ( .A1(n3713), .A2(n3710), .ZN(n3734) );
  INV_X1 U4159 ( .A(n5171), .ZN(n5059) );
  AND2_X1 U4160 ( .A1(n4230), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4231)
         );
  INV_X1 U4161 ( .A(n4122), .ZN(n3975) );
  NOR2_X1 U4162 ( .A1(n4057), .A2(n3973), .ZN(n4036) );
  AND2_X1 U4163 ( .A1(n3813), .A2(n3812), .ZN(n6014) );
  INV_X1 U4164 ( .A(n4886), .ZN(n3795) );
  AND2_X1 U4165 ( .A1(n3778), .A2(n3777), .ZN(n4466) );
  AND2_X1 U4166 ( .A1(n3687), .A2(n3686), .ZN(n3736) );
  INV_X1 U4167 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4489) );
  NAND2_X1 U4168 ( .A1(n4328), .A2(STATE2_REG_0__SCAN_IN), .ZN(n5177) );
  INV_X1 U4169 ( .A(n4189), .ZN(n4188) );
  AND2_X1 U4170 ( .A1(n5396), .A2(n5395), .ZN(n5378) );
  AND2_X1 U4171 ( .A1(n5657), .A2(n5454), .ZN(n5473) );
  INV_X1 U4172 ( .A(n3971), .ZN(n3972) );
  AND2_X1 U4173 ( .A1(n3781), .A2(n3780), .ZN(n5534) );
  INV_X1 U4174 ( .A(n3755), .ZN(n4328) );
  OAI21_X1 U4175 ( .B1(n6078), .B2(n6077), .A(n6076), .ZN(n6100) );
  NAND2_X1 U4176 ( .A1(n3528), .A2(n3527), .ZN(n4780) );
  XNOR2_X1 U4177 ( .A(n3551), .B(n3550), .ZN(n4387) );
  AND2_X1 U4178 ( .A1(n3524), .A2(n4425), .ZN(n6249) );
  INV_X1 U4179 ( .A(n6206), .ZN(n6312) );
  NAND2_X1 U4180 ( .A1(n5060), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5185)
         );
  NOR2_X1 U4181 ( .A1(n4107), .A2(n6401), .ZN(n4100) );
  OR2_X1 U4182 ( .A1(n3992), .A2(n5769), .ZN(n4137) );
  NAND2_X1 U4183 ( .A1(n4074), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4057)
         );
  AND2_X1 U4184 ( .A1(n3826), .A2(n3825), .ZN(n5442) );
  NAND2_X1 U4185 ( .A1(n6072), .A2(n3912), .ZN(n6103) );
  AND2_X1 U4186 ( .A1(n4670), .A2(n4669), .ZN(n6072) );
  INV_X1 U4187 ( .A(n4815), .ZN(n4653) );
  AND2_X1 U4188 ( .A1(n4904), .A2(n4903), .ZN(n4934) );
  INV_X1 U4189 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6302) );
  NAND2_X1 U4190 ( .A1(n4853), .A2(n4852), .ZN(n6295) );
  OR2_X1 U4191 ( .A1(n4424), .A2(n5266), .ZN(n6723) );
  AND2_X1 U4192 ( .A1(n4513), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3757) );
  OR2_X1 U4193 ( .A1(n4286), .A2(n6736), .ZN(n5039) );
  NAND2_X1 U4194 ( .A1(n5054), .A2(n5053), .ZN(n5055) );
  INV_X1 U4195 ( .A(n5605), .ZN(n6477) );
  INV_X1 U4196 ( .A(n5664), .ZN(n5658) );
  OR2_X2 U4197 ( .A1(n5040), .A2(n4335), .ZN(n6557) );
  AND2_X1 U4198 ( .A1(n5398), .A2(n5397), .ZN(n5754) );
  AND2_X1 U4199 ( .A1(n5441), .A2(n5440), .ZN(n5783) );
  AND2_X1 U4200 ( .A1(n5586), .A2(n5585), .ZN(n6392) );
  NAND2_X1 U4201 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n3933), .ZN(n3948)
         );
  OR2_X1 U4202 ( .A1(n5929), .A2(n5983), .ZN(n6032) );
  INV_X1 U4203 ( .A(n6103), .ZN(n4710) );
  INV_X1 U4204 ( .A(n6107), .ZN(n6142) );
  AND2_X1 U4205 ( .A1(n4853), .A2(n4624), .ZN(n4815) );
  AND2_X1 U4206 ( .A1(n4853), .A2(n4602), .ZN(n6150) );
  INV_X1 U4207 ( .A(n4742), .ZN(n6146) );
  AND3_X1 U4208 ( .A1(n3119), .A2(n3912), .A3(n6203), .ZN(n6151) );
  OAI21_X1 U4209 ( .B1(n4432), .B2(n4605), .A(n4618), .ZN(n4455) );
  AND2_X1 U4210 ( .A1(n3119), .A2(n6246), .ZN(n4937) );
  INV_X1 U4211 ( .A(n6732), .ZN(n6242) );
  NAND2_X1 U4212 ( .A1(n4583), .A2(n6056), .ZN(n6665) );
  OAI21_X1 U4213 ( .B1(n4849), .B2(n4848), .A(n4847), .ZN(n4875) );
  AND2_X1 U4214 ( .A1(n4853), .A2(n4850), .ZN(n6309) );
  AND2_X1 U4215 ( .A1(n4257), .A2(n6663), .ZN(n5839) );
  INV_X1 U4216 ( .A(n4707), .ZN(n4428) );
  INV_X1 U4217 ( .A(n5858), .ZN(n6594) );
  INV_X1 U4218 ( .A(n6478), .ZN(n6471) );
  INV_X1 U4219 ( .A(n5754), .ZN(n5639) );
  INV_X1 U4220 ( .A(n5783), .ZN(n5649) );
  INV_X1 U4221 ( .A(n6392), .ZN(n5663) );
  NAND2_X1 U4222 ( .A1(n6556), .A2(n4725), .ZN(n5664) );
  INV_X1 U4223 ( .A(n6812), .ZN(n6506) );
  OR2_X1 U4224 ( .A1(n4715), .A2(n4530), .ZN(n6561) );
  INV_X1 U4225 ( .A(n6557), .ZN(n6523) );
  INV_X1 U4226 ( .A(n4246), .ZN(n4247) );
  INV_X1 U4227 ( .A(n5839), .ZN(n5858) );
  NAND2_X1 U4228 ( .A1(n5853), .A2(n4345), .ZN(n6599) );
  NAND2_X1 U4229 ( .A1(n6032), .A2(n3885), .ZN(n5962) );
  INV_X1 U4230 ( .A(n6653), .ZN(n6638) );
  INV_X1 U4231 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4474) );
  NOR2_X1 U4232 ( .A1(n4675), .A2(n4674), .ZN(n4713) );
  AOI22_X1 U4233 ( .A1(n6070), .A2(n6077), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6074), .ZN(n6106) );
  INV_X1 U4234 ( .A(n6109), .ZN(n6145) );
  INV_X1 U4235 ( .A(n4779), .ZN(n4818) );
  AOI21_X1 U4236 ( .B1(n4620), .B2(n4622), .A(n4619), .ZN(n4658) );
  INV_X1 U4237 ( .A(n4937), .ZN(n4461) );
  OR2_X1 U4238 ( .A1(n6665), .A2(n4891), .ZN(n6199) );
  AOI22_X1 U4239 ( .A1(n6162), .A2(n6167), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6161), .ZN(n6202) );
  AOI21_X1 U4240 ( .B1(n6209), .B2(n6668), .A(n6208), .ZN(n6245) );
  OR2_X1 U4241 ( .A1(n6665), .A2(n6204), .ZN(n6732) );
  OR2_X1 U4242 ( .A1(n6665), .A2(n6247), .ZN(n6725) );
  INV_X1 U4243 ( .A(n6704), .ZN(n6335) );
  INV_X1 U4244 ( .A(n6309), .ZN(n6359) );
  INV_X1 U4245 ( .A(n6354), .ZN(n4431) );
  AOI22_X1 U4246 ( .A1(n4075), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3487), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3296) );
  AOI22_X1 U4247 ( .A1(n5116), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3486), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3295) );
  AND2_X4 U4248 ( .A1(n3299), .A2(n4314), .ZN(n3488) );
  AOI22_X1 U4249 ( .A1(n3488), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3535), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3294) );
  AOI22_X1 U4250 ( .A1(n3489), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3087), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3293) );
  NAND4_X1 U4251 ( .A1(n3296), .A2(n3295), .A3(n3294), .A4(n3293), .ZN(n3305)
         );
  AOI22_X1 U4252 ( .A1(n3498), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3485), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3303) );
  AOI22_X1 U4253 ( .A1(n3460), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3467), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3302) );
  AND2_X2 U4254 ( .A1(n4319), .A2(n3298), .ZN(n3495) );
  AOI22_X1 U4255 ( .A1(n3495), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3497), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3301) );
  AOI22_X1 U4256 ( .A1(n3484), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3490), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3300) );
  NAND4_X1 U4257 ( .A1(n3303), .A2(n3302), .A3(n3301), .A4(n3300), .ZN(n3304)
         );
  AOI22_X1 U4258 ( .A1(n5116), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4075), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3309) );
  AOI22_X1 U4259 ( .A1(n3467), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3489), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3308) );
  AOI22_X1 U4260 ( .A1(n3484), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3087), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3307) );
  AOI22_X1 U4261 ( .A1(n3498), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3306) );
  AOI22_X1 U4262 ( .A1(n3495), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3486), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3313) );
  AOI22_X1 U4263 ( .A1(n3485), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3535), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3312) );
  AOI22_X1 U4264 ( .A1(n3488), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3497), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3311) );
  AOI22_X1 U4265 ( .A1(n3487), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3490), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3310) );
  INV_X2 U4266 ( .A(n3384), .ZN(n3387) );
  NAND2_X2 U4267 ( .A1(n3398), .A2(n3387), .ZN(n4373) );
  NAND2_X1 U4268 ( .A1(n5116), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3318)
         );
  NAND2_X1 U4269 ( .A1(n3495), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3317) );
  NAND2_X1 U4270 ( .A1(n3498), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3316)
         );
  NAND2_X1 U4271 ( .A1(n3088), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3315) );
  NAND2_X1 U4272 ( .A1(n3484), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3322) );
  NAND2_X1 U4273 ( .A1(n3460), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3321) );
  NAND2_X1 U4274 ( .A1(n4075), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3320)
         );
  NAND2_X1 U4275 ( .A1(n3497), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3319) );
  NAND2_X1 U4276 ( .A1(n3486), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3326)
         );
  NAND2_X1 U4277 ( .A1(n3485), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3325) );
  NAND2_X1 U4278 ( .A1(n3487), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3324) );
  NAND2_X1 U4279 ( .A1(n3490), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3323)
         );
  NAND2_X1 U4280 ( .A1(n3467), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3330) );
  NAND2_X1 U4281 ( .A1(n3488), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3329) );
  NAND2_X1 U4282 ( .A1(n3489), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3328) );
  NAND2_X1 U4283 ( .A1(n3535), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3327)
         );
  NAND4_X4 U4284 ( .A1(n3334), .A2(n3333), .A3(n3332), .A4(n3331), .ZN(n3405)
         );
  AOI22_X1 U4285 ( .A1(n3498), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3338) );
  AOI22_X1 U4286 ( .A1(n5116), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4075), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3337) );
  AOI22_X1 U4287 ( .A1(n3467), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3489), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3336) );
  AOI22_X1 U4288 ( .A1(n3484), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3089), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3335) );
  NAND4_X1 U4289 ( .A1(n3338), .A2(n3337), .A3(n3336), .A4(n3335), .ZN(n3344)
         );
  AOI22_X1 U4290 ( .A1(n3495), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3486), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3342) );
  AOI22_X1 U4291 ( .A1(n3485), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3535), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3341) );
  AOI22_X1 U4292 ( .A1(n3488), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3497), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3340) );
  AOI22_X1 U4293 ( .A1(n3487), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3490), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3339) );
  NAND4_X1 U4294 ( .A1(n3342), .A2(n3341), .A3(n3340), .A4(n3339), .ZN(n3343)
         );
  INV_X1 U4295 ( .A(n3401), .ZN(n3345) );
  AOI22_X1 U4296 ( .A1(n5116), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4075), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3348) );
  AOI22_X1 U4297 ( .A1(n3467), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3489), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3347) );
  AOI22_X1 U4298 ( .A1(n3484), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3087), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3346) );
  AOI22_X1 U4299 ( .A1(n3495), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3486), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3353) );
  AOI22_X1 U4300 ( .A1(n3485), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3535), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3352) );
  AOI22_X1 U4301 ( .A1(n3488), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3497), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3351) );
  AOI22_X1 U4302 ( .A1(n3487), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3490), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3350) );
  AOI22_X1 U4303 ( .A1(n5116), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3087), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3357) );
  AOI22_X1 U4304 ( .A1(n3460), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3486), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3356) );
  AOI22_X1 U4305 ( .A1(n3495), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4075), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3355) );
  AOI22_X1 U4306 ( .A1(n3485), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3535), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3354) );
  NAND4_X1 U4307 ( .A1(n3357), .A2(n3356), .A3(n3355), .A4(n3354), .ZN(n3363)
         );
  AOI22_X1 U4308 ( .A1(n3498), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3487), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3361) );
  AOI22_X1 U4309 ( .A1(n3484), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3467), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3360) );
  AOI22_X1 U4310 ( .A1(n3488), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3497), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3359) );
  AOI22_X1 U4311 ( .A1(n3489), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3490), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3358) );
  NAND4_X1 U4312 ( .A1(n3361), .A2(n3360), .A3(n3359), .A4(n3358), .ZN(n3362)
         );
  OR2_X2 U4313 ( .A1(n3404), .A2(n4406), .ZN(n3411) );
  NAND2_X1 U4314 ( .A1(n4402), .A2(n3400), .ZN(n3867) );
  AOI22_X1 U4315 ( .A1(n3495), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4075), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3367) );
  AOI22_X1 U4316 ( .A1(n3484), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3467), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3366) );
  AOI22_X1 U4317 ( .A1(n5116), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3497), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3365) );
  AOI22_X1 U4318 ( .A1(n3488), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3535), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3364) );
  NAND4_X1 U4319 ( .A1(n3367), .A2(n3366), .A3(n3365), .A4(n3364), .ZN(n3373)
         );
  AOI22_X1 U4320 ( .A1(n3498), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3371) );
  AOI22_X1 U4321 ( .A1(n3485), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3489), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3370) );
  AOI22_X1 U4322 ( .A1(n3460), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3486), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3369) );
  AOI22_X1 U4323 ( .A1(n3487), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3490), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3368) );
  NAND4_X1 U4324 ( .A1(n3371), .A2(n3370), .A3(n3369), .A4(n3368), .ZN(n3372)
         );
  OR2_X4 U4325 ( .A1(n3373), .A2(n3372), .ZN(n5200) );
  AOI22_X1 U4326 ( .A1(n3498), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3378) );
  AOI22_X1 U4327 ( .A1(n3484), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3089), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3377) );
  AOI22_X1 U4328 ( .A1(n3467), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3489), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3376) );
  AOI22_X1 U4329 ( .A1(n5116), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4075), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3375) );
  AOI22_X1 U4330 ( .A1(n3495), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3486), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3382) );
  AOI22_X1 U4331 ( .A1(n3485), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3535), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3381) );
  AOI22_X1 U4332 ( .A1(n3488), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3497), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3380) );
  AOI22_X1 U4333 ( .A1(n3487), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3490), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3379) );
  NAND2_X2 U4334 ( .A1(n3752), .A2(n4413), .ZN(n4721) );
  CLKBUF_X3 U4335 ( .A(n3384), .Z(n3745) );
  NOR2_X1 U4336 ( .A1(n3848), .A2(n3745), .ZN(n3385) );
  XNOR2_X1 U4337 ( .A(STATE_REG_1__SCAN_IN), .B(STATE_REG_2__SCAN_IN), .ZN(
        n3676) );
  NAND2_X1 U4338 ( .A1(n4413), .A2(n3676), .ZN(n3393) );
  AND2_X2 U4339 ( .A1(n3410), .A2(n4413), .ZN(n4279) );
  NAND2_X1 U4340 ( .A1(n3398), .A2(n3400), .ZN(n3894) );
  NAND2_X1 U4341 ( .A1(n4721), .A2(n3388), .ZN(n3389) );
  NAND2_X1 U4342 ( .A1(n3389), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3421) );
  INV_X1 U4343 ( .A(n3421), .ZN(n3390) );
  NOR2_X1 U4344 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n4948) );
  NAND2_X1 U4345 ( .A1(n4948), .A2(n4531), .ZN(n6805) );
  XNOR2_X1 U4346 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6301) );
  INV_X1 U4347 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n4513) );
  OAI22_X1 U4348 ( .A1(n6805), .A2(n6301), .B1(n3757), .B2(n4839), .ZN(n3418)
         );
  NAND2_X1 U4349 ( .A1(n3390), .A2(n3112), .ZN(n3446) );
  NAND2_X1 U4350 ( .A1(n3404), .A2(n4717), .ZN(n3392) );
  NAND2_X1 U4351 ( .A1(n3393), .A2(n3387), .ZN(n3394) );
  NAND2_X1 U4352 ( .A1(n3410), .A2(n3396), .ZN(n3842) );
  NAND2_X1 U4353 ( .A1(n3749), .A2(n5197), .ZN(n3397) );
  OAI21_X1 U4354 ( .B1(n3387), .B2(n3851), .A(n3398), .ZN(n3399) );
  NAND2_X1 U4355 ( .A1(n3399), .A2(n3292), .ZN(n3403) );
  OAI22_X1 U4356 ( .A1(n3401), .A2(n3387), .B1(n5266), .B2(n3851), .ZN(n3402)
         );
  NAND3_X1 U4357 ( .A1(n3403), .A2(n3411), .A3(n3402), .ZN(n3409) );
  MUX2_X1 U4358 ( .A(n3757), .B(n6805), .S(n6304), .Z(n3408) );
  NAND2_X1 U4359 ( .A1(n3409), .A2(n4279), .ZN(n3857) );
  INV_X1 U4360 ( .A(n3867), .ZN(n3913) );
  NAND2_X1 U4361 ( .A1(n4948), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6737) );
  AOI21_X1 U4362 ( .B1(n3860), .B2(n3913), .A(n6737), .ZN(n3414) );
  NAND2_X1 U4363 ( .A1(n3411), .A2(n5197), .ZN(n3413) );
  INV_X1 U4364 ( .A(n3842), .ZN(n5516) );
  AND2_X1 U4365 ( .A1(n5200), .A2(n3851), .ZN(n3412) );
  AOI21_X1 U4366 ( .B1(n5516), .B2(n3759), .A(n3412), .ZN(n3854) );
  OAI21_X1 U4367 ( .B1(n3404), .B2(n4717), .A(n3519), .ZN(n3415) );
  OAI21_X1 U4368 ( .B1(n3850), .B2(n3415), .A(n3396), .ZN(n3416) );
  NAND4_X1 U4369 ( .A1(n3857), .A2(n3417), .A3(n3106), .A4(n3416), .ZN(n3480)
         );
  NAND2_X1 U4370 ( .A1(n3446), .A2(n3483), .ZN(n3422) );
  INV_X1 U4371 ( .A(n3418), .ZN(n3420) );
  NAND2_X1 U4372 ( .A1(n3423), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3419) );
  NAND3_X1 U4373 ( .A1(n3421), .A2(n3420), .A3(n3419), .ZN(n3447) );
  AND2_X1 U4374 ( .A1(n4489), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6210)
         );
  NAND2_X1 U4375 ( .A1(n6210), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3426) );
  NAND2_X1 U4376 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3424) );
  NAND2_X1 U4377 ( .A1(n3424), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3425) );
  NAND2_X1 U4378 ( .A1(n3426), .A2(n3425), .ZN(n4608) );
  INV_X1 U4379 ( .A(n6805), .ZN(n3526) );
  NAND2_X1 U4380 ( .A1(n4608), .A2(n3526), .ZN(n3427) );
  OAI21_X1 U4381 ( .B1(n3757), .B2(n4489), .A(n3427), .ZN(n3428) );
  INV_X1 U4382 ( .A(n3429), .ZN(n3430) );
  AOI22_X1 U4383 ( .A1(n5121), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n5107), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3435) );
  AOI22_X1 U4384 ( .A1(n5116), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5124), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3434) );
  AOI22_X1 U4385 ( .A1(n3468), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3433) );
  AOI22_X1 U4386 ( .A1(n5122), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3087), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3432) );
  NAND4_X1 U4387 ( .A1(n3435), .A2(n3434), .A3(n3433), .A4(n3432), .ZN(n3442)
         );
  BUF_X1 U4388 ( .A(n3486), .Z(n3436) );
  AOI22_X1 U4389 ( .A1(n3496), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3440) );
  AOI22_X1 U4390 ( .A1(n5123), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n5114), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3439) );
  AOI22_X1 U4391 ( .A1(n3462), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n5115), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3438) );
  AOI22_X1 U4392 ( .A1(n3086), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3437) );
  NAND4_X1 U4393 ( .A1(n3440), .A2(n3439), .A3(n3438), .A4(n3437), .ZN(n3441)
         );
  INV_X1 U4394 ( .A(n3530), .ZN(n3443) );
  AOI22_X1 U4395 ( .A1(n3713), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3443), 
        .B2(n3518), .ZN(n3444) );
  INV_X1 U4396 ( .A(n3483), .ZN(n3448) );
  INV_X1 U4397 ( .A(n3529), .ZN(n3514) );
  AOI22_X1 U4398 ( .A1(n5107), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n5124), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3452) );
  BUF_X2 U4399 ( .A(n3485), .Z(n5123) );
  AOI22_X1 U4400 ( .A1(n5123), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4401 ( .A1(n5116), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n5114), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U4402 ( .A1(n5122), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3089), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3449) );
  NAND4_X1 U4403 ( .A1(n3452), .A2(n3451), .A3(n3450), .A4(n3449), .ZN(n3458)
         );
  BUF_X2 U4404 ( .A(n3498), .Z(n5121) );
  AOI22_X1 U4405 ( .A1(n3496), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5121), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3456) );
  AOI22_X1 U4406 ( .A1(n3086), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3455) );
  AOI22_X1 U4407 ( .A1(n3462), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n5115), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3454) );
  AOI22_X1 U4408 ( .A1(n3468), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3453) );
  NAND4_X1 U4409 ( .A1(n3456), .A2(n3455), .A3(n3454), .A4(n3453), .ZN(n3457)
         );
  NAND2_X1 U4410 ( .A1(n3514), .A2(n3553), .ZN(n3459) );
  INV_X1 U4411 ( .A(n3553), .ZN(n3478) );
  NAND2_X1 U4412 ( .A1(n3713), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3477) );
  AOI22_X1 U4413 ( .A1(n5122), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5107), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3466) );
  AOI22_X1 U4414 ( .A1(n3436), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3465) );
  AOI22_X1 U4415 ( .A1(n5124), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3464) );
  BUF_X1 U4416 ( .A(n3488), .Z(n3462) );
  AOI22_X1 U4417 ( .A1(n3462), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n5115), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3463) );
  NAND4_X1 U4418 ( .A1(n3466), .A2(n3465), .A3(n3464), .A4(n3463), .ZN(n3475)
         );
  AOI22_X1 U4420 ( .A1(n5123), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3468), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3473) );
  AOI22_X1 U4421 ( .A1(n5116), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5114), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3472) );
  AOI22_X1 U4422 ( .A1(n5121), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3087), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3471) );
  BUF_X1 U4423 ( .A(n3490), .Z(n3469) );
  AOI22_X1 U4424 ( .A1(n3496), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3470) );
  NAND4_X1 U4425 ( .A1(n3473), .A2(n3472), .A3(n3471), .A4(n3470), .ZN(n3474)
         );
  NOR2_X1 U4426 ( .A1(n3529), .A2(n3654), .ZN(n3506) );
  INV_X1 U4427 ( .A(n3506), .ZN(n3476) );
  OAI211_X1 U4428 ( .C1(n3478), .C2(n3530), .A(n3477), .B(n3476), .ZN(n3548)
         );
  INV_X1 U4429 ( .A(n3479), .ZN(n3482) );
  INV_X1 U4430 ( .A(n3480), .ZN(n3481) );
  AOI22_X1 U4431 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n5122), .B1(n5123), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3494) );
  AOI22_X1 U4432 ( .A1(n5107), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3493) );
  AOI22_X1 U4433 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n3086), .B1(n3462), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3492) );
  AOI22_X1 U4434 ( .A1(n3461), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3491) );
  NAND4_X1 U4435 ( .A1(n3494), .A2(n3493), .A3(n3492), .A4(n3491), .ZN(n3504)
         );
  AOI22_X1 U4436 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n3496), .B1(n4075), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3502) );
  AOI22_X1 U4437 ( .A1(n4192), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3468), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3501) );
  AOI22_X1 U4438 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n5114), .B1(n5115), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3500) );
  AOI22_X1 U4439 ( .A1(n5121), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3499) );
  NAND4_X1 U4440 ( .A1(n3502), .A2(n3501), .A3(n3500), .A4(n3499), .ZN(n3503)
         );
  INV_X1 U4441 ( .A(n3562), .ZN(n3505) );
  NAND2_X1 U4442 ( .A1(n3505), .A2(n4717), .ZN(n3507) );
  NAND2_X1 U4443 ( .A1(n3506), .A2(n3562), .ZN(n3557) );
  NAND2_X1 U4444 ( .A1(n3713), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3513) );
  OAI21_X1 U4445 ( .B1(n3562), .B2(n4531), .A(n3701), .ZN(n3511) );
  NAND2_X1 U4446 ( .A1(n4717), .A2(n3654), .ZN(n3510) );
  AND2_X1 U4447 ( .A1(n3511), .A2(n3510), .ZN(n3512) );
  NAND2_X1 U4448 ( .A1(n3513), .A2(n3512), .ZN(n3556) );
  NAND2_X1 U4449 ( .A1(n3514), .A2(n3654), .ZN(n3515) );
  NAND2_X1 U4450 ( .A1(n3560), .A2(n3515), .ZN(n3551) );
  OAI21_X1 U4451 ( .B1(n3549), .B2(n3548), .A(n3551), .ZN(n3517) );
  NAND2_X1 U4452 ( .A1(n3549), .A2(n3548), .ZN(n3516) );
  NAND2_X1 U4453 ( .A1(n3562), .A2(n3553), .ZN(n3552) );
  XNOR2_X1 U4454 ( .A(n3552), .B(n3518), .ZN(n3520) );
  INV_X1 U4455 ( .A(n5197), .ZN(n3750) );
  OAI21_X1 U4456 ( .B1(n3520), .B2(n3750), .A(n3561), .ZN(n3521) );
  INV_X1 U4457 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3522) );
  OAI21_X1 U4458 ( .B1(n6578), .B2(n6579), .A(n3522), .ZN(n3523) );
  NAND2_X1 U4459 ( .A1(n3423), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3528) );
  AND3_X1 U4460 ( .A1(n6302), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4605) );
  NAND2_X1 U4461 ( .A1(n4605), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4456) );
  NAND2_X1 U4462 ( .A1(n4456), .A2(n6302), .ZN(n3524) );
  AND2_X1 U4463 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4840) );
  AND2_X1 U4464 ( .A1(n4840), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6305)
         );
  NAND2_X1 U4465 ( .A1(n6305), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4425) );
  NOR2_X1 U4466 ( .A1(n3757), .A2(n6302), .ZN(n3525) );
  AOI21_X1 U4467 ( .B1(n6249), .B2(n3526), .A(n3525), .ZN(n3527) );
  AOI22_X1 U4468 ( .A1(n5121), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n5107), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3534) );
  INV_X1 U4469 ( .A(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n7027) );
  AOI22_X1 U4470 ( .A1(n4192), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4075), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3533) );
  AOI22_X1 U4471 ( .A1(n3468), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3532) );
  AOI22_X1 U4472 ( .A1(n5122), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3087), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3531) );
  NAND4_X1 U4473 ( .A1(n3534), .A2(n3533), .A3(n3532), .A4(n3531), .ZN(n3541)
         );
  AOI22_X1 U4474 ( .A1(n3496), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3539) );
  AOI22_X1 U4475 ( .A1(n5123), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n5114), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3538) );
  AOI22_X1 U4476 ( .A1(n3462), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n5115), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3537) );
  AOI22_X1 U4477 ( .A1(n3086), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3536) );
  NAND4_X1 U4478 ( .A1(n3539), .A2(n3538), .A3(n3537), .A4(n3536), .ZN(n3540)
         );
  AOI22_X1 U4479 ( .A1(n3730), .A2(n3587), .B1(n3713), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3542) );
  NAND2_X1 U4480 ( .A1(n3552), .A2(n3543), .ZN(n3588) );
  INV_X1 U4481 ( .A(n3587), .ZN(n3544) );
  XNOR2_X1 U4482 ( .A(n3588), .B(n3544), .ZN(n3545) );
  AOI21_X2 U4483 ( .B1(n4542), .B2(n3710), .A(n3291), .ZN(n3547) );
  INV_X1 U4484 ( .A(n6578), .ZN(n3546) );
  NAND3_X1 U4485 ( .A1(n3546), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3573) );
  INV_X1 U4486 ( .A(n3547), .ZN(n6582) );
  XNOR2_X1 U4487 ( .A(n3549), .B(n3548), .ZN(n3550) );
  NAND2_X1 U4488 ( .A1(n4387), .A2(n3710), .ZN(n4955) );
  OAI21_X1 U4489 ( .B1(n3553), .B2(n3562), .A(n3552), .ZN(n3554) );
  OAI211_X1 U4490 ( .C1(n3554), .C2(n3750), .A(n3264), .B(n3745), .ZN(n3555)
         );
  INV_X1 U4491 ( .A(n3555), .ZN(n4954) );
  INV_X1 U4492 ( .A(n3556), .ZN(n3558) );
  NAND2_X1 U4493 ( .A1(n3558), .A2(n3557), .ZN(n3559) );
  NAND2_X2 U4494 ( .A1(n3560), .A2(n3559), .ZN(n3912) );
  NAND2_X1 U4495 ( .A1(n6071), .A2(n3710), .ZN(n3567) );
  OAI21_X1 U4496 ( .B1(n3750), .B2(n3562), .A(n3561), .ZN(n3563) );
  INV_X1 U4497 ( .A(n3563), .ZN(n3565) );
  NAND2_X1 U4498 ( .A1(n3567), .A2(n3565), .ZN(n4340) );
  AND2_X1 U4499 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4595) );
  NAND2_X1 U4500 ( .A1(n4340), .A2(n4595), .ZN(n4957) );
  AND2_X1 U4501 ( .A1(n4954), .A2(n4957), .ZN(n3564) );
  NAND2_X1 U4502 ( .A1(n4955), .A2(n3564), .ZN(n3570) );
  INV_X1 U4503 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4592) );
  AND2_X1 U4504 ( .A1(n3565), .A2(n4592), .ZN(n3566) );
  NAND2_X1 U4505 ( .A1(n3567), .A2(n3566), .ZN(n3569) );
  OR2_X1 U4506 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3568) );
  AND2_X1 U4507 ( .A1(n3569), .A2(n3568), .ZN(n4956) );
  AND2_X1 U4508 ( .A1(n3570), .A2(n4956), .ZN(n4588) );
  INV_X1 U4509 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6579) );
  NAND2_X1 U4510 ( .A1(n6578), .A2(n6579), .ZN(n3571) );
  AOI22_X1 U4511 ( .A1(n5122), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n5121), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3578) );
  AOI22_X1 U4512 ( .A1(n3496), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n5123), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3577) );
  AOI22_X1 U4513 ( .A1(n3468), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3576) );
  AOI22_X1 U4514 ( .A1(n3488), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3575) );
  NAND4_X1 U4515 ( .A1(n3578), .A2(n3577), .A3(n3576), .A4(n3575), .ZN(n3584)
         );
  AOI22_X1 U4516 ( .A1(n5107), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3582) );
  AOI22_X1 U4517 ( .A1(n5124), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3581) );
  AOI22_X1 U4518 ( .A1(n5115), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n5114), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4519 ( .A1(n4192), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3087), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3579) );
  NAND4_X1 U4520 ( .A1(n3582), .A2(n3581), .A3(n3580), .A4(n3579), .ZN(n3583)
         );
  NAND2_X1 U4521 ( .A1(n3730), .A2(n3634), .ZN(n3586) );
  NAND2_X1 U4522 ( .A1(n3713), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3585) );
  NAND2_X1 U4523 ( .A1(n3586), .A2(n3585), .ZN(n3617) );
  NAND2_X1 U4524 ( .A1(n3890), .A2(n3710), .ZN(n3591) );
  NAND2_X1 U4525 ( .A1(n3588), .A2(n3587), .ZN(n3636) );
  XNOR2_X1 U4526 ( .A(n3636), .B(n3634), .ZN(n3589) );
  NAND2_X1 U4527 ( .A1(n3589), .A2(n5197), .ZN(n3590) );
  INV_X1 U4528 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6648) );
  NAND2_X1 U4529 ( .A1(n3592), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3593)
         );
  NAND2_X1 U4530 ( .A1(n4660), .A2(n3593), .ZN(n6571) );
  NAND2_X1 U4532 ( .A1(n3208), .A2(n3617), .ZN(n3607) );
  AOI22_X1 U4533 ( .A1(n5121), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n5107), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3598) );
  AOI22_X1 U4534 ( .A1(n4192), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4075), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3597) );
  AOI22_X1 U4535 ( .A1(n3468), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3596) );
  AOI22_X1 U4536 ( .A1(n5122), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3087), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3595) );
  NAND4_X1 U4537 ( .A1(n3598), .A2(n3597), .A3(n3596), .A4(n3595), .ZN(n3604)
         );
  AOI22_X1 U4538 ( .A1(n3496), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3602) );
  AOI22_X1 U4539 ( .A1(n5123), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n5114), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3601) );
  INV_X1 U4540 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n7095) );
  AOI22_X1 U4541 ( .A1(n3488), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n5115), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3600) );
  AOI22_X1 U4542 ( .A1(n3086), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3599) );
  NAND4_X1 U4543 ( .A1(n3602), .A2(n3601), .A3(n3600), .A4(n3599), .ZN(n3603)
         );
  NAND2_X1 U4544 ( .A1(n3730), .A2(n3633), .ZN(n3606) );
  NAND2_X1 U4545 ( .A1(n3713), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3605) );
  NAND2_X1 U4546 ( .A1(n3606), .A2(n3605), .ZN(n3616) );
  XNOR2_X1 U4547 ( .A(n3607), .B(n3616), .ZN(n3932) );
  NAND2_X1 U4548 ( .A1(n3932), .A2(n3710), .ZN(n3612) );
  INV_X1 U4549 ( .A(n3636), .ZN(n3608) );
  NAND2_X1 U4550 ( .A1(n3608), .A2(n3634), .ZN(n3609) );
  XNOR2_X1 U4551 ( .A(n3609), .B(n3633), .ZN(n3610) );
  NAND2_X1 U4552 ( .A1(n3610), .A2(n5197), .ZN(n3611) );
  NAND2_X1 U4553 ( .A1(n3612), .A2(n3611), .ZN(n3613) );
  INV_X1 U4554 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3871) );
  XNOR2_X1 U4555 ( .A(n3613), .B(n3871), .ZN(n6570) );
  NAND2_X1 U4556 ( .A1(n3613), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3614)
         );
  AOI22_X1 U4557 ( .A1(n5121), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n5107), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3622) );
  AOI22_X1 U4558 ( .A1(n4192), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4075), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3621) );
  AOI22_X1 U4559 ( .A1(n3468), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3620) );
  AOI22_X1 U4560 ( .A1(n5122), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3619) );
  NAND4_X1 U4561 ( .A1(n3622), .A2(n3621), .A3(n3620), .A4(n3619), .ZN(n3628)
         );
  AOI22_X1 U4562 ( .A1(n3496), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3626) );
  AOI22_X1 U4563 ( .A1(n5123), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n5114), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3625) );
  AOI22_X1 U4564 ( .A1(n3488), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n5115), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3624) );
  AOI22_X1 U4565 ( .A1(n3086), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3623) );
  NAND4_X1 U4566 ( .A1(n3626), .A2(n3625), .A3(n3624), .A4(n3623), .ZN(n3627)
         );
  NAND2_X1 U4567 ( .A1(n3730), .A2(n3643), .ZN(n3630) );
  NAND2_X1 U4568 ( .A1(n3713), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3629) );
  NAND2_X1 U4569 ( .A1(n3632), .A2(n3631), .ZN(n3939) );
  NAND3_X1 U4570 ( .A1(n3653), .A2(n3939), .A3(n3710), .ZN(n3639) );
  NAND2_X1 U4571 ( .A1(n3634), .A2(n3633), .ZN(n3635) );
  OR2_X1 U4572 ( .A1(n3636), .A2(n3635), .ZN(n3642) );
  XNOR2_X1 U4573 ( .A(n3642), .B(n3643), .ZN(n3637) );
  NAND2_X1 U4574 ( .A1(n3637), .A2(n5197), .ZN(n3638) );
  NAND2_X1 U4575 ( .A1(n3639), .A2(n3638), .ZN(n4820) );
  NAND2_X1 U4576 ( .A1(n3730), .A2(n3654), .ZN(n3641) );
  NAND2_X1 U4577 ( .A1(n3713), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3640) );
  INV_X1 U4578 ( .A(n3642), .ZN(n3644) );
  NAND2_X1 U4579 ( .A1(n3644), .A2(n3643), .ZN(n3656) );
  XNOR2_X1 U4580 ( .A(n3656), .B(n3654), .ZN(n3645) );
  NAND2_X1 U4581 ( .A1(n3645), .A2(n5197), .ZN(n3646) );
  XNOR2_X1 U4582 ( .A(n3650), .B(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6562)
         );
  NOR2_X1 U4583 ( .A1(n4820), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3648)
         );
  NOR2_X1 U4584 ( .A1(n6562), .A2(n3648), .ZN(n3649) );
  NAND2_X1 U4585 ( .A1(n3650), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3651)
         );
  AND2_X1 U4586 ( .A1(n3710), .A2(n3654), .ZN(n3652) );
  INV_X1 U4587 ( .A(n3654), .ZN(n3655) );
  OR3_X1 U4588 ( .A1(n3656), .A2(n3655), .A3(n3750), .ZN(n3657) );
  NAND2_X1 U4589 ( .A1(n3659), .A2(n3657), .ZN(n3658) );
  INV_X1 U4590 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6616) );
  XNOR2_X1 U4591 ( .A(n3658), .B(n6616), .ZN(n5849) );
  NAND2_X1 U4592 ( .A1(n3658), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5841)
         );
  INV_X1 U4593 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n7064) );
  OR2_X1 U4594 ( .A1(n3659), .A2(n7064), .ZN(n5843) );
  INV_X1 U4595 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5811) );
  INV_X1 U4596 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6031) );
  INV_X1 U4597 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6021) );
  AND3_X1 U4598 ( .A1(n5811), .A2(n6031), .A3(n6021), .ZN(n3660) );
  OR2_X1 U4599 ( .A1(n5815), .A2(n3660), .ZN(n3661) );
  NAND2_X1 U4600 ( .A1(n5824), .A2(n7064), .ZN(n5842) );
  NAND2_X1 U4601 ( .A1(n5824), .A2(n6021), .ZN(n5814) );
  NAND2_X1 U4602 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3663) );
  NAND2_X1 U4603 ( .A1(n5824), .A2(n3663), .ZN(n3664) );
  XNOR2_X1 U4604 ( .A(n5824), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5801)
         );
  INV_X1 U4605 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U4606 ( .A1(n5824), .A2(n5986), .ZN(n3667) );
  INV_X1 U4607 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5994) );
  NAND2_X1 U4608 ( .A1(n5813), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3669) );
  INV_X1 U4609 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n7023) );
  NAND2_X1 U4610 ( .A1(n5815), .A2(n7023), .ZN(n3670) );
  INV_X1 U4611 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n7058) );
  INV_X1 U4612 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5930) );
  INV_X1 U4613 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5950) );
  NAND3_X1 U4614 ( .A1(n7058), .A2(n5930), .A3(n5950), .ZN(n3671) );
  NAND2_X1 U4615 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3886) );
  INV_X1 U4616 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5935) );
  INV_X1 U4617 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5738) );
  XNOR2_X1 U4618 ( .A(n5824), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5730)
         );
  AND2_X1 U4619 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5217) );
  NAND4_X1 U4620 ( .A1(n5746), .A2(n5217), .A3(INSTADDRPOINTER_REG_20__SCAN_IN), .A4(n5824), .ZN(n3675) );
  INV_X1 U4621 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5032) );
  NOR2_X1 U4622 ( .A1(n3676), .A2(STATE_REG_0__SCAN_IN), .ZN(n4472) );
  INV_X1 U4623 ( .A(n4472), .ZN(n6798) );
  NAND2_X1 U4624 ( .A1(n3396), .A2(n6798), .ZN(n3697) );
  XNOR2_X1 U4625 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3688) );
  NAND2_X1 U4626 ( .A1(n3688), .A2(n3700), .ZN(n3678) );
  NAND2_X1 U4627 ( .A1(n4839), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3677) );
  NAND2_X1 U4628 ( .A1(n3678), .A2(n3677), .ZN(n3693) );
  XNOR2_X1 U4629 ( .A(n4952), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3692)
         );
  INV_X1 U4630 ( .A(n3692), .ZN(n3679) );
  NAND2_X1 U4631 ( .A1(n3693), .A2(n3679), .ZN(n3681) );
  NAND2_X1 U4632 ( .A1(n4489), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3680) );
  NAND2_X1 U4633 ( .A1(n3681), .A2(n3680), .ZN(n3691) );
  XNOR2_X1 U4634 ( .A(n4495), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3690)
         );
  INV_X1 U4635 ( .A(n3690), .ZN(n3682) );
  NAND2_X1 U4636 ( .A1(n3691), .A2(n3682), .ZN(n3684) );
  NAND2_X1 U4637 ( .A1(n6302), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3683) );
  NAND2_X1 U4638 ( .A1(n3684), .A2(n3683), .ZN(n3694) );
  INV_X1 U4639 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6659) );
  AND2_X1 U4640 ( .A1(n6659), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3685)
         );
  OR2_X1 U4641 ( .A1(n3694), .A2(n3685), .ZN(n3687) );
  INV_X1 U4642 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4512) );
  NAND2_X1 U4643 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n4512), .ZN(n3686) );
  INV_X1 U4644 ( .A(n3736), .ZN(n3696) );
  INV_X1 U4645 ( .A(n3700), .ZN(n3689) );
  XNOR2_X1 U4646 ( .A(n3689), .B(n3688), .ZN(n3711) );
  XNOR2_X1 U4647 ( .A(n3691), .B(n3690), .ZN(n3721) );
  XNOR2_X1 U4648 ( .A(n3693), .B(n3692), .ZN(n3715) );
  NAND4_X1 U4649 ( .A1(n3711), .A2(n3721), .A3(n3715), .A4(n3733), .ZN(n3695)
         );
  NAND2_X1 U4650 ( .A1(n3696), .A2(n3695), .ZN(n4293) );
  NOR2_X1 U4651 ( .A1(READY_N), .A2(n4293), .ZN(n4716) );
  NAND2_X1 U4652 ( .A1(n3697), .A2(n4716), .ZN(n3744) );
  NAND2_X1 U4653 ( .A1(n3730), .A2(n3396), .ZN(n3698) );
  NAND2_X1 U4654 ( .A1(n3698), .A2(n3745), .ZN(n3705) );
  AND2_X1 U4655 ( .A1(n3711), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3706) );
  NOR2_X1 U4656 ( .A1(n3700), .A2(n3699), .ZN(n3704) );
  AOI21_X1 U4657 ( .B1(n3759), .B2(n3704), .A(n3701), .ZN(n3703) );
  INV_X2 U4658 ( .A(n4279), .ZN(n5515) );
  NAND2_X1 U4659 ( .A1(n4413), .A2(n3745), .ZN(n3702) );
  NAND2_X1 U4660 ( .A1(n5515), .A2(n3702), .ZN(n3718) );
  OAI22_X1 U4661 ( .A1(n3705), .A2(n3706), .B1(n3703), .B2(n3718), .ZN(n3712)
         );
  NAND2_X1 U4662 ( .A1(n3730), .A2(n3704), .ZN(n3709) );
  INV_X1 U4663 ( .A(n3705), .ZN(n3708) );
  INV_X1 U4664 ( .A(n3706), .ZN(n3707) );
  NAND2_X1 U4665 ( .A1(n3730), .A2(n3715), .ZN(n3717) );
  INV_X1 U4666 ( .A(n3718), .ZN(n3714) );
  OAI211_X1 U4667 ( .C1(n3715), .C2(n3727), .A(n3717), .B(n3714), .ZN(n3716)
         );
  INV_X1 U4668 ( .A(n3717), .ZN(n3719) );
  NAND2_X1 U4669 ( .A1(n3719), .A2(n3718), .ZN(n3720) );
  INV_X1 U4670 ( .A(n3721), .ZN(n3723) );
  NAND2_X1 U4671 ( .A1(n3727), .A2(n3723), .ZN(n3722) );
  NAND2_X1 U4672 ( .A1(n3737), .A2(n3723), .ZN(n3724) );
  NAND2_X1 U4673 ( .A1(n3725), .A2(n3724), .ZN(n3729) );
  INV_X1 U4674 ( .A(n3733), .ZN(n3726) );
  NAND2_X1 U4675 ( .A1(n3727), .A2(n3726), .ZN(n3728) );
  NAND2_X1 U4676 ( .A1(n3730), .A2(n3736), .ZN(n3732) );
  NAND2_X1 U4677 ( .A1(n4531), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3731) );
  OAI211_X1 U4678 ( .C1(n3734), .C2(n3733), .A(n3732), .B(n3731), .ZN(n3735)
         );
  INV_X1 U4679 ( .A(READY_N), .ZN(n6800) );
  NAND2_X1 U4680 ( .A1(n3396), .A2(n6800), .ZN(n4334) );
  NAND2_X1 U4681 ( .A1(n4472), .A2(n6800), .ZN(n3740) );
  NAND2_X1 U4682 ( .A1(n4334), .A2(n3740), .ZN(n5189) );
  NAND2_X1 U4683 ( .A1(n3739), .A2(n5189), .ZN(n3741) );
  NAND3_X1 U4684 ( .A1(n3741), .A2(n5200), .A3(n3894), .ZN(n3742) );
  NAND2_X1 U4685 ( .A1(n4376), .A2(n3742), .ZN(n3743) );
  NAND2_X1 U4686 ( .A1(n3405), .A2(n3745), .ZN(n3746) );
  OR2_X1 U4687 ( .A1(n3867), .A2(n3746), .ZN(n3755) );
  NAND2_X1 U4688 ( .A1(n3748), .A2(n3747), .ZN(n3760) );
  NAND2_X1 U4689 ( .A1(n3749), .A2(n5200), .ZN(n3751) );
  MUX2_X1 U4690 ( .A(n3751), .B(n3750), .S(n3404), .Z(n3856) );
  INV_X1 U4691 ( .A(n3856), .ZN(n3754) );
  INV_X1 U4692 ( .A(n3752), .ZN(n3753) );
  OAI21_X1 U4693 ( .B1(n3760), .B2(n3754), .A(n3753), .ZN(n3843) );
  NAND2_X1 U4694 ( .A1(n4328), .A2(n3396), .ZN(n3844) );
  NAND3_X1 U4695 ( .A1(n3756), .A2(n3843), .A3(n4307), .ZN(n3758) );
  AND2_X1 U4696 ( .A1(n3757), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4737) );
  AND2_X2 U4697 ( .A1(n3758), .A2(n4737), .ZN(n3870) );
  OR2_X1 U4698 ( .A1(n3760), .A2(n5515), .ZN(n4714) );
  OR2_X1 U4699 ( .A1(n3760), .A2(n3759), .ZN(n4516) );
  AND2_X1 U4700 ( .A1(n4714), .A2(n4516), .ZN(n4291) );
  AOI22_X1 U4701 ( .A1(n4991), .A2(n3739), .B1(n3839), .B2(n3405), .ZN(n3761)
         );
  NAND3_X1 U4702 ( .A1(n4291), .A2(n3761), .A3(n4721), .ZN(n3762) );
  NAND2_X1 U4703 ( .A1(n3889), .A2(n6653), .ZN(n3888) );
  MUX2_X1 U4704 ( .A(n4980), .B(n3771), .S(EBX_REG_19__SCAN_IN), .Z(n3766) );
  NAND2_X1 U4705 ( .A1(n3764), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3765) );
  INV_X1 U4706 ( .A(n3771), .ZN(n3767) );
  NAND2_X1 U4707 ( .A1(n3767), .A2(n3764), .ZN(n3783) );
  NAND2_X1 U4708 ( .A1(n3764), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3768)
         );
  AND2_X1 U4709 ( .A1(n3783), .A2(n3768), .ZN(n3769) );
  NAND2_X1 U4710 ( .A1(n3771), .A2(EBX_REG_0__SCAN_IN), .ZN(n3773) );
  INV_X1 U4711 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4385) );
  NAND2_X1 U4712 ( .A1(n5050), .A2(n4385), .ZN(n3772) );
  NAND2_X1 U4713 ( .A1(n3773), .A2(n3772), .ZN(n4353) );
  XNOR2_X1 U4714 ( .A(n3774), .B(n4353), .ZN(n4382) );
  NAND2_X1 U4715 ( .A1(n4381), .A2(n3774), .ZN(n4467) );
  INV_X1 U4716 ( .A(EBX_REG_2__SCAN_IN), .ZN(n6468) );
  NAND2_X1 U4717 ( .A1(n3763), .A2(n6468), .ZN(n3778) );
  NAND2_X1 U4718 ( .A1(n3771), .A2(n6579), .ZN(n3776) );
  NAND2_X1 U4719 ( .A1(n4991), .A2(n6468), .ZN(n3775) );
  INV_X1 U4720 ( .A(EBX_REG_3__SCAN_IN), .ZN(n6992) );
  NAND2_X1 U4721 ( .A1(n3098), .A2(n6992), .ZN(n3781) );
  NAND2_X1 U4722 ( .A1(n5050), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3779)
         );
  OAI211_X1 U4723 ( .C1(n3764), .C2(EBX_REG_3__SCAN_IN), .A(n3771), .B(n3779), 
        .ZN(n3780) );
  NAND2_X1 U4724 ( .A1(n4468), .A2(n5534), .ZN(n5536) );
  MUX2_X1 U4725 ( .A(n4980), .B(n3771), .S(EBX_REG_4__SCAN_IN), .Z(n3785) );
  NAND2_X1 U4726 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n3764), .ZN(n3782)
         );
  AND2_X1 U4727 ( .A1(n3783), .A2(n3782), .ZN(n3784) );
  INV_X1 U4728 ( .A(n4537), .ZN(n3786) );
  INV_X1 U4729 ( .A(EBX_REG_6__SCAN_IN), .ZN(n3788) );
  NAND2_X1 U4730 ( .A1(n3763), .A2(n3788), .ZN(n3792) );
  INV_X1 U4731 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4819) );
  NAND2_X1 U4732 ( .A1(n3771), .A2(n4819), .ZN(n3790) );
  NAND2_X1 U4733 ( .A1(n4991), .A2(n3788), .ZN(n3789) );
  NAND2_X1 U4734 ( .A1(n3792), .A2(n3791), .ZN(n4775) );
  OAI211_X1 U4735 ( .C1(n3764), .C2(EBX_REG_7__SCAN_IN), .A(n3771), .B(n3793), 
        .ZN(n3794) );
  OAI21_X1 U4736 ( .B1(n4987), .B2(EBX_REG_7__SCAN_IN), .A(n3794), .ZN(n4886)
         );
  INV_X1 U4737 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6408) );
  NAND2_X1 U4738 ( .A1(n3763), .A2(n6408), .ZN(n3800) );
  NAND2_X1 U4739 ( .A1(n3771), .A2(n6616), .ZN(n3798) );
  NAND2_X1 U4740 ( .A1(n4991), .A2(n6408), .ZN(n3797) );
  NAND2_X1 U4741 ( .A1(n5050), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3801)
         );
  OAI211_X1 U4742 ( .C1(n3764), .C2(EBX_REG_9__SCAN_IN), .A(n3771), .B(n3801), 
        .ZN(n3802) );
  OAI21_X1 U4743 ( .B1(n4987), .B2(EBX_REG_9__SCAN_IN), .A(n3802), .ZN(n5596)
         );
  INV_X1 U4744 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5590) );
  NAND2_X1 U4745 ( .A1(n3763), .A2(n5590), .ZN(n3806) );
  NAND2_X1 U4746 ( .A1(n3771), .A2(n5811), .ZN(n3804) );
  NAND2_X1 U4747 ( .A1(n4991), .A2(n5590), .ZN(n3803) );
  NAND2_X1 U4748 ( .A1(n3806), .A2(n3805), .ZN(n5587) );
  INV_X1 U4749 ( .A(n3807), .ZN(n3809) );
  NOR2_X1 U4750 ( .A1(n4993), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3808)
         );
  NOR2_X1 U4751 ( .A1(n3809), .A2(n3808), .ZN(n5506) );
  INV_X1 U4752 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6475) );
  NAND2_X1 U4753 ( .A1(n3763), .A2(n6475), .ZN(n3813) );
  NAND2_X1 U4754 ( .A1(n3771), .A2(n6021), .ZN(n3811) );
  NAND2_X1 U4755 ( .A1(n4991), .A2(n6475), .ZN(n3810) );
  INV_X1 U4756 ( .A(n3814), .ZN(n5493) );
  NAND2_X1 U4757 ( .A1(n3815), .A2(n3286), .ZN(n5492) );
  OAI21_X1 U4758 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n4993), .A(n3816), 
        .ZN(n3817) );
  INV_X1 U4759 ( .A(n3817), .ZN(n5459) );
  INV_X1 U4760 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U4761 ( .A1(n3763), .A2(n5578), .ZN(n3821) );
  NAND2_X1 U4762 ( .A1(n3771), .A2(n5994), .ZN(n3819) );
  NAND2_X1 U4763 ( .A1(n4991), .A2(n5578), .ZN(n3818) );
  NAND2_X1 U4764 ( .A1(n3821), .A2(n3820), .ZN(n5478) );
  OAI21_X1 U4765 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n4993), .A(n3822), 
        .ZN(n5427) );
  INV_X1 U4766 ( .A(EBX_REG_16__SCAN_IN), .ZN(n3823) );
  NAND2_X1 U4767 ( .A1(n3763), .A2(n3823), .ZN(n3826) );
  NAND2_X1 U4768 ( .A1(n3771), .A2(n7058), .ZN(n3824) );
  INV_X1 U4769 ( .A(n4993), .ZN(n3847) );
  NOR2_X1 U4770 ( .A1(n3764), .A2(EBX_REG_20__SCAN_IN), .ZN(n3827) );
  AOI21_X1 U4771 ( .B1(n3847), .B2(n5738), .A(n3827), .ZN(n5381) );
  OR2_X1 U4772 ( .A1(n4993), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3828)
         );
  INV_X1 U4773 ( .A(EBX_REG_18__SCAN_IN), .ZN(n7101) );
  NAND2_X1 U4774 ( .A1(n4991), .A2(n7101), .ZN(n5390) );
  NAND2_X1 U4775 ( .A1(n3828), .A2(n5390), .ZN(n5391) );
  NAND2_X1 U4776 ( .A1(n5389), .A2(EBX_REG_20__SCAN_IN), .ZN(n3830) );
  NAND2_X1 U4777 ( .A1(n5391), .A2(n5050), .ZN(n3829) );
  OAI211_X1 U4778 ( .C1(n5381), .C2(n5391), .A(n3830), .B(n3829), .ZN(n3831)
         );
  INV_X1 U4779 ( .A(n3831), .ZN(n3832) );
  MUX2_X1 U4780 ( .A(n4980), .B(n3771), .S(EBX_REG_21__SCAN_IN), .Z(n3834) );
  NAND2_X1 U4781 ( .A1(n3764), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3833) );
  NAND2_X1 U4782 ( .A1(n3834), .A2(n3833), .ZN(n5372) );
  MUX2_X1 U4783 ( .A(n4987), .B(n5050), .S(EBX_REG_22__SCAN_IN), .Z(n3835) );
  OAI21_X1 U4784 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n4993), .A(n3835), 
        .ZN(n3836) );
  INV_X1 U4785 ( .A(n3836), .ZN(n5350) );
  MUX2_X1 U4786 ( .A(n4980), .B(n3771), .S(EBX_REG_23__SCAN_IN), .Z(n3838) );
  NAND2_X1 U4787 ( .A1(n3764), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3837) );
  NAND2_X1 U4788 ( .A1(n3838), .A2(n3837), .ZN(n5026) );
  XNOR2_X1 U4789 ( .A(n5349), .B(n5026), .ZN(n5569) );
  NAND2_X1 U4790 ( .A1(n3739), .A2(n5197), .ZN(n4530) );
  NAND2_X1 U4791 ( .A1(n3839), .A2(n4717), .ZN(n3840) );
  NAND2_X1 U4792 ( .A1(n4530), .A2(n3840), .ZN(n3841) );
  OR2_X1 U4793 ( .A1(n3842), .A2(n3851), .ZN(n3846) );
  NAND2_X1 U4794 ( .A1(n3843), .A2(n3846), .ZN(n4304) );
  INV_X1 U4795 ( .A(n4473), .ZN(n3845) );
  NAND2_X1 U4796 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6037) );
  NAND2_X1 U4797 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6036) );
  NOR2_X1 U4798 ( .A1(n6037), .A2(n6036), .ZN(n3872) );
  AOI21_X1 U4799 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6644) );
  NAND2_X1 U4800 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6645) );
  NOR2_X1 U4801 ( .A1(n6644), .A2(n6645), .ZN(n6624) );
  NAND2_X1 U4802 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6624), .ZN(n4829)
         );
  NOR2_X1 U4803 ( .A1(n4819), .A2(n4829), .ZN(n6039) );
  AND2_X1 U4804 ( .A1(n3872), .A2(n6039), .ZN(n3883) );
  NAND2_X1 U4805 ( .A1(n3847), .A2(n3846), .ZN(n3849) );
  NAND2_X1 U4806 ( .A1(n3849), .A2(n3848), .ZN(n3855) );
  NAND2_X1 U4807 ( .A1(n3850), .A2(n5389), .ZN(n3853) );
  NAND2_X1 U4808 ( .A1(n3894), .A2(n3851), .ZN(n3852) );
  AND4_X1 U4809 ( .A1(n3855), .A2(n3854), .A3(n3853), .A4(n3852), .ZN(n3858)
         );
  AND3_X1 U4810 ( .A1(n3858), .A2(n3857), .A3(n3856), .ZN(n4313) );
  NAND2_X1 U4811 ( .A1(n4328), .A2(n3860), .ZN(n4500) );
  INV_X1 U4812 ( .A(n4719), .ZN(n3861) );
  NAND2_X1 U4813 ( .A1(n3861), .A2(n3913), .ZN(n3862) );
  OAI211_X1 U4814 ( .C1(n3859), .C2(n5200), .A(n4500), .B(n3862), .ZN(n3863)
         );
  INV_X1 U4815 ( .A(n3863), .ZN(n3864) );
  NAND2_X1 U4816 ( .A1(n4313), .A2(n3864), .ZN(n3865) );
  NAND2_X1 U4817 ( .A1(n3870), .A2(n3865), .ZN(n4352) );
  OR2_X1 U4818 ( .A1(n4352), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3866)
         );
  OR2_X1 U4819 ( .A1(n6805), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6639) );
  OR2_X1 U4820 ( .A1(n3870), .A2(n6577), .ZN(n4355) );
  NAND2_X1 U4821 ( .A1(n3866), .A2(n4355), .ZN(n6043) );
  INV_X1 U4822 ( .A(n6043), .ZN(n3874) );
  NAND2_X1 U4823 ( .A1(n5516), .A2(n3867), .ZN(n3868) );
  NOR2_X1 U4824 ( .A1(n3869), .A2(n3868), .ZN(n4498) );
  NAND2_X1 U4825 ( .A1(n3870), .A2(n4498), .ZN(n6004) );
  NAND4_X1 U4826 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(INSTADDRPOINTER_REG_3__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6627) );
  NOR3_X1 U4827 ( .A1(n3871), .A2(n4819), .A3(n6627), .ZN(n6040) );
  NAND2_X1 U4828 ( .A1(n6040), .A2(n3872), .ZN(n6003) );
  INV_X1 U4829 ( .A(n6003), .ZN(n5984) );
  OR2_X1 U4830 ( .A1(n6041), .A2(n5984), .ZN(n3873) );
  OAI211_X1 U4831 ( .C1(n6038), .C2(n3883), .A(n3874), .B(n3873), .ZN(n6026)
         );
  AND2_X1 U4832 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U4833 ( .A1(n5990), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U4834 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3875) );
  NOR2_X1 U4835 ( .A1(n5968), .A2(n3875), .ZN(n5963) );
  NAND2_X1 U4836 ( .A1(n5963), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3884) );
  AND2_X1 U4837 ( .A1(n5967), .A2(n3884), .ZN(n3876) );
  INV_X1 U4838 ( .A(n3886), .ZN(n3877) );
  AND2_X1 U4839 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5925) );
  NAND2_X1 U4840 ( .A1(n3877), .A2(n5925), .ZN(n3878) );
  AND2_X1 U4841 ( .A1(n5967), .A2(n3878), .ZN(n3879) );
  NOR2_X1 U4842 ( .A1(n5959), .A2(n3879), .ZN(n5906) );
  INV_X1 U4843 ( .A(n5217), .ZN(n5911) );
  NAND2_X1 U4844 ( .A1(n5967), .A2(n5911), .ZN(n3880) );
  NAND2_X1 U4845 ( .A1(n5906), .A2(n3880), .ZN(n5030) );
  NAND2_X1 U4846 ( .A1(n5030), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3881) );
  NAND2_X1 U4847 ( .A1(n6577), .A2(REIP_REG_23__SCAN_IN), .ZN(n4240) );
  NAND2_X1 U4848 ( .A1(n3881), .A2(n4240), .ZN(n3882) );
  AOI21_X1 U4849 ( .B1(n5569), .B2(n6651), .A(n3882), .ZN(n3887) );
  INV_X1 U4850 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6838) );
  NAND2_X1 U4851 ( .A1(n6838), .A2(n6004), .ZN(n4960) );
  NOR2_X1 U4852 ( .A1(n6628), .A2(n6003), .ZN(n5929) );
  INV_X1 U4853 ( .A(n3884), .ZN(n3885) );
  NAND2_X1 U4854 ( .A1(n5936), .A2(n5925), .ZN(n5923) );
  NAND2_X1 U4855 ( .A1(n3888), .A2(n3284), .ZN(U2995) );
  NOR2_X2 U4856 ( .A1(n3398), .A2(n6673), .ZN(n4116) );
  NAND2_X1 U4857 ( .A1(n3890), .A2(n4116), .ZN(n3899) );
  OR2_X1 U4858 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n5165) );
  INV_X1 U4859 ( .A(n3900), .ZN(n3893) );
  INV_X1 U4860 ( .A(n3933), .ZN(n3892) );
  OAI21_X1 U4861 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n3893), .A(n3892), 
        .ZN(n5527) );
  INV_X1 U4862 ( .A(n3894), .ZN(n4728) );
  AND2_X1 U4863 ( .A1(n4728), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3916) );
  INV_X1 U4864 ( .A(n3916), .ZN(n3925) );
  NAND2_X1 U4865 ( .A1(n4168), .A2(EAX_REG_4__SCAN_IN), .ZN(n3896) );
  INV_X1 U4866 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6361) );
  OAI21_X1 U4867 ( .B1(n6361), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6673), 
        .ZN(n3895) );
  OAI211_X1 U4868 ( .C1(n3925), .C2(n4512), .A(n3896), .B(n3895), .ZN(n3897)
         );
  OAI21_X1 U4869 ( .B1(n5165), .B2(n5527), .A(n3897), .ZN(n3898) );
  NAND2_X1 U4870 ( .A1(n3899), .A2(n3898), .ZN(n4533) );
  NAND2_X1 U4871 ( .A1(n4542), .A2(n4116), .ZN(n3906) );
  INV_X2 U4872 ( .A(n5165), .ZN(n5182) );
  OAI21_X1 U4873 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3901), .A(n3900), 
        .ZN(n6588) );
  AND2_X1 U4874 ( .A1(n6673), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5245) );
  AOI22_X1 U4875 ( .A1(n5182), .A2(n6588), .B1(n5245), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3903) );
  NAND2_X1 U4876 ( .A1(n4168), .A2(EAX_REG_3__SCAN_IN), .ZN(n3902) );
  OAI211_X1 U4877 ( .C1(n3925), .C2(n4495), .A(n3903), .B(n3902), .ZN(n3904)
         );
  INV_X1 U4878 ( .A(n3904), .ZN(n3905) );
  NAND2_X1 U4879 ( .A1(n3906), .A2(n3905), .ZN(n4883) );
  NAND2_X1 U4880 ( .A1(n4387), .A2(n4116), .ZN(n3911) );
  AOI22_X1 U4881 ( .A1(n4168), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6673), .ZN(n3909) );
  NAND2_X1 U4882 ( .A1(n3916), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3908) );
  AND2_X1 U4883 ( .A1(n3909), .A2(n3908), .ZN(n3910) );
  NAND2_X1 U4884 ( .A1(n3911), .A2(n3910), .ZN(n4380) );
  NAND2_X1 U4885 ( .A1(n3912), .A2(n3913), .ZN(n3914) );
  NAND2_X1 U4886 ( .A1(n3914), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4342) );
  INV_X1 U4887 ( .A(n4116), .ZN(n3970) );
  OR2_X1 U4888 ( .A1(n3915), .A2(n3970), .ZN(n3920) );
  AOI22_X1 U4889 ( .A1(n4168), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6673), .ZN(n3918) );
  NAND2_X1 U4890 ( .A1(n3916), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3917) );
  AND2_X1 U4891 ( .A1(n3918), .A2(n3917), .ZN(n3919) );
  NAND2_X1 U4892 ( .A1(n4341), .A2(n5182), .ZN(n3921) );
  NAND2_X1 U4893 ( .A1(n4344), .A2(n3921), .ZN(n4379) );
  NAND2_X1 U4894 ( .A1(n4380), .A2(n4379), .ZN(n4378) );
  NAND2_X1 U4895 ( .A1(n3926), .A2(n4378), .ZN(n4464) );
  OAI21_X1 U4896 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3922), .ZN(n6598) );
  AOI22_X1 U4897 ( .A1(n5245), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n5182), 
        .B2(n6598), .ZN(n3924) );
  NAND2_X1 U4898 ( .A1(n4168), .A2(EAX_REG_2__SCAN_IN), .ZN(n3923) );
  OAI211_X1 U4899 ( .C1(n3925), .C2(n4952), .A(n3924), .B(n3923), .ZN(n4463)
         );
  NAND2_X1 U4900 ( .A1(n4464), .A2(n4463), .ZN(n3930) );
  INV_X1 U4901 ( .A(n4378), .ZN(n3928) );
  INV_X1 U4902 ( .A(n3926), .ZN(n3927) );
  NAND2_X1 U4903 ( .A1(n3928), .A2(n3927), .ZN(n3929) );
  NAND2_X1 U4904 ( .A1(n3932), .A2(n4116), .ZN(n3938) );
  INV_X1 U4905 ( .A(n5245), .ZN(n3954) );
  INV_X1 U4906 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3935) );
  OAI21_X1 U4907 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n3933), .A(n3948), 
        .ZN(n6576) );
  NAND2_X1 U4908 ( .A1(n6576), .A2(n5182), .ZN(n3934) );
  OAI21_X1 U4909 ( .B1(n3954), .B2(n3935), .A(n3934), .ZN(n3936) );
  AOI21_X1 U4910 ( .B1(n4168), .B2(EAX_REG_5__SCAN_IN), .A(n3936), .ZN(n3937)
         );
  NAND2_X1 U4911 ( .A1(n3939), .A2(n4116), .ZN(n3945) );
  INV_X1 U4912 ( .A(EAX_REG_6__SCAN_IN), .ZN(n3941) );
  OAI21_X1 U4913 ( .B1(n6361), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6673), 
        .ZN(n3940) );
  OAI21_X1 U4914 ( .B1(n3290), .B2(n3941), .A(n3940), .ZN(n3943) );
  XNOR2_X1 U4915 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .B(n3948), .ZN(n6428) );
  NAND2_X1 U4916 ( .A1(n6428), .A2(n5182), .ZN(n3942) );
  NAND2_X1 U4917 ( .A1(n3943), .A2(n3942), .ZN(n3944) );
  NAND2_X1 U4918 ( .A1(n3945), .A2(n3944), .ZN(n4771) );
  INV_X1 U4919 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3953) );
  OR2_X1 U4920 ( .A1(n3949), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3950) );
  NAND2_X1 U4921 ( .A1(n3950), .A2(n3971), .ZN(n6569) );
  NAND2_X1 U4922 ( .A1(n6569), .A2(n5182), .ZN(n3952) );
  NAND2_X1 U4923 ( .A1(n4168), .A2(EAX_REG_7__SCAN_IN), .ZN(n3951) );
  OAI211_X1 U4924 ( .C1(n3954), .C2(n3953), .A(n3952), .B(n3951), .ZN(n3955)
         );
  AOI22_X1 U4925 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n3496), .B1(n5116), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U4926 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n5124), .B1(n5107), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3958) );
  AOI22_X1 U4927 ( .A1(n5122), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3087), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U4928 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n3488), .B1(n5114), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3956) );
  NAND4_X1 U4929 ( .A1(n3959), .A2(n3958), .A3(n3957), .A4(n3956), .ZN(n3965)
         );
  AOI22_X1 U4930 ( .A1(n5121), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3468), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U4931 ( .A1(n5123), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3486), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3962) );
  AOI22_X1 U4932 ( .A1(n3461), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n5115), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U4933 ( .A1(n3086), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3960) );
  NAND4_X1 U4934 ( .A1(n3963), .A2(n3962), .A3(n3961), .A4(n3960), .ZN(n3964)
         );
  NOR2_X1 U4935 ( .A1(n3965), .A2(n3964), .ZN(n3969) );
  XNOR2_X1 U4936 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3971), .ZN(n6411) );
  INV_X1 U4937 ( .A(n6411), .ZN(n3966) );
  AOI22_X1 U4938 ( .A1(n5245), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n5182), 
        .B2(n3966), .ZN(n3968) );
  NAND2_X1 U4939 ( .A1(n4168), .A2(EAX_REG_8__SCAN_IN), .ZN(n3967) );
  OAI211_X1 U4940 ( .C1(n3970), .C2(n3969), .A(n3968), .B(n3967), .ZN(n5600)
         );
  INV_X1 U4941 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6401) );
  NAND2_X1 U4942 ( .A1(PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3973) );
  AND2_X1 U4943 ( .A1(PHYADDRPOINTER_REG_14__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3974) );
  INV_X1 U4944 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5769) );
  INV_X1 U4945 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5760) );
  INV_X1 U4946 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3976) );
  OAI21_X1 U4947 ( .B1(n4137), .B2(n5760), .A(n3976), .ZN(n3978) );
  NAND2_X1 U4948 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3977) );
  NAND2_X1 U4949 ( .A1(n3978), .A2(n4155), .ZN(n5752) );
  AOI22_X1 U4950 ( .A1(n4192), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3468), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3982) );
  AOI22_X1 U4951 ( .A1(n5123), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U4952 ( .A1(n3462), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n5114), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3980) );
  AOI22_X1 U4953 ( .A1(n3461), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3087), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3979) );
  NAND4_X1 U4954 ( .A1(n3982), .A2(n3981), .A3(n3980), .A4(n3979), .ZN(n3988)
         );
  AOI22_X1 U4955 ( .A1(n5107), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5124), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3986) );
  AOI22_X1 U4956 ( .A1(n5121), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3985) );
  AOI22_X1 U4957 ( .A1(n5122), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n5115), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3984) );
  AOI22_X1 U4958 ( .A1(n3496), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3983) );
  NAND4_X1 U4959 ( .A1(n3986), .A2(n3985), .A3(n3984), .A4(n3983), .ZN(n3987)
         );
  NOR2_X1 U4960 ( .A1(n3988), .A2(n3987), .ZN(n3990) );
  AOI22_X1 U4961 ( .A1(n4168), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6673), .ZN(n3989) );
  OAI21_X1 U4962 ( .B1(n5177), .B2(n3990), .A(n3989), .ZN(n3991) );
  MUX2_X1 U4963 ( .A(n5752), .B(n3991), .S(n5165), .Z(n5396) );
  NAND2_X1 U4964 ( .A1(n3992), .A2(n5769), .ZN(n3993) );
  AND2_X1 U4965 ( .A1(n4137), .A2(n3993), .ZN(n5771) );
  INV_X1 U4966 ( .A(n5177), .ZN(n5155) );
  AOI22_X1 U4967 ( .A1(n5121), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n5107), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3997) );
  AOI22_X1 U4968 ( .A1(n4192), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3468), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U4969 ( .A1(n5123), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U4970 ( .A1(n5122), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3994) );
  NAND4_X1 U4971 ( .A1(n3997), .A2(n3996), .A3(n3995), .A4(n3994), .ZN(n4003)
         );
  AOI22_X1 U4972 ( .A1(n3086), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4001) );
  AOI22_X1 U4973 ( .A1(n3496), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U4974 ( .A1(n5115), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n5114), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U4975 ( .A1(n5124), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3087), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3998) );
  NAND4_X1 U4976 ( .A1(n4001), .A2(n4000), .A3(n3999), .A4(n3998), .ZN(n4002)
         );
  OR2_X1 U4977 ( .A1(n4003), .A2(n4002), .ZN(n4006) );
  INV_X1 U4978 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4004) );
  OAI22_X1 U4979 ( .A1(n3290), .A2(n4004), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5769), .ZN(n4005) );
  AOI21_X1 U4980 ( .B1(n5155), .B2(n4006), .A(n4005), .ZN(n4007) );
  MUX2_X1 U4981 ( .A(n5771), .B(n4007), .S(n5165), .Z(n4008) );
  INV_X1 U4982 ( .A(n4008), .ZN(n5425) );
  NAND2_X1 U4983 ( .A1(n4036), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4009)
         );
  INV_X1 U4984 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5462) );
  XNOR2_X1 U4985 ( .A(n4009), .B(n5462), .ZN(n5789) );
  AOI22_X1 U4986 ( .A1(n5107), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5124), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U4987 ( .A1(n3086), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U4988 ( .A1(n5115), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n5114), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U4989 ( .A1(n4192), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3089), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4010) );
  NAND4_X1 U4990 ( .A1(n4013), .A2(n4012), .A3(n4011), .A4(n4010), .ZN(n4019)
         );
  AOI22_X1 U4991 ( .A1(n5122), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5121), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U4992 ( .A1(n3496), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5123), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4016) );
  AOI22_X1 U4993 ( .A1(n3436), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3468), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U4994 ( .A1(n3488), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4014) );
  NAND4_X1 U4995 ( .A1(n4017), .A2(n4016), .A3(n4015), .A4(n4014), .ZN(n4018)
         );
  OAI21_X1 U4996 ( .B1(n4019), .B2(n4018), .A(n4116), .ZN(n4022) );
  NAND2_X1 U4997 ( .A1(n4168), .A2(EAX_REG_15__SCAN_IN), .ZN(n4021) );
  NAND2_X1 U4998 ( .A1(n5245), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4020)
         );
  NAND3_X1 U4999 ( .A1(n4022), .A2(n4021), .A3(n4020), .ZN(n4023) );
  AOI21_X1 U5000 ( .B1(n5789), .B2(n5182), .A(n4023), .ZN(n5457) );
  AOI22_X1 U5001 ( .A1(n5121), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n5123), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4027) );
  AOI22_X1 U5002 ( .A1(n3086), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3468), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4026) );
  AOI22_X1 U5003 ( .A1(n3462), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n5114), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4025) );
  AOI22_X1 U5004 ( .A1(n5124), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n5115), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4024) );
  NAND4_X1 U5005 ( .A1(n4027), .A2(n4026), .A3(n4025), .A4(n4024), .ZN(n4033)
         );
  AOI22_X1 U5006 ( .A1(n5122), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n5107), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U5007 ( .A1(n3496), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4030) );
  AOI22_X1 U5008 ( .A1(n4192), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4029) );
  AOI22_X1 U5009 ( .A1(n3469), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3087), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4028) );
  NAND4_X1 U5010 ( .A1(n4031), .A2(n4030), .A3(n4029), .A4(n4028), .ZN(n4032)
         );
  OR2_X1 U5011 ( .A1(n4033), .A2(n4032), .ZN(n4034) );
  AND2_X1 U5012 ( .A1(n4116), .A2(n4034), .ZN(n5490) );
  INV_X1 U5013 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5818) );
  INV_X1 U5014 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4035) );
  OAI21_X1 U5015 ( .B1(n4057), .B2(n5818), .A(n4035), .ZN(n4037) );
  INV_X1 U5016 ( .A(n4036), .ZN(n4041) );
  NAND2_X1 U5017 ( .A1(n4037), .A2(n4041), .ZN(n5804) );
  NAND2_X1 U5018 ( .A1(n5804), .A2(n5182), .ZN(n4039) );
  AOI22_X1 U5019 ( .A1(n4168), .A2(EAX_REG_13__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n5245), .ZN(n4038) );
  NAND2_X1 U5020 ( .A1(n4039), .A2(n4038), .ZN(n5454) );
  INV_X1 U5021 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4040) );
  XNOR2_X1 U5022 ( .A(n4041), .B(n4040), .ZN(n5796) );
  NAND2_X1 U5023 ( .A1(n5796), .A2(n5182), .ZN(n4055) );
  AOI22_X1 U5024 ( .A1(n5121), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4045) );
  AOI22_X1 U5025 ( .A1(n5124), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U5026 ( .A1(n3461), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3089), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U5027 ( .A1(n5114), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4042) );
  NAND4_X1 U5028 ( .A1(n4045), .A2(n4044), .A3(n4043), .A4(n4042), .ZN(n4051)
         );
  AOI22_X1 U5029 ( .A1(n5107), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3468), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4049) );
  AOI22_X1 U5030 ( .A1(n4192), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5123), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4048) );
  AOI22_X1 U5031 ( .A1(n3496), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4047) );
  AOI22_X1 U5032 ( .A1(n5122), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5115), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4046) );
  NAND4_X1 U5033 ( .A1(n4049), .A2(n4048), .A3(n4047), .A4(n4046), .ZN(n4050)
         );
  OAI21_X1 U5034 ( .B1(n4051), .B2(n4050), .A(n4116), .ZN(n4054) );
  NAND2_X1 U5035 ( .A1(n4168), .A2(EAX_REG_14__SCAN_IN), .ZN(n4053) );
  NAND2_X1 U5036 ( .A1(n5245), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4052)
         );
  NAND2_X1 U5037 ( .A1(n4055), .A2(n3285), .ZN(n5472) );
  OAI21_X1 U5038 ( .B1(n5490), .B2(n5454), .A(n5472), .ZN(n4056) );
  NOR2_X1 U5039 ( .A1(n5457), .A2(n4056), .ZN(n4106) );
  XNOR2_X1 U5040 ( .A(n4057), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6378)
         );
  NAND2_X1 U5041 ( .A1(n6378), .A2(n5182), .ZN(n4061) );
  INV_X1 U5042 ( .A(EAX_REG_12__SCAN_IN), .ZN(n4059) );
  OAI21_X1 U5043 ( .B1(PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n6361), .A(n6673), 
        .ZN(n4058) );
  OAI21_X1 U5044 ( .B1(n3290), .B2(n4059), .A(n4058), .ZN(n4060) );
  NAND2_X1 U5045 ( .A1(n4061), .A2(n4060), .ZN(n4073) );
  AOI22_X1 U5046 ( .A1(n5123), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4075), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U5047 ( .A1(n5122), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4064) );
  AOI22_X1 U5048 ( .A1(n5121), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4063) );
  AOI22_X1 U5049 ( .A1(n5114), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4062) );
  NAND4_X1 U5050 ( .A1(n4065), .A2(n4064), .A3(n4063), .A4(n4062), .ZN(n4071)
         );
  AOI22_X1 U5051 ( .A1(n4192), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n5107), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4069) );
  AOI22_X1 U5052 ( .A1(n3496), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4068) );
  AOI22_X1 U5053 ( .A1(n3468), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4067) );
  AOI22_X1 U5054 ( .A1(n3462), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n5115), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4066) );
  NAND4_X1 U5055 ( .A1(n4069), .A2(n4068), .A3(n4067), .A4(n4066), .ZN(n4070)
         );
  OAI21_X1 U5056 ( .B1(n4071), .B2(n4070), .A(n4116), .ZN(n4072) );
  NAND2_X1 U5057 ( .A1(n4073), .A2(n4072), .ZN(n5654) );
  INV_X1 U5058 ( .A(n5654), .ZN(n4105) );
  XNOR2_X1 U5059 ( .A(n4074), .B(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5828)
         );
  AOI22_X1 U5060 ( .A1(n5107), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4075), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4079) );
  AOI22_X1 U5061 ( .A1(n3468), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4078) );
  AOI22_X1 U5062 ( .A1(n4192), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3087), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4077) );
  AOI22_X1 U5063 ( .A1(n3436), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4076) );
  NAND4_X1 U5064 ( .A1(n4079), .A2(n4078), .A3(n4077), .A4(n4076), .ZN(n4085)
         );
  AOI22_X1 U5065 ( .A1(n5122), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4083) );
  AOI22_X1 U5066 ( .A1(n5123), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4082) );
  AOI22_X1 U5067 ( .A1(n5121), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n5114), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4081) );
  AOI22_X1 U5068 ( .A1(n3496), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5115), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4080) );
  NAND4_X1 U5069 ( .A1(n4083), .A2(n4082), .A3(n4081), .A4(n4080), .ZN(n4084)
         );
  OAI21_X1 U5070 ( .B1(n4085), .B2(n4084), .A(n4116), .ZN(n4088) );
  NAND2_X1 U5071 ( .A1(n4168), .A2(EAX_REG_11__SCAN_IN), .ZN(n4087) );
  NAND2_X1 U5072 ( .A1(n5245), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4086)
         );
  NAND3_X1 U5073 ( .A1(n4088), .A2(n4087), .A3(n4086), .ZN(n4089) );
  AOI21_X1 U5074 ( .B1(n5828), .B2(n5182), .A(n4089), .ZN(n5503) );
  AOI22_X1 U5075 ( .A1(n3496), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5116), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4093) );
  AOI22_X1 U5076 ( .A1(n5107), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3468), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4092) );
  AOI22_X1 U5077 ( .A1(n5122), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4091) );
  AOI22_X1 U5078 ( .A1(n5114), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4090) );
  NAND4_X1 U5079 ( .A1(n4093), .A2(n4092), .A3(n4091), .A4(n4090), .ZN(n4099)
         );
  AOI22_X1 U5080 ( .A1(n5124), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4097) );
  AOI22_X1 U5081 ( .A1(n5123), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4096) );
  AOI22_X1 U5082 ( .A1(n5121), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4095) );
  AOI22_X1 U5083 ( .A1(n3462), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n5115), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4094) );
  NAND4_X1 U5084 ( .A1(n4097), .A2(n4096), .A3(n4095), .A4(n4094), .ZN(n4098)
         );
  OAI21_X1 U5085 ( .B1(n4099), .B2(n4098), .A(n4116), .ZN(n4104) );
  INV_X1 U5086 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4101) );
  XNOR2_X1 U5087 ( .A(n4101), .B(n4100), .ZN(n6385) );
  INV_X1 U5088 ( .A(n6385), .ZN(n5837) );
  AOI22_X1 U5089 ( .A1(PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n5245), .B1(n5182), 
        .B2(n5837), .ZN(n4103) );
  NAND2_X1 U5090 ( .A1(n4168), .A2(EAX_REG_10__SCAN_IN), .ZN(n4102) );
  AND3_X1 U5091 ( .A1(n4104), .A2(n4103), .A3(n4102), .ZN(n5584) );
  OR2_X1 U5092 ( .A1(n5503), .A2(n5584), .ZN(n5502) );
  NOR2_X1 U5093 ( .A1(n4105), .A2(n5502), .ZN(n5451) );
  AND2_X1 U5094 ( .A1(n4106), .A2(n5451), .ZN(n4121) );
  XNOR2_X1 U5095 ( .A(n4107), .B(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6399) );
  AOI22_X1 U5096 ( .A1(n4168), .A2(EAX_REG_9__SCAN_IN), .B1(n5245), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4120) );
  AOI22_X1 U5097 ( .A1(n5121), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n5107), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4111) );
  AOI22_X1 U5098 ( .A1(n4192), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5114), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4110) );
  AOI22_X1 U5099 ( .A1(n5122), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3089), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4109) );
  AOI22_X1 U5100 ( .A1(n3436), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4108) );
  NAND4_X1 U5101 ( .A1(n4111), .A2(n4110), .A3(n4109), .A4(n4108), .ZN(n4118)
         );
  AOI22_X1 U5102 ( .A1(n3496), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3468), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4115) );
  AOI22_X1 U5103 ( .A1(n5123), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4114) );
  AOI22_X1 U5104 ( .A1(n5124), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4113) );
  AOI22_X1 U5105 ( .A1(n3462), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n5115), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4112) );
  NAND4_X1 U5106 ( .A1(n4115), .A2(n4114), .A3(n4113), .A4(n4112), .ZN(n4117)
         );
  OAI21_X1 U5107 ( .B1(n4118), .B2(n4117), .A(n4116), .ZN(n4119) );
  OAI211_X1 U5108 ( .C1(n6399), .C2(n5165), .A(n4120), .B(n4119), .ZN(n5594)
         );
  AND2_X1 U5109 ( .A1(n4121), .A2(n5594), .ZN(n5438) );
  INV_X1 U5110 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5778) );
  XNOR2_X1 U5111 ( .A(n4122), .B(n5778), .ZN(n5781) );
  AOI22_X1 U5112 ( .A1(n5123), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4126) );
  AOI22_X1 U5113 ( .A1(n3086), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3488), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4125) );
  AOI22_X1 U5114 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n5122), .B1(n5114), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4124) );
  AOI22_X1 U5115 ( .A1(n5121), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3087), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4123) );
  NAND4_X1 U5116 ( .A1(n4126), .A2(n4125), .A3(n4124), .A4(n4123), .ZN(n4132)
         );
  AOI22_X1 U5117 ( .A1(n5107), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n5124), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4130) );
  AOI22_X1 U5118 ( .A1(n3496), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4129) );
  AOI22_X1 U5119 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n3467), .B1(n5115), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4128) );
  AOI22_X1 U5120 ( .A1(n4192), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4127) );
  NAND4_X1 U5121 ( .A1(n4130), .A2(n4129), .A3(n4128), .A4(n4127), .ZN(n4131)
         );
  NOR2_X1 U5122 ( .A1(n4132), .A2(n4131), .ZN(n4134) );
  AOI22_X1 U5123 ( .A1(n4168), .A2(EAX_REG_16__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n5245), .ZN(n4133) );
  OAI21_X1 U5124 ( .B1(n5177), .B2(n4134), .A(n4133), .ZN(n4135) );
  AOI21_X1 U5125 ( .B1(n5781), .B2(n5182), .A(n4135), .ZN(n5439) );
  INV_X1 U5126 ( .A(n5439), .ZN(n4136) );
  AND2_X1 U5127 ( .A1(n5438), .A2(n4136), .ZN(n5423) );
  XNOR2_X1 U5128 ( .A(n4137), .B(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5758)
         );
  NAND2_X1 U5129 ( .A1(n5758), .A2(n5182), .ZN(n4152) );
  AOI22_X1 U5130 ( .A1(n5121), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n5107), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4141) );
  AOI22_X1 U5131 ( .A1(n4192), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n5124), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4140) );
  AOI22_X1 U5132 ( .A1(n3467), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4139) );
  AOI22_X1 U5133 ( .A1(n5122), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4138) );
  NAND4_X1 U5134 ( .A1(n4141), .A2(n4140), .A3(n4139), .A4(n4138), .ZN(n4147)
         );
  AOI22_X1 U5135 ( .A1(n3496), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4145) );
  AOI22_X1 U5136 ( .A1(n5123), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n5114), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4144) );
  AOI22_X1 U5137 ( .A1(n3462), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n5115), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4143) );
  AOI22_X1 U5138 ( .A1(n3086), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4142) );
  NAND4_X1 U5139 ( .A1(n4145), .A2(n4144), .A3(n4143), .A4(n4142), .ZN(n4146)
         );
  NOR2_X1 U5140 ( .A1(n4147), .A2(n4146), .ZN(n4150) );
  AOI21_X1 U5141 ( .B1(n5760), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4148) );
  AOI21_X1 U5142 ( .B1(n4168), .B2(EAX_REG_18__SCAN_IN), .A(n4148), .ZN(n4149)
         );
  OAI21_X1 U5143 ( .B1(n5177), .B2(n4150), .A(n4149), .ZN(n4151) );
  NAND2_X1 U5144 ( .A1(n4152), .A2(n4151), .ZN(n5412) );
  INV_X1 U5145 ( .A(n5412), .ZN(n4153) );
  INV_X1 U5146 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6966) );
  NAND2_X1 U5147 ( .A1(n4155), .A2(n6966), .ZN(n4156) );
  NAND2_X1 U5148 ( .A1(n4189), .A2(n4156), .ZN(n5742) );
  OR2_X1 U5149 ( .A1(n5742), .A2(n5165), .ZN(n4172) );
  AOI22_X1 U5150 ( .A1(n5121), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n5107), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4160) );
  AOI22_X1 U5151 ( .A1(n4192), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n5124), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4159) );
  AOI22_X1 U5152 ( .A1(n3468), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4158) );
  AOI22_X1 U5153 ( .A1(n5122), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3089), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4157) );
  NAND4_X1 U5154 ( .A1(n4160), .A2(n4159), .A3(n4158), .A4(n4157), .ZN(n4166)
         );
  AOI22_X1 U5155 ( .A1(n3496), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3486), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4164) );
  AOI22_X1 U5156 ( .A1(n5123), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n5114), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4163) );
  AOI22_X1 U5157 ( .A1(n3462), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n5115), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4162) );
  AOI22_X1 U5158 ( .A1(n3086), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4161) );
  NAND4_X1 U5159 ( .A1(n4164), .A2(n4163), .A3(n4162), .A4(n4161), .ZN(n4165)
         );
  NOR2_X1 U5160 ( .A1(n4166), .A2(n4165), .ZN(n4170) );
  AOI21_X1 U5161 ( .B1(n6966), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4167) );
  AOI21_X1 U5162 ( .B1(n4168), .B2(EAX_REG_20__SCAN_IN), .A(n4167), .ZN(n4169)
         );
  OAI21_X1 U5163 ( .B1(n5177), .B2(n4170), .A(n4169), .ZN(n4171) );
  NAND2_X1 U5164 ( .A1(n4172), .A2(n4171), .ZN(n5379) );
  INV_X1 U5165 ( .A(n5379), .ZN(n4173) );
  AOI22_X1 U5166 ( .A1(n5122), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5107), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4178) );
  AOI22_X1 U5167 ( .A1(n4192), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n5124), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4177) );
  AOI22_X1 U5168 ( .A1(n3496), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3486), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4176) );
  AOI22_X1 U5169 ( .A1(n5123), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4175) );
  NAND4_X1 U5170 ( .A1(n4178), .A2(n4177), .A3(n4176), .A4(n4175), .ZN(n4184)
         );
  AOI22_X1 U5171 ( .A1(n5121), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n5114), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4182) );
  AOI22_X1 U5172 ( .A1(n3468), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n5115), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4181) );
  AOI22_X1 U5173 ( .A1(n3461), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3087), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4180) );
  AOI22_X1 U5174 ( .A1(n3086), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3490), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4179) );
  NAND4_X1 U5175 ( .A1(n4182), .A2(n4181), .A3(n4180), .A4(n4179), .ZN(n4183)
         );
  OR2_X1 U5176 ( .A1(n4184), .A2(n4183), .ZN(n4187) );
  INV_X1 U5177 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4185) );
  INV_X1 U5178 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6953) );
  OAI22_X1 U5179 ( .A1(n3290), .A2(n4185), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6953), .ZN(n4186) );
  AOI21_X1 U5180 ( .B1(n5155), .B2(n4187), .A(n4186), .ZN(n4191) );
  NAND2_X1 U5181 ( .A1(n4189), .A2(n6953), .ZN(n4190) );
  AND2_X1 U5182 ( .A1(n4229), .A2(n4190), .ZN(n5734) );
  MUX2_X1 U5183 ( .A(n4191), .B(n5734), .S(n5182), .Z(n5364) );
  AOI22_X1 U5184 ( .A1(n4192), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n5107), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4196) );
  AOI22_X1 U5185 ( .A1(n5124), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3468), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4195) );
  AOI22_X1 U5186 ( .A1(n3086), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4194) );
  AOI22_X1 U5187 ( .A1(n3496), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5114), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4193) );
  NAND4_X1 U5188 ( .A1(n4196), .A2(n4195), .A3(n4194), .A4(n4193), .ZN(n4202)
         );
  AOI22_X1 U5189 ( .A1(n5122), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3486), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4200) );
  AOI22_X1 U5190 ( .A1(n3461), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n5115), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4199) );
  AOI22_X1 U5191 ( .A1(n5121), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3087), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4198) );
  AOI22_X1 U5192 ( .A1(n5123), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3490), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4197) );
  NAND4_X1 U5193 ( .A1(n4200), .A2(n4199), .A3(n4198), .A4(n4197), .ZN(n4201)
         );
  NOR2_X1 U5194 ( .A1(n4202), .A2(n4201), .ZN(n4204) );
  AOI22_X1 U5195 ( .A1(n4168), .A2(EAX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6673), .ZN(n4203) );
  OAI21_X1 U5196 ( .B1(n5177), .B2(n4204), .A(n4203), .ZN(n4206) );
  INV_X1 U5197 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4205) );
  XNOR2_X1 U5198 ( .A(n4229), .B(n4205), .ZN(n5725) );
  MUX2_X1 U5199 ( .A(n4206), .B(n5725), .S(n5182), .Z(n5351) );
  AOI22_X1 U5200 ( .A1(n5122), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3468), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4210) );
  AOI22_X1 U5201 ( .A1(n3488), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5115), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4209) );
  AOI22_X1 U5202 ( .A1(n5121), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3089), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4208) );
  AOI22_X1 U5203 ( .A1(n3461), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4207) );
  NAND4_X1 U5204 ( .A1(n4210), .A2(n4209), .A3(n4208), .A4(n4207), .ZN(n4216)
         );
  AOI22_X1 U5205 ( .A1(n4192), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n5107), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4214) );
  AOI22_X1 U5206 ( .A1(n5124), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4213) );
  AOI22_X1 U5207 ( .A1(n5123), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4212) );
  AOI22_X1 U5208 ( .A1(n3496), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5114), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4211) );
  NAND4_X1 U5209 ( .A1(n4214), .A2(n4213), .A3(n4212), .A4(n4211), .ZN(n4215)
         );
  NOR2_X1 U5210 ( .A1(n4216), .A2(n4215), .ZN(n5005) );
  AOI22_X1 U5211 ( .A1(n5122), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n5107), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4220) );
  AOI22_X1 U5212 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n4192), .B1(n5121), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4219) );
  AOI22_X1 U5213 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n3467), .B1(n3486), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4218) );
  AOI22_X1 U5214 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n5124), .B1(n3461), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4217) );
  NAND4_X1 U5215 ( .A1(n4220), .A2(n4219), .A3(n4218), .A4(n4217), .ZN(n4226)
         );
  AOI22_X1 U5216 ( .A1(n5123), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n5114), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4224) );
  AOI22_X1 U5217 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n3462), .B1(n5115), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4223) );
  AOI22_X1 U5218 ( .A1(n3496), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3087), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4222) );
  AOI22_X1 U5219 ( .A1(n3086), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4221) );
  NAND4_X1 U5220 ( .A1(n4224), .A2(n4223), .A3(n4222), .A4(n4221), .ZN(n4225)
         );
  NOR2_X1 U5221 ( .A1(n4226), .A2(n4225), .ZN(n5006) );
  XNOR2_X1 U5222 ( .A(n5005), .B(n5006), .ZN(n4228) );
  AOI22_X1 U5223 ( .A1(n4168), .A2(EAX_REG_23__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n6673), .ZN(n4227) );
  OAI21_X1 U5224 ( .B1(n5177), .B2(n4228), .A(n4227), .ZN(n4235) );
  INV_X1 U5225 ( .A(n4229), .ZN(n4230) );
  INV_X1 U5226 ( .A(n4231), .ZN(n4233) );
  INV_X1 U5227 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4232) );
  NAND2_X1 U5228 ( .A1(n4233), .A2(n4232), .ZN(n4234) );
  NAND2_X1 U5229 ( .A1(n5057), .A2(n4234), .ZN(n5346) );
  MUX2_X1 U5230 ( .A(n4235), .B(n5346), .S(n5182), .Z(n4236) );
  OR2_X1 U5231 ( .A1(n5353), .A2(n4236), .ZN(n4237) );
  NAND2_X1 U5232 ( .A1(n5021), .A2(n4237), .ZN(n5628) );
  NAND2_X1 U5233 ( .A1(n4531), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5041) );
  NOR2_X1 U5234 ( .A1(n5041), .A2(n6361), .ZN(n4257) );
  INV_X1 U5235 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6260) );
  NAND2_X1 U5236 ( .A1(n6673), .A2(n6260), .ZN(n6804) );
  NAND2_X1 U5237 ( .A1(n6805), .A2(n6804), .ZN(n4238) );
  NAND2_X1 U5238 ( .A1(n4238), .A2(n4531), .ZN(n4239) );
  INV_X1 U5239 ( .A(n4240), .ZN(n4244) );
  NAND2_X1 U5240 ( .A1(n4531), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4242) );
  NAND2_X1 U5241 ( .A1(n6361), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4241) );
  NAND2_X1 U5242 ( .A1(n4242), .A2(n4241), .ZN(n4345) );
  NOR2_X1 U5243 ( .A1(n5346), .A2(n6599), .ZN(n4243) );
  AOI211_X1 U5244 ( .C1(PHYADDRPOINTER_REG_23__SCAN_IN), .C2(n6591), .A(n4244), 
        .B(n4243), .ZN(n4245) );
  NAND2_X1 U5245 ( .A1(n4248), .A2(n4247), .ZN(U2963) );
  AOI221_X1 U5246 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6800), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n4249) );
  INV_X1 U5247 ( .A(STATE_REG_0__SCAN_IN), .ZN(n4250) );
  AOI221_X1 U5248 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n4249), .C2(HOLD), .A(n4250), .ZN(n4253) );
  INV_X1 U5249 ( .A(NA_N), .ZN(n4251) );
  AOI221_X1 U5250 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n4251), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n4264) );
  AOI22_X1 U5251 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n4270) );
  INV_X1 U5252 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n4265) );
  NOR2_X1 U5253 ( .A1(n4250), .A2(n4265), .ZN(n4255) );
  AND2_X1 U5254 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n4269) );
  AOI21_X1 U5255 ( .B1(n4251), .B2(n4255), .A(n4269), .ZN(n4252) );
  OAI22_X1 U5256 ( .A1(n4253), .A2(n4264), .B1(n4270), .B2(n4252), .ZN(U3183)
         );
  INV_X1 U5257 ( .A(STATE_REG_1__SCAN_IN), .ZN(n4276) );
  AND2_X1 U5258 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n4266) );
  NAND2_X1 U5259 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n4254) );
  OAI21_X1 U5260 ( .B1(n4255), .B2(n4266), .A(n4254), .ZN(n4256) );
  OAI211_X1 U5261 ( .C1(n6800), .C2(n4276), .A(n6798), .B(n4256), .ZN(U3182)
         );
  NOR2_X1 U5262 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6803) );
  INV_X1 U5263 ( .A(n6803), .ZN(n4732) );
  OAI21_X1 U5264 ( .B1(n4531), .B2(READY_N), .A(n6673), .ZN(n4258) );
  AOI21_X1 U5265 ( .B1(n4732), .B2(n4258), .A(n4257), .ZN(n4260) );
  NAND2_X1 U5266 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n6050) );
  INV_X1 U5267 ( .A(n6050), .ZN(n4392) );
  NAND2_X1 U5268 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4392), .ZN(n4741) );
  INV_X1 U5269 ( .A(n4741), .ZN(n4259) );
  NOR2_X1 U5270 ( .A1(n4260), .A2(n4259), .ZN(U3150) );
  INV_X1 U5271 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n4262) );
  NAND2_X1 U5272 ( .A1(n4250), .A2(STATE_REG_1__SCAN_IN), .ZN(n6774) );
  NAND2_X1 U5273 ( .A1(BE_N_REG_3__SCAN_IN), .A2(n6774), .ZN(n4261) );
  OAI21_X1 U5274 ( .B1(n4262), .B2(n6774), .A(n4261), .ZN(U3445) );
  NOR2_X1 U5275 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6360) );
  OAI21_X1 U5276 ( .B1(n6360), .B2(D_C_N_REG_SCAN_IN), .A(n6774), .ZN(n4263)
         );
  OAI21_X1 U5277 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6774), .A(n4263), .ZN(
        U2791) );
  INV_X1 U5278 ( .A(n4264), .ZN(n4268) );
  OAI21_X1 U5279 ( .B1(n4266), .B2(n4265), .A(n6774), .ZN(n4267) );
  OAI211_X1 U5280 ( .C1(n4270), .C2(n4269), .A(n4268), .B(n4267), .ZN(U3181)
         );
  INV_X1 U5281 ( .A(n6774), .ZN(n6751) );
  INV_X1 U5282 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n6991) );
  NAND2_X1 U5283 ( .A1(BYTEENABLE_REG_0__SCAN_IN), .A2(n6751), .ZN(n4271) );
  OAI21_X1 U5284 ( .B1(n6751), .B2(n6991), .A(n4271), .ZN(U3448) );
  NAND2_X1 U5285 ( .A1(n6780), .A2(W_R_N_REG_SCAN_IN), .ZN(n4272) );
  OAI21_X1 U5286 ( .B1(n6780), .B2(READREQUEST_REG_SCAN_IN), .A(n4272), .ZN(
        U3470) );
  INV_X1 U5287 ( .A(STATE_REG_2__SCAN_IN), .ZN(n4273) );
  OR2_X1 U5288 ( .A1(n6774), .A2(n4273), .ZN(n6783) );
  INV_X1 U5289 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6770) );
  INV_X1 U5290 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n6849) );
  INV_X1 U5291 ( .A(REIP_REG_21__SCAN_IN), .ZN(n5732) );
  OR2_X1 U5292 ( .A1(n6774), .A2(STATE_REG_2__SCAN_IN), .ZN(n6778) );
  OAI222_X1 U5293 ( .A1(n6783), .A2(n6770), .B1(n6751), .B2(n6849), .C1(n5732), 
        .C2(n6778), .ZN(U3203) );
  INV_X1 U5294 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n6816) );
  INV_X1 U5295 ( .A(REIP_REG_22__SCAN_IN), .ZN(n5723) );
  OAI222_X1 U5296 ( .A1(n6783), .A2(n5732), .B1(n6751), .B2(n6816), .C1(n5723), 
        .C2(n6778), .ZN(U3204) );
  INV_X1 U5297 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n6829) );
  INV_X1 U5298 ( .A(REIP_REG_23__SCAN_IN), .ZN(n4274) );
  OAI222_X1 U5299 ( .A1(n6783), .A2(n5723), .B1(n6751), .B2(n6829), .C1(n6778), 
        .C2(n4274), .ZN(U3205) );
  INV_X1 U5300 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6952) );
  INV_X1 U5301 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n6874) );
  INV_X1 U5302 ( .A(REIP_REG_30__SCAN_IN), .ZN(n5259) );
  OAI222_X1 U5303 ( .A1(n6783), .A2(n6952), .B1(n6751), .B2(n6874), .C1(n5259), 
        .C2(n6778), .ZN(U3212) );
  INV_X1 U5304 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n6995) );
  INV_X1 U5305 ( .A(REIP_REG_31__SCAN_IN), .ZN(n4275) );
  OAI222_X1 U5306 ( .A1(n6783), .A2(n5259), .B1(n6751), .B2(n6995), .C1(n4275), 
        .C2(n6778), .ZN(U3213) );
  INV_X1 U5307 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6748) );
  INV_X1 U5308 ( .A(REIP_REG_3__SCAN_IN), .ZN(n7085) );
  INV_X1 U5309 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n6830) );
  OAI222_X1 U5310 ( .A1(n6778), .A2(n6748), .B1(n6783), .B2(n7085), .C1(n6830), 
        .C2(n6751), .ZN(U3186) );
  INV_X1 U5311 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6609) );
  INV_X1 U5312 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6753) );
  INV_X1 U5313 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n6876) );
  OAI222_X1 U5314 ( .A1(n6778), .A2(n6609), .B1(n6783), .B2(n6753), .C1(n6751), 
        .C2(n6876), .ZN(U3190) );
  INV_X1 U5315 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6784) );
  INV_X1 U5316 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n7104) );
  INV_X1 U5317 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6779) );
  OAI222_X1 U5318 ( .A1(n6778), .A2(n6784), .B1(n6751), .B2(n7104), .C1(n6779), 
        .C2(n6783), .ZN(U3210) );
  INV_X1 U5319 ( .A(ADS_N_REG_SCAN_IN), .ZN(n4278) );
  OAI21_X1 U5320 ( .B1(n4276), .B2(STATE_REG_2__SCAN_IN), .A(
        STATE_REG_0__SCAN_IN), .ZN(n4277) );
  AND2_X1 U5321 ( .A1(n4277), .A2(n6774), .ZN(n6788) );
  INV_X1 U5322 ( .A(n6788), .ZN(n6786) );
  OAI21_X1 U5323 ( .B1(n6751), .B2(n4278), .A(n6786), .ZN(U2789) );
  NOR2_X1 U5324 ( .A1(n6804), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5400) );
  INV_X1 U5325 ( .A(n5400), .ZN(n4285) );
  OR2_X1 U5326 ( .A1(n4376), .A2(n4279), .ZN(n4283) );
  INV_X1 U5327 ( .A(n4293), .ZN(n4280) );
  NAND2_X1 U5328 ( .A1(n3752), .A2(n4280), .ZN(n4286) );
  INV_X1 U5329 ( .A(n4281), .ZN(n4290) );
  NAND2_X1 U5330 ( .A1(n4286), .A2(n4290), .ZN(n4282) );
  NAND2_X1 U5331 ( .A1(n4283), .A2(n4282), .ZN(n4289) );
  INV_X1 U5332 ( .A(n4737), .ZN(n6736) );
  OAI21_X1 U5333 ( .B1(n4289), .B2(n6736), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n4284) );
  OAI21_X1 U5334 ( .B1(n4285), .B2(n4531), .A(n4284), .ZN(U2790) );
  AOI21_X1 U5335 ( .B1(n5039), .B2(MEMORYFETCH_REG_SCAN_IN), .A(n5400), .ZN(
        n4287) );
  NAND2_X1 U5336 ( .A1(n5040), .A2(n4287), .ZN(U2788) );
  INV_X1 U5337 ( .A(MORE_REG_SCAN_IN), .ZN(n6897) );
  AND2_X1 U5338 ( .A1(n5515), .A2(n3764), .ZN(n6797) );
  AOI21_X1 U5339 ( .B1(n6797), .B2(n6798), .A(READY_N), .ZN(n4288) );
  OR2_X1 U5340 ( .A1(n4289), .A2(n4288), .ZN(n4518) );
  AND2_X1 U5341 ( .A1(n4518), .A2(n4737), .ZN(n6363) );
  AND2_X1 U5342 ( .A1(n4291), .A2(n4290), .ZN(n4292) );
  MUX2_X1 U5343 ( .A(n4292), .B(n4473), .S(n4376), .Z(n4295) );
  NAND2_X1 U5344 ( .A1(n3752), .A2(n4293), .ZN(n4294) );
  AND2_X1 U5345 ( .A1(n4295), .A2(n4294), .ZN(n4517) );
  INV_X1 U5346 ( .A(n4517), .ZN(n4296) );
  NAND2_X1 U5347 ( .A1(n4296), .A2(n6363), .ZN(n4297) );
  OAI21_X1 U5348 ( .B1(n6897), .B2(n6363), .A(n4297), .ZN(U3471) );
  NAND2_X1 U5349 ( .A1(n4498), .A2(n4472), .ZN(n4299) );
  OAI21_X1 U5350 ( .B1(n4472), .B2(n4991), .A(n3739), .ZN(n4298) );
  NAND2_X1 U5351 ( .A1(n4299), .A2(n4298), .ZN(n4300) );
  NAND2_X1 U5352 ( .A1(n4300), .A2(n6800), .ZN(n4301) );
  NAND2_X1 U5353 ( .A1(n4301), .A2(n4714), .ZN(n4306) );
  INV_X1 U5354 ( .A(n4716), .ZN(n4302) );
  NOR2_X1 U5355 ( .A1(n4721), .A2(n4302), .ZN(n4303) );
  OR2_X1 U5356 ( .A1(n4304), .A2(n4303), .ZN(n4305) );
  AOI21_X1 U5357 ( .B1(n4376), .B2(n4306), .A(n4305), .ZN(n4308) );
  NAND2_X1 U5358 ( .A1(n4308), .A2(n4307), .ZN(n4511) );
  INV_X1 U5359 ( .A(FLUSH_REG_SCAN_IN), .ZN(n4525) );
  NOR2_X1 U5360 ( .A1(n4525), .A2(n4741), .ZN(n4309) );
  AOI21_X1 U5361 ( .B1(n4511), .B2(n4737), .A(n4309), .ZN(n4326) );
  OAI21_X1 U5362 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n6260), .A(n4326), .ZN(
        n6065) );
  OAI21_X1 U5363 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6061), .A(n6065), 
        .ZN(n4332) );
  INV_X1 U5364 ( .A(n4332), .ZN(n4322) );
  NAND2_X1 U5365 ( .A1(n4719), .A2(n3859), .ZN(n4311) );
  NOR2_X1 U5366 ( .A1(n3739), .A2(n4311), .ZN(n4312) );
  NAND3_X1 U5367 ( .A1(n4313), .A2(n4312), .A3(n4721), .ZN(n4490) );
  NAND2_X1 U5368 ( .A1(n4310), .A2(n4490), .ZN(n4318) );
  NOR2_X1 U5369 ( .A1(n4314), .A2(n4943), .ZN(n4316) );
  AOI22_X1 U5370 ( .A1(n4498), .A2(n4474), .B1(n4316), .B2(n4328), .ZN(n4317)
         );
  NAND2_X1 U5371 ( .A1(n4318), .A2(n4317), .ZN(n4484) );
  NAND2_X1 U5372 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        STATE2_REG_1__SCAN_IN), .ZN(n4944) );
  INV_X1 U5373 ( .A(n4944), .ZN(n4320) );
  INV_X1 U5374 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5240) );
  AOI22_X1 U5375 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5240), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4592), .ZN(n4945) );
  INV_X1 U5376 ( .A(n6061), .ZN(n4942) );
  AOI222_X1 U5377 ( .A1(n4484), .A2(n4948), .B1(n4320), .B2(n4945), .C1(n4319), 
        .C2(n4942), .ZN(n4321) );
  INV_X1 U5378 ( .A(n6065), .ZN(n4951) );
  OAI22_X1 U5379 ( .A1(n4322), .A2(n4474), .B1(n4321), .B2(n4951), .ZN(U3460)
         );
  INV_X1 U5380 ( .A(n4780), .ZN(n4323) );
  NOR2_X1 U5381 ( .A1(n4324), .A2(n4323), .ZN(n4325) );
  XNOR2_X1 U5382 ( .A(n4325), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5526)
         );
  INV_X1 U5383 ( .A(n4948), .ZN(n6063) );
  OR4_X1 U5384 ( .A1(n5526), .A2(n4326), .A3(n4721), .A4(n6063), .ZN(n4327) );
  OAI21_X1 U5385 ( .B1(n6065), .B2(n4512), .A(n4327), .ZN(U3455) );
  NAND2_X1 U5386 ( .A1(n4498), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4481) );
  INV_X1 U5387 ( .A(n4490), .ZN(n4480) );
  OR2_X1 U5388 ( .A1(n3915), .A2(n4480), .ZN(n4330) );
  AND2_X1 U5389 ( .A1(n4330), .A2(n4329), .ZN(n4483) );
  OAI22_X1 U5390 ( .A1(n4483), .A2(n6063), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n4513), .ZN(n4331) );
  OAI22_X1 U5391 ( .A1(n4332), .A2(n4331), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6065), .ZN(n4333) );
  OAI21_X1 U5392 ( .B1(n4481), .B2(n6063), .A(n4333), .ZN(U3461) );
  INV_X1 U5393 ( .A(DATAI_15_), .ZN(n4337) );
  NOR2_X1 U5394 ( .A1(n5197), .A2(n6800), .ZN(n4335) );
  INV_X1 U5395 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n6818) );
  INV_X1 U5396 ( .A(EAX_REG_15__SCAN_IN), .ZN(n4336) );
  OAI222_X1 U5397 ( .A1(n4337), .A2(n6556), .B1(n6523), .B2(n6818), .C1(n4336), 
        .C2(n6561), .ZN(U2954) );
  INV_X1 U5398 ( .A(UWORD_REG_14__SCAN_IN), .ZN(n7012) );
  INV_X2 U5399 ( .A(n6561), .ZN(n6553) );
  NAND2_X1 U5400 ( .A1(n6553), .A2(EAX_REG_30__SCAN_IN), .ZN(n4339) );
  INV_X1 U5401 ( .A(DATAI_14_), .ZN(n4338) );
  OR2_X1 U5402 ( .A1(n6556), .A2(n4338), .ZN(n6559) );
  OAI211_X1 U5403 ( .C1(n6523), .C2(n7012), .A(n4339), .B(n6559), .ZN(U2938)
         );
  XNOR2_X1 U5404 ( .A(n4340), .B(n6838), .ZN(n4358) );
  INV_X1 U5405 ( .A(n4358), .ZN(n4351) );
  NAND2_X1 U5406 ( .A1(n4342), .A2(n4341), .ZN(n4343) );
  NAND2_X1 U5407 ( .A1(n4344), .A2(n4343), .ZN(n5560) );
  INV_X1 U5408 ( .A(n5560), .ZN(n4349) );
  INV_X1 U5409 ( .A(REIP_REG_0__SCAN_IN), .ZN(n7076) );
  NOR2_X1 U5410 ( .A1(n6639), .A2(n7076), .ZN(n4357) );
  INV_X1 U5411 ( .A(n4345), .ZN(n4347) );
  INV_X1 U5412 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n4346) );
  AOI21_X1 U5413 ( .B1(n5853), .B2(n4347), .A(n4346), .ZN(n4348) );
  AOI211_X1 U5414 ( .C1(n4349), .C2(n6594), .A(n4357), .B(n4348), .ZN(n4350)
         );
  OAI21_X1 U5415 ( .B1(n4351), .B2(n6362), .A(n4350), .ZN(U2986) );
  INV_X1 U5416 ( .A(n4352), .ZN(n5985) );
  NOR2_X1 U5417 ( .A1(n5985), .A2(n6636), .ZN(n5991) );
  OR2_X1 U5418 ( .A1(n4993), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4354)
         );
  AND2_X1 U5419 ( .A1(n4354), .A2(n4353), .ZN(n5553) );
  AOI21_X1 U5420 ( .B1(n6004), .B2(n4355), .A(n6838), .ZN(n4356) );
  AOI211_X1 U5421 ( .C1(n5553), .C2(n6651), .A(n4357), .B(n4356), .ZN(n4360)
         );
  NAND2_X1 U5422 ( .A1(n4358), .A2(n6653), .ZN(n4359) );
  OAI211_X1 U5423 ( .C1(INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n5991), .A(n4360), 
        .B(n4359), .ZN(U3018) );
  INV_X1 U5424 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4365) );
  INV_X1 U5425 ( .A(n4498), .ZN(n4361) );
  OR2_X1 U5426 ( .A1(n4715), .A2(n4361), .ZN(n4362) );
  NAND2_X1 U5427 ( .A1(n6561), .A2(n4362), .ZN(n4363) );
  NAND2_X1 U5428 ( .A1(n6814), .A2(n5200), .ZN(n6481) );
  NOR2_X2 U5429 ( .A1(n6050), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6813) );
  NOR2_X4 U5430 ( .A1(n6814), .A2(n6813), .ZN(n6812) );
  AOI22_X1 U5431 ( .A1(n6813), .A2(UWORD_REG_4__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4364) );
  OAI21_X1 U5432 ( .B1(n4365), .B2(n6481), .A(n4364), .ZN(U2903) );
  INV_X1 U5433 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4367) );
  AOI22_X1 U5434 ( .A1(n6813), .A2(UWORD_REG_12__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4366) );
  OAI21_X1 U5435 ( .B1(n4367), .B2(n6481), .A(n4366), .ZN(U2895) );
  AOI22_X1 U5436 ( .A1(n6813), .A2(UWORD_REG_1__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4368) );
  OAI21_X1 U5437 ( .B1(n4004), .B2(n6481), .A(n4368), .ZN(U2906) );
  INV_X1 U5438 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4370) );
  AOI22_X1 U5439 ( .A1(n6813), .A2(UWORD_REG_3__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4369) );
  OAI21_X1 U5440 ( .B1(n4370), .B2(n6481), .A(n4369), .ZN(U2904) );
  AOI22_X1 U5441 ( .A1(n6813), .A2(UWORD_REG_5__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4371) );
  OAI21_X1 U5442 ( .B1(n4185), .B2(n6481), .A(n4371), .ZN(U2902) );
  INV_X1 U5443 ( .A(EAX_REG_23__SCAN_IN), .ZN(n6833) );
  AOI22_X1 U5444 ( .A1(n6813), .A2(UWORD_REG_7__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4372) );
  OAI21_X1 U5445 ( .B1(n6833), .B2(n6481), .A(n4372), .ZN(U2900) );
  OR2_X1 U5446 ( .A1(n4373), .A2(n3764), .ZN(n4374) );
  OAI22_X1 U5447 ( .A1(n4376), .A2(n4473), .B1(n4375), .B2(n4374), .ZN(n4377)
         );
  NAND2_X1 U5448 ( .A1(n6480), .A2(n3400), .ZN(n5599) );
  OAI21_X1 U5449 ( .B1(n4380), .B2(n4379), .A(n4378), .ZN(n5551) );
  INV_X1 U5450 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4384) );
  OAI21_X1 U5451 ( .B1(n4382), .B2(n4991), .A(n4381), .ZN(n5544) );
  INV_X1 U5452 ( .A(n5544), .ZN(n4383) );
  OAI222_X1 U5453 ( .A1(n5599), .A2(n5551), .B1(n6480), .B2(n4384), .C1(n5605), 
        .C2(n4383), .ZN(U2858) );
  INV_X1 U5454 ( .A(n5553), .ZN(n4386) );
  INV_X1 U5455 ( .A(n5599), .ZN(n6478) );
  OAI222_X1 U5456 ( .A1(n4386), .A2(n5605), .B1(n4385), .B2(n6480), .C1(n5560), 
        .C2(n6471), .ZN(U2859) );
  AND2_X1 U5457 ( .A1(n3091), .A2(n3912), .ZN(n6354) );
  NAND2_X1 U5458 ( .A1(n6594), .A2(DATAI_29_), .ZN(n6714) );
  OR2_X1 U5459 ( .A1(n6804), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6108) );
  OAI21_X1 U5460 ( .B1(n3091), .B2(n5858), .A(n6108), .ZN(n4391) );
  INV_X1 U5461 ( .A(n6455), .ZN(n4388) );
  NAND2_X1 U5462 ( .A1(n4388), .A2(n4310), .ZN(n6311) );
  INV_X1 U5463 ( .A(n6311), .ZN(n4390) );
  INV_X1 U5464 ( .A(n3915), .ZN(n6667) );
  AND2_X1 U5465 ( .A1(n4491), .A2(n6667), .ZN(n6159) );
  INV_X1 U5466 ( .A(n4425), .ZN(n4389) );
  AOI21_X1 U5467 ( .B1(n4390), .B2(n6159), .A(n4389), .ZN(n4397) );
  NAND2_X1 U5468 ( .A1(n4391), .A2(n4397), .ZN(n4396) );
  OR2_X1 U5469 ( .A1(n6803), .A2(n4392), .ZN(n4393) );
  NAND2_X1 U5470 ( .A1(n6304), .A2(STATE2_REG_3__SCAN_IN), .ZN(n4395) );
  NAND2_X1 U5471 ( .A1(n4673), .A2(n4395), .ZN(n6164) );
  INV_X1 U5472 ( .A(n6164), .ZN(n4618) );
  OAI211_X1 U5473 ( .C1(n6305), .C2(n6663), .A(n4396), .B(n4618), .ZN(n4423)
         );
  NAND2_X1 U5474 ( .A1(n4423), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4401)
         );
  NAND2_X1 U5475 ( .A1(n3091), .A2(n6071), .ZN(n4707) );
  AND2_X1 U5476 ( .A1(n5839), .A2(DATAI_21_), .ZN(n6342) );
  INV_X1 U5477 ( .A(n4397), .ZN(n4398) );
  AOI22_X1 U5478 ( .A1(n4398), .A2(n6663), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6305), .ZN(n4426) );
  AND2_X1 U5479 ( .A1(n4673), .A2(DATAI_5_), .ZN(n6711) );
  OR2_X1 U5480 ( .A1(n4424), .A2(n3387), .ZN(n6708) );
  OAI22_X1 U5481 ( .A1(n4426), .A2(n6340), .B1(n4425), .B2(n6708), .ZN(n4399)
         );
  AOI21_X1 U5482 ( .B1(n4428), .B2(n6342), .A(n4399), .ZN(n4400) );
  OAI211_X1 U5483 ( .C1(n4431), .C2(n6714), .A(n4401), .B(n4400), .ZN(U3145)
         );
  NAND2_X1 U5484 ( .A1(n6594), .A2(DATAI_30_), .ZN(n6721) );
  NAND2_X1 U5485 ( .A1(n4423), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4405)
         );
  AND2_X1 U5486 ( .A1(n5839), .A2(DATAI_22_), .ZN(n6347) );
  AND2_X1 U5487 ( .A1(n4673), .A2(DATAI_6_), .ZN(n6718) );
  OR2_X1 U5488 ( .A1(n4424), .A2(n4402), .ZN(n6715) );
  OAI22_X1 U5489 ( .A1(n4426), .A2(n6345), .B1(n4425), .B2(n6715), .ZN(n4403)
         );
  AOI21_X1 U5490 ( .B1(n4428), .B2(n6347), .A(n4403), .ZN(n4404) );
  OAI211_X1 U5491 ( .C1(n4431), .C2(n6721), .A(n4405), .B(n4404), .ZN(U3146)
         );
  NAND2_X1 U5492 ( .A1(n6594), .A2(DATAI_27_), .ZN(n6695) );
  NAND2_X1 U5493 ( .A1(n4423), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4409)
         );
  NAND2_X1 U5494 ( .A1(n6594), .A2(DATAI_19_), .ZN(n6700) );
  INV_X1 U5495 ( .A(n6700), .ZN(n6332) );
  AND2_X1 U5496 ( .A1(n4673), .A2(DATAI_3_), .ZN(n6697) );
  OR2_X1 U5497 ( .A1(n4424), .A2(n4406), .ZN(n6694) );
  OAI22_X1 U5498 ( .A1(n4426), .A2(n6330), .B1(n4425), .B2(n6694), .ZN(n4407)
         );
  AOI21_X1 U5499 ( .B1(n4428), .B2(n6332), .A(n4407), .ZN(n4408) );
  OAI211_X1 U5500 ( .C1(n4431), .C2(n6695), .A(n4409), .B(n4408), .ZN(U3143)
         );
  NAND2_X1 U5501 ( .A1(n6594), .A2(DATAI_28_), .ZN(n6707) );
  NAND2_X1 U5502 ( .A1(n4423), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4412)
         );
  AND2_X1 U5503 ( .A1(n5839), .A2(DATAI_20_), .ZN(n6337) );
  AND2_X1 U5504 ( .A1(n4673), .A2(DATAI_4_), .ZN(n6704) );
  OR2_X1 U5505 ( .A1(n4424), .A2(n4717), .ZN(n6701) );
  OAI22_X1 U5506 ( .A1(n4426), .A2(n6335), .B1(n4425), .B2(n6701), .ZN(n4410)
         );
  AOI21_X1 U5507 ( .B1(n4428), .B2(n6337), .A(n4410), .ZN(n4411) );
  OAI211_X1 U5508 ( .C1(n4431), .C2(n6707), .A(n4412), .B(n4411), .ZN(U3144)
         );
  NAND2_X1 U5509 ( .A1(n6594), .A2(DATAI_25_), .ZN(n6681) );
  NAND2_X1 U5510 ( .A1(n4423), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4416)
         );
  NAND2_X1 U5511 ( .A1(n5839), .A2(DATAI_17_), .ZN(n6686) );
  INV_X1 U5512 ( .A(n6686), .ZN(n6322) );
  AND2_X1 U5513 ( .A1(n4673), .A2(DATAI_1_), .ZN(n6683) );
  OR2_X1 U5514 ( .A1(n4424), .A2(n4413), .ZN(n6680) );
  OAI22_X1 U5515 ( .A1(n4426), .A2(n6320), .B1(n4425), .B2(n6680), .ZN(n4414)
         );
  AOI21_X1 U5516 ( .B1(n4428), .B2(n6322), .A(n4414), .ZN(n4415) );
  OAI211_X1 U5517 ( .C1(n4431), .C2(n6681), .A(n4416), .B(n4415), .ZN(U3141)
         );
  NAND2_X1 U5518 ( .A1(n6594), .A2(DATAI_26_), .ZN(n6693) );
  NAND2_X1 U5519 ( .A1(n4423), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4419)
         );
  AND2_X1 U5520 ( .A1(n5839), .A2(DATAI_18_), .ZN(n6327) );
  AND2_X1 U5521 ( .A1(n4673), .A2(DATAI_2_), .ZN(n6690) );
  OAI22_X1 U5522 ( .A1(n4426), .A2(n6325), .B1(n4425), .B2(n6687), .ZN(n4417)
         );
  AOI21_X1 U5523 ( .B1(n4428), .B2(n6327), .A(n4417), .ZN(n4418) );
  OAI211_X1 U5524 ( .C1(n4431), .C2(n6693), .A(n4419), .B(n4418), .ZN(U3142)
         );
  NAND2_X1 U5525 ( .A1(n6594), .A2(DATAI_31_), .ZN(n6733) );
  NAND2_X1 U5526 ( .A1(n4423), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4422)
         );
  AND2_X1 U5527 ( .A1(n5839), .A2(DATAI_23_), .ZN(n6355) );
  AND2_X1 U5528 ( .A1(n4673), .A2(DATAI_7_), .ZN(n6728) );
  OAI22_X1 U5529 ( .A1(n4426), .A2(n6351), .B1(n4425), .B2(n6723), .ZN(n4420)
         );
  AOI21_X1 U5530 ( .B1(n4428), .B2(n6355), .A(n4420), .ZN(n4421) );
  OAI211_X1 U5531 ( .C1(n4431), .C2(n6733), .A(n4422), .B(n4421), .ZN(U3147)
         );
  NAND2_X1 U5532 ( .A1(n5839), .A2(DATAI_24_), .ZN(n6679) );
  NAND2_X1 U5533 ( .A1(n4423), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4430)
         );
  AND2_X1 U5534 ( .A1(n5839), .A2(DATAI_16_), .ZN(n6308) );
  AND2_X1 U5535 ( .A1(n4673), .A2(DATAI_0_), .ZN(n6676) );
  OAI22_X1 U5536 ( .A1(n4426), .A2(n6306), .B1(n4425), .B2(n6660), .ZN(n4427)
         );
  AOI21_X1 U5537 ( .B1(n4428), .B2(n6308), .A(n4427), .ZN(n4429) );
  OAI211_X1 U5538 ( .C1(n4431), .C2(n6679), .A(n4430), .B(n4429), .ZN(U3140)
         );
  INV_X1 U5539 ( .A(n6347), .ZN(n6716) );
  NAND2_X1 U5540 ( .A1(n6203), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6664) );
  INV_X1 U5541 ( .A(n6664), .ZN(n4539) );
  NAND2_X1 U5542 ( .A1(n3119), .A2(n4539), .ZN(n4582) );
  NOR2_X1 U5543 ( .A1(n4582), .A2(n6804), .ZN(n4432) );
  NAND2_X1 U5544 ( .A1(n4455), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4436) );
  INV_X1 U5545 ( .A(n6721), .ZN(n4906) );
  OR2_X1 U5546 ( .A1(n6206), .A2(n6311), .ZN(n4610) );
  OAI21_X1 U5547 ( .B1(n4610), .B2(n3915), .A(n4456), .ZN(n4433) );
  AOI22_X1 U5548 ( .A1(n4433), .A2(n6663), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4605), .ZN(n4457) );
  OAI22_X1 U5549 ( .A1(n4457), .A2(n6345), .B1(n4456), .B2(n6715), .ZN(n4434)
         );
  AOI21_X1 U5550 ( .B1(n6151), .B2(n4906), .A(n4434), .ZN(n4435) );
  OAI211_X1 U5551 ( .C1(n4461), .C2(n6716), .A(n4436), .B(n4435), .ZN(U3082)
         );
  INV_X1 U5552 ( .A(n6327), .ZN(n6688) );
  NAND2_X1 U5553 ( .A1(n4455), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4439) );
  INV_X1 U5554 ( .A(n6693), .ZN(n4914) );
  OAI22_X1 U5555 ( .A1(n4457), .A2(n6325), .B1(n4456), .B2(n6687), .ZN(n4437)
         );
  AOI21_X1 U5556 ( .B1(n6151), .B2(n4914), .A(n4437), .ZN(n4438) );
  OAI211_X1 U5557 ( .C1(n4461), .C2(n6688), .A(n4439), .B(n4438), .ZN(U3078)
         );
  INV_X1 U5558 ( .A(n6342), .ZN(n6709) );
  NAND2_X1 U5559 ( .A1(n4455), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4442) );
  INV_X1 U5560 ( .A(n6714), .ZN(n4922) );
  OAI22_X1 U5561 ( .A1(n4457), .A2(n6340), .B1(n4456), .B2(n6708), .ZN(n4440)
         );
  AOI21_X1 U5562 ( .B1(n6151), .B2(n4922), .A(n4440), .ZN(n4441) );
  OAI211_X1 U5563 ( .C1(n4461), .C2(n6709), .A(n4442), .B(n4441), .ZN(U3081)
         );
  NAND2_X1 U5564 ( .A1(n4455), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4445) );
  INV_X1 U5565 ( .A(n6695), .ZN(n4918) );
  OAI22_X1 U5566 ( .A1(n4457), .A2(n6330), .B1(n4456), .B2(n6694), .ZN(n4443)
         );
  AOI21_X1 U5567 ( .B1(n6151), .B2(n4918), .A(n4443), .ZN(n4444) );
  OAI211_X1 U5568 ( .C1(n4461), .C2(n6700), .A(n4445), .B(n4444), .ZN(U3079)
         );
  INV_X1 U5569 ( .A(n6355), .ZN(n6724) );
  NAND2_X1 U5570 ( .A1(n4455), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4448) );
  INV_X1 U5571 ( .A(n6733), .ZN(n4910) );
  OAI22_X1 U5572 ( .A1(n4457), .A2(n6351), .B1(n4456), .B2(n6723), .ZN(n4446)
         );
  AOI21_X1 U5573 ( .B1(n6151), .B2(n4910), .A(n4446), .ZN(n4447) );
  OAI211_X1 U5574 ( .C1(n4461), .C2(n6724), .A(n4448), .B(n4447), .ZN(U3083)
         );
  INV_X1 U5575 ( .A(n6308), .ZN(n6661) );
  NAND2_X1 U5576 ( .A1(n4455), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4451) );
  INV_X1 U5577 ( .A(n6679), .ZN(n6149) );
  OAI22_X1 U5578 ( .A1(n4457), .A2(n6306), .B1(n4456), .B2(n6660), .ZN(n4449)
         );
  AOI21_X1 U5579 ( .B1(n6151), .B2(n6149), .A(n4449), .ZN(n4450) );
  OAI211_X1 U5580 ( .C1(n4461), .C2(n6661), .A(n4451), .B(n4450), .ZN(U3076)
         );
  NAND2_X1 U5581 ( .A1(n4455), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4454) );
  INV_X1 U5582 ( .A(n6681), .ZN(n4929) );
  OAI22_X1 U5583 ( .A1(n4457), .A2(n6320), .B1(n4456), .B2(n6680), .ZN(n4452)
         );
  AOI21_X1 U5584 ( .B1(n6151), .B2(n4929), .A(n4452), .ZN(n4453) );
  OAI211_X1 U5585 ( .C1(n4461), .C2(n6686), .A(n4454), .B(n4453), .ZN(U3077)
         );
  INV_X1 U5586 ( .A(n6337), .ZN(n6702) );
  NAND2_X1 U5587 ( .A1(n4455), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4460) );
  INV_X1 U5588 ( .A(n6707), .ZN(n4936) );
  OAI22_X1 U5589 ( .A1(n4457), .A2(n6335), .B1(n4456), .B2(n6701), .ZN(n4458)
         );
  AOI21_X1 U5590 ( .B1(n6151), .B2(n4936), .A(n4458), .ZN(n4459) );
  OAI211_X1 U5591 ( .C1(n4461), .C2(n6702), .A(n4460), .B(n4459), .ZN(U3080)
         );
  NOR2_X1 U5592 ( .A1(n4464), .A2(n4463), .ZN(n4465) );
  NOR2_X1 U5593 ( .A1(n4462), .A2(n4465), .ZN(n6595) );
  INV_X1 U5594 ( .A(n6595), .ZN(n4882) );
  AND2_X1 U5595 ( .A1(n4467), .A2(n4466), .ZN(n4469) );
  OR2_X1 U5596 ( .A1(n4469), .A2(n4468), .ZN(n4591) );
  INV_X1 U5597 ( .A(n4591), .ZN(n6450) );
  INV_X1 U5598 ( .A(n6480), .ZN(n5597) );
  AOI22_X1 U5599 ( .A1(n6477), .A2(n6450), .B1(EBX_REG_2__SCAN_IN), .B2(n5597), 
        .ZN(n4470) );
  OAI21_X1 U5600 ( .B1(n4882), .B2(n6471), .A(n4470), .ZN(U2857) );
  NAND2_X1 U5601 ( .A1(n6800), .A2(n6361), .ZN(n5198) );
  INV_X1 U5602 ( .A(n5198), .ZN(n4471) );
  NAND2_X1 U5603 ( .A1(n4472), .A2(n4471), .ZN(n5196) );
  NAND2_X1 U5604 ( .A1(n4473), .A2(n4714), .ZN(n4503) );
  XNOR2_X1 U5605 ( .A(n4943), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4478)
         );
  XNOR2_X1 U5606 ( .A(n4474), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4475)
         );
  NAND2_X1 U5607 ( .A1(n4498), .A2(n4475), .ZN(n4476) );
  OAI21_X1 U5608 ( .B1(n4478), .B2(n4500), .A(n4476), .ZN(n4477) );
  AOI21_X1 U5609 ( .B1(n4503), .B2(n4478), .A(n4477), .ZN(n4479) );
  OAI21_X1 U5610 ( .B1(n6455), .B2(n4480), .A(n4479), .ZN(n4949) );
  MUX2_X1 U5611 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n4949), .S(n4511), 
        .Z(n4523) );
  AND2_X1 U5612 ( .A1(n4481), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4482)
         );
  NAND2_X1 U5613 ( .A1(n4483), .A2(n4482), .ZN(n4485) );
  INV_X1 U5614 ( .A(n4485), .ZN(n4487) );
  OAI211_X1 U5615 ( .C1(n4485), .C2(n4839), .A(n4511), .B(n4484), .ZN(n4486)
         );
  OAI21_X1 U5616 ( .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n4487), .A(n4486), 
        .ZN(n4488) );
  AOI21_X1 U5617 ( .B1(n4523), .B2(n4489), .A(n4488), .ZN(n4507) );
  NOR2_X1 U5618 ( .A1(n4523), .A2(n4489), .ZN(n4506) );
  NAND2_X1 U5619 ( .A1(n4491), .A2(n4490), .ZN(n4505) );
  MUX2_X1 U5620 ( .A(n4492), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4943), 
        .Z(n4493) );
  AOI21_X1 U5621 ( .B1(n4943), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n4495), 
        .ZN(n4494) );
  NOR2_X1 U5622 ( .A1(n3086), .A2(n4494), .ZN(n6062) );
  XNOR2_X1 U5623 ( .A(n4496), .B(n4495), .ZN(n4497) );
  NAND2_X1 U5624 ( .A1(n4498), .A2(n4497), .ZN(n4499) );
  OAI21_X1 U5625 ( .B1(n6062), .B2(n4500), .A(n4499), .ZN(n4501) );
  AOI21_X1 U5626 ( .B1(n4503), .B2(n4502), .A(n4501), .ZN(n4504) );
  NAND2_X1 U5627 ( .A1(n4505), .A2(n4504), .ZN(n6060) );
  MUX2_X1 U5628 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6060), .S(n4511), 
        .Z(n4524) );
  INV_X1 U5629 ( .A(n4524), .ZN(n4508) );
  OAI22_X1 U5630 ( .A1(n4507), .A2(n4506), .B1(n4508), .B2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4510) );
  NAND2_X1 U5631 ( .A1(n4508), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4509) );
  NAND3_X1 U5632 ( .A1(n4510), .A2(n6659), .A3(n4509), .ZN(n4522) );
  NOR2_X1 U5633 ( .A1(n4512), .A2(FLUSH_REG_SCAN_IN), .ZN(n4515) );
  OAI22_X1 U5634 ( .A1(n5526), .A2(n4721), .B1(n4512), .B2(n4511), .ZN(n4514)
         );
  MUX2_X1 U5635 ( .A(n4515), .B(n4514), .S(n4513), .Z(n4576) );
  NOR2_X1 U5636 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n4519) );
  OAI211_X1 U5637 ( .C1(n4519), .C2(n4518), .A(n4517), .B(n4516), .ZN(n4520)
         );
  NOR2_X1 U5638 ( .A1(n4576), .A2(n4520), .ZN(n4521) );
  AND2_X1 U5639 ( .A1(n4522), .A2(n4521), .ZN(n4528) );
  NAND2_X1 U5640 ( .A1(n4524), .A2(n4523), .ZN(n4527) );
  MUX2_X1 U5641 ( .A(n4527), .B(n4526), .S(STATE2_REG_1__SCAN_IN), .Z(n4578)
         );
  NAND2_X1 U5642 ( .A1(n4528), .A2(n4578), .ZN(n4738) );
  INV_X1 U5643 ( .A(n6813), .ZN(n6806) );
  OAI22_X1 U5644 ( .A1(n4738), .A2(n6736), .B1(n6800), .B2(n6806), .ZN(n4529)
         );
  OAI21_X1 U5645 ( .B1(n5196), .B2(n4530), .A(n4529), .ZN(n6741) );
  INV_X1 U5646 ( .A(n6741), .ZN(n4733) );
  OAI21_X1 U5647 ( .B1(n4733), .B2(n4531), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n4532) );
  NAND2_X1 U5648 ( .A1(n4532), .A2(n4741), .ZN(U3453) );
  NAND2_X1 U5649 ( .A1(n4462), .A2(n4883), .ZN(n4535) );
  INV_X1 U5650 ( .A(n4533), .ZN(n4534) );
  NAND2_X1 U5651 ( .A1(n4535), .A2(n4534), .ZN(n4536) );
  NAND2_X1 U5652 ( .A1(n4536), .A2(n4769), .ZN(n5532) );
  INV_X1 U5653 ( .A(EBX_REG_4__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U5654 ( .A1(n5536), .A2(n4537), .ZN(n4538) );
  NAND2_X1 U5655 ( .A1(n4666), .A2(n4538), .ZN(n6641) );
  OAI222_X1 U5656 ( .A1(n5532), .A2(n6471), .B1(n6480), .B2(n5520), .C1(n6641), 
        .C2(n5605), .ZN(U2855) );
  AOI21_X1 U5657 ( .B1(n6056), .B2(n4539), .A(n6804), .ZN(n4546) );
  AND2_X1 U5658 ( .A1(n6455), .A2(n4310), .ZN(n6207) );
  NAND2_X1 U5659 ( .A1(n6312), .A2(n6207), .ZN(n6113) );
  OR2_X1 U5660 ( .A1(n6113), .A2(n3915), .ZN(n4540) );
  NAND2_X1 U5661 ( .A1(n6210), .A2(n6302), .ZN(n6111) );
  OR2_X1 U5662 ( .A1(n6111), .A2(n6304), .ZN(n4570) );
  NAND2_X1 U5663 ( .A1(n4540), .A2(n4570), .ZN(n4548) );
  INV_X1 U5664 ( .A(n6111), .ZN(n4541) );
  AOI22_X1 U5665 ( .A1(n4546), .A2(n4548), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4541), .ZN(n4575) );
  AND2_X1 U5666 ( .A1(n6056), .A2(n6246), .ZN(n4543) );
  INV_X1 U5667 ( .A(n4583), .ZN(n4670) );
  NAND3_X1 U5668 ( .A1(n6056), .A2(n3912), .A3(n6203), .ZN(n4544) );
  OAI22_X1 U5669 ( .A1(n6107), .A2(n6714), .B1(n6708), .B2(n4570), .ZN(n4545)
         );
  AOI21_X1 U5670 ( .B1(n6342), .B2(n4779), .A(n4545), .ZN(n4551) );
  INV_X1 U5671 ( .A(n4546), .ZN(n4549) );
  INV_X1 U5672 ( .A(n6210), .ZN(n4547) );
  AOI21_X1 U5673 ( .B1(n4547), .B2(n6804), .A(n6164), .ZN(n6669) );
  OAI211_X1 U5674 ( .C1(n4549), .C2(n4548), .A(n6669), .B(n6302), .ZN(n4572)
         );
  NAND2_X1 U5675 ( .A1(n4572), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4550) );
  OAI211_X1 U5676 ( .C1(n4575), .C2(n6340), .A(n4551), .B(n4550), .ZN(U3049)
         );
  OAI22_X1 U5677 ( .A1(n6107), .A2(n6679), .B1(n6660), .B2(n4570), .ZN(n4552)
         );
  AOI21_X1 U5678 ( .B1(n6308), .B2(n4779), .A(n4552), .ZN(n4554) );
  NAND2_X1 U5679 ( .A1(n4572), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4553) );
  OAI211_X1 U5680 ( .C1(n4575), .C2(n6306), .A(n4554), .B(n4553), .ZN(U3044)
         );
  OAI22_X1 U5681 ( .A1(n6107), .A2(n6707), .B1(n6701), .B2(n4570), .ZN(n4555)
         );
  AOI21_X1 U5682 ( .B1(n6337), .B2(n4779), .A(n4555), .ZN(n4557) );
  NAND2_X1 U5683 ( .A1(n4572), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4556) );
  OAI211_X1 U5684 ( .C1(n4575), .C2(n6335), .A(n4557), .B(n4556), .ZN(U3048)
         );
  OAI22_X1 U5685 ( .A1(n6107), .A2(n6695), .B1(n6694), .B2(n4570), .ZN(n4558)
         );
  AOI21_X1 U5686 ( .B1(n6332), .B2(n4779), .A(n4558), .ZN(n4560) );
  NAND2_X1 U5687 ( .A1(n4572), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4559) );
  OAI211_X1 U5688 ( .C1(n4575), .C2(n6330), .A(n4560), .B(n4559), .ZN(U3047)
         );
  OAI22_X1 U5689 ( .A1(n6107), .A2(n6733), .B1(n6723), .B2(n4570), .ZN(n4561)
         );
  AOI21_X1 U5690 ( .B1(n6355), .B2(n4779), .A(n4561), .ZN(n4563) );
  NAND2_X1 U5691 ( .A1(n4572), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4562) );
  OAI211_X1 U5692 ( .C1(n4575), .C2(n6351), .A(n4563), .B(n4562), .ZN(U3051)
         );
  OAI22_X1 U5693 ( .A1(n6107), .A2(n6681), .B1(n6680), .B2(n4570), .ZN(n4564)
         );
  AOI21_X1 U5694 ( .B1(n6322), .B2(n4779), .A(n4564), .ZN(n4566) );
  NAND2_X1 U5695 ( .A1(n4572), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4565) );
  OAI211_X1 U5696 ( .C1(n4575), .C2(n6320), .A(n4566), .B(n4565), .ZN(U3045)
         );
  OAI22_X1 U5697 ( .A1(n6107), .A2(n6721), .B1(n6715), .B2(n4570), .ZN(n4567)
         );
  AOI21_X1 U5698 ( .B1(n6347), .B2(n4779), .A(n4567), .ZN(n4569) );
  NAND2_X1 U5699 ( .A1(n4572), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4568) );
  OAI211_X1 U5700 ( .C1(n4575), .C2(n6345), .A(n4569), .B(n4568), .ZN(U3050)
         );
  OAI22_X1 U5701 ( .A1(n6107), .A2(n6693), .B1(n6687), .B2(n4570), .ZN(n4571)
         );
  AOI21_X1 U5702 ( .B1(n6327), .B2(n4779), .A(n4571), .ZN(n4574) );
  NAND2_X1 U5703 ( .A1(n4572), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4573) );
  OAI211_X1 U5704 ( .C1(n4575), .C2(n6325), .A(n4574), .B(n4573), .ZN(U3046)
         );
  INV_X1 U5705 ( .A(n4576), .ZN(n4577) );
  OAI21_X1 U5706 ( .B1(n4578), .B2(n4314), .A(n4577), .ZN(n6051) );
  NOR2_X1 U5707 ( .A1(n6051), .A2(FLUSH_REG_SCAN_IN), .ZN(n4580) );
  INV_X1 U5708 ( .A(n4673), .ZN(n4579) );
  OAI21_X1 U5709 ( .B1(n4580), .B2(n4741), .A(n4579), .ZN(n6658) );
  INV_X1 U5710 ( .A(n6658), .ZN(n4587) );
  INV_X1 U5711 ( .A(n6203), .ZN(n6156) );
  NAND3_X1 U5712 ( .A1(n4853), .A2(STATEBS16_REG_SCAN_IN), .A3(n4581), .ZN(
        n4837) );
  NAND3_X1 U5713 ( .A1(n4837), .A2(n6665), .A3(n4582), .ZN(n4584) );
  NAND2_X1 U5714 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6260), .ZN(n6049) );
  INV_X1 U5715 ( .A(n6108), .ZN(n4894) );
  AOI222_X1 U5716 ( .A1(n4584), .A2(n6663), .B1(n6206), .B2(n6049), .C1(n4583), 
        .C2(n4894), .ZN(n4586) );
  NAND2_X1 U5717 ( .A1(n4587), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4585) );
  OAI21_X1 U5718 ( .B1(n4587), .B2(n4586), .A(n4585), .ZN(U3462) );
  XNOR2_X1 U5719 ( .A(n6578), .B(n6579), .ZN(n4589) );
  XNOR2_X1 U5720 ( .A(n4589), .B(n4588), .ZN(n6593) );
  NAND2_X1 U5721 ( .A1(n6577), .A2(REIP_REG_2__SCAN_IN), .ZN(n6589) );
  NAND2_X1 U5722 ( .A1(n6636), .A2(n6644), .ZN(n4590) );
  OAI211_X1 U5723 ( .C1(n6640), .C2(n4591), .A(n6589), .B(n4590), .ZN(n4600)
         );
  NOR2_X1 U5724 ( .A1(n4592), .A2(n6628), .ZN(n4598) );
  NAND2_X1 U5725 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4828) );
  AOI21_X1 U5726 ( .B1(n4593), .B2(n4828), .A(n6043), .ZN(n4594) );
  INV_X1 U5727 ( .A(n4594), .ZN(n6635) );
  AOI21_X1 U5728 ( .B1(n6636), .B2(n4595), .A(n6635), .ZN(n4596) );
  INV_X1 U5729 ( .A(n4596), .ZN(n4597) );
  MUX2_X1 U5730 ( .A(n4598), .B(n4597), .S(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .Z(n4599) );
  AOI211_X1 U5731 ( .C1(n6653), .C2(n6593), .A(n4600), .B(n4599), .ZN(n4601)
         );
  INV_X1 U5732 ( .A(n4601), .ZN(U3016) );
  AND2_X1 U5733 ( .A1(n4851), .A2(n6071), .ZN(n4602) );
  OAI21_X1 U5734 ( .B1(n6151), .B2(n6150), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4603) );
  NAND3_X1 U5735 ( .A1(n4603), .A2(n6663), .A3(n4610), .ZN(n4607) );
  NAND2_X1 U5736 ( .A1(n6301), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4604) );
  NAND2_X1 U5737 ( .A1(n4605), .A2(n6304), .ZN(n4611) );
  AOI21_X1 U5738 ( .B1(n4611), .B2(STATE2_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4606) );
  NOR2_X1 U5739 ( .A1(n4608), .A2(n6673), .ZN(n6262) );
  INV_X1 U5740 ( .A(n6262), .ZN(n6315) );
  INV_X1 U5741 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4615) );
  INV_X1 U5742 ( .A(n6151), .ZN(n4765) );
  NAND2_X1 U5743 ( .A1(n4608), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6300) );
  INV_X1 U5744 ( .A(n6300), .ZN(n6213) );
  INV_X1 U5745 ( .A(n6301), .ZN(n4786) );
  NAND3_X1 U5746 ( .A1(n6213), .A2(n4786), .A3(n6302), .ZN(n4609) );
  OAI21_X1 U5747 ( .B1(n4610), .B2(n6804), .A(n4609), .ZN(n6148) );
  INV_X1 U5748 ( .A(n6680), .ZN(n6172) );
  INV_X1 U5749 ( .A(n4611), .ZN(n6147) );
  AOI22_X1 U5750 ( .A1(n6683), .A2(n6148), .B1(n6172), .B2(n6147), .ZN(n4612)
         );
  OAI21_X1 U5751 ( .B1(n4765), .B2(n6686), .A(n4612), .ZN(n4613) );
  AOI21_X1 U5752 ( .B1(n4929), .B2(n6150), .A(n4613), .ZN(n4614) );
  OAI21_X1 U5753 ( .B1(n4742), .B2(n4615), .A(n4614), .ZN(U3069) );
  NAND3_X1 U5754 ( .A1(n4853), .A2(n4851), .A3(STATEBS16_REG_SCAN_IN), .ZN(
        n4616) );
  NAND2_X1 U5755 ( .A1(n4616), .A2(n6663), .ZN(n4623) );
  INV_X1 U5756 ( .A(n4623), .ZN(n4620) );
  NOR2_X1 U5757 ( .A1(n6455), .A2(n4310), .ZN(n4838) );
  NOR2_X1 U5758 ( .A1(n3915), .A2(n4780), .ZN(n4617) );
  NAND2_X1 U5759 ( .A1(n4839), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4843) );
  OR2_X1 U5760 ( .A1(n4843), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4621)
         );
  NOR2_X1 U5761 ( .A1(n4621), .A2(n6304), .ZN(n4651) );
  AOI21_X1 U5762 ( .B1(n4838), .B2(n4617), .A(n4651), .ZN(n4622) );
  INV_X1 U5763 ( .A(n4621), .ZN(n4782) );
  OAI21_X1 U5764 ( .B1(n6663), .B2(n4782), .A(n4618), .ZN(n4619) );
  INV_X1 U5765 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4628) );
  OAI22_X1 U5766 ( .A1(n4623), .A2(n4622), .B1(n6673), .B2(n4621), .ZN(n4655)
         );
  AND2_X1 U5767 ( .A1(n4851), .A2(n3912), .ZN(n4624) );
  AOI22_X1 U5768 ( .A1(n6150), .A2(n6327), .B1(n3152), .B2(n4651), .ZN(n4625)
         );
  OAI21_X1 U5769 ( .B1(n6693), .B2(n4653), .A(n4625), .ZN(n4626) );
  AOI21_X1 U5770 ( .B1(n6690), .B2(n4655), .A(n4626), .ZN(n4627) );
  OAI21_X1 U5771 ( .B1(n4658), .B2(n4628), .A(n4627), .ZN(U3062) );
  INV_X1 U5772 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4632) );
  AOI22_X1 U5773 ( .A1(n6150), .A2(n6322), .B1(n6172), .B2(n4651), .ZN(n4629)
         );
  OAI21_X1 U5774 ( .B1(n6681), .B2(n4653), .A(n4629), .ZN(n4630) );
  AOI21_X1 U5775 ( .B1(n6683), .B2(n4655), .A(n4630), .ZN(n4631) );
  OAI21_X1 U5776 ( .B1(n4658), .B2(n4632), .A(n4631), .ZN(U3061) );
  INV_X1 U5777 ( .A(n6701), .ZN(n6183) );
  AOI22_X1 U5778 ( .A1(n6150), .A2(n6337), .B1(n6183), .B2(n4651), .ZN(n4633)
         );
  OAI21_X1 U5779 ( .B1(n6707), .B2(n4653), .A(n4633), .ZN(n4634) );
  AOI21_X1 U5780 ( .B1(n6704), .B2(n4655), .A(n4634), .ZN(n4635) );
  OAI21_X1 U5781 ( .B1(n4658), .B2(n6889), .A(n4635), .ZN(U3064) );
  INV_X1 U5782 ( .A(n6708), .ZN(n6187) );
  AOI22_X1 U5783 ( .A1(n6150), .A2(n6342), .B1(n6187), .B2(n4651), .ZN(n4636)
         );
  OAI21_X1 U5784 ( .B1(n6714), .B2(n4653), .A(n4636), .ZN(n4637) );
  AOI21_X1 U5785 ( .B1(n6711), .B2(n4655), .A(n4637), .ZN(n4638) );
  OAI21_X1 U5786 ( .B1(n4658), .B2(n7095), .A(n4638), .ZN(U3065) );
  INV_X1 U5787 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4642) );
  INV_X1 U5788 ( .A(n6715), .ZN(n6191) );
  AOI22_X1 U5789 ( .A1(n6150), .A2(n6347), .B1(n6191), .B2(n4651), .ZN(n4639)
         );
  OAI21_X1 U5790 ( .B1(n6721), .B2(n4653), .A(n4639), .ZN(n4640) );
  AOI21_X1 U5791 ( .B1(n6718), .B2(n4655), .A(n4640), .ZN(n4641) );
  OAI21_X1 U5792 ( .B1(n4658), .B2(n4642), .A(n4641), .ZN(U3066) );
  INV_X1 U5793 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4646) );
  INV_X1 U5794 ( .A(n6723), .ZN(n6197) );
  AOI22_X1 U5795 ( .A1(n6150), .A2(n6355), .B1(n6197), .B2(n4651), .ZN(n4643)
         );
  OAI21_X1 U5796 ( .B1(n6733), .B2(n4653), .A(n4643), .ZN(n4644) );
  AOI21_X1 U5797 ( .B1(n6728), .B2(n4655), .A(n4644), .ZN(n4645) );
  OAI21_X1 U5798 ( .B1(n4658), .B2(n4646), .A(n4645), .ZN(U3067) );
  INV_X1 U5799 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4650) );
  AOI22_X1 U5800 ( .A1(n6150), .A2(n6308), .B1(n3171), .B2(n4651), .ZN(n4647)
         );
  OAI21_X1 U5801 ( .B1(n6679), .B2(n4653), .A(n4647), .ZN(n4648) );
  AOI21_X1 U5802 ( .B1(n6676), .B2(n4655), .A(n4648), .ZN(n4649) );
  OAI21_X1 U5803 ( .B1(n4658), .B2(n4650), .A(n4649), .ZN(U3060) );
  INV_X1 U5804 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4657) );
  INV_X1 U5805 ( .A(n6694), .ZN(n6179) );
  AOI22_X1 U5806 ( .A1(n6150), .A2(n6332), .B1(n6179), .B2(n4651), .ZN(n4652)
         );
  OAI21_X1 U5807 ( .B1(n6695), .B2(n4653), .A(n4652), .ZN(n4654) );
  AOI21_X1 U5808 ( .B1(n6697), .B2(n4655), .A(n4654), .ZN(n4656) );
  OAI21_X1 U5809 ( .B1(n4658), .B2(n4657), .A(n4656), .ZN(U3063) );
  OAI21_X1 U5810 ( .B1(n4661), .B2(n4659), .A(n4660), .ZN(n6637) );
  INV_X1 U5811 ( .A(n5532), .ZN(n4664) );
  AOI22_X1 U5812 ( .A1(n6591), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .B1(n6577), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n4662) );
  OAI21_X1 U5813 ( .B1(n5527), .B2(n6599), .A(n4662), .ZN(n4663) );
  AOI21_X1 U5814 ( .B1(n4664), .B2(n6594), .A(n4663), .ZN(n4665) );
  OAI21_X1 U5815 ( .B1(n6362), .B2(n6637), .A(n4665), .ZN(U2982) );
  XNOR2_X1 U5816 ( .A(n4769), .B(n4768), .ZN(n6573) );
  INV_X1 U5817 ( .A(n6573), .ZN(n4731) );
  AOI21_X1 U5818 ( .B1(n4667), .B2(n4666), .A(n4776), .ZN(n6626) );
  AOI22_X1 U5819 ( .A1(n6626), .A2(n6477), .B1(EBX_REG_5__SCAN_IN), .B2(n5597), 
        .ZN(n4668) );
  OAI21_X1 U5820 ( .B1(n4731), .B2(n6471), .A(n4668), .ZN(U2854) );
  NAND3_X1 U5821 ( .A1(n6103), .A2(n6663), .A3(n4707), .ZN(n4671) );
  INV_X1 U5822 ( .A(n4310), .ZN(n6054) );
  NAND2_X1 U5823 ( .A1(n6054), .A2(n6455), .ZN(n4893) );
  NOR2_X1 U5824 ( .A1(n6206), .A2(n4893), .ZN(n6068) );
  AOI21_X1 U5825 ( .B1(n4671), .B2(n6108), .A(n6068), .ZN(n4675) );
  NOR2_X1 U5826 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4898) );
  AND2_X1 U5827 ( .A1(n4898), .A2(n6302), .ZN(n6074) );
  AND2_X1 U5828 ( .A1(n6074), .A2(n6304), .ZN(n4676) );
  NAND2_X1 U5829 ( .A1(n4786), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4672) );
  NAND2_X1 U5830 ( .A1(n4673), .A2(n4672), .ZN(n4897) );
  AOI21_X1 U5831 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6249), .A(n4897), .ZN(
        n4784) );
  OAI211_X1 U5832 ( .C1(n4676), .C2(n6260), .A(n4784), .B(n6300), .ZN(n4674)
         );
  INV_X1 U5833 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4680) );
  AND2_X1 U5834 ( .A1(n6262), .A2(n6301), .ZN(n4902) );
  INV_X1 U5835 ( .A(n6249), .ZN(n4787) );
  AOI22_X1 U5836 ( .A1(n6068), .A2(n6663), .B1(n4902), .B2(n4787), .ZN(n4706)
         );
  INV_X1 U5837 ( .A(n4676), .ZN(n4705) );
  OAI22_X1 U5838 ( .A1(n4706), .A2(n6351), .B1(n6723), .B2(n4705), .ZN(n4678)
         );
  NOR2_X1 U5839 ( .A1(n4707), .A2(n6733), .ZN(n4677) );
  AOI211_X1 U5840 ( .C1(n4710), .C2(n6355), .A(n4678), .B(n4677), .ZN(n4679)
         );
  OAI21_X1 U5841 ( .B1(n4713), .B2(n4680), .A(n4679), .ZN(U3027) );
  INV_X1 U5842 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4684) );
  OAI22_X1 U5843 ( .A1(n4706), .A2(n6335), .B1(n6701), .B2(n4705), .ZN(n4682)
         );
  NOR2_X1 U5844 ( .A1(n4707), .A2(n6707), .ZN(n4681) );
  AOI211_X1 U5845 ( .C1(n4710), .C2(n6337), .A(n4682), .B(n4681), .ZN(n4683)
         );
  OAI21_X1 U5846 ( .B1(n4713), .B2(n4684), .A(n4683), .ZN(U3024) );
  INV_X1 U5847 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4688) );
  OAI22_X1 U5848 ( .A1(n4706), .A2(n6306), .B1(n6660), .B2(n4705), .ZN(n4686)
         );
  NOR2_X1 U5849 ( .A1(n4707), .A2(n6679), .ZN(n4685) );
  AOI211_X1 U5850 ( .C1(n4710), .C2(n6308), .A(n4686), .B(n4685), .ZN(n4687)
         );
  OAI21_X1 U5851 ( .B1(n4713), .B2(n4688), .A(n4687), .ZN(U3020) );
  INV_X1 U5852 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4692) );
  OAI22_X1 U5853 ( .A1(n4706), .A2(n6345), .B1(n6715), .B2(n4705), .ZN(n4690)
         );
  NOR2_X1 U5854 ( .A1(n4707), .A2(n6721), .ZN(n4689) );
  AOI211_X1 U5855 ( .C1(n4710), .C2(n6347), .A(n4690), .B(n4689), .ZN(n4691)
         );
  OAI21_X1 U5856 ( .B1(n4713), .B2(n4692), .A(n4691), .ZN(U3026) );
  INV_X1 U5857 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4696) );
  OAI22_X1 U5858 ( .A1(n4706), .A2(n6325), .B1(n6687), .B2(n4705), .ZN(n4694)
         );
  NOR2_X1 U5859 ( .A1(n4707), .A2(n6693), .ZN(n4693) );
  AOI211_X1 U5860 ( .C1(n4710), .C2(n6327), .A(n4694), .B(n4693), .ZN(n4695)
         );
  OAI21_X1 U5861 ( .B1(n4713), .B2(n4696), .A(n4695), .ZN(U3022) );
  INV_X1 U5862 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4700) );
  OAI22_X1 U5863 ( .A1(n4706), .A2(n6330), .B1(n6694), .B2(n4705), .ZN(n4698)
         );
  NOR2_X1 U5864 ( .A1(n4707), .A2(n6695), .ZN(n4697) );
  AOI211_X1 U5865 ( .C1(n4710), .C2(n6332), .A(n4698), .B(n4697), .ZN(n4699)
         );
  OAI21_X1 U5866 ( .B1(n4713), .B2(n4700), .A(n4699), .ZN(U3023) );
  INV_X1 U5867 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4704) );
  OAI22_X1 U5868 ( .A1(n4706), .A2(n6320), .B1(n6680), .B2(n4705), .ZN(n4702)
         );
  NOR2_X1 U5869 ( .A1(n4707), .A2(n6681), .ZN(n4701) );
  AOI211_X1 U5870 ( .C1(n4710), .C2(n6322), .A(n4702), .B(n4701), .ZN(n4703)
         );
  OAI21_X1 U5871 ( .B1(n4713), .B2(n4704), .A(n4703), .ZN(U3021) );
  INV_X1 U5872 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4712) );
  OAI22_X1 U5873 ( .A1(n4706), .A2(n6340), .B1(n6708), .B2(n4705), .ZN(n4709)
         );
  NOR2_X1 U5874 ( .A1(n4707), .A2(n6714), .ZN(n4708) );
  AOI211_X1 U5875 ( .C1(n4710), .C2(n6342), .A(n4709), .B(n4708), .ZN(n4711)
         );
  OAI21_X1 U5876 ( .B1(n4713), .B2(n4712), .A(n4711), .ZN(U3025) );
  OR2_X1 U5877 ( .A1(n4715), .A2(n4714), .ZN(n4724) );
  NAND2_X1 U5878 ( .A1(n4737), .A2(n4716), .ZN(n4720) );
  NAND4_X1 U5879 ( .A1(n5266), .A2(n4717), .A3(n4737), .A4(n3398), .ZN(n4718)
         );
  OAI22_X1 U5880 ( .A1(n4721), .A2(n4720), .B1(n4719), .B2(n4718), .ZN(n4722)
         );
  INV_X1 U5881 ( .A(n4722), .ZN(n4723) );
  NAND2_X1 U5882 ( .A1(n4726), .A2(n3400), .ZN(n4727) );
  NAND2_X2 U5883 ( .A1(n5664), .A2(n4727), .ZN(n5662) );
  INV_X1 U5884 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4730) );
  INV_X1 U5885 ( .A(DATAI_5_), .ZN(n6540) );
  AND2_X1 U5886 ( .A1(n3387), .A2(n3400), .ZN(n4729) );
  OAI222_X1 U5887 ( .A1(n5662), .A2(n4731), .B1(n5664), .B2(n4730), .C1(n6540), 
        .C2(n5665), .ZN(U2886) );
  OAI21_X1 U5888 ( .B1(n4732), .B2(n6061), .A(n6741), .ZN(n4734) );
  AOI21_X1 U5889 ( .B1(n6673), .B2(READY_N), .A(n4733), .ZN(n6734) );
  MUX2_X1 U5890 ( .A(n4734), .B(n6734), .S(STATE2_REG_0__SCAN_IN), .Z(n4740)
         );
  AND2_X1 U5891 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n4735) );
  NAND2_X1 U5892 ( .A1(n6803), .A2(n4735), .ZN(n5043) );
  INV_X1 U5893 ( .A(n5043), .ZN(n4736) );
  AOI21_X1 U5894 ( .B1(n4738), .B2(n4737), .A(n4736), .ZN(n4739) );
  OAI211_X1 U5895 ( .C1(n4741), .C2(n6051), .A(n4740), .B(n4739), .ZN(U3148)
         );
  AOI22_X1 U5896 ( .A1(n6711), .A2(n6148), .B1(n6187), .B2(n6147), .ZN(n4744)
         );
  NAND2_X1 U5897 ( .A1(n6150), .A2(n4922), .ZN(n4743) );
  OAI211_X1 U5898 ( .C1(n4765), .C2(n6709), .A(n4744), .B(n4743), .ZN(n4745)
         );
  AOI21_X1 U5899 ( .B1(n6146), .B2(INSTQUEUE_REG_6__5__SCAN_IN), .A(n4745), 
        .ZN(n4746) );
  INV_X1 U5900 ( .A(n4746), .ZN(U3073) );
  AOI22_X1 U5901 ( .A1(n6697), .A2(n6148), .B1(n6179), .B2(n6147), .ZN(n4748)
         );
  NAND2_X1 U5902 ( .A1(n6150), .A2(n4918), .ZN(n4747) );
  OAI211_X1 U5903 ( .C1(n4765), .C2(n6700), .A(n4748), .B(n4747), .ZN(n4749)
         );
  AOI21_X1 U5904 ( .B1(n6146), .B2(INSTQUEUE_REG_6__3__SCAN_IN), .A(n4749), 
        .ZN(n4750) );
  INV_X1 U5905 ( .A(n4750), .ZN(U3071) );
  AOI22_X1 U5906 ( .A1(n6728), .A2(n6148), .B1(n6197), .B2(n6147), .ZN(n4752)
         );
  NAND2_X1 U5907 ( .A1(n6150), .A2(n4910), .ZN(n4751) );
  OAI211_X1 U5908 ( .C1(n4765), .C2(n6724), .A(n4752), .B(n4751), .ZN(n4753)
         );
  AOI21_X1 U5909 ( .B1(n6146), .B2(INSTQUEUE_REG_6__7__SCAN_IN), .A(n4753), 
        .ZN(n4754) );
  INV_X1 U5910 ( .A(n4754), .ZN(U3075) );
  AOI22_X1 U5911 ( .A1(n6718), .A2(n6148), .B1(n6191), .B2(n6147), .ZN(n4756)
         );
  NAND2_X1 U5912 ( .A1(n6150), .A2(n4906), .ZN(n4755) );
  OAI211_X1 U5913 ( .C1(n4765), .C2(n6716), .A(n4756), .B(n4755), .ZN(n4757)
         );
  AOI21_X1 U5914 ( .B1(n6146), .B2(INSTQUEUE_REG_6__6__SCAN_IN), .A(n4757), 
        .ZN(n4758) );
  INV_X1 U5915 ( .A(n4758), .ZN(U3074) );
  AOI22_X1 U5916 ( .A1(n6690), .A2(n6148), .B1(n3152), .B2(n6147), .ZN(n4760)
         );
  NAND2_X1 U5917 ( .A1(n6150), .A2(n4914), .ZN(n4759) );
  OAI211_X1 U5918 ( .C1(n4765), .C2(n6688), .A(n4760), .B(n4759), .ZN(n4761)
         );
  AOI21_X1 U5919 ( .B1(n6146), .B2(INSTQUEUE_REG_6__2__SCAN_IN), .A(n4761), 
        .ZN(n4762) );
  INV_X1 U5920 ( .A(n4762), .ZN(U3070) );
  AOI22_X1 U5921 ( .A1(n6704), .A2(n6148), .B1(n6183), .B2(n6147), .ZN(n4764)
         );
  NAND2_X1 U5922 ( .A1(n6150), .A2(n4936), .ZN(n4763) );
  OAI211_X1 U5923 ( .C1(n4765), .C2(n6702), .A(n4764), .B(n4763), .ZN(n4766)
         );
  AOI21_X1 U5924 ( .B1(n6146), .B2(INSTQUEUE_REG_6__4__SCAN_IN), .A(n4766), 
        .ZN(n4767) );
  INV_X1 U5925 ( .A(n4767), .ZN(U3072) );
  INV_X1 U5926 ( .A(n4768), .ZN(n4770) );
  OR2_X1 U5927 ( .A1(n4770), .A2(n4769), .ZN(n4773) );
  INV_X1 U5928 ( .A(n4771), .ZN(n4772) );
  NAND2_X1 U5929 ( .A1(n4773), .A2(n4772), .ZN(n4774) );
  AND2_X1 U5930 ( .A1(n4774), .A2(n4884), .ZN(n4826) );
  OR2_X1 U5931 ( .A1(n4776), .A2(n4775), .ZN(n4777) );
  NAND2_X1 U5932 ( .A1(n4887), .A2(n4777), .ZN(n6439) );
  INV_X1 U5933 ( .A(n6439), .ZN(n4834) );
  AOI22_X1 U5934 ( .A1(n6477), .A2(n4834), .B1(EBX_REG_6__SCAN_IN), .B2(n5597), 
        .ZN(n4778) );
  OAI21_X1 U5935 ( .B1(n6434), .B2(n6471), .A(n4778), .ZN(U2853) );
  NOR3_X1 U5936 ( .A1(n4779), .A2(n4815), .A3(n6804), .ZN(n4781) );
  INV_X1 U5937 ( .A(n4838), .ZN(n6257) );
  OAI22_X1 U5938 ( .A1(n4781), .A2(n4894), .B1(n4780), .B2(n6257), .ZN(n4785)
         );
  NAND2_X1 U5939 ( .A1(n4782), .A2(n6304), .ZN(n4812) );
  AOI21_X1 U5940 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n4812), .A(n6262), .ZN(
        n4783) );
  NAND3_X1 U5941 ( .A1(n4785), .A2(n4784), .A3(n4783), .ZN(n4811) );
  NAND2_X1 U5942 ( .A1(n4811), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4792) );
  NAND2_X1 U5943 ( .A1(n4838), .A2(n6663), .ZN(n6248) );
  OR2_X1 U5944 ( .A1(n6248), .A2(n6206), .ZN(n4789) );
  NOR2_X1 U5945 ( .A1(n6300), .A2(n4786), .ZN(n6250) );
  NAND2_X1 U5946 ( .A1(n4787), .A2(n6250), .ZN(n4788) );
  OAI22_X1 U5947 ( .A1(n4813), .A2(n6335), .B1(n6701), .B2(n4812), .ZN(n4790)
         );
  AOI21_X1 U5948 ( .B1(n4815), .B2(n6337), .A(n4790), .ZN(n4791) );
  OAI211_X1 U5949 ( .C1(n4818), .C2(n6707), .A(n4792), .B(n4791), .ZN(U3056)
         );
  NAND2_X1 U5950 ( .A1(n4811), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4795) );
  OAI22_X1 U5951 ( .A1(n4813), .A2(n6345), .B1(n6715), .B2(n4812), .ZN(n4793)
         );
  AOI21_X1 U5952 ( .B1(n4815), .B2(n6347), .A(n4793), .ZN(n4794) );
  OAI211_X1 U5953 ( .C1(n4818), .C2(n6721), .A(n4795), .B(n4794), .ZN(U3058)
         );
  NAND2_X1 U5954 ( .A1(n4811), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4798) );
  OAI22_X1 U5955 ( .A1(n4813), .A2(n6320), .B1(n6680), .B2(n4812), .ZN(n4796)
         );
  AOI21_X1 U5956 ( .B1(n4815), .B2(n6322), .A(n4796), .ZN(n4797) );
  OAI211_X1 U5957 ( .C1(n4818), .C2(n6681), .A(n4798), .B(n4797), .ZN(U3053)
         );
  NAND2_X1 U5958 ( .A1(n4811), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4801) );
  OAI22_X1 U5959 ( .A1(n4813), .A2(n6351), .B1(n6723), .B2(n4812), .ZN(n4799)
         );
  AOI21_X1 U5960 ( .B1(n4815), .B2(n6355), .A(n4799), .ZN(n4800) );
  OAI211_X1 U5961 ( .C1(n4818), .C2(n6733), .A(n4801), .B(n4800), .ZN(U3059)
         );
  NAND2_X1 U5962 ( .A1(n4811), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4804) );
  OAI22_X1 U5963 ( .A1(n4813), .A2(n6330), .B1(n6694), .B2(n4812), .ZN(n4802)
         );
  AOI21_X1 U5964 ( .B1(n4815), .B2(n6332), .A(n4802), .ZN(n4803) );
  OAI211_X1 U5965 ( .C1(n4818), .C2(n6695), .A(n4804), .B(n4803), .ZN(U3055)
         );
  NAND2_X1 U5966 ( .A1(n4811), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4807) );
  OAI22_X1 U5967 ( .A1(n4813), .A2(n6325), .B1(n6687), .B2(n4812), .ZN(n4805)
         );
  AOI21_X1 U5968 ( .B1(n4815), .B2(n6327), .A(n4805), .ZN(n4806) );
  OAI211_X1 U5969 ( .C1(n4818), .C2(n6693), .A(n4807), .B(n4806), .ZN(U3054)
         );
  NAND2_X1 U5970 ( .A1(n4811), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4810) );
  OAI22_X1 U5971 ( .A1(n4813), .A2(n6306), .B1(n6660), .B2(n4812), .ZN(n4808)
         );
  AOI21_X1 U5972 ( .B1(n4815), .B2(n6308), .A(n4808), .ZN(n4809) );
  OAI211_X1 U5973 ( .C1(n4818), .C2(n6679), .A(n4810), .B(n4809), .ZN(U3052)
         );
  NAND2_X1 U5974 ( .A1(n4811), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4817) );
  OAI22_X1 U5975 ( .A1(n4813), .A2(n6340), .B1(n6708), .B2(n4812), .ZN(n4814)
         );
  AOI21_X1 U5976 ( .B1(n4815), .B2(n6342), .A(n4814), .ZN(n4816) );
  OAI211_X1 U5977 ( .C1(n4818), .C2(n6714), .A(n4817), .B(n4816), .ZN(U3057)
         );
  XNOR2_X1 U5978 ( .A(n4820), .B(n4819), .ZN(n4821) );
  INV_X1 U5979 ( .A(n6428), .ZN(n4824) );
  INV_X1 U5980 ( .A(REIP_REG_6__SCAN_IN), .ZN(n4822) );
  NOR2_X1 U5981 ( .A1(n6639), .A2(n4822), .ZN(n4833) );
  AOI21_X1 U5982 ( .B1(n6591), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n4833), 
        .ZN(n4823) );
  OAI21_X1 U5983 ( .B1(n4824), .B2(n6599), .A(n4823), .ZN(n4825) );
  AOI21_X1 U5984 ( .B1(n4826), .B2(n6594), .A(n4825), .ZN(n4827) );
  OAI21_X1 U5985 ( .B1(n4836), .B2(n6362), .A(n4827), .ZN(U2980) );
  OAI21_X1 U5986 ( .B1(n6628), .B2(n4828), .A(n6038), .ZN(n6035) );
  INV_X1 U5987 ( .A(n6035), .ZN(n6643) );
  NOR2_X1 U5988 ( .A1(n4829), .A2(n6643), .ZN(n4831) );
  AOI21_X1 U5989 ( .B1(n4829), .B2(n5967), .A(n6635), .ZN(n6634) );
  INV_X1 U5990 ( .A(n6634), .ZN(n4830) );
  MUX2_X1 U5991 ( .A(n4831), .B(n4830), .S(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .Z(n4832) );
  AOI211_X1 U5992 ( .C1(n6651), .C2(n4834), .A(n4833), .B(n4832), .ZN(n4835)
         );
  OAI21_X1 U5993 ( .B1(n6638), .B2(n4836), .A(n4835), .ZN(U3012) );
  NAND2_X1 U5994 ( .A1(n4837), .A2(n6663), .ZN(n4849) );
  NAND2_X1 U5995 ( .A1(n6159), .A2(n4838), .ZN(n4842) );
  NAND2_X1 U5996 ( .A1(n4840), .A2(n4839), .ZN(n6253) );
  INV_X1 U5997 ( .A(n6253), .ZN(n4841) );
  NAND2_X1 U5998 ( .A1(n4841), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4876) );
  NAND2_X1 U5999 ( .A1(n4842), .A2(n4876), .ZN(n4848) );
  INV_X1 U6000 ( .A(n4848), .ZN(n4845) );
  NAND2_X1 U6001 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4844) );
  OAI22_X1 U6002 ( .A1(n4849), .A2(n4845), .B1(n4844), .B2(n4843), .ZN(n4846)
         );
  AOI21_X1 U6003 ( .B1(n6804), .B2(n6253), .A(n6164), .ZN(n4847) );
  NAND2_X1 U6004 ( .A1(n4875), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4856)
         );
  NOR2_X1 U6005 ( .A1(n4851), .A2(n3912), .ZN(n4850) );
  NOR2_X1 U6006 ( .A1(n4851), .A2(n6071), .ZN(n4852) );
  OAI22_X1 U6007 ( .A1(n6295), .A2(n6695), .B1(n4876), .B2(n6694), .ZN(n4854)
         );
  AOI21_X1 U6008 ( .B1(n6309), .B2(n6332), .A(n4854), .ZN(n4855) );
  OAI211_X1 U6009 ( .C1(n4880), .C2(n6330), .A(n4856), .B(n4855), .ZN(U3127)
         );
  NAND2_X1 U6010 ( .A1(n4875), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4859)
         );
  OAI22_X1 U6011 ( .A1(n6295), .A2(n6693), .B1(n4876), .B2(n6687), .ZN(n4857)
         );
  AOI21_X1 U6012 ( .B1(n6309), .B2(n6327), .A(n4857), .ZN(n4858) );
  OAI211_X1 U6013 ( .C1(n4880), .C2(n6325), .A(n4859), .B(n4858), .ZN(U3126)
         );
  NAND2_X1 U6014 ( .A1(n4875), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4862)
         );
  OAI22_X1 U6015 ( .A1(n6295), .A2(n6681), .B1(n4876), .B2(n6680), .ZN(n4860)
         );
  AOI21_X1 U6016 ( .B1(n6309), .B2(n6322), .A(n4860), .ZN(n4861) );
  OAI211_X1 U6017 ( .C1(n4880), .C2(n6320), .A(n4862), .B(n4861), .ZN(U3125)
         );
  NAND2_X1 U6018 ( .A1(n4875), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4865)
         );
  OAI22_X1 U6019 ( .A1(n6295), .A2(n6679), .B1(n4876), .B2(n6660), .ZN(n4863)
         );
  AOI21_X1 U6020 ( .B1(n6308), .B2(n6309), .A(n4863), .ZN(n4864) );
  OAI211_X1 U6021 ( .C1(n4880), .C2(n6306), .A(n4865), .B(n4864), .ZN(U3124)
         );
  NAND2_X1 U6022 ( .A1(n4875), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4868)
         );
  OAI22_X1 U6023 ( .A1(n6295), .A2(n6714), .B1(n4876), .B2(n6708), .ZN(n4866)
         );
  AOI21_X1 U6024 ( .B1(n6309), .B2(n6342), .A(n4866), .ZN(n4867) );
  OAI211_X1 U6025 ( .C1(n4880), .C2(n6340), .A(n4868), .B(n4867), .ZN(U3129)
         );
  NAND2_X1 U6026 ( .A1(n4875), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4871)
         );
  OAI22_X1 U6027 ( .A1(n6295), .A2(n6733), .B1(n4876), .B2(n6723), .ZN(n4869)
         );
  AOI21_X1 U6028 ( .B1(n6309), .B2(n6355), .A(n4869), .ZN(n4870) );
  OAI211_X1 U6029 ( .C1(n4880), .C2(n6351), .A(n4871), .B(n4870), .ZN(U3131)
         );
  NAND2_X1 U6030 ( .A1(n4875), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4874)
         );
  OAI22_X1 U6031 ( .A1(n6295), .A2(n6721), .B1(n4876), .B2(n6715), .ZN(n4872)
         );
  AOI21_X1 U6032 ( .B1(n6309), .B2(n6347), .A(n4872), .ZN(n4873) );
  OAI211_X1 U6033 ( .C1(n4880), .C2(n6345), .A(n4874), .B(n4873), .ZN(U3130)
         );
  NAND2_X1 U6034 ( .A1(n4875), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4879)
         );
  OAI22_X1 U6035 ( .A1(n6295), .A2(n6707), .B1(n4876), .B2(n6701), .ZN(n4877)
         );
  AOI21_X1 U6036 ( .B1(n6309), .B2(n6337), .A(n4877), .ZN(n4878) );
  OAI211_X1 U6037 ( .C1(n4880), .C2(n6335), .A(n4879), .B(n4878), .ZN(U3128)
         );
  INV_X1 U6038 ( .A(DATAI_4_), .ZN(n6538) );
  INV_X1 U6039 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6505) );
  OAI222_X1 U6040 ( .A1(n5532), .A2(n5662), .B1(n5665), .B2(n6538), .C1(n5664), 
        .C2(n6505), .ZN(U2887) );
  INV_X1 U6041 ( .A(DATAI_0_), .ZN(n6531) );
  INV_X1 U6042 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6513) );
  OAI222_X1 U6043 ( .A1(n5560), .A2(n5662), .B1(n5665), .B2(n6531), .C1(n5664), 
        .C2(n6513), .ZN(U2891) );
  INV_X1 U6044 ( .A(DATAI_1_), .ZN(n6835) );
  INV_X1 U6045 ( .A(EAX_REG_1__SCAN_IN), .ZN(n4881) );
  OAI222_X1 U6046 ( .A1(n5551), .A2(n5662), .B1(n5665), .B2(n6835), .C1(n5664), 
        .C2(n4881), .ZN(U2890) );
  INV_X1 U6047 ( .A(DATAI_2_), .ZN(n6534) );
  INV_X1 U6048 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6509) );
  OAI222_X1 U6049 ( .A1(n4882), .A2(n5662), .B1(n5665), .B2(n6534), .C1(n5664), 
        .C2(n6509), .ZN(U2889) );
  INV_X1 U6050 ( .A(DATAI_6_), .ZN(n6542) );
  OAI222_X1 U6051 ( .A1(n6434), .A2(n5662), .B1(n5665), .B2(n6542), .C1(n5664), 
        .C2(n3941), .ZN(U2885) );
  XNOR2_X1 U6052 ( .A(n4462), .B(n4883), .ZN(n6476) );
  INV_X1 U6053 ( .A(DATAI_3_), .ZN(n6536) );
  INV_X1 U6054 ( .A(EAX_REG_3__SCAN_IN), .ZN(n7108) );
  OAI222_X1 U6055 ( .A1(n6476), .A2(n5662), .B1(n5665), .B2(n6536), .C1(n5664), 
        .C2(n7108), .ZN(U2888) );
  XOR2_X1 U6056 ( .A(n4885), .B(n4884), .Z(n6566) );
  INV_X1 U6057 ( .A(n6566), .ZN(n4940) );
  NAND2_X1 U6058 ( .A1(n4887), .A2(n4886), .ZN(n4888) );
  NAND2_X1 U6059 ( .A1(n5603), .A2(n4888), .ZN(n6617) );
  INV_X1 U6060 ( .A(EBX_REG_7__SCAN_IN), .ZN(n6936) );
  OAI22_X1 U6061 ( .A1(n6617), .A2(n5605), .B1(n6936), .B2(n6480), .ZN(n4889)
         );
  INV_X1 U6062 ( .A(n4889), .ZN(n4890) );
  OAI21_X1 U6063 ( .B1(n4940), .B2(n6471), .A(n4890), .ZN(U2852) );
  OR2_X1 U6064 ( .A1(n6203), .A2(n6071), .ZN(n4891) );
  INV_X1 U6065 ( .A(n6199), .ZN(n4892) );
  NOR3_X1 U6066 ( .A1(n4892), .A2(n4937), .A3(n6804), .ZN(n4895) );
  INV_X1 U6067 ( .A(n4893), .ZN(n6158) );
  NAND2_X1 U6068 ( .A1(n6158), .A2(n6206), .ZN(n4901) );
  OAI21_X1 U6069 ( .B1(n4895), .B2(n4894), .A(n4901), .ZN(n4900) );
  NOR2_X1 U6070 ( .A1(n6249), .A2(n6673), .ZN(n4896) );
  NOR2_X1 U6071 ( .A1(n4897), .A2(n4896), .ZN(n6259) );
  NAND2_X1 U6072 ( .A1(n4898), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6165) );
  OR2_X1 U6073 ( .A1(n6165), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4933)
         );
  AOI21_X1 U6074 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n4933), .A(n6213), .ZN(
        n4899) );
  NAND3_X1 U6075 ( .A1(n4900), .A2(n6259), .A3(n4899), .ZN(n4932) );
  NAND2_X1 U6076 ( .A1(n4932), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4908) );
  OR2_X1 U6077 ( .A1(n4901), .A2(n6804), .ZN(n4904) );
  NAND2_X1 U6078 ( .A1(n4902), .A2(n6249), .ZN(n4903) );
  OAI22_X1 U6079 ( .A1(n4934), .A2(n6345), .B1(n6715), .B2(n4933), .ZN(n4905)
         );
  AOI21_X1 U6080 ( .B1(n4937), .B2(n4906), .A(n4905), .ZN(n4907) );
  OAI211_X1 U6081 ( .C1(n6199), .C2(n6716), .A(n4908), .B(n4907), .ZN(U3090)
         );
  NAND2_X1 U6082 ( .A1(n4932), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4912) );
  OAI22_X1 U6083 ( .A1(n4934), .A2(n6351), .B1(n6723), .B2(n4933), .ZN(n4909)
         );
  AOI21_X1 U6084 ( .B1(n4937), .B2(n4910), .A(n4909), .ZN(n4911) );
  OAI211_X1 U6085 ( .C1(n6199), .C2(n6724), .A(n4912), .B(n4911), .ZN(U3091)
         );
  NAND2_X1 U6086 ( .A1(n4932), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4916) );
  OAI22_X1 U6087 ( .A1(n4934), .A2(n6325), .B1(n6687), .B2(n4933), .ZN(n4913)
         );
  AOI21_X1 U6088 ( .B1(n4937), .B2(n4914), .A(n4913), .ZN(n4915) );
  OAI211_X1 U6089 ( .C1(n6199), .C2(n6688), .A(n4916), .B(n4915), .ZN(U3086)
         );
  NAND2_X1 U6090 ( .A1(n4932), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4920) );
  OAI22_X1 U6091 ( .A1(n4934), .A2(n6330), .B1(n6694), .B2(n4933), .ZN(n4917)
         );
  AOI21_X1 U6092 ( .B1(n4937), .B2(n4918), .A(n4917), .ZN(n4919) );
  OAI211_X1 U6093 ( .C1(n6199), .C2(n6700), .A(n4920), .B(n4919), .ZN(U3087)
         );
  NAND2_X1 U6094 ( .A1(n4932), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4924) );
  OAI22_X1 U6095 ( .A1(n4934), .A2(n6340), .B1(n6708), .B2(n4933), .ZN(n4921)
         );
  AOI21_X1 U6096 ( .B1(n4937), .B2(n4922), .A(n4921), .ZN(n4923) );
  OAI211_X1 U6097 ( .C1(n6199), .C2(n6709), .A(n4924), .B(n4923), .ZN(U3089)
         );
  NAND2_X1 U6098 ( .A1(n4932), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4927) );
  OAI22_X1 U6099 ( .A1(n4934), .A2(n6306), .B1(n6660), .B2(n4933), .ZN(n4925)
         );
  AOI21_X1 U6100 ( .B1(n4937), .B2(n6149), .A(n4925), .ZN(n4926) );
  OAI211_X1 U6101 ( .C1(n6199), .C2(n6661), .A(n4927), .B(n4926), .ZN(U3084)
         );
  NAND2_X1 U6102 ( .A1(n4932), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4931) );
  OAI22_X1 U6103 ( .A1(n4934), .A2(n6320), .B1(n6680), .B2(n4933), .ZN(n4928)
         );
  AOI21_X1 U6104 ( .B1(n4937), .B2(n4929), .A(n4928), .ZN(n4930) );
  OAI211_X1 U6105 ( .C1(n6199), .C2(n6686), .A(n4931), .B(n4930), .ZN(U3085)
         );
  NAND2_X1 U6106 ( .A1(n4932), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4939) );
  OAI22_X1 U6107 ( .A1(n4934), .A2(n6335), .B1(n6701), .B2(n4933), .ZN(n4935)
         );
  AOI21_X1 U6108 ( .B1(n4937), .B2(n4936), .A(n4935), .ZN(n4938) );
  OAI211_X1 U6109 ( .C1(n6199), .C2(n6702), .A(n4939), .B(n4938), .ZN(U3088)
         );
  INV_X1 U6110 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6501) );
  INV_X1 U6111 ( .A(DATAI_7_), .ZN(n6544) );
  OAI222_X1 U6112 ( .A1(n5662), .A2(n4940), .B1(n5664), .B2(n6501), .C1(n6544), 
        .C2(n5665), .ZN(U2884) );
  INV_X1 U6113 ( .A(n4943), .ZN(n4941) );
  AOI21_X1 U6114 ( .B1(n4942), .B2(n4941), .A(n4951), .ZN(n4953) );
  NAND2_X1 U6115 ( .A1(n4943), .A2(n4952), .ZN(n4946) );
  OAI22_X1 U6116 ( .A1(n6061), .A2(n4946), .B1(n4945), .B2(n4944), .ZN(n4947)
         );
  AOI21_X1 U6117 ( .B1(n4949), .B2(n4948), .A(n4947), .ZN(n4950) );
  OAI22_X1 U6118 ( .A1(n4953), .A2(n4952), .B1(n4951), .B2(n4950), .ZN(U3459)
         );
  NAND2_X1 U6119 ( .A1(n4955), .A2(n4954), .ZN(n4959) );
  AND2_X1 U6120 ( .A1(n4957), .A2(n4956), .ZN(n4958) );
  XNOR2_X1 U6121 ( .A(n4959), .B(n4958), .ZN(n4969) );
  NAND2_X1 U6122 ( .A1(n5967), .A2(n4960), .ZN(n4962) );
  AOI21_X1 U6123 ( .B1(n6636), .B2(n6838), .A(n6043), .ZN(n4961) );
  MUX2_X1 U6124 ( .A(n4962), .B(n4961), .S(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .Z(n4964) );
  INV_X1 U6125 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6792) );
  NOR2_X1 U6126 ( .A1(n6639), .A2(n6792), .ZN(n4966) );
  AOI21_X1 U6127 ( .B1(n6651), .B2(n5544), .A(n4966), .ZN(n4963) );
  OAI211_X1 U6128 ( .C1(n4969), .C2(n6638), .A(n4964), .B(n4963), .ZN(U3017)
         );
  INV_X1 U6129 ( .A(n5551), .ZN(n4967) );
  MUX2_X1 U6130 ( .A(n5855), .B(n6591), .S(PHYADDRPOINTER_REG_1__SCAN_IN), .Z(
        n4965) );
  AOI211_X1 U6131 ( .C1(n4967), .C2(n6594), .A(n4966), .B(n4965), .ZN(n4968)
         );
  OAI21_X1 U6132 ( .B1(n4969), .B2(n6362), .A(n4968), .ZN(U2985) );
  NAND2_X1 U6133 ( .A1(n4993), .A2(EBX_REG_30__SCAN_IN), .ZN(n4971) );
  NAND2_X1 U6134 ( .A1(n3764), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4970) );
  AND2_X1 U6135 ( .A1(n4971), .A2(n4970), .ZN(n5049) );
  OAI21_X1 U6136 ( .B1(INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n4993), .A(n4972), 
        .ZN(n5027) );
  INV_X1 U6137 ( .A(n5027), .ZN(n4973) );
  INV_X1 U6138 ( .A(EBX_REG_25__SCAN_IN), .ZN(n6832) );
  NAND2_X1 U6139 ( .A1(n3763), .A2(n6832), .ZN(n4976) );
  INV_X1 U6140 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n7061) );
  NAND2_X1 U6141 ( .A1(n3771), .A2(n7061), .ZN(n4974) );
  OAI211_X1 U6142 ( .C1(EBX_REG_25__SCAN_IN), .C2(n3764), .A(n4974), .B(n5050), 
        .ZN(n4975) );
  AND2_X1 U6143 ( .A1(n4976), .A2(n4975), .ZN(n5319) );
  INV_X1 U6144 ( .A(EBX_REG_26__SCAN_IN), .ZN(n7040) );
  NAND2_X1 U6145 ( .A1(n3098), .A2(n7040), .ZN(n4979) );
  OAI211_X1 U6146 ( .C1(n3764), .C2(EBX_REG_26__SCAN_IN), .A(n3771), .B(n4977), 
        .ZN(n4978) );
  AND2_X1 U6147 ( .A1(n4979), .A2(n4978), .ZN(n5304) );
  MUX2_X1 U6148 ( .A(n4980), .B(n3771), .S(EBX_REG_27__SCAN_IN), .Z(n4982) );
  NAND2_X1 U6149 ( .A1(n3764), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4981) );
  NAND2_X1 U6150 ( .A1(n4982), .A2(n4981), .ZN(n5299) );
  INV_X1 U6151 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U6152 ( .A1(n3098), .A2(n5564), .ZN(n4985) );
  NAND2_X1 U6153 ( .A1(n5050), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4983) );
  OAI211_X1 U6154 ( .C1(n3764), .C2(EBX_REG_28__SCAN_IN), .A(n3771), .B(n4983), 
        .ZN(n4984) );
  AND2_X1 U6155 ( .A1(n4985), .A2(n4984), .ZN(n5283) );
  AND2_X1 U6156 ( .A1(n5299), .A2(n5283), .ZN(n4986) );
  NOR2_X1 U6157 ( .A1(n4993), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4992)
         );
  MUX2_X1 U6158 ( .A(EBX_REG_29__SCAN_IN), .B(n4992), .S(n5050), .Z(n4989) );
  NOR2_X1 U6159 ( .A1(n4987), .A2(EBX_REG_29__SCAN_IN), .ZN(n4988) );
  NOR2_X1 U6160 ( .A1(n4989), .A2(n4988), .ZN(n5275) );
  INV_X1 U6161 ( .A(EBX_REG_29__SCAN_IN), .ZN(n4990) );
  AOI22_X1 U6162 ( .A1(n4993), .A2(EBX_REG_31__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n3764), .ZN(n4994) );
  INV_X1 U6163 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5199) );
  OAI22_X1 U6164 ( .A1(n5265), .A2(n5605), .B1(n6480), .B2(n5199), .ZN(U2828)
         );
  INV_X1 U6165 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5034) );
  NAND4_X1 U6166 ( .A1(n5824), .A2(n5217), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .A4(n5034), .ZN(n4996) );
  OAI21_X1 U6167 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5034), .A(n4996), 
        .ZN(n5003) );
  NOR2_X1 U6168 ( .A1(n5720), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4997)
         );
  AND2_X1 U6169 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5216) );
  AOI21_X1 U6170 ( .B1(n4997), .B2(n5034), .A(n5216), .ZN(n5001) );
  INV_X1 U6171 ( .A(n4997), .ZN(n4999) );
  NAND3_X1 U6172 ( .A1(n5815), .A2(n5217), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4998) );
  NAND3_X1 U6173 ( .A1(n4999), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .A3(n4998), .ZN(n5000) );
  OAI21_X1 U6174 ( .B1(n5729), .B2(n5001), .A(n5000), .ZN(n5002) );
  AOI21_X1 U6175 ( .B1(n5729), .B2(n5003), .A(n5002), .ZN(n5038) );
  INV_X1 U6176 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5004) );
  XNOR2_X1 U6177 ( .A(n5057), .B(n5004), .ZN(n5338) );
  NOR2_X1 U6178 ( .A1(n5006), .A2(n5005), .ZN(n5092) );
  AOI22_X1 U6179 ( .A1(n5121), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n5107), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5011) );
  AOI22_X1 U6180 ( .A1(n5116), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n5124), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n5010) );
  AOI22_X1 U6181 ( .A1(n3467), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5009) );
  AOI22_X1 U6182 ( .A1(n5122), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5008) );
  NAND4_X1 U6183 ( .A1(n5011), .A2(n5010), .A3(n5009), .A4(n5008), .ZN(n5017)
         );
  AOI22_X1 U6184 ( .A1(n3496), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3486), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5015) );
  AOI22_X1 U6185 ( .A1(n5123), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n5114), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5014) );
  AOI22_X1 U6186 ( .A1(n3462), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5115), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n5013) );
  AOI22_X1 U6187 ( .A1(n3086), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n5012) );
  NAND4_X1 U6188 ( .A1(n5015), .A2(n5014), .A3(n5013), .A4(n5012), .ZN(n5016)
         );
  OR2_X1 U6189 ( .A1(n5017), .A2(n5016), .ZN(n5091) );
  XNOR2_X1 U6190 ( .A(n5092), .B(n5091), .ZN(n5019) );
  AOI22_X1 U6191 ( .A1(n4168), .A2(EAX_REG_24__SCAN_IN), .B1(n5245), .B2(
        PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5018) );
  OAI21_X1 U6192 ( .B1(n5019), .B2(n5177), .A(n5018), .ZN(n5020) );
  AOI21_X1 U6193 ( .B1(n5338), .B2(n5182), .A(n5020), .ZN(n5022) );
  OR2_X2 U6194 ( .A1(n5021), .A2(n5022), .ZN(n5148) );
  INV_X1 U6195 ( .A(n5148), .ZN(n5326) );
  AOI21_X1 U6196 ( .B1(n5022), .B2(n5021), .A(n5326), .ZN(n5566) );
  INV_X1 U6197 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6773) );
  NOR2_X1 U6198 ( .A1(n6639), .A2(n6773), .ZN(n5036) );
  AOI21_X1 U6199 ( .B1(n6591), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5036), 
        .ZN(n5023) );
  OAI21_X1 U6200 ( .B1(n5338), .B2(n6599), .A(n5023), .ZN(n5024) );
  AOI21_X1 U6201 ( .B1(n5566), .B2(n5839), .A(n5024), .ZN(n5025) );
  OAI21_X1 U6202 ( .B1(n5038), .B2(n6362), .A(n5025), .ZN(U2962) );
  INV_X1 U6203 ( .A(n5026), .ZN(n5028) );
  OAI21_X1 U6204 ( .B1(n5349), .B2(n5028), .A(n5027), .ZN(n5029) );
  AND2_X1 U6205 ( .A1(n5029), .A2(n5320), .ZN(n5567) );
  NAND2_X1 U6206 ( .A1(n6628), .A2(n6038), .ZN(n5031) );
  INV_X1 U6207 ( .A(n5216), .ZN(n5230) );
  AOI21_X1 U6208 ( .B1(n5031), .B2(n5230), .A(n5030), .ZN(n5899) );
  NAND2_X1 U6209 ( .A1(n5032), .A2(n5034), .ZN(n5707) );
  INV_X1 U6210 ( .A(n5707), .ZN(n5033) );
  AOI211_X1 U6211 ( .C1(n5231), .C2(n5034), .A(n5899), .B(n5033), .ZN(n5035)
         );
  AOI211_X1 U6212 ( .C1(n6651), .C2(n5567), .A(n5036), .B(n5035), .ZN(n5037)
         );
  OAI21_X1 U6213 ( .B1(n5038), .B2(n6638), .A(n5037), .ZN(U2994) );
  INV_X1 U6214 ( .A(n5041), .ZN(n5042) );
  NAND2_X1 U6215 ( .A1(n5042), .A2(n5182), .ZN(n6738) );
  NAND2_X1 U6216 ( .A1(n6738), .A2(n5043), .ZN(n5044) );
  NAND2_X1 U6217 ( .A1(n5198), .A2(EBX_REG_31__SCAN_IN), .ZN(n5045) );
  NOR2_X1 U6218 ( .A1(n3764), .A2(n5045), .ZN(n5046) );
  INV_X1 U6219 ( .A(n5049), .ZN(n5047) );
  INV_X1 U6220 ( .A(n5048), .ZN(n5054) );
  OAI21_X1 U6221 ( .B1(n5051), .B2(n5050), .A(n5049), .ZN(n5052) );
  INV_X1 U6222 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5701) );
  INV_X1 U6223 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5158) );
  XNOR2_X1 U6224 ( .A(n5185), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5666)
         );
  AOI22_X1 U6225 ( .A1(n5121), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n5107), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5064) );
  AOI22_X1 U6226 ( .A1(n3496), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n5123), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n5063) );
  AOI22_X1 U6227 ( .A1(n5124), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3486), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5062) );
  AOI22_X1 U6228 ( .A1(n3462), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3490), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5061) );
  NAND4_X1 U6229 ( .A1(n5064), .A2(n5063), .A3(n5062), .A4(n5061), .ZN(n5070)
         );
  AOI22_X1 U6230 ( .A1(n5122), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3468), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5068) );
  AOI22_X1 U6231 ( .A1(n3086), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5067) );
  AOI22_X1 U6232 ( .A1(n5115), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5114), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5066) );
  AOI22_X1 U6233 ( .A1(n5116), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3089), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5065) );
  NAND4_X1 U6234 ( .A1(n5068), .A2(n5067), .A3(n5066), .A4(n5065), .ZN(n5069)
         );
  NOR2_X1 U6235 ( .A1(n5070), .A2(n5069), .ZN(n5175) );
  AOI22_X1 U6236 ( .A1(n5122), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n5107), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5074) );
  AOI22_X1 U6237 ( .A1(n3467), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5073) );
  AOI22_X1 U6238 ( .A1(n3086), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n5114), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5072) );
  AOI22_X1 U6239 ( .A1(n3462), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n5115), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n5071) );
  NAND4_X1 U6240 ( .A1(n5074), .A2(n5073), .A3(n5072), .A4(n5071), .ZN(n5080)
         );
  AOI22_X1 U6241 ( .A1(n5123), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n5124), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n5078) );
  AOI22_X1 U6242 ( .A1(n5116), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5077) );
  AOI22_X1 U6243 ( .A1(n5121), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3087), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5076) );
  AOI22_X1 U6244 ( .A1(n3496), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3490), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n5075) );
  NAND4_X1 U6245 ( .A1(n5078), .A2(n5077), .A3(n5076), .A4(n5075), .ZN(n5079)
         );
  NOR2_X1 U6246 ( .A1(n5080), .A2(n5079), .ZN(n5162) );
  AOI22_X1 U6247 ( .A1(n5122), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n5084) );
  AOI22_X1 U6248 ( .A1(n5123), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5083) );
  AOI22_X1 U6249 ( .A1(n5116), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5082) );
  AOI22_X1 U6250 ( .A1(n3467), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3490), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n5081) );
  NAND4_X1 U6251 ( .A1(n5084), .A2(n5083), .A3(n5082), .A4(n5081), .ZN(n5090)
         );
  AOI22_X1 U6252 ( .A1(n5121), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n5107), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5088) );
  AOI22_X1 U6253 ( .A1(n5124), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5087) );
  AOI22_X1 U6254 ( .A1(n3486), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n5114), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5086) );
  AOI22_X1 U6255 ( .A1(n3496), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n5115), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n5085) );
  NAND4_X1 U6256 ( .A1(n5088), .A2(n5087), .A3(n5086), .A4(n5085), .ZN(n5089)
         );
  NOR2_X1 U6257 ( .A1(n5090), .A2(n5089), .ZN(n5138) );
  NAND2_X1 U6258 ( .A1(n5092), .A2(n5091), .ZN(n5139) );
  NOR2_X1 U6259 ( .A1(n5138), .A2(n5139), .ZN(n5151) );
  AOI22_X1 U6260 ( .A1(n5121), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n5107), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5096) );
  AOI22_X1 U6261 ( .A1(n5116), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n5124), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n5095) );
  AOI22_X1 U6262 ( .A1(n3468), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5094) );
  AOI22_X1 U6263 ( .A1(n5122), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3089), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5093) );
  NAND4_X1 U6264 ( .A1(n5096), .A2(n5095), .A3(n5094), .A4(n5093), .ZN(n5102)
         );
  AOI22_X1 U6265 ( .A1(n3496), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5100) );
  AOI22_X1 U6266 ( .A1(n5123), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n5114), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5099) );
  AOI22_X1 U6267 ( .A1(n3462), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n5115), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n5098) );
  AOI22_X1 U6268 ( .A1(n3086), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3490), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n5097) );
  NAND4_X1 U6269 ( .A1(n5100), .A2(n5099), .A3(n5098), .A4(n5097), .ZN(n5101)
         );
  OR2_X1 U6270 ( .A1(n5102), .A2(n5101), .ZN(n5149) );
  NAND2_X1 U6271 ( .A1(n5151), .A2(n5149), .ZN(n5161) );
  NOR2_X1 U6272 ( .A1(n5162), .A2(n5161), .ZN(n5168) );
  AOI22_X1 U6273 ( .A1(n3496), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5106) );
  AOI22_X1 U6274 ( .A1(n5123), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n5114), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5105) );
  AOI22_X1 U6275 ( .A1(n3488), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5115), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n5104) );
  AOI22_X1 U6276 ( .A1(n3086), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3490), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n5103) );
  NAND4_X1 U6277 ( .A1(n5106), .A2(n5105), .A3(n5104), .A4(n5103), .ZN(n5113)
         );
  AOI22_X1 U6278 ( .A1(n5121), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n5107), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5111) );
  AOI22_X1 U6279 ( .A1(n5116), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n5124), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n5110) );
  AOI22_X1 U6280 ( .A1(n3467), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5109) );
  AOI22_X1 U6281 ( .A1(n5122), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5108) );
  NAND4_X1 U6282 ( .A1(n5111), .A2(n5110), .A3(n5109), .A4(n5108), .ZN(n5112)
         );
  OR2_X1 U6283 ( .A1(n5113), .A2(n5112), .ZN(n5167) );
  NAND2_X1 U6284 ( .A1(n5168), .A2(n5167), .ZN(n5174) );
  NOR2_X1 U6285 ( .A1(n5175), .A2(n5174), .ZN(n5132) );
  AOI22_X1 U6286 ( .A1(n5107), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5114), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5120) );
  AOI22_X1 U6287 ( .A1(n3462), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5115), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n5119) );
  AOI22_X1 U6288 ( .A1(n5116), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3087), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5118) );
  AOI22_X1 U6289 ( .A1(n3436), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3490), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5117) );
  NAND4_X1 U6290 ( .A1(n5120), .A2(n5119), .A3(n5118), .A4(n5117), .ZN(n5130)
         );
  AOI22_X1 U6291 ( .A1(n5122), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n5121), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5128) );
  AOI22_X1 U6292 ( .A1(n3496), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3467), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5127) );
  AOI22_X1 U6293 ( .A1(n5123), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n5126) );
  AOI22_X1 U6294 ( .A1(n5124), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5125) );
  NAND4_X1 U6295 ( .A1(n5128), .A2(n5127), .A3(n5126), .A4(n5125), .ZN(n5129)
         );
  NOR2_X1 U6296 ( .A1(n5130), .A2(n5129), .ZN(n5131) );
  XNOR2_X1 U6297 ( .A(n5132), .B(n5131), .ZN(n5136) );
  INV_X1 U6298 ( .A(EAX_REG_30__SCAN_IN), .ZN(n5134) );
  OAI21_X1 U6299 ( .B1(n6361), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n6673), 
        .ZN(n5133) );
  OAI21_X1 U6300 ( .B1(n3290), .B2(n5134), .A(n5133), .ZN(n5135) );
  AOI21_X1 U6301 ( .B1(n5136), .B2(n5155), .A(n5135), .ZN(n5137) );
  AOI21_X1 U6302 ( .B1(n5666), .B2(n5182), .A(n5137), .ZN(n5246) );
  XNOR2_X1 U6303 ( .A(n5139), .B(n5138), .ZN(n5141) );
  AOI22_X1 U6304 ( .A1(n4168), .A2(EAX_REG_25__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6673), .ZN(n5140) );
  OAI21_X1 U6305 ( .B1(n5141), .B2(n5177), .A(n5140), .ZN(n5146) );
  INV_X1 U6306 ( .A(n5142), .ZN(n5144) );
  INV_X1 U6307 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5143) );
  NAND2_X1 U6308 ( .A1(n5144), .A2(n5143), .ZN(n5145) );
  NAND2_X1 U6309 ( .A1(n5159), .A2(n5145), .ZN(n5716) );
  MUX2_X1 U6310 ( .A(n5146), .B(n5716), .S(n5182), .Z(n5325) );
  XNOR2_X1 U6311 ( .A(n5159), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5705)
         );
  INV_X1 U6312 ( .A(n5149), .ZN(n5150) );
  XNOR2_X1 U6313 ( .A(n5151), .B(n5150), .ZN(n5156) );
  INV_X1 U6314 ( .A(EAX_REG_26__SCAN_IN), .ZN(n5153) );
  OAI21_X1 U6315 ( .B1(n6361), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n6673), 
        .ZN(n5152) );
  OAI21_X1 U6316 ( .B1(n3290), .B2(n5153), .A(n5152), .ZN(n5154) );
  AOI21_X1 U6317 ( .B1(n5156), .B2(n5155), .A(n5154), .ZN(n5157) );
  AOI21_X1 U6318 ( .B1(n5705), .B2(n5182), .A(n5157), .ZN(n5309) );
  OAI21_X1 U6319 ( .B1(n5159), .B2(n5701), .A(n5158), .ZN(n5160) );
  NAND2_X1 U6320 ( .A1(n5160), .A2(n5171), .ZN(n5689) );
  XNOR2_X1 U6321 ( .A(n5162), .B(n5161), .ZN(n5164) );
  AOI22_X1 U6322 ( .A1(n4168), .A2(EAX_REG_27__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6673), .ZN(n5163) );
  OAI21_X1 U6323 ( .B1(n5164), .B2(n5177), .A(n5163), .ZN(n5166) );
  MUX2_X1 U6324 ( .A(n5689), .B(n5166), .S(n5165), .Z(n5296) );
  XNOR2_X1 U6325 ( .A(n5168), .B(n5167), .ZN(n5170) );
  AOI22_X1 U6326 ( .A1(n4168), .A2(EAX_REG_28__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6673), .ZN(n5169) );
  OAI21_X1 U6327 ( .B1(n5170), .B2(n5177), .A(n5169), .ZN(n5173) );
  INV_X1 U6328 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n6861) );
  NAND2_X1 U6329 ( .A1(n5171), .A2(n6861), .ZN(n5172) );
  NAND2_X1 U6330 ( .A1(n5180), .A2(n5172), .ZN(n5684) );
  MUX2_X1 U6331 ( .A(n5173), .B(n5684), .S(n5182), .Z(n5282) );
  XNOR2_X1 U6332 ( .A(n5175), .B(n5174), .ZN(n5178) );
  AOI22_X1 U6333 ( .A1(n4168), .A2(EAX_REG_29__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6673), .ZN(n5176) );
  OAI21_X1 U6334 ( .B1(n5178), .B2(n5177), .A(n5176), .ZN(n5183) );
  INV_X1 U6335 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5179) );
  NAND2_X1 U6336 ( .A1(n5180), .A2(n5179), .ZN(n5181) );
  NAND2_X1 U6337 ( .A1(n5185), .A2(n5181), .ZN(n5677) );
  MUX2_X1 U6338 ( .A(n5183), .B(n5677), .S(n5182), .Z(n5184) );
  XOR2_X1 U6339 ( .A(n5246), .B(n5273), .Z(n5671) );
  INV_X1 U6340 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5669) );
  INV_X1 U6341 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5258) );
  NAND2_X1 U6342 ( .A1(n6423), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5187) );
  NAND2_X1 U6343 ( .A1(n5671), .A2(n6422), .ZN(n5215) );
  INV_X1 U6344 ( .A(n5187), .ZN(n5188) );
  AND2_X1 U6345 ( .A1(n5200), .A2(n6361), .ZN(n6799) );
  AND2_X1 U6346 ( .A1(n5189), .A2(n6799), .ZN(n5190) );
  NAND2_X1 U6347 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5194) );
  INV_X1 U6348 ( .A(n6423), .ZN(n6458) );
  NOR2_X1 U6349 ( .A1(n6459), .A2(n6458), .ZN(n5556) );
  NAND3_X1 U6350 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .ZN(n5208) );
  NAND3_X1 U6351 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .ZN(n5191) );
  INV_X1 U6352 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6750) );
  NAND3_X1 U6353 ( .A1(REIP_REG_3__SCAN_IN), .A2(REIP_REG_1__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5518) );
  NOR3_X1 U6354 ( .A1(n6750), .A2(n6748), .A3(n5518), .ZN(n6430) );
  NAND2_X1 U6355 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6430), .ZN(n6417) );
  NOR2_X1 U6356 ( .A1(n6753), .A2(n6417), .ZN(n6407) );
  NAND2_X1 U6357 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6407), .ZN(n5205) );
  NAND4_X1 U6358 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .A3(
        REIP_REG_19__SCAN_IN), .A4(n5399), .ZN(n5355) );
  NAND3_X1 U6359 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n5210) );
  NOR2_X1 U6360 ( .A1(n5355), .A2(n5210), .ZN(n5192) );
  AND2_X1 U6361 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5311) );
  NAND2_X1 U6362 ( .A1(n5311), .A2(REIP_REG_26__SCAN_IN), .ZN(n5211) );
  NAND2_X1 U6363 ( .A1(n6459), .A2(n5211), .ZN(n5193) );
  AOI21_X1 U6364 ( .B1(n6459), .B2(n6952), .A(n5195), .ZN(n5255) );
  AND2_X1 U6365 ( .A1(n5197), .A2(n5196), .ZN(n5256) );
  INV_X1 U6366 ( .A(n5256), .ZN(n5202) );
  NAND3_X1 U6367 ( .A1(n5200), .A2(n5199), .A3(n5198), .ZN(n5201) );
  NAND2_X1 U6368 ( .A1(n5202), .A2(n5201), .ZN(n5203) );
  AOI22_X1 U6369 ( .A1(n6441), .A2(EBX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6452), .ZN(n5204) );
  OAI21_X1 U6370 ( .B1(n5255), .B2(n5259), .A(n5204), .ZN(n5213) );
  INV_X1 U6371 ( .A(n5205), .ZN(n5206) );
  AND3_X1 U6372 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_11__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .ZN(n5207) );
  NAND2_X1 U6373 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .ZN(
        n5498) );
  NAND2_X1 U6374 ( .A1(REIP_REG_18__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .ZN(
        n5209) );
  NAND3_X1 U6375 ( .A1(n3101), .A2(REIP_REG_27__SCAN_IN), .A3(
        REIP_REG_28__SCAN_IN), .ZN(n5279) );
  NOR3_X1 U6376 ( .A1(n5279), .A2(REIP_REG_30__SCAN_IN), .A3(n6952), .ZN(n5212) );
  AOI211_X1 U6377 ( .C1(n5666), .C2(n6427), .A(n5213), .B(n5212), .ZN(n5214)
         );
  OAI211_X1 U6378 ( .C1(n6440), .C2(n5270), .A(n5215), .B(n5214), .ZN(U2797)
         );
  NAND3_X1 U6379 ( .A1(n5217), .A2(n5925), .A3(n5216), .ZN(n5710) );
  INV_X1 U6380 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5219) );
  INV_X1 U6381 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5218) );
  NAND2_X1 U6382 ( .A1(n5219), .A2(n5218), .ZN(n5910) );
  NAND2_X1 U6383 ( .A1(n5935), .A2(n5738), .ZN(n5924) );
  NOR4_X1 U6384 ( .A1(n5910), .A2(n5707), .A3(n5924), .A4(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5220) );
  MUX2_X1 U6385 ( .A(n5220), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .S(n5824), 
        .Z(n5221) );
  NAND2_X1 U6386 ( .A1(n5824), .A2(n7061), .ZN(n5223) );
  NOR2_X1 U6387 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5235) );
  INV_X1 U6388 ( .A(n5235), .ZN(n5222) );
  NOR3_X2 U6389 ( .A1(n5699), .A2(n5697), .A3(n5222), .ZN(n5674) );
  INV_X1 U6390 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5864) );
  AND2_X1 U6391 ( .A1(n5824), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5698)
         );
  NAND3_X1 U6392 ( .A1(n5698), .A2(n3115), .A3(n5223), .ZN(n5224) );
  AND2_X1 U6393 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5682) );
  XOR2_X1 U6394 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .B(n5225), .Z(n5673) );
  INV_X1 U6395 ( .A(n5967), .ZN(n6044) );
  AND2_X1 U6396 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5232) );
  INV_X1 U6397 ( .A(n5232), .ZN(n5894) );
  NAND2_X1 U6398 ( .A1(n5967), .A2(n5894), .ZN(n5226) );
  INV_X1 U6399 ( .A(n5682), .ZN(n5227) );
  NAND2_X1 U6400 ( .A1(n5967), .A2(n5227), .ZN(n5228) );
  OAI21_X1 U6401 ( .B1(n6044), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5861), 
        .ZN(n5237) );
  NAND2_X1 U6402 ( .A1(n6577), .A2(REIP_REG_30__SCAN_IN), .ZN(n5667) );
  INV_X1 U6403 ( .A(n5667), .ZN(n5229) );
  AND2_X2 U6404 ( .A1(n5871), .A2(n5682), .ZN(n5865) );
  INV_X1 U6405 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5238) );
  NAND3_X1 U6406 ( .A1(n5865), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5238), .ZN(n5233) );
  OAI211_X1 U6407 ( .C1(n5673), .C2(n6638), .A(n5234), .B(n5233), .ZN(U2988)
         );
  AOI21_X1 U6408 ( .B1(n5967), .B2(n5238), .A(n5237), .ZN(n5241) );
  NAND4_X1 U6409 ( .A1(n5865), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n5240), .ZN(n5239) );
  NAND2_X1 U6410 ( .A1(n6577), .A2(REIP_REG_31__SCAN_IN), .ZN(n5250) );
  OAI211_X1 U6411 ( .C1(n5241), .C2(n5240), .A(n5239), .B(n5250), .ZN(n5242)
         );
  AOI21_X1 U6412 ( .B1(n5243), .B2(n6651), .A(n5242), .ZN(n5244) );
  OAI21_X1 U6413 ( .B1(n5254), .B2(n6638), .A(n5244), .ZN(U2987) );
  AOI22_X1 U6414 ( .A1(n4168), .A2(EAX_REG_31__SCAN_IN), .B1(n5245), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5248) );
  NAND2_X1 U6415 ( .A1(n5273), .A2(n5246), .ZN(n5247) );
  XOR2_X1 U6416 ( .A(n5248), .B(n5247), .Z(n5267) );
  NAND2_X1 U6417 ( .A1(n6591), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5249)
         );
  OAI211_X1 U6418 ( .C1(n5251), .C2(n6599), .A(n5250), .B(n5249), .ZN(n5252)
         );
  OAI21_X1 U6419 ( .B1(n5254), .B2(n6362), .A(n5253), .ZN(U2955) );
  NAND2_X1 U6420 ( .A1(n5267), .A2(n6422), .ZN(n5264) );
  INV_X1 U6421 ( .A(n6459), .ZN(n6424) );
  OAI21_X1 U6422 ( .B1(REIP_REG_30__SCAN_IN), .B2(n6424), .A(n5255), .ZN(n5262) );
  NAND3_X1 U6423 ( .A1(n5517), .A2(EBX_REG_31__SCAN_IN), .A3(n5256), .ZN(n5257) );
  OAI21_X1 U6424 ( .B1(n6444), .B2(n5258), .A(n5257), .ZN(n5261) );
  NOR4_X1 U6425 ( .A1(n5279), .A2(REIP_REG_31__SCAN_IN), .A3(n5259), .A4(n6952), .ZN(n5260) );
  AOI211_X1 U6426 ( .C1(REIP_REG_31__SCAN_IN), .C2(n5262), .A(n5261), .B(n5260), .ZN(n5263) );
  OAI211_X1 U6427 ( .C1(n5265), .C2(n6440), .A(n5264), .B(n5263), .ZN(U2796)
         );
  NAND3_X1 U6428 ( .A1(n5267), .A2(n5266), .A3(n5664), .ZN(n5269) );
  AOI22_X1 U6429 ( .A1(n5645), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n5658), .ZN(n5268) );
  NAND2_X1 U6430 ( .A1(n5269), .A2(n5268), .ZN(U2860) );
  INV_X1 U6431 ( .A(n5671), .ZN(n5610) );
  INV_X1 U6432 ( .A(EBX_REG_30__SCAN_IN), .ZN(n6910) );
  OAI222_X1 U6433 ( .A1(n5599), .A2(n5610), .B1(n6910), .B2(n6480), .C1(n5270), 
        .C2(n5605), .ZN(U2829) );
  OR2_X1 U6434 ( .A1(n5400), .A2(READREQUEST_REG_SCAN_IN), .ZN(n5272) );
  INV_X1 U6435 ( .A(n6797), .ZN(n5271) );
  MUX2_X1 U6436 ( .A(n5272), .B(n5271), .S(n6808), .Z(U3474) );
  MUX2_X1 U6437 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6780), .Z(U3473) );
  AOI21_X1 U6438 ( .B1(n5274), .B2(n5281), .A(n5273), .ZN(n5679) );
  INV_X1 U6439 ( .A(n5679), .ZN(n5613) );
  INV_X1 U6440 ( .A(n5275), .ZN(n5276) );
  AND2_X1 U6441 ( .A1(n5286), .A2(n5276), .ZN(n5277) );
  AOI22_X1 U6442 ( .A1(n6441), .A2(EBX_REG_29__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6452), .ZN(n5280) );
  OAI21_X1 U6443 ( .B1(n5294), .B2(n5282), .A(n5281), .ZN(n5688) );
  NAND2_X1 U6444 ( .A1(n5306), .A2(n5299), .ZN(n5285) );
  INV_X1 U6445 ( .A(n5283), .ZN(n5284) );
  NAND2_X1 U6446 ( .A1(n5285), .A2(n5284), .ZN(n5287) );
  NAND2_X1 U6447 ( .A1(n5287), .A2(n5286), .ZN(n5563) );
  INV_X1 U6448 ( .A(n5563), .ZN(n5873) );
  NAND2_X1 U6449 ( .A1(n3101), .A2(REIP_REG_27__SCAN_IN), .ZN(n5289) );
  MUX2_X1 U6450 ( .A(n5289), .B(n5288), .S(REIP_REG_28__SCAN_IN), .Z(n5291) );
  AOI22_X1 U6451 ( .A1(n6441), .A2(EBX_REG_28__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6452), .ZN(n5290) );
  OAI211_X1 U6452 ( .C1(n6462), .C2(n5684), .A(n5291), .B(n5290), .ZN(n5292)
         );
  AOI21_X1 U6453 ( .B1(n5873), .B2(n6451), .A(n5292), .ZN(n5293) );
  OAI21_X1 U6454 ( .B1(n5688), .B2(n6435), .A(n5293), .ZN(U2799) );
  INV_X1 U6455 ( .A(n5294), .ZN(n5295) );
  OAI21_X1 U6456 ( .B1(n5307), .B2(n5296), .A(n5295), .ZN(n5696) );
  AOI22_X1 U6457 ( .A1(n6441), .A2(EBX_REG_27__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6452), .ZN(n5298) );
  NAND2_X1 U6458 ( .A1(n5312), .A2(REIP_REG_27__SCAN_IN), .ZN(n5297) );
  OAI211_X1 U6459 ( .C1(n6462), .C2(n5689), .A(n5298), .B(n5297), .ZN(n5301)
         );
  XNOR2_X1 U6460 ( .A(n5306), .B(n5299), .ZN(n5882) );
  NOR2_X1 U6461 ( .A1(n5882), .A2(n6440), .ZN(n5300) );
  AOI211_X1 U6462 ( .C1(n3101), .C2(n6779), .A(n5301), .B(n5300), .ZN(n5302)
         );
  OAI21_X1 U6463 ( .B1(n5696), .B2(n6435), .A(n5302), .ZN(U2800) );
  NOR2_X1 U6464 ( .A1(n5303), .A2(n5304), .ZN(n5305) );
  OR2_X1 U6465 ( .A1(n5306), .A2(n5305), .ZN(n5889) );
  OAI21_X1 U6466 ( .B1(n5309), .B2(n5323), .A(n5308), .ZN(n5702) );
  INV_X1 U6467 ( .A(n5702), .ZN(n5310) );
  NAND2_X1 U6468 ( .A1(n5310), .A2(n6422), .ZN(n5318) );
  OAI22_X1 U6469 ( .A1(n6467), .A2(n7040), .B1(n5701), .B2(n6444), .ZN(n5316)
         );
  AOI21_X1 U6470 ( .B1(n3217), .B2(n5311), .A(REIP_REG_26__SCAN_IN), .ZN(n5314) );
  INV_X1 U6471 ( .A(n5312), .ZN(n5313) );
  NOR2_X1 U6472 ( .A1(n5314), .A2(n5313), .ZN(n5315) );
  AOI211_X1 U6473 ( .C1(n3090), .C2(n5705), .A(n5316), .B(n5315), .ZN(n5317)
         );
  OAI211_X1 U6474 ( .C1(n6440), .C2(n5889), .A(n5318), .B(n5317), .ZN(U2801)
         );
  INV_X1 U6475 ( .A(n5303), .ZN(n5322) );
  NAND2_X1 U6476 ( .A1(n5320), .A2(n5319), .ZN(n5321) );
  NAND2_X1 U6477 ( .A1(n5322), .A2(n5321), .ZN(n5900) );
  INV_X1 U6478 ( .A(n5323), .ZN(n5324) );
  OAI21_X1 U6479 ( .B1(n5326), .B2(n5325), .A(n5324), .ZN(n5622) );
  INV_X1 U6480 ( .A(n5622), .ZN(n5718) );
  NAND2_X1 U6481 ( .A1(n5718), .A2(n6422), .ZN(n5333) );
  XOR2_X1 U6482 ( .A(REIP_REG_24__SCAN_IN), .B(REIP_REG_25__SCAN_IN), .Z(n5331) );
  INV_X1 U6483 ( .A(REIP_REG_25__SCAN_IN), .ZN(n5328) );
  AOI22_X1 U6484 ( .A1(n6441), .A2(EBX_REG_25__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6452), .ZN(n5327) );
  OAI21_X1 U6485 ( .B1(n5341), .B2(n5328), .A(n5327), .ZN(n5330) );
  NOR2_X1 U6486 ( .A1(n6462), .A2(n5716), .ZN(n5329) );
  AOI211_X1 U6487 ( .C1(n3217), .C2(n5331), .A(n5330), .B(n5329), .ZN(n5332)
         );
  OAI211_X1 U6488 ( .C1(n5900), .C2(n6440), .A(n5333), .B(n5332), .ZN(U2802)
         );
  NAND2_X1 U6489 ( .A1(n5567), .A2(n6451), .ZN(n5337) );
  AOI22_X1 U6490 ( .A1(n6441), .A2(EBX_REG_24__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n6452), .ZN(n5334) );
  OAI21_X1 U6491 ( .B1(n5341), .B2(n6773), .A(n5334), .ZN(n5335) );
  AOI21_X1 U6492 ( .B1(n3217), .B2(n6773), .A(n5335), .ZN(n5336) );
  OAI211_X1 U6493 ( .C1(n6462), .C2(n5338), .A(n5337), .B(n5336), .ZN(n5339)
         );
  AOI21_X1 U6494 ( .B1(n5566), .B2(n6422), .A(n5339), .ZN(n5340) );
  INV_X1 U6495 ( .A(n5340), .ZN(U2803) );
  NOR3_X1 U6496 ( .A1(n5369), .A2(n5723), .A3(n5732), .ZN(n5343) );
  INV_X1 U6497 ( .A(n5341), .ZN(n5342) );
  OAI21_X1 U6498 ( .B1(n5343), .B2(REIP_REG_23__SCAN_IN), .A(n5342), .ZN(n5345) );
  AOI22_X1 U6499 ( .A1(n6441), .A2(EBX_REG_23__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n6452), .ZN(n5344) );
  OAI211_X1 U6500 ( .C1(n6462), .C2(n5346), .A(n5345), .B(n5344), .ZN(n5347)
         );
  AOI21_X1 U6501 ( .B1(n5569), .B2(n6451), .A(n5347), .ZN(n5348) );
  OAI21_X1 U6502 ( .B1(n5628), .B2(n6435), .A(n5348), .ZN(U2804) );
  OAI21_X1 U6503 ( .B1(n5370), .B2(n5350), .A(n5349), .ZN(n5907) );
  INV_X1 U6504 ( .A(n5351), .ZN(n5354) );
  INV_X1 U6505 ( .A(n5352), .ZN(n5365) );
  AOI21_X1 U6506 ( .B1(n5354), .B2(n5365), .A(n5353), .ZN(n5727) );
  NAND2_X1 U6507 ( .A1(n5727), .A2(n6422), .ZN(n5363) );
  INV_X1 U6508 ( .A(n5369), .ZN(n5361) );
  XOR2_X1 U6509 ( .A(REIP_REG_22__SCAN_IN), .B(REIP_REG_21__SCAN_IN), .Z(n5360) );
  INV_X1 U6510 ( .A(n5355), .ZN(n5356) );
  OR2_X1 U6511 ( .A1(n5556), .A2(n5356), .ZN(n5366) );
  AOI22_X1 U6512 ( .A1(n6441), .A2(EBX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6452), .ZN(n5357) );
  OAI21_X1 U6513 ( .B1(n5366), .B2(n5723), .A(n5357), .ZN(n5359) );
  NOR2_X1 U6514 ( .A1(n6462), .A2(n5725), .ZN(n5358) );
  AOI211_X1 U6515 ( .C1(n5361), .C2(n5360), .A(n5359), .B(n5358), .ZN(n5362)
         );
  OAI211_X1 U6516 ( .C1(n6440), .C2(n5907), .A(n5363), .B(n5362), .ZN(U2805)
         );
  OAI21_X1 U6517 ( .B1(n3117), .B2(n3232), .A(n5365), .ZN(n5737) );
  AOI22_X1 U6518 ( .A1(n6441), .A2(EBX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6452), .ZN(n5368) );
  INV_X1 U6519 ( .A(n5366), .ZN(n5383) );
  NAND2_X1 U6520 ( .A1(n5383), .A2(REIP_REG_21__SCAN_IN), .ZN(n5367) );
  OAI211_X1 U6521 ( .C1(n5369), .C2(REIP_REG_21__SCAN_IN), .A(n5368), .B(n5367), .ZN(n5375) );
  INV_X1 U6522 ( .A(n5370), .ZN(n5371) );
  OAI21_X1 U6523 ( .B1(n5373), .B2(n5372), .A(n5371), .ZN(n5917) );
  NOR2_X1 U6524 ( .A1(n5917), .A2(n6440), .ZN(n5374) );
  AOI211_X1 U6525 ( .C1(n3090), .C2(n5734), .A(n5375), .B(n5374), .ZN(n5376)
         );
  OAI21_X1 U6526 ( .B1(n5737), .B2(n6435), .A(n5376), .ZN(U2806) );
  NAND2_X1 U6527 ( .A1(n3085), .A2(n5378), .ZN(n5397) );
  AOI21_X1 U6528 ( .B1(n5379), .B2(n5397), .A(n3117), .ZN(n5744) );
  INV_X1 U6529 ( .A(n5744), .ZN(n5636) );
  XNOR2_X1 U6530 ( .A(n5382), .B(n5381), .ZN(n5931) );
  AOI22_X1 U6531 ( .A1(n6441), .A2(EBX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6452), .ZN(n5386) );
  OAI21_X1 U6532 ( .B1(n5384), .B2(REIP_REG_20__SCAN_IN), .A(n5383), .ZN(n5385) );
  OAI211_X1 U6533 ( .C1(n6462), .C2(n5742), .A(n5386), .B(n5385), .ZN(n5387)
         );
  AOI21_X1 U6534 ( .B1(n5931), .B2(n6451), .A(n5387), .ZN(n5388) );
  OAI21_X1 U6535 ( .B1(n5636), .B2(n6435), .A(n5388), .ZN(U2807) );
  INV_X1 U6536 ( .A(n5428), .ZN(n5393) );
  MUX2_X1 U6537 ( .A(n5391), .B(n5390), .S(n5389), .Z(n5413) );
  INV_X1 U6538 ( .A(n5413), .ZN(n5392) );
  NAND2_X1 U6539 ( .A1(n5393), .A2(n5392), .ZN(n5415) );
  XNOR2_X1 U6540 ( .A(n5415), .B(n5394), .ZN(n5939) );
  AND2_X1 U6541 ( .A1(n3085), .A2(n5395), .ZN(n5411) );
  OR2_X1 U6542 ( .A1(n5411), .A2(n5396), .ZN(n5398) );
  NAND2_X1 U6543 ( .A1(n5754), .A2(n6422), .ZN(n5409) );
  INV_X1 U6544 ( .A(n5752), .ZN(n5407) );
  INV_X1 U6545 ( .A(REIP_REG_19__SCAN_IN), .ZN(n5403) );
  OR2_X1 U6546 ( .A1(n5556), .A2(n5399), .ZN(n5430) );
  NAND2_X1 U6547 ( .A1(n6423), .A2(n5400), .ZN(n6442) );
  INV_X1 U6548 ( .A(n6442), .ZN(n6429) );
  INV_X1 U6549 ( .A(EBX_REG_19__SCAN_IN), .ZN(n6912) );
  NOR2_X1 U6550 ( .A1(n6467), .A2(n6912), .ZN(n5401) );
  AOI211_X1 U6551 ( .C1(n6452), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n6429), 
        .B(n5401), .ZN(n5402) );
  OAI21_X1 U6552 ( .B1(n5403), .B2(n5430), .A(n5402), .ZN(n5406) );
  XNOR2_X1 U6553 ( .A(REIP_REG_18__SCAN_IN), .B(REIP_REG_19__SCAN_IN), .ZN(
        n5404) );
  NOR2_X1 U6554 ( .A1(n5420), .A2(n5404), .ZN(n5405) );
  AOI211_X1 U6555 ( .C1(n6427), .C2(n5407), .A(n5406), .B(n5405), .ZN(n5408)
         );
  OAI211_X1 U6556 ( .C1(n5939), .C2(n6440), .A(n5409), .B(n5408), .ZN(U2808)
         );
  NAND2_X1 U6557 ( .A1(n3085), .A2(n5410), .ZN(n5424) );
  AOI21_X1 U6558 ( .B1(n5412), .B2(n5424), .A(n5411), .ZN(n5762) );
  INV_X1 U6559 ( .A(n5762), .ZN(n5642) );
  NAND2_X1 U6560 ( .A1(n5428), .A2(n5413), .ZN(n5414) );
  AND2_X1 U6561 ( .A1(n5415), .A2(n5414), .ZN(n5947) );
  NAND2_X1 U6562 ( .A1(n6427), .A2(n5758), .ZN(n5419) );
  OAI21_X1 U6563 ( .B1(n6444), .B2(n5760), .A(n6442), .ZN(n5417) );
  INV_X1 U6564 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6862) );
  NOR2_X1 U6565 ( .A1(n5430), .A2(n6862), .ZN(n5416) );
  AOI211_X1 U6566 ( .C1(EBX_REG_18__SCAN_IN), .C2(n6441), .A(n5417), .B(n5416), 
        .ZN(n5418) );
  OAI211_X1 U6567 ( .C1(REIP_REG_18__SCAN_IN), .C2(n5420), .A(n5419), .B(n5418), .ZN(n5421) );
  AOI21_X1 U6568 ( .B1(n5947), .B2(n6451), .A(n5421), .ZN(n5422) );
  OAI21_X1 U6569 ( .B1(n5642), .B2(n6435), .A(n5422), .ZN(U2809) );
  NAND2_X1 U6570 ( .A1(n3085), .A2(n5423), .ZN(n5441) );
  INV_X1 U6571 ( .A(n5441), .ZN(n5426) );
  OAI21_X1 U6572 ( .B1(n5426), .B2(n5425), .A(n5424), .ZN(n5774) );
  OAI21_X1 U6573 ( .B1(n5461), .B2(n5442), .A(n5427), .ZN(n5429) );
  NAND2_X1 U6574 ( .A1(n5429), .A2(n5428), .ZN(n5956) );
  NOR2_X1 U6575 ( .A1(n5956), .A2(n6440), .ZN(n5436) );
  AND2_X1 U6576 ( .A1(n3090), .A2(n5771), .ZN(n5435) );
  INV_X1 U6577 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5777) );
  INV_X1 U6578 ( .A(REIP_REG_15__SCAN_IN), .ZN(n5787) );
  OR3_X1 U6579 ( .A1(n5448), .A2(n5777), .A3(n5787), .ZN(n5431) );
  INV_X1 U6580 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6766) );
  AOI21_X1 U6581 ( .B1(n5431), .B2(n6766), .A(n5430), .ZN(n5434) );
  NAND2_X1 U6582 ( .A1(n6441), .A2(EBX_REG_17__SCAN_IN), .ZN(n5432) );
  OAI211_X1 U6583 ( .C1(n6444), .C2(n5769), .A(n5432), .B(n6442), .ZN(n5433)
         );
  NOR4_X1 U6584 ( .A1(n5436), .A2(n5435), .A3(n5434), .A4(n5433), .ZN(n5437)
         );
  OAI21_X1 U6585 ( .B1(n5774), .B2(n6435), .A(n5437), .ZN(U2810) );
  NAND2_X1 U6586 ( .A1(n3085), .A2(n5438), .ZN(n5455) );
  NAND2_X1 U6587 ( .A1(n5455), .A2(n5439), .ZN(n5440) );
  XOR2_X1 U6588 ( .A(n5442), .B(n5461), .Z(n5966) );
  OAI21_X1 U6589 ( .B1(n6444), .B2(n5778), .A(n6442), .ZN(n5444) );
  NOR3_X1 U6590 ( .A1(n5448), .A2(REIP_REG_16__SCAN_IN), .A3(n5787), .ZN(n5443) );
  AOI211_X1 U6591 ( .C1(EBX_REG_16__SCAN_IN), .C2(n6441), .A(n5444), .B(n5443), 
        .ZN(n5445) );
  OAI21_X1 U6592 ( .B1(n5781), .B2(n6462), .A(n5445), .ZN(n5446) );
  AOI21_X1 U6593 ( .B1(n6451), .B2(n5966), .A(n5446), .ZN(n5450) );
  INV_X1 U6594 ( .A(n5556), .ZN(n6387) );
  NAND2_X1 U6595 ( .A1(n5447), .A2(n6387), .ZN(n5470) );
  INV_X1 U6596 ( .A(n5470), .ZN(n5484) );
  NOR2_X1 U6597 ( .A1(n5448), .A2(REIP_REG_15__SCAN_IN), .ZN(n5463) );
  OAI21_X1 U6598 ( .B1(n5484), .B2(n5463), .A(REIP_REG_16__SCAN_IN), .ZN(n5449) );
  OAI211_X1 U6599 ( .C1(n5649), .C2(n6435), .A(n5450), .B(n5449), .ZN(U2811)
         );
  INV_X1 U6600 ( .A(n5490), .ZN(n5453) );
  OAI21_X1 U6601 ( .B1(n5487), .B2(n5473), .A(n5472), .ZN(n5471) );
  INV_X1 U6602 ( .A(n5455), .ZN(n5456) );
  AOI21_X1 U6603 ( .B1(n5471), .B2(n5457), .A(n5456), .ZN(n5791) );
  NAND2_X1 U6604 ( .A1(n5791), .A2(n6422), .ZN(n5469) );
  INV_X1 U6605 ( .A(n5789), .ZN(n5467) );
  AND2_X1 U6606 ( .A1(n5458), .A2(n5478), .ZN(n5480) );
  OR2_X1 U6607 ( .A1(n5480), .A2(n5459), .ZN(n5460) );
  NAND2_X1 U6608 ( .A1(n5461), .A2(n5460), .ZN(n5974) );
  OAI21_X1 U6609 ( .B1(n6444), .B2(n5462), .A(n6442), .ZN(n5464) );
  AOI211_X1 U6610 ( .C1(EBX_REG_15__SCAN_IN), .C2(n6441), .A(n5464), .B(n5463), 
        .ZN(n5465) );
  OAI21_X1 U6611 ( .B1(n6440), .B2(n5974), .A(n5465), .ZN(n5466) );
  AOI21_X1 U6612 ( .B1(n5467), .B2(n3090), .A(n5466), .ZN(n5468) );
  OAI211_X1 U6613 ( .C1(n5787), .C2(n5470), .A(n5469), .B(n5468), .ZN(U2812)
         );
  INV_X1 U6614 ( .A(n5471), .ZN(n5475) );
  NOR3_X1 U6615 ( .A1(n5487), .A2(n5473), .A3(n5472), .ZN(n5474) );
  NOR2_X1 U6616 ( .A1(n5475), .A2(n5474), .ZN(n5798) );
  INV_X1 U6617 ( .A(n5798), .ZN(n5653) );
  INV_X1 U6618 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6763) );
  AOI21_X1 U6619 ( .B1(n5476), .B2(n6763), .A(n6429), .ZN(n5477) );
  OAI21_X1 U6620 ( .B1(n6462), .B2(n5796), .A(n5477), .ZN(n5483) );
  NOR2_X1 U6621 ( .A1(n5458), .A2(n5478), .ZN(n5479) );
  OR2_X1 U6622 ( .A1(n5480), .A2(n5479), .ZN(n5982) );
  AOI22_X1 U6623 ( .A1(EBX_REG_14__SCAN_IN), .A2(n6441), .B1(
        PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n6452), .ZN(n5481) );
  OAI21_X1 U6624 ( .B1(n6440), .B2(n5982), .A(n5481), .ZN(n5482) );
  AOI211_X1 U6625 ( .C1(n5484), .C2(REIP_REG_14__SCAN_IN), .A(n5483), .B(n5482), .ZN(n5485) );
  OAI21_X1 U6626 ( .B1(n5653), .B2(n6435), .A(n5485), .ZN(U2813) );
  INV_X1 U6627 ( .A(n5486), .ZN(n5489) );
  INV_X1 U6628 ( .A(n5487), .ZN(n5488) );
  NOR2_X1 U6629 ( .A1(n5556), .A2(n5491), .ZN(n6377) );
  AOI21_X1 U6630 ( .B1(n5493), .B2(n5492), .A(n5458), .ZN(n6010) );
  INV_X1 U6631 ( .A(n6010), .ZN(n5581) );
  AOI22_X1 U6632 ( .A1(EBX_REG_13__SCAN_IN), .A2(n6441), .B1(
        PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n6452), .ZN(n5494) );
  OAI21_X1 U6633 ( .B1(n6440), .B2(n5581), .A(n5494), .ZN(n5496) );
  OAI21_X1 U6634 ( .B1(n6462), .B2(n5804), .A(n6442), .ZN(n5495) );
  AOI211_X1 U6635 ( .C1(n6377), .C2(REIP_REG_13__SCAN_IN), .A(n5496), .B(n5495), .ZN(n5501) );
  INV_X1 U6636 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6761) );
  INV_X1 U6637 ( .A(REIP_REG_12__SCAN_IN), .ZN(n5497) );
  AOI21_X1 U6638 ( .B1(n6761), .B2(n5497), .A(n6384), .ZN(n5499) );
  NAND2_X1 U6639 ( .A1(n5499), .A2(n5498), .ZN(n5500) );
  OAI211_X1 U6640 ( .C1(n5802), .C2(n6435), .A(n5501), .B(n5500), .ZN(U2814)
         );
  NAND2_X1 U6641 ( .A1(n3085), .A2(n5594), .ZN(n5593) );
  OR2_X1 U6642 ( .A1(n5593), .A2(n5584), .ZN(n5586) );
  NOR2_X1 U6643 ( .A1(n5593), .A2(n5502), .ZN(n5655) );
  AOI21_X1 U6644 ( .B1(n5503), .B2(n5586), .A(n5655), .ZN(n5830) );
  INV_X1 U6645 ( .A(n5830), .ZN(n5661) );
  INV_X1 U6646 ( .A(n6389), .ZN(n5505) );
  NAND2_X1 U6647 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n5504) );
  INV_X1 U6648 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6997) );
  OAI21_X1 U6649 ( .B1(n5505), .B2(n5504), .A(n6997), .ZN(n5512) );
  INV_X1 U6650 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5508) );
  OR2_X1 U6651 ( .A1(n5589), .A2(n5506), .ZN(n5507) );
  NAND2_X1 U6652 ( .A1(n6016), .A2(n5507), .ZN(n6029) );
  OAI22_X1 U6653 ( .A1(n5508), .A2(n6444), .B1(n6440), .B2(n6029), .ZN(n5509)
         );
  AOI211_X1 U6654 ( .C1(n6441), .C2(EBX_REG_11__SCAN_IN), .A(n5509), .B(n6429), 
        .ZN(n5510) );
  OAI21_X1 U6655 ( .B1(n6462), .B2(n5828), .A(n5510), .ZN(n5511) );
  AOI21_X1 U6656 ( .B1(n6377), .B2(n5512), .A(n5511), .ZN(n5513) );
  OAI21_X1 U6657 ( .B1(n5661), .B2(n6435), .A(n5513), .ZN(U2816) );
  INV_X1 U6658 ( .A(n5517), .ZN(n5514) );
  OAI21_X1 U6659 ( .B1(n5515), .B2(n5514), .A(n6435), .ZN(n6464) );
  INV_X1 U6660 ( .A(n6464), .ZN(n5561) );
  AOI21_X1 U6661 ( .B1(n6459), .B2(n5518), .A(n6458), .ZN(n5540) );
  INV_X1 U6662 ( .A(n5540), .ZN(n5530) );
  NAND2_X1 U6663 ( .A1(n5517), .A2(n5516), .ZN(n6456) );
  INV_X1 U6664 ( .A(n5518), .ZN(n5519) );
  AND2_X1 U6665 ( .A1(n6459), .A2(n5519), .ZN(n6447) );
  NAND2_X1 U6666 ( .A1(n6447), .A2(n6748), .ZN(n5525) );
  OAI22_X1 U6667 ( .A1(n5520), .A2(n6467), .B1(n6440), .B2(n6641), .ZN(n5521)
         );
  INV_X1 U6668 ( .A(n5521), .ZN(n5522) );
  NAND2_X1 U6669 ( .A1(n6442), .A2(n5522), .ZN(n5523) );
  AOI21_X1 U6670 ( .B1(n6452), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n5523), 
        .ZN(n5524) );
  OAI211_X1 U6671 ( .C1(n6456), .C2(n5526), .A(n5525), .B(n5524), .ZN(n5529)
         );
  NOR2_X1 U6672 ( .A1(n6462), .A2(n5527), .ZN(n5528) );
  AOI211_X1 U6673 ( .C1(REIP_REG_4__SCAN_IN), .C2(n5530), .A(n5529), .B(n5528), 
        .ZN(n5531) );
  OAI21_X1 U6674 ( .B1(n5561), .B2(n5532), .A(n5531), .ZN(U2823) );
  INV_X1 U6675 ( .A(n6588), .ZN(n5542) );
  INV_X1 U6676 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6746) );
  NOR2_X1 U6677 ( .A1(n6746), .A2(n6792), .ZN(n5533) );
  AOI21_X1 U6678 ( .B1(n6423), .B2(n5533), .A(REIP_REG_3__SCAN_IN), .ZN(n5539)
         );
  INV_X1 U6679 ( .A(n6456), .ZN(n5552) );
  AOI22_X1 U6680 ( .A1(n5552), .A2(n6206), .B1(n6452), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5538) );
  OR2_X1 U6681 ( .A1(n4468), .A2(n5534), .ZN(n5535) );
  AND2_X1 U6682 ( .A1(n5536), .A2(n5535), .ZN(n6650) );
  AOI22_X1 U6683 ( .A1(n6451), .A2(n6650), .B1(n6441), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n5537) );
  OAI211_X1 U6684 ( .C1(n5540), .C2(n5539), .A(n5538), .B(n5537), .ZN(n5541)
         );
  AOI21_X1 U6685 ( .B1(n6427), .B2(n5542), .A(n5541), .ZN(n5543) );
  OAI21_X1 U6686 ( .B1(n5561), .B2(n6476), .A(n5543), .ZN(U2824) );
  INV_X1 U6687 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5549) );
  OAI22_X1 U6688 ( .A1(n4384), .A2(n6467), .B1(n6424), .B2(REIP_REG_1__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U6689 ( .A1(n6451), .A2(n5544), .ZN(n5546) );
  AOI22_X1 U6690 ( .A1(n6452), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6458), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n5545) );
  OAI211_X1 U6691 ( .C1(n6456), .C2(n6054), .A(n5546), .B(n5545), .ZN(n5547)
         );
  AOI211_X1 U6692 ( .C1(n3090), .C2(n5549), .A(n5548), .B(n5547), .ZN(n5550)
         );
  OAI21_X1 U6693 ( .B1(n5561), .B2(n5551), .A(n5550), .ZN(U2826) );
  NAND2_X1 U6694 ( .A1(n6462), .A2(n6444), .ZN(n5558) );
  AOI22_X1 U6695 ( .A1(n6667), .A2(n5552), .B1(n6441), .B2(EBX_REG_0__SCAN_IN), 
        .ZN(n5555) );
  NAND2_X1 U6696 ( .A1(n6451), .A2(n5553), .ZN(n5554) );
  OAI211_X1 U6697 ( .C1(n5556), .C2(n7076), .A(n5555), .B(n5554), .ZN(n5557)
         );
  AOI21_X1 U6698 ( .B1(n5558), .B2(PHYADDRPOINTER_REG_0__SCAN_IN), .A(n5557), 
        .ZN(n5559) );
  OAI21_X1 U6699 ( .B1(n5561), .B2(n5560), .A(n5559), .ZN(U2827) );
  AOI22_X1 U6700 ( .A1(n5863), .A2(n6477), .B1(EBX_REG_29__SCAN_IN), .B2(n5597), .ZN(n5562) );
  OAI21_X1 U6701 ( .B1(n5613), .B2(n6471), .A(n5562), .ZN(U2830) );
  OAI222_X1 U6702 ( .A1(n5688), .A2(n5599), .B1(n5564), .B2(n6480), .C1(n5563), 
        .C2(n5605), .ZN(U2831) );
  INV_X1 U6703 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5565) );
  OAI222_X1 U6704 ( .A1(n5696), .A2(n5599), .B1(n5565), .B2(n6480), .C1(n5605), 
        .C2(n5882), .ZN(U2832) );
  OAI222_X1 U6705 ( .A1(n5599), .A2(n5702), .B1(n7040), .B2(n6480), .C1(n5889), 
        .C2(n5605), .ZN(U2833) );
  OAI222_X1 U6706 ( .A1(n5622), .A2(n5599), .B1(n6832), .B2(n6480), .C1(n5900), 
        .C2(n5605), .ZN(U2834) );
  INV_X1 U6707 ( .A(n5566), .ZN(n5625) );
  AOI22_X1 U6708 ( .A1(n5567), .A2(n6477), .B1(EBX_REG_24__SCAN_IN), .B2(n5597), .ZN(n5568) );
  OAI21_X1 U6709 ( .B1(n5625), .B2(n6471), .A(n5568), .ZN(U2835) );
  AOI22_X1 U6710 ( .A1(n5569), .A2(n6477), .B1(EBX_REG_23__SCAN_IN), .B2(n5597), .ZN(n5570) );
  OAI21_X1 U6711 ( .B1(n5628), .B2(n6471), .A(n5570), .ZN(U2836) );
  INV_X1 U6712 ( .A(n5727), .ZN(n5631) );
  INV_X1 U6713 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5571) );
  OAI222_X1 U6714 ( .A1(n5599), .A2(n5631), .B1(n5571), .B2(n6480), .C1(n5907), 
        .C2(n5605), .ZN(U2837) );
  INV_X1 U6715 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5572) );
  OAI222_X1 U6716 ( .A1(n5737), .A2(n5599), .B1(n5572), .B2(n6480), .C1(n5917), 
        .C2(n5605), .ZN(U2838) );
  INV_X1 U6717 ( .A(EBX_REG_20__SCAN_IN), .ZN(n6820) );
  INV_X1 U6718 ( .A(n5931), .ZN(n5573) );
  OAI222_X1 U6719 ( .A1(n5636), .A2(n5599), .B1(n6820), .B2(n6480), .C1(n5605), 
        .C2(n5573), .ZN(U2839) );
  OAI222_X1 U6720 ( .A1(n5639), .A2(n5599), .B1(n6912), .B2(n6480), .C1(n5605), 
        .C2(n5939), .ZN(U2840) );
  INV_X1 U6721 ( .A(n5947), .ZN(n5574) );
  OAI222_X1 U6722 ( .A1(n5642), .A2(n5599), .B1(n7101), .B2(n6480), .C1(n5574), 
        .C2(n5605), .ZN(U2841) );
  INV_X1 U6723 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5575) );
  OAI222_X1 U6724 ( .A1(n5774), .A2(n6471), .B1(n5575), .B2(n6480), .C1(n5956), 
        .C2(n5605), .ZN(U2842) );
  AOI22_X1 U6725 ( .A1(n5966), .A2(n6477), .B1(EBX_REG_16__SCAN_IN), .B2(n5597), .ZN(n5576) );
  OAI21_X1 U6726 ( .B1(n5649), .B2(n6471), .A(n5576), .ZN(U2843) );
  INV_X1 U6727 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5577) );
  INV_X1 U6728 ( .A(n5791), .ZN(n5651) );
  OAI222_X1 U6729 ( .A1(n5974), .A2(n5605), .B1(n5577), .B2(n6480), .C1(n5651), 
        .C2(n6471), .ZN(U2844) );
  OAI22_X1 U6730 ( .A1(n5982), .A2(n5605), .B1(n5578), .B2(n6480), .ZN(n5579)
         );
  INV_X1 U6731 ( .A(n5579), .ZN(n5580) );
  OAI21_X1 U6732 ( .B1(n5653), .B2(n6471), .A(n5580), .ZN(U2845) );
  INV_X1 U6733 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5582) );
  OAI222_X1 U6734 ( .A1(n5802), .A2(n5599), .B1(n6480), .B2(n5582), .C1(n5581), 
        .C2(n5605), .ZN(U2846) );
  INV_X1 U6735 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5583) );
  OAI222_X1 U6736 ( .A1(n5661), .A2(n5599), .B1(n6480), .B2(n5583), .C1(n6029), 
        .C2(n5605), .ZN(U2848) );
  NAND2_X1 U6737 ( .A1(n5593), .A2(n5584), .ZN(n5585) );
  NOR2_X1 U6738 ( .A1(n5595), .A2(n5587), .ZN(n5588) );
  OR2_X1 U6739 ( .A1(n5589), .A2(n5588), .ZN(n6398) );
  OAI22_X1 U6740 ( .A1(n6398), .A2(n5605), .B1(n5590), .B2(n6480), .ZN(n5591)
         );
  INV_X1 U6741 ( .A(n5591), .ZN(n5592) );
  OAI21_X1 U6742 ( .B1(n5663), .B2(n6471), .A(n5592), .ZN(U2849) );
  OAI21_X1 U6743 ( .B1(n3085), .B2(n5594), .A(n5593), .ZN(n6402) );
  AOI21_X1 U6744 ( .B1(n3246), .B2(n5596), .A(n5595), .ZN(n6603) );
  AOI22_X1 U6745 ( .A1(n6603), .A2(n6477), .B1(EBX_REG_9__SCAN_IN), .B2(n5597), 
        .ZN(n5598) );
  OAI21_X1 U6746 ( .B1(n6402), .B2(n5599), .A(n5598), .ZN(U2850) );
  NOR2_X1 U6747 ( .A1(n3104), .A2(n5600), .ZN(n5601) );
  OR2_X1 U6748 ( .A1(n3085), .A2(n5601), .ZN(n6410) );
  NAND2_X1 U6749 ( .A1(n5603), .A2(n5602), .ZN(n5604) );
  NAND2_X1 U6750 ( .A1(n3246), .A2(n5604), .ZN(n6610) );
  OAI22_X1 U6751 ( .A1(n6610), .A2(n5605), .B1(n6408), .B2(n6480), .ZN(n5606)
         );
  INV_X1 U6752 ( .A(n5606), .ZN(n5607) );
  OAI21_X1 U6753 ( .B1(n6410), .B2(n6471), .A(n5607), .ZN(U2851) );
  AOI22_X1 U6754 ( .A1(n5645), .A2(DATAI_30_), .B1(n5658), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U6755 ( .A1(n5646), .A2(DATAI_14_), .ZN(n5608) );
  OAI211_X1 U6756 ( .C1(n5610), .C2(n5662), .A(n5609), .B(n5608), .ZN(U2861)
         );
  AOI22_X1 U6757 ( .A1(n5645), .A2(DATAI_29_), .B1(n5658), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5612) );
  NAND2_X1 U6758 ( .A1(n5646), .A2(DATAI_13_), .ZN(n5611) );
  OAI211_X1 U6759 ( .C1(n5613), .C2(n5662), .A(n5612), .B(n5611), .ZN(U2862)
         );
  AOI22_X1 U6760 ( .A1(n5645), .A2(DATAI_28_), .B1(n5658), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5615) );
  NAND2_X1 U6761 ( .A1(n5646), .A2(DATAI_12_), .ZN(n5614) );
  OAI211_X1 U6762 ( .C1(n5688), .C2(n5662), .A(n5615), .B(n5614), .ZN(U2863)
         );
  AOI22_X1 U6763 ( .A1(n5645), .A2(DATAI_27_), .B1(n5658), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U6764 ( .A1(n5646), .A2(DATAI_11_), .ZN(n5616) );
  OAI211_X1 U6765 ( .C1(n5696), .C2(n5662), .A(n5617), .B(n5616), .ZN(U2864)
         );
  AOI22_X1 U6766 ( .A1(n5645), .A2(DATAI_26_), .B1(n5658), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5619) );
  NAND2_X1 U6767 ( .A1(n5646), .A2(DATAI_10_), .ZN(n5618) );
  OAI211_X1 U6768 ( .C1(n5702), .C2(n5662), .A(n5619), .B(n5618), .ZN(U2865)
         );
  AOI22_X1 U6769 ( .A1(n5645), .A2(DATAI_25_), .B1(n5658), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5621) );
  NAND2_X1 U6770 ( .A1(n5646), .A2(DATAI_9_), .ZN(n5620) );
  OAI211_X1 U6771 ( .C1(n5622), .C2(n5662), .A(n5621), .B(n5620), .ZN(U2866)
         );
  AOI22_X1 U6772 ( .A1(n5645), .A2(DATAI_24_), .B1(n5658), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5624) );
  NAND2_X1 U6773 ( .A1(n5646), .A2(DATAI_8_), .ZN(n5623) );
  OAI211_X1 U6774 ( .C1(n5625), .C2(n5662), .A(n5624), .B(n5623), .ZN(U2867)
         );
  AOI22_X1 U6775 ( .A1(n5645), .A2(DATAI_23_), .B1(n5658), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5627) );
  NAND2_X1 U6776 ( .A1(n5646), .A2(DATAI_7_), .ZN(n5626) );
  OAI211_X1 U6777 ( .C1(n5628), .C2(n5662), .A(n5627), .B(n5626), .ZN(U2868)
         );
  AOI22_X1 U6778 ( .A1(n5645), .A2(DATAI_22_), .B1(n5658), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5630) );
  NAND2_X1 U6779 ( .A1(n5646), .A2(DATAI_6_), .ZN(n5629) );
  OAI211_X1 U6780 ( .C1(n5631), .C2(n5662), .A(n5630), .B(n5629), .ZN(U2869)
         );
  AOI22_X1 U6781 ( .A1(n5645), .A2(DATAI_21_), .B1(n5658), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5633) );
  NAND2_X1 U6782 ( .A1(n5646), .A2(DATAI_5_), .ZN(n5632) );
  OAI211_X1 U6783 ( .C1(n5737), .C2(n5662), .A(n5633), .B(n5632), .ZN(U2870)
         );
  AOI22_X1 U6784 ( .A1(n5645), .A2(DATAI_20_), .B1(n5658), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5635) );
  NAND2_X1 U6785 ( .A1(n5646), .A2(DATAI_4_), .ZN(n5634) );
  OAI211_X1 U6786 ( .C1(n5636), .C2(n5662), .A(n5635), .B(n5634), .ZN(U2871)
         );
  AOI22_X1 U6787 ( .A1(n5645), .A2(DATAI_19_), .B1(n5658), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U6788 ( .A1(n5646), .A2(DATAI_3_), .ZN(n5637) );
  OAI211_X1 U6789 ( .C1(n5639), .C2(n5662), .A(n5638), .B(n5637), .ZN(U2872)
         );
  AOI22_X1 U6790 ( .A1(n5645), .A2(DATAI_18_), .B1(n5658), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5641) );
  NAND2_X1 U6791 ( .A1(n5646), .A2(DATAI_2_), .ZN(n5640) );
  OAI211_X1 U6792 ( .C1(n5642), .C2(n5662), .A(n5641), .B(n5640), .ZN(U2873)
         );
  AOI22_X1 U6793 ( .A1(n5645), .A2(DATAI_17_), .B1(n5658), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5644) );
  NAND2_X1 U6794 ( .A1(n5646), .A2(DATAI_1_), .ZN(n5643) );
  OAI211_X1 U6795 ( .C1(n5774), .C2(n5662), .A(n5644), .B(n5643), .ZN(U2874)
         );
  AOI22_X1 U6796 ( .A1(n5645), .A2(DATAI_16_), .B1(n5658), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U6797 ( .A1(n5646), .A2(DATAI_0_), .ZN(n5647) );
  OAI211_X1 U6798 ( .C1(n5649), .C2(n5662), .A(n5648), .B(n5647), .ZN(U2875)
         );
  AOI22_X1 U6799 ( .A1(n5659), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n5658), .ZN(n5650) );
  OAI21_X1 U6800 ( .B1(n5651), .B2(n5662), .A(n5650), .ZN(U2876) );
  AOI22_X1 U6801 ( .A1(n5659), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n5658), .ZN(n5652) );
  OAI21_X1 U6802 ( .B1(n5653), .B2(n5662), .A(n5652), .ZN(U2877) );
  INV_X1 U6803 ( .A(DATAI_13_), .ZN(n6555) );
  INV_X1 U6804 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6495) );
  OAI222_X1 U6805 ( .A1(n5802), .A2(n5662), .B1(n5665), .B2(n6555), .C1(n5664), 
        .C2(n6495), .ZN(U2878) );
  NOR2_X1 U6806 ( .A1(n5655), .A2(n5654), .ZN(n5656) );
  INV_X1 U6807 ( .A(DATAI_12_), .ZN(n6949) );
  OAI222_X1 U6808 ( .A1(n6472), .A2(n5662), .B1(n5665), .B2(n6949), .C1(n5664), 
        .C2(n4059), .ZN(U2879) );
  AOI22_X1 U6809 ( .A1(n5659), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n5658), .ZN(n5660) );
  OAI21_X1 U6810 ( .B1(n5661), .B2(n5662), .A(n5660), .ZN(U2880) );
  INV_X1 U6811 ( .A(DATAI_10_), .ZN(n6549) );
  INV_X1 U6812 ( .A(EAX_REG_10__SCAN_IN), .ZN(n7092) );
  OAI222_X1 U6813 ( .A1(n5663), .A2(n5662), .B1(n5665), .B2(n6549), .C1(n5664), 
        .C2(n7092), .ZN(U2881) );
  INV_X1 U6814 ( .A(DATAI_9_), .ZN(n6547) );
  INV_X1 U6815 ( .A(EAX_REG_9__SCAN_IN), .ZN(n7025) );
  OAI222_X1 U6816 ( .A1(n6402), .A2(n5662), .B1(n5665), .B2(n6547), .C1(n5664), 
        .C2(n7025), .ZN(U2882) );
  INV_X1 U6817 ( .A(DATAI_8_), .ZN(n6848) );
  INV_X1 U6818 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6879) );
  OAI222_X1 U6819 ( .A1(n6410), .A2(n5662), .B1(n5665), .B2(n6848), .C1(n5664), 
        .C2(n6879), .ZN(U2883) );
  NAND2_X1 U6820 ( .A1(n5666), .A2(n5855), .ZN(n5668) );
  OAI211_X1 U6821 ( .C1(n5669), .C2(n5853), .A(n5668), .B(n5667), .ZN(n5670)
         );
  AOI21_X1 U6822 ( .B1(n5671), .B2(n5839), .A(n5670), .ZN(n5672) );
  OAI21_X1 U6823 ( .B1(n5673), .B2(n6362), .A(n5672), .ZN(U2956) );
  INV_X1 U6824 ( .A(n5681), .ZN(n5691) );
  AOI21_X1 U6825 ( .B1(n5682), .B2(n5691), .A(n5674), .ZN(n5675) );
  XNOR2_X1 U6826 ( .A(n5675), .B(n5864), .ZN(n5868) );
  NOR2_X1 U6827 ( .A1(n6639), .A2(n6952), .ZN(n5859) );
  AOI21_X1 U6828 ( .B1(n6591), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5859), 
        .ZN(n5676) );
  OAI21_X1 U6829 ( .B1(n5677), .B2(n6599), .A(n5676), .ZN(n5678) );
  AOI21_X1 U6830 ( .B1(n5679), .B2(n5839), .A(n5678), .ZN(n5680) );
  OAI21_X1 U6831 ( .B1(n5868), .B2(n6362), .A(n5680), .ZN(U2957) );
  INV_X1 U6832 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5870) );
  NAND2_X1 U6833 ( .A1(n5870), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U6834 ( .A1(n5879), .A2(n6592), .ZN(n5687) );
  NOR2_X1 U6835 ( .A1(n6639), .A2(n6784), .ZN(n5872) );
  NOR2_X1 U6836 ( .A1(n5684), .A2(n6599), .ZN(n5685) );
  AOI211_X1 U6837 ( .C1(PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n6591), .A(n5872), 
        .B(n5685), .ZN(n5686) );
  OAI211_X1 U6838 ( .C1(n5858), .C2(n5688), .A(n5687), .B(n5686), .ZN(U2958)
         );
  NOR2_X1 U6839 ( .A1(n6639), .A2(n6779), .ZN(n5884) );
  NOR2_X1 U6840 ( .A1(n5689), .A2(n6599), .ZN(n5690) );
  AOI211_X1 U6841 ( .C1(PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n6591), .A(n5884), 
        .B(n5690), .ZN(n5695) );
  XNOR2_X1 U6842 ( .A(n5693), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5880)
         );
  NAND2_X1 U6843 ( .A1(n5880), .A2(n6592), .ZN(n5694) );
  OAI211_X1 U6844 ( .C1(n5696), .C2(n5858), .A(n5695), .B(n5694), .ZN(U2959)
         );
  NOR2_X1 U6845 ( .A1(n3214), .A2(n5698), .ZN(n5700) );
  XOR2_X1 U6846 ( .A(n5700), .B(n5699), .Z(n5897) );
  NAND2_X1 U6847 ( .A1(n6577), .A2(REIP_REG_26__SCAN_IN), .ZN(n5890) );
  OAI21_X1 U6848 ( .B1(n5853), .B2(n5701), .A(n5890), .ZN(n5704) );
  NOR2_X1 U6849 ( .A1(n5702), .A2(n5858), .ZN(n5703) );
  AOI211_X1 U6850 ( .C1(n5705), .C2(n5855), .A(n5704), .B(n5703), .ZN(n5706)
         );
  NOR3_X1 U6851 ( .A1(n5910), .A2(n5707), .A3(n5924), .ZN(n5709) );
  XNOR2_X1 U6852 ( .A(n5815), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5708)
         );
  AOI21_X1 U6853 ( .B1(n5747), .B2(n5709), .A(n5708), .ZN(n5714) );
  OAI21_X1 U6854 ( .B1(n5747), .B2(n5710), .A(n5815), .ZN(n5713) );
  INV_X1 U6855 ( .A(n5711), .ZN(n5712) );
  AOI21_X1 U6856 ( .B1(n5714), .B2(n5713), .A(n5712), .ZN(n5905) );
  NAND2_X1 U6857 ( .A1(n6577), .A2(REIP_REG_25__SCAN_IN), .ZN(n5898) );
  NAND2_X1 U6858 ( .A1(n6591), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5715)
         );
  OAI211_X1 U6859 ( .C1(n5716), .C2(n6599), .A(n5898), .B(n5715), .ZN(n5717)
         );
  AOI21_X1 U6860 ( .B1(n5718), .B2(n5839), .A(n5717), .ZN(n5719) );
  OAI21_X1 U6861 ( .B1(n5905), .B2(n6362), .A(n5719), .ZN(U2961) );
  OAI21_X1 U6862 ( .B1(n5813), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5729), 
        .ZN(n5722) );
  AOI21_X1 U6863 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5815), .A(n3279), 
        .ZN(n5721) );
  XNOR2_X1 U6864 ( .A(n5722), .B(n5721), .ZN(n5915) );
  NOR2_X1 U6865 ( .A1(n6639), .A2(n5723), .ZN(n5909) );
  AOI21_X1 U6866 ( .B1(n6591), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5909), 
        .ZN(n5724) );
  OAI21_X1 U6867 ( .B1(n5725), .B2(n6599), .A(n5724), .ZN(n5726) );
  AOI21_X1 U6868 ( .B1(n5727), .B2(n5839), .A(n5726), .ZN(n5728) );
  OAI21_X1 U6869 ( .B1(n5915), .B2(n6362), .A(n5728), .ZN(U2964) );
  OAI21_X1 U6870 ( .B1(n5731), .B2(n5730), .A(n5729), .ZN(n5916) );
  NAND2_X1 U6871 ( .A1(n5916), .A2(n6592), .ZN(n5736) );
  NOR2_X1 U6872 ( .A1(n6639), .A2(n5732), .ZN(n5919) );
  NOR2_X1 U6873 ( .A1(n5853), .A2(n6953), .ZN(n5733) );
  AOI211_X1 U6874 ( .C1(n5855), .C2(n5734), .A(n5919), .B(n5733), .ZN(n5735)
         );
  OAI211_X1 U6875 ( .C1(n5858), .C2(n5737), .A(n5736), .B(n5735), .ZN(U2965)
         );
  XNOR2_X1 U6876 ( .A(n5815), .B(n5738), .ZN(n5739) );
  XNOR2_X1 U6877 ( .A(n5740), .B(n5739), .ZN(n5934) );
  NOR2_X1 U6878 ( .A1(n6639), .A2(n6770), .ZN(n5927) );
  AOI21_X1 U6879 ( .B1(n6591), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n5927), 
        .ZN(n5741) );
  OAI21_X1 U6880 ( .B1(n5742), .B2(n6599), .A(n5741), .ZN(n5743) );
  AOI21_X1 U6881 ( .B1(n5744), .B2(n5839), .A(n5743), .ZN(n5745) );
  OAI21_X1 U6882 ( .B1(n5934), .B2(n6362), .A(n5745), .ZN(U2966) );
  INV_X1 U6883 ( .A(n5747), .ZN(n5749) );
  XNOR2_X1 U6884 ( .A(n5824), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5748)
         );
  OAI22_X1 U6885 ( .A1(n3282), .A2(n5750), .B1(n5749), .B2(n5748), .ZN(n5943)
         );
  NAND2_X1 U6886 ( .A1(n6577), .A2(REIP_REG_19__SCAN_IN), .ZN(n5937) );
  NAND2_X1 U6887 ( .A1(n6591), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5751)
         );
  OAI211_X1 U6888 ( .C1(n6599), .C2(n5752), .A(n5937), .B(n5751), .ZN(n5753)
         );
  AOI21_X1 U6889 ( .B1(n5754), .B2(n5839), .A(n5753), .ZN(n5755) );
  OAI21_X1 U6890 ( .B1(n5943), .B2(n6362), .A(n5755), .ZN(U2967) );
  NAND2_X1 U6891 ( .A1(n5813), .A2(n7058), .ZN(n5765) );
  NOR3_X1 U6892 ( .A1(n5756), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5765), 
        .ZN(n5766) );
  NOR2_X1 U6893 ( .A1(n5768), .A2(n5766), .ZN(n5757) );
  XNOR2_X1 U6894 ( .A(n5757), .B(n5950), .ZN(n5954) );
  NAND2_X1 U6895 ( .A1(n5855), .A2(n5758), .ZN(n5759) );
  NAND2_X1 U6896 ( .A1(n6577), .A2(REIP_REG_18__SCAN_IN), .ZN(n5945) );
  OAI211_X1 U6897 ( .C1(n5853), .C2(n5760), .A(n5759), .B(n5945), .ZN(n5761)
         );
  AOI21_X1 U6898 ( .B1(n5762), .B2(n5839), .A(n5761), .ZN(n5763) );
  OAI21_X1 U6899 ( .B1(n5954), .B2(n6362), .A(n5763), .ZN(U2968) );
  INV_X1 U6900 ( .A(n5766), .ZN(n5767) );
  NAND2_X1 U6901 ( .A1(n5955), .A2(n6592), .ZN(n5773) );
  NOR2_X1 U6902 ( .A1(n6639), .A2(n6766), .ZN(n5958) );
  NOR2_X1 U6903 ( .A1(n5853), .A2(n5769), .ZN(n5770) );
  AOI211_X1 U6904 ( .C1(n5855), .C2(n5771), .A(n5958), .B(n5770), .ZN(n5772)
         );
  XNOR2_X1 U6905 ( .A(n5824), .B(n7058), .ZN(n5775) );
  XNOR2_X1 U6906 ( .A(n5776), .B(n5775), .ZN(n5973) );
  NOR2_X1 U6907 ( .A1(n6639), .A2(n5777), .ZN(n5965) );
  INV_X1 U6908 ( .A(n5965), .ZN(n5780) );
  OR2_X1 U6909 ( .A1(n5853), .A2(n5778), .ZN(n5779) );
  OAI211_X1 U6910 ( .C1(n6599), .C2(n5781), .A(n5780), .B(n5779), .ZN(n5782)
         );
  AOI21_X1 U6911 ( .B1(n5783), .B2(n6594), .A(n5782), .ZN(n5784) );
  OAI21_X1 U6912 ( .B1(n5973), .B2(n6362), .A(n5784), .ZN(U2970) );
  XNOR2_X1 U6913 ( .A(n5824), .B(n7023), .ZN(n5785) );
  XNOR2_X1 U6914 ( .A(n5786), .B(n5785), .ZN(n5981) );
  NOR2_X1 U6915 ( .A1(n6639), .A2(n5787), .ZN(n5976) );
  AOI21_X1 U6916 ( .B1(n6591), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5976), 
        .ZN(n5788) );
  OAI21_X1 U6917 ( .B1(n5789), .B2(n6599), .A(n5788), .ZN(n5790) );
  AOI21_X1 U6918 ( .B1(n5791), .B2(n5839), .A(n5790), .ZN(n5792) );
  OAI21_X1 U6919 ( .B1(n5981), .B2(n6362), .A(n5792), .ZN(U2971) );
  XNOR2_X1 U6920 ( .A(n5824), .B(n5994), .ZN(n5794) );
  XNOR2_X1 U6921 ( .A(n5793), .B(n5794), .ZN(n6000) );
  NAND2_X1 U6922 ( .A1(n6577), .A2(REIP_REG_14__SCAN_IN), .ZN(n5993) );
  NAND2_X1 U6923 ( .A1(n6591), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5795)
         );
  OAI211_X1 U6924 ( .C1(n6599), .C2(n5796), .A(n5993), .B(n5795), .ZN(n5797)
         );
  AOI21_X1 U6925 ( .B1(n5798), .B2(n5839), .A(n5797), .ZN(n5799) );
  OAI21_X1 U6926 ( .B1(n6362), .B2(n6000), .A(n5799), .ZN(U2972) );
  XOR2_X1 U6927 ( .A(n5801), .B(n5800), .Z(n6012) );
  INV_X1 U6928 ( .A(n5802), .ZN(n5806) );
  NAND2_X1 U6929 ( .A1(n6577), .A2(REIP_REG_13__SCAN_IN), .ZN(n6005) );
  NAND2_X1 U6930 ( .A1(n6591), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5803)
         );
  OAI211_X1 U6931 ( .C1(n6599), .C2(n5804), .A(n6005), .B(n5803), .ZN(n5805)
         );
  AOI21_X1 U6932 ( .B1(n5806), .B2(n5839), .A(n5805), .ZN(n5807) );
  OAI21_X1 U6933 ( .B1(n6362), .B2(n6012), .A(n5807), .ZN(U2973) );
  NOR2_X1 U6934 ( .A1(n5815), .A2(n5811), .ZN(n5822) );
  NAND2_X1 U6935 ( .A1(n5808), .A2(n5809), .ZN(n5810) );
  NAND2_X1 U6936 ( .A1(n5824), .A2(n5811), .ZN(n5832) );
  NAND2_X1 U6937 ( .A1(n5834), .A2(n5832), .ZN(n5823) );
  AOI21_X1 U6938 ( .B1(n5815), .B2(n6031), .A(n5823), .ZN(n5812) );
  AOI211_X1 U6939 ( .C1(INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n5813), .A(n5822), .B(n5812), .ZN(n5817) );
  OAI21_X1 U6940 ( .B1(n5815), .B2(n6021), .A(n5814), .ZN(n5816) );
  XNOR2_X1 U6941 ( .A(n5817), .B(n5816), .ZN(n6025) );
  NAND2_X1 U6942 ( .A1(n6577), .A2(REIP_REG_12__SCAN_IN), .ZN(n6017) );
  OAI21_X1 U6943 ( .B1(n5853), .B2(n5818), .A(n6017), .ZN(n5820) );
  NOR2_X1 U6944 ( .A1(n6472), .A2(n5858), .ZN(n5819) );
  AOI211_X1 U6945 ( .C1(n5855), .C2(n6378), .A(n5820), .B(n5819), .ZN(n5821)
         );
  OAI21_X1 U6946 ( .B1(n6025), .B2(n6362), .A(n5821), .ZN(U2974) );
  INV_X1 U6947 ( .A(n5822), .ZN(n5833) );
  NAND2_X1 U6948 ( .A1(n5823), .A2(n5833), .ZN(n5826) );
  XNOR2_X1 U6949 ( .A(n5824), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5825)
         );
  XNOR2_X1 U6950 ( .A(n5826), .B(n5825), .ZN(n6034) );
  NAND2_X1 U6951 ( .A1(n6577), .A2(REIP_REG_11__SCAN_IN), .ZN(n6028) );
  NAND2_X1 U6952 ( .A1(n6591), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5827)
         );
  OAI211_X1 U6953 ( .C1(n6599), .C2(n5828), .A(n6028), .B(n5827), .ZN(n5829)
         );
  AOI21_X1 U6954 ( .B1(n5830), .B2(n5839), .A(n5829), .ZN(n5831) );
  OAI21_X1 U6955 ( .B1(n6034), .B2(n6362), .A(n5831), .ZN(U2975) );
  NAND2_X1 U6956 ( .A1(n5833), .A2(n5832), .ZN(n5835) );
  XOR2_X1 U6957 ( .A(n5835), .B(n5834), .Z(n6048) );
  AOI22_X1 U6958 ( .A1(n6591), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6577), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5836) );
  OAI21_X1 U6959 ( .B1(n5837), .B2(n6599), .A(n5836), .ZN(n5838) );
  AOI21_X1 U6960 ( .B1(n6392), .B2(n5839), .A(n5838), .ZN(n5840) );
  OAI21_X1 U6961 ( .B1(n6048), .B2(n6362), .A(n5840), .ZN(U2976) );
  NAND2_X1 U6962 ( .A1(n5808), .A2(n5841), .ZN(n5845) );
  NAND2_X1 U6963 ( .A1(n5843), .A2(n5842), .ZN(n5844) );
  XNOR2_X1 U6964 ( .A(n5845), .B(n5844), .ZN(n6605) );
  NAND2_X1 U6965 ( .A1(n6605), .A2(n6592), .ZN(n5848) );
  NAND2_X1 U6966 ( .A1(n6577), .A2(REIP_REG_9__SCAN_IN), .ZN(n6601) );
  OAI21_X1 U6967 ( .B1(n5853), .B2(n6401), .A(n6601), .ZN(n5846) );
  AOI21_X1 U6968 ( .B1(n5855), .B2(n6399), .A(n5846), .ZN(n5847) );
  OAI211_X1 U6969 ( .C1(n5858), .C2(n6402), .A(n5848), .B(n5847), .ZN(U2977)
         );
  OAI21_X1 U6970 ( .B1(n5850), .B2(n5849), .A(n5808), .ZN(n5851) );
  INV_X1 U6971 ( .A(n5851), .ZN(n6614) );
  NAND2_X1 U6972 ( .A1(n6614), .A2(n6592), .ZN(n5857) );
  INV_X1 U6973 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5852) );
  OAI22_X1 U6974 ( .A1(n5853), .A2(n5852), .B1(n6639), .B2(n6609), .ZN(n5854)
         );
  AOI21_X1 U6975 ( .B1(n5855), .B2(n6411), .A(n5854), .ZN(n5856) );
  OAI211_X1 U6976 ( .C1(n5858), .C2(n6410), .A(n5857), .B(n5856), .ZN(U2978)
         );
  INV_X1 U6977 ( .A(n5859), .ZN(n5860) );
  OAI21_X1 U6978 ( .B1(n5861), .B2(n5864), .A(n5860), .ZN(n5862) );
  AOI21_X1 U6979 ( .B1(n5863), .B2(n6651), .A(n5862), .ZN(n5867) );
  NAND2_X1 U6980 ( .A1(n5865), .A2(n5864), .ZN(n5866) );
  OAI211_X1 U6981 ( .C1(n5868), .C2(n6638), .A(n5867), .B(n5866), .ZN(U2989)
         );
  INV_X1 U6982 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5869) );
  NAND2_X1 U6983 ( .A1(n5871), .A2(n5869), .ZN(n5886) );
  AOI21_X1 U6984 ( .B1(n5886), .B2(n5881), .A(n5870), .ZN(n5878) );
  INV_X1 U6985 ( .A(n5871), .ZN(n5876) );
  AOI21_X1 U6986 ( .B1(n5873), .B2(n6651), .A(n5872), .ZN(n5874) );
  OAI21_X1 U6987 ( .B1(n5876), .B2(n5875), .A(n5874), .ZN(n5877) );
  INV_X1 U6988 ( .A(n5880), .ZN(n5888) );
  INV_X1 U6989 ( .A(n5881), .ZN(n5885) );
  NOR2_X1 U6990 ( .A1(n5882), .A2(n6640), .ZN(n5883) );
  AOI211_X1 U6991 ( .C1(INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n5885), .A(n5884), .B(n5883), .ZN(n5887) );
  OAI211_X1 U6992 ( .C1(n5888), .C2(n6638), .A(n5887), .B(n5886), .ZN(U2991)
         );
  INV_X1 U6993 ( .A(n5889), .ZN(n5893) );
  INV_X1 U6994 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5891) );
  OAI21_X1 U6995 ( .B1(n5899), .B2(n5891), .A(n5890), .ZN(n5892) );
  AOI21_X1 U6996 ( .B1(n5893), .B2(n6651), .A(n5892), .ZN(n5896) );
  OAI211_X1 U6997 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5903), .B(n5894), .ZN(n5895) );
  OAI211_X1 U6998 ( .C1(n5897), .C2(n6638), .A(n5896), .B(n5895), .ZN(U2992)
         );
  OAI21_X1 U6999 ( .B1(n5899), .B2(n7061), .A(n5898), .ZN(n5902) );
  NOR2_X1 U7000 ( .A1(n5900), .A2(n6640), .ZN(n5901) );
  AOI211_X1 U7001 ( .C1(n5903), .C2(n7061), .A(n5902), .B(n5901), .ZN(n5904)
         );
  OAI21_X1 U7002 ( .B1(n5905), .B2(n6638), .A(n5904), .ZN(U2993) );
  INV_X1 U7003 ( .A(n5906), .ZN(n5920) );
  NOR2_X1 U7004 ( .A1(n5907), .A2(n6640), .ZN(n5908) );
  AOI211_X1 U7005 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5920), .A(n5909), .B(n5908), .ZN(n5914) );
  INV_X1 U7006 ( .A(n5923), .ZN(n5912) );
  NAND3_X1 U7007 ( .A1(n5912), .A2(n5911), .A3(n5910), .ZN(n5913) );
  OAI211_X1 U7008 ( .C1(n5915), .C2(n6638), .A(n5914), .B(n5913), .ZN(U2996)
         );
  NAND2_X1 U7009 ( .A1(n5916), .A2(n6653), .ZN(n5922) );
  NOR2_X1 U7010 ( .A1(n5917), .A2(n6640), .ZN(n5918) );
  AOI211_X1 U7011 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5920), .A(n5919), .B(n5918), .ZN(n5921) );
  OAI211_X1 U7012 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5923), .A(n5922), .B(n5921), .ZN(U2997) );
  INV_X1 U7013 ( .A(n5924), .ZN(n5926) );
  NOR2_X1 U7014 ( .A1(n5926), .A2(n5925), .ZN(n5928) );
  AOI21_X1 U7015 ( .B1(n5936), .B2(n5928), .A(n5927), .ZN(n5933) );
  OR2_X1 U7016 ( .A1(n5929), .A2(n6636), .ZN(n6013) );
  AOI21_X1 U7017 ( .B1(n6013), .B2(n5930), .A(n5959), .ZN(n5951) );
  OAI21_X1 U7018 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n6044), .A(n5951), 
        .ZN(n5941) );
  AOI22_X1 U7019 ( .A1(n5941), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(n5931), .B2(n6651), .ZN(n5932) );
  OAI211_X1 U7020 ( .C1(n5934), .C2(n6638), .A(n5933), .B(n5932), .ZN(U2998)
         );
  NAND2_X1 U7021 ( .A1(n5936), .A2(n5935), .ZN(n5938) );
  OAI211_X1 U7022 ( .C1(n5939), .C2(n6640), .A(n5938), .B(n5937), .ZN(n5940)
         );
  AOI21_X1 U7023 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n5941), .A(n5940), 
        .ZN(n5942) );
  OAI21_X1 U7024 ( .B1(n5943), .B2(n6638), .A(n5942), .ZN(U2999) );
  INV_X1 U7025 ( .A(n5962), .ZN(n5944) );
  NAND3_X1 U7026 ( .A1(n5944), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5950), .ZN(n5949) );
  INV_X1 U7027 ( .A(n5945), .ZN(n5946) );
  AOI21_X1 U7028 ( .B1(n5947), .B2(n6651), .A(n5946), .ZN(n5948) );
  OAI211_X1 U7029 ( .C1(n5951), .C2(n5950), .A(n5949), .B(n5948), .ZN(n5952)
         );
  INV_X1 U7030 ( .A(n5952), .ZN(n5953) );
  OAI21_X1 U7031 ( .B1(n5954), .B2(n6638), .A(n5953), .ZN(U3000) );
  NOR2_X1 U7032 ( .A1(n5956), .A2(n6640), .ZN(n5957) );
  AOI211_X1 U7033 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5959), .A(n5958), .B(n5957), .ZN(n5960) );
  OAI211_X1 U7034 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5962), .A(n5961), .B(n5960), .ZN(U3001) );
  AND3_X1 U7035 ( .A1(n6032), .A2(n5963), .A3(n7058), .ZN(n5964) );
  AOI211_X1 U7036 ( .C1(n6651), .C2(n5966), .A(n5965), .B(n5964), .ZN(n5972)
         );
  INV_X1 U7037 ( .A(n5968), .ZN(n5989) );
  NAND2_X1 U7038 ( .A1(n6032), .A2(n5989), .ZN(n5995) );
  NOR3_X1 U7039 ( .A1(n5995), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .A3(n5994), 
        .ZN(n5978) );
  INV_X1 U7040 ( .A(n6026), .ZN(n5970) );
  OAI21_X1 U7041 ( .B1(n5968), .B2(n5994), .A(n5967), .ZN(n5969) );
  NAND2_X1 U7042 ( .A1(n5970), .A2(n5969), .ZN(n5977) );
  OAI21_X1 U7043 ( .B1(n5978), .B2(n5977), .A(INSTADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n5971) );
  OAI211_X1 U7044 ( .C1(n5973), .C2(n6638), .A(n5972), .B(n5971), .ZN(U3002)
         );
  NOR2_X1 U7045 ( .A1(n5974), .A2(n6640), .ZN(n5975) );
  AOI211_X1 U7046 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n5977), .A(n5976), .B(n5975), .ZN(n5980) );
  INV_X1 U7047 ( .A(n5978), .ZN(n5979) );
  OAI211_X1 U7048 ( .C1(n5981), .C2(n6638), .A(n5980), .B(n5979), .ZN(U3003)
         );
  INV_X1 U7049 ( .A(n5982), .ZN(n5998) );
  INV_X1 U7050 ( .A(n5983), .ZN(n5988) );
  NAND3_X1 U7051 ( .A1(n5985), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .A3(n5984), 
        .ZN(n5987) );
  NAND2_X1 U7052 ( .A1(n5990), .A2(n5986), .ZN(n6002) );
  AOI21_X1 U7053 ( .B1(n5988), .B2(n5987), .A(n6002), .ZN(n6001) );
  OAI22_X1 U7054 ( .A1(n5991), .A2(n5990), .B1(n5989), .B2(n6004), .ZN(n5992)
         );
  NOR3_X1 U7055 ( .A1(n6001), .A2(n5992), .A3(n6026), .ZN(n6008) );
  OAI21_X1 U7056 ( .B1(n6008), .B2(n5994), .A(n5993), .ZN(n5997) );
  NOR2_X1 U7057 ( .A1(n5995), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5996)
         );
  AOI211_X1 U7058 ( .C1(n6651), .C2(n5998), .A(n5997), .B(n5996), .ZN(n5999)
         );
  OAI21_X1 U7059 ( .B1(n6000), .B2(n6638), .A(n5999), .ZN(U3004) );
  NOR2_X1 U7060 ( .A1(n6001), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6007)
         );
  OR3_X1 U7061 ( .A1(n6004), .A2(n6003), .A3(n6002), .ZN(n6006) );
  OAI211_X1 U7062 ( .C1(n6008), .C2(n6007), .A(n6006), .B(n6005), .ZN(n6009)
         );
  AOI21_X1 U7063 ( .B1(n6651), .B2(n6010), .A(n6009), .ZN(n6011) );
  OAI21_X1 U7064 ( .B1(n6012), .B2(n6638), .A(n6011), .ZN(U3005) );
  AOI21_X1 U7065 ( .B1(n6013), .B2(n6031), .A(n6026), .ZN(n6022) );
  INV_X1 U7066 ( .A(n6014), .ZN(n6015) );
  XNOR2_X1 U7067 ( .A(n6016), .B(n6015), .ZN(n6469) );
  INV_X1 U7068 ( .A(n6017), .ZN(n6018) );
  AOI21_X1 U7069 ( .B1(n6469), .B2(n6651), .A(n6018), .ZN(n6020) );
  NAND3_X1 U7070 ( .A1(n6032), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n6021), .ZN(n6019) );
  OAI211_X1 U7071 ( .C1(n6022), .C2(n6021), .A(n6020), .B(n6019), .ZN(n6023)
         );
  INV_X1 U7072 ( .A(n6023), .ZN(n6024) );
  OAI21_X1 U7073 ( .B1(n6025), .B2(n6638), .A(n6024), .ZN(U3006) );
  NAND2_X1 U7074 ( .A1(n6026), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6027) );
  OAI211_X1 U7075 ( .C1(n6029), .C2(n6640), .A(n6028), .B(n6027), .ZN(n6030)
         );
  AOI21_X1 U7076 ( .B1(n6032), .B2(n6031), .A(n6030), .ZN(n6033) );
  OAI21_X1 U7077 ( .B1(n6034), .B2(n6638), .A(n6033), .ZN(U3007) );
  NAND2_X1 U7078 ( .A1(n6039), .A2(n6035), .ZN(n6623) );
  NOR2_X1 U7079 ( .A1(n6037), .A2(n6623), .ZN(n6604) );
  OAI211_X1 U7080 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6604), .B(n6036), .ZN(n6047) );
  INV_X1 U7081 ( .A(n6037), .ZN(n6611) );
  OAI22_X1 U7082 ( .A1(n6041), .A2(n6040), .B1(n6039), .B2(n6038), .ZN(n6042)
         );
  NOR2_X1 U7083 ( .A1(n6043), .A2(n6042), .ZN(n6621) );
  OAI21_X1 U7084 ( .B1(n6611), .B2(n6044), .A(n6621), .ZN(n6600) );
  INV_X1 U7085 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6965) );
  OAI22_X1 U7086 ( .A1(n6398), .A2(n6640), .B1(n6965), .B2(n6639), .ZN(n6045)
         );
  AOI21_X1 U7087 ( .B1(n6600), .B2(INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6045), 
        .ZN(n6046) );
  OAI211_X1 U7088 ( .C1(n6048), .C2(n6638), .A(n6047), .B(n6046), .ZN(U3008)
         );
  INV_X1 U7089 ( .A(n6049), .ZN(n6057) );
  OAI222_X1 U7090 ( .A1(n6804), .A2(n3912), .B1(n6051), .B2(n6050), .C1(n3915), 
        .C2(n6057), .ZN(n6052) );
  MUX2_X1 U7091 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n6052), .S(n6658), 
        .Z(U3465) );
  OAI211_X1 U7092 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6203), .A(n6664), .B(
        n6663), .ZN(n6053) );
  OAI21_X1 U7093 ( .B1(n6054), .B2(n6057), .A(n6053), .ZN(n6055) );
  MUX2_X1 U7094 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n6055), .S(n6658), 
        .Z(U3464) );
  XNOR2_X1 U7095 ( .A(n6056), .B(n6664), .ZN(n6058) );
  OAI22_X1 U7096 ( .A1(n6058), .A2(n6804), .B1(n6455), .B2(n6057), .ZN(n6059)
         );
  MUX2_X1 U7097 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n6059), .S(n6658), 
        .Z(U3463) );
  INV_X1 U7098 ( .A(n6060), .ZN(n6064) );
  OAI22_X1 U7099 ( .A1(n6064), .A2(n6063), .B1(n6062), .B2(n6061), .ZN(n6066)
         );
  MUX2_X1 U7100 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6066), .S(n6065), 
        .Z(U3456) );
  INV_X1 U7101 ( .A(n6072), .ZN(n6067) );
  OAI21_X1 U7102 ( .B1(n6067), .B2(n6361), .A(n6663), .ZN(n6078) );
  INV_X1 U7103 ( .A(n6078), .ZN(n6070) );
  NAND2_X1 U7104 ( .A1(n6068), .A2(n6667), .ZN(n6069) );
  NAND2_X1 U7105 ( .A1(n6074), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6073) );
  NAND2_X1 U7106 ( .A1(n6069), .A2(n6073), .ZN(n6077) );
  AND2_X1 U7107 ( .A1(n6072), .A2(n6071), .ZN(n6109) );
  INV_X1 U7108 ( .A(n6073), .ZN(n6101) );
  INV_X1 U7109 ( .A(n6074), .ZN(n6075) );
  AOI21_X1 U7110 ( .B1(n6804), .B2(n6075), .A(n6164), .ZN(n6076) );
  AOI22_X1 U7111 ( .A1(n3171), .A2(n6101), .B1(INSTQUEUE_REG_1__0__SCAN_IN), 
        .B2(n6100), .ZN(n6079) );
  OAI21_X1 U7112 ( .B1(n6103), .B2(n6679), .A(n6079), .ZN(n6080) );
  AOI21_X1 U7113 ( .B1(n6308), .B2(n6109), .A(n6080), .ZN(n6081) );
  OAI21_X1 U7114 ( .B1(n6106), .B2(n6306), .A(n6081), .ZN(U3028) );
  AOI22_X1 U7115 ( .A1(n6172), .A2(n6101), .B1(INSTQUEUE_REG_1__1__SCAN_IN), 
        .B2(n6100), .ZN(n6082) );
  OAI21_X1 U7116 ( .B1(n6103), .B2(n6681), .A(n6082), .ZN(n6083) );
  AOI21_X1 U7117 ( .B1(n6322), .B2(n6109), .A(n6083), .ZN(n6084) );
  OAI21_X1 U7118 ( .B1(n6106), .B2(n6320), .A(n6084), .ZN(U3029) );
  AOI22_X1 U7119 ( .A1(n3152), .A2(n6101), .B1(INSTQUEUE_REG_1__2__SCAN_IN), 
        .B2(n6100), .ZN(n6085) );
  OAI21_X1 U7120 ( .B1(n6103), .B2(n6693), .A(n6085), .ZN(n6086) );
  AOI21_X1 U7121 ( .B1(n6327), .B2(n6109), .A(n6086), .ZN(n6087) );
  OAI21_X1 U7122 ( .B1(n6106), .B2(n6325), .A(n6087), .ZN(U3030) );
  AOI22_X1 U7123 ( .A1(n6179), .A2(n6101), .B1(INSTQUEUE_REG_1__3__SCAN_IN), 
        .B2(n6100), .ZN(n6088) );
  OAI21_X1 U7124 ( .B1(n6103), .B2(n6695), .A(n6088), .ZN(n6089) );
  AOI21_X1 U7125 ( .B1(n6332), .B2(n6109), .A(n6089), .ZN(n6090) );
  OAI21_X1 U7126 ( .B1(n6106), .B2(n6330), .A(n6090), .ZN(U3031) );
  AOI22_X1 U7127 ( .A1(n6183), .A2(n6101), .B1(INSTQUEUE_REG_1__4__SCAN_IN), 
        .B2(n6100), .ZN(n6091) );
  OAI21_X1 U7128 ( .B1(n6103), .B2(n6707), .A(n6091), .ZN(n6092) );
  AOI21_X1 U7129 ( .B1(n6337), .B2(n6109), .A(n6092), .ZN(n6093) );
  OAI21_X1 U7130 ( .B1(n6106), .B2(n6335), .A(n6093), .ZN(U3032) );
  AOI22_X1 U7131 ( .A1(n6187), .A2(n6101), .B1(INSTQUEUE_REG_1__5__SCAN_IN), 
        .B2(n6100), .ZN(n6094) );
  OAI21_X1 U7132 ( .B1(n6103), .B2(n6714), .A(n6094), .ZN(n6095) );
  AOI21_X1 U7133 ( .B1(n6342), .B2(n6109), .A(n6095), .ZN(n6096) );
  OAI21_X1 U7134 ( .B1(n6106), .B2(n6340), .A(n6096), .ZN(U3033) );
  AOI22_X1 U7135 ( .A1(n6191), .A2(n6101), .B1(INSTQUEUE_REG_1__6__SCAN_IN), 
        .B2(n6100), .ZN(n6097) );
  OAI21_X1 U7136 ( .B1(n6103), .B2(n6721), .A(n6097), .ZN(n6098) );
  AOI21_X1 U7137 ( .B1(n6347), .B2(n6109), .A(n6098), .ZN(n6099) );
  OAI21_X1 U7138 ( .B1(n6106), .B2(n6345), .A(n6099), .ZN(U3034) );
  AOI22_X1 U7139 ( .A1(n6197), .A2(n6101), .B1(INSTQUEUE_REG_1__7__SCAN_IN), 
        .B2(n6100), .ZN(n6102) );
  OAI21_X1 U7140 ( .B1(n6103), .B2(n6733), .A(n6102), .ZN(n6104) );
  AOI21_X1 U7141 ( .B1(n6355), .B2(n6109), .A(n6104), .ZN(n6105) );
  OAI21_X1 U7142 ( .B1(n6106), .B2(n6351), .A(n6105), .ZN(U3035) );
  OAI21_X1 U7143 ( .B1(n6109), .B2(n6142), .A(n6108), .ZN(n6110) );
  AOI21_X1 U7144 ( .B1(n6110), .B2(n6113), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n6112) );
  NOR2_X1 U7145 ( .A1(n6111), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6116)
         );
  NAND2_X1 U7146 ( .A1(n6138), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n6119) );
  INV_X1 U7147 ( .A(n6113), .ZN(n6115) );
  NOR3_X1 U7148 ( .A1(n6315), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6301), 
        .ZN(n6114) );
  AOI21_X1 U7149 ( .B1(n6115), .B2(n6663), .A(n6114), .ZN(n6140) );
  INV_X1 U7150 ( .A(n6116), .ZN(n6139) );
  OAI22_X1 U7151 ( .A1(n6140), .A2(n6306), .B1(n6660), .B2(n6139), .ZN(n6117)
         );
  AOI21_X1 U7152 ( .B1(n6142), .B2(n6308), .A(n6117), .ZN(n6118) );
  OAI211_X1 U7153 ( .C1(n6145), .C2(n6679), .A(n6119), .B(n6118), .ZN(U3036)
         );
  NAND2_X1 U7154 ( .A1(n6138), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n6122) );
  OAI22_X1 U7155 ( .A1(n6140), .A2(n6320), .B1(n6680), .B2(n6139), .ZN(n6120)
         );
  AOI21_X1 U7156 ( .B1(n6142), .B2(n6322), .A(n6120), .ZN(n6121) );
  OAI211_X1 U7157 ( .C1(n6145), .C2(n6681), .A(n6122), .B(n6121), .ZN(U3037)
         );
  NAND2_X1 U7158 ( .A1(n6138), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n6125) );
  OAI22_X1 U7159 ( .A1(n6140), .A2(n6325), .B1(n6687), .B2(n6139), .ZN(n6123)
         );
  AOI21_X1 U7160 ( .B1(n6142), .B2(n6327), .A(n6123), .ZN(n6124) );
  OAI211_X1 U7161 ( .C1(n6145), .C2(n6693), .A(n6125), .B(n6124), .ZN(U3038)
         );
  NAND2_X1 U7162 ( .A1(n6138), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n6128) );
  OAI22_X1 U7163 ( .A1(n6140), .A2(n6330), .B1(n6694), .B2(n6139), .ZN(n6126)
         );
  AOI21_X1 U7164 ( .B1(n6142), .B2(n6332), .A(n6126), .ZN(n6127) );
  OAI211_X1 U7165 ( .C1(n6145), .C2(n6695), .A(n6128), .B(n6127), .ZN(U3039)
         );
  NAND2_X1 U7166 ( .A1(n6138), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n6131) );
  OAI22_X1 U7167 ( .A1(n6140), .A2(n6335), .B1(n6701), .B2(n6139), .ZN(n6129)
         );
  AOI21_X1 U7168 ( .B1(n6142), .B2(n6337), .A(n6129), .ZN(n6130) );
  OAI211_X1 U7169 ( .C1(n6145), .C2(n6707), .A(n6131), .B(n6130), .ZN(U3040)
         );
  NAND2_X1 U7170 ( .A1(n6138), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n6134) );
  OAI22_X1 U7171 ( .A1(n6140), .A2(n6340), .B1(n6708), .B2(n6139), .ZN(n6132)
         );
  AOI21_X1 U7172 ( .B1(n6142), .B2(n6342), .A(n6132), .ZN(n6133) );
  OAI211_X1 U7173 ( .C1(n6145), .C2(n6714), .A(n6134), .B(n6133), .ZN(U3041)
         );
  NAND2_X1 U7174 ( .A1(n6138), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n6137) );
  OAI22_X1 U7175 ( .A1(n6140), .A2(n6345), .B1(n6715), .B2(n6139), .ZN(n6135)
         );
  AOI21_X1 U7176 ( .B1(n6142), .B2(n6347), .A(n6135), .ZN(n6136) );
  OAI211_X1 U7177 ( .C1(n6145), .C2(n6721), .A(n6137), .B(n6136), .ZN(U3042)
         );
  NAND2_X1 U7178 ( .A1(n6138), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n6144) );
  OAI22_X1 U7179 ( .A1(n6140), .A2(n6351), .B1(n6723), .B2(n6139), .ZN(n6141)
         );
  AOI21_X1 U7180 ( .B1(n6142), .B2(n6355), .A(n6141), .ZN(n6143) );
  OAI211_X1 U7181 ( .C1(n6145), .C2(n6733), .A(n6144), .B(n6143), .ZN(U3043)
         );
  NAND2_X1 U7182 ( .A1(n6146), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n6155) );
  AOI22_X1 U7183 ( .A1(n6676), .A2(n6148), .B1(n3171), .B2(n6147), .ZN(n6154)
         );
  NAND2_X1 U7184 ( .A1(n6150), .A2(n6149), .ZN(n6153) );
  NAND2_X1 U7185 ( .A1(n6151), .A2(n6308), .ZN(n6152) );
  NAND4_X1 U7186 ( .A1(n6155), .A2(n6154), .A3(n6153), .A4(n6152), .ZN(U3068)
         );
  NAND2_X1 U7187 ( .A1(n6156), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6157) );
  OAI21_X1 U7188 ( .B1(n6665), .B2(n6157), .A(n6663), .ZN(n6168) );
  INV_X1 U7189 ( .A(n6168), .ZN(n6162) );
  NAND2_X1 U7190 ( .A1(n6159), .A2(n6158), .ZN(n6160) );
  OR2_X1 U7191 ( .A1(n6165), .A2(n6304), .ZN(n6163) );
  NAND2_X1 U7192 ( .A1(n6160), .A2(n6163), .ZN(n6167) );
  INV_X1 U7193 ( .A(n6165), .ZN(n6161) );
  NOR3_X2 U7194 ( .A1(n6665), .A2(n3912), .A3(n6203), .ZN(n6216) );
  INV_X1 U7195 ( .A(n6163), .ZN(n6196) );
  AOI21_X1 U7196 ( .B1(n6804), .B2(n6165), .A(n6164), .ZN(n6166) );
  OAI21_X1 U7197 ( .B1(n6168), .B2(n6167), .A(n6166), .ZN(n6195) );
  AOI22_X1 U7198 ( .A1(n3171), .A2(n6196), .B1(INSTQUEUE_REG_9__0__SCAN_IN), 
        .B2(n6195), .ZN(n6169) );
  OAI21_X1 U7199 ( .B1(n6199), .B2(n6679), .A(n6169), .ZN(n6170) );
  AOI21_X1 U7200 ( .B1(n6216), .B2(n6308), .A(n6170), .ZN(n6171) );
  OAI21_X1 U7201 ( .B1(n6202), .B2(n6306), .A(n6171), .ZN(U3092) );
  AOI22_X1 U7202 ( .A1(n6172), .A2(n6196), .B1(INSTQUEUE_REG_9__1__SCAN_IN), 
        .B2(n6195), .ZN(n6173) );
  OAI21_X1 U7203 ( .B1(n6199), .B2(n6681), .A(n6173), .ZN(n6174) );
  AOI21_X1 U7204 ( .B1(n6216), .B2(n6322), .A(n6174), .ZN(n6175) );
  OAI21_X1 U7205 ( .B1(n6202), .B2(n6320), .A(n6175), .ZN(U3093) );
  AOI22_X1 U7206 ( .A1(n3152), .A2(n6196), .B1(INSTQUEUE_REG_9__2__SCAN_IN), 
        .B2(n6195), .ZN(n6176) );
  OAI21_X1 U7207 ( .B1(n6199), .B2(n6693), .A(n6176), .ZN(n6177) );
  AOI21_X1 U7208 ( .B1(n6216), .B2(n6327), .A(n6177), .ZN(n6178) );
  OAI21_X1 U7209 ( .B1(n6202), .B2(n6325), .A(n6178), .ZN(U3094) );
  AOI22_X1 U7210 ( .A1(n6179), .A2(n6196), .B1(INSTQUEUE_REG_9__3__SCAN_IN), 
        .B2(n6195), .ZN(n6180) );
  OAI21_X1 U7211 ( .B1(n6199), .B2(n6695), .A(n6180), .ZN(n6181) );
  AOI21_X1 U7212 ( .B1(n6216), .B2(n6332), .A(n6181), .ZN(n6182) );
  OAI21_X1 U7213 ( .B1(n6202), .B2(n6330), .A(n6182), .ZN(U3095) );
  AOI22_X1 U7214 ( .A1(n6183), .A2(n6196), .B1(INSTQUEUE_REG_9__4__SCAN_IN), 
        .B2(n6195), .ZN(n6184) );
  OAI21_X1 U7215 ( .B1(n6199), .B2(n6707), .A(n6184), .ZN(n6185) );
  AOI21_X1 U7216 ( .B1(n6216), .B2(n6337), .A(n6185), .ZN(n6186) );
  OAI21_X1 U7217 ( .B1(n6202), .B2(n6335), .A(n6186), .ZN(U3096) );
  AOI22_X1 U7218 ( .A1(n6187), .A2(n6196), .B1(INSTQUEUE_REG_9__5__SCAN_IN), 
        .B2(n6195), .ZN(n6188) );
  OAI21_X1 U7219 ( .B1(n6199), .B2(n6714), .A(n6188), .ZN(n6189) );
  AOI21_X1 U7220 ( .B1(n6216), .B2(n6342), .A(n6189), .ZN(n6190) );
  OAI21_X1 U7221 ( .B1(n6202), .B2(n6340), .A(n6190), .ZN(U3097) );
  AOI22_X1 U7222 ( .A1(n6191), .A2(n6196), .B1(INSTQUEUE_REG_9__6__SCAN_IN), 
        .B2(n6195), .ZN(n6192) );
  OAI21_X1 U7223 ( .B1(n6199), .B2(n6721), .A(n6192), .ZN(n6193) );
  AOI21_X1 U7224 ( .B1(n6216), .B2(n6347), .A(n6193), .ZN(n6194) );
  OAI21_X1 U7225 ( .B1(n6202), .B2(n6345), .A(n6194), .ZN(U3098) );
  AOI22_X1 U7226 ( .A1(n6197), .A2(n6196), .B1(INSTQUEUE_REG_9__7__SCAN_IN), 
        .B2(n6195), .ZN(n6198) );
  OAI21_X1 U7227 ( .B1(n6199), .B2(n6733), .A(n6198), .ZN(n6200) );
  AOI21_X1 U7228 ( .B1(n6216), .B2(n6355), .A(n6200), .ZN(n6201) );
  OAI21_X1 U7229 ( .B1(n6202), .B2(n6351), .A(n6201), .ZN(U3099) );
  NAND2_X1 U7230 ( .A1(n6203), .A2(n3912), .ZN(n6204) );
  OAI21_X1 U7231 ( .B1(n6216), .B2(n6242), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6205) );
  NAND2_X1 U7232 ( .A1(n6205), .A2(n6663), .ZN(n6215) );
  INV_X1 U7233 ( .A(n6215), .ZN(n6209) );
  AND2_X1 U7234 ( .A1(n6207), .A2(n6206), .ZN(n6668) );
  NOR3_X1 U7235 ( .A1(n6315), .A2(n6301), .A3(n6302), .ZN(n6208) );
  AND2_X1 U7236 ( .A1(n6210), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6671)
         );
  NAND2_X1 U7237 ( .A1(n6671), .A2(n6304), .ZN(n6239) );
  NAND2_X1 U7238 ( .A1(n6302), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6211) );
  NAND2_X1 U7239 ( .A1(n6212), .A2(n6211), .ZN(n6313) );
  AOI211_X1 U7240 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6239), .A(n6213), .B(
        n6313), .ZN(n6214) );
  NAND2_X1 U7241 ( .A1(n6238), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n6219)
         );
  INV_X1 U7242 ( .A(n6216), .ZN(n6240) );
  OAI22_X1 U7243 ( .A1(n6240), .A2(n6679), .B1(n6660), .B2(n6239), .ZN(n6217)
         );
  AOI21_X1 U7244 ( .B1(n6308), .B2(n6242), .A(n6217), .ZN(n6218) );
  OAI211_X1 U7245 ( .C1(n6245), .C2(n6306), .A(n6219), .B(n6218), .ZN(U3100)
         );
  NAND2_X1 U7246 ( .A1(n6238), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n6222)
         );
  OAI22_X1 U7247 ( .A1(n6240), .A2(n6681), .B1(n6680), .B2(n6239), .ZN(n6220)
         );
  AOI21_X1 U7248 ( .B1(n6322), .B2(n6242), .A(n6220), .ZN(n6221) );
  OAI211_X1 U7249 ( .C1(n6245), .C2(n6320), .A(n6222), .B(n6221), .ZN(U3101)
         );
  NAND2_X1 U7250 ( .A1(n6238), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n6225)
         );
  OAI22_X1 U7251 ( .A1(n6240), .A2(n6693), .B1(n6687), .B2(n6239), .ZN(n6223)
         );
  AOI21_X1 U7252 ( .B1(n6327), .B2(n6242), .A(n6223), .ZN(n6224) );
  OAI211_X1 U7253 ( .C1(n6245), .C2(n6325), .A(n6225), .B(n6224), .ZN(U3102)
         );
  NAND2_X1 U7254 ( .A1(n6238), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n6228)
         );
  OAI22_X1 U7255 ( .A1(n6240), .A2(n6695), .B1(n6694), .B2(n6239), .ZN(n6226)
         );
  AOI21_X1 U7256 ( .B1(n6332), .B2(n6242), .A(n6226), .ZN(n6227) );
  OAI211_X1 U7257 ( .C1(n6245), .C2(n6330), .A(n6228), .B(n6227), .ZN(U3103)
         );
  NAND2_X1 U7258 ( .A1(n6238), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n6231)
         );
  OAI22_X1 U7259 ( .A1(n6240), .A2(n6707), .B1(n6701), .B2(n6239), .ZN(n6229)
         );
  AOI21_X1 U7260 ( .B1(n6337), .B2(n6242), .A(n6229), .ZN(n6230) );
  OAI211_X1 U7261 ( .C1(n6245), .C2(n6335), .A(n6231), .B(n6230), .ZN(U3104)
         );
  NAND2_X1 U7262 ( .A1(n6238), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n6234)
         );
  OAI22_X1 U7263 ( .A1(n6240), .A2(n6714), .B1(n6708), .B2(n6239), .ZN(n6232)
         );
  AOI21_X1 U7264 ( .B1(n6342), .B2(n6242), .A(n6232), .ZN(n6233) );
  OAI211_X1 U7265 ( .C1(n6245), .C2(n6340), .A(n6234), .B(n6233), .ZN(U3105)
         );
  NAND2_X1 U7266 ( .A1(n6238), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n6237)
         );
  OAI22_X1 U7267 ( .A1(n6240), .A2(n6721), .B1(n6715), .B2(n6239), .ZN(n6235)
         );
  AOI21_X1 U7268 ( .B1(n6347), .B2(n6242), .A(n6235), .ZN(n6236) );
  OAI211_X1 U7269 ( .C1(n6245), .C2(n6345), .A(n6237), .B(n6236), .ZN(U3106)
         );
  NAND2_X1 U7270 ( .A1(n6238), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n6244)
         );
  OAI22_X1 U7271 ( .A1(n6240), .A2(n6733), .B1(n6723), .B2(n6239), .ZN(n6241)
         );
  AOI21_X1 U7272 ( .B1(n6355), .B2(n6242), .A(n6241), .ZN(n6243) );
  OAI211_X1 U7273 ( .C1(n6245), .C2(n6351), .A(n6244), .B(n6243), .ZN(U3107)
         );
  INV_X1 U7274 ( .A(n6246), .ZN(n6247) );
  OR2_X1 U7275 ( .A1(n6248), .A2(n6312), .ZN(n6252) );
  NAND2_X1 U7276 ( .A1(n6250), .A2(n6249), .ZN(n6251) );
  NAND2_X1 U7277 ( .A1(n6252), .A2(n6251), .ZN(n6298) );
  NOR2_X1 U7278 ( .A1(n6253), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6261)
         );
  INV_X1 U7279 ( .A(n6261), .ZN(n6294) );
  INV_X1 U7280 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n6264) );
  INV_X1 U7281 ( .A(n6295), .ZN(n6255) );
  INV_X1 U7282 ( .A(n6725), .ZN(n6254) );
  OAI21_X1 U7283 ( .B1(n6255), .B2(n6254), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6256) );
  OAI211_X1 U7284 ( .C1(n6312), .C2(n6257), .A(n6663), .B(n6256), .ZN(n6258)
         );
  OAI211_X1 U7285 ( .C1(n6261), .C2(n6260), .A(n6259), .B(n6258), .ZN(n6263)
         );
  OAI22_X1 U7286 ( .A1(n6660), .A2(n6294), .B1(n6264), .B2(n6292), .ZN(n6266)
         );
  NOR2_X1 U7287 ( .A1(n6295), .A2(n6661), .ZN(n6265) );
  AOI211_X1 U7288 ( .C1(n6676), .C2(n6298), .A(n6266), .B(n6265), .ZN(n6267)
         );
  OAI21_X1 U7289 ( .B1(n6679), .B2(n6725), .A(n6267), .ZN(U3116) );
  INV_X1 U7290 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n6268) );
  OAI22_X1 U7291 ( .A1(n6680), .A2(n6294), .B1(n6268), .B2(n6292), .ZN(n6270)
         );
  NOR2_X1 U7292 ( .A1(n6295), .A2(n6686), .ZN(n6269) );
  AOI211_X1 U7293 ( .C1(n6683), .C2(n6298), .A(n6270), .B(n6269), .ZN(n6271)
         );
  OAI21_X1 U7294 ( .B1(n6681), .B2(n6725), .A(n6271), .ZN(U3117) );
  INV_X1 U7295 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n6272) );
  OAI22_X1 U7296 ( .A1(n6687), .A2(n6294), .B1(n6272), .B2(n6292), .ZN(n6274)
         );
  NOR2_X1 U7297 ( .A1(n6295), .A2(n6688), .ZN(n6273) );
  AOI211_X1 U7298 ( .C1(n6690), .C2(n6298), .A(n6274), .B(n6273), .ZN(n6275)
         );
  OAI21_X1 U7299 ( .B1(n6693), .B2(n6725), .A(n6275), .ZN(U3118) );
  INV_X1 U7300 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n6276) );
  OAI22_X1 U7301 ( .A1(n6694), .A2(n6294), .B1(n6276), .B2(n6292), .ZN(n6278)
         );
  NOR2_X1 U7302 ( .A1(n6295), .A2(n6700), .ZN(n6277) );
  AOI211_X1 U7303 ( .C1(n6697), .C2(n6298), .A(n6278), .B(n6277), .ZN(n6279)
         );
  OAI21_X1 U7304 ( .B1(n6695), .B2(n6725), .A(n6279), .ZN(U3119) );
  INV_X1 U7305 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n6280) );
  OAI22_X1 U7306 ( .A1(n6701), .A2(n6294), .B1(n6280), .B2(n6292), .ZN(n6282)
         );
  NOR2_X1 U7307 ( .A1(n6295), .A2(n6702), .ZN(n6281) );
  AOI211_X1 U7308 ( .C1(n6704), .C2(n6298), .A(n6282), .B(n6281), .ZN(n6283)
         );
  OAI21_X1 U7309 ( .B1(n6707), .B2(n6725), .A(n6283), .ZN(U3120) );
  INV_X1 U7310 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n6284) );
  OAI22_X1 U7311 ( .A1(n6708), .A2(n6294), .B1(n6284), .B2(n6292), .ZN(n6286)
         );
  NOR2_X1 U7312 ( .A1(n6295), .A2(n6709), .ZN(n6285) );
  AOI211_X1 U7313 ( .C1(n6711), .C2(n6298), .A(n6286), .B(n6285), .ZN(n6287)
         );
  OAI21_X1 U7314 ( .B1(n6714), .B2(n6725), .A(n6287), .ZN(U3121) );
  INV_X1 U7315 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n6288) );
  OAI22_X1 U7316 ( .A1(n6715), .A2(n6294), .B1(n6288), .B2(n6292), .ZN(n6290)
         );
  NOR2_X1 U7317 ( .A1(n6295), .A2(n6716), .ZN(n6289) );
  AOI211_X1 U7318 ( .C1(n6718), .C2(n6298), .A(n6290), .B(n6289), .ZN(n6291)
         );
  OAI21_X1 U7319 ( .B1(n6721), .B2(n6725), .A(n6291), .ZN(U3122) );
  INV_X1 U7320 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n6293) );
  OAI22_X1 U7321 ( .A1(n6723), .A2(n6294), .B1(n6293), .B2(n6292), .ZN(n6297)
         );
  NOR2_X1 U7322 ( .A1(n6295), .A2(n6724), .ZN(n6296) );
  AOI211_X1 U7323 ( .C1(n6728), .C2(n6298), .A(n6297), .B(n6296), .ZN(n6299)
         );
  OAI21_X1 U7324 ( .B1(n6733), .B2(n6725), .A(n6299), .ZN(U3123) );
  OAI33_X1 U7325 ( .A1(n6302), .A2(n6301), .A3(n6300), .B1(n6311), .B2(n6804), 
        .B3(n6312), .ZN(n6303) );
  INV_X1 U7326 ( .A(n6303), .ZN(n6352) );
  NAND2_X1 U7327 ( .A1(n6305), .A2(n6304), .ZN(n6350) );
  OAI22_X1 U7328 ( .A1(n6352), .A2(n6306), .B1(n6660), .B2(n6350), .ZN(n6307)
         );
  AOI21_X1 U7329 ( .B1(n6308), .B2(n6354), .A(n6307), .ZN(n6319) );
  OAI21_X1 U7330 ( .B1(n6354), .B2(n6309), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6310) );
  OAI211_X1 U7331 ( .C1(n6312), .C2(n6311), .A(n6310), .B(n6663), .ZN(n6317)
         );
  INV_X1 U7332 ( .A(n6313), .ZN(n6316) );
  NAND2_X1 U7333 ( .A1(n6350), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6314) );
  NAND4_X1 U7334 ( .A1(n6317), .A2(n6316), .A3(n6315), .A4(n6314), .ZN(n6356)
         );
  NAND2_X1 U7335 ( .A1(n6356), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n6318)
         );
  OAI211_X1 U7336 ( .C1(n6679), .C2(n6359), .A(n6319), .B(n6318), .ZN(U3132)
         );
  OAI22_X1 U7337 ( .A1(n6352), .A2(n6320), .B1(n6680), .B2(n6350), .ZN(n6321)
         );
  AOI21_X1 U7338 ( .B1(n6322), .B2(n6354), .A(n6321), .ZN(n6324) );
  NAND2_X1 U7339 ( .A1(n6356), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n6323)
         );
  OAI211_X1 U7340 ( .C1(n6681), .C2(n6359), .A(n6324), .B(n6323), .ZN(U3133)
         );
  OAI22_X1 U7341 ( .A1(n6352), .A2(n6325), .B1(n6687), .B2(n6350), .ZN(n6326)
         );
  AOI21_X1 U7342 ( .B1(n6327), .B2(n6354), .A(n6326), .ZN(n6329) );
  NAND2_X1 U7343 ( .A1(n6356), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n6328)
         );
  OAI211_X1 U7344 ( .C1(n6693), .C2(n6359), .A(n6329), .B(n6328), .ZN(U3134)
         );
  OAI22_X1 U7345 ( .A1(n6352), .A2(n6330), .B1(n6694), .B2(n6350), .ZN(n6331)
         );
  AOI21_X1 U7346 ( .B1(n6332), .B2(n6354), .A(n6331), .ZN(n6334) );
  NAND2_X1 U7347 ( .A1(n6356), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n6333)
         );
  OAI211_X1 U7348 ( .C1(n6695), .C2(n6359), .A(n6334), .B(n6333), .ZN(U3135)
         );
  OAI22_X1 U7349 ( .A1(n6352), .A2(n6335), .B1(n6701), .B2(n6350), .ZN(n6336)
         );
  AOI21_X1 U7350 ( .B1(n6337), .B2(n6354), .A(n6336), .ZN(n6339) );
  NAND2_X1 U7351 ( .A1(n6356), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n6338)
         );
  OAI211_X1 U7352 ( .C1(n6707), .C2(n6359), .A(n6339), .B(n6338), .ZN(U3136)
         );
  OAI22_X1 U7353 ( .A1(n6352), .A2(n6340), .B1(n6708), .B2(n6350), .ZN(n6341)
         );
  AOI21_X1 U7354 ( .B1(n6342), .B2(n6354), .A(n6341), .ZN(n6344) );
  NAND2_X1 U7355 ( .A1(n6356), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n6343)
         );
  OAI211_X1 U7356 ( .C1(n6714), .C2(n6359), .A(n6344), .B(n6343), .ZN(U3137)
         );
  OAI22_X1 U7357 ( .A1(n6352), .A2(n6345), .B1(n6715), .B2(n6350), .ZN(n6346)
         );
  AOI21_X1 U7358 ( .B1(n6347), .B2(n6354), .A(n6346), .ZN(n6349) );
  NAND2_X1 U7359 ( .A1(n6356), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n6348)
         );
  OAI211_X1 U7360 ( .C1(n6721), .C2(n6359), .A(n6349), .B(n6348), .ZN(U3138)
         );
  OAI22_X1 U7361 ( .A1(n6352), .A2(n6351), .B1(n6723), .B2(n6350), .ZN(n6353)
         );
  AOI21_X1 U7362 ( .B1(n6355), .B2(n6354), .A(n6353), .ZN(n6358) );
  NAND2_X1 U7363 ( .A1(n6356), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n6357)
         );
  OAI211_X1 U7364 ( .C1(n6733), .C2(n6359), .A(n6358), .B(n6357), .ZN(U3139)
         );
  MUX2_X1 U7365 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6780), .Z(U3447) );
  MUX2_X1 U7366 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6780), .Z(U3446) );
  INV_X1 U7367 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n7078) );
  NOR2_X1 U7368 ( .A1(n7078), .A2(n6506), .ZN(U2892) );
  OAI21_X1 U7369 ( .B1(n6360), .B2(BS16_N), .A(n6788), .ZN(n6787) );
  OAI21_X1 U7370 ( .B1(n6788), .B2(n6361), .A(n6787), .ZN(U2792) );
  OAI21_X1 U7371 ( .B1(n6363), .B2(n4525), .A(n6362), .ZN(U2793) );
  NOR4_X1 U7372 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_17__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n6948) );
  AOI211_X1 U7373 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_6__SCAN_IN), .B(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n6372) );
  NOR4_X1 U7374 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_8__SCAN_IN), .ZN(
        n6364) );
  INV_X1 U7375 ( .A(DATAWIDTH_REG_12__SCAN_IN), .ZN(n7010) );
  INV_X1 U7376 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n7038) );
  NAND3_X1 U7377 ( .A1(n6364), .A2(n7010), .A3(n7038), .ZN(n6370) );
  NOR4_X1 U7378 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_15__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n6368) );
  NOR4_X1 U7379 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(DATAWIDTH_REG_9__SCAN_IN), .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6367)
         );
  NOR4_X1 U7380 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(
        DATAWIDTH_REG_27__SCAN_IN), .A3(DATAWIDTH_REG_28__SCAN_IN), .A4(
        DATAWIDTH_REG_29__SCAN_IN), .ZN(n6366) );
  NOR4_X1 U7381 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6365) );
  NAND4_X1 U7382 ( .A1(n6368), .A2(n6367), .A3(n6366), .A4(n6365), .ZN(n6369)
         );
  NOR4_X1 U7383 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(DATAWIDTH_REG_2__SCAN_IN), .A3(n6370), .A4(n6369), .ZN(n6371) );
  NAND3_X1 U7384 ( .A1(n6948), .A2(n6372), .A3(n6371), .ZN(n6375) );
  INV_X1 U7385 ( .A(n6375), .ZN(n6796) );
  NAND2_X1 U7386 ( .A1(n6796), .A2(n7076), .ZN(n6791) );
  NOR3_X1 U7387 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(n6791), .ZN(n6374) );
  AOI21_X1 U7388 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(n6375), .A(n6374), .ZN(
        n6373) );
  OAI21_X1 U7389 ( .B1(n6792), .B2(n6375), .A(n6373), .ZN(U2794) );
  NAND2_X1 U7390 ( .A1(n6796), .A2(n6792), .ZN(n6789) );
  AOI21_X1 U7391 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(n6375), .A(n6374), .ZN(
        n6376) );
  OAI21_X1 U7392 ( .B1(DATAWIDTH_REG_1__SCAN_IN), .B2(n6789), .A(n6376), .ZN(
        U2795) );
  AOI22_X1 U7393 ( .A1(n6378), .A2(n3090), .B1(REIP_REG_12__SCAN_IN), .B2(
        n6377), .ZN(n6383) );
  INV_X1 U7394 ( .A(n6472), .ZN(n6381) );
  AOI22_X1 U7395 ( .A1(PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n6452), .B1(n6451), 
        .B2(n6469), .ZN(n6379) );
  OAI211_X1 U7396 ( .C1(n6467), .C2(n6475), .A(n6379), .B(n6442), .ZN(n6380)
         );
  AOI21_X1 U7397 ( .B1(n6381), .B2(n6422), .A(n6380), .ZN(n6382) );
  OAI211_X1 U7398 ( .C1(REIP_REG_12__SCAN_IN), .C2(n6384), .A(n6383), .B(n6382), .ZN(U2815) );
  AOI22_X1 U7399 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6441), .B1(n6385), .B2(n6427), .ZN(n6397) );
  NAND2_X1 U7400 ( .A1(n6387), .A2(n6386), .ZN(n6415) );
  INV_X1 U7401 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6756) );
  NAND2_X1 U7402 ( .A1(n6389), .A2(n6756), .ZN(n6400) );
  AOI21_X1 U7403 ( .B1(n6415), .B2(n6400), .A(n6965), .ZN(n6388) );
  INV_X1 U7404 ( .A(n6388), .ZN(n6395) );
  NAND3_X1 U7405 ( .A1(n6389), .A2(REIP_REG_9__SCAN_IN), .A3(n6965), .ZN(n6390) );
  NAND2_X1 U7406 ( .A1(n6442), .A2(n6390), .ZN(n6391) );
  AOI21_X1 U7407 ( .B1(n6452), .B2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6391), 
        .ZN(n6394) );
  NAND2_X1 U7408 ( .A1(n6392), .A2(n6422), .ZN(n6393) );
  AND3_X1 U7409 ( .A1(n6395), .A2(n6394), .A3(n6393), .ZN(n6396) );
  OAI211_X1 U7410 ( .C1(n6440), .C2(n6398), .A(n6397), .B(n6396), .ZN(U2817)
         );
  INV_X1 U7411 ( .A(EBX_REG_9__SCAN_IN), .ZN(n7028) );
  AOI22_X1 U7412 ( .A1(n6399), .A2(n6427), .B1(n6451), .B2(n6603), .ZN(n6406)
         );
  OAI211_X1 U7413 ( .C1(n6444), .C2(n6401), .A(n6442), .B(n6400), .ZN(n6404)
         );
  OAI22_X1 U7414 ( .A1(n6402), .A2(n6435), .B1(n6756), .B2(n6415), .ZN(n6403)
         );
  NOR2_X1 U7415 ( .A1(n6404), .A2(n6403), .ZN(n6405) );
  OAI211_X1 U7416 ( .C1(n7028), .C2(n6467), .A(n6406), .B(n6405), .ZN(U2818)
         );
  AOI21_X1 U7417 ( .B1(n6459), .B2(n6407), .A(REIP_REG_8__SCAN_IN), .ZN(n6416)
         );
  OAI22_X1 U7418 ( .A1(n6408), .A2(n6467), .B1(n6440), .B2(n6610), .ZN(n6409)
         );
  AOI211_X1 U7419 ( .C1(n6452), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6429), 
        .B(n6409), .ZN(n6414) );
  INV_X1 U7420 ( .A(n6410), .ZN(n6412) );
  AOI22_X1 U7421 ( .A1(n6412), .A2(n6422), .B1(n3090), .B2(n6411), .ZN(n6413)
         );
  OAI211_X1 U7422 ( .C1(n6416), .C2(n6415), .A(n6414), .B(n6413), .ZN(U2819)
         );
  NOR3_X1 U7423 ( .A1(n6424), .A2(REIP_REG_7__SCAN_IN), .A3(n6417), .ZN(n6421)
         );
  OAI22_X1 U7424 ( .A1(n6936), .A2(n6467), .B1(n6440), .B2(n6617), .ZN(n6418)
         );
  AOI211_X1 U7425 ( .C1(n6452), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6418), 
        .B(n6429), .ZN(n6419) );
  INV_X1 U7426 ( .A(n6419), .ZN(n6420) );
  AOI211_X1 U7427 ( .C1(n6566), .C2(n6422), .A(n6421), .B(n6420), .ZN(n6426)
         );
  OAI21_X1 U7428 ( .B1(n6424), .B2(n6430), .A(n6423), .ZN(n6446) );
  NOR2_X1 U7429 ( .A1(n6424), .A2(REIP_REG_6__SCAN_IN), .ZN(n6431) );
  OAI21_X1 U7430 ( .B1(n6446), .B2(n6431), .A(REIP_REG_7__SCAN_IN), .ZN(n6425)
         );
  OAI211_X1 U7431 ( .C1(n6462), .C2(n6569), .A(n6426), .B(n6425), .ZN(U2820)
         );
  AOI22_X1 U7432 ( .A1(EBX_REG_6__SCAN_IN), .A2(n6441), .B1(n6428), .B2(n3090), 
        .ZN(n6438) );
  AOI21_X1 U7433 ( .B1(n6452), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6429), 
        .ZN(n6433) );
  NAND2_X1 U7434 ( .A1(n6431), .A2(n6430), .ZN(n6432) );
  OAI211_X1 U7435 ( .C1(n6435), .C2(n6434), .A(n6433), .B(n6432), .ZN(n6436)
         );
  AOI21_X1 U7436 ( .B1(REIP_REG_6__SCAN_IN), .B2(n6446), .A(n6436), .ZN(n6437)
         );
  OAI211_X1 U7437 ( .C1(n6440), .C2(n6439), .A(n6438), .B(n6437), .ZN(U2821)
         );
  AOI22_X1 U7438 ( .A1(EBX_REG_5__SCAN_IN), .A2(n6441), .B1(n6451), .B2(n6626), 
        .ZN(n6443) );
  OAI211_X1 U7439 ( .C1(n6444), .C2(n3935), .A(n6443), .B(n6442), .ZN(n6445)
         );
  AOI21_X1 U7440 ( .B1(n6464), .B2(n6573), .A(n6445), .ZN(n6449) );
  OAI221_X1 U7441 ( .B1(REIP_REG_5__SCAN_IN), .B2(REIP_REG_4__SCAN_IN), .C1(
        REIP_REG_5__SCAN_IN), .C2(n6447), .A(n6446), .ZN(n6448) );
  OAI211_X1 U7442 ( .C1(n6462), .C2(n6576), .A(n6449), .B(n6448), .ZN(U2822)
         );
  NAND2_X1 U7443 ( .A1(n6451), .A2(n6450), .ZN(n6454) );
  NAND2_X1 U7444 ( .A1(n6452), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6453)
         );
  OAI211_X1 U7445 ( .C1(n6456), .C2(n6455), .A(n6454), .B(n6453), .ZN(n6457)
         );
  INV_X1 U7446 ( .A(n6457), .ZN(n6466) );
  AOI211_X1 U7447 ( .C1(n6459), .C2(n6792), .A(n6458), .B(n6746), .ZN(n6461)
         );
  AOI21_X1 U7448 ( .B1(n6459), .B2(REIP_REG_1__SCAN_IN), .A(
        REIP_REG_2__SCAN_IN), .ZN(n6460) );
  OAI22_X1 U7449 ( .A1(n6462), .A2(n6598), .B1(n6461), .B2(n6460), .ZN(n6463)
         );
  AOI21_X1 U7450 ( .B1(n6595), .B2(n6464), .A(n6463), .ZN(n6465) );
  OAI211_X1 U7451 ( .C1(n6468), .C2(n6467), .A(n6466), .B(n6465), .ZN(U2825)
         );
  INV_X1 U7452 ( .A(n6469), .ZN(n6470) );
  OAI22_X1 U7453 ( .A1(n6472), .A2(n6471), .B1(n6470), .B2(n5605), .ZN(n6473)
         );
  INV_X1 U7454 ( .A(n6473), .ZN(n6474) );
  OAI21_X1 U7455 ( .B1(n6475), .B2(n6480), .A(n6474), .ZN(U2847) );
  INV_X1 U7456 ( .A(n6476), .ZN(n6585) );
  AOI22_X1 U7457 ( .A1(n6585), .A2(n6478), .B1(n6477), .B2(n6650), .ZN(n6479)
         );
  OAI21_X1 U7458 ( .B1(n6992), .B2(n6480), .A(n6479), .ZN(U2856) );
  AOI22_X1 U7459 ( .A1(n6812), .A2(DATAO_REG_30__SCAN_IN), .B1(n6490), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n6482) );
  OAI21_X1 U7460 ( .B1(n6806), .B2(n7012), .A(n6482), .ZN(U2893) );
  INV_X1 U7461 ( .A(UWORD_REG_13__SCAN_IN), .ZN(n7056) );
  AOI22_X1 U7462 ( .A1(n6812), .A2(DATAO_REG_29__SCAN_IN), .B1(n6490), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n6483) );
  OAI21_X1 U7463 ( .B1(n6806), .B2(n7056), .A(n6483), .ZN(U2894) );
  INV_X1 U7464 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n7107) );
  AOI22_X1 U7465 ( .A1(n6490), .A2(EAX_REG_27__SCAN_IN), .B1(n6813), .B2(
        UWORD_REG_11__SCAN_IN), .ZN(n6484) );
  OAI21_X1 U7466 ( .B1(n7107), .B2(n6506), .A(n6484), .ZN(U2896) );
  INV_X1 U7467 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n7062) );
  AOI22_X1 U7468 ( .A1(n6490), .A2(EAX_REG_26__SCAN_IN), .B1(n6813), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n6485) );
  OAI21_X1 U7469 ( .B1(n7062), .B2(n6506), .A(n6485), .ZN(U2897) );
  INV_X1 U7470 ( .A(UWORD_REG_9__SCAN_IN), .ZN(n7091) );
  AOI22_X1 U7471 ( .A1(n6812), .A2(DATAO_REG_25__SCAN_IN), .B1(n6490), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n6486) );
  OAI21_X1 U7472 ( .B1(n6806), .B2(n7091), .A(n6486), .ZN(U2898) );
  INV_X1 U7473 ( .A(UWORD_REG_8__SCAN_IN), .ZN(n6888) );
  AOI22_X1 U7474 ( .A1(n6812), .A2(DATAO_REG_24__SCAN_IN), .B1(n6490), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n6487) );
  OAI21_X1 U7475 ( .B1(n6806), .B2(n6888), .A(n6487), .ZN(U2899) );
  INV_X1 U7476 ( .A(UWORD_REG_6__SCAN_IN), .ZN(n6898) );
  AOI22_X1 U7477 ( .A1(n6812), .A2(DATAO_REG_22__SCAN_IN), .B1(n6490), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n6488) );
  OAI21_X1 U7478 ( .B1(n6806), .B2(n6898), .A(n6488), .ZN(U2901) );
  INV_X1 U7479 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n7007) );
  AOI22_X1 U7480 ( .A1(n6490), .A2(EAX_REG_18__SCAN_IN), .B1(n6813), .B2(
        UWORD_REG_2__SCAN_IN), .ZN(n6489) );
  OAI21_X1 U7481 ( .B1(n7007), .B2(n6506), .A(n6489), .ZN(U2905) );
  INV_X1 U7482 ( .A(UWORD_REG_0__SCAN_IN), .ZN(n6945) );
  AOI22_X1 U7483 ( .A1(n6812), .A2(DATAO_REG_16__SCAN_IN), .B1(n6490), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6491) );
  OAI21_X1 U7484 ( .B1(n6806), .B2(n6945), .A(n6491), .ZN(U2907) );
  AOI22_X1 U7485 ( .A1(EAX_REG_15__SCAN_IN), .A2(n6814), .B1(n6812), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6492) );
  OAI21_X1 U7486 ( .B1(n6806), .B2(n6818), .A(n6492), .ZN(U2908) );
  INV_X1 U7487 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n7088) );
  INV_X1 U7488 ( .A(n6814), .ZN(n6512) );
  INV_X1 U7489 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6954) );
  INV_X1 U7490 ( .A(LWORD_REG_14__SCAN_IN), .ZN(n6493) );
  OAI222_X1 U7491 ( .A1(n6506), .A2(n7088), .B1(n6512), .B2(n6954), .C1(n6806), 
        .C2(n6493), .ZN(U2909) );
  AOI22_X1 U7492 ( .A1(n6813), .A2(LWORD_REG_13__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6494) );
  OAI21_X1 U7493 ( .B1(n6495), .B2(n6512), .A(n6494), .ZN(U2910) );
  INV_X1 U7494 ( .A(LWORD_REG_12__SCAN_IN), .ZN(n6903) );
  AOI22_X1 U7495 ( .A1(EAX_REG_12__SCAN_IN), .A2(n6814), .B1(n6812), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6496) );
  OAI21_X1 U7496 ( .B1(n6806), .B2(n6903), .A(n6496), .ZN(U2911) );
  AOI22_X1 U7497 ( .A1(n6813), .A2(LWORD_REG_10__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6497) );
  OAI21_X1 U7498 ( .B1(n7092), .B2(n6512), .A(n6497), .ZN(U2913) );
  AOI22_X1 U7499 ( .A1(n6813), .A2(LWORD_REG_9__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6498) );
  OAI21_X1 U7500 ( .B1(n7025), .B2(n6512), .A(n6498), .ZN(U2914) );
  INV_X1 U7501 ( .A(LWORD_REG_8__SCAN_IN), .ZN(n7016) );
  AOI22_X1 U7502 ( .A1(EAX_REG_8__SCAN_IN), .A2(n6814), .B1(n6812), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6499) );
  OAI21_X1 U7503 ( .B1(n6806), .B2(n7016), .A(n6499), .ZN(U2915) );
  INV_X1 U7504 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n7086) );
  INV_X1 U7505 ( .A(LWORD_REG_7__SCAN_IN), .ZN(n6500) );
  OAI222_X1 U7506 ( .A1(n6506), .A2(n7086), .B1(n6512), .B2(n6501), .C1(n6806), 
        .C2(n6500), .ZN(U2916) );
  INV_X1 U7507 ( .A(LWORD_REG_6__SCAN_IN), .ZN(n6955) );
  AOI22_X1 U7508 ( .A1(EAX_REG_6__SCAN_IN), .A2(n6814), .B1(n6812), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6502) );
  OAI21_X1 U7509 ( .B1(n6806), .B2(n6955), .A(n6502), .ZN(U2917) );
  INV_X1 U7510 ( .A(LWORD_REG_5__SCAN_IN), .ZN(n6994) );
  AOI22_X1 U7511 ( .A1(EAX_REG_5__SCAN_IN), .A2(n6814), .B1(n6812), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6503) );
  OAI21_X1 U7512 ( .B1(n6806), .B2(n6994), .A(n6503), .ZN(U2918) );
  INV_X1 U7513 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n7013) );
  INV_X1 U7514 ( .A(LWORD_REG_4__SCAN_IN), .ZN(n6504) );
  OAI222_X1 U7515 ( .A1(n6506), .A2(n7013), .B1(n6512), .B2(n6505), .C1(n6806), 
        .C2(n6504), .ZN(U2919) );
  AOI22_X1 U7516 ( .A1(n6813), .A2(LWORD_REG_3__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6507) );
  OAI21_X1 U7517 ( .B1(n7108), .B2(n6512), .A(n6507), .ZN(U2920) );
  AOI22_X1 U7518 ( .A1(n6813), .A2(LWORD_REG_2__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6508) );
  OAI21_X1 U7519 ( .B1(n6509), .B2(n6512), .A(n6508), .ZN(U2921) );
  INV_X1 U7520 ( .A(LWORD_REG_1__SCAN_IN), .ZN(n6909) );
  AOI22_X1 U7521 ( .A1(EAX_REG_1__SCAN_IN), .A2(n6814), .B1(n6812), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6510) );
  OAI21_X1 U7522 ( .B1(n6806), .B2(n6909), .A(n6510), .ZN(U2922) );
  AOI22_X1 U7523 ( .A1(n6813), .A2(LWORD_REG_0__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6511) );
  OAI21_X1 U7524 ( .B1(n6513), .B2(n6512), .A(n6511), .ZN(U2923) );
  AOI22_X1 U7525 ( .A1(UWORD_REG_0__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6514) );
  OAI21_X1 U7526 ( .B1(n6556), .B2(n6531), .A(n6514), .ZN(U2924) );
  AOI22_X1 U7527 ( .A1(UWORD_REG_1__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6515) );
  OAI21_X1 U7528 ( .B1(n6556), .B2(n6835), .A(n6515), .ZN(U2925) );
  AOI22_X1 U7529 ( .A1(UWORD_REG_2__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6516) );
  OAI21_X1 U7530 ( .B1(n6556), .B2(n6534), .A(n6516), .ZN(U2926) );
  AOI22_X1 U7531 ( .A1(UWORD_REG_3__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n6517) );
  OAI21_X1 U7532 ( .B1(n6556), .B2(n6536), .A(n6517), .ZN(U2927) );
  AOI22_X1 U7533 ( .A1(UWORD_REG_4__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6518) );
  OAI21_X1 U7534 ( .B1(n6556), .B2(n6538), .A(n6518), .ZN(U2928) );
  AOI22_X1 U7535 ( .A1(UWORD_REG_5__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n6519) );
  OAI21_X1 U7536 ( .B1(n6556), .B2(n6540), .A(n6519), .ZN(U2929) );
  AOI22_X1 U7537 ( .A1(UWORD_REG_6__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n6520) );
  OAI21_X1 U7538 ( .B1(n6556), .B2(n6542), .A(n6520), .ZN(U2930) );
  AOI22_X1 U7539 ( .A1(UWORD_REG_7__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n6521) );
  OAI21_X1 U7540 ( .B1(n6556), .B2(n6544), .A(n6521), .ZN(U2931) );
  AOI22_X1 U7541 ( .A1(UWORD_REG_8__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n6522) );
  OAI21_X1 U7542 ( .B1(n6556), .B2(n6848), .A(n6522), .ZN(U2932) );
  AOI22_X1 U7543 ( .A1(UWORD_REG_9__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n6524) );
  OAI21_X1 U7544 ( .B1(n6556), .B2(n6547), .A(n6524), .ZN(U2933) );
  AOI22_X1 U7545 ( .A1(UWORD_REG_10__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n6525) );
  OAI21_X1 U7546 ( .B1(n6556), .B2(n6549), .A(n6525), .ZN(U2934) );
  AOI22_X1 U7547 ( .A1(UWORD_REG_11__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n6527) );
  INV_X1 U7548 ( .A(n6556), .ZN(n6526) );
  NAND2_X1 U7549 ( .A1(n6526), .A2(DATAI_11_), .ZN(n6550) );
  NAND2_X1 U7550 ( .A1(n6527), .A2(n6550), .ZN(U2935) );
  AOI22_X1 U7551 ( .A1(UWORD_REG_12__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n6528) );
  OAI21_X1 U7552 ( .B1(n6556), .B2(n6949), .A(n6528), .ZN(U2936) );
  AOI22_X1 U7553 ( .A1(UWORD_REG_13__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n6529) );
  OAI21_X1 U7554 ( .B1(n6556), .B2(n6555), .A(n6529), .ZN(U2937) );
  AOI22_X1 U7555 ( .A1(LWORD_REG_0__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_0__SCAN_IN), .ZN(n6530) );
  OAI21_X1 U7556 ( .B1(n6556), .B2(n6531), .A(n6530), .ZN(U2939) );
  AOI22_X1 U7557 ( .A1(LWORD_REG_1__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_1__SCAN_IN), .ZN(n6532) );
  OAI21_X1 U7558 ( .B1(n6556), .B2(n6835), .A(n6532), .ZN(U2940) );
  AOI22_X1 U7559 ( .A1(LWORD_REG_2__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_2__SCAN_IN), .ZN(n6533) );
  OAI21_X1 U7560 ( .B1(n6556), .B2(n6534), .A(n6533), .ZN(U2941) );
  AOI22_X1 U7561 ( .A1(LWORD_REG_3__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_3__SCAN_IN), .ZN(n6535) );
  OAI21_X1 U7562 ( .B1(n6556), .B2(n6536), .A(n6535), .ZN(U2942) );
  AOI22_X1 U7563 ( .A1(LWORD_REG_4__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_4__SCAN_IN), .ZN(n6537) );
  OAI21_X1 U7564 ( .B1(n6556), .B2(n6538), .A(n6537), .ZN(U2943) );
  AOI22_X1 U7565 ( .A1(LWORD_REG_5__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_5__SCAN_IN), .ZN(n6539) );
  OAI21_X1 U7566 ( .B1(n6556), .B2(n6540), .A(n6539), .ZN(U2944) );
  AOI22_X1 U7567 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_6__SCAN_IN), .ZN(n6541) );
  OAI21_X1 U7568 ( .B1(n6556), .B2(n6542), .A(n6541), .ZN(U2945) );
  AOI22_X1 U7569 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n6543) );
  OAI21_X1 U7570 ( .B1(n6556), .B2(n6544), .A(n6543), .ZN(U2946) );
  AOI22_X1 U7571 ( .A1(LWORD_REG_8__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n6545) );
  OAI21_X1 U7572 ( .B1(n6556), .B2(n6848), .A(n6545), .ZN(U2947) );
  AOI22_X1 U7573 ( .A1(LWORD_REG_9__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n6546) );
  OAI21_X1 U7574 ( .B1(n6556), .B2(n6547), .A(n6546), .ZN(U2948) );
  AOI22_X1 U7575 ( .A1(LWORD_REG_10__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n6548) );
  OAI21_X1 U7576 ( .B1(n6556), .B2(n6549), .A(n6548), .ZN(U2949) );
  AOI22_X1 U7577 ( .A1(LWORD_REG_11__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n6551) );
  NAND2_X1 U7578 ( .A1(n6551), .A2(n6550), .ZN(U2950) );
  AOI22_X1 U7579 ( .A1(LWORD_REG_12__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n6552) );
  OAI21_X1 U7580 ( .B1(n6556), .B2(n6949), .A(n6552), .ZN(U2951) );
  AOI22_X1 U7581 ( .A1(LWORD_REG_13__SCAN_IN), .A2(n6557), .B1(n6553), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n6554) );
  OAI21_X1 U7582 ( .B1(n6556), .B2(n6555), .A(n6554), .ZN(U2952) );
  NAND2_X1 U7583 ( .A1(n6557), .A2(LWORD_REG_14__SCAN_IN), .ZN(n6558) );
  AND2_X1 U7584 ( .A1(n6559), .A2(n6558), .ZN(n6560) );
  OAI21_X1 U7585 ( .B1(n6954), .B2(n6561), .A(n6560), .ZN(U2953) );
  AOI22_X1 U7586 ( .A1(n6591), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .B1(n6577), 
        .B2(REIP_REG_7__SCAN_IN), .ZN(n6568) );
  NAND3_X1 U7587 ( .A1(n6563), .A2(n6562), .A3(n3124), .ZN(n6564) );
  AND2_X1 U7588 ( .A1(n6565), .A2(n6564), .ZN(n6619) );
  AOI22_X1 U7589 ( .A1(n6619), .A2(n6592), .B1(n6594), .B2(n6566), .ZN(n6567)
         );
  OAI211_X1 U7590 ( .C1(n6599), .C2(n6569), .A(n6568), .B(n6567), .ZN(U2979)
         );
  AND2_X1 U7591 ( .A1(n6577), .A2(REIP_REG_5__SCAN_IN), .ZN(n6625) );
  AOI21_X1 U7592 ( .B1(n6591), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n6625), 
        .ZN(n6575) );
  INV_X1 U7593 ( .A(n6572), .ZN(n6630) );
  AOI22_X1 U7594 ( .A1(n6630), .A2(n6592), .B1(n6594), .B2(n6573), .ZN(n6574)
         );
  OAI211_X1 U7595 ( .C1(n6599), .C2(n6576), .A(n6575), .B(n6574), .ZN(U2981)
         );
  AND2_X1 U7596 ( .A1(n6577), .A2(REIP_REG_3__SCAN_IN), .ZN(n6649) );
  AOI21_X1 U7597 ( .B1(n6591), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n6649), 
        .ZN(n6587) );
  INV_X1 U7598 ( .A(n4588), .ZN(n6580) );
  OAI21_X1 U7599 ( .B1(n6580), .B2(n6579), .A(n6578), .ZN(n6581) );
  OAI21_X1 U7600 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n4588), .A(n6581), 
        .ZN(n6584) );
  XNOR2_X1 U7601 ( .A(n3547), .B(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6583)
         );
  XNOR2_X1 U7602 ( .A(n6584), .B(n6583), .ZN(n6652) );
  AOI22_X1 U7603 ( .A1(n6594), .A2(n6585), .B1(n6652), .B2(n6592), .ZN(n6586)
         );
  OAI211_X1 U7604 ( .C1(n6599), .C2(n6588), .A(n6587), .B(n6586), .ZN(U2983)
         );
  INV_X1 U7605 ( .A(n6589), .ZN(n6590) );
  AOI21_X1 U7606 ( .B1(n6591), .B2(PHYADDRPOINTER_REG_2__SCAN_IN), .A(n6590), 
        .ZN(n6597) );
  AOI22_X1 U7607 ( .A1(n6595), .A2(n6594), .B1(n6593), .B2(n6592), .ZN(n6596)
         );
  OAI211_X1 U7608 ( .C1(n6599), .C2(n6598), .A(n6597), .B(n6596), .ZN(U2984)
         );
  INV_X1 U7609 ( .A(n6600), .ZN(n6608) );
  INV_X1 U7610 ( .A(n6601), .ZN(n6602) );
  AOI21_X1 U7611 ( .B1(n6603), .B2(n6651), .A(n6602), .ZN(n6607) );
  AOI22_X1 U7612 ( .A1(n6605), .A2(n6653), .B1(n6604), .B2(n7064), .ZN(n6606)
         );
  OAI211_X1 U7613 ( .C1(n6608), .C2(n7064), .A(n6607), .B(n6606), .ZN(U3009)
         );
  OAI22_X1 U7614 ( .A1(n6640), .A2(n6610), .B1(n6609), .B2(n6639), .ZN(n6613)
         );
  INV_X1 U7615 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6622) );
  AOI211_X1 U7616 ( .C1(n6622), .C2(n6616), .A(n6611), .B(n6623), .ZN(n6612)
         );
  AOI211_X1 U7617 ( .C1(n6614), .C2(n6653), .A(n6613), .B(n6612), .ZN(n6615)
         );
  OAI21_X1 U7618 ( .B1(n6621), .B2(n6616), .A(n6615), .ZN(U3010) );
  OAI22_X1 U7619 ( .A1(n6640), .A2(n6617), .B1(n6753), .B2(n6639), .ZN(n6618)
         );
  AOI21_X1 U7620 ( .B1(n6619), .B2(n6653), .A(n6618), .ZN(n6620) );
  OAI221_X1 U7621 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n6623), .C1(n6622), .C2(n6621), .A(n6620), .ZN(U3011) );
  AOI21_X1 U7622 ( .B1(n6636), .B2(n6624), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n6633) );
  AOI21_X1 U7623 ( .B1(n6651), .B2(n6626), .A(n6625), .ZN(n6632) );
  NOR3_X1 U7624 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6628), .A3(n6627), 
        .ZN(n6629) );
  AOI21_X1 U7625 ( .B1(n6630), .B2(n6653), .A(n6629), .ZN(n6631) );
  OAI211_X1 U7626 ( .C1(n6634), .C2(n6633), .A(n6632), .B(n6631), .ZN(U3013)
         );
  AOI21_X1 U7627 ( .B1(n6636), .B2(n6644), .A(n6635), .ZN(n6657) );
  OAI222_X1 U7628 ( .A1(n6641), .A2(n6640), .B1(n6639), .B2(n6748), .C1(n6638), 
        .C2(n6637), .ZN(n6642) );
  INV_X1 U7629 ( .A(n6642), .ZN(n6647) );
  NOR2_X1 U7630 ( .A1(n6644), .A2(n6643), .ZN(n6654) );
  OAI211_X1 U7631 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6654), .B(n6645), .ZN(n6646) );
  OAI211_X1 U7632 ( .C1(n6657), .C2(n6648), .A(n6647), .B(n6646), .ZN(U3014)
         );
  AOI21_X1 U7633 ( .B1(n6651), .B2(n6650), .A(n6649), .ZN(n6656) );
  AOI22_X1 U7634 ( .A1(n6654), .A2(n3522), .B1(n6653), .B2(n6652), .ZN(n6655)
         );
  OAI211_X1 U7635 ( .C1(n6657), .C2(n3522), .A(n6656), .B(n6655), .ZN(U3015)
         );
  NOR2_X1 U7636 ( .A1(n6659), .A2(n6658), .ZN(U3019) );
  AND2_X1 U7637 ( .A1(n6671), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6666)
         );
  INV_X1 U7638 ( .A(n6666), .ZN(n6722) );
  OAI22_X1 U7639 ( .A1(n6725), .A2(n6661), .B1(n6660), .B2(n6722), .ZN(n6662)
         );
  INV_X1 U7640 ( .A(n6662), .ZN(n6678) );
  OAI21_X1 U7641 ( .B1(n6665), .B2(n6664), .A(n6663), .ZN(n6675) );
  AOI21_X1 U7642 ( .B1(n6668), .B2(n6667), .A(n6666), .ZN(n6674) );
  INV_X1 U7643 ( .A(n6674), .ZN(n6670) );
  OAI211_X1 U7644 ( .C1(n6675), .C2(n6670), .A(n6669), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6729) );
  INV_X1 U7645 ( .A(n6671), .ZN(n6672) );
  OAI22_X1 U7646 ( .A1(n6675), .A2(n6674), .B1(n6673), .B2(n6672), .ZN(n6727)
         );
  AOI22_X1 U7647 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6729), .B1(n6676), 
        .B2(n6727), .ZN(n6677) );
  OAI211_X1 U7648 ( .C1(n6679), .C2(n6732), .A(n6678), .B(n6677), .ZN(U3108)
         );
  OAI22_X1 U7649 ( .A1(n6732), .A2(n6681), .B1(n6680), .B2(n6722), .ZN(n6682)
         );
  INV_X1 U7650 ( .A(n6682), .ZN(n6685) );
  AOI22_X1 U7651 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6729), .B1(n6683), 
        .B2(n6727), .ZN(n6684) );
  OAI211_X1 U7652 ( .C1(n6686), .C2(n6725), .A(n6685), .B(n6684), .ZN(U3109)
         );
  OAI22_X1 U7653 ( .A1(n6725), .A2(n6688), .B1(n6687), .B2(n6722), .ZN(n6689)
         );
  INV_X1 U7654 ( .A(n6689), .ZN(n6692) );
  AOI22_X1 U7655 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6729), .B1(n6690), 
        .B2(n6727), .ZN(n6691) );
  OAI211_X1 U7656 ( .C1(n6693), .C2(n6732), .A(n6692), .B(n6691), .ZN(U3110)
         );
  OAI22_X1 U7657 ( .A1(n6732), .A2(n6695), .B1(n6694), .B2(n6722), .ZN(n6696)
         );
  INV_X1 U7658 ( .A(n6696), .ZN(n6699) );
  AOI22_X1 U7659 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6729), .B1(n6697), 
        .B2(n6727), .ZN(n6698) );
  OAI211_X1 U7660 ( .C1(n6700), .C2(n6725), .A(n6699), .B(n6698), .ZN(U3111)
         );
  OAI22_X1 U7661 ( .A1(n6725), .A2(n6702), .B1(n6701), .B2(n6722), .ZN(n6703)
         );
  INV_X1 U7662 ( .A(n6703), .ZN(n6706) );
  AOI22_X1 U7663 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6729), .B1(n6704), 
        .B2(n6727), .ZN(n6705) );
  OAI211_X1 U7664 ( .C1(n6707), .C2(n6732), .A(n6706), .B(n6705), .ZN(U3112)
         );
  OAI22_X1 U7665 ( .A1(n6725), .A2(n6709), .B1(n6708), .B2(n6722), .ZN(n6710)
         );
  INV_X1 U7666 ( .A(n6710), .ZN(n6713) );
  AOI22_X1 U7667 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6729), .B1(n6711), 
        .B2(n6727), .ZN(n6712) );
  OAI211_X1 U7668 ( .C1(n6714), .C2(n6732), .A(n6713), .B(n6712), .ZN(U3113)
         );
  OAI22_X1 U7669 ( .A1(n6725), .A2(n6716), .B1(n6715), .B2(n6722), .ZN(n6717)
         );
  INV_X1 U7670 ( .A(n6717), .ZN(n6720) );
  AOI22_X1 U7671 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6729), .B1(n6718), 
        .B2(n6727), .ZN(n6719) );
  OAI211_X1 U7672 ( .C1(n6721), .C2(n6732), .A(n6720), .B(n6719), .ZN(U3114)
         );
  OAI22_X1 U7673 ( .A1(n6725), .A2(n6724), .B1(n6723), .B2(n6722), .ZN(n6726)
         );
  INV_X1 U7674 ( .A(n6726), .ZN(n6731) );
  AOI22_X1 U7675 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6729), .B1(n6728), 
        .B2(n6727), .ZN(n6730) );
  OAI211_X1 U7676 ( .C1(n6733), .C2(n6732), .A(n6731), .B(n6730), .ZN(U3115)
         );
  INV_X1 U7677 ( .A(n6734), .ZN(n6735) );
  OAI211_X1 U7678 ( .C1(STATE2_REG_0__SCAN_IN), .C2(STATE2_REG_2__SCAN_IN), 
        .A(n6735), .B(STATE2_REG_1__SCAN_IN), .ZN(n6743) );
  OAI21_X1 U7679 ( .B1(READY_N), .B2(n6737), .A(n6736), .ZN(n6740) );
  INV_X1 U7680 ( .A(n6738), .ZN(n6739) );
  AOI21_X1 U7681 ( .B1(n6741), .B2(n6740), .A(n6739), .ZN(n6742) );
  NAND2_X1 U7682 ( .A1(n6743), .A2(n6742), .ZN(U3149) );
  AND2_X1 U7683 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6786), .ZN(U3151) );
  INV_X1 U7684 ( .A(DATAWIDTH_REG_30__SCAN_IN), .ZN(n6877) );
  NOR2_X1 U7685 ( .A1(n6788), .A2(n6877), .ZN(U3152) );
  AND2_X1 U7686 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6786), .ZN(U3153) );
  AND2_X1 U7687 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6786), .ZN(U3154) );
  AND2_X1 U7688 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6786), .ZN(U3155) );
  AND2_X1 U7689 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6786), .ZN(U3156) );
  AND2_X1 U7690 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6786), .ZN(U3157) );
  AND2_X1 U7691 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6786), .ZN(U3158) );
  INV_X1 U7692 ( .A(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6915) );
  NOR2_X1 U7693 ( .A1(n6788), .A2(n6915), .ZN(U3159) );
  AND2_X1 U7694 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6786), .ZN(U3160) );
  INV_X1 U7695 ( .A(DATAWIDTH_REG_21__SCAN_IN), .ZN(n7065) );
  NOR2_X1 U7696 ( .A1(n6788), .A2(n7065), .ZN(U3161) );
  INV_X1 U7697 ( .A(DATAWIDTH_REG_20__SCAN_IN), .ZN(n7105) );
  NOR2_X1 U7698 ( .A1(n6788), .A2(n7105), .ZN(U3162) );
  INV_X1 U7699 ( .A(DATAWIDTH_REG_19__SCAN_IN), .ZN(n7059) );
  NOR2_X1 U7700 ( .A1(n6788), .A2(n7059), .ZN(U3163) );
  AND2_X1 U7701 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6786), .ZN(U3164) );
  INV_X1 U7702 ( .A(DATAWIDTH_REG_17__SCAN_IN), .ZN(n6852) );
  NOR2_X1 U7703 ( .A1(n6788), .A2(n6852), .ZN(U3165) );
  AND2_X1 U7704 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6786), .ZN(U3166) );
  AND2_X1 U7705 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6786), .ZN(U3167) );
  AND2_X1 U7706 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6786), .ZN(U3168) );
  AND2_X1 U7707 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6786), .ZN(U3169) );
  NOR2_X1 U7708 ( .A1(n6788), .A2(n7010), .ZN(U3170) );
  AND2_X1 U7709 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6786), .ZN(U3171) );
  AND2_X1 U7710 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6786), .ZN(U3172) );
  AND2_X1 U7711 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6786), .ZN(U3173) );
  AND2_X1 U7712 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6786), .ZN(U3174) );
  AND2_X1 U7713 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6786), .ZN(U3175) );
  INV_X1 U7714 ( .A(DATAWIDTH_REG_6__SCAN_IN), .ZN(n6999) );
  NOR2_X1 U7715 ( .A1(n6788), .A2(n6999), .ZN(U3176) );
  NOR2_X1 U7716 ( .A1(n6788), .A2(n7038), .ZN(U3177) );
  AND2_X1 U7717 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6786), .ZN(U3178) );
  AND2_X1 U7718 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6786), .ZN(U3179) );
  AND2_X1 U7719 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6786), .ZN(U3180) );
  INV_X1 U7720 ( .A(n6778), .ZN(n6781) );
  AOI22_X1 U7721 ( .A1(n6781), .A2(REIP_REG_2__SCAN_IN), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6780), .ZN(n6744) );
  OAI21_X1 U7722 ( .B1(n6792), .B2(n6783), .A(n6744), .ZN(U3184) );
  AOI22_X1 U7723 ( .A1(n6781), .A2(REIP_REG_3__SCAN_IN), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6780), .ZN(n6745) );
  OAI21_X1 U7724 ( .B1(n6746), .B2(n6783), .A(n6745), .ZN(U3185) );
  AOI22_X1 U7725 ( .A1(n6781), .A2(REIP_REG_5__SCAN_IN), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6774), .ZN(n6747) );
  OAI21_X1 U7726 ( .B1(n6748), .B2(n6783), .A(n6747), .ZN(U3187) );
  AOI22_X1 U7727 ( .A1(n6781), .A2(REIP_REG_6__SCAN_IN), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6774), .ZN(n6749) );
  OAI21_X1 U7728 ( .B1(n6750), .B2(n6783), .A(n6749), .ZN(U3188) );
  INV_X1 U7729 ( .A(n6783), .ZN(n6776) );
  INV_X1 U7730 ( .A(n6751), .ZN(n6780) );
  AOI22_X1 U7731 ( .A1(n6776), .A2(REIP_REG_6__SCAN_IN), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6780), .ZN(n6752) );
  OAI21_X1 U7732 ( .B1(n6753), .B2(n6778), .A(n6752), .ZN(U3189) );
  AOI22_X1 U7733 ( .A1(n6776), .A2(REIP_REG_8__SCAN_IN), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6780), .ZN(n6754) );
  OAI21_X1 U7734 ( .B1(n6756), .B2(n6778), .A(n6754), .ZN(U3191) );
  AOI22_X1 U7735 ( .A1(n6781), .A2(REIP_REG_10__SCAN_IN), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6780), .ZN(n6755) );
  OAI21_X1 U7736 ( .B1(n6756), .B2(n6783), .A(n6755), .ZN(U3192) );
  AOI22_X1 U7737 ( .A1(n6781), .A2(REIP_REG_11__SCAN_IN), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6780), .ZN(n6757) );
  OAI21_X1 U7738 ( .B1(n6965), .B2(n6783), .A(n6757), .ZN(U3193) );
  AOI22_X1 U7739 ( .A1(n6781), .A2(REIP_REG_12__SCAN_IN), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6780), .ZN(n6758) );
  OAI21_X1 U7740 ( .B1(n6997), .B2(n6783), .A(n6758), .ZN(U3194) );
  AOI22_X1 U7741 ( .A1(n6776), .A2(REIP_REG_12__SCAN_IN), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6780), .ZN(n6759) );
  OAI21_X1 U7742 ( .B1(n6761), .B2(n6778), .A(n6759), .ZN(U3195) );
  AOI22_X1 U7743 ( .A1(n6781), .A2(REIP_REG_14__SCAN_IN), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6780), .ZN(n6760) );
  OAI21_X1 U7744 ( .B1(n6761), .B2(n6783), .A(n6760), .ZN(U3196) );
  AOI22_X1 U7745 ( .A1(n6781), .A2(REIP_REG_15__SCAN_IN), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6780), .ZN(n6762) );
  OAI21_X1 U7746 ( .B1(n6763), .B2(n6783), .A(n6762), .ZN(U3197) );
  AOI22_X1 U7747 ( .A1(n6781), .A2(REIP_REG_16__SCAN_IN), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6780), .ZN(n6764) );
  OAI21_X1 U7748 ( .B1(n5787), .B2(n6783), .A(n6764), .ZN(U3198) );
  AOI22_X1 U7749 ( .A1(n6776), .A2(REIP_REG_16__SCAN_IN), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6780), .ZN(n6765) );
  OAI21_X1 U7750 ( .B1(n6766), .B2(n6778), .A(n6765), .ZN(U3199) );
  AOI22_X1 U7751 ( .A1(n6776), .A2(REIP_REG_17__SCAN_IN), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6780), .ZN(n6767) );
  OAI21_X1 U7752 ( .B1(n6862), .B2(n6778), .A(n6767), .ZN(U3200) );
  AOI22_X1 U7753 ( .A1(n6781), .A2(REIP_REG_19__SCAN_IN), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6774), .ZN(n6768) );
  OAI21_X1 U7754 ( .B1(n6862), .B2(n6783), .A(n6768), .ZN(U3201) );
  AOI22_X1 U7755 ( .A1(n6776), .A2(REIP_REG_19__SCAN_IN), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6774), .ZN(n6769) );
  OAI21_X1 U7756 ( .B1(n6770), .B2(n6778), .A(n6769), .ZN(U3202) );
  AOI22_X1 U7757 ( .A1(n6776), .A2(REIP_REG_23__SCAN_IN), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6774), .ZN(n6771) );
  OAI21_X1 U7758 ( .B1(n6773), .B2(n6778), .A(n6771), .ZN(U3206) );
  AOI22_X1 U7759 ( .A1(n6781), .A2(REIP_REG_25__SCAN_IN), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6774), .ZN(n6772) );
  OAI21_X1 U7760 ( .B1(n6773), .B2(n6783), .A(n6772), .ZN(U3207) );
  INV_X1 U7761 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6856) );
  AOI22_X1 U7762 ( .A1(n6776), .A2(REIP_REG_25__SCAN_IN), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6774), .ZN(n6775) );
  OAI21_X1 U7763 ( .B1(n6856), .B2(n6778), .A(n6775), .ZN(U3208) );
  AOI22_X1 U7764 ( .A1(n6776), .A2(REIP_REG_26__SCAN_IN), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6780), .ZN(n6777) );
  OAI21_X1 U7765 ( .B1(n6779), .B2(n6778), .A(n6777), .ZN(U3209) );
  AOI22_X1 U7766 ( .A1(n6781), .A2(REIP_REG_29__SCAN_IN), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6780), .ZN(n6782) );
  OAI21_X1 U7767 ( .B1(n6784), .B2(n6783), .A(n6782), .ZN(U3211) );
  INV_X1 U7768 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6931) );
  INV_X1 U7769 ( .A(n6787), .ZN(n6785) );
  AOI21_X1 U7770 ( .B1(n6931), .B2(n6786), .A(n6785), .ZN(U3451) );
  INV_X1 U7771 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6790) );
  OAI21_X1 U7772 ( .B1(n6788), .B2(n6790), .A(n6787), .ZN(U3452) );
  AOI221_X1 U7773 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n7076), .C1(n6931), 
        .C2(n6790), .A(n6789), .ZN(n6794) );
  OAI22_X1 U7774 ( .A1(n6796), .A2(BYTEENABLE_REG_2__SCAN_IN), .B1(n6792), 
        .B2(n6791), .ZN(n6793) );
  NOR2_X1 U7775 ( .A1(n6794), .A2(n6793), .ZN(U3468) );
  INV_X1 U7776 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n7022) );
  OAI21_X1 U7777 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6796), .ZN(n6795) );
  OAI21_X1 U7778 ( .B1(n6796), .B2(n7022), .A(n6795), .ZN(U3469) );
  OAI21_X1 U7779 ( .B1(n6799), .B2(n6798), .A(n6797), .ZN(n6801) );
  NAND3_X1 U7780 ( .A1(n6801), .A2(n6800), .A3(STATE2_REG_2__SCAN_IN), .ZN(
        n6802) );
  OAI21_X1 U7781 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n6803), .A(n6802), .ZN(
        n6811) );
  OAI211_X1 U7782 ( .C1(READY_N), .C2(n6806), .A(n6805), .B(n6804), .ZN(n6807)
         );
  NOR2_X1 U7783 ( .A1(n6808), .A2(n6807), .ZN(n6810) );
  NAND2_X1 U7784 ( .A1(n6810), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6809) );
  OAI21_X1 U7785 ( .B1(n6811), .B2(n6810), .A(n6809), .ZN(U3472) );
  AOI222_X1 U7786 ( .A1(EAX_REG_11__SCAN_IN), .A2(n6814), .B1(n6813), .B2(
        LWORD_REG_11__SCAN_IN), .C1(n6812), .C2(DATAO_REG_11__SCAN_IN), .ZN(
        n7127) );
  AOI22_X1 U7787 ( .A1(n6955), .A2(keyinput23), .B1(keyinput115), .B2(n6816), 
        .ZN(n6815) );
  OAI221_X1 U7788 ( .B1(n6955), .B2(keyinput23), .C1(n6816), .C2(keyinput115), 
        .A(n6815), .ZN(n6827) );
  AOI22_X1 U7789 ( .A1(n6818), .A2(keyinput54), .B1(n6953), .B2(keyinput106), 
        .ZN(n6817) );
  OAI221_X1 U7790 ( .B1(n6818), .B2(keyinput54), .C1(n6953), .C2(keyinput106), 
        .A(n6817), .ZN(n6826) );
  INV_X1 U7791 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n6821) );
  AOI22_X1 U7792 ( .A1(n6821), .A2(keyinput70), .B1(keyinput19), .B2(n6820), 
        .ZN(n6819) );
  OAI221_X1 U7793 ( .B1(n6821), .B2(keyinput70), .C1(n6820), .C2(keyinput19), 
        .A(n6819), .ZN(n6825) );
  XOR2_X1 U7794 ( .A(n6954), .B(keyinput67), .Z(n6823) );
  XNOR2_X1 U7795 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(keyinput94), .ZN(
        n6822) );
  NAND2_X1 U7796 ( .A1(n6823), .A2(n6822), .ZN(n6824) );
  NOR4_X1 U7797 ( .A1(n6827), .A2(n6826), .A3(n6825), .A4(n6824), .ZN(n7125)
         );
  NAND2_X1 U7798 ( .A1(n6829), .A2(keyinput83), .ZN(n6828) );
  OAI221_X1 U7799 ( .B1(n6830), .B2(keyinput31), .C1(n6829), .C2(keyinput83), 
        .A(n6828), .ZN(n6843) );
  AOI22_X1 U7800 ( .A1(n6833), .A2(keyinput18), .B1(n6832), .B2(keyinput44), 
        .ZN(n6831) );
  OAI221_X1 U7801 ( .B1(n6833), .B2(keyinput18), .C1(n6832), .C2(keyinput44), 
        .A(n6831), .ZN(n6842) );
  INV_X1 U7802 ( .A(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n6836) );
  AOI22_X1 U7803 ( .A1(n6836), .A2(keyinput84), .B1(keyinput10), .B2(n6835), 
        .ZN(n6834) );
  OAI221_X1 U7804 ( .B1(n6836), .B2(keyinput84), .C1(n6835), .C2(keyinput10), 
        .A(n6834), .ZN(n6841) );
  INV_X1 U7805 ( .A(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n6839) );
  AOI22_X1 U7806 ( .A1(n6839), .A2(keyinput11), .B1(keyinput63), .B2(n6838), 
        .ZN(n6837) );
  OAI221_X1 U7807 ( .B1(n6839), .B2(keyinput11), .C1(n6838), .C2(keyinput63), 
        .A(n6837), .ZN(n6840) );
  NOR4_X1 U7808 ( .A1(n6843), .A2(n6842), .A3(n6841), .A4(n6840), .ZN(n7124)
         );
  INV_X1 U7809 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n6846) );
  INV_X1 U7810 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n6845) );
  AOI22_X1 U7811 ( .A1(n6846), .A2(keyinput35), .B1(keyinput85), .B2(n6845), 
        .ZN(n6844) );
  OAI221_X1 U7812 ( .B1(n6846), .B2(keyinput35), .C1(n6845), .C2(keyinput85), 
        .A(n6844), .ZN(n6930) );
  AOI22_X1 U7813 ( .A1(n6849), .A2(keyinput66), .B1(n6848), .B2(keyinput105), 
        .ZN(n6847) );
  OAI221_X1 U7814 ( .B1(n6849), .B2(keyinput66), .C1(n6848), .C2(keyinput105), 
        .A(n6847), .ZN(n6929) );
  INV_X1 U7815 ( .A(LWORD_REG_11__SCAN_IN), .ZN(n6851) );
  OAI22_X1 U7816 ( .A1(n6852), .A2(keyinput72), .B1(n6851), .B2(keyinput122), 
        .ZN(n6850) );
  AOI221_X1 U7817 ( .B1(n6852), .B2(keyinput72), .C1(keyinput122), .C2(n6851), 
        .A(n6850), .ZN(n6869) );
  OAI22_X1 U7818 ( .A1(n4692), .A2(keyinput109), .B1(n6952), .B2(keyinput12), 
        .ZN(n6853) );
  AOI221_X1 U7819 ( .B1(n4692), .B2(keyinput109), .C1(keyinput12), .C2(n6952), 
        .A(n6853), .ZN(n6868) );
  INV_X1 U7820 ( .A(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n6951) );
  AOI22_X1 U7821 ( .A1(n6949), .A2(keyinput36), .B1(n6951), .B2(keyinput97), 
        .ZN(n6854) );
  OAI221_X1 U7822 ( .B1(n6949), .B2(keyinput36), .C1(n6951), .C2(keyinput97), 
        .A(n6854), .ZN(n6866) );
  INV_X1 U7823 ( .A(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n6950) );
  AOI22_X1 U7824 ( .A1(n6950), .A2(keyinput39), .B1(keyinput24), .B2(n6856), 
        .ZN(n6855) );
  OAI221_X1 U7825 ( .B1(n6950), .B2(keyinput39), .C1(n6856), .C2(keyinput24), 
        .A(n6855), .ZN(n6865) );
  INV_X1 U7826 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n6859) );
  INV_X1 U7827 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n6858) );
  AOI22_X1 U7828 ( .A1(n6859), .A2(keyinput1), .B1(keyinput56), .B2(n6858), 
        .ZN(n6857) );
  OAI221_X1 U7829 ( .B1(n6859), .B2(keyinput1), .C1(n6858), .C2(keyinput56), 
        .A(n6857), .ZN(n6864) );
  AOI22_X1 U7830 ( .A1(n6862), .A2(keyinput65), .B1(n6861), .B2(keyinput112), 
        .ZN(n6860) );
  OAI221_X1 U7831 ( .B1(n6862), .B2(keyinput65), .C1(n6861), .C2(keyinput112), 
        .A(n6860), .ZN(n6863) );
  NOR4_X1 U7832 ( .A1(n6866), .A2(n6865), .A3(n6864), .A4(n6863), .ZN(n6867)
         );
  NAND3_X1 U7833 ( .A1(n6869), .A2(n6868), .A3(n6867), .ZN(n6928) );
  INV_X1 U7834 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6872) );
  INV_X1 U7835 ( .A(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n6871) );
  AOI22_X1 U7836 ( .A1(n6872), .A2(keyinput27), .B1(n6871), .B2(keyinput95), 
        .ZN(n6870) );
  OAI221_X1 U7837 ( .B1(n6872), .B2(keyinput27), .C1(n6871), .C2(keyinput95), 
        .A(n6870), .ZN(n6883) );
  INV_X1 U7838 ( .A(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n6932) );
  AOI22_X1 U7839 ( .A1(n6874), .A2(keyinput117), .B1(n6932), .B2(keyinput88), 
        .ZN(n6873) );
  OAI221_X1 U7840 ( .B1(n6874), .B2(keyinput117), .C1(n6932), .C2(keyinput88), 
        .A(n6873), .ZN(n6882) );
  AOI22_X1 U7841 ( .A1(n6877), .A2(keyinput26), .B1(keyinput37), .B2(n6876), 
        .ZN(n6875) );
  OAI221_X1 U7842 ( .B1(n6877), .B2(keyinput26), .C1(n6876), .C2(keyinput37), 
        .A(n6875), .ZN(n6881) );
  AOI22_X1 U7843 ( .A1(n6879), .A2(keyinput34), .B1(keyinput28), .B2(n4059), 
        .ZN(n6878) );
  OAI221_X1 U7844 ( .B1(n6879), .B2(keyinput34), .C1(n4059), .C2(keyinput28), 
        .A(n6878), .ZN(n6880) );
  NOR4_X1 U7845 ( .A1(n6883), .A2(n6882), .A3(n6881), .A4(n6880), .ZN(n6926)
         );
  INV_X1 U7846 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n6885) );
  AOI22_X1 U7847 ( .A1(n6885), .A2(keyinput48), .B1(keyinput17), .B2(n6931), 
        .ZN(n6884) );
  OAI221_X1 U7848 ( .B1(n6885), .B2(keyinput48), .C1(n6931), .C2(keyinput17), 
        .A(n6884), .ZN(n6895) );
  AOI22_X1 U7849 ( .A1(n5158), .A2(keyinput33), .B1(n6936), .B2(keyinput87), 
        .ZN(n6886) );
  OAI221_X1 U7850 ( .B1(n5158), .B2(keyinput33), .C1(n6936), .C2(keyinput87), 
        .A(n6886), .ZN(n6894) );
  INV_X1 U7851 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n6889) );
  AOI22_X1 U7852 ( .A1(n6889), .A2(keyinput98), .B1(keyinput55), .B2(n6888), 
        .ZN(n6887) );
  OAI221_X1 U7853 ( .B1(n6889), .B2(keyinput98), .C1(n6888), .C2(keyinput55), 
        .A(n6887), .ZN(n6893) );
  INV_X1 U7854 ( .A(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n6937) );
  XOR2_X1 U7855 ( .A(n6937), .B(keyinput101), .Z(n6891) );
  XNOR2_X1 U7856 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .B(keyinput64), .ZN(n6890) );
  NAND2_X1 U7857 ( .A1(n6891), .A2(n6890), .ZN(n6892) );
  NOR4_X1 U7858 ( .A1(n6895), .A2(n6894), .A3(n6893), .A4(n6892), .ZN(n6925)
         );
  AOI22_X1 U7859 ( .A1(n6898), .A2(keyinput82), .B1(n6897), .B2(keyinput81), 
        .ZN(n6896) );
  OAI221_X1 U7860 ( .B1(n6898), .B2(keyinput82), .C1(n6897), .C2(keyinput81), 
        .A(n6896), .ZN(n6907) );
  INV_X1 U7861 ( .A(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n6934) );
  AOI22_X1 U7862 ( .A1(n6945), .A2(keyinput89), .B1(n6934), .B2(keyinput68), 
        .ZN(n6899) );
  OAI221_X1 U7863 ( .B1(n6945), .B2(keyinput89), .C1(n6934), .C2(keyinput68), 
        .A(n6899), .ZN(n6906) );
  INV_X1 U7864 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n6901) );
  AOI22_X1 U7865 ( .A1(n6966), .A2(keyinput45), .B1(n6901), .B2(keyinput40), 
        .ZN(n6900) );
  OAI221_X1 U7866 ( .B1(n6966), .B2(keyinput45), .C1(n6901), .C2(keyinput40), 
        .A(n6900), .ZN(n6905) );
  AOI22_X1 U7867 ( .A1(n6903), .A2(keyinput111), .B1(n6965), .B2(keyinput93), 
        .ZN(n6902) );
  OAI221_X1 U7868 ( .B1(n6903), .B2(keyinput111), .C1(n6965), .C2(keyinput93), 
        .A(n6902), .ZN(n6904) );
  NOR4_X1 U7869 ( .A1(n6907), .A2(n6906), .A3(n6905), .A4(n6904), .ZN(n6924)
         );
  AOI22_X1 U7870 ( .A1(n6910), .A2(keyinput86), .B1(keyinput25), .B2(n6909), 
        .ZN(n6908) );
  OAI221_X1 U7871 ( .B1(n6910), .B2(keyinput86), .C1(n6909), .C2(keyinput25), 
        .A(n6908), .ZN(n6922) );
  INV_X1 U7872 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n6938) );
  AOI22_X1 U7873 ( .A1(n6938), .A2(keyinput6), .B1(keyinput49), .B2(n6912), 
        .ZN(n6911) );
  OAI221_X1 U7874 ( .B1(n6938), .B2(keyinput6), .C1(n6912), .C2(keyinput49), 
        .A(n6911), .ZN(n6921) );
  INV_X1 U7875 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n6914) );
  AOI22_X1 U7876 ( .A1(n6915), .A2(keyinput114), .B1(n6914), .B2(keyinput57), 
        .ZN(n6913) );
  OAI221_X1 U7877 ( .B1(n6915), .B2(keyinput114), .C1(n6914), .C2(keyinput57), 
        .A(n6913), .ZN(n6920) );
  INV_X1 U7878 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n6918) );
  INV_X1 U7879 ( .A(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n6917) );
  AOI22_X1 U7880 ( .A1(n6918), .A2(keyinput43), .B1(n6917), .B2(keyinput0), 
        .ZN(n6916) );
  OAI221_X1 U7881 ( .B1(n6918), .B2(keyinput43), .C1(n6917), .C2(keyinput0), 
        .A(n6916), .ZN(n6919) );
  NOR4_X1 U7882 ( .A1(n6922), .A2(n6921), .A3(n6920), .A4(n6919), .ZN(n6923)
         );
  NAND4_X1 U7883 ( .A1(n6926), .A2(n6925), .A3(n6924), .A4(n6923), .ZN(n6927)
         );
  NOR4_X1 U7884 ( .A1(n6930), .A2(n6929), .A3(n6928), .A4(n6927), .ZN(n7123)
         );
  NAND4_X1 U7885 ( .A1(INSTQUEUE_REG_6__3__SCAN_IN), .A2(
        ADDRESS_REG_28__SCAN_IN), .A3(n6932), .A4(n6931), .ZN(n6933) );
  NOR3_X1 U7886 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(EAX_REG_29__SCAN_IN), 
        .A3(n6933), .ZN(n6947) );
  NOR4_X1 U7887 ( .A1(UWORD_REG_6__SCAN_IN), .A2(MORE_REG_SCAN_IN), .A3(
        LWORD_REG_12__SCAN_IN), .A4(n6934), .ZN(n6935) );
  NAND3_X1 U7888 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(n6935), .ZN(n6944) );
  NOR4_X1 U7889 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(n6937), .A3(n6936), 
        .A4(n5158), .ZN(n6942) );
  NOR4_X1 U7890 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(
        INSTQUEUE_REG_4__1__SCAN_IN), .A3(PHYADDRPOINTER_REG_28__SCAN_IN), 
        .A4(REIP_REG_18__SCAN_IN), .ZN(n6941) );
  NOR4_X1 U7891 ( .A1(INSTQUEUE_REG_14__2__SCAN_IN), .A2(EBX_REG_30__SCAN_IN), 
        .A3(EBX_REG_19__SCAN_IN), .A4(LWORD_REG_1__SCAN_IN), .ZN(n6940) );
  NOR4_X1 U7892 ( .A1(EAX_REG_12__SCAN_IN), .A2(EAX_REG_8__SCAN_IN), .A3(
        ADDRESS_REG_6__SCAN_IN), .A4(n6938), .ZN(n6939) );
  NAND4_X1 U7893 ( .A1(n6942), .A2(n6941), .A3(n6940), .A4(n6939), .ZN(n6943)
         );
  NOR4_X1 U7894 ( .A1(INSTQUEUE_REG_2__6__SCAN_IN), .A2(n6945), .A3(n6944), 
        .A4(n6943), .ZN(n6946) );
  NAND4_X1 U7895 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(UWORD_REG_8__SCAN_IN), 
        .A3(n6947), .A4(n6946), .ZN(n6989) );
  INV_X1 U7896 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n7110) );
  NAND4_X1 U7897 ( .A1(EBX_REG_25__SCAN_IN), .A2(EAX_REG_23__SCAN_IN), .A3(
        n6948), .A4(n7110), .ZN(n6963) );
  NAND4_X1 U7898 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6951), .A3(n6950), .A4(
        n6949), .ZN(n6962) );
  NAND4_X1 U7899 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(
        LWORD_REG_11__SCAN_IN), .A3(n4692), .A4(n6952), .ZN(n6961) );
  NOR4_X1 U7900 ( .A1(DATAI_1_), .A2(LWORD_REG_15__SCAN_IN), .A3(n6954), .A4(
        n6953), .ZN(n6959) );
  NOR4_X1 U7901 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(
        INSTQUEUE_REG_7__5__SCAN_IN), .A3(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .A4(ADDRESS_REG_21__SCAN_IN), .ZN(n6958) );
  NOR4_X1 U7902 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(DATAI_8_), .A3(
        ADDRESS_REG_20__SCAN_IN), .A4(ADDRESS_REG_19__SCAN_IN), .ZN(n6957) );
  NOR4_X1 U7903 ( .A1(INSTQUEUE_REG_15__2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(EBX_REG_20__SCAN_IN), .A4(n6955), 
        .ZN(n6956) );
  NAND4_X1 U7904 ( .A1(n6959), .A2(n6958), .A3(n6957), .A4(n6956), .ZN(n6960)
         );
  NOR4_X1 U7905 ( .A1(n6963), .A2(n6962), .A3(n6961), .A4(n6960), .ZN(n6987)
         );
  INV_X1 U7906 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n7006) );
  NOR4_X1 U7907 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTQUEUE_REG_10__1__SCAN_IN), .A3(DATAWIDTH_REG_12__SCAN_IN), .A4(
        n7006), .ZN(n6964) );
  NAND3_X1 U7908 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(DATAO_REG_18__SCAN_IN), 
        .A3(n6964), .ZN(n6975) );
  INV_X1 U7909 ( .A(DATAI_21_), .ZN(n7041) );
  NOR4_X1 U7910 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(
        DATAWIDTH_REG_5__SCAN_IN), .A3(n7040), .A4(n7041), .ZN(n6973) );
  NOR4_X1 U7911 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A3(BYTEENABLE_REG_0__SCAN_IN), .A4(
        n7025), .ZN(n6972) );
  NAND4_X1 U7912 ( .A1(BE_N_REG_0__SCAN_IN), .A2(REIP_REG_11__SCAN_IN), .A3(
        LWORD_REG_5__SCAN_IN), .A4(n6995), .ZN(n6970) );
  NAND4_X1 U7913 ( .A1(INSTQUEUE_REG_4__5__SCAN_IN), .A2(n6966), .A3(n6992), 
        .A4(n6965), .ZN(n6969) );
  NAND4_X1 U7914 ( .A1(INSTQUEUE_REG_0__5__SCAN_IN), .A2(
        INSTQUEUE_REG_11__3__SCAN_IN), .A3(INSTQUEUE_REG_0__3__SCAN_IN), .A4(
        INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n6968) );
  NAND4_X1 U7915 ( .A1(EBX_REG_9__SCAN_IN), .A2(INSTQUEUE_REG_9__2__SCAN_IN), 
        .A3(LWORD_REG_8__SCAN_IN), .A4(n7012), .ZN(n6967) );
  NOR4_X1 U7916 ( .A1(n6970), .A2(n6969), .A3(n6968), .A4(n6967), .ZN(n6971)
         );
  NAND3_X1 U7917 ( .A1(n6973), .A2(n6972), .A3(n6971), .ZN(n6974) );
  NOR4_X1 U7918 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(DATAO_REG_4__SCAN_IN), 
        .A3(n6975), .A4(n6974), .ZN(n6986) );
  NAND4_X1 U7919 ( .A1(n7095), .A2(n7092), .A3(n7088), .A4(n7091), .ZN(n6979)
         );
  INV_X1 U7920 ( .A(BE_N_REG_3__SCAN_IN), .ZN(n7089) );
  NAND4_X1 U7921 ( .A1(DATAO_REG_31__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        n7086), .A4(n7089), .ZN(n6978) );
  NAND4_X1 U7922 ( .A1(ADDRESS_REG_26__SCAN_IN), .A2(DATAO_REG_27__SCAN_IN), 
        .A3(n5571), .A4(n7108), .ZN(n6977) );
  INV_X1 U7923 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n7102) );
  NAND4_X1 U7924 ( .A1(INSTQUEUE_REG_6__6__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(n7102), .A4(n7101), .ZN(n6976) );
  NOR4_X1 U7925 ( .A1(n6979), .A2(n6978), .A3(n6977), .A4(n6976), .ZN(n6985)
         );
  INV_X1 U7926 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n7055) );
  NAND4_X1 U7927 ( .A1(DATAO_REG_26__SCAN_IN), .A2(n7055), .A3(n7061), .A4(
        n7058), .ZN(n6983) );
  NAND4_X1 U7928 ( .A1(INSTQUEUE_REG_0__2__SCAN_IN), .A2(DATAI_25_), .A3(
        CODEFETCH_REG_SCAN_IN), .A4(UWORD_REG_13__SCAN_IN), .ZN(n6982) );
  NAND4_X1 U7929 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(
        INSTQUEUE_REG_10__0__SCAN_IN), .A3(REIP_REG_0__SCAN_IN), .A4(n3935), 
        .ZN(n6981) );
  NAND4_X1 U7930 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(EBX_REG_17__SCAN_IN), 
        .A3(LWORD_REG_0__SCAN_IN), .A4(n7064), .ZN(n6980) );
  NOR4_X1 U7931 ( .A1(n6983), .A2(n6982), .A3(n6981), .A4(n6980), .ZN(n6984)
         );
  NAND4_X1 U7932 ( .A1(n6987), .A2(n6986), .A3(n6985), .A4(n6984), .ZN(n6988)
         );
  OAI21_X1 U7933 ( .B1(n6989), .B2(n6988), .A(ADDRESS_REG_2__SCAN_IN), .ZN(
        n7121) );
  AOI22_X1 U7934 ( .A1(n6992), .A2(keyinput62), .B1(keyinput125), .B2(n6991), 
        .ZN(n6990) );
  OAI221_X1 U7935 ( .B1(n6992), .B2(keyinput62), .C1(n6991), .C2(keyinput125), 
        .A(n6990), .ZN(n7004) );
  AOI22_X1 U7936 ( .A1(n6995), .A2(keyinput104), .B1(keyinput8), .B2(n6994), 
        .ZN(n6993) );
  OAI221_X1 U7937 ( .B1(n6995), .B2(keyinput104), .C1(n6994), .C2(keyinput8), 
        .A(n6993), .ZN(n7003) );
  AOI22_X1 U7938 ( .A1(n6997), .A2(keyinput108), .B1(n3953), .B2(keyinput74), 
        .ZN(n6996) );
  OAI221_X1 U7939 ( .B1(n6997), .B2(keyinput108), .C1(n3953), .C2(keyinput74), 
        .A(n6996), .ZN(n7002) );
  INV_X1 U7940 ( .A(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n7000) );
  AOI22_X1 U7941 ( .A1(n7000), .A2(keyinput5), .B1(keyinput16), .B2(n6999), 
        .ZN(n6998) );
  OAI221_X1 U7942 ( .B1(n7000), .B2(keyinput5), .C1(n6999), .C2(keyinput16), 
        .A(n6998), .ZN(n7001) );
  NOR4_X1 U7943 ( .A1(n7004), .A2(n7003), .A3(n7002), .A4(n7001), .ZN(n7053)
         );
  AOI22_X1 U7944 ( .A1(n7007), .A2(keyinput99), .B1(n7006), .B2(keyinput110), 
        .ZN(n7005) );
  OAI221_X1 U7945 ( .B1(n7007), .B2(keyinput99), .C1(n7006), .C2(keyinput110), 
        .A(n7005), .ZN(n7020) );
  INV_X1 U7946 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n7009) );
  AOI22_X1 U7947 ( .A1(n7010), .A2(keyinput50), .B1(n7009), .B2(keyinput14), 
        .ZN(n7008) );
  OAI221_X1 U7948 ( .B1(n7010), .B2(keyinput50), .C1(n7009), .C2(keyinput14), 
        .A(n7008), .ZN(n7019) );
  AOI22_X1 U7949 ( .A1(n7013), .A2(keyinput38), .B1(keyinput120), .B2(n7012), 
        .ZN(n7011) );
  OAI221_X1 U7950 ( .B1(n7013), .B2(keyinput38), .C1(n7012), .C2(keyinput120), 
        .A(n7011), .ZN(n7018) );
  INV_X1 U7951 ( .A(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n7015) );
  AOI22_X1 U7952 ( .A1(n7016), .A2(keyinput59), .B1(n7015), .B2(keyinput7), 
        .ZN(n7014) );
  OAI221_X1 U7953 ( .B1(n7016), .B2(keyinput59), .C1(n7015), .C2(keyinput7), 
        .A(n7014), .ZN(n7017) );
  NOR4_X1 U7954 ( .A1(n7020), .A2(n7019), .A3(n7018), .A4(n7017), .ZN(n7052)
         );
  AOI22_X1 U7955 ( .A1(n7023), .A2(keyinput32), .B1(keyinput127), .B2(n7022), 
        .ZN(n7021) );
  OAI221_X1 U7956 ( .B1(n7023), .B2(keyinput32), .C1(n7022), .C2(keyinput127), 
        .A(n7021), .ZN(n7035) );
  AOI22_X1 U7957 ( .A1(n4700), .A2(keyinput4), .B1(keyinput102), .B2(n7025), 
        .ZN(n7024) );
  OAI221_X1 U7958 ( .B1(n4700), .B2(keyinput4), .C1(n7025), .C2(keyinput102), 
        .A(n7024), .ZN(n7034) );
  AOI22_X1 U7959 ( .A1(n7028), .A2(keyinput103), .B1(n7027), .B2(keyinput77), 
        .ZN(n7026) );
  OAI221_X1 U7960 ( .B1(n7028), .B2(keyinput103), .C1(n7027), .C2(keyinput77), 
        .A(n7026), .ZN(n7033) );
  INV_X1 U7961 ( .A(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n7029) );
  XOR2_X1 U7962 ( .A(n7029), .B(keyinput41), .Z(n7031) );
  XNOR2_X1 U7963 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .B(keyinput73), .ZN(n7030)
         );
  NAND2_X1 U7964 ( .A1(n7031), .A2(n7030), .ZN(n7032) );
  NOR4_X1 U7965 ( .A1(n7035), .A2(n7034), .A3(n7033), .A4(n7032), .ZN(n7051)
         );
  INV_X1 U7966 ( .A(DATAI_25_), .ZN(n7037) );
  AOI22_X1 U7967 ( .A1(n7038), .A2(keyinput15), .B1(n7037), .B2(keyinput47), 
        .ZN(n7036) );
  OAI221_X1 U7968 ( .B1(n7038), .B2(keyinput15), .C1(n7037), .C2(keyinput47), 
        .A(n7036), .ZN(n7049) );
  AOI22_X1 U7969 ( .A1(n5870), .A2(keyinput119), .B1(keyinput60), .B2(n7040), 
        .ZN(n7039) );
  OAI221_X1 U7970 ( .B1(n5870), .B2(keyinput119), .C1(n7040), .C2(keyinput60), 
        .A(n7039), .ZN(n7048) );
  XOR2_X1 U7971 ( .A(n7041), .B(keyinput9), .Z(n7046) );
  INV_X1 U7972 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n7042) );
  XOR2_X1 U7973 ( .A(n7042), .B(keyinput80), .Z(n7045) );
  XNOR2_X1 U7974 ( .A(INSTQUEUE_REG_9__1__SCAN_IN), .B(keyinput71), .ZN(n7044)
         );
  XNOR2_X1 U7975 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .B(keyinput116), .ZN(n7043) );
  NAND4_X1 U7976 ( .A1(n7046), .A2(n7045), .A3(n7044), .A4(n7043), .ZN(n7047)
         );
  NOR3_X1 U7977 ( .A1(n7049), .A2(n7048), .A3(n7047), .ZN(n7050) );
  NAND4_X1 U7978 ( .A1(n7053), .A2(n7052), .A3(n7051), .A4(n7050), .ZN(n7120)
         );
  AOI22_X1 U7979 ( .A1(n7056), .A2(keyinput75), .B1(n7055), .B2(keyinput46), 
        .ZN(n7054) );
  OAI221_X1 U7980 ( .B1(n7056), .B2(keyinput75), .C1(n7055), .C2(keyinput46), 
        .A(n7054), .ZN(n7069) );
  AOI22_X1 U7981 ( .A1(n7059), .A2(keyinput100), .B1(n7058), .B2(keyinput79), 
        .ZN(n7057) );
  OAI221_X1 U7982 ( .B1(n7059), .B2(keyinput100), .C1(n7058), .C2(keyinput79), 
        .A(n7057), .ZN(n7068) );
  AOI22_X1 U7983 ( .A1(n7062), .A2(keyinput22), .B1(n7061), .B2(keyinput42), 
        .ZN(n7060) );
  OAI221_X1 U7984 ( .B1(n7062), .B2(keyinput22), .C1(n7061), .C2(keyinput42), 
        .A(n7060), .ZN(n7067) );
  AOI22_X1 U7985 ( .A1(n7065), .A2(keyinput20), .B1(n7064), .B2(keyinput78), 
        .ZN(n7063) );
  OAI221_X1 U7986 ( .B1(n7065), .B2(keyinput20), .C1(n7064), .C2(keyinput78), 
        .A(n7063), .ZN(n7066) );
  NOR4_X1 U7987 ( .A1(n7069), .A2(n7068), .A3(n7067), .A4(n7066), .ZN(n7118)
         );
  INV_X1 U7988 ( .A(LWORD_REG_0__SCAN_IN), .ZN(n7071) );
  AOI22_X1 U7989 ( .A1(n7071), .A2(keyinput29), .B1(n5575), .B2(keyinput51), 
        .ZN(n7070) );
  OAI221_X1 U7990 ( .B1(n7071), .B2(keyinput29), .C1(n5575), .C2(keyinput51), 
        .A(n7070), .ZN(n7083) );
  INV_X1 U7991 ( .A(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n7074) );
  INV_X1 U7992 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n7073) );
  AOI22_X1 U7993 ( .A1(n7074), .A2(keyinput96), .B1(keyinput3), .B2(n7073), 
        .ZN(n7072) );
  OAI221_X1 U7994 ( .B1(n7074), .B2(keyinput96), .C1(n7073), .C2(keyinput3), 
        .A(n7072), .ZN(n7082) );
  AOI22_X1 U7995 ( .A1(n7076), .A2(keyinput90), .B1(n3935), .B2(keyinput91), 
        .ZN(n7075) );
  OAI221_X1 U7996 ( .B1(n7076), .B2(keyinput90), .C1(n3935), .C2(keyinput91), 
        .A(n7075), .ZN(n7081) );
  INV_X1 U7997 ( .A(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n7079) );
  AOI22_X1 U7998 ( .A1(n7079), .A2(keyinput124), .B1(keyinput126), .B2(n7078), 
        .ZN(n7077) );
  OAI221_X1 U7999 ( .B1(n7079), .B2(keyinput124), .C1(n7078), .C2(keyinput126), 
        .A(n7077), .ZN(n7080) );
  NOR4_X1 U8000 ( .A1(n7083), .A2(n7082), .A3(n7081), .A4(n7080), .ZN(n7117)
         );
  AOI22_X1 U8001 ( .A1(n7086), .A2(keyinput2), .B1(n7085), .B2(keyinput61), 
        .ZN(n7084) );
  OAI221_X1 U8002 ( .B1(n7086), .B2(keyinput2), .C1(n7085), .C2(keyinput61), 
        .A(n7084), .ZN(n7099) );
  AOI22_X1 U8003 ( .A1(n7089), .A2(keyinput58), .B1(keyinput69), .B2(n7088), 
        .ZN(n7087) );
  OAI221_X1 U8004 ( .B1(n7089), .B2(keyinput58), .C1(n7088), .C2(keyinput69), 
        .A(n7087), .ZN(n7098) );
  AOI22_X1 U8005 ( .A1(n7092), .A2(keyinput113), .B1(keyinput52), .B2(n7091), 
        .ZN(n7090) );
  OAI221_X1 U8006 ( .B1(n7092), .B2(keyinput113), .C1(n7091), .C2(keyinput52), 
        .A(n7090), .ZN(n7097) );
  INV_X1 U8007 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n7094) );
  AOI22_X1 U8008 ( .A1(n7095), .A2(keyinput123), .B1(keyinput13), .B2(n7094), 
        .ZN(n7093) );
  OAI221_X1 U8009 ( .B1(n7095), .B2(keyinput123), .C1(n7094), .C2(keyinput13), 
        .A(n7093), .ZN(n7096) );
  NOR4_X1 U8010 ( .A1(n7099), .A2(n7098), .A3(n7097), .A4(n7096), .ZN(n7116)
         );
  AOI22_X1 U8011 ( .A1(n7102), .A2(keyinput107), .B1(keyinput30), .B2(n7101), 
        .ZN(n7100) );
  OAI221_X1 U8012 ( .B1(n7102), .B2(keyinput107), .C1(n7101), .C2(keyinput30), 
        .A(n7100), .ZN(n7114) );
  AOI22_X1 U8013 ( .A1(n7105), .A2(keyinput76), .B1(keyinput53), .B2(n7104), 
        .ZN(n7103) );
  OAI221_X1 U8014 ( .B1(n7105), .B2(keyinput76), .C1(n7104), .C2(keyinput53), 
        .A(n7103), .ZN(n7113) );
  AOI22_X1 U8015 ( .A1(n7108), .A2(keyinput21), .B1(keyinput118), .B2(n7107), 
        .ZN(n7106) );
  OAI221_X1 U8016 ( .B1(n7108), .B2(keyinput21), .C1(n7107), .C2(keyinput118), 
        .A(n7106), .ZN(n7112) );
  AOI22_X1 U8017 ( .A1(n5571), .A2(keyinput92), .B1(n7110), .B2(keyinput121), 
        .ZN(n7109) );
  OAI221_X1 U8018 ( .B1(n5571), .B2(keyinput92), .C1(n7110), .C2(keyinput121), 
        .A(n7109), .ZN(n7111) );
  NOR4_X1 U8019 ( .A1(n7114), .A2(n7113), .A3(n7112), .A4(n7111), .ZN(n7115)
         );
  NAND4_X1 U8020 ( .A1(n7118), .A2(n7117), .A3(n7116), .A4(n7115), .ZN(n7119)
         );
  AOI211_X1 U8021 ( .C1(keyinput31), .C2(n7121), .A(n7120), .B(n7119), .ZN(
        n7122) );
  NAND4_X1 U8022 ( .A1(n7125), .A2(n7124), .A3(n7123), .A4(n7122), .ZN(n7126)
         );
  XOR2_X1 U8023 ( .A(n7127), .B(n7126), .Z(U2912) );
  CLKBUF_X1 U3538 ( .A(n3467), .Z(n3468) );
  CLKBUF_X3 U3550 ( .A(n5007), .Z(n3089) );
  NAND2_X1 U3554 ( .A1(n3591), .A2(n3590), .ZN(n3592) );
  CLKBUF_X1 U3558 ( .A(n4387), .Z(n6203) );
  CLKBUF_X1 U3995 ( .A(n5377), .Z(n3085) );
  XNOR2_X1 U4419 ( .A(n3592), .B(n6648), .ZN(n4661) );
endmodule

