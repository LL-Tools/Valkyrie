

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10288, n10289, n10290,
         n10291, n10292, n10293, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576;

  NAND2_X1 U4886 ( .A1(n7194), .A2(n7213), .ZN(n6527) );
  NAND2_X1 U4887 ( .A1(n5515), .A2(n5514), .ZN(n8535) );
  INV_X1 U4888 ( .A(n6591), .ZN(n7759) );
  CLKBUF_X1 U4889 ( .A(n6199), .Z(n4389) );
  INV_X1 U4890 ( .A(n7847), .ZN(n8189) );
  INV_X1 U4891 ( .A(n8861), .ZN(n8004) );
  INV_X1 U4892 ( .A(n8193), .ZN(n4944) );
  AND2_X2 U4893 ( .A1(n9626), .A2(n6164), .ZN(n7169) );
  MUX2_X1 U4894 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5058), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n7061) );
  AND2_X1 U4895 ( .A1(n5186), .A2(n5185), .ZN(n9990) );
  AOI21_X1 U4896 ( .B1(n9410), .B2(n7363), .A(n6350), .ZN(n9379) );
  BUF_X1 U4897 ( .A(n6446), .Z(n4387) );
  OR2_X1 U4898 ( .A1(n9235), .A2(n9498), .ZN(n4409) );
  INV_X1 U4899 ( .A(n5524), .ZN(n5800) );
  INV_X1 U4900 ( .A(n8865), .ZN(n8874) );
  NAND2_X1 U4901 ( .A1(n8080), .A2(n8286), .ZN(n8317) );
  INV_X1 U4902 ( .A(n8250), .ZN(n7051) );
  INV_X1 U4903 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5148) );
  XNOR2_X1 U4904 ( .A(n5237), .B(n5228), .ZN(n5460) );
  INV_X2 U4905 ( .A(n7759), .ZN(n6670) );
  BUF_X1 U4906 ( .A(n6228), .Z(n6558) );
  INV_X1 U4907 ( .A(n9228), .ZN(n4994) );
  OR2_X1 U4908 ( .A1(n4383), .A2(n4944), .ZN(n6584) );
  AOI21_X1 U4909 ( .B1(n9806), .B2(n8874), .A(n7789), .ZN(n8930) );
  INV_X2 U4910 ( .A(n8836), .ZN(n8872) );
  NAND2_X1 U4911 ( .A1(n10156), .A2(n8789), .ZN(n5905) );
  NAND2_X1 U4912 ( .A1(n10193), .A2(n10072), .ZN(n10065) );
  BUF_X1 U4913 ( .A(n5407), .Z(n5620) );
  INV_X1 U4914 ( .A(n7959), .ZN(n10380) );
  AND2_X1 U4915 ( .A1(n6421), .A2(n6420), .ZN(n9264) );
  NAND2_X1 U4916 ( .A1(n6456), .A2(n6455), .ZN(n9498) );
  CLKBUF_X3 U4917 ( .A(n5225), .Z(n7388) );
  CLKBUF_X3 U4918 ( .A(n6574), .Z(n4384) );
  NAND2_X2 U4920 ( .A1(n4830), .A2(n4829), .ZN(n9882) );
  NAND2_X2 U4921 ( .A1(n9918), .A2(n7040), .ZN(n4830) );
  INV_X1 U4922 ( .A(n5225), .ZN(n4382) );
  NAND2_X2 U4923 ( .A1(n5031), .A2(n7061), .ZN(n7812) );
  NOR2_X4 U4924 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5062) );
  NAND2_X2 U4925 ( .A1(n6119), .A2(n6157), .ZN(n6563) );
  INV_X2 U4926 ( .A(n9122), .ZN(n7218) );
  NOR2_X2 U4927 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5053) );
  AND2_X4 U4928 ( .A1(n4939), .A2(n4938), .ZN(n5225) );
  INV_X2 U4929 ( .A(n5225), .ZN(n5398) );
  BUF_X8 U4930 ( .A(n7389), .Z(n4522) );
  NOR2_X2 U4931 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5052) );
  NAND4_X2 U4932 ( .A1(n6192), .A2(n6191), .A3(n6190), .A4(n6189), .ZN(n6592)
         );
  NAND2_X2 U4933 ( .A1(n4439), .A2(n5038), .ZN(n5076) );
  OR2_X2 U4934 ( .A1(n5362), .A2(n5143), .ZN(n4777) );
  NAND2_X2 U4935 ( .A1(n4943), .A2(n6585), .ZN(n6594) );
  NOR2_X2 U4936 ( .A1(n7637), .A2(n4482), .ZN(n7859) );
  AND3_X2 U4937 ( .A1(n5063), .A2(n5055), .A3(n6914), .ZN(n5038) );
  BUF_X1 U4939 ( .A(n6574), .Z(n4383) );
  XNOR2_X2 U4940 ( .A(n5571), .B(n5034), .ZN(n7419) );
  NAND2_X2 U4941 ( .A1(n8003), .A2(n8002), .ZN(n8237) );
  NAND2_X2 U4942 ( .A1(n6266), .A2(n6265), .ZN(n9587) );
  AND2_X1 U4943 ( .A1(n9626), .A2(n6164), .ZN(n4385) );
  AND2_X1 U4944 ( .A1(n9626), .A2(n6164), .ZN(n4386) );
  OR2_X1 U4945 ( .A1(n5225), .A2(n5226), .ZN(n5227) );
  AND2_X2 U4946 ( .A1(n7792), .A2(n7793), .ZN(n7798) );
  AND2_X4 U4947 ( .A1(n5378), .A2(n5377), .ZN(n4402) );
  INV_X1 U4948 ( .A(n5465), .ZN(n5766) );
  AOI21_X2 U4949 ( .B1(n7164), .B2(n7163), .A(n7162), .ZN(n8907) );
  XNOR2_X2 U4950 ( .A(n5756), .B(n5755), .ZN(n8573) );
  NAND2_X2 U4951 ( .A1(n5159), .A2(n7686), .ZN(n5407) );
  NAND2_X2 U4952 ( .A1(n6114), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6117) );
  CLKBUF_X3 U4953 ( .A(n6446), .Z(n4388) );
  BUF_X1 U4954 ( .A(n6233), .Z(n6446) );
  AOI211_X1 U4955 ( .C1(n5812), .C2(n5811), .A(n5810), .B(n5809), .ZN(n5831)
         );
  NOR2_X2 U4956 ( .A1(n7546), .A2(n6047), .ZN(n7593) );
  NAND2_X1 U4957 ( .A1(n9249), .A2(n7297), .ZN(n9229) );
  NAND2_X1 U4958 ( .A1(n9330), .A2(n9338), .ZN(n9331) );
  NAND2_X1 U4959 ( .A1(n4945), .A2(n4946), .ZN(n9010) );
  NAND2_X1 U4960 ( .A1(n5527), .A2(n5526), .ZN(n10181) );
  NAND2_X1 U4961 ( .A1(n8317), .A2(n5976), .ZN(n8076) );
  NAND2_X1 U4962 ( .A1(n6316), .A2(n6315), .ZN(n6570) );
  NAND2_X1 U4963 ( .A1(n5491), .A2(n5490), .ZN(n5976) );
  NAND2_X1 U4964 ( .A1(n5917), .A2(n7933), .ZN(n7936) );
  NAND2_X1 U4965 ( .A1(n9802), .A2(n10401), .ZN(n7102) );
  INV_X1 U4966 ( .A(n9796), .ZN(n8510) );
  NAND2_X1 U4967 ( .A1(n5971), .A2(n5864), .ZN(n7938) );
  INV_X1 U4968 ( .A(n8246), .ZN(n10401) );
  AND4_X1 U4969 ( .A1(n5581), .A2(n5580), .A3(n5579), .A4(n5578), .ZN(n8533)
         );
  INV_X1 U4970 ( .A(n7089), .ZN(n5854) );
  NAND2_X1 U4971 ( .A1(n8250), .A2(n7941), .ZN(n7620) );
  CLKBUF_X3 U4972 ( .A(n7091), .Z(n9806) );
  CLKBUF_X2 U4973 ( .A(n7090), .Z(n8925) );
  INV_X1 U4974 ( .A(n9801), .ZN(n8011) );
  AND4_X1 U4975 ( .A1(n5438), .A2(n5437), .A3(n5436), .A4(n5435), .ZN(n7097)
         );
  AND4_X1 U4976 ( .A1(n5418), .A2(n5417), .A3(n5416), .A4(n5415), .ZN(n7090)
         );
  INV_X1 U4977 ( .A(n9123), .ZN(n7923) );
  INV_X1 U4978 ( .A(n7982), .ZN(n7972) );
  INV_X1 U4979 ( .A(n6199), .ZN(n7924) );
  INV_X1 U4980 ( .A(n6592), .ZN(n7774) );
  INV_X4 U4981 ( .A(n5464), .ZN(n5762) );
  INV_X1 U4982 ( .A(n7339), .ZN(n7340) );
  NAND2_X1 U4983 ( .A1(n6554), .A2(n7981), .ZN(n6585) );
  INV_X1 U4984 ( .A(n7998), .ZN(n6554) );
  NAND2_X2 U4985 ( .A1(n6563), .A2(n8695), .ZN(n6197) );
  OR2_X1 U4986 ( .A1(n10121), .A2(n4831), .ZN(n10207) );
  NOR2_X1 U4987 ( .A1(n4435), .A2(n4524), .ZN(n4523) );
  AND2_X1 U4988 ( .A1(n8895), .A2(n7048), .ZN(n8947) );
  NAND2_X1 U4989 ( .A1(n10103), .A2(n8937), .ZN(n10111) );
  NAND2_X1 U4990 ( .A1(n4536), .A2(n7149), .ZN(n8895) );
  OR2_X1 U4991 ( .A1(n8936), .A2(n8935), .ZN(n8937) );
  NAND2_X1 U4992 ( .A1(n4680), .A2(n4677), .ZN(n5892) );
  AOI21_X1 U4993 ( .B1(n8914), .B2(n9385), .A(n8913), .ZN(n9485) );
  AOI21_X1 U4994 ( .B1(n4988), .B2(n4987), .A(n4985), .ZN(n7183) );
  OAI21_X1 U4995 ( .B1(n5853), .B2(n4679), .A(n5948), .ZN(n4678) );
  AND2_X1 U4996 ( .A1(n8905), .A2(n4440), .ZN(n9491) );
  AND2_X1 U4997 ( .A1(n4997), .A2(n7308), .ZN(n9218) );
  AND2_X1 U4998 ( .A1(n5777), .A2(n5776), .ZN(n5808) );
  NAND2_X1 U4999 ( .A1(n9229), .A2(n9228), .ZN(n4997) );
  AND2_X1 U5000 ( .A1(n6747), .A2(n6746), .ZN(n8900) );
  AND2_X1 U5001 ( .A1(n9859), .A2(n9639), .ZN(n8938) );
  NAND2_X1 U5002 ( .A1(n5817), .A2(n5816), .ZN(n10107) );
  AND2_X1 U5003 ( .A1(n9277), .A2(n9340), .ZN(n9326) );
  NAND2_X1 U5004 ( .A1(n8582), .A2(n8583), .ZN(n4873) );
  NAND2_X1 U5005 ( .A1(n5814), .A2(n5813), .ZN(n5387) );
  OAI21_X1 U5006 ( .B1(n9010), .B2(n6674), .A(n6673), .ZN(n9015) );
  NAND2_X1 U5007 ( .A1(n6482), .A2(n6481), .ZN(n9220) );
  NAND2_X1 U5008 ( .A1(n5758), .A2(n5757), .ZN(n10123) );
  NOR2_X1 U5009 ( .A1(n7031), .A2(n4839), .ZN(n4838) );
  OR2_X1 U5010 ( .A1(n9943), .A2(n7035), .ZN(n7031) );
  CLKBUF_X1 U5011 ( .A(n7348), .Z(n4518) );
  NAND2_X1 U5012 ( .A1(n5723), .A2(n5722), .ZN(n10134) );
  NAND2_X1 U5013 ( .A1(n6424), .A2(n6423), .ZN(n9520) );
  AND2_X1 U5014 ( .A1(n8581), .A2(n8580), .ZN(n8582) );
  NAND2_X1 U5015 ( .A1(n6402), .A2(n6401), .ZN(n9523) );
  OR2_X1 U5016 ( .A1(n8464), .A2(n8463), .ZN(n8580) );
  AND2_X1 U5017 ( .A1(n9429), .A2(n8676), .ZN(n8671) );
  AND2_X1 U5018 ( .A1(n8446), .A2(n8447), .ZN(n8463) );
  INV_X1 U5019 ( .A(n9264), .ZN(n4390) );
  OR2_X1 U5020 ( .A1(n9146), .A2(n6074), .ZN(n6075) );
  NAND2_X1 U5021 ( .A1(n5612), .A2(n5611), .ZN(n7028) );
  XNOR2_X1 U5022 ( .A(n6074), .B(n6073), .ZN(n9141) );
  NAND2_X1 U5023 ( .A1(n6396), .A2(n6395), .ZN(n9528) );
  NAND2_X1 U5024 ( .A1(n6373), .A2(n6372), .ZN(n9539) );
  NAND2_X1 U5025 ( .A1(n5691), .A2(n5690), .ZN(n5304) );
  NAND2_X2 U5026 ( .A1(n5605), .A2(n5604), .ZN(n10165) );
  NAND2_X1 U5027 ( .A1(n7122), .A2(n7120), .ZN(n10170) );
  XNOR2_X1 U5028 ( .A(n5650), .B(n5615), .ZN(n7704) );
  NAND2_X1 U5029 ( .A1(n8480), .A2(n6061), .ZN(n8708) );
  AND2_X1 U5030 ( .A1(n7015), .A2(n5921), .ZN(n8319) );
  NAND2_X1 U5031 ( .A1(n6305), .A2(n6304), .ZN(n9565) );
  OR2_X1 U5032 ( .A1(n10427), .A2(n8386), .ZN(n7015) );
  AND2_X1 U5033 ( .A1(n7235), .A2(n7228), .ZN(n8544) );
  NAND2_X2 U5034 ( .A1(n5548), .A2(n5547), .ZN(n10193) );
  AND2_X1 U5035 ( .A1(n7623), .A2(n7622), .ZN(n7627) );
  NAND2_X1 U5036 ( .A1(n4544), .A2(n6281), .ZN(n9580) );
  NAND2_X1 U5037 ( .A1(n9119), .A2(n8554), .ZN(n7235) );
  XNOR2_X1 U5038 ( .A(n4521), .B(n5503), .ZN(n7421) );
  AOI22_X1 U5039 ( .A1(n8004), .A2(n7982), .B1(n7624), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n7622) );
  AND2_X1 U5040 ( .A1(n8262), .A2(n7102), .ZN(n8061) );
  INV_X1 U5041 ( .A(n8260), .ZN(n8346) );
  NAND2_X1 U5042 ( .A1(n6329), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6356) );
  CLKBUF_X2 U5043 ( .A(n8861), .Z(n4401) );
  NAND2_X1 U5044 ( .A1(n5463), .A2(n5462), .ZN(n8260) );
  INV_X1 U5045 ( .A(n9806), .ZN(n8087) );
  AND4_X1 U5046 ( .A1(n5554), .A2(n5553), .A3(n5552), .A4(n5551), .ZN(n10072)
         );
  BUF_X4 U5047 ( .A(n8439), .Z(n8785) );
  NAND4_X2 U5048 ( .A1(n5451), .A2(n5450), .A3(n5449), .A4(n5448), .ZN(n9802)
         );
  NAND2_X1 U5049 ( .A1(n6526), .A2(n7211), .ZN(n6525) );
  INV_X1 U5050 ( .A(n7873), .ZN(n8092) );
  NAND4_X1 U5051 ( .A1(n5393), .A2(n5394), .A3(n5392), .A4(n5391), .ZN(n7091)
         );
  NAND2_X1 U5052 ( .A1(n10457), .A2(n7196), .ZN(n7352) );
  CLKBUF_X1 U5053 ( .A(n7720), .Z(n4495) );
  INV_X1 U5054 ( .A(n7922), .ZN(n9460) );
  INV_X1 U5055 ( .A(n5469), .ZN(n5367) );
  CLKBUF_X1 U5056 ( .A(n6600), .Z(n9445) );
  NAND2_X1 U5057 ( .A1(n4726), .A2(n4449), .ZN(n9440) );
  NAND2_X1 U5058 ( .A1(n9468), .A2(n7740), .ZN(n7196) );
  NAND4_X1 U5059 ( .A1(n6209), .A2(n6208), .A3(n6207), .A4(n6206), .ZN(n9123)
         );
  AOI21_X1 U5060 ( .B1(P2_REG2_REG_4__SCAN_IN), .B2(n6210), .A(n7598), .ZN(
        n7548) );
  NAND4_X1 U5061 ( .A1(n6223), .A2(n6222), .A3(n6221), .A4(n6220), .ZN(n9443)
         );
  NAND4_X1 U5062 ( .A1(n6174), .A2(n6173), .A3(n6172), .A4(n6171), .ZN(n6199)
         );
  INV_X1 U5063 ( .A(n5378), .ZN(n10235) );
  CLKBUF_X1 U5064 ( .A(n4388), .Z(n7177) );
  OR2_X1 U5065 ( .A1(n7187), .A2(n7378), .ZN(n6591) );
  AOI21_X1 U5066 ( .B1(n4920), .B2(n4925), .A(n4459), .ZN(n4919) );
  AND2_X1 U5067 ( .A1(n7993), .A2(n8059), .ZN(n7941) );
  NAND2_X2 U5068 ( .A1(n4384), .A2(n7189), .ZN(n7339) );
  AND2_X1 U5069 ( .A1(n4922), .A2(n5555), .ZN(n4920) );
  AND2_X2 U5070 ( .A1(n5363), .A2(n10227), .ZN(n5378) );
  INV_X1 U5071 ( .A(n7169), .ZN(n6228) );
  XNOR2_X1 U5072 ( .A(n4863), .B(P1_IR_REG_26__SCAN_IN), .ZN(n7082) );
  MUX2_X1 U5073 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5361), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5363) );
  NAND2_X1 U5074 ( .A1(n5088), .A2(n5360), .ZN(n7686) );
  XNOR2_X1 U5075 ( .A(n6513), .B(n6512), .ZN(n7981) );
  NAND2_X1 U5076 ( .A1(n7065), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4863) );
  MUX2_X1 U5077 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6113), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n6115) );
  MUX2_X1 U5078 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5087), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n5088) );
  NAND2_X1 U5079 ( .A1(n6125), .A2(n6124), .ZN(n8695) );
  MUX2_X1 U5080 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5082), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5085) );
  AND2_X1 U5081 ( .A1(n6158), .A2(n9619), .ZN(n6163) );
  INV_X2 U5082 ( .A(n9621), .ZN(n9624) );
  MUX2_X1 U5083 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6123), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n6125) );
  INV_X2 U5084 ( .A(n8330), .ZN(n4391) );
  NAND2_X1 U5085 ( .A1(n5253), .A2(n5252), .ZN(n5256) );
  XNOR2_X1 U5086 ( .A(n5231), .B(SI_5_), .ZN(n5452) );
  OAI21_X1 U5087 ( .B1(n5398), .B2(P1_DATAO_REG_8__SCAN_IN), .A(n4531), .ZN(
        n5234) );
  MUX2_X1 U5088 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6156), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n6158) );
  NAND2_X2 U5089 ( .A1(n7388), .A2(P1_U3084), .ZN(n10238) );
  AND2_X1 U5090 ( .A1(n4672), .A2(n5079), .ZN(n5138) );
  NAND2_X1 U5091 ( .A1(n6085), .A2(n4466), .ZN(n6511) );
  BUF_X2 U5092 ( .A(n6101), .Z(n6085) );
  AND2_X1 U5093 ( .A1(n6011), .A2(n6010), .ZN(n6041) );
  AND4_X1 U5094 ( .A1(n4525), .A2(n5113), .A3(n5127), .A4(n5116), .ZN(n5050)
         );
  AND4_X1 U5095 ( .A1(n6009), .A2(n6018), .A3(n6065), .A4(n6026), .ZN(n4735)
         );
  AND4_X1 U5096 ( .A1(n6016), .A2(n4613), .A3(n4612), .A4(n4611), .ZN(n4736)
         );
  INV_X1 U5097 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5127) );
  INV_X1 U5098 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5197) );
  INV_X1 U5099 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6097) );
  NOR2_X1 U5100 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n4613) );
  NAND3_X2 U5101 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n6226) );
  NOR2_X1 U5102 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n4612) );
  INV_X4 U5103 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U5104 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5113) );
  NOR2_X1 U5105 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5049) );
  INV_X1 U5106 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6096) );
  NOR2_X1 U5107 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n4525) );
  INV_X1 U5108 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6026) );
  NOR2_X1 U5109 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6011) );
  INV_X1 U5110 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5090) );
  NOR2_X1 U5111 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6010) );
  INV_X4 U5112 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U5113 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6065) );
  INV_X1 U5114 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6018) );
  INV_X1 U5115 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5108) );
  NAND2_X1 U5116 ( .A1(n7774), .A2(n10489), .ZN(n10457) );
  OAI21_X1 U5117 ( .B1(n7389), .B2(n7409), .A(n5227), .ZN(n5237) );
  OR2_X2 U5118 ( .A1(n9764), .A2(n4899), .ZN(n4898) );
  INV_X1 U5119 ( .A(n7619), .ZN(n7723) );
  OAI21_X1 U5120 ( .B1(n9010), .B2(n6674), .A(n6673), .ZN(n4392) );
  OR2_X1 U5121 ( .A1(n9034), .A2(n9035), .ZN(n4393) );
  NAND2_X1 U5122 ( .A1(n4393), .A2(n9031), .ZN(n6699) );
  OAI21_X1 U5123 ( .B1(n7737), .B2(n7738), .A(n6599), .ZN(n4394) );
  AND2_X1 U5124 ( .A1(n6702), .A2(n6700), .ZN(n9031) );
  AND2_X1 U5125 ( .A1(n6699), .A2(n5035), .ZN(n6706) );
  OAI21_X1 U5126 ( .B1(n7737), .B2(n7738), .A(n6599), .ZN(n7921) );
  NAND2_X1 U5127 ( .A1(n8559), .A2(n4398), .ZN(n4395) );
  AND2_X2 U5128 ( .A1(n4395), .A2(n4396), .ZN(n8741) );
  OR2_X1 U5129 ( .A1(n4397), .A2(n4821), .ZN(n4396) );
  INV_X1 U5130 ( .A(n7023), .ZN(n4397) );
  AND2_X1 U5131 ( .A1(n4824), .A2(n7023), .ZN(n4398) );
  NOR2_X2 U5132 ( .A1(n7845), .A2(n9460), .ZN(n7780) );
  AOI21_X2 U5133 ( .B1(n8759), .B2(n4412), .A(n4470), .ZN(n4865) );
  INV_X4 U5134 ( .A(n5766), .ZN(n5803) );
  NAND2_X1 U5135 ( .A1(n4823), .A2(n4821), .ZN(n4399) );
  AND2_X2 U5136 ( .A1(n5377), .A2(n10235), .ZN(n5465) );
  AND4_X2 U5137 ( .A1(n5062), .A2(n5054), .A3(n5053), .A4(n5052), .ZN(n4439)
         );
  NAND2_X1 U5138 ( .A1(n9626), .A2(n8955), .ZN(n6258) );
  NAND2_X2 U5139 ( .A1(n5423), .A2(n5965), .ZN(n5917) );
  AND2_X1 U5140 ( .A1(n7082), .A2(n4862), .ZN(n5031) );
  XNOR2_X1 U5141 ( .A(n7091), .B(n7153), .ZN(n5872) );
  AOI21_X2 U5142 ( .B1(n9722), .B2(n9721), .A(n9720), .ZN(n9724) );
  XOR2_X2 U5143 ( .A(n8180), .B(n7218), .Z(n4422) );
  NAND2_X1 U5144 ( .A1(n8024), .A2(n4480), .ZN(n4874) );
  INV_X4 U5145 ( .A(n5367), .ZN(n5763) );
  BUF_X1 U5146 ( .A(n9500), .Z(n4400) );
  INV_X2 U5147 ( .A(n5076), .ZN(n5081) );
  NAND2_X2 U5148 ( .A1(n4874), .A2(n4875), .ZN(n8462) );
  NAND2_X1 U5149 ( .A1(n7723), .A2(n7812), .ZN(n8861) );
  INV_X1 U5150 ( .A(n10234), .ZN(n5377) );
  INV_X2 U5151 ( .A(n6197), .ZN(n6382) );
  NAND2_X4 U5152 ( .A1(n8439), .A2(n7620), .ZN(n8865) );
  AND2_X4 U5153 ( .A1(n7619), .A2(n7812), .ZN(n8439) );
  NOR2_X2 U5154 ( .A1(n7798), .A2(n7797), .ZN(n7868) );
  OR2_X1 U5155 ( .A1(n9881), .A2(n5854), .ZN(n4698) );
  INV_X1 U5156 ( .A(n5452), .ZN(n5224) );
  NAND2_X1 U5157 ( .A1(n7411), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4577) );
  INV_X1 U5158 ( .A(n4620), .ZN(n4619) );
  OAI22_X1 U5159 ( .A1(n4926), .A2(n4621), .B1(n9351), .B2(n9026), .ZN(n4620)
         );
  INV_X1 U5160 ( .A(n9515), .ZN(n9266) );
  OR2_X1 U5161 ( .A1(n10107), .A2(n9634), .ZN(n5893) );
  NOR2_X1 U5162 ( .A1(n7144), .A2(n4762), .ZN(n4761) );
  INV_X1 U5163 ( .A(n4764), .ZN(n4762) );
  INV_X1 U5164 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5011) );
  AND2_X1 U5165 ( .A1(n4667), .A2(n5786), .ZN(n4666) );
  NAND2_X1 U5166 ( .A1(n5755), .A2(n5330), .ZN(n4667) );
  AOI21_X1 U5167 ( .B1(n9209), .B2(n4917), .A(n4455), .ZN(n4916) );
  INV_X1 U5168 ( .A(n6470), .ZN(n4917) );
  AOI21_X1 U5169 ( .B1(n4904), .B2(n4716), .A(n4430), .ZN(n4903) );
  INV_X1 U5170 ( .A(n4423), .ZN(n6264) );
  MUX2_X1 U5171 ( .A(n7356), .B(n7357), .S(n7339), .Z(n7214) );
  AND2_X1 U5172 ( .A1(n7123), .A2(n5613), .ZN(n4501) );
  OAI21_X1 U5173 ( .B1(n5773), .B2(n5719), .A(n4695), .ZN(n4701) );
  NAND2_X1 U5174 ( .A1(n4699), .A2(n4688), .ZN(n4687) );
  INV_X1 U5175 ( .A(n4695), .ZN(n4688) );
  AOI21_X1 U5176 ( .B1(n9791), .B2(n5858), .A(n7089), .ZN(n4806) );
  NAND2_X1 U5177 ( .A1(n9849), .A2(n10116), .ZN(n4804) );
  NOR2_X1 U5178 ( .A1(n5589), .A2(n4937), .ZN(n4936) );
  INV_X1 U5179 ( .A(n5271), .ZN(n4937) );
  NAND2_X1 U5180 ( .A1(n5274), .A2(n5273), .ZN(n5277) );
  INV_X1 U5181 ( .A(n6713), .ZN(n4961) );
  INV_X1 U5182 ( .A(n8352), .ZN(n4569) );
  AND2_X1 U5183 ( .A1(n7317), .A2(n7320), .ZN(n7163) );
  NAND2_X1 U5184 ( .A1(n4457), .A2(n6371), .ZN(n4621) );
  OR2_X1 U5185 ( .A1(n9392), .A2(n9105), .ZN(n7268) );
  OR2_X1 U5186 ( .A1(n6337), .A2(n9420), .ZN(n7257) );
  INV_X1 U5187 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6095) );
  NAND2_X1 U5188 ( .A1(n5943), .A2(n10092), .ZN(n4679) );
  OR2_X1 U5189 ( .A1(n10129), .A2(n9887), .ZN(n9881) );
  NAND2_X1 U5190 ( .A1(n7106), .A2(n7105), .ZN(n7107) );
  AND2_X1 U5191 ( .A1(n9806), .A2(n7153), .ZN(n7929) );
  NAND2_X1 U5192 ( .A1(n4499), .A2(n4498), .ZN(n4497) );
  NAND2_X1 U5193 ( .A1(n5387), .A2(n5386), .ZN(n5834) );
  AND2_X1 U5194 ( .A1(n5794), .A2(n5334), .ZN(n5786) );
  NOR2_X1 U5195 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5054) );
  OR2_X1 U5196 ( .A1(n5298), .A2(n5297), .ZN(n5651) );
  AND2_X1 U5197 ( .A1(n5632), .A2(n5296), .ZN(n5297) );
  NAND2_X1 U5198 ( .A1(n5299), .A2(n5287), .ZN(n5653) );
  AOI21_X1 U5199 ( .B1(n4936), .B2(n5272), .A(n4935), .ZN(n4934) );
  INV_X1 U5200 ( .A(n5277), .ZN(n4935) );
  AND2_X1 U5201 ( .A1(n5616), .A2(n5282), .ZN(n5615) );
  NAND2_X1 U5202 ( .A1(n4579), .A2(n4934), .ZN(n5650) );
  NAND2_X1 U5203 ( .A1(n5523), .A2(n4936), .ZN(n4579) );
  INV_X1 U5204 ( .A(n5522), .ZN(n5272) );
  NAND2_X1 U5205 ( .A1(n5268), .A2(n5267), .ZN(n5523) );
  NAND2_X1 U5206 ( .A1(n5479), .A2(n5478), .ZN(n5500) );
  NAND2_X1 U5207 ( .A1(n4958), .A2(n4954), .ZN(n4957) );
  OR2_X1 U5208 ( .A1(n6675), .A2(n6676), .ZN(n4534) );
  AND2_X1 U5209 ( .A1(n7679), .A2(n7176), .ZN(n6349) );
  INV_X1 U5210 ( .A(n6486), .ZN(n6561) );
  INV_X1 U5211 ( .A(n6257), .ZN(n6489) );
  INV_X2 U5212 ( .A(n6258), .ZN(n6555) );
  NAND2_X1 U5213 ( .A1(n6473), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6484) );
  INV_X1 U5214 ( .A(n6475), .ZN(n6473) );
  NOR2_X1 U5215 ( .A1(n9483), .A2(n8916), .ZN(n8915) );
  NAND2_X1 U5216 ( .A1(n9220), .A2(n9446), .ZN(n6564) );
  INV_X1 U5217 ( .A(n9498), .ZN(n6469) );
  OR2_X1 U5218 ( .A1(n9237), .A2(n9252), .ZN(n6454) );
  INV_X1 U5219 ( .A(n9219), .ZN(n9214) );
  INV_X1 U5220 ( .A(n5037), .ZN(n4905) );
  AND2_X1 U5221 ( .A1(n6197), .A2(n4522), .ZN(n6233) );
  INV_X1 U5222 ( .A(n8900), .ZN(n7182) );
  INV_X1 U5223 ( .A(n10507), .ZN(n9588) );
  AND2_X1 U5224 ( .A1(n9638), .A2(n4463), .ZN(n4897) );
  NAND2_X1 U5225 ( .A1(n8756), .A2(n8757), .ZN(n9640) );
  NOR2_X1 U5226 ( .A1(n10083), .A2(n9837), .ZN(n5947) );
  INV_X1 U5227 ( .A(n5762), .ZN(n5824) );
  INV_X1 U5228 ( .A(n4402), .ZN(n5821) );
  XNOR2_X1 U5229 ( .A(n7396), .B(n4588), .ZN(n7437) );
  INV_X1 U5230 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n4588) );
  INV_X1 U5231 ( .A(n7470), .ZN(n4607) );
  INV_X1 U5232 ( .A(n9814), .ZN(n4608) );
  OR2_X1 U5233 ( .A1(n10123), .A2(n9888), .ZN(n9849) );
  OR2_X1 U5234 ( .A1(n5760), .A2(n5759), .ZN(n5778) );
  AOI21_X1 U5235 ( .B1(n7143), .B2(n4765), .A(n4446), .ZN(n4764) );
  INV_X1 U5236 ( .A(n7141), .ZN(n4765) );
  NAND2_X1 U5237 ( .A1(n9905), .A2(n10068), .ZN(n4514) );
  AOI21_X1 U5238 ( .B1(n4792), .B2(n4790), .A(n4452), .ZN(n4789) );
  INV_X1 U5239 ( .A(n4792), .ZN(n4791) );
  NAND2_X1 U5240 ( .A1(n8619), .A2(n4767), .ZN(n4770) );
  AOI21_X1 U5241 ( .B1(n4773), .B2(n7117), .A(n4772), .ZN(n4769) );
  NOR2_X1 U5242 ( .A1(n10061), .A2(n9794), .ZN(n4772) );
  NOR2_X1 U5243 ( .A1(n4774), .A2(n7119), .ZN(n4773) );
  INV_X1 U5244 ( .A(n7118), .ZN(n4774) );
  NAND2_X1 U5245 ( .A1(n4784), .A2(n4780), .ZN(n10103) );
  INV_X1 U5246 ( .A(n4781), .ZN(n4780) );
  OAI211_X1 U5247 ( .C1(n4783), .C2(n4782), .A(n8935), .B(n4787), .ZN(n4781)
         );
  AND2_X1 U5248 ( .A1(n7065), .A2(n5057), .ZN(n4862) );
  AND2_X1 U5249 ( .A1(n5742), .A2(n5318), .ZN(n5731) );
  NAND2_X1 U5250 ( .A1(n8691), .A2(n7176), .ZN(n6472) );
  NAND2_X2 U5251 ( .A1(n6706), .A2(n6705), .ZN(n9084) );
  NAND2_X1 U5252 ( .A1(n9033), .A2(n6704), .ZN(n6705) );
  OR2_X1 U5253 ( .A1(n9488), .A2(n9204), .ZN(n8904) );
  INV_X1 U5254 ( .A(n8912), .ZN(n8913) );
  AOI22_X1 U5255 ( .A1(n9204), .A2(n9446), .B1(n8911), .B2(n9112), .ZN(n8912)
         );
  NOR3_X1 U5256 ( .A1(n7208), .A2(n6525), .A3(n7214), .ZN(n7209) );
  MUX2_X1 U5257 ( .A(n7207), .B(n7206), .S(n7339), .Z(n7208) );
  AND2_X1 U5258 ( .A1(n4725), .A2(n7339), .ZN(n4720) );
  AOI21_X1 U5259 ( .B1(n4517), .B2(n7240), .A(n7239), .ZN(n7249) );
  NAND2_X1 U5260 ( .A1(n5443), .A2(n5444), .ZN(n5474) );
  OAI21_X1 U5261 ( .B1(n8101), .B2(n5972), .A(n7089), .ZN(n5444) );
  NAND2_X1 U5262 ( .A1(n4685), .A2(n7089), .ZN(n4684) );
  INV_X1 U5263 ( .A(n8262), .ZN(n4685) );
  AND2_X1 U5264 ( .A1(n7101), .A2(n5919), .ZN(n4686) );
  OR2_X1 U5265 ( .A1(n7249), .A2(n7242), .ZN(n7246) );
  OR2_X1 U5266 ( .A1(n7247), .A2(n6540), .ZN(n7242) );
  NOR2_X1 U5267 ( .A1(n9279), .A2(n7282), .ZN(n4718) );
  AND2_X1 U5268 ( .A1(n4730), .A2(n4729), .ZN(n4728) );
  NAND2_X1 U5269 ( .A1(n4429), .A2(n4502), .ZN(n5776) );
  NOR2_X1 U5270 ( .A1(n4734), .A2(n4733), .ZN(n7324) );
  OR2_X1 U5271 ( .A1(n7319), .A2(n7321), .ZN(n4733) );
  INV_X1 U5272 ( .A(n7107), .ZN(n4798) );
  INV_X1 U5273 ( .A(n7109), .ZN(n4801) );
  NAND2_X1 U5274 ( .A1(n5285), .A2(n5284), .ZN(n5299) );
  NAND2_X1 U5275 ( .A1(n5260), .A2(n5259), .ZN(n5263) );
  OAI21_X1 U5276 ( .B1(n5398), .B2(n4539), .A(n4538), .ZN(n5480) );
  NAND2_X1 U5277 ( .A1(n4382), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n4538) );
  OAI21_X1 U5278 ( .B1(n5398), .B2(n5219), .A(n5218), .ZN(n5221) );
  NAND2_X1 U5279 ( .A1(n5398), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5218) );
  NAND2_X1 U5280 ( .A1(n6680), .A2(n6681), .ZN(n4976) );
  NAND2_X1 U5281 ( .A1(n7168), .A2(n7370), .ZN(n4989) );
  NOR2_X1 U5282 ( .A1(n7998), .A2(n4944), .ZN(n7189) );
  AND2_X1 U5283 ( .A1(n4564), .A2(n4562), .ZN(n7535) );
  INV_X1 U5284 ( .A(n7574), .ZN(n4562) );
  NAND2_X1 U5285 ( .A1(n7576), .A2(n7575), .ZN(n4564) );
  AOI22_X1 U5286 ( .A1(n9126), .A2(n9127), .B1(n6332), .B2(n9133), .ZN(n6074)
         );
  AND2_X1 U5287 ( .A1(n9483), .A2(n7165), .ZN(n7166) );
  NOR2_X1 U5288 ( .A1(n9483), .A2(n7165), .ZN(n7330) );
  OR2_X1 U5289 ( .A1(n9493), .A2(n9498), .ZN(n4860) );
  OR2_X1 U5290 ( .A1(n9498), .A2(n6468), .ZN(n7309) );
  NOR2_X1 U5291 ( .A1(n4855), .A2(n9520), .ZN(n4853) );
  NOR2_X1 U5292 ( .A1(n6549), .A2(n6548), .ZN(n6550) );
  NAND2_X1 U5293 ( .A1(n4619), .A2(n4621), .ZN(n4618) );
  NAND2_X1 U5294 ( .A1(n6573), .A2(n4856), .ZN(n4855) );
  NAND2_X1 U5295 ( .A1(n9321), .A2(n4431), .ZN(n4910) );
  AND2_X1 U5296 ( .A1(n9278), .A2(n7281), .ZN(n7365) );
  AND2_X1 U5297 ( .A1(n4549), .A2(n7274), .ZN(n4546) );
  AOI21_X1 U5298 ( .B1(n4549), .B2(n7269), .A(n4548), .ZN(n4547) );
  INV_X1 U5299 ( .A(n9371), .ZN(n4548) );
  AND2_X1 U5300 ( .A1(n9357), .A2(n9367), .ZN(n4926) );
  NOR2_X1 U5301 ( .A1(n6356), .A2(n6355), .ZN(n4542) );
  NAND2_X1 U5302 ( .A1(n6289), .A2(n8299), .ZN(n6279) );
  NAND2_X1 U5303 ( .A1(n9443), .A2(n8196), .ZN(n7213) );
  NAND2_X1 U5304 ( .A1(n7923), .A2(n9440), .ZN(n7188) );
  NAND2_X1 U5305 ( .A1(n6600), .A2(n7922), .ZN(n7211) );
  NAND2_X1 U5306 ( .A1(n7924), .A2(n8189), .ZN(n7197) );
  OAI22_X1 U5307 ( .A1(n8925), .A2(n4401), .B1(n8092), .B2(n8012), .ZN(n7788)
         );
  INV_X1 U5308 ( .A(n9775), .ZN(n4869) );
  INV_X1 U5309 ( .A(n7890), .ZN(n4640) );
  OR3_X1 U5310 ( .A1(n5818), .A2(n9633), .A3(n8880), .ZN(n5819) );
  INV_X1 U5311 ( .A(n5724), .ZN(n5375) );
  NOR2_X1 U5312 ( .A1(n9902), .A2(n4700), .ZN(n4829) );
  OR2_X1 U5313 ( .A1(n10127), .A2(n9871), .ZN(n5935) );
  AND2_X1 U5314 ( .A1(n5859), .A2(n7039), .ZN(n7139) );
  NOR2_X1 U5315 ( .A1(n10156), .A2(n10159), .ZN(n5023) );
  INV_X1 U5316 ( .A(n10165), .ZN(n5612) );
  NAND2_X1 U5317 ( .A1(n10165), .A2(n10041), .ZN(n7029) );
  NAND2_X1 U5318 ( .A1(n8559), .A2(n7021), .ZN(n8624) );
  AOI21_X1 U5319 ( .B1(n4824), .B2(n4827), .A(n4822), .ZN(n4821) );
  NAND2_X1 U5320 ( .A1(n8559), .A2(n4824), .ZN(n4823) );
  INV_X1 U5321 ( .A(n7022), .ZN(n4827) );
  OR2_X1 U5322 ( .A1(n10193), .A2(n10072), .ZN(n5861) );
  INV_X1 U5323 ( .A(n8076), .ZN(n7101) );
  NAND2_X1 U5324 ( .A1(n8101), .A2(n4426), .ZN(n8068) );
  NAND2_X1 U5325 ( .A1(n5655), .A2(n7399), .ZN(n4675) );
  INV_X1 U5326 ( .A(n7148), .ZN(n4782) );
  INV_X1 U5327 ( .A(n5330), .ZN(n4664) );
  INV_X1 U5328 ( .A(n5794), .ZN(n4663) );
  NOR2_X1 U5329 ( .A1(n4665), .A2(n4660), .ZN(n4659) );
  INV_X1 U5330 ( .A(n5324), .ZN(n4660) );
  INV_X1 U5331 ( .A(n4666), .ZN(n4665) );
  INV_X1 U5332 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4756) );
  NAND2_X1 U5333 ( .A1(n4647), .A2(n5731), .ZN(n4646) );
  NAND2_X1 U5334 ( .A1(n4650), .A2(n4652), .ZN(n4647) );
  NAND2_X1 U5335 ( .A1(n5310), .A2(n5309), .ZN(n5313) );
  NOR2_X1 U5336 ( .A1(n5308), .A2(n4655), .ZN(n4654) );
  INV_X1 U5337 ( .A(n5303), .ZN(n4655) );
  INV_X1 U5338 ( .A(n5706), .ZN(n5308) );
  XNOR2_X1 U5339 ( .A(n5305), .B(SI_21_), .ZN(n5706) );
  NAND2_X1 U5340 ( .A1(n4530), .A2(n4528), .ZN(n5691) );
  NOR2_X1 U5341 ( .A1(n4442), .A2(n4529), .ZN(n4528) );
  NAND2_X1 U5342 ( .A1(n5650), .A2(n5289), .ZN(n4530) );
  INV_X1 U5343 ( .A(n5299), .ZN(n4529) );
  AND2_X1 U5344 ( .A1(n5303), .A2(n5302), .ZN(n5690) );
  AND2_X1 U5345 ( .A1(n5615), .A2(n5291), .ZN(n5634) );
  OR2_X1 U5346 ( .A1(n5294), .A2(n5293), .ZN(n5632) );
  AND2_X1 U5347 ( .A1(n5616), .A2(n5618), .ZN(n5293) );
  INV_X1 U5348 ( .A(n4936), .ZN(n4932) );
  INV_X1 U5349 ( .A(n5615), .ZN(n4931) );
  NOR2_X1 U5350 ( .A1(n4933), .A2(n4929), .ZN(n4928) );
  INV_X1 U5351 ( .A(n5267), .ZN(n4929) );
  INV_X1 U5352 ( .A(n4934), .ZN(n4933) );
  AOI21_X1 U5353 ( .B1(n5034), .B2(n4924), .A(n4923), .ZN(n4922) );
  INV_X1 U5354 ( .A(n5250), .ZN(n4924) );
  INV_X1 U5355 ( .A(n5256), .ZN(n4923) );
  INV_X1 U5356 ( .A(n5034), .ZN(n4925) );
  AND3_X1 U5357 ( .A1(n4453), .A2(n5242), .A3(n5240), .ZN(n4537) );
  NAND2_X1 U5358 ( .A1(n5244), .A2(n5236), .ZN(n5503) );
  INV_X1 U5359 ( .A(n5234), .ZN(n5235) );
  NOR2_X2 U5360 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5118) );
  NAND2_X1 U5361 ( .A1(n5217), .A2(n5216), .ZN(n5439) );
  OR2_X1 U5362 ( .A1(n5118), .A2(n5143), .ZN(n5122) );
  OR2_X1 U5363 ( .A1(n6319), .A2(n6307), .ZN(n6330) );
  INV_X1 U5364 ( .A(n7391), .ZN(n4616) );
  AOI21_X1 U5365 ( .B1(n4960), .B2(n4962), .A(n4959), .ZN(n4958) );
  INV_X1 U5366 ( .A(n6727), .ZN(n4959) );
  NAND2_X1 U5367 ( .A1(n6239), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6270) );
  INV_X1 U5368 ( .A(n6241), .ZN(n6239) );
  NAND2_X1 U5369 ( .A1(n6306), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6319) );
  INV_X1 U5370 ( .A(n6317), .ZN(n6306) );
  OR2_X1 U5371 ( .A1(n9009), .A2(n9011), .ZN(n6672) );
  NAND2_X1 U5372 ( .A1(n4540), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6282) );
  INV_X1 U5373 ( .A(n6272), .ZN(n4540) );
  INV_X1 U5374 ( .A(n8975), .ZN(n4967) );
  NAND2_X1 U5375 ( .A1(n4969), .A2(n4976), .ZN(n4968) );
  INV_X1 U5376 ( .A(n4974), .ZN(n4969) );
  AOI21_X1 U5377 ( .B1(n9024), .B2(n4977), .A(n4975), .ZN(n4974) );
  INV_X1 U5378 ( .A(n9077), .ZN(n4975) );
  NOR2_X1 U5379 ( .A1(n4967), .A2(n4972), .ZN(n4964) );
  NAND2_X1 U5380 ( .A1(n6224), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6241) );
  INV_X1 U5381 ( .A(n6226), .ZN(n6224) );
  INV_X1 U5382 ( .A(n9443), .ZN(n7915) );
  NOR2_X1 U5383 ( .A1(n6736), .A2(n10472), .ZN(n6734) );
  OAI21_X1 U5385 ( .B1(n6175), .B2(P2_REG1_REG_2__SCAN_IN), .A(n4563), .ZN(
        n7574) );
  NAND2_X1 U5386 ( .A1(n6175), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4563) );
  INV_X1 U5387 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6029) );
  NAND2_X1 U5388 ( .A1(n7596), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4752) );
  OAI22_X1 U5389 ( .A1(n7593), .A2(n4751), .B1(n7638), .B2(n4752), .ZN(n7637)
         );
  OR2_X1 U5390 ( .A1(n7592), .A2(n7638), .ZN(n4751) );
  OR2_X1 U5391 ( .A1(n7593), .A2(n7592), .ZN(n4753) );
  NAND2_X1 U5392 ( .A1(n4574), .A2(n4577), .ZN(n4571) );
  NAND2_X1 U5393 ( .A1(n4576), .A2(n4577), .ZN(n4572) );
  OR2_X1 U5394 ( .A1(n8708), .A2(n8709), .ZN(n4750) );
  AND2_X1 U5395 ( .A1(n8720), .A2(n4481), .ZN(n4749) );
  NAND2_X1 U5396 ( .A1(n9141), .A2(n9140), .ZN(n9139) );
  AND2_X1 U5397 ( .A1(n6141), .A2(n6140), .ZN(n9171) );
  MUX2_X1 U5398 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6118), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n6119) );
  OR2_X1 U5399 ( .A1(n7998), .A2(n4384), .ZN(n6728) );
  AND2_X1 U5400 ( .A1(n4914), .A2(n7369), .ZN(n4913) );
  NAND2_X1 U5401 ( .A1(n4916), .A2(n4992), .ZN(n4914) );
  NAND2_X1 U5402 ( .A1(n4990), .A2(n4656), .ZN(n7164) );
  AND2_X1 U5403 ( .A1(n4657), .A2(n7318), .ZN(n4656) );
  NAND2_X1 U5404 ( .A1(n9229), .A2(n4991), .ZN(n4990) );
  INV_X1 U5405 ( .A(n7163), .ZN(n7369) );
  AND2_X1 U5406 ( .A1(n7309), .A2(n7311), .ZN(n9219) );
  AND2_X1 U5407 ( .A1(n9219), .A2(n7308), .ZN(n4996) );
  NAND2_X1 U5408 ( .A1(n6458), .A2(n6457), .ZN(n6475) );
  NAND2_X1 U5409 ( .A1(n4903), .A2(n4902), .ZN(n4901) );
  OR2_X1 U5410 ( .A1(n9266), .A2(n9070), .ZN(n5037) );
  NAND2_X1 U5411 ( .A1(n6424), .A2(n6422), .ZN(n7293) );
  NOR2_X1 U5412 ( .A1(n9261), .A2(n5003), .ZN(n5002) );
  INV_X1 U5413 ( .A(n7293), .ZN(n5003) );
  NAND2_X1 U5414 ( .A1(n9259), .A2(n9261), .ZN(n9258) );
  NAND2_X1 U5415 ( .A1(n6551), .A2(n6550), .ZN(n9280) );
  NAND2_X1 U5416 ( .A1(n4912), .A2(n4404), .ZN(n4911) );
  AND2_X1 U5417 ( .A1(n4550), .A2(n7268), .ZN(n4549) );
  OR2_X1 U5418 ( .A1(n7269), .A2(n7264), .ZN(n4550) );
  NAND2_X1 U5419 ( .A1(n7274), .A2(n7275), .ZN(n9357) );
  NAND2_X2 U5420 ( .A1(n4506), .A2(n6352), .ZN(n9392) );
  NAND2_X1 U5421 ( .A1(n7704), .A2(n7176), .ZN(n4506) );
  AND2_X1 U5422 ( .A1(n6339), .A2(n6338), .ZN(n6340) );
  OR2_X1 U5423 ( .A1(n6337), .A2(n9400), .ZN(n6338) );
  AND2_X1 U5424 ( .A1(n7264), .A2(n7263), .ZN(n9409) );
  INV_X1 U5425 ( .A(n9119), .ZN(n8209) );
  INV_X1 U5426 ( .A(n9385), .ZN(n9263) );
  INV_X1 U5427 ( .A(n9418), .ZN(n9446) );
  INV_X1 U5428 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7564) );
  INV_X1 U5429 ( .A(n9263), .ZN(n10460) );
  NAND2_X1 U5430 ( .A1(n7179), .A2(n7178), .ZN(n9478) );
  NAND2_X1 U5431 ( .A1(n6495), .A2(n6494), .ZN(n9488) );
  NAND2_X1 U5432 ( .A1(n6384), .A2(n6383), .ZN(n9535) );
  NAND2_X1 U5433 ( .A1(n6294), .A2(n6293), .ZN(n9574) );
  INV_X1 U5434 ( .A(n9440), .ZN(n10494) );
  OR2_X1 U5435 ( .A1(n7187), .A2(n7355), .ZN(n10508) );
  NAND2_X1 U5436 ( .A1(n6518), .A2(n6517), .ZN(n7674) );
  NOR2_X1 U5437 ( .A1(n6759), .A2(n6758), .ZN(n7676) );
  NAND2_X1 U5438 ( .A1(n6738), .A2(n10487), .ZN(n10472) );
  AND3_X1 U5439 ( .A1(n6101), .A2(n5005), .A3(n6100), .ZN(n6159) );
  AND2_X1 U5440 ( .A1(n5008), .A2(n5006), .ZN(n5005) );
  INV_X1 U5441 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5006) );
  XNOR2_X1 U5442 ( .A(n4560), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6210) );
  OR2_X1 U5443 ( .A1(n6041), .A2(n6033), .ZN(n4560) );
  NAND2_X1 U5444 ( .A1(n7564), .A2(n4737), .ZN(n6039) );
  INV_X1 U5445 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4737) );
  NOR2_X1 U5446 ( .A1(n9630), .A2(n9631), .ZN(n4896) );
  INV_X1 U5447 ( .A(n4877), .ZN(n4876) );
  OAI21_X1 U5448 ( .B1(n8338), .B2(n4878), .A(n8276), .ZN(n4877) );
  NAND2_X1 U5449 ( .A1(n5373), .A2(n4818), .ZN(n5624) );
  NAND2_X1 U5450 ( .A1(n8780), .A2(n4884), .ZN(n4883) );
  NOR2_X1 U5451 ( .A1(n8798), .A2(n4885), .ZN(n4884) );
  INV_X1 U5452 ( .A(n8779), .ZN(n4885) );
  NOR2_X1 U5453 ( .A1(n8598), .A2(n4872), .ZN(n4871) );
  INV_X1 U5454 ( .A(n8587), .ZN(n4872) );
  OR2_X1 U5455 ( .A1(n5711), .A2(n5710), .ZN(n5724) );
  NAND2_X1 U5456 ( .A1(n5375), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5735) );
  NOR2_X1 U5457 ( .A1(n8822), .A2(n4880), .ZN(n4879) );
  INV_X1 U5458 ( .A(n8817), .ZN(n4880) );
  AND2_X1 U5459 ( .A1(n10225), .A2(n7813), .ZN(n7615) );
  OR2_X1 U5460 ( .A1(n9762), .A2(n9763), .ZN(n4899) );
  NAND2_X1 U5461 ( .A1(n8759), .A2(n8758), .ZN(n9641) );
  NAND2_X1 U5462 ( .A1(n9640), .A2(n9643), .ZN(n4870) );
  NAND2_X1 U5463 ( .A1(n5469), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5391) );
  NOR2_X1 U5464 ( .A1(n7438), .A2(n4434), .ZN(n10308) );
  NOR2_X1 U5465 ( .A1(n10307), .A2(n10308), .ZN(n10306) );
  NAND2_X1 U5466 ( .A1(n4599), .A2(n4597), .ZN(n7455) );
  AOI21_X1 U5467 ( .B1(n4601), .B2(n4600), .A(n4598), .ZN(n4597) );
  NAND2_X1 U5468 ( .A1(n4596), .A2(n4595), .ZN(n4599) );
  AND2_X1 U5469 ( .A1(n9812), .A2(n9811), .ZN(n9809) );
  INV_X1 U5470 ( .A(n5165), .ZN(n4610) );
  OAI21_X1 U5471 ( .B1(n9809), .B2(n7490), .A(n7491), .ZN(n7489) );
  NAND2_X1 U5472 ( .A1(n7523), .A2(n4641), .ZN(n7520) );
  NOR2_X1 U5473 ( .A1(n4643), .A2(n4642), .ZN(n4641) );
  INV_X1 U5474 ( .A(n7522), .ZN(n4643) );
  INV_X1 U5475 ( .A(n7521), .ZN(n4642) );
  NAND2_X1 U5476 ( .A1(n4636), .A2(n4640), .ZN(n4635) );
  INV_X1 U5477 ( .A(n4637), .ZN(n4636) );
  AOI21_X1 U5478 ( .B1(n7653), .B2(n7654), .A(n4638), .ZN(n4637) );
  INV_X1 U5479 ( .A(n7891), .ZN(n4638) );
  OAI21_X1 U5480 ( .B1(n7655), .B2(n7654), .A(n7653), .ZN(n7892) );
  AND2_X1 U5481 ( .A1(n4640), .A2(n7653), .ZN(n4634) );
  NAND2_X1 U5482 ( .A1(n7655), .A2(n4634), .ZN(n4633) );
  OR2_X1 U5483 ( .A1(n7887), .A2(n4594), .ZN(n4593) );
  AND2_X1 U5484 ( .A1(n7896), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4594) );
  XNOR2_X1 U5485 ( .A(n5156), .B(n5173), .ZN(n10319) );
  NOR2_X1 U5486 ( .A1(n8426), .A2(n4644), .ZN(n5156) );
  AND2_X1 U5487 ( .A1(n8425), .A2(n5155), .ZN(n4644) );
  NAND2_X1 U5488 ( .A1(n10319), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n10318) );
  NOR2_X1 U5489 ( .A1(n8423), .A2(n5172), .ZN(n5174) );
  INV_X1 U5490 ( .A(n5020), .ZN(n9842) );
  NAND2_X1 U5491 ( .A1(n5390), .A2(n5389), .ZN(n10093) );
  AND2_X1 U5492 ( .A1(n4416), .A2(n9877), .ZN(n5024) );
  AOI21_X1 U5493 ( .B1(n4761), .B2(n4766), .A(n4454), .ZN(n4759) );
  NAND2_X1 U5494 ( .A1(n5375), .A2(n4814), .ZN(n5748) );
  AND2_X1 U5495 ( .A1(n5769), .A2(n5768), .ZN(n9888) );
  NAND2_X1 U5496 ( .A1(n5935), .A2(n9868), .ZN(n9886) );
  INV_X1 U5497 ( .A(n7143), .ZN(n4766) );
  NAND2_X1 U5498 ( .A1(n9925), .A2(n7039), .ZN(n9918) );
  NAND2_X1 U5499 ( .A1(n9931), .A2(n9916), .ZN(n9910) );
  NOR2_X1 U5500 ( .A1(n7138), .A2(n4796), .ZN(n4795) );
  INV_X1 U5501 ( .A(n7135), .ZN(n4796) );
  OR2_X1 U5502 ( .A1(n10146), .A2(n9970), .ZN(n7137) );
  NOR2_X1 U5503 ( .A1(n7139), .A2(n4793), .ZN(n4792) );
  INV_X1 U5504 ( .A(n7137), .ZN(n4793) );
  NAND2_X1 U5505 ( .A1(n5067), .A2(n5055), .ZN(n5185) );
  INV_X1 U5506 ( .A(n5183), .ZN(n5067) );
  NAND2_X1 U5507 ( .A1(n10025), .A2(n7128), .ZN(n9995) );
  OR2_X1 U5508 ( .A1(n7114), .A2(n8620), .ZN(n7116) );
  OR2_X1 U5509 ( .A1(n8323), .A2(n10427), .ZN(n8379) );
  NAND2_X1 U5510 ( .A1(n8316), .A2(n8315), .ZN(n8314) );
  NAND2_X1 U5511 ( .A1(n6236), .A2(n5800), .ZN(n5482) );
  OAI211_X1 U5512 ( .C1(n7931), .C2(n7093), .A(n7092), .B(n7938), .ZN(n7934)
         );
  AND2_X1 U5513 ( .A1(n9808), .A2(n7982), .ZN(n7724) );
  INV_X1 U5514 ( .A(n5872), .ZN(n7726) );
  NAND2_X1 U5515 ( .A1(n5847), .A2(n5846), .ZN(n10083) );
  NAND2_X1 U5516 ( .A1(n5789), .A2(n5788), .ZN(n10116) );
  OR2_X1 U5517 ( .A1(n7971), .A2(n7941), .ZN(n10400) );
  OR2_X1 U5518 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n5359) );
  XNOR2_X1 U5519 ( .A(n5787), .B(n5786), .ZN(n8685) );
  OAI21_X1 U5520 ( .B1(n5756), .B2(n5755), .A(n5330), .ZN(n5787) );
  NAND2_X1 U5521 ( .A1(n4653), .A2(n5307), .ZN(n4652) );
  INV_X1 U5522 ( .A(n5720), .ZN(n4653) );
  INV_X1 U5523 ( .A(n4651), .ZN(n4650) );
  OAI21_X1 U5524 ( .B1(n4654), .B2(n4652), .A(n5313), .ZN(n4651) );
  XNOR2_X1 U5525 ( .A(n5707), .B(n5706), .ZN(n7996) );
  NAND2_X1 U5526 ( .A1(n5304), .A2(n5303), .ZN(n5707) );
  OAI21_X1 U5527 ( .B1(n5523), .B2(n5272), .A(n5271), .ZN(n5588) );
  NAND2_X1 U5528 ( .A1(n6364), .A2(n6363), .ZN(n9545) );
  NAND2_X1 U5529 ( .A1(n6437), .A2(n6436), .ZN(n9508) );
  NAND2_X1 U5530 ( .A1(n9045), .A2(n6611), .ZN(n4980) );
  AND2_X1 U5531 ( .A1(n6739), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9102) );
  NAND2_X1 U5532 ( .A1(n6623), .A2(n6621), .ZN(n7913) );
  INV_X1 U5533 ( .A(n9092), .ZN(n9106) );
  INV_X1 U5534 ( .A(n4520), .ZN(n4519) );
  OAI21_X1 U5535 ( .B1(n7346), .B2(n10488), .A(n7981), .ZN(n4520) );
  OR2_X1 U5536 ( .A1(n8964), .A2(n6561), .ZN(n6482) );
  NAND2_X1 U5537 ( .A1(n6453), .A2(n6452), .ZN(n9252) );
  NAND2_X1 U5538 ( .A1(n6445), .A2(n6444), .ZN(n9114) );
  XNOR2_X1 U5539 ( .A(n7568), .B(n6037), .ZN(n7561) );
  INV_X1 U5540 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6037) );
  NOR2_X1 U5541 ( .A1(n9183), .A2(n9182), .ZN(n9181) );
  NAND2_X1 U5542 ( .A1(n4739), .A2(n4738), .ZN(n6147) );
  NAND2_X1 U5543 ( .A1(n6150), .A2(n9169), .ZN(n4738) );
  NAND2_X1 U5544 ( .A1(n6148), .A2(n9163), .ZN(n4739) );
  OR2_X1 U5545 ( .A1(n6484), .A2(n6483), .ZN(n8918) );
  AOI21_X1 U5546 ( .B1(n4553), .B2(n9385), .A(n4551), .ZN(n9495) );
  INV_X1 U5547 ( .A(n4552), .ZN(n4551) );
  XNOR2_X1 U5548 ( .A(n4554), .B(n4992), .ZN(n4553) );
  AOI22_X1 U5549 ( .A1(n9204), .A2(n9444), .B1(n9446), .B2(n9203), .ZN(n4552)
         );
  NAND2_X1 U5550 ( .A1(n9210), .A2(n9209), .ZN(n9208) );
  NAND2_X1 U5551 ( .A1(n6427), .A2(n6426), .ZN(n9515) );
  NAND2_X1 U5552 ( .A1(n6577), .A2(n9290), .ZN(n9457) );
  OAI211_X1 U5553 ( .C1(n9486), .C2(n9579), .A(n9485), .B(n4671), .ZN(n9596)
         );
  NOR2_X1 U5554 ( .A1(n4411), .A2(n4441), .ZN(n4671) );
  INV_X1 U5555 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6033) );
  NOR2_X1 U5556 ( .A1(n4891), .A2(n4889), .ZN(n4888) );
  INV_X1 U5557 ( .A(n4896), .ZN(n4889) );
  NAND2_X1 U5558 ( .A1(n4895), .A2(n9630), .ZN(n4894) );
  INV_X1 U5559 ( .A(n4899), .ZN(n4895) );
  NAND2_X1 U5560 ( .A1(n9630), .A2(n9631), .ZN(n4893) );
  NAND2_X1 U5561 ( .A1(n5734), .A2(n5733), .ZN(n10129) );
  INV_X1 U5562 ( .A(n9903), .ZN(n9930) );
  INV_X1 U5563 ( .A(n9905), .ZN(n9871) );
  OR2_X1 U5564 ( .A1(n7819), .A2(n7616), .ZN(n9683) );
  NAND2_X1 U5565 ( .A1(n5785), .A2(n5784), .ZN(n9791) );
  OR2_X1 U5566 ( .A1(n9863), .A2(n5821), .ZN(n5785) );
  NOR2_X1 U5567 ( .A1(n7511), .A2(n4589), .ZN(n7652) );
  AND2_X1 U5568 ( .A1(n7425), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4589) );
  NAND2_X1 U5569 ( .A1(n7652), .A2(n7651), .ZN(n7650) );
  NOR2_X1 U5570 ( .A1(n7889), .A2(n7888), .ZN(n7887) );
  XNOR2_X1 U5571 ( .A(n4626), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n5188) );
  NAND2_X1 U5572 ( .A1(n4628), .A2(n4627), .ZN(n4626) );
  NAND2_X1 U5573 ( .A1(n9827), .A2(n5644), .ZN(n4627) );
  INV_X1 U5574 ( .A(n8950), .ZN(n4494) );
  NAND2_X1 U5575 ( .A1(n4778), .A2(n4444), .ZN(n8936) );
  NAND2_X1 U5576 ( .A1(n4835), .A2(n4833), .ZN(n10121) );
  INV_X1 U5577 ( .A(n4834), .ZN(n4833) );
  NAND2_X1 U5578 ( .A1(n4836), .A2(n10074), .ZN(n4835) );
  OAI22_X1 U5579 ( .A1(n9872), .A2(n10040), .B1(n10071), .B2(n9871), .ZN(n4834) );
  AOI21_X1 U5580 ( .B1(n9904), .B2(n10074), .A(n4512), .ZN(n10132) );
  NAND2_X1 U5581 ( .A1(n4514), .A2(n4513), .ZN(n4512) );
  NAND2_X1 U5582 ( .A1(n9903), .A2(n10011), .ZN(n4513) );
  NAND2_X1 U5583 ( .A1(n7142), .A2(n7141), .ZN(n9894) );
  NAND3_X1 U5584 ( .A1(n10184), .A2(n10225), .A3(n5946), .ZN(n10049) );
  OR2_X1 U5585 ( .A1(n10020), .A2(n7943), .ZN(n10063) );
  NAND2_X1 U5586 ( .A1(n10078), .A2(n7613), .ZN(n9999) );
  INV_X1 U5587 ( .A(n10063), .ZN(n10007) );
  OR2_X1 U5588 ( .A1(n7216), .A2(n7339), .ZN(n4724) );
  AND2_X1 U5589 ( .A1(n4686), .A2(n4683), .ZN(n4682) );
  NAND2_X1 U5590 ( .A1(n4425), .A2(n5854), .ZN(n4683) );
  AND2_X1 U5591 ( .A1(n7246), .A2(n7245), .ZN(n7261) );
  INV_X1 U5592 ( .A(n9357), .ZN(n7273) );
  INV_X1 U5593 ( .A(n7278), .ZN(n4730) );
  AND2_X1 U5594 ( .A1(n4711), .A2(n4472), .ZN(n4710) );
  INV_X1 U5595 ( .A(n7283), .ZN(n4712) );
  AOI21_X1 U5596 ( .B1(n4710), .B2(n4713), .A(n4709), .ZN(n4708) );
  INV_X1 U5597 ( .A(n4718), .ZN(n4713) );
  AOI21_X1 U5598 ( .B1(n4708), .B2(n4706), .A(n7339), .ZN(n4705) );
  INV_X1 U5599 ( .A(n4710), .ZN(n4706) );
  AND2_X1 U5600 ( .A1(n7292), .A2(n4714), .ZN(n4703) );
  NOR2_X1 U5601 ( .A1(n4709), .A2(n4715), .ZN(n4714) );
  NAND2_X1 U5602 ( .A1(n4518), .A2(n7339), .ZN(n4715) );
  AND2_X1 U5603 ( .A1(n4702), .A2(n4696), .ZN(n4695) );
  NAND2_X1 U5604 ( .A1(n7039), .A2(n4697), .ZN(n4696) );
  INV_X1 U5605 ( .A(n5899), .ZN(n4702) );
  AND2_X1 U5606 ( .A1(n5703), .A2(n5702), .ZN(n5704) );
  NAND2_X1 U5607 ( .A1(n4693), .A2(n4692), .ZN(n4691) );
  NAND2_X1 U5608 ( .A1(n4694), .A2(n5934), .ZN(n4693) );
  INV_X1 U5609 ( .A(n4698), .ZN(n4694) );
  NAND2_X1 U5610 ( .A1(n4805), .A2(n4803), .ZN(n5807) );
  NAND2_X1 U5611 ( .A1(n7048), .A2(n4806), .ZN(n4805) );
  NOR2_X1 U5612 ( .A1(n8544), .A2(n8538), .ZN(n6289) );
  OR2_X1 U5613 ( .A1(n6251), .A2(n8116), .ZN(n6253) );
  AND2_X1 U5614 ( .A1(n10471), .A2(n6510), .ZN(n6721) );
  NOR2_X1 U5615 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n4611) );
  AOI21_X1 U5616 ( .B1(n7022), .B2(n4826), .A(n4825), .ZN(n4824) );
  INV_X1 U5617 ( .A(n7021), .ZN(n4826) );
  INV_X1 U5618 ( .A(n5387), .ZN(n4499) );
  INV_X1 U5619 ( .A(n5356), .ZN(n4498) );
  AND2_X1 U5620 ( .A1(n5649), .A2(n5288), .ZN(n5289) );
  INV_X1 U5621 ( .A(SI_10_), .ZN(n5252) );
  INV_X1 U5622 ( .A(n5480), .ZN(n5230) );
  NAND2_X1 U5623 ( .A1(n7389), .A2(n7422), .ZN(n4531) );
  INV_X1 U5624 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4940) );
  INV_X1 U5625 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4941) );
  INV_X1 U5626 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4942) );
  NOR2_X1 U5627 ( .A1(n6404), .A2(n6403), .ZN(n4541) );
  INV_X1 U5628 ( .A(n6691), .ZN(n6694) );
  OR3_X1 U5629 ( .A1(n6721), .A2(n7674), .A3(n6757), .ZN(n6736) );
  AOI21_X1 U5630 ( .B1(n7336), .B2(n7335), .A(n7334), .ZN(n7338) );
  AOI211_X1 U5631 ( .C1(n7329), .C2(n7328), .A(n7327), .B(n7326), .ZN(n7345)
         );
  OR2_X1 U5632 ( .A1(n6228), .A2(n9459), .ZN(n6165) );
  AND2_X1 U5633 ( .A1(n4993), .A2(n4992), .ZN(n4991) );
  AOI21_X1 U5634 ( .B1(n4996), .B2(n4994), .A(n7303), .ZN(n4993) );
  INV_X1 U5635 ( .A(n4996), .ZN(n4995) );
  INV_X1 U5636 ( .A(n9220), .ZN(n7315) );
  NAND2_X1 U5637 ( .A1(n9523), .A2(n9071), .ZN(n7348) );
  INV_X1 U5638 ( .A(n4541), .ZN(n6414) );
  OR2_X1 U5639 ( .A1(n9528), .A2(n8987), .ZN(n9278) );
  NAND2_X1 U5640 ( .A1(n6385), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6404) );
  INV_X1 U5641 ( .A(n6387), .ZN(n6385) );
  OR2_X1 U5642 ( .A1(n6375), .A2(n6374), .ZN(n6387) );
  NAND2_X1 U5643 ( .A1(n4542), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6375) );
  OR2_X1 U5644 ( .A1(n6349), .A2(n6346), .ZN(n7264) );
  NAND2_X1 U5645 ( .A1(n9118), .A2(n4543), .ZN(n7233) );
  NOR2_X1 U5646 ( .A1(n9580), .A2(n9587), .ZN(n4843) );
  OR2_X1 U5647 ( .A1(n8308), .A2(n8545), .ZN(n7225) );
  NAND2_X1 U5648 ( .A1(n7915), .A2(n7747), .ZN(n7194) );
  NAND2_X1 U5649 ( .A1(n8715), .A2(n7176), .ZN(n6495) );
  NOR2_X1 U5650 ( .A1(n9331), .A2(n4851), .ZN(n9287) );
  INV_X1 U5651 ( .A(n4853), .ZN(n4851) );
  NOR2_X1 U5652 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n5008) );
  NAND2_X1 U5653 ( .A1(n6117), .A2(n6769), .ZN(n6109) );
  OR2_X1 U5654 ( .A1(n6025), .A2(n6014), .ZN(n6048) );
  INV_X1 U5655 ( .A(n5484), .ZN(n4816) );
  NAND2_X1 U5656 ( .A1(n8747), .A2(n8746), .ZN(n8756) );
  NOR2_X1 U5657 ( .A1(n5658), .A2(n4812), .ZN(n4811) );
  NAND2_X1 U5658 ( .A1(n8780), .A2(n8779), .ZN(n9666) );
  NOR2_X1 U5659 ( .A1(n5446), .A2(n4802), .ZN(n5445) );
  NAND2_X1 U5660 ( .A1(n9852), .A2(n7150), .ZN(n5941) );
  NOR2_X1 U5661 ( .A1(n10277), .A2(n7452), .ZN(n4595) );
  OR2_X1 U5662 ( .A1(n4602), .A2(n4410), .ZN(n4601) );
  NAND2_X1 U5663 ( .A1(n4807), .A2(n9639), .ZN(n7048) );
  AND2_X1 U5664 ( .A1(n5938), .A2(n9849), .ZN(n7045) );
  NOR2_X1 U5665 ( .A1(n4815), .A2(n9745), .ZN(n4814) );
  NOR2_X1 U5666 ( .A1(n10129), .A2(n10134), .ZN(n5026) );
  INV_X1 U5667 ( .A(n4795), .ZN(n4790) );
  OR2_X1 U5668 ( .A1(n10134), .A2(n9930), .ZN(n7040) );
  INV_X1 U5669 ( .A(n7029), .ZN(n4839) );
  NAND2_X1 U5670 ( .A1(n9964), .A2(n9969), .ZN(n4587) );
  NOR2_X1 U5671 ( .A1(n4819), .A2(n5590), .ZN(n4818) );
  INV_X1 U5672 ( .A(n5591), .ZN(n5373) );
  INV_X1 U5673 ( .A(n5640), .ZN(n5374) );
  NAND2_X1 U5674 ( .A1(n7027), .A2(n4841), .ZN(n4840) );
  NOR2_X1 U5675 ( .A1(n7030), .A2(n4842), .ZN(n4841) );
  INV_X1 U5676 ( .A(n7026), .ZN(n4842) );
  NOR2_X1 U5677 ( .A1(n10196), .A2(n8641), .ZN(n5018) );
  OR2_X1 U5678 ( .A1(n8641), .A2(n8533), .ZN(n7019) );
  NAND2_X1 U5679 ( .A1(n4462), .A2(n7110), .ZN(n4800) );
  INV_X1 U5680 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7526) );
  INV_X1 U5681 ( .A(n8286), .ZN(n5490) );
  NAND2_X1 U5682 ( .A1(n8101), .A2(n7096), .ZN(n8053) );
  NAND2_X1 U5683 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5446) );
  INV_X1 U5684 ( .A(n5946), .ZN(n7720) );
  INV_X1 U5685 ( .A(n4785), .ZN(n4783) );
  AND2_X1 U5686 ( .A1(n10017), .A2(n4418), .ZN(n9950) );
  INV_X1 U5687 ( .A(n5009), .ZN(n7154) );
  NOR2_X1 U5688 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n4754) );
  AND2_X1 U5689 ( .A1(n5079), .A2(n5078), .ZN(n4755) );
  NAND2_X1 U5690 ( .A1(n5270), .A2(SI_14_), .ZN(n5271) );
  NAND2_X1 U5691 ( .A1(n5277), .A2(n5276), .ZN(n5589) );
  NAND2_X1 U5692 ( .A1(n5263), .A2(n5262), .ZN(n5545) );
  NAND2_X1 U5693 ( .A1(n5247), .A2(n5246), .ZN(n5250) );
  NAND2_X1 U5694 ( .A1(n5223), .A2(n5222), .ZN(n5453) );
  OAI21_X1 U5695 ( .B1(n5225), .B2(P2_DATAO_REG_3__SCAN_IN), .A(n4508), .ZN(
        n5214) );
  NAND2_X1 U5696 ( .A1(n5225), .A2(n7387), .ZN(n4508) );
  AND2_X1 U5697 ( .A1(n6712), .A2(n9088), .ZN(n6713) );
  NAND2_X1 U5698 ( .A1(n4541), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6428) );
  OR2_X1 U5699 ( .A1(n6428), .A2(n8969), .ZN(n6438) );
  OAI21_X1 U5700 ( .B1(n9035), .B2(n9114), .A(n9032), .ZN(n6703) );
  XNOR2_X1 U5701 ( .A(n9508), .B(n6719), .ZN(n9035) );
  NAND2_X1 U5702 ( .A1(n6254), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6272) );
  INV_X1 U5703 ( .A(n6270), .ZN(n6254) );
  NAND2_X1 U5704 ( .A1(n6295), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6317) );
  INV_X1 U5705 ( .A(n6297), .ZN(n6295) );
  OR2_X1 U5706 ( .A1(n6282), .A2(n8353), .ZN(n6297) );
  NAND2_X1 U5707 ( .A1(n6677), .A2(n4978), .ZN(n4977) );
  INV_X1 U5708 ( .A(n6678), .ZN(n4978) );
  AOI21_X1 U5709 ( .B1(n4407), .B2(n8372), .A(n4947), .ZN(n4946) );
  INV_X1 U5710 ( .A(n6669), .ZN(n4947) );
  AND2_X1 U5711 ( .A1(n7374), .A2(n7168), .ZN(n4987) );
  OAI21_X1 U5712 ( .B1(n4460), .B2(n4986), .A(n7372), .ZN(n4985) );
  INV_X1 U5713 ( .A(n7374), .ZN(n4986) );
  NOR2_X1 U5714 ( .A1(n7532), .A2(n6045), .ZN(n7600) );
  NAND2_X1 U5715 ( .A1(n4561), .A2(n6134), .ZN(n7604) );
  OR2_X1 U5716 ( .A1(n7535), .A2(n7536), .ZN(n4561) );
  OAI21_X1 U5717 ( .B1(n6210), .B2(P2_REG1_REG_4__SCAN_IN), .A(n4559), .ZN(
        n7602) );
  NAND2_X1 U5718 ( .A1(n6210), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4559) );
  NOR2_X1 U5719 ( .A1(n7600), .A2(n7599), .ZN(n7598) );
  AOI21_X1 U5720 ( .B1(n7604), .B2(n7603), .A(n7602), .ZN(n7606) );
  NOR2_X1 U5721 ( .A1(n7857), .A2(n6050), .ZN(n8045) );
  NOR2_X1 U5722 ( .A1(n8045), .A2(n8044), .ZN(n8043) );
  INV_X1 U5723 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8353) );
  AOI21_X1 U5724 ( .B1(n7411), .B2(P2_REG2_REG_9__SCAN_IN), .A(n8043), .ZN(
        n8359) );
  NOR2_X1 U5725 ( .A1(n8359), .A2(n8358), .ZN(n8357) );
  AOI21_X1 U5726 ( .B1(n4433), .B2(n4572), .A(n4421), .ZN(n4567) );
  AND2_X1 U5727 ( .A1(n8701), .A2(n8702), .ZN(n8723) );
  NAND2_X1 U5728 ( .A1(n9128), .A2(n4558), .ZN(n4557) );
  NAND2_X1 U5729 ( .A1(n9133), .A2(n6911), .ZN(n4558) );
  NAND2_X1 U5730 ( .A1(n4556), .A2(n4555), .ZN(n9158) );
  OR2_X1 U5731 ( .A1(n4557), .A2(n6073), .ZN(n4555) );
  NAND2_X1 U5732 ( .A1(n9138), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n4556) );
  XNOR2_X1 U5733 ( .A(n4741), .B(n4740), .ZN(n6148) );
  INV_X1 U5734 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n4740) );
  NAND2_X1 U5735 ( .A1(n4742), .A2(n4427), .ZN(n4741) );
  XNOR2_X1 U5736 ( .A(n4565), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n6150) );
  OR2_X1 U5737 ( .A1(n9181), .A2(n4566), .ZN(n4565) );
  NOR2_X1 U5738 ( .A1(n9192), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n4566) );
  AND2_X1 U5739 ( .A1(n8918), .A2(n6485), .ZN(n6740) );
  NAND2_X1 U5740 ( .A1(n9234), .A2(n4857), .ZN(n8916) );
  NOR2_X1 U5741 ( .A1(n4860), .A2(n4858), .ZN(n4857) );
  OR2_X1 U5742 ( .A1(n9488), .A2(n9237), .ZN(n4858) );
  OAI21_X1 U5743 ( .B1(n9229), .B2(n4995), .A(n4993), .ZN(n4554) );
  NOR2_X1 U5744 ( .A1(n5000), .A2(n6552), .ZN(n4999) );
  NAND2_X1 U5745 ( .A1(n9266), .A2(n4853), .ZN(n4852) );
  INV_X1 U5746 ( .A(n4907), .ZN(n4906) );
  INV_X1 U5747 ( .A(n4910), .ZN(n4909) );
  NOR2_X1 U5748 ( .A1(n7351), .A2(n9311), .ZN(n9340) );
  NAND2_X1 U5749 ( .A1(n4545), .A2(n4414), .ZN(n9345) );
  NOR2_X1 U5750 ( .A1(n9390), .A2(n9545), .ZN(n9361) );
  INV_X1 U5751 ( .A(n4542), .ZN(n6365) );
  INV_X1 U5752 ( .A(n6330), .ZN(n6329) );
  OR2_X1 U5753 ( .A1(n9388), .A2(n9392), .ZN(n9390) );
  NAND2_X1 U5754 ( .A1(n7257), .A2(n7258), .ZN(n8680) );
  NAND2_X1 U5755 ( .A1(n9415), .A2(n4998), .ZN(n8669) );
  AND2_X1 U5756 ( .A1(n6544), .A2(n7253), .ZN(n4998) );
  AND2_X1 U5757 ( .A1(n7243), .A2(n7253), .ZN(n9424) );
  INV_X1 U5758 ( .A(n8660), .ZN(n6572) );
  AND2_X1 U5759 ( .A1(n6569), .A2(n4843), .ZN(n8229) );
  INV_X1 U5760 ( .A(n9117), .ZN(n8655) );
  AND3_X1 U5761 ( .A1(n4847), .A2(n6568), .A3(n4844), .ZN(n8306) );
  AND2_X1 U5762 ( .A1(n4845), .A2(n8196), .ZN(n4844) );
  AND2_X1 U5763 ( .A1(n7225), .A2(n8541), .ZN(n8299) );
  NAND2_X1 U5764 ( .A1(n4846), .A2(n4847), .ZN(n8176) );
  INV_X1 U5765 ( .A(n7748), .ZN(n4846) );
  OR2_X1 U5766 ( .A1(n6532), .A2(n6531), .ZN(n6533) );
  OAI21_X1 U5767 ( .B1(n7839), .B2(n7836), .A(n6201), .ZN(n7776) );
  NAND2_X1 U5768 ( .A1(n7846), .A2(n7847), .ZN(n7845) );
  AND2_X1 U5769 ( .A1(n6586), .A2(n10463), .ZN(n7846) );
  NAND2_X1 U5770 ( .A1(n6745), .A2(n6744), .ZN(n9483) );
  NAND2_X1 U5771 ( .A1(n6328), .A2(n6327), .ZN(n6337) );
  INV_X1 U5772 ( .A(n10508), .ZN(n9589) );
  INV_X1 U5773 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5007) );
  OR2_X1 U5774 ( .A1(n6109), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n6111) );
  AND2_X1 U5775 ( .A1(n4983), .A2(n6084), .ZN(n4982) );
  NOR2_X1 U5776 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n4983) );
  INV_X1 U5777 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4981) );
  XNOR2_X1 U5778 ( .A(n6034), .B(P2_IR_REG_2__SCAN_IN), .ZN(n6175) );
  OR2_X1 U5779 ( .A1(n5516), .A2(n7526), .ZN(n5575) );
  NAND2_X1 U5780 ( .A1(n4816), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U5781 ( .A1(n8824), .A2(n9741), .ZN(n9655) );
  NAND2_X1 U5782 ( .A1(n5373), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5606) );
  NOR2_X1 U5783 ( .A1(n8762), .A2(n4869), .ZN(n4866) );
  NAND2_X1 U5784 ( .A1(n8280), .A2(n8279), .ZN(n8281) );
  NAND2_X1 U5785 ( .A1(n10427), .A2(n8785), .ZN(n8280) );
  OR2_X1 U5786 ( .A1(n8386), .A2(n4401), .ZN(n8279) );
  NAND2_X1 U5787 ( .A1(n8400), .A2(n8401), .ZN(n8521) );
  NAND2_X1 U5788 ( .A1(n5374), .A2(n4811), .ZN(n5694) );
  NAND2_X1 U5789 ( .A1(n4810), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5550) );
  INV_X1 U5790 ( .A(n5560), .ZN(n4810) );
  NAND2_X1 U5791 ( .A1(n4461), .A2(n8434), .ZN(n8446) );
  NAND2_X1 U5792 ( .A1(n5372), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5577) );
  INV_X1 U5793 ( .A(n5575), .ZN(n5372) );
  OR2_X1 U5794 ( .A1(n5577), .A2(n7658), .ZN(n5560) );
  INV_X1 U5795 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7658) );
  NAND2_X1 U5796 ( .A1(n5445), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5484) );
  AOI21_X1 U5797 ( .B1(n4678), .B2(n7089), .A(n5947), .ZN(n4677) );
  OAI21_X1 U5798 ( .B1(n5996), .B2(n9837), .A(n10083), .ZN(n5948) );
  AND2_X1 U5799 ( .A1(n6000), .A2(n5999), .ZN(n6004) );
  AND2_X1 U5800 ( .A1(n5647), .A2(n5646), .ZN(n8789) );
  AND2_X1 U5801 ( .A1(n7437), .A2(n4469), .ZN(n7438) );
  NOR2_X1 U5802 ( .A1(n10306), .A2(n5027), .ZN(n10278) );
  NOR2_X1 U5803 ( .A1(n10276), .A2(n4601), .ZN(n7692) );
  AND2_X1 U5804 ( .A1(n9818), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5165) );
  NOR2_X1 U5805 ( .A1(n9815), .A2(n9814), .ZN(n9813) );
  NAND2_X1 U5806 ( .A1(n7489), .A2(n4437), .ZN(n7523) );
  NAND2_X1 U5807 ( .A1(n4591), .A2(n4590), .ZN(n5171) );
  OR2_X1 U5808 ( .A1(n8140), .A2(n6829), .ZN(n4590) );
  NAND2_X1 U5809 ( .A1(n4593), .A2(n4592), .ZN(n4591) );
  INV_X1 U5810 ( .A(n8137), .ZN(n4592) );
  OR2_X1 U5811 ( .A1(n9824), .A2(n9825), .ZN(n4628) );
  NAND2_X1 U5812 ( .A1(n9859), .A2(n4445), .ZN(n5020) );
  NOR2_X1 U5813 ( .A1(n10093), .A2(n10107), .ZN(n5019) );
  NAND2_X1 U5814 ( .A1(n8938), .A2(n8945), .ZN(n8939) );
  INV_X1 U5815 ( .A(n8935), .ZN(n8948) );
  NOR2_X1 U5816 ( .A1(n7149), .A2(n4786), .ZN(n4785) );
  INV_X1 U5817 ( .A(n7147), .ZN(n4786) );
  NAND2_X1 U5818 ( .A1(n4787), .A2(n4782), .ZN(n4779) );
  AND2_X1 U5819 ( .A1(n5827), .A2(n5826), .ZN(n9634) );
  OR2_X1 U5820 ( .A1(n8942), .A2(n5821), .ZN(n5827) );
  XNOR2_X1 U5821 ( .A(n5818), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9637) );
  NAND2_X1 U5822 ( .A1(n5376), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5818) );
  INV_X1 U5823 ( .A(n5778), .ZN(n5376) );
  INV_X1 U5824 ( .A(n9791), .ZN(n9872) );
  XNOR2_X1 U5825 ( .A(n9870), .B(n4837), .ZN(n4836) );
  INV_X1 U5826 ( .A(n9869), .ZN(n4837) );
  AND2_X1 U5827 ( .A1(n9885), .A2(n9886), .ZN(n4586) );
  NAND2_X1 U5828 ( .A1(n9931), .A2(n5026), .ZN(n9895) );
  AND2_X1 U5829 ( .A1(n7040), .A2(n7041), .ZN(n9917) );
  AND2_X1 U5830 ( .A1(n5718), .A2(n5717), .ZN(n9948) );
  NAND2_X1 U5831 ( .A1(n4587), .A2(n5931), .ZN(n9944) );
  OR2_X1 U5832 ( .A1(n7032), .A2(n7033), .ZN(n9964) );
  INV_X1 U5833 ( .A(n4587), .ZN(n9965) );
  NAND2_X1 U5834 ( .A1(n10017), .A2(n5023), .ZN(n9986) );
  NAND2_X1 U5835 ( .A1(n10017), .A2(n4408), .ZN(n9958) );
  AND2_X1 U5836 ( .A1(n5896), .A2(n5931), .ZN(n9969) );
  NAND2_X1 U5837 ( .A1(n5373), .A2(n4817), .ZN(n5640) );
  AND2_X1 U5838 ( .A1(n4818), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n4817) );
  NAND2_X1 U5839 ( .A1(n5374), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5659) );
  NAND2_X1 U5840 ( .A1(n4840), .A2(n7029), .ZN(n10002) );
  AND2_X1 U5841 ( .A1(n5904), .A2(n9978), .ZN(n10001) );
  NOR2_X1 U5842 ( .A1(n7123), .A2(n10026), .ZN(n4510) );
  NAND2_X1 U5843 ( .A1(n4809), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5540) );
  INV_X1 U5844 ( .A(n5550), .ZN(n4809) );
  NAND2_X1 U5845 ( .A1(n4808), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5591) );
  INV_X1 U5846 ( .A(n5540), .ZN(n4808) );
  NAND2_X1 U5847 ( .A1(n8624), .A2(n7022), .ZN(n10066) );
  NAND2_X1 U5848 ( .A1(n5538), .A2(n5537), .ZN(n10061) );
  AND2_X1 U5849 ( .A1(n8631), .A2(n10186), .ZN(n10057) );
  NAND2_X1 U5850 ( .A1(n8506), .A2(n5018), .ZN(n8632) );
  NAND2_X1 U5851 ( .A1(n8506), .A2(n8507), .ZN(n8565) );
  NAND2_X1 U5852 ( .A1(n5015), .A2(n5013), .ZN(n8323) );
  NOR2_X1 U5853 ( .A1(n5014), .A2(n8246), .ZN(n5013) );
  NAND2_X1 U5854 ( .A1(n5015), .A2(n5012), .ZN(n8259) );
  NOR2_X1 U5855 ( .A1(n8246), .A2(n8260), .ZN(n5012) );
  NAND2_X1 U5856 ( .A1(n4828), .A2(n7101), .ZN(n8318) );
  NOR2_X1 U5857 ( .A1(n5016), .A2(n8246), .ZN(n8257) );
  OAI21_X1 U5858 ( .B1(n5524), .B2(n4676), .A(n4675), .ZN(n4674) );
  INV_X1 U5859 ( .A(n10068), .ZN(n10040) );
  INV_X1 U5860 ( .A(n10011), .ZN(n10071) );
  AND2_X1 U5861 ( .A1(n7055), .A2(n7684), .ZN(n10068) );
  AND2_X1 U5862 ( .A1(n7089), .A2(n7993), .ZN(n10184) );
  INV_X1 U5863 ( .A(n10413), .ZN(n10429) );
  OR2_X1 U5864 ( .A1(n5407), .A2(n5010), .ZN(n5401) );
  NAND2_X1 U5865 ( .A1(n7087), .A2(n7086), .ZN(n7975) );
  XNOR2_X1 U5866 ( .A(n5843), .B(n5842), .ZN(n9617) );
  OAI21_X1 U5867 ( .B1(n5840), .B2(n5839), .A(n5838), .ZN(n5843) );
  XNOR2_X1 U5868 ( .A(n5840), .B(SI_30_), .ZN(n8953) );
  XNOR2_X1 U5869 ( .A(n5834), .B(n5833), .ZN(n9623) );
  AND2_X1 U5870 ( .A1(n5340), .A2(n5796), .ZN(n5814) );
  NAND2_X1 U5871 ( .A1(n4661), .A2(n4666), .ZN(n5795) );
  AND2_X1 U5872 ( .A1(n5386), .A2(n5344), .ZN(n5813) );
  CLKBUF_X1 U5873 ( .A(n5159), .Z(n7684) );
  XNOR2_X1 U5874 ( .A(n5799), .B(n5798), .ZN(n8691) );
  NAND2_X1 U5875 ( .A1(n4658), .A2(n4662), .ZN(n5799) );
  AOI21_X1 U5876 ( .B1(n4666), .B2(n4664), .A(n4663), .ZN(n4662) );
  NAND2_X1 U5877 ( .A1(n5144), .A2(n5056), .ZN(n7065) );
  XNOR2_X1 U5878 ( .A(n5745), .B(n5744), .ZN(n8477) );
  INV_X1 U5879 ( .A(n4648), .ZN(n5721) );
  AOI21_X1 U5880 ( .B1(n5304), .B2(n4654), .A(n4649), .ZN(n4648) );
  INV_X1 U5881 ( .A(n5307), .ZN(n4649) );
  INV_X1 U5882 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5954) );
  XNOR2_X1 U5883 ( .A(n5654), .B(n5653), .ZN(n7883) );
  XNOR2_X1 U5884 ( .A(n5636), .B(n5635), .ZN(n7879) );
  AOI21_X1 U5885 ( .B1(n5650), .B2(n5634), .A(n5633), .ZN(n5636) );
  XNOR2_X1 U5886 ( .A(n5619), .B(n5618), .ZN(n7832) );
  NAND2_X1 U5887 ( .A1(n4927), .A2(n4930), .ZN(n5617) );
  AOI21_X1 U5888 ( .B1(n4934), .B2(n4932), .A(n4931), .ZN(n4930) );
  AND2_X1 U5889 ( .A1(n5107), .A2(n5106), .ZN(n5525) );
  NAND2_X1 U5890 ( .A1(n4921), .A2(n4922), .ZN(n5556) );
  OR2_X1 U5891 ( .A1(n5251), .A2(n4925), .ZN(n4921) );
  AND2_X2 U5892 ( .A1(n5051), .A2(n5050), .ZN(n4672) );
  NAND2_X1 U5893 ( .A1(n5502), .A2(n5501), .ZN(n4521) );
  XNOR2_X1 U5894 ( .A(n5500), .B(n5498), .ZN(n6236) );
  XNOR2_X1 U5895 ( .A(n5214), .B(SI_3_), .ZN(n5429) );
  XNOR2_X1 U5896 ( .A(n5122), .B(P1_IR_REG_2__SCAN_IN), .ZN(n7399) );
  NOR2_X1 U5897 ( .A1(n10559), .A2(n10254), .ZN(n10255) );
  NOR2_X1 U5898 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10558), .ZN(n10254) );
  NAND2_X1 U5899 ( .A1(n4948), .A2(n4407), .ZN(n8607) );
  AND2_X1 U5900 ( .A1(n4948), .A2(n4432), .ZN(n8608) );
  NAND2_X1 U5901 ( .A1(n4949), .A2(n6663), .ZN(n4948) );
  AND3_X1 U5902 ( .A1(n6169), .A2(n4615), .A3(n4614), .ZN(n7922) );
  NAND2_X1 U5903 ( .A1(n4423), .A2(n4616), .ZN(n4615) );
  NAND2_X1 U5904 ( .A1(n6382), .A2(n7537), .ZN(n4614) );
  NAND2_X1 U5905 ( .A1(n8976), .A2(n8975), .ZN(n8974) );
  NAND2_X1 U5906 ( .A1(n4970), .A2(n4968), .ZN(n8976) );
  NAND2_X1 U5907 ( .A1(n4511), .A2(n4971), .ZN(n4970) );
  NOR2_X1 U5908 ( .A1(n6732), .A2(n4954), .ZN(n4951) );
  NOR2_X1 U5909 ( .A1(n4956), .A2(n4953), .ZN(n4952) );
  NOR3_X1 U5910 ( .A1(n4954), .A2(n6732), .A3(n8962), .ZN(n4953) );
  NAND2_X1 U5911 ( .A1(n4957), .A2(n6731), .ZN(n4956) );
  INV_X1 U5912 ( .A(n4958), .ZN(n4955) );
  AND2_X1 U5914 ( .A1(n8615), .A2(n9446), .ZN(n9103) );
  INV_X1 U5915 ( .A(n4966), .ZN(n4965) );
  OAI21_X1 U5916 ( .B1(n4968), .B2(n4967), .A(n6685), .ZN(n4966) );
  AND2_X1 U5917 ( .A1(n6734), .A2(n6733), .ZN(n8615) );
  INV_X1 U5918 ( .A(n9110), .ZN(n9048) );
  NAND2_X1 U5919 ( .A1(n4973), .A2(n4977), .ZN(n9078) );
  OR2_X1 U5920 ( .A1(n4511), .A2(n9024), .ZN(n4973) );
  NAND2_X1 U5921 ( .A1(n4533), .A2(n9085), .ZN(n9086) );
  NAND2_X1 U5922 ( .A1(n9084), .A2(n9087), .ZN(n4533) );
  OR2_X1 U5923 ( .A1(n6349), .A2(n6348), .ZN(n9556) );
  OR2_X1 U5924 ( .A1(n9224), .A2(n6561), .ZN(n6467) );
  NAND4_X1 U5925 ( .A1(n6263), .A2(n6262), .A3(n6261), .A4(n6260), .ZN(n9119)
         );
  NAND4_X1 U5926 ( .A1(n6247), .A2(n6246), .A3(n6245), .A4(n6244), .ZN(n9121)
         );
  AOI21_X1 U5927 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n6175), .A(n7571), .ZN(
        n7534) );
  NOR2_X1 U5928 ( .A1(n7534), .A2(n7533), .ZN(n7532) );
  AND2_X1 U5929 ( .A1(n6032), .A2(n6031), .ZN(n7596) );
  NAND2_X1 U5930 ( .A1(n4573), .A2(n4576), .ZN(n8038) );
  NAND2_X1 U5931 ( .A1(n4570), .A2(n4571), .ZN(n8351) );
  NOR2_X1 U5932 ( .A1(n8357), .A2(n6056), .ZN(n8482) );
  AND2_X1 U5933 ( .A1(n6280), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6056) );
  NAND2_X1 U5934 ( .A1(n4750), .A2(n4749), .ZN(n8719) );
  AOI21_X1 U5935 ( .B1(n4749), .B2(n8709), .A(n4484), .ZN(n4748) );
  XNOR2_X1 U5936 ( .A(n4557), .B(n9146), .ZN(n9138) );
  AND3_X1 U5937 ( .A1(n9139), .A2(n4745), .A3(n6075), .ZN(n9150) );
  NOR2_X1 U5938 ( .A1(n4746), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4744) );
  NAND2_X1 U5939 ( .A1(n9168), .A2(n4490), .ZN(n9183) );
  OAI21_X1 U5940 ( .B1(n9213), .B2(n4992), .A(n4916), .ZN(n6497) );
  AOI21_X1 U5941 ( .B1(n6567), .B2(n10460), .A(n6566), .ZN(n9490) );
  NAND2_X1 U5942 ( .A1(n6565), .A2(n6564), .ZN(n6566) );
  NAND2_X1 U5943 ( .A1(n9113), .A2(n9444), .ZN(n6565) );
  AOI21_X1 U5944 ( .B1(n9492), .B2(n9472), .A(n9212), .ZN(n4624) );
  NAND2_X1 U5945 ( .A1(n4997), .A2(n4996), .ZN(n9217) );
  OAI21_X1 U5946 ( .B1(n9259), .B2(n4902), .A(n4903), .ZN(n9233) );
  INV_X1 U5947 ( .A(n9508), .ZN(n9248) );
  NAND2_X1 U5948 ( .A1(n9258), .A2(n5037), .ZN(n9243) );
  NAND2_X1 U5949 ( .A1(n9280), .A2(n7293), .ZN(n9260) );
  INV_X1 U5950 ( .A(n9523), .ZN(n6573) );
  AND2_X1 U5951 ( .A1(n4911), .A2(n4431), .ZN(n9322) );
  NAND2_X1 U5952 ( .A1(n9368), .A2(n6371), .ZN(n9353) );
  OAI21_X1 U5953 ( .B1(n9399), .B2(n7269), .A(n4549), .ZN(n9358) );
  NAND2_X1 U5954 ( .A1(n4423), .A2(n7393), .ZN(n4726) );
  OR2_X1 U5955 ( .A1(n10472), .A2(n6756), .ZN(n9290) );
  OR2_X1 U5956 ( .A1(n10461), .A2(n6578), .ZN(n10464) );
  INV_X1 U5957 ( .A(n9290), .ZN(n10462) );
  OAI211_X1 U5958 ( .C1(n8903), .C2(n10508), .A(n9480), .B(n6755), .ZN(n9482)
         );
  AND2_X2 U5959 ( .A1(n7676), .A2(n7675), .ZN(n10526) );
  INV_X1 U5960 ( .A(n9211), .ZN(n9496) );
  AND2_X1 U5961 ( .A1(n6737), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10487) );
  INV_X1 U5962 ( .A(n10481), .ZN(n10484) );
  INV_X1 U5963 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n6160) );
  INV_X1 U5964 ( .A(n6163), .ZN(n9626) );
  XNOR2_X1 U5965 ( .A(n6088), .B(P2_IR_REG_24__SCAN_IN), .ZN(n8493) );
  NAND2_X1 U5966 ( .A1(n6111), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6088) );
  INV_X1 U5967 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7886) );
  INV_X1 U5968 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7680) );
  INV_X1 U5969 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7513) );
  INV_X1 U5970 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7477) );
  INV_X1 U5971 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7430) );
  INV_X1 U5972 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7420) );
  INV_X1 U5973 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7412) );
  NAND2_X1 U5974 ( .A1(n6036), .A2(n6039), .ZN(n7568) );
  MUX2_X1 U5975 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6035), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n6036) );
  NAND2_X1 U5976 ( .A1(n8024), .A2(n8338), .ZN(n8278) );
  NAND2_X1 U5977 ( .A1(n4876), .A2(n4878), .ZN(n4875) );
  NAND2_X1 U5978 ( .A1(n8809), .A2(n9730), .ZN(n9680) );
  AND2_X1 U5979 ( .A1(n8797), .A2(n8804), .ZN(n4882) );
  NAND2_X1 U5980 ( .A1(n5709), .A2(n5708), .ZN(n10141) );
  AND3_X1 U5981 ( .A1(n5610), .A2(n5609), .A3(n5608), .ZN(n10041) );
  NAND2_X1 U5982 ( .A1(n4883), .A2(n8797), .ZN(n9734) );
  NAND2_X1 U5983 ( .A1(n4873), .A2(n8587), .ZN(n8597) );
  NAND2_X1 U5984 ( .A1(n7822), .A2(n7821), .ZN(n9778) );
  AND2_X1 U5985 ( .A1(n7817), .A2(n7615), .ZN(n8347) );
  INV_X1 U5986 ( .A(n10116), .ZN(n9858) );
  INV_X1 U5987 ( .A(n9683), .ZN(n9780) );
  NAND2_X1 U5988 ( .A1(n4867), .A2(n8763), .ZN(n9777) );
  AND2_X1 U5989 ( .A1(n8347), .A2(n10428), .ZN(n9784) );
  INV_X1 U5990 ( .A(n9888), .ZN(n9792) );
  NAND2_X1 U5991 ( .A1(n5754), .A2(n5753), .ZN(n9905) );
  OR2_X1 U5992 ( .A1(n9889), .A2(n5821), .ZN(n5754) );
  NAND2_X1 U5993 ( .A1(n5741), .A2(n5740), .ZN(n9919) );
  OR2_X1 U5994 ( .A1(n9897), .A2(n5821), .ZN(n5741) );
  NAND2_X1 U5995 ( .A1(n5730), .A2(n5729), .ZN(n9903) );
  OR2_X1 U5996 ( .A1(n9913), .A2(n5821), .ZN(n5730) );
  INV_X1 U5997 ( .A(n10041), .ZN(n5611) );
  NOR2_X1 U5998 ( .A1(n9813), .A2(n4609), .ZN(n7485) );
  AOI21_X1 U5999 ( .B1(n4605), .B2(n4609), .A(n4604), .ZN(n4603) );
  INV_X1 U6000 ( .A(n7471), .ZN(n4604) );
  AOI21_X1 U6001 ( .B1(n7516), .B2(n7500), .A(n7499), .ZN(n7511) );
  OR2_X1 U6002 ( .A1(n7519), .A2(n7518), .ZN(n7516) );
  NAND2_X1 U6003 ( .A1(n7650), .A2(n5029), .ZN(n7889) );
  NAND2_X1 U6004 ( .A1(n4633), .A2(n4635), .ZN(n7894) );
  OAI21_X1 U6005 ( .B1(n7655), .B2(n4632), .A(n4629), .ZN(n4639) );
  AOI21_X1 U6006 ( .B1(n4631), .B2(n4630), .A(n8135), .ZN(n4629) );
  INV_X1 U6007 ( .A(n4634), .ZN(n4630) );
  INV_X1 U6008 ( .A(n4593), .ZN(n8136) );
  XNOR2_X1 U6009 ( .A(n5171), .B(n5525), .ZN(n8424) );
  NAND2_X1 U6010 ( .A1(n10318), .A2(n5157), .ZN(n10331) );
  OAI21_X1 U6011 ( .B1(n10326), .B2(n5176), .A(n10332), .ZN(n10350) );
  INV_X1 U6012 ( .A(n4628), .ZN(n9823) );
  NAND2_X1 U6013 ( .A1(n5188), .A2(n10344), .ZN(n5189) );
  INV_X1 U6014 ( .A(n10087), .ZN(n9843) );
  AND2_X1 U6015 ( .A1(n5021), .A2(n5020), .ZN(n10098) );
  AOI21_X1 U6016 ( .B1(n8939), .B2(n10093), .A(n10413), .ZN(n5021) );
  NAND2_X1 U6017 ( .A1(n4788), .A2(n7147), .ZN(n8889) );
  OR2_X1 U6018 ( .A1(n9855), .A2(n7148), .ZN(n4788) );
  AND2_X1 U6019 ( .A1(n5778), .A2(n5761), .ZN(n9874) );
  NAND2_X1 U6020 ( .A1(n4585), .A2(n4583), .ZN(n10125) );
  INV_X1 U6021 ( .A(n4584), .ZN(n4583) );
  OAI21_X1 U6022 ( .B1(n9884), .B2(n4586), .A(n10074), .ZN(n4585) );
  OAI22_X1 U6023 ( .A1(n9888), .A2(n10040), .B1(n10071), .B2(n9887), .ZN(n4584) );
  NAND2_X1 U6024 ( .A1(n4763), .A2(n4764), .ZN(n9880) );
  OR2_X1 U6025 ( .A1(n7142), .A2(n4766), .ZN(n4763) );
  NAND2_X1 U6026 ( .A1(n4794), .A2(n4792), .ZN(n9937) );
  NAND2_X1 U6027 ( .A1(n7136), .A2(n4795), .ZN(n4794) );
  NAND2_X1 U6028 ( .A1(n7136), .A2(n7135), .ZN(n9942) );
  NAND2_X1 U6029 ( .A1(n4771), .A2(n7117), .ZN(n10055) );
  OR2_X1 U6030 ( .A1(n8619), .A2(n7118), .ZN(n4771) );
  NAND2_X1 U6031 ( .A1(n8314), .A2(n7109), .ZN(n8378) );
  NAND2_X1 U6032 ( .A1(n5620), .A2(n10239), .ZN(n5412) );
  INV_X1 U6033 ( .A(n9999), .ZN(n10060) );
  OAI21_X1 U6034 ( .B1(n10124), .B2(n10102), .A(n4415), .ZN(n4831) );
  AND2_X1 U6035 ( .A1(n10123), .A2(n10428), .ZN(n4832) );
  OAI211_X1 U6036 ( .C1(n10128), .C2(n10102), .A(n4582), .B(n4580), .ZN(n10208) );
  NOR2_X1 U6037 ( .A1(n10126), .A2(n4581), .ZN(n4580) );
  INV_X1 U6038 ( .A(n10125), .ZN(n4582) );
  AND2_X1 U6039 ( .A1(n10127), .A2(n10428), .ZN(n4581) );
  NOR2_X1 U6040 ( .A1(n10355), .A2(n10354), .ZN(n10367) );
  AND2_X1 U6041 ( .A1(n7812), .A2(n5952), .ZN(n10225) );
  INV_X1 U6042 ( .A(n7975), .ZN(n10226) );
  INV_X1 U6043 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n4776) );
  XNOR2_X1 U6044 ( .A(n5814), .B(n5813), .ZN(n8715) );
  OAI21_X1 U6045 ( .B1(n5304), .B2(n4652), .A(n4650), .ZN(n5732) );
  INV_X1 U6046 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7884) );
  INV_X1 U6047 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7835) );
  INV_X1 U6048 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7515) );
  INV_X1 U6049 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7498) );
  INV_X1 U6050 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7480) );
  INV_X1 U6051 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n7436) );
  INV_X1 U6052 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n7415) );
  INV_X1 U6053 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n7422) );
  NOR2_X1 U6054 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10265), .ZN(n10563) );
  NOR2_X1 U6055 ( .A1(n10564), .A2(n10562), .ZN(n10555) );
  NOR2_X1 U6056 ( .A1(n10555), .A2(n10554), .ZN(n10553) );
  AOI21_X1 U6057 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10553), .ZN(n10552) );
  NOR2_X1 U6058 ( .A1(n10552), .A2(n10551), .ZN(n10550) );
  AOI21_X1 U6059 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10550), .ZN(n10549) );
  OAI21_X1 U6060 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10547), .ZN(n10545) );
  INV_X1 U6061 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n10270) );
  NAND2_X1 U6062 ( .A1(n4980), .A2(n6616), .ZN(n7912) );
  NAND2_X1 U6063 ( .A1(n4731), .A2(n8273), .ZN(n4507) );
  AOI21_X1 U6064 ( .B1(n6147), .B2(n4944), .A(n6146), .ZN(n6155) );
  OR2_X1 U6065 ( .A1(n6153), .A2(n4944), .ZN(n6154) );
  NAND2_X1 U6066 ( .A1(n4623), .A2(n4622), .ZN(P2_U3269) );
  NAND2_X1 U6067 ( .A1(n9211), .A2(n10467), .ZN(n4622) );
  AND2_X1 U6068 ( .A1(n4625), .A2(n4624), .ZN(n4623) );
  OR2_X1 U6069 ( .A1(n9495), .A2(n10461), .ZN(n4625) );
  OR2_X1 U6070 ( .A1(n10526), .A2(n4849), .ZN(n4848) );
  NAND2_X1 U6071 ( .A1(n9596), .A2(n10526), .ZN(n4850) );
  INV_X1 U6072 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n4849) );
  OR2_X1 U6073 ( .A1(n10516), .A2(n4669), .ZN(n4668) );
  NAND2_X1 U6074 ( .A1(n9596), .A2(n10516), .ZN(n4670) );
  INV_X1 U6075 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n4669) );
  OAI21_X1 U6076 ( .B1(n4417), .B2(n4406), .A(n4892), .ZN(n4887) );
  OR2_X1 U6077 ( .A1(n4894), .A2(n4891), .ZN(n4890) );
  INV_X1 U6078 ( .A(n4515), .ZN(n8952) );
  OAI21_X1 U6079 ( .B1(n10110), .B2(n10020), .A(n4516), .ZN(n4515) );
  AOI21_X1 U6080 ( .B1(n10108), .B2(n10007), .A(n8951), .ZN(n4516) );
  NOR2_X1 U6081 ( .A1(n10132), .A2(n10020), .ZN(n9906) );
  AND4_X1 U6082 ( .A1(n4755), .A2(n5080), .A3(n4754), .A4(n4758), .ZN(n4403)
         );
  NAND2_X1 U6083 ( .A1(n9535), .A2(n9346), .ZN(n4404) );
  NOR2_X1 U6084 ( .A1(n7150), .A2(n4807), .ZN(n4405) );
  AND2_X1 U6085 ( .A1(n4896), .A2(n4899), .ZN(n4406) );
  AND2_X1 U6086 ( .A1(n8609), .A2(n4432), .ZN(n4407) );
  AOI21_X1 U6087 ( .B1(n9637), .B2(n4402), .A(n5806), .ZN(n9852) );
  INV_X1 U6088 ( .A(n9852), .ZN(n4807) );
  INV_X1 U6089 ( .A(n6527), .ZN(n7752) );
  AND2_X1 U6090 ( .A1(n5023), .A2(n9962), .ZN(n4408) );
  INV_X1 U6091 ( .A(n8196), .ZN(n7747) );
  AOI21_X1 U6092 ( .B1(n8962), .B2(n4961), .A(n6718), .ZN(n4960) );
  INV_X1 U6093 ( .A(n4960), .ZN(n4954) );
  AND2_X1 U6094 ( .A1(n7390), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4410) );
  NOR2_X1 U6095 ( .A1(n4700), .A2(n5854), .ZN(n4699) );
  NOR2_X1 U6096 ( .A1(n9199), .A2(n7431), .ZN(n7325) );
  AND2_X1 U6097 ( .A1(n9484), .A2(n9589), .ZN(n4411) );
  OR2_X1 U6098 ( .A1(n9545), .A2(n6370), .ZN(n7274) );
  AND2_X1 U6099 ( .A1(n4868), .A2(n8758), .ZN(n4412) );
  AND2_X1 U6100 ( .A1(n7273), .A2(n7272), .ZN(n4413) );
  OR2_X1 U6101 ( .A1(n4547), .A2(n6545), .ZN(n4414) );
  NOR2_X1 U6102 ( .A1(n10122), .A2(n4832), .ZN(n4415) );
  AND2_X1 U6103 ( .A1(n5026), .A2(n5025), .ZN(n4416) );
  NAND2_X1 U6104 ( .A1(n4893), .A2(n4897), .ZN(n4417) );
  NAND2_X1 U6105 ( .A1(n7295), .A2(n7294), .ZN(n9261) );
  INV_X1 U6106 ( .A(n9261), .ZN(n4716) );
  AND2_X1 U6107 ( .A1(n4408), .A2(n5022), .ZN(n4418) );
  AND2_X1 U6108 ( .A1(n5018), .A2(n5017), .ZN(n4419) );
  NAND2_X1 U6109 ( .A1(n9528), .A2(n9328), .ZN(n4420) );
  AND2_X1 U6110 ( .A1(n6057), .A2(n6055), .ZN(n6280) );
  AND2_X1 U6111 ( .A1(n6280), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4421) );
  NAND2_X2 U6112 ( .A1(n6235), .A2(n6234), .ZN(n8180) );
  INV_X1 U6113 ( .A(n8180), .ZN(n4847) );
  OAI211_X2 U6114 ( .C1(n5524), .C2(n7398), .A(n5402), .B(n5401), .ZN(n7153)
         );
  NAND2_X1 U6115 ( .A1(n4770), .A2(n4769), .ZN(n8733) );
  AND2_X2 U6116 ( .A1(n6197), .A2(n7388), .ZN(n4423) );
  INV_X1 U6117 ( .A(n9209), .ZN(n4992) );
  AND2_X1 U6118 ( .A1(n9361), .A2(n9351), .ZN(n9330) );
  AND2_X1 U6119 ( .A1(n7028), .A2(n7029), .ZN(n7123) );
  NAND2_X1 U6120 ( .A1(n4911), .A2(n4909), .ZN(n9323) );
  INV_X1 U6121 ( .A(n5430), .ZN(n5535) );
  AND2_X1 U6122 ( .A1(n9931), .A2(n4416), .ZN(n4424) );
  AND2_X1 U6123 ( .A1(n8264), .A2(n4684), .ZN(n4425) );
  AND2_X1 U6124 ( .A1(n5975), .A2(n7096), .ZN(n4426) );
  OR2_X1 U6125 ( .A1(n6083), .A2(n6082), .ZN(n4427) );
  NAND2_X1 U6126 ( .A1(n5358), .A2(n5357), .ZN(n10087) );
  INV_X1 U6127 ( .A(n4902), .ZN(n4904) );
  OR2_X1 U6128 ( .A1(n4905), .A2(n9250), .ZN(n4902) );
  XNOR2_X1 U6129 ( .A(n8281), .B(n8872), .ZN(n8525) );
  INV_X1 U6130 ( .A(n4405), .ZN(n4787) );
  AND3_X1 U6131 ( .A1(n4861), .A2(n7869), .A3(n8930), .ZN(n4428) );
  AND3_X1 U6132 ( .A1(n4689), .A2(n4687), .A3(n4698), .ZN(n4429) );
  NOR2_X1 U6133 ( .A1(n9508), .A2(n9114), .ZN(n4430) );
  OR2_X1 U6134 ( .A1(n9535), .A2(n9346), .ZN(n4431) );
  NAND2_X1 U6135 ( .A1(n6662), .A2(n6661), .ZN(n4432) );
  AND2_X1 U6136 ( .A1(n4571), .A2(n4569), .ZN(n4433) );
  INV_X1 U6137 ( .A(n7041), .ZN(n4700) );
  INV_X1 U6138 ( .A(n8962), .ZN(n4962) );
  NOR2_X1 U6139 ( .A1(n7330), .A2(n7166), .ZN(n8908) );
  AND2_X1 U6140 ( .A1(n7396), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4434) );
  NOR3_X1 U6141 ( .A1(n10103), .A2(n10091), .A3(n10102), .ZN(n4435) );
  AND2_X1 U6142 ( .A1(n7188), .A2(n7750), .ZN(n6528) );
  INV_X1 U6143 ( .A(n5535), .ZN(n5845) );
  INV_X1 U6144 ( .A(n7291), .ZN(n4709) );
  OR2_X1 U6145 ( .A1(n9237), .A2(n9039), .ZN(n7308) );
  AND3_X1 U6146 ( .A1(n7377), .A2(n4984), .A3(n7376), .ZN(n4436) );
  AND3_X1 U6147 ( .A1(n5132), .A2(n7463), .A3(n7522), .ZN(n4437) );
  NAND2_X1 U6148 ( .A1(n7127), .A2(n10027), .ZN(n4438) );
  OR2_X1 U6149 ( .A1(n6497), .A2(n7369), .ZN(n4440) );
  AND2_X1 U6150 ( .A1(n9483), .A2(n9588), .ZN(n4441) );
  INV_X1 U6151 ( .A(n8277), .ZN(n4878) );
  OR2_X1 U6152 ( .A1(n10146), .A2(n9929), .ZN(n7036) );
  INV_X1 U6153 ( .A(n7036), .ZN(n4697) );
  NOR2_X1 U6154 ( .A1(n5653), .A2(n5651), .ZN(n4442) );
  AND2_X1 U6155 ( .A1(n8338), .A2(n4878), .ZN(n4443) );
  OR2_X1 U6156 ( .A1(n4785), .A2(n4405), .ZN(n4444) );
  NAND2_X1 U6157 ( .A1(n5802), .A2(n5801), .ZN(n7150) );
  NAND2_X1 U6158 ( .A1(n5623), .A2(n5622), .ZN(n10159) );
  AND2_X1 U6159 ( .A1(n5019), .A2(n9639), .ZN(n4445) );
  NAND2_X1 U6160 ( .A1(n7484), .A2(n4610), .ZN(n4609) );
  AND2_X1 U6161 ( .A1(n10129), .A2(n9919), .ZN(n4446) );
  AND2_X1 U6162 ( .A1(n4794), .A2(n7137), .ZN(n4447) );
  INV_X1 U6163 ( .A(n7149), .ZN(n8892) );
  AND2_X1 U6164 ( .A1(n7048), .A2(n5941), .ZN(n7149) );
  AND4_X1 U6165 ( .A1(n5489), .A2(n5488), .A3(n5487), .A4(n5486), .ZN(n8286)
         );
  XOR2_X1 U6166 ( .A(n7151), .B(n10091), .Z(n4448) );
  INV_X1 U6167 ( .A(n4859), .ZN(n6575) );
  NOR2_X1 U6168 ( .A1(n9235), .A2(n4860), .ZN(n4859) );
  AND2_X1 U6169 ( .A1(n7293), .A2(n7291), .ZN(n9275) );
  INV_X1 U6170 ( .A(n9275), .ZN(n6549) );
  AND2_X1 U6171 ( .A1(n6212), .A2(n6211), .ZN(n4449) );
  NAND2_X1 U6172 ( .A1(n9498), .A2(n6468), .ZN(n7311) );
  NAND2_X1 U6173 ( .A1(n6253), .A2(n6252), .ZN(n4450) );
  NOR2_X1 U6174 ( .A1(n9331), .A2(n9528), .ZN(n9301) );
  OR2_X1 U6175 ( .A1(n7293), .A2(n7340), .ZN(n4451) );
  AND2_X1 U6176 ( .A1(n10141), .A2(n9921), .ZN(n4452) );
  INV_X1 U6177 ( .A(n4854), .ZN(n9302) );
  NOR2_X1 U6178 ( .A1(n9331), .A2(n4855), .ZN(n4854) );
  AND2_X1 U6179 ( .A1(n5241), .A2(n5501), .ZN(n4453) );
  NOR2_X1 U6180 ( .A1(n10127), .A2(n9905), .ZN(n4454) );
  NAND2_X1 U6181 ( .A1(n9366), .A2(n4926), .ZN(n9368) );
  INV_X1 U6182 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6255) );
  INV_X1 U6183 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6785) );
  INV_X1 U6184 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6512) );
  NOR2_X1 U6185 ( .A1(n9493), .A2(n9220), .ZN(n4455) );
  NAND2_X1 U6186 ( .A1(n8677), .A2(n8680), .ZN(n4456) );
  OR2_X1 U6187 ( .A1(n9539), .A2(n9359), .ZN(n4457) );
  INV_X1 U6188 ( .A(n4972), .ZN(n4971) );
  NAND2_X1 U6189 ( .A1(n4977), .A2(n4976), .ZN(n4972) );
  AND2_X1 U6190 ( .A1(n7296), .A2(n9250), .ZN(n4458) );
  NAND2_X1 U6191 ( .A1(n5482), .A2(n5481), .ZN(n8080) );
  AND2_X1 U6192 ( .A1(n5258), .A2(SI_11_), .ZN(n4459) );
  AND2_X1 U6193 ( .A1(n7175), .A2(n4989), .ZN(n4460) );
  INV_X1 U6194 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7424) );
  AND2_X1 U6195 ( .A1(n10017), .A2(n10000), .ZN(n9985) );
  AND2_X1 U6196 ( .A1(n9931), .A2(n5024), .ZN(n9857) );
  NAND2_X1 U6197 ( .A1(n8437), .A2(n8436), .ZN(n4461) );
  OAI21_X1 U6198 ( .B1(n9366), .B2(n4621), .A(n4619), .ZN(n9339) );
  OAI21_X1 U6199 ( .B1(n4575), .B2(n4578), .A(n8039), .ZN(n4574) );
  OR2_X1 U6200 ( .A1(n4801), .A2(n7111), .ZN(n4462) );
  OR2_X1 U6201 ( .A1(n9639), .A2(n9771), .ZN(n4463) );
  OR2_X1 U6202 ( .A1(n7267), .A2(n9378), .ZN(n4464) );
  NOR2_X1 U6203 ( .A1(n10012), .A2(n7121), .ZN(n4465) );
  AND2_X1 U6204 ( .A1(n6084), .A2(n4981), .ZN(n4466) );
  AND2_X1 U6205 ( .A1(n5921), .A2(n5866), .ZN(n4467) );
  AND2_X1 U6206 ( .A1(n4868), .A2(n9643), .ZN(n4468) );
  AND2_X1 U6207 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n4469) );
  AND2_X1 U6208 ( .A1(n4868), .A2(n4866), .ZN(n4470) );
  AND2_X1 U6209 ( .A1(n4699), .A2(n5934), .ZN(n4471) );
  INV_X1 U6210 ( .A(n9237), .ZN(n9503) );
  NAND2_X1 U6211 ( .A1(n6448), .A2(n6447), .ZN(n9237) );
  AND2_X1 U6212 ( .A1(n7293), .A2(n7349), .ZN(n4472) );
  INV_X1 U6213 ( .A(n7452), .ZN(n4600) );
  AND2_X1 U6214 ( .A1(n4843), .A2(n8233), .ZN(n4473) );
  XNOR2_X1 U6215 ( .A(n5257), .B(SI_11_), .ZN(n5555) );
  INV_X1 U6216 ( .A(n9493), .ZN(n9207) );
  NAND2_X1 U6217 ( .A1(n6472), .A2(n6471), .ZN(n9493) );
  AND2_X1 U6218 ( .A1(n8948), .A2(n7048), .ZN(n4474) );
  OAI21_X1 U6219 ( .B1(n8900), .B2(n7173), .A(n7332), .ZN(n7167) );
  AND2_X1 U6220 ( .A1(n9280), .A2(n5002), .ZN(n4475) );
  INV_X1 U6221 ( .A(n4606), .ZN(n4605) );
  OAI21_X1 U6222 ( .B1(n4609), .B2(n4608), .A(n4607), .ZN(n4606) );
  AND2_X1 U6223 ( .A1(n6279), .A2(n6278), .ZN(n4476) );
  AND2_X1 U6224 ( .A1(n4716), .A2(n4451), .ZN(n4477) );
  INV_X1 U6225 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5079) );
  NOR2_X1 U6226 ( .A1(n7856), .A2(n6828), .ZN(n4478) );
  AND2_X1 U6227 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n4479) );
  OR2_X1 U6228 ( .A1(n4876), .A2(n4443), .ZN(n4480) );
  INV_X1 U6229 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5143) );
  AND2_X1 U6230 ( .A1(n7308), .A2(n7301), .ZN(n9228) );
  INV_X2 U6231 ( .A(n10078), .ZN(n10020) );
  NAND2_X1 U6232 ( .A1(n7156), .A2(n10049), .ZN(n10078) );
  INV_X1 U6233 ( .A(n9411), .ZN(n10467) );
  AND2_X1 U6234 ( .A1(n8506), .A2(n4419), .ZN(n8631) );
  INV_X1 U6235 ( .A(n9760), .ZN(n9772) );
  NAND2_X1 U6236 ( .A1(n6569), .A2(n8554), .ZN(n8213) );
  NAND2_X1 U6237 ( .A1(n7476), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4481) );
  AND2_X1 U6238 ( .A1(n9399), .A2(n7264), .ZN(n9376) );
  AND2_X1 U6239 ( .A1(n7640), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4482) );
  INV_X1 U6240 ( .A(n9528), .ZN(n4856) );
  NAND2_X1 U6241 ( .A1(n5747), .A2(n5746), .ZN(n10127) );
  INV_X1 U6242 ( .A(n10127), .ZN(n5025) );
  NAND2_X1 U6243 ( .A1(n5693), .A2(n5692), .ZN(n10146) );
  INV_X1 U6244 ( .A(n10146), .ZN(n5022) );
  NAND2_X1 U6245 ( .A1(n9415), .A2(n7253), .ZN(n8667) );
  AND2_X1 U6246 ( .A1(n4775), .A2(n4438), .ZN(n10025) );
  INV_X1 U6247 ( .A(n10065), .ZN(n4825) );
  XNOR2_X1 U6248 ( .A(n9237), .B(n6719), .ZN(n9087) );
  NAND2_X1 U6249 ( .A1(n5384), .A2(n5383), .ZN(n10092) );
  INV_X1 U6250 ( .A(n10064), .ZN(n4822) );
  INV_X1 U6251 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n4802) );
  AND2_X1 U6252 ( .A1(n4633), .A2(n4631), .ZN(n4483) );
  NOR2_X1 U6253 ( .A1(n7482), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4484) );
  INV_X1 U6254 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8139) );
  NOR2_X1 U6255 ( .A1(n5059), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4509) );
  INV_X1 U6256 ( .A(n4632), .ZN(n4631) );
  NAND2_X1 U6257 ( .A1(n4635), .A2(n5154), .ZN(n4632) );
  INV_X1 U6258 ( .A(n4892), .ZN(n4891) );
  NAND2_X1 U6259 ( .A1(n4897), .A2(n9760), .ZN(n4892) );
  AND2_X1 U6260 ( .A1(n4811), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n4485) );
  OR2_X1 U6261 ( .A1(n4745), .A2(n4746), .ZN(n4486) );
  AND2_X1 U6262 ( .A1(n4750), .A2(n4481), .ZN(n4487) );
  OR2_X1 U6263 ( .A1(n6728), .A2(n6562), .ZN(n9419) );
  INV_X1 U6264 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n4812) );
  OR2_X1 U6265 ( .A1(n8107), .A2(n8109), .ZN(n5016) );
  INV_X1 U6266 ( .A(n5016), .ZN(n5015) );
  NAND2_X1 U6267 ( .A1(n6238), .A2(n6237), .ZN(n8126) );
  INV_X1 U6268 ( .A(n8126), .ZN(n4845) );
  INV_X1 U6269 ( .A(n9580), .ZN(n4543) );
  NOR2_X1 U6270 ( .A1(n7153), .A2(n7982), .ZN(n7732) );
  INV_X1 U6271 ( .A(n10074), .ZN(n10044) );
  NAND2_X1 U6272 ( .A1(n7053), .A2(n7052), .ZN(n10074) );
  NOR2_X1 U6273 ( .A1(n7645), .A2(n6137), .ZN(n4488) );
  INV_X1 U6274 ( .A(n10193), .ZN(n5017) );
  NOR2_X1 U6275 ( .A1(n10276), .A2(n4410), .ZN(n4489) );
  OR2_X1 U6276 ( .A1(n9177), .A2(n6369), .ZN(n4490) );
  INV_X1 U6277 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n4813) );
  NAND2_X1 U6278 ( .A1(n4980), .A2(n4979), .ZN(n7910) );
  NAND2_X1 U6279 ( .A1(n6568), .A2(n8196), .ZN(n7748) );
  INV_X1 U6280 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4758) );
  AND2_X1 U6281 ( .A1(n4814), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n4491) );
  AND2_X1 U6282 ( .A1(n4753), .A2(n4752), .ZN(n4492) );
  INV_X1 U6283 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4757) );
  INV_X1 U6284 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n4539) );
  INV_X1 U6285 ( .A(n7384), .ZN(n4676) );
  NAND2_X1 U6286 ( .A1(n6115), .A2(n6114), .ZN(n7998) );
  OR2_X1 U6287 ( .A1(n9813), .A2(n5165), .ZN(n4493) );
  INV_X1 U6288 ( .A(n7396), .ZN(n5010) );
  AND2_X1 U6289 ( .A1(n6043), .A2(n6042), .ZN(n7537) );
  INV_X1 U6290 ( .A(n9152), .ZN(n4745) );
  NAND2_X1 U6291 ( .A1(n9416), .A2(n9424), .ZN(n9415) );
  NAND2_X1 U6292 ( .A1(n9399), .A2(n4546), .ZN(n4545) );
  NAND2_X1 U6293 ( .A1(n9345), .A2(n9352), .ZN(n9344) );
  NAND2_X1 U6294 ( .A1(n8669), .A2(n7257), .ZN(n9398) );
  NOR3_X1 U6295 ( .A1(n9326), .A2(n9311), .A3(n9321), .ZN(n9310) );
  AOI21_X1 U6296 ( .B1(n7777), .B2(n7778), .A(n7192), .ZN(n9442) );
  OAI22_X2 U6297 ( .A1(n7904), .A2(n7903), .B1(n6625), .B2(n6624), .ZN(n7986)
         );
  NAND2_X1 U6298 ( .A1(n4963), .A2(n4965), .ZN(n9055) );
  NAND2_X1 U6299 ( .A1(n9015), .A2(n4534), .ZN(n9025) );
  AOI21_X1 U6300 ( .B1(n8165), .B2(n8166), .A(n6652), .ZN(n8994) );
  AOI21_X2 U6301 ( .B1(n8949), .B2(n10074), .A(n4494), .ZN(n10110) );
  NAND2_X1 U6302 ( .A1(n7018), .A2(n7017), .ZN(n8509) );
  NAND2_X1 U6303 ( .A1(n4535), .A2(n7037), .ZN(n9927) );
  NAND2_X1 U6304 ( .A1(n7725), .A2(n5872), .ZN(n5414) );
  NAND2_X1 U6305 ( .A1(n4523), .A2(n10106), .ZN(n10203) );
  NAND2_X1 U6306 ( .A1(n5413), .A2(n5414), .ZN(n5962) );
  NAND2_X2 U6307 ( .A1(n5505), .A2(n5504), .ZN(n10427) );
  INV_X1 U6308 ( .A(n4674), .ZN(n4673) );
  OAI21_X2 U6309 ( .B1(n4428), .B2(n4496), .A(n7951), .ZN(n7954) );
  OAI21_X2 U6310 ( .B1(n8237), .B2(n8019), .A(n8018), .ZN(n8024) );
  INV_X4 U6311 ( .A(n5407), .ZN(n5655) );
  NAND2_X1 U6312 ( .A1(n7803), .A2(n7950), .ZN(n4496) );
  NAND2_X1 U6313 ( .A1(n5148), .A2(n5108), .ZN(n5102) );
  NAND2_X2 U6314 ( .A1(n7720), .A2(n7993), .ZN(n7619) );
  OAI21_X1 U6315 ( .B1(n9691), .B2(n9764), .A(n9772), .ZN(n9695) );
  NAND2_X1 U6316 ( .A1(n7868), .A2(n7869), .ZN(n7803) );
  NAND2_X1 U6317 ( .A1(n7809), .A2(n7810), .ZN(n8003) );
  OAI21_X2 U6318 ( .B1(n9883), .B2(n7047), .A(n7046), .ZN(n8893) );
  NAND2_X1 U6319 ( .A1(n5962), .A2(n8090), .ZN(n5423) );
  NAND2_X1 U6320 ( .A1(n7038), .A2(n7139), .ZN(n9925) );
  NAND2_X1 U6321 ( .A1(n5795), .A2(n5337), .ZN(n5340) );
  NAND2_X1 U6322 ( .A1(n5855), .A2(n5856), .ZN(n4680) );
  NAND3_X1 U6323 ( .A1(n5354), .A2(n5355), .A3(n4497), .ZN(n5840) );
  AOI21_X1 U6324 ( .B1(n5304), .B2(n4650), .A(n4646), .ZN(n4645) );
  NAND2_X1 U6325 ( .A1(n5756), .A2(n5330), .ZN(n4661) );
  NAND2_X1 U6326 ( .A1(n4500), .A2(n5043), .ZN(n5705) );
  NAND2_X1 U6327 ( .A1(n5614), .A2(n4501), .ZN(n4500) );
  OAI21_X1 U6328 ( .B1(n5774), .B2(n9886), .A(n4503), .ZN(n4502) );
  OR2_X1 U6329 ( .A1(n5775), .A2(n7089), .ZN(n4503) );
  NAND2_X1 U6330 ( .A1(n4504), .A2(n4527), .ZN(n4526) );
  NAND2_X1 U6331 ( .A1(n4505), .A2(n4467), .ZN(n4504) );
  NAND2_X1 U6332 ( .A1(n5583), .A2(n7015), .ZN(n4505) );
  NAND2_X1 U6333 ( .A1(n5474), .A2(n5868), .ZN(n5457) );
  NAND2_X2 U6334 ( .A1(n7936), .A2(n5971), .ZN(n8101) );
  OAI21_X1 U6335 ( .B1(n5493), .B2(n5476), .A(n5867), .ZN(n5492) );
  NAND2_X1 U6336 ( .A1(n6361), .A2(n7268), .ZN(n9378) );
  INV_X4 U6337 ( .A(n5225), .ZN(n7389) );
  NAND2_X1 U6338 ( .A1(n4413), .A2(n4464), .ZN(n4729) );
  OAI21_X1 U6339 ( .B1(n4436), .B2(n4507), .A(n7382), .ZN(P2_U3244) );
  INV_X1 U6340 ( .A(n7288), .ZN(n7285) );
  OAI21_X2 U6341 ( .B1(n5546), .B2(n5545), .A(n5263), .ZN(n5534) );
  NAND2_X1 U6342 ( .A1(n4918), .A2(n4919), .ZN(n5546) );
  NAND2_X1 U6343 ( .A1(n7060), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5058) );
  INV_X1 U6344 ( .A(n4509), .ZN(n7060) );
  NAND2_X2 U6345 ( .A1(n8849), .A2(n8848), .ZN(n9764) );
  NAND2_X1 U6346 ( .A1(n10105), .A2(n10104), .ZN(n4524) );
  NAND3_X1 U6347 ( .A1(n4770), .A2(n4769), .A3(n4510), .ZN(n4775) );
  OAI21_X2 U6348 ( .B1(n7136), .B2(n4791), .A(n4789), .ZN(n9909) );
  OR2_X1 U6349 ( .A1(n6632), .A2(n6631), .ZN(n6634) );
  NAND2_X1 U6350 ( .A1(n8963), .A2(n8962), .ZN(n8961) );
  NAND2_X1 U6351 ( .A1(n7419), .A2(n7176), .ZN(n4544) );
  NAND2_X2 U6352 ( .A1(n7020), .A2(n7019), .ZN(n8559) );
  NAND2_X1 U6353 ( .A1(n4830), .A2(n7041), .ZN(n9901) );
  NAND3_X1 U6354 ( .A1(n7227), .A2(n7226), .A3(n7228), .ZN(n4517) );
  NAND2_X1 U6355 ( .A1(n4727), .A2(n4728), .ZN(n7288) );
  NAND2_X1 U6356 ( .A1(n4760), .A2(n4759), .ZN(n9867) );
  NOR2_X1 U6357 ( .A1(n4768), .A2(n7119), .ZN(n4767) );
  NAND3_X1 U6358 ( .A1(n7347), .A2(n4984), .A3(n4519), .ZN(n4731) );
  NAND2_X1 U6359 ( .A1(n4873), .A2(n4871), .ZN(n8747) );
  NAND2_X1 U6360 ( .A1(n9632), .A2(n8878), .ZN(n8879) );
  NAND2_X1 U6361 ( .A1(n8946), .A2(n7049), .ZN(n7050) );
  AOI21_X2 U6362 ( .B1(n7059), .B2(n10074), .A(n7058), .ZN(n10106) );
  NAND2_X1 U6363 ( .A1(n5513), .A2(n5039), .ZN(n5251) );
  NAND2_X1 U6364 ( .A1(n5534), .A2(n5040), .ZN(n5268) );
  XNOR2_X1 U6365 ( .A(n5221), .B(SI_4_), .ZN(n5440) );
  NOR2_X1 U6366 ( .A1(n9944), .A2(n7035), .ZN(n5045) );
  OAI211_X1 U6367 ( .C1(n10111), .C2(n10102), .A(n10110), .B(n10109), .ZN(
        n10204) );
  OAI211_X1 U6368 ( .C1(n5603), .C2(n5602), .A(n4526), .B(n5601), .ZN(n5614)
         );
  AND2_X1 U6369 ( .A1(n5582), .A2(n5032), .ZN(n4527) );
  INV_X1 U6370 ( .A(n5892), .ZN(n5891) );
  AOI21_X1 U6371 ( .B1(n4701), .B2(n4471), .A(n4691), .ZN(n5770) );
  NAND3_X1 U6372 ( .A1(n4900), .A2(n4901), .A3(n4994), .ZN(n9232) );
  NAND2_X1 U6373 ( .A1(n4915), .A2(n4913), .ZN(n8905) );
  NAND2_X1 U6374 ( .A1(n8224), .A2(n6303), .ZN(n8662) );
  NAND2_X1 U6375 ( .A1(n4670), .A2(n4668), .ZN(P2_U3517) );
  NAND2_X1 U6376 ( .A1(n4850), .A2(n4848), .ZN(P2_U3549) );
  AOI21_X2 U6377 ( .B1(n9305), .B2(n6412), .A(n4532), .ZN(n9276) );
  AND2_X1 U6378 ( .A1(n9523), .A2(n9314), .ZN(n4532) );
  NAND2_X1 U6379 ( .A1(n4908), .A2(n4906), .ZN(n9305) );
  OAI21_X1 U6380 ( .B1(n8291), .B2(n6292), .A(n6291), .ZN(n8225) );
  NAND2_X1 U6381 ( .A1(n9047), .A2(n9046), .ZN(n9045) );
  OAI22_X2 U6382 ( .A1(n9055), .A2(n9054), .B1(n6689), .B2(n6688), .ZN(n8984)
         );
  NAND2_X1 U6383 ( .A1(n9680), .A2(n9679), .ZN(n4881) );
  AND2_X2 U6384 ( .A1(n4898), .A2(n4896), .ZN(n9632) );
  NAND2_X1 U6385 ( .A1(n4865), .A2(n4864), .ZN(n9696) );
  NOR2_X2 U6386 ( .A1(n5360), .A2(n5359), .ZN(n5362) );
  NAND2_X1 U6387 ( .A1(n4838), .A2(n4840), .ZN(n4535) );
  NAND2_X1 U6388 ( .A1(n8895), .A2(n4474), .ZN(n8946) );
  INV_X1 U6389 ( .A(n8893), .ZN(n4536) );
  OAI21_X1 U6390 ( .B1(n5459), .B2(n5243), .A(n4537), .ZN(n5245) );
  NAND2_X1 U6391 ( .A1(n4732), .A2(n7323), .ZN(n7336) );
  INV_X1 U6392 ( .A(n4708), .ZN(n4707) );
  NAND2_X1 U6393 ( .A1(n4718), .A2(n4712), .ZN(n4711) );
  NAND2_X1 U6394 ( .A1(n4717), .A2(n4477), .ZN(n4704) );
  OAI21_X1 U6395 ( .B1(n4704), .B2(n4703), .A(n4458), .ZN(n7300) );
  INV_X1 U6396 ( .A(n7324), .ZN(n4732) );
  OAI21_X1 U6397 ( .B1(n7284), .B2(n4707), .A(n4705), .ZN(n4717) );
  AOI21_X1 U6398 ( .B1(n7314), .B2(n7313), .A(n5041), .ZN(n4734) );
  OR2_X1 U6399 ( .A1(n7645), .A2(n4572), .ZN(n4570) );
  NAND2_X1 U6400 ( .A1(n4568), .A2(n4567), .ZN(n8483) );
  NAND2_X1 U6401 ( .A1(n7645), .A2(n4433), .ZN(n4568) );
  NAND2_X1 U6402 ( .A1(n7645), .A2(n4578), .ZN(n4573) );
  INV_X1 U6403 ( .A(n4576), .ZN(n4575) );
  AOI21_X1 U6404 ( .B1(n6137), .B2(n4578), .A(n4478), .ZN(n4576) );
  INV_X1 U6405 ( .A(n7853), .ZN(n4578) );
  NAND2_X2 U6406 ( .A1(n9882), .A2(n7043), .ZN(n9883) );
  NOR2_X1 U6407 ( .A1(n10278), .A2(n10277), .ZN(n10276) );
  INV_X1 U6408 ( .A(n10278), .ZN(n4596) );
  INV_X1 U6409 ( .A(n7694), .ZN(n4602) );
  INV_X1 U6410 ( .A(n7453), .ZN(n4598) );
  OAI21_X1 U6411 ( .B1(n9815), .B2(n4606), .A(n4603), .ZN(n7469) );
  NOR2_X2 U6412 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n6016) );
  NAND2_X1 U6413 ( .A1(n9366), .A2(n4619), .ZN(n4617) );
  NAND3_X1 U6414 ( .A1(n4617), .A2(n4618), .A3(n4909), .ZN(n4908) );
  OAI21_X2 U6415 ( .B1(n8662), .B2(n4456), .A(n6340), .ZN(n9410) );
  NAND2_X1 U6416 ( .A1(n7746), .A2(n6527), .ZN(n7745) );
  AOI21_X1 U6417 ( .B1(n7745), .B2(n6249), .A(n4450), .ZN(n8291) );
  INV_X1 U6418 ( .A(n4639), .ZN(n8134) );
  INV_X1 U6419 ( .A(n4645), .ZN(n5743) );
  NAND3_X1 U6420 ( .A1(n4993), .A2(n4992), .A3(n4995), .ZN(n4657) );
  NAND2_X1 U6421 ( .A1(n5325), .A2(n5324), .ZN(n5756) );
  NAND2_X1 U6422 ( .A1(n5325), .A2(n4659), .ZN(n4658) );
  OR2_X1 U6423 ( .A1(n4672), .A2(n5143), .ZN(n5133) );
  NAND3_X1 U6424 ( .A1(n5081), .A2(n4672), .A3(n4403), .ZN(n5086) );
  NAND4_X2 U6425 ( .A1(n5081), .A2(n4672), .A3(n4403), .A4(n5011), .ZN(n5360)
         );
  NAND2_X1 U6426 ( .A1(n5066), .A2(n4672), .ZN(n5183) );
  NAND2_X2 U6427 ( .A1(n4673), .A2(n5422), .ZN(n7873) );
  NAND2_X1 U6428 ( .A1(n5457), .A2(n4425), .ZN(n4681) );
  OAI21_X1 U6429 ( .B1(n5457), .B2(n5854), .A(n4425), .ZN(n5493) );
  NAND2_X1 U6430 ( .A1(n4681), .A2(n4682), .ZN(n5495) );
  NAND3_X1 U6431 ( .A1(n4690), .A2(n4699), .A3(n7039), .ZN(n4689) );
  INV_X1 U6432 ( .A(n5773), .ZN(n4690) );
  INV_X1 U6433 ( .A(n9886), .ZN(n4692) );
  NAND2_X1 U6434 ( .A1(n7209), .A2(n4725), .ZN(n4721) );
  NAND2_X1 U6435 ( .A1(n7210), .A2(n4720), .ZN(n4719) );
  NAND3_X1 U6436 ( .A1(n4721), .A2(n4724), .A3(n4719), .ZN(n4723) );
  NAND2_X1 U6437 ( .A1(n4722), .A2(n7224), .ZN(n7227) );
  NAND2_X1 U6438 ( .A1(n4723), .A2(n7221), .ZN(n4722) );
  INV_X1 U6439 ( .A(n7217), .ZN(n4725) );
  NAND3_X1 U6440 ( .A1(n7262), .A2(n9409), .A3(n4413), .ZN(n4727) );
  NAND3_X1 U6441 ( .A1(n6100), .A2(n6101), .A3(n5007), .ZN(n6124) );
  AND3_X2 U6442 ( .A1(n4736), .A2(n6041), .A3(n4735), .ZN(n6101) );
  NOR2_X2 U6443 ( .A1(n6099), .A2(n6098), .ZN(n6100) );
  NAND4_X1 U6444 ( .A1(n6091), .A2(n6092), .A3(n6090), .A4(n6089), .ZN(n6099)
         );
  INV_X1 U6445 ( .A(n9185), .ZN(n4742) );
  NAND2_X1 U6446 ( .A1(n9141), .A2(n4744), .ZN(n4743) );
  OAI211_X1 U6447 ( .C1(n6075), .C2(n4746), .A(n4743), .B(n4486), .ZN(n9167)
         );
  NAND2_X1 U6448 ( .A1(n9139), .A2(n6075), .ZN(n9151) );
  AND2_X1 U6449 ( .A1(n6351), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4746) );
  NAND2_X1 U6450 ( .A1(n8708), .A2(n4749), .ZN(n4747) );
  NAND2_X1 U6451 ( .A1(n4747), .A2(n4748), .ZN(n9126) );
  INV_X1 U6452 ( .A(n4750), .ZN(n8707) );
  INV_X1 U6453 ( .A(n4753), .ZN(n7591) );
  NAND3_X1 U6454 ( .A1(n4756), .A2(n4758), .A3(n4757), .ZN(n5077) );
  NAND2_X1 U6455 ( .A1(n7142), .A2(n4761), .ZN(n4760) );
  INV_X1 U6456 ( .A(n7117), .ZN(n4768) );
  NAND2_X1 U6457 ( .A1(n5378), .A2(n10234), .ZN(n5464) );
  XNOR2_X2 U6458 ( .A(n4777), .B(n4776), .ZN(n10234) );
  OR2_X1 U6459 ( .A1(n9855), .A2(n4779), .ZN(n4778) );
  NAND2_X1 U6460 ( .A1(n9855), .A2(n4785), .ZN(n4784) );
  OAI21_X1 U6461 ( .B1(n4797), .B2(n7108), .A(n4800), .ZN(n4799) );
  NAND3_X1 U6462 ( .A1(n4798), .A2(n8315), .A3(n7110), .ZN(n4797) );
  NOR2_X1 U6463 ( .A1(n7108), .A2(n7107), .ZN(n8316) );
  INV_X1 U6464 ( .A(n4799), .ZN(n8504) );
  NOR2_X1 U6465 ( .A1(n8075), .A2(n7101), .ZN(n7108) );
  INV_X1 U6466 ( .A(n8109), .ZN(n10388) );
  NAND2_X1 U6467 ( .A1(n9803), .A2(n10388), .ZN(n7096) );
  INV_X1 U6468 ( .A(n7097), .ZN(n9803) );
  NAND2_X1 U6469 ( .A1(n7724), .A2(n7726), .ZN(n7931) );
  NAND3_X1 U6470 ( .A1(n5941), .A2(n7089), .A3(n4804), .ZN(n4803) );
  NAND2_X1 U6471 ( .A1(n5374), .A2(n4485), .ZN(n5711) );
  NAND2_X1 U6472 ( .A1(n5375), .A2(n4491), .ZN(n5760) );
  INV_X1 U6473 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n4815) );
  NAND2_X1 U6474 ( .A1(n4816), .A2(n4479), .ZN(n5516) );
  INV_X1 U6475 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n4819) );
  NAND2_X1 U6476 ( .A1(n4820), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6477 ( .A1(n5085), .A2(n4820), .ZN(n5159) );
  NAND2_X1 U6478 ( .A1(n5084), .A2(n5083), .ZN(n4820) );
  NAND2_X1 U6479 ( .A1(n8068), .A2(n8067), .ZN(n4828) );
  NAND2_X1 U6480 ( .A1(n7027), .A2(n7026), .ZN(n10010) );
  NAND2_X1 U6481 ( .A1(n6100), .A2(n6101), .ZN(n6122) );
  NAND2_X1 U6482 ( .A1(n6569), .A2(n4473), .ZN(n8660) );
  NAND2_X1 U6483 ( .A1(n8306), .A2(n8364), .ZN(n8305) );
  NOR2_X2 U6484 ( .A1(n9331), .A2(n4852), .ZN(n9244) );
  NAND2_X1 U6485 ( .A1(n9234), .A2(n9503), .ZN(n9235) );
  INV_X1 U6486 ( .A(n4861), .ZN(n7867) );
  NAND2_X1 U6487 ( .A1(n7798), .A2(n7797), .ZN(n4861) );
  NAND2_X1 U6488 ( .A1(n9640), .A2(n4468), .ZN(n4864) );
  NAND2_X1 U6489 ( .A1(n4870), .A2(n9641), .ZN(n4867) );
  NAND2_X1 U6490 ( .A1(n8762), .A2(n4869), .ZN(n4868) );
  NAND2_X1 U6491 ( .A1(n9776), .A2(n9775), .ZN(n9773) );
  NAND3_X1 U6492 ( .A1(n4870), .A2(n9641), .A3(n8762), .ZN(n9776) );
  NAND2_X1 U6493 ( .A1(n4881), .A2(n8817), .ZN(n8823) );
  NAND2_X1 U6494 ( .A1(n4881), .A2(n4879), .ZN(n9742) );
  NAND2_X1 U6495 ( .A1(n4883), .A2(n4882), .ZN(n8809) );
  NAND2_X1 U6496 ( .A1(n9764), .A2(n4888), .ZN(n4886) );
  OAI211_X1 U6497 ( .C1(n9764), .C2(n4890), .A(n4886), .B(n4887), .ZN(P1_U3212) );
  NAND2_X1 U6498 ( .A1(n9259), .A2(n4903), .ZN(n4900) );
  INV_X1 U6499 ( .A(n9339), .ZN(n4912) );
  OAI21_X1 U6500 ( .B1(n4910), .B2(n4404), .A(n4420), .ZN(n4907) );
  NAND2_X1 U6501 ( .A1(n9213), .A2(n4916), .ZN(n4915) );
  NAND2_X1 U6502 ( .A1(n9213), .A2(n6470), .ZN(n9210) );
  NAND2_X1 U6503 ( .A1(n5251), .A2(n4920), .ZN(n4918) );
  NAND2_X1 U6504 ( .A1(n5251), .A2(n5250), .ZN(n5571) );
  NAND2_X1 U6505 ( .A1(n5268), .A2(n4928), .ZN(n4927) );
  NAND3_X1 U6506 ( .A1(n5197), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4938) );
  NAND3_X1 U6507 ( .A1(n4942), .A2(n4941), .A3(n4940), .ZN(n4939) );
  INV_X1 U6508 ( .A(n4384), .ZN(n6553) );
  NAND3_X1 U6509 ( .A1(n6584), .A2(n7187), .A3(n7998), .ZN(n4943) );
  NAND2_X1 U6510 ( .A1(n8373), .A2(n4407), .ZN(n4945) );
  INV_X1 U6511 ( .A(n8373), .ZN(n4949) );
  NAND2_X1 U6512 ( .A1(n6714), .A2(n4951), .ZN(n4950) );
  OAI211_X1 U6513 ( .C1(n6714), .C2(n4955), .A(n4952), .B(n4950), .ZN(n6743)
         );
  NAND2_X1 U6514 ( .A1(n6714), .A2(n6713), .ZN(n8963) );
  NAND2_X1 U6515 ( .A1(n9025), .A2(n4964), .ZN(n4963) );
  AND2_X1 U6516 ( .A1(n6622), .A2(n6616), .ZN(n4979) );
  NAND2_X1 U6517 ( .A1(n6085), .A2(n4982), .ZN(n6112) );
  NAND2_X1 U6518 ( .A1(n6101), .A2(n6084), .ZN(n6142) );
  INV_X1 U6519 ( .A(n6112), .ZN(n6087) );
  NAND2_X1 U6520 ( .A1(n7186), .A2(n5036), .ZN(n4984) );
  INV_X1 U6521 ( .A(n8907), .ZN(n4988) );
  NAND2_X1 U6522 ( .A1(n8907), .A2(n8908), .ZN(n8910) );
  NAND2_X1 U6523 ( .A1(n6551), .A2(n4999), .ZN(n5001) );
  INV_X1 U6524 ( .A(n6550), .ZN(n5000) );
  OAI21_X1 U6525 ( .B1(n5002), .B2(n6552), .A(n5001), .ZN(n9251) );
  NAND3_X1 U6526 ( .A1(n6534), .A2(n6533), .A3(n4422), .ZN(n8172) );
  AND2_X1 U6527 ( .A1(n6534), .A2(n6533), .ZN(n5004) );
  OAI21_X1 U6528 ( .B1(n4422), .B2(n5004), .A(n8172), .ZN(n8173) );
  NAND3_X1 U6529 ( .A1(n6101), .A2(n6100), .A3(n5008), .ZN(n6157) );
  NAND2_X1 U6530 ( .A1(n8093), .A2(n5009), .ZN(n10375) );
  NAND2_X1 U6531 ( .A1(n7732), .A2(n8092), .ZN(n5009) );
  NAND2_X1 U6532 ( .A1(n5491), .A2(n8346), .ZN(n5014) );
  BUF_X4 U6533 ( .A(n8004), .Z(n8869) );
  NAND2_X1 U6534 ( .A1(n9198), .A2(n6748), .ZN(n8903) );
  NAND2_X1 U6535 ( .A1(n6572), .A2(n6571), .ZN(n9430) );
  OR2_X1 U6536 ( .A1(n8915), .A2(n8900), .ZN(n6748) );
  OR2_X1 U6537 ( .A1(n6197), .A2(n7568), .ZN(n6185) );
  AND2_X1 U6538 ( .A1(n9252), .A2(n6670), .ZN(n9001) );
  AND2_X1 U6539 ( .A1(n9114), .A2(n6670), .ZN(n9034) );
  INV_X1 U6540 ( .A(n6525), .ZN(n7777) );
  NAND2_X1 U6542 ( .A1(n8053), .A2(n5854), .ZN(n5443) );
  INV_X1 U6543 ( .A(n9301), .ZN(n9317) );
  NAND2_X1 U6544 ( .A1(n7154), .A2(n10380), .ZN(n8107) );
  NAND4_X1 U6545 ( .A1(n6183), .A2(n6182), .A3(n6181), .A4(n6180), .ZN(n6198)
         );
  OR2_X1 U6546 ( .A1(n5464), .A2(n10440), .ZN(n5416) );
  OR2_X1 U6547 ( .A1(n5464), .A2(n5124), .ZN(n5404) );
  OR2_X1 U6548 ( .A1(n5464), .A2(n10438), .ZN(n5393) );
  AND2_X1 U6549 ( .A1(n7399), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5027) );
  AND2_X1 U6550 ( .A1(n6742), .A2(n6741), .ZN(n5028) );
  INV_X1 U6551 ( .A(n9146), .ZN(n6073) );
  OR2_X1 U6552 ( .A1(n7659), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5029) );
  INV_X1 U6553 ( .A(n10316), .ZN(n5173) );
  AND3_X1 U6554 ( .A1(n6007), .A2(n6006), .A3(n6005), .ZN(n5030) );
  AND3_X1 U6555 ( .A1(n7019), .A2(n7017), .A3(n5854), .ZN(n5032) );
  INV_X1 U6556 ( .A(n7371), .ZN(n7174) );
  XOR2_X1 U6557 ( .A(n7375), .B(n4944), .Z(n5033) );
  AND2_X1 U6558 ( .A1(n5256), .A2(n5255), .ZN(n5034) );
  OR2_X1 U6559 ( .A1(n6698), .A2(n6697), .ZN(n5035) );
  OR2_X1 U6560 ( .A1(n7759), .A2(n7185), .ZN(n5036) );
  INV_X1 U6561 ( .A(n9192), .ZN(n6082) );
  INV_X1 U6562 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5219) );
  AND2_X1 U6563 ( .A1(n5250), .A2(n5249), .ZN(n5039) );
  AND2_X1 U6564 ( .A1(n5267), .A2(n5266), .ZN(n5040) );
  INV_X1 U6565 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6089) );
  OR2_X1 U6566 ( .A1(n9209), .A2(n7312), .ZN(n5041) );
  INV_X1 U6567 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5055) );
  OR2_X1 U6568 ( .A1(n7223), .A2(n7222), .ZN(n5042) );
  INV_X1 U6569 ( .A(n7219), .ZN(n8121) );
  XNOR2_X1 U6570 ( .A(n8126), .B(n9121), .ZN(n7219) );
  AND3_X1 U6571 ( .A1(n10001), .A2(n5673), .A3(n5672), .ZN(n5043) );
  OR2_X1 U6572 ( .A1(n10106), .A2(n10020), .ZN(n5044) );
  INV_X1 U6573 ( .A(n6570), .ZN(n6571) );
  OR2_X1 U6574 ( .A1(n6570), .A2(n9417), .ZN(n6539) );
  NAND2_X1 U6575 ( .A1(n7780), .A2(n10494), .ZN(n9438) );
  INV_X1 U6576 ( .A(n9438), .ZN(n6568) );
  AND3_X1 U6577 ( .A1(n6693), .A2(n6692), .A3(n4390), .ZN(n5046) );
  INV_X1 U6578 ( .A(n7139), .ZN(n9938) );
  AND2_X1 U6579 ( .A1(n9089), .A2(n6707), .ZN(n5047) );
  AND3_X1 U6580 ( .A1(n8884), .A2(n9772), .A3(n8883), .ZN(n5048) );
  AND2_X1 U6581 ( .A1(n8299), .A2(n5042), .ZN(n7224) );
  NAND2_X1 U6582 ( .A1(n6539), .A2(n7339), .ZN(n7244) );
  NOR2_X1 U6583 ( .A1(n7244), .A2(n7251), .ZN(n7245) );
  INV_X1 U6584 ( .A(n7271), .ZN(n7272) );
  INV_X1 U6585 ( .A(n9946), .ZN(n5702) );
  NOR2_X1 U6586 ( .A1(n7311), .A2(n7339), .ZN(n7312) );
  INV_X1 U6587 ( .A(n7320), .ZN(n7321) );
  NOR2_X1 U6588 ( .A1(n7322), .A2(n7321), .ZN(n7323) );
  NAND2_X1 U6589 ( .A1(n7213), .A2(n6527), .ZN(n6530) );
  OR2_X1 U6590 ( .A1(n9087), .A2(n9001), .ZN(n6707) );
  NAND2_X1 U6591 ( .A1(n6547), .A2(n4518), .ZN(n6548) );
  INV_X1 U6592 ( .A(n9203), .ZN(n6468) );
  INV_X1 U6593 ( .A(n8439), .ZN(n8012) );
  INV_X1 U6594 ( .A(SI_6_), .ZN(n5228) );
  INV_X1 U6595 ( .A(n6703), .ZN(n6704) );
  AND2_X1 U6596 ( .A1(n6362), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6080) );
  INV_X1 U6597 ( .A(n6460), .ZN(n6458) );
  INV_X1 U6598 ( .A(n7045), .ZN(n7047) );
  AND2_X1 U6599 ( .A1(n5634), .A2(n5290), .ZN(n5649) );
  INV_X1 U6600 ( .A(SI_13_), .ZN(n6990) );
  NOR2_X1 U6601 ( .A1(n6694), .A2(n5046), .ZN(n6695) );
  AND2_X1 U6602 ( .A1(n9013), .A2(n6672), .ZN(n6673) );
  INV_X1 U6603 ( .A(n6600), .ZN(n6202) );
  NAND2_X1 U6604 ( .A1(n5033), .A2(n7998), .ZN(n7376) );
  NOR2_X1 U6605 ( .A1(n6044), .A2(n9459), .ZN(n6045) );
  AND2_X1 U6606 ( .A1(n7550), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6047) );
  AND2_X1 U6607 ( .A1(n6267), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6050) );
  AOI21_X1 U6608 ( .B1(n7841), .B2(n7837), .A(n6200), .ZN(n6201) );
  INV_X1 U6609 ( .A(n7350), .ZN(n9311) );
  NAND2_X1 U6610 ( .A1(n9708), .A2(n8774), .ZN(n8780) );
  INV_X1 U6611 ( .A(n7123), .ZN(n7127) );
  AOI22_X1 U6612 ( .A1(n10092), .A2(n10068), .B1(n10011), .B2(n4807), .ZN(
        n8950) );
  INV_X1 U6613 ( .A(n5632), .ZN(n5633) );
  NAND2_X1 U6614 ( .A1(n5264), .A2(n6990), .ZN(n5267) );
  INV_X1 U6615 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5080) );
  INV_X1 U6616 ( .A(n6700), .ZN(n6701) );
  MUX2_X1 U6617 ( .A(n6593), .B(n6594), .S(n10463), .Z(n7768) );
  INV_X1 U6618 ( .A(n9252), .ZN(n9039) );
  INV_X1 U6619 ( .A(n9282), .ZN(n9070) );
  INV_X1 U6620 ( .A(n9102), .ZN(n9095) );
  OR2_X1 U6621 ( .A1(n6258), .A2(n6170), .ZN(n6174) );
  INV_X1 U6622 ( .A(n7568), .ZN(n6132) );
  NAND2_X1 U6623 ( .A1(n8482), .A2(n8481), .ZN(n8480) );
  INV_X1 U6624 ( .A(n7365), .ZN(n9321) );
  INV_X1 U6625 ( .A(n8680), .ZN(n6544) );
  NAND2_X1 U6626 ( .A1(n4476), .A2(n8220), .ZN(n6292) );
  AND3_X2 U6627 ( .A1(n6187), .A2(n6186), .A3(n6185), .ZN(n6586) );
  INV_X1 U6628 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6760) );
  AND2_X1 U6629 ( .A1(n7279), .A2(n7287), .ZN(n9352) );
  OR2_X1 U6630 ( .A1(n7187), .A2(n6733), .ZN(n10507) );
  OR3_X1 U6631 ( .A1(n6721), .A2(n6735), .A3(n10472), .ZN(n6759) );
  NAND2_X1 U6632 ( .A1(n6085), .A2(n6097), .ZN(n6093) );
  OR2_X1 U6633 ( .A1(n5464), .A2(n10442), .ZN(n5426) );
  OR2_X1 U6634 ( .A1(n5181), .A2(n5180), .ZN(n10339) );
  NAND2_X1 U6635 ( .A1(n5893), .A2(n7049), .ZN(n8935) );
  INV_X1 U6636 ( .A(n9919), .ZN(n9887) );
  OR2_X1 U6637 ( .A1(n10156), .A2(n8789), .ZN(n5860) );
  AND2_X1 U6638 ( .A1(n5910), .A2(n7023), .ZN(n10064) );
  INV_X1 U6639 ( .A(n10400), .ZN(n10428) );
  AND2_X1 U6640 ( .A1(n7017), .A2(n5866), .ZN(n8384) );
  AND2_X1 U6641 ( .A1(n7722), .A2(n7721), .ZN(n10090) );
  NAND2_X1 U6642 ( .A1(n5313), .A2(n5312), .ZN(n5720) );
  XNOR2_X1 U6643 ( .A(n5269), .B(SI_14_), .ZN(n5522) );
  INV_X1 U6644 ( .A(n5460), .ZN(n5461) );
  AND2_X1 U6645 ( .A1(n8615), .A2(n9444), .ZN(n9092) );
  INV_X1 U6646 ( .A(n9023), .ZN(n9108) );
  OR2_X1 U6647 ( .A1(n6258), .A2(n6219), .ZN(n6220) );
  INV_X1 U6648 ( .A(n9196), .ZN(n9169) );
  AND2_X1 U6649 ( .A1(n6149), .A2(n6128), .ZN(n9163) );
  OAI21_X1 U6650 ( .B1(n9190), .B2(n10270), .A(n8978), .ZN(n6146) );
  XNOR2_X1 U6651 ( .A(n9508), .B(n9114), .ZN(n9250) );
  INV_X1 U6652 ( .A(n9419), .ZN(n9444) );
  INV_X1 U6653 ( .A(n10464), .ZN(n9469) );
  AND2_X1 U6654 ( .A1(n9425), .A2(n9594), .ZN(n9579) );
  AND2_X1 U6655 ( .A1(n4384), .A2(n6521), .ZN(n9552) );
  INV_X1 U6656 ( .A(n9579), .ZN(n10512) );
  AND2_X1 U6657 ( .A1(n6500), .A2(n6516), .ZN(n10471) );
  AND2_X1 U6658 ( .A1(n6071), .A2(n6070), .ZN(n6326) );
  XNOR2_X1 U6659 ( .A(n6046), .B(P2_IR_REG_5__SCAN_IN), .ZN(n7550) );
  INV_X1 U6660 ( .A(n9782), .ZN(n9713) );
  OR2_X1 U6661 ( .A1(n5464), .A2(n10448), .ZN(n5473) );
  XNOR2_X1 U6662 ( .A(n5174), .B(n5173), .ZN(n10321) );
  AND2_X1 U6663 ( .A1(n5179), .A2(n5178), .ZN(n10348) );
  NAND2_X1 U6664 ( .A1(n9849), .A2(n5858), .ZN(n9869) );
  AND2_X1 U6665 ( .A1(n7055), .A2(n7690), .ZN(n10011) );
  OR2_X1 U6666 ( .A1(n7971), .A2(n7155), .ZN(n10413) );
  AOI21_X1 U6667 ( .B1(n10100), .B2(n10099), .A(n10098), .ZN(n10104) );
  OR2_X1 U6668 ( .A1(n7965), .A2(n7964), .ZN(n7976) );
  AND2_X1 U6669 ( .A1(n7068), .A2(n7067), .ZN(n10355) );
  AND2_X1 U6670 ( .A1(n5151), .A2(n5150), .ZN(n7896) );
  INV_X1 U6671 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5116) );
  AND2_X1 U6672 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10253), .ZN(n10558) );
  OAI21_X1 U6673 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10532), .ZN(n10567) );
  INV_X1 U6674 ( .A(n9190), .ZN(n9174) );
  INV_X1 U6675 ( .A(n9103), .ZN(n9072) );
  AND2_X1 U6676 ( .A1(n6723), .A2(n9290), .ZN(n9023) );
  NAND2_X1 U6677 ( .A1(n6734), .A2(n6729), .ZN(n9110) );
  INV_X1 U6678 ( .A(n9163), .ZN(n9184) );
  OR2_X1 U6679 ( .A1(n6129), .A2(n6749), .ZN(n9196) );
  XNOR2_X1 U6680 ( .A(n8906), .B(n8908), .ZN(n9486) );
  AND2_X1 U6681 ( .A1(n9316), .A2(n9315), .ZN(n9533) );
  INV_X2 U6682 ( .A(n9457), .ZN(n10461) );
  OR2_X1 U6683 ( .A1(n10461), .A2(n6524), .ZN(n9411) );
  INV_X1 U6684 ( .A(n9457), .ZN(n10470) );
  INV_X1 U6685 ( .A(n10526), .ZN(n10523) );
  INV_X1 U6686 ( .A(n10516), .ZN(n10514) );
  AND2_X2 U6687 ( .A1(n7676), .A2(n7674), .ZN(n10516) );
  NOR2_X1 U6688 ( .A1(n10472), .A2(n10471), .ZN(n10481) );
  INV_X1 U6689 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7483) );
  INV_X1 U6690 ( .A(n7150), .ZN(n9639) );
  INV_X1 U6691 ( .A(n7153), .ZN(n8934) );
  AND2_X1 U6692 ( .A1(n7818), .A2(n7817), .ZN(n9782) );
  INV_X1 U6693 ( .A(n10061), .ZN(n10186) );
  OR2_X1 U6694 ( .A1(n7628), .A2(n7618), .ZN(n9760) );
  INV_X1 U6695 ( .A(n9784), .ZN(n9771) );
  INV_X1 U6696 ( .A(n9634), .ZN(n9790) );
  INV_X1 U6697 ( .A(n8789), .ZN(n10003) );
  INV_X1 U6698 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10245) );
  INV_X1 U6699 ( .A(n10348), .ZN(n10305) );
  AOI21_X1 U6700 ( .B1(n5194), .B2(n8059), .A(n5193), .ZN(n5195) );
  NAND2_X1 U6701 ( .A1(n4448), .A2(n10030), .ZN(n7161) );
  NAND2_X1 U6702 ( .A1(n10078), .A2(n7152), .ZN(n10009) );
  INV_X1 U6703 ( .A(n10455), .ZN(n10452) );
  OR3_X1 U6704 ( .A1(n10190), .A2(n10189), .A3(n10188), .ZN(n10221) );
  INV_X1 U6705 ( .A(n10437), .ZN(n10435) );
  INV_X1 U6706 ( .A(n10367), .ZN(n10364) );
  INV_X1 U6707 ( .A(n9990), .ZN(n8059) );
  INV_X1 U6708 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7682) );
  INV_X1 U6709 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n7427) );
  NOR2_X1 U6710 ( .A1(n10563), .A2(n10565), .ZN(n10562) );
  INV_X1 U6711 ( .A(n10561), .ZN(n10564) );
  OAI21_X1 U6712 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10544), .ZN(n10542) );
  NAND2_X1 U6713 ( .A1(n6154), .A2(n6155), .ZN(P2_U3264) );
  NAND2_X1 U6714 ( .A1(n5196), .A2(n5195), .ZN(P1_U3260) );
  NAND2_X1 U6715 ( .A1(n5118), .A2(n5049), .ZN(n5110) );
  INV_X1 U6716 ( .A(n5110), .ZN(n5051) );
  AND2_X2 U6717 ( .A1(n5138), .A2(n5080), .ZN(n5144) );
  NOR2_X2 U6718 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5063) );
  NOR2_X1 U6719 ( .A1(n5076), .A2(n5077), .ZN(n5056) );
  XNOR2_X1 U6720 ( .A(n5143), .B(P1_IR_REG_25__SCAN_IN), .ZN(n5057) );
  NAND2_X1 U6721 ( .A1(n5144), .A2(n5081), .ZN(n5059) );
  INV_X1 U6722 ( .A(n7812), .ZN(n7624) );
  NAND2_X1 U6723 ( .A1(n5059), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5060) );
  XNOR2_X1 U6724 ( .A(n5060), .B(n4758), .ZN(n7811) );
  NAND2_X1 U6725 ( .A1(n7624), .A2(n7811), .ZN(n7383) );
  INV_X1 U6726 ( .A(n5102), .ZN(n5061) );
  NAND4_X1 U6727 ( .A1(n5062), .A2(n5061), .A3(n5080), .A4(n5079), .ZN(n5065)
         );
  NAND3_X1 U6728 ( .A1(n5063), .A2(n5090), .A3(n6914), .ZN(n5064) );
  NOR2_X1 U6729 ( .A1(n5065), .A2(n5064), .ZN(n5066) );
  NAND2_X2 U6730 ( .A1(n5185), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5953) );
  NAND2_X1 U6731 ( .A1(n5953), .A2(n5954), .ZN(n5068) );
  NAND2_X2 U6732 ( .A1(n5068), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5073) );
  INV_X1 U6733 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5072) );
  NAND2_X1 U6734 ( .A1(n5073), .A2(n5072), .ZN(n5069) );
  NAND2_X1 U6735 ( .A1(n5069), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5071) );
  INV_X1 U6736 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5070) );
  XNOR2_X2 U6737 ( .A(n5071), .B(n5070), .ZN(n8250) );
  XNOR2_X2 U6738 ( .A(n5073), .B(n5072), .ZN(n5946) );
  NAND2_X1 U6739 ( .A1(n7051), .A2(n4495), .ZN(n7617) );
  INV_X1 U6740 ( .A(n7811), .ZN(n5074) );
  OR2_X1 U6741 ( .A1(n7617), .A2(n5074), .ZN(n5075) );
  NAND2_X1 U6742 ( .A1(n7383), .A2(n5075), .ZN(n5181) );
  INV_X1 U6743 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5078) );
  NAND2_X1 U6744 ( .A1(n5360), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5082) );
  INV_X1 U6745 ( .A(n5360), .ZN(n5084) );
  INV_X1 U6746 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5083) );
  NAND2_X1 U6747 ( .A1(n5086), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5087) );
  OR2_X1 U6748 ( .A1(n5181), .A2(n5655), .ZN(n5089) );
  NAND2_X1 U6749 ( .A1(n5089), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  NAND2_X1 U6750 ( .A1(n5144), .A2(n5090), .ZN(n5101) );
  INV_X1 U6751 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5092) );
  INV_X1 U6752 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5091) );
  NAND4_X1 U6753 ( .A1(n5092), .A2(n5108), .A3(n5148), .A4(n5091), .ZN(n5093)
         );
  OR2_X1 U6754 ( .A1(n5101), .A2(n5093), .ZN(n5099) );
  OAI21_X1 U6755 ( .B1(n5099), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5096) );
  INV_X1 U6756 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U6757 ( .A1(n5096), .A2(n5095), .ZN(n5098) );
  NAND2_X1 U6758 ( .A1(n5098), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5094) );
  XNOR2_X1 U6759 ( .A(n5094), .B(P1_IR_REG_18__SCAN_IN), .ZN(n5637) );
  INV_X1 U6760 ( .A(n5637), .ZN(n9827) );
  INV_X1 U6761 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n5644) );
  AOI22_X1 U6762 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n9827), .B1(n5637), .B2(
        n5644), .ZN(n9825) );
  OR2_X1 U6763 ( .A1(n5096), .A2(n5095), .ZN(n5097) );
  NAND2_X1 U6764 ( .A1(n5098), .A2(n5097), .ZN(n10338) );
  INV_X1 U6765 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n5628) );
  XNOR2_X1 U6766 ( .A(n10338), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n10346) );
  NAND2_X1 U6767 ( .A1(n5099), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5100) );
  XNOR2_X1 U6768 ( .A(n5100), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7705) );
  INV_X1 U6769 ( .A(n7705), .ZN(n10326) );
  INV_X1 U6770 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n5158) );
  XOR2_X1 U6771 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n7705), .Z(n10330) );
  NAND2_X1 U6772 ( .A1(n5101), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5149) );
  NAND2_X1 U6773 ( .A1(n5102), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5103) );
  NAND2_X1 U6774 ( .A1(n5149), .A2(n5103), .ZN(n5105) );
  OR2_X1 U6775 ( .A1(n5105), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5107) );
  NAND2_X1 U6776 ( .A1(n5107), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5104) );
  XNOR2_X1 U6777 ( .A(n5104), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10316) );
  NAND2_X1 U6778 ( .A1(n5105), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5106) );
  INV_X1 U6779 ( .A(n5525), .ZN(n8425) );
  INV_X1 U6780 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n5155) );
  INV_X1 U6781 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6940) );
  NAND2_X1 U6782 ( .A1(n5149), .A2(n5148), .ZN(n5151) );
  NAND2_X1 U6783 ( .A1(n5151), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5109) );
  XNOR2_X1 U6784 ( .A(n5109), .B(n5108), .ZN(n8140) );
  NOR2_X1 U6785 ( .A1(n5110), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5114) );
  INV_X1 U6786 ( .A(n5114), .ZN(n5111) );
  NAND2_X1 U6787 ( .A1(n5111), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5112) );
  MUX2_X1 U6788 ( .A(n5112), .B(P1_IR_REG_31__SCAN_IN), .S(n5113), .Z(n5115)
         );
  NAND2_X1 U6789 ( .A1(n5114), .A2(n5113), .ZN(n5126) );
  NAND2_X1 U6790 ( .A1(n5115), .A2(n5126), .ZN(n7451) );
  INV_X1 U6791 ( .A(n7451), .ZN(n5454) );
  NAND2_X1 U6792 ( .A1(n5110), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5117) );
  XNOR2_X1 U6793 ( .A(n5117), .B(n5116), .ZN(n7701) );
  INV_X1 U6794 ( .A(n7701), .ZN(n5163) );
  INV_X1 U6795 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5119) );
  NAND2_X1 U6796 ( .A1(n5122), .A2(n5119), .ZN(n5120) );
  NAND2_X1 U6797 ( .A1(n5120), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5121) );
  XNOR2_X1 U6798 ( .A(n5121), .B(P1_IR_REG_3__SCAN_IN), .ZN(n7390) );
  INV_X1 U6799 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10440) );
  NAND2_X1 U6800 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5123) );
  XNOR2_X1 U6801 ( .A(n5123), .B(P1_IR_REG_1__SCAN_IN), .ZN(n7396) );
  INV_X1 U6802 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10438) );
  MUX2_X1 U6803 ( .A(n10438), .B(P1_REG1_REG_1__SCAN_IN), .S(n7396), .Z(n7442)
         );
  INV_X1 U6804 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5124) );
  INV_X1 U6805 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10289) );
  NOR3_X1 U6806 ( .A1(n7442), .A2(n5124), .A3(n10289), .ZN(n7440) );
  AOI21_X1 U6807 ( .B1(n7396), .B2(P1_REG1_REG_1__SCAN_IN), .A(n7440), .ZN(
        n10303) );
  MUX2_X1 U6808 ( .A(n10440), .B(P1_REG1_REG_2__SCAN_IN), .S(n7399), .Z(n10302) );
  NOR2_X1 U6809 ( .A1(n10303), .A2(n10302), .ZN(n10301) );
  AOI21_X1 U6810 ( .B1(n7399), .B2(P1_REG1_REG_2__SCAN_IN), .A(n10301), .ZN(
        n10282) );
  INV_X1 U6811 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10442) );
  MUX2_X1 U6812 ( .A(n10442), .B(P1_REG1_REG_3__SCAN_IN), .S(n7390), .Z(n10281) );
  NOR2_X1 U6813 ( .A1(n10282), .A2(n10281), .ZN(n10280) );
  AOI21_X1 U6814 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n7390), .A(n10280), .ZN(
        n7697) );
  INV_X1 U6815 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10444) );
  MUX2_X1 U6816 ( .A(n10444), .B(P1_REG1_REG_4__SCAN_IN), .S(n7701), .Z(n7696)
         );
  NAND2_X1 U6817 ( .A1(n7697), .A2(n7696), .ZN(n7695) );
  OAI21_X1 U6818 ( .B1(n5163), .B2(P1_REG1_REG_4__SCAN_IN), .A(n7695), .ZN(
        n7450) );
  INV_X1 U6819 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10446) );
  MUX2_X1 U6820 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10446), .S(n7451), .Z(n7449)
         );
  NOR2_X1 U6821 ( .A1(n7450), .A2(n7449), .ZN(n7448) );
  AOI21_X1 U6822 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n5454), .A(n7448), .ZN(
        n9812) );
  INV_X1 U6823 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10448) );
  NAND2_X1 U6824 ( .A1(n5126), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5125) );
  XNOR2_X1 U6825 ( .A(n5125), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9818) );
  MUX2_X1 U6826 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10448), .S(n9818), .Z(n9811)
         );
  NOR2_X1 U6827 ( .A1(n9818), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7490) );
  INV_X1 U6828 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10450) );
  INV_X1 U6829 ( .A(n5126), .ZN(n5128) );
  NAND2_X1 U6830 ( .A1(n5128), .A2(n5127), .ZN(n5130) );
  NAND2_X1 U6831 ( .A1(n5130), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5129) );
  XNOR2_X1 U6832 ( .A(n5129), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7488) );
  MUX2_X1 U6833 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n10450), .S(n7488), .Z(n7491)
         );
  OAI21_X1 U6834 ( .B1(n5130), .B2(P1_IR_REG_7__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5131) );
  XNOR2_X1 U6835 ( .A(n5131), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7462) );
  NAND2_X1 U6836 ( .A1(n7462), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7522) );
  OR2_X1 U6837 ( .A1(n7462), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5132) );
  OR2_X1 U6838 ( .A1(n7488), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7463) );
  MUX2_X1 U6839 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5133), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n5135) );
  INV_X1 U6840 ( .A(n5138), .ZN(n5134) );
  NAND2_X1 U6841 ( .A1(n5135), .A2(n5134), .ZN(n7413) );
  INV_X1 U6842 ( .A(n7413), .ZN(n7527) );
  NAND2_X1 U6843 ( .A1(n7527), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5137) );
  INV_X1 U6844 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5136) );
  NAND2_X1 U6845 ( .A1(n7413), .A2(n5136), .ZN(n7504) );
  AND2_X1 U6846 ( .A1(n5137), .A2(n7504), .ZN(n7521) );
  NOR2_X1 U6847 ( .A1(n5138), .A2(n5143), .ZN(n5139) );
  MUX2_X1 U6848 ( .A(n5143), .B(n5139), .S(P1_IR_REG_10__SCAN_IN), .Z(n5140)
         );
  NOR2_X1 U6849 ( .A1(n5140), .A2(n5144), .ZN(n7425) );
  OR2_X1 U6850 ( .A1(n7425), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5142) );
  NAND2_X1 U6851 ( .A1(n7425), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5141) );
  NAND2_X1 U6852 ( .A1(n5142), .A2(n5141), .ZN(n7503) );
  AOI21_X1 U6853 ( .B1(n7520), .B2(n7504), .A(n7503), .ZN(n7655) );
  INV_X1 U6854 ( .A(n5142), .ZN(n7654) );
  OR2_X1 U6855 ( .A1(n5144), .A2(n5143), .ZN(n5145) );
  XNOR2_X1 U6856 ( .A(n5145), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7659) );
  INV_X1 U6857 ( .A(n7659), .ZN(n7434) );
  INV_X1 U6858 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n5146) );
  NAND2_X1 U6859 ( .A1(n7434), .A2(n5146), .ZN(n7891) );
  NAND2_X1 U6860 ( .A1(n7659), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5147) );
  AND2_X1 U6861 ( .A1(n7891), .A2(n5147), .ZN(n7653) );
  OR2_X1 U6862 ( .A1(n5149), .A2(n5148), .ZN(n5150) );
  INV_X1 U6863 ( .A(n7896), .ZN(n7478) );
  INV_X1 U6864 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5152) );
  NAND2_X1 U6865 ( .A1(n7478), .A2(n5152), .ZN(n5154) );
  NAND2_X1 U6866 ( .A1(n7896), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5153) );
  NAND2_X1 U6867 ( .A1(n5154), .A2(n5153), .ZN(n7890) );
  XOR2_X1 U6868 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n8140), .Z(n8135) );
  AOI21_X1 U6869 ( .B1(n6940), .B2(n8140), .A(n8134), .ZN(n8428) );
  AOI22_X1 U6870 ( .A1(n5525), .A2(n5155), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n8425), .ZN(n8427) );
  NOR2_X1 U6871 ( .A1(n8428), .A2(n8427), .ZN(n8426) );
  NAND2_X1 U6872 ( .A1(n10316), .A2(n5156), .ZN(n5157) );
  NAND2_X1 U6873 ( .A1(n10330), .A2(n10331), .ZN(n10329) );
  OAI21_X1 U6874 ( .B1(n10326), .B2(n5158), .A(n10329), .ZN(n10345) );
  NAND2_X1 U6875 ( .A1(n10346), .A2(n10345), .ZN(n10343) );
  OAI21_X1 U6876 ( .B1(n10338), .B2(n5628), .A(n10343), .ZN(n9824) );
  NOR2_X1 U6877 ( .A1(n7684), .A2(P1_U3084), .ZN(n8697) );
  NAND2_X1 U6878 ( .A1(n8697), .A2(n7686), .ZN(n5160) );
  OR2_X1 U6879 ( .A1(n5181), .A2(n5160), .ZN(n10300) );
  INV_X1 U6880 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n6892) );
  XNOR2_X1 U6881 ( .A(n9827), .B(P1_REG2_REG_18__SCAN_IN), .ZN(n9831) );
  INV_X1 U6882 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n6923) );
  MUX2_X1 U6883 ( .A(n6923), .B(P1_REG2_REG_17__SCAN_IN), .S(n10338), .Z(
        n10349) );
  INV_X1 U6884 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n5176) );
  MUX2_X1 U6885 ( .A(P1_REG2_REG_16__SCAN_IN), .B(n5176), .S(n7705), .Z(n10333) );
  INV_X1 U6886 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6829) );
  INV_X1 U6887 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5161) );
  MUX2_X1 U6888 ( .A(n5161), .B(P1_REG2_REG_2__SCAN_IN), .S(n7399), .Z(n10307)
         );
  INV_X1 U6889 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7944) );
  MUX2_X1 U6890 ( .A(n7944), .B(P1_REG2_REG_3__SCAN_IN), .S(n7390), .Z(n10277)
         );
  INV_X1 U6891 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5162) );
  MUX2_X1 U6892 ( .A(n5162), .B(P1_REG2_REG_4__SCAN_IN), .S(n7701), .Z(n7694)
         );
  NOR2_X1 U6893 ( .A1(n5163), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7452) );
  INV_X1 U6894 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n8063) );
  MUX2_X1 U6895 ( .A(n8063), .B(P1_REG2_REG_5__SCAN_IN), .S(n7451), .Z(n7453)
         );
  OAI21_X1 U6896 ( .B1(n5454), .B2(P1_REG2_REG_5__SCAN_IN), .A(n7455), .ZN(
        n9815) );
  INV_X1 U6897 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5164) );
  MUX2_X1 U6898 ( .A(n5164), .B(P1_REG2_REG_6__SCAN_IN), .S(n9818), .Z(n9814)
         );
  INV_X1 U6899 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n5166) );
  MUX2_X1 U6900 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n5166), .S(n7488), .Z(n7484)
         );
  NOR2_X1 U6901 ( .A1(n7488), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7470) );
  INV_X1 U6902 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5167) );
  MUX2_X1 U6903 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n5167), .S(n7462), .Z(n7471)
         );
  OAI21_X1 U6904 ( .B1(n7462), .B2(P1_REG2_REG_8__SCAN_IN), .A(n7469), .ZN(
        n7519) );
  INV_X1 U6905 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n5168) );
  MUX2_X1 U6906 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n5168), .S(n7413), .Z(n7518)
         );
  NAND2_X1 U6907 ( .A1(n7527), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7500) );
  INV_X1 U6908 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6852) );
  MUX2_X1 U6909 ( .A(n6852), .B(P1_REG2_REG_10__SCAN_IN), .S(n7425), .Z(n7499)
         );
  INV_X1 U6910 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n5169) );
  MUX2_X1 U6911 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n5169), .S(n7659), .Z(n7651)
         );
  INV_X1 U6912 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n5170) );
  MUX2_X1 U6913 ( .A(n5170), .B(P1_REG2_REG_12__SCAN_IN), .S(n7896), .Z(n7888)
         );
  MUX2_X1 U6914 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n6829), .S(n8140), .Z(n8137)
         );
  NOR2_X1 U6915 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(n8424), .ZN(n8423) );
  NOR2_X1 U6916 ( .A1(n5525), .A2(n5171), .ZN(n5172) );
  NAND2_X1 U6917 ( .A1(n10316), .A2(n5174), .ZN(n5175) );
  NAND2_X1 U6918 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n10321), .ZN(n10320) );
  NAND2_X1 U6919 ( .A1(n5175), .A2(n10320), .ZN(n10334) );
  NAND2_X1 U6920 ( .A1(n10333), .A2(n10334), .ZN(n10332) );
  NAND2_X1 U6921 ( .A1(n10349), .A2(n10350), .ZN(n10347) );
  OAI21_X1 U6922 ( .B1(n10338), .B2(n6923), .A(n10347), .ZN(n9830) );
  NAND2_X1 U6923 ( .A1(n9831), .A2(n9830), .ZN(n9829) );
  OAI21_X1 U6924 ( .B1(n9827), .B2(n6892), .A(n9829), .ZN(n5177) );
  XNOR2_X1 U6925 ( .A(n5177), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n5190) );
  INV_X1 U6926 ( .A(n5181), .ZN(n5179) );
  INV_X1 U6927 ( .A(n7686), .ZN(n10288) );
  AND2_X1 U6928 ( .A1(n8697), .A2(n10288), .ZN(n5178) );
  NAND2_X1 U6929 ( .A1(n5190), .A2(n10348), .ZN(n5182) );
  NOR2_X1 U6930 ( .A1(n7686), .A2(P1_U3084), .ZN(n8692) );
  NAND2_X1 U6931 ( .A1(n8692), .A2(n7684), .ZN(n5180) );
  OAI211_X1 U6932 ( .C1(n5188), .C2(n10300), .A(n5182), .B(n10339), .ZN(n5187)
         );
  NAND2_X1 U6933 ( .A1(n5183), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5184) );
  MUX2_X1 U6934 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5184), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n5186) );
  NAND2_X1 U6935 ( .A1(n5187), .A2(n9990), .ZN(n5196) );
  INV_X1 U6936 ( .A(n10300), .ZN(n10344) );
  OAI21_X1 U6937 ( .B1(n5190), .B2(n10305), .A(n5189), .ZN(n5194) );
  INV_X1 U6938 ( .A(n7383), .ZN(n5191) );
  NOR2_X2 U6939 ( .A1(P1_U3083), .A2(n5191), .ZN(n10342) );
  AND2_X1 U6940 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9673) );
  AOI21_X1 U6941 ( .B1(n10342), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n9673), .ZN(
        n5192) );
  INV_X1 U6942 ( .A(n5192), .ZN(n5193) );
  INV_X1 U6943 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n7385) );
  NAND2_X1 U6944 ( .A1(n4382), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5199) );
  INV_X1 U6945 ( .A(SI_2_), .ZN(n5198) );
  OAI211_X1 U6946 ( .C1(n5398), .C2(n7385), .A(n5199), .B(n5198), .ZN(n5210)
         );
  NOR2_X1 U6947 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(SI_1_), .ZN(n5202) );
  AND2_X1 U6948 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5395) );
  INV_X1 U6949 ( .A(n5395), .ZN(n5201) );
  NAND2_X1 U6950 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(SI_1_), .ZN(n5200) );
  OAI21_X1 U6951 ( .B1(n5202), .B2(n5201), .A(n5200), .ZN(n5203) );
  NAND2_X1 U6952 ( .A1(n4382), .A2(n5203), .ZN(n5209) );
  NOR2_X1 U6953 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5206) );
  AND2_X1 U6954 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5396) );
  INV_X1 U6955 ( .A(n5396), .ZN(n5205) );
  NAND2_X1 U6956 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5204) );
  OAI21_X1 U6957 ( .B1(n5206), .B2(n5205), .A(n5204), .ZN(n5207) );
  NAND2_X1 U6958 ( .A1(n5225), .A2(n5207), .ZN(n5208) );
  NAND2_X1 U6959 ( .A1(n5209), .A2(n5208), .ZN(n5419) );
  NAND2_X1 U6960 ( .A1(n5210), .A2(n5419), .ZN(n5213) );
  INV_X1 U6961 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7400) );
  NAND2_X1 U6962 ( .A1(n7389), .A2(n7400), .ZN(n5211) );
  OAI211_X1 U6963 ( .C1(n7389), .C2(P1_DATAO_REG_2__SCAN_IN), .A(n5211), .B(
        SI_2_), .ZN(n5212) );
  NAND2_X1 U6964 ( .A1(n5213), .A2(n5212), .ZN(n5428) );
  INV_X1 U6965 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7392) );
  INV_X1 U6966 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n7387) );
  NAND2_X1 U6967 ( .A1(n5428), .A2(n5429), .ZN(n5217) );
  INV_X1 U6968 ( .A(n5214), .ZN(n5215) );
  NAND2_X1 U6969 ( .A1(n5215), .A2(SI_3_), .ZN(n5216) );
  INV_X1 U6970 ( .A(n5440), .ZN(n5220) );
  NAND2_X1 U6971 ( .A1(n5439), .A2(n5220), .ZN(n5223) );
  NAND2_X1 U6972 ( .A1(n5221), .A2(SI_4_), .ZN(n5222) );
  MUX2_X1 U6973 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n7389), .Z(n5231) );
  NAND2_X1 U6974 ( .A1(n5453), .A2(n5224), .ZN(n5459) );
  INV_X1 U6975 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n5226) );
  INV_X1 U6976 ( .A(SI_7_), .ZN(n5229) );
  NAND2_X1 U6977 ( .A1(n5230), .A2(n5229), .ZN(n5238) );
  NAND2_X1 U6978 ( .A1(n5460), .A2(n5238), .ZN(n5243) );
  NAND2_X1 U6979 ( .A1(n5231), .A2(SI_5_), .ZN(n5458) );
  INV_X1 U6980 ( .A(n5458), .ZN(n5232) );
  NAND3_X1 U6981 ( .A1(n5232), .A2(n5238), .A3(n5460), .ZN(n5242) );
  INV_X1 U6982 ( .A(SI_8_), .ZN(n5233) );
  NAND2_X1 U6983 ( .A1(n5234), .A2(n5233), .ZN(n5244) );
  NAND2_X1 U6984 ( .A1(n5235), .A2(SI_8_), .ZN(n5236) );
  INV_X1 U6985 ( .A(n5503), .ZN(n5241) );
  NAND2_X1 U6986 ( .A1(n5480), .A2(SI_7_), .ZN(n5501) );
  NAND2_X1 U6987 ( .A1(n5237), .A2(SI_6_), .ZN(n5478) );
  INV_X1 U6988 ( .A(n5478), .ZN(n5239) );
  NAND2_X1 U6989 ( .A1(n5239), .A2(n5238), .ZN(n5240) );
  NAND2_X1 U6990 ( .A1(n5245), .A2(n5244), .ZN(n5513) );
  MUX2_X1 U6991 ( .A(n7412), .B(n7415), .S(n4522), .Z(n5247) );
  INV_X1 U6992 ( .A(SI_9_), .ZN(n5246) );
  INV_X1 U6993 ( .A(n5247), .ZN(n5248) );
  NAND2_X1 U6994 ( .A1(n5248), .A2(SI_9_), .ZN(n5249) );
  MUX2_X1 U6995 ( .A(n7420), .B(n7427), .S(n4382), .Z(n5253) );
  INV_X1 U6996 ( .A(n5253), .ZN(n5254) );
  NAND2_X1 U6997 ( .A1(n5254), .A2(SI_10_), .ZN(n5255) );
  MUX2_X1 U6998 ( .A(n7430), .B(n7436), .S(n4522), .Z(n5257) );
  INV_X1 U6999 ( .A(n5257), .ZN(n5258) );
  MUX2_X1 U7000 ( .A(n7477), .B(n7480), .S(n4522), .Z(n5260) );
  INV_X1 U7001 ( .A(SI_12_), .ZN(n5259) );
  INV_X1 U7002 ( .A(n5260), .ZN(n5261) );
  NAND2_X1 U7003 ( .A1(n5261), .A2(SI_12_), .ZN(n5262) );
  MUX2_X1 U7004 ( .A(n7483), .B(n7498), .S(n4522), .Z(n5264) );
  INV_X1 U7005 ( .A(n5264), .ZN(n5265) );
  NAND2_X1 U7006 ( .A1(n5265), .A2(SI_13_), .ZN(n5266) );
  MUX2_X1 U7007 ( .A(n7513), .B(n7515), .S(n4522), .Z(n5269) );
  INV_X1 U7008 ( .A(n5269), .ZN(n5270) );
  MUX2_X1 U7009 ( .A(n7680), .B(n7682), .S(n4522), .Z(n5274) );
  INV_X1 U7010 ( .A(SI_15_), .ZN(n5273) );
  INV_X1 U7011 ( .A(n5274), .ZN(n5275) );
  NAND2_X1 U7012 ( .A1(n5275), .A2(SI_15_), .ZN(n5276) );
  INV_X1 U7013 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7717) );
  INV_X1 U7014 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5278) );
  MUX2_X1 U7015 ( .A(n7717), .B(n5278), .S(n4522), .Z(n5280) );
  INV_X1 U7016 ( .A(SI_16_), .ZN(n5279) );
  NAND2_X1 U7017 ( .A1(n5280), .A2(n5279), .ZN(n5616) );
  INV_X1 U7018 ( .A(n5280), .ZN(n5281) );
  NAND2_X1 U7019 ( .A1(n5281), .A2(SI_16_), .ZN(n5282) );
  INV_X1 U7020 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7833) );
  MUX2_X1 U7021 ( .A(n7833), .B(n7835), .S(n4522), .Z(n5292) );
  INV_X1 U7022 ( .A(n5292), .ZN(n5283) );
  NAND2_X1 U7023 ( .A1(n5283), .A2(SI_17_), .ZN(n5291) );
  MUX2_X1 U7024 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4522), .Z(n5295) );
  NAND2_X1 U7025 ( .A1(n5295), .A2(SI_18_), .ZN(n5290) );
  MUX2_X1 U7026 ( .A(n7886), .B(n7884), .S(n4522), .Z(n5285) );
  INV_X1 U7027 ( .A(SI_19_), .ZN(n5284) );
  INV_X1 U7028 ( .A(n5285), .ZN(n5286) );
  NAND2_X1 U7029 ( .A1(n5286), .A2(SI_19_), .ZN(n5287) );
  INV_X1 U7030 ( .A(n5653), .ZN(n5288) );
  INV_X1 U7031 ( .A(n5290), .ZN(n5298) );
  INV_X1 U7032 ( .A(n5291), .ZN(n5294) );
  XNOR2_X1 U7033 ( .A(n5292), .B(SI_17_), .ZN(n5618) );
  XNOR2_X1 U7034 ( .A(n5295), .B(SI_18_), .ZN(n5635) );
  INV_X1 U7035 ( .A(n5635), .ZN(n5296) );
  INV_X1 U7036 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7980) );
  INV_X1 U7037 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7995) );
  MUX2_X1 U7038 ( .A(n7980), .B(n7995), .S(n4522), .Z(n5300) );
  INV_X1 U7039 ( .A(SI_20_), .ZN(n6831) );
  NAND2_X1 U7040 ( .A1(n5300), .A2(n6831), .ZN(n5303) );
  INV_X1 U7041 ( .A(n5300), .ZN(n5301) );
  NAND2_X1 U7042 ( .A1(n5301), .A2(SI_20_), .ZN(n5302) );
  INV_X1 U7043 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7997) );
  INV_X1 U7044 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8958) );
  MUX2_X1 U7045 ( .A(n7997), .B(n8958), .S(n4522), .Z(n5305) );
  INV_X1 U7046 ( .A(n5305), .ZN(n5306) );
  NAND2_X1 U7047 ( .A1(n5306), .A2(SI_21_), .ZN(n5307) );
  INV_X1 U7048 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8960) );
  INV_X1 U7049 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8251) );
  MUX2_X1 U7050 ( .A(n8960), .B(n8251), .S(n4522), .Z(n5310) );
  INV_X1 U7051 ( .A(SI_22_), .ZN(n5309) );
  INV_X1 U7052 ( .A(n5310), .ZN(n5311) );
  NAND2_X1 U7053 ( .A1(n5311), .A2(SI_22_), .ZN(n5312) );
  INV_X1 U7054 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5314) );
  INV_X1 U7055 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8334) );
  MUX2_X1 U7056 ( .A(n5314), .B(n8334), .S(n4522), .Z(n5316) );
  INV_X1 U7057 ( .A(SI_23_), .ZN(n5315) );
  NAND2_X1 U7058 ( .A1(n5316), .A2(n5315), .ZN(n5742) );
  INV_X1 U7059 ( .A(n5316), .ZN(n5317) );
  NAND2_X1 U7060 ( .A1(n5317), .A2(SI_23_), .ZN(n5318) );
  INV_X1 U7061 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8496) );
  INV_X1 U7062 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8478) );
  MUX2_X1 U7063 ( .A(n8496), .B(n8478), .S(n4522), .Z(n5322) );
  XNOR2_X1 U7064 ( .A(n5322), .B(SI_24_), .ZN(n5744) );
  INV_X1 U7065 ( .A(n5744), .ZN(n5320) );
  INV_X1 U7066 ( .A(n5742), .ZN(n5319) );
  NOR2_X1 U7067 ( .A1(n5320), .A2(n5319), .ZN(n5321) );
  NAND2_X1 U7068 ( .A1(n5743), .A2(n5321), .ZN(n5325) );
  INV_X1 U7069 ( .A(n5322), .ZN(n5323) );
  NAND2_X1 U7070 ( .A1(n5323), .A2(SI_24_), .ZN(n5324) );
  INV_X1 U7071 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8578) );
  INV_X1 U7072 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8575) );
  MUX2_X1 U7073 ( .A(n8578), .B(n8575), .S(n4522), .Z(n5327) );
  INV_X1 U7074 ( .A(SI_25_), .ZN(n5326) );
  NAND2_X1 U7075 ( .A1(n5327), .A2(n5326), .ZN(n5330) );
  INV_X1 U7076 ( .A(n5327), .ZN(n5328) );
  NAND2_X1 U7077 ( .A1(n5328), .A2(SI_25_), .ZN(n5329) );
  NAND2_X1 U7078 ( .A1(n5330), .A2(n5329), .ZN(n5755) );
  INV_X1 U7079 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8686) );
  INV_X1 U7080 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8688) );
  MUX2_X1 U7081 ( .A(n8686), .B(n8688), .S(n4522), .Z(n5332) );
  INV_X1 U7082 ( .A(SI_26_), .ZN(n5331) );
  NAND2_X1 U7083 ( .A1(n5332), .A2(n5331), .ZN(n5794) );
  INV_X1 U7084 ( .A(n5332), .ZN(n5333) );
  NAND2_X1 U7085 ( .A1(n5333), .A2(SI_26_), .ZN(n5334) );
  INV_X1 U7086 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8694) );
  INV_X1 U7087 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5335) );
  MUX2_X1 U7088 ( .A(n8694), .B(n5335), .S(n4522), .Z(n5338) );
  INV_X1 U7089 ( .A(SI_27_), .ZN(n5336) );
  NAND2_X1 U7090 ( .A1(n5338), .A2(n5336), .ZN(n5797) );
  AND2_X1 U7091 ( .A1(n5794), .A2(n5797), .ZN(n5337) );
  INV_X1 U7092 ( .A(n5338), .ZN(n5339) );
  NAND2_X1 U7093 ( .A1(n5339), .A2(SI_27_), .ZN(n5796) );
  INV_X1 U7094 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8718) );
  INV_X1 U7095 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n6917) );
  MUX2_X1 U7096 ( .A(n8718), .B(n6917), .S(n7389), .Z(n5342) );
  INV_X1 U7097 ( .A(SI_28_), .ZN(n5341) );
  NAND2_X1 U7098 ( .A1(n5342), .A2(n5341), .ZN(n5386) );
  INV_X1 U7099 ( .A(n5342), .ZN(n5343) );
  NAND2_X1 U7100 ( .A1(n5343), .A2(SI_28_), .ZN(n5344) );
  INV_X1 U7101 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10237) );
  INV_X1 U7102 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9625) );
  MUX2_X1 U7103 ( .A(n10237), .B(n9625), .S(n7388), .Z(n5347) );
  INV_X1 U7104 ( .A(n5347), .ZN(n5345) );
  NAND2_X1 U7105 ( .A1(n5345), .A2(SI_29_), .ZN(n5388) );
  MUX2_X1 U7106 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n7388), .Z(n5836) );
  INV_X1 U7107 ( .A(n5836), .ZN(n5348) );
  NAND2_X1 U7108 ( .A1(n5388), .A2(n5348), .ZN(n5356) );
  INV_X1 U7109 ( .A(SI_29_), .ZN(n5346) );
  NAND2_X1 U7110 ( .A1(n5347), .A2(n5346), .ZN(n5835) );
  INV_X1 U7111 ( .A(n5835), .ZN(n5349) );
  NAND2_X1 U7112 ( .A1(n5349), .A2(n5348), .ZN(n5352) );
  INV_X1 U7113 ( .A(n5388), .ZN(n5350) );
  NAND2_X1 U7114 ( .A1(n5350), .A2(n5836), .ZN(n5351) );
  OAI211_X1 U7115 ( .C1(n5356), .C2(n5386), .A(n5352), .B(n5351), .ZN(n5353)
         );
  INV_X1 U7116 ( .A(n5353), .ZN(n5355) );
  NAND4_X1 U7117 ( .A1(n5387), .A2(n5836), .A3(n5386), .A4(n5835), .ZN(n5354)
         );
  NAND2_X2 U7118 ( .A1(n5407), .A2(n4522), .ZN(n5524) );
  INV_X1 U7119 ( .A(n5524), .ZN(n5844) );
  NAND2_X1 U7120 ( .A1(n8953), .A2(n5844), .ZN(n5358) );
  AND2_X2 U7121 ( .A1(n5407), .A2(n7388), .ZN(n5430) );
  INV_X2 U7122 ( .A(n5535), .ZN(n5815) );
  NAND2_X1 U7123 ( .A1(n5815), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n5357) );
  INV_X1 U7124 ( .A(n5362), .ZN(n10227) );
  NAND2_X1 U7125 ( .A1(n5762), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5366) );
  NAND2_X1 U7126 ( .A1(n5803), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5365) );
  AND2_X2 U7127 ( .A1(n10235), .A2(n10234), .ZN(n5469) );
  NAND2_X1 U7128 ( .A1(n5763), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5364) );
  AND3_X1 U7129 ( .A1(n5366), .A2(n5365), .A3(n5364), .ZN(n7057) );
  INV_X1 U7130 ( .A(n7057), .ZN(n9789) );
  NAND2_X1 U7131 ( .A1(n5762), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5370) );
  NAND2_X1 U7132 ( .A1(n5803), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5369) );
  NAND2_X1 U7133 ( .A1(n5763), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5368) );
  NAND3_X1 U7134 ( .A1(n5370), .A2(n5369), .A3(n5368), .ZN(n9788) );
  NAND2_X1 U7135 ( .A1(n9789), .A2(n9788), .ZN(n5371) );
  AND2_X1 U7136 ( .A1(n10087), .A2(n5371), .ZN(n5851) );
  INV_X1 U7137 ( .A(n5851), .ZN(n5943) );
  INV_X1 U7138 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5528) );
  INV_X1 U7139 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9714) );
  INV_X1 U7140 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5658) );
  INV_X1 U7141 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5710) );
  INV_X1 U7142 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9725) );
  INV_X1 U7143 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5759) );
  INV_X1 U7144 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9633) );
  INV_X1 U7145 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8880) );
  INV_X1 U7146 ( .A(n5819), .ZN(n7157) );
  NAND2_X1 U7147 ( .A1(n7157), .A2(n4402), .ZN(n5384) );
  INV_X1 U7148 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5381) );
  NAND2_X1 U7149 ( .A1(n5803), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5380) );
  NAND2_X1 U7150 ( .A1(n5763), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5379) );
  OAI211_X1 U7151 ( .C1(n5824), .C2(n5381), .A(n5380), .B(n5379), .ZN(n5382)
         );
  INV_X1 U7152 ( .A(n5382), .ZN(n5383) );
  AND2_X2 U7153 ( .A1(n8250), .A2(n9990), .ZN(n7089) );
  AND2_X1 U7154 ( .A1(n10092), .A2(n5854), .ZN(n5385) );
  AND2_X1 U7155 ( .A1(n5943), .A2(n5385), .ZN(n5850) );
  AND2_X1 U7156 ( .A1(n5835), .A2(n5388), .ZN(n5833) );
  NAND2_X1 U7157 ( .A1(n9623), .A2(n5844), .ZN(n5390) );
  NAND2_X1 U7158 ( .A1(n5845), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5389) );
  NOR3_X1 U7159 ( .A1(n5851), .A2(n10093), .A3(n10092), .ZN(n5832) );
  NAND2_X1 U7160 ( .A1(n4402), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5394) );
  NAND2_X1 U7161 ( .A1(n5465), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5392) );
  NAND2_X1 U7162 ( .A1(n5398), .A2(n5395), .ZN(n5410) );
  NAND2_X1 U7163 ( .A1(n7388), .A2(n5396), .ZN(n6195) );
  NAND2_X1 U7164 ( .A1(n5410), .A2(n6195), .ZN(n5397) );
  XNOR2_X1 U7165 ( .A(n5397), .B(SI_1_), .ZN(n5400) );
  MUX2_X1 U7166 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n7389), .Z(n5399) );
  XNOR2_X1 U7167 ( .A(n5400), .B(n5399), .ZN(n6184) );
  INV_X1 U7168 ( .A(n6184), .ZN(n7398) );
  NAND2_X1 U7169 ( .A1(n5430), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5402) );
  NAND2_X1 U7170 ( .A1(n4402), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5406) );
  NAND2_X1 U7171 ( .A1(n5465), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U7172 ( .A1(n5469), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5403) );
  NAND4_X2 U7173 ( .A1(n5406), .A2(n5405), .A3(n5404), .A4(n5403), .ZN(n9808)
         );
  INV_X1 U7174 ( .A(SI_0_), .ZN(n5409) );
  INV_X1 U7175 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5408) );
  OAI21_X1 U7176 ( .B1(n7388), .B2(n5409), .A(n5408), .ZN(n5411) );
  AND2_X1 U7177 ( .A1(n5411), .A2(n5410), .ZN(n10239) );
  OAI21_X2 U7178 ( .B1(n5620), .B2(n10289), .A(n5412), .ZN(n7982) );
  NOR2_X2 U7179 ( .A1(n9808), .A2(n7972), .ZN(n7725) );
  NAND2_X1 U7180 ( .A1(n8087), .A2(n7153), .ZN(n5413) );
  NAND2_X1 U7181 ( .A1(n4402), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5418) );
  NAND2_X1 U7182 ( .A1(n5465), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5417) );
  NAND2_X1 U7183 ( .A1(n5469), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5415) );
  INV_X1 U7184 ( .A(n7090), .ZN(n9805) );
  XNOR2_X1 U7185 ( .A(n5419), .B(SI_2_), .ZN(n5421) );
  MUX2_X1 U7186 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n4522), .Z(n5420) );
  XNOR2_X1 U7187 ( .A(n5421), .B(n5420), .ZN(n7384) );
  NAND2_X1 U7188 ( .A1(n5430), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5422) );
  XNOR2_X2 U7189 ( .A(n9805), .B(n7873), .ZN(n8090) );
  NAND2_X1 U7190 ( .A1(n8925), .A2(n7873), .ZN(n5965) );
  NAND2_X1 U7191 ( .A1(n5465), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5427) );
  INV_X1 U7192 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6789) );
  NAND2_X1 U7193 ( .A1(n4402), .A2(n6789), .ZN(n5425) );
  NAND2_X1 U7194 ( .A1(n5469), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5424) );
  AND4_X2 U7195 ( .A1(n5427), .A2(n5426), .A3(n5425), .A4(n5424), .ZN(n7094)
         );
  XNOR2_X1 U7196 ( .A(n5429), .B(n5428), .ZN(n7391) );
  NAND2_X1 U7197 ( .A1(n5430), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5432) );
  NAND2_X1 U7198 ( .A1(n5655), .A2(n7390), .ZN(n5431) );
  OAI211_X1 U7199 ( .C1(n5524), .C2(n7391), .A(n5432), .B(n5431), .ZN(n7959)
         );
  NAND2_X1 U7200 ( .A1(n7094), .A2(n7959), .ZN(n5971) );
  INV_X1 U7201 ( .A(n7094), .ZN(n9804) );
  NAND2_X1 U7202 ( .A1(n9804), .A2(n10380), .ZN(n5864) );
  INV_X1 U7203 ( .A(n7938), .ZN(n7933) );
  NAND2_X1 U7204 ( .A1(n5465), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5438) );
  INV_X1 U7205 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5433) );
  NAND2_X1 U7206 ( .A1(n5433), .A2(n6789), .ZN(n5434) );
  AND2_X1 U7207 ( .A1(n5434), .A2(n5446), .ZN(n8110) );
  NAND2_X1 U7208 ( .A1(n4402), .A2(n8110), .ZN(n5437) );
  NAND2_X1 U7209 ( .A1(n5762), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U7210 ( .A1(n5469), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5435) );
  XNOR2_X1 U7211 ( .A(n5439), .B(n5440), .ZN(n7393) );
  NAND2_X1 U7212 ( .A1(n7393), .A2(n5800), .ZN(n5442) );
  NAND2_X1 U7213 ( .A1(n5815), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5441) );
  OAI211_X1 U7214 ( .C1(n5620), .C2(n7701), .A(n5442), .B(n5441), .ZN(n8109)
         );
  NAND2_X1 U7215 ( .A1(n7097), .A2(n8109), .ZN(n8052) );
  INV_X1 U7216 ( .A(n8052), .ZN(n5972) );
  NAND2_X1 U7217 ( .A1(n5465), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5451) );
  INV_X1 U7218 ( .A(n5445), .ZN(n5467) );
  NAND2_X1 U7219 ( .A1(n5446), .A2(n4802), .ZN(n5447) );
  AND2_X1 U7220 ( .A1(n5467), .A2(n5447), .ZN(n8051) );
  NAND2_X1 U7221 ( .A1(n4402), .A2(n8051), .ZN(n5450) );
  NAND2_X1 U7222 ( .A1(n5762), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5449) );
  NAND2_X1 U7223 ( .A1(n5469), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5448) );
  XNOR2_X1 U7224 ( .A(n5453), .B(n5452), .ZN(n7401) );
  NAND2_X1 U7225 ( .A1(n7401), .A2(n5800), .ZN(n5456) );
  AOI22_X1 U7226 ( .A1(n5430), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n5655), .B2(
        n5454), .ZN(n5455) );
  NAND2_X1 U7227 ( .A1(n5456), .A2(n5455), .ZN(n8246) );
  AND2_X1 U7228 ( .A1(n7102), .A2(n7096), .ZN(n5868) );
  INV_X1 U7229 ( .A(n9802), .ZN(n8343) );
  NAND2_X1 U7230 ( .A1(n8343), .A2(n8246), .ZN(n8262) );
  NAND2_X1 U7231 ( .A1(n5459), .A2(n5458), .ZN(n5477) );
  XNOR2_X1 U7232 ( .A(n5477), .B(n5461), .ZN(n7403) );
  NAND2_X1 U7233 ( .A1(n7403), .A2(n5800), .ZN(n5463) );
  AOI22_X1 U7234 ( .A1(n5430), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5655), .B2(
        n9818), .ZN(n5462) );
  NAND2_X1 U7235 ( .A1(n5465), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5472) );
  INV_X1 U7236 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5466) );
  NAND2_X1 U7237 ( .A1(n5467), .A2(n5466), .ZN(n5468) );
  AND2_X1 U7238 ( .A1(n5484), .A2(n5468), .ZN(n8345) );
  NAND2_X1 U7239 ( .A1(n4402), .A2(n8345), .ZN(n5471) );
  NAND2_X1 U7240 ( .A1(n5469), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5470) );
  NAND4_X1 U7241 ( .A1(n5473), .A2(n5472), .A3(n5471), .A4(n5470), .ZN(n9801)
         );
  NAND2_X1 U7242 ( .A1(n8346), .A2(n9801), .ZN(n5919) );
  NAND2_X1 U7243 ( .A1(n8260), .A2(n8011), .ZN(n5867) );
  NAND2_X1 U7244 ( .A1(n5919), .A2(n5867), .ZN(n8255) );
  INV_X1 U7245 ( .A(n8255), .ZN(n8264) );
  NAND3_X1 U7246 ( .A1(n5474), .A2(n8052), .A3(n8262), .ZN(n5475) );
  NAND2_X1 U7247 ( .A1(n5475), .A2(n7102), .ZN(n5476) );
  NAND2_X1 U7248 ( .A1(n5477), .A2(n5460), .ZN(n5479) );
  XNOR2_X1 U7249 ( .A(n5480), .B(SI_7_), .ZN(n5498) );
  AOI22_X1 U7250 ( .A1(n5815), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5655), .B2(
        n7488), .ZN(n5481) );
  INV_X1 U7251 ( .A(n8080), .ZN(n5491) );
  NAND2_X1 U7252 ( .A1(n5762), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5489) );
  NAND2_X1 U7253 ( .A1(n5803), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5488) );
  INV_X1 U7254 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5483) );
  NAND2_X1 U7255 ( .A1(n5484), .A2(n5483), .ZN(n5485) );
  AND2_X1 U7256 ( .A1(n5507), .A2(n5485), .ZN(n8079) );
  NAND2_X1 U7257 ( .A1(n4402), .A2(n8079), .ZN(n5487) );
  NAND2_X1 U7258 ( .A1(n5763), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5486) );
  NAND3_X1 U7259 ( .A1(n5492), .A2(n5976), .A3(n5854), .ZN(n5497) );
  XNOR2_X1 U7260 ( .A(n8317), .B(n7089), .ZN(n5494) );
  NAND2_X1 U7261 ( .A1(n5495), .A2(n5494), .ZN(n5496) );
  NAND2_X1 U7262 ( .A1(n5497), .A2(n5496), .ZN(n5583) );
  INV_X1 U7263 ( .A(n5498), .ZN(n5499) );
  NAND2_X1 U7264 ( .A1(n5500), .A2(n5499), .ZN(n5502) );
  NAND2_X1 U7265 ( .A1(n7421), .A2(n5800), .ZN(n5505) );
  AOI22_X1 U7266 ( .A1(n5815), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5655), .B2(
        n7462), .ZN(n5504) );
  NAND2_X1 U7267 ( .A1(n5803), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5512) );
  INV_X1 U7268 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5506) );
  NAND2_X1 U7269 ( .A1(n5507), .A2(n5506), .ZN(n5508) );
  AND2_X1 U7270 ( .A1(n5516), .A2(n5508), .ZN(n8324) );
  NAND2_X1 U7271 ( .A1(n4402), .A2(n8324), .ZN(n5511) );
  NAND2_X1 U7272 ( .A1(n5762), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U7273 ( .A1(n5763), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5509) );
  AND4_X2 U7274 ( .A1(n5512), .A2(n5511), .A3(n5510), .A4(n5509), .ZN(n8386)
         );
  NAND2_X1 U7275 ( .A1(n10427), .A2(n8386), .ZN(n5921) );
  XNOR2_X1 U7276 ( .A(n5513), .B(n5039), .ZN(n7410) );
  NAND2_X1 U7277 ( .A1(n7410), .A2(n5800), .ZN(n5515) );
  AOI22_X1 U7278 ( .A1(n5845), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5655), .B2(
        n7527), .ZN(n5514) );
  NAND2_X1 U7279 ( .A1(n5465), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U7280 ( .A1(n5762), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U7281 ( .A1(n5516), .A2(n7526), .ZN(n5517) );
  AND2_X1 U7282 ( .A1(n5575), .A2(n5517), .ZN(n8529) );
  NAND2_X1 U7283 ( .A1(n4402), .A2(n8529), .ZN(n5519) );
  NAND2_X1 U7284 ( .A1(n5763), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5518) );
  NAND4_X1 U7285 ( .A1(n5521), .A2(n5520), .A3(n5519), .A4(n5518), .ZN(n9798)
         );
  INV_X1 U7286 ( .A(n9798), .ZN(n8511) );
  OR2_X1 U7287 ( .A1(n8535), .A2(n8511), .ZN(n7017) );
  NAND2_X1 U7288 ( .A1(n7015), .A2(n7017), .ZN(n5907) );
  AOI21_X1 U7289 ( .B1(n5583), .B2(n5921), .A(n5907), .ZN(n5603) );
  XNOR2_X1 U7290 ( .A(n5523), .B(n5522), .ZN(n7512) );
  NAND2_X1 U7291 ( .A1(n7512), .A2(n5844), .ZN(n5527) );
  AOI22_X1 U7292 ( .A1(n5815), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5525), .B2(
        n5655), .ZN(n5526) );
  NAND2_X1 U7293 ( .A1(n5540), .A2(n5528), .ZN(n5529) );
  NAND2_X1 U7294 ( .A1(n5591), .A2(n5529), .ZN(n9648) );
  NAND2_X1 U7295 ( .A1(n5803), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U7296 ( .A1(n5763), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5530) );
  AND2_X1 U7297 ( .A1(n5531), .A2(n5530), .ZN(n5533) );
  NAND2_X1 U7298 ( .A1(n5762), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5532) );
  OAI211_X1 U7299 ( .C1(n5821), .C2(n9648), .A(n5533), .B(n5532), .ZN(n10069)
         );
  INV_X1 U7300 ( .A(n10069), .ZN(n10039) );
  NAND2_X1 U7301 ( .A1(n10181), .A2(n10039), .ZN(n5595) );
  XNOR2_X1 U7302 ( .A(n5534), .B(n5040), .ZN(n7481) );
  NAND2_X1 U7303 ( .A1(n7481), .A2(n5844), .ZN(n5538) );
  OAI22_X1 U7304 ( .A1(n8140), .A2(n5620), .B1(n5535), .B2(n7498), .ZN(n5536)
         );
  INV_X1 U7305 ( .A(n5536), .ZN(n5537) );
  NAND2_X1 U7306 ( .A1(n5762), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U7307 ( .A1(n5803), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5543) );
  NAND2_X1 U7308 ( .A1(n5550), .A2(n8139), .ZN(n5539) );
  AND2_X1 U7309 ( .A1(n5540), .A2(n5539), .ZN(n10058) );
  NAND2_X1 U7310 ( .A1(n4402), .A2(n10058), .ZN(n5542) );
  NAND2_X1 U7311 ( .A1(n5763), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5541) );
  NAND4_X1 U7312 ( .A1(n5544), .A2(n5543), .A3(n5542), .A4(n5541), .ZN(n9794)
         );
  INV_X1 U7313 ( .A(n9794), .ZN(n9645) );
  NAND2_X1 U7314 ( .A1(n10061), .A2(n9645), .ZN(n7023) );
  NAND2_X1 U7315 ( .A1(n5595), .A2(n7023), .ZN(n5925) );
  XNOR2_X1 U7316 ( .A(n5546), .B(n5545), .ZN(n6314) );
  NAND2_X1 U7317 ( .A1(n6314), .A2(n5800), .ZN(n5548) );
  AOI22_X1 U7318 ( .A1(n5845), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5655), .B2(
        n7896), .ZN(n5547) );
  NAND2_X1 U7319 ( .A1(n5762), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5554) );
  NAND2_X1 U7320 ( .A1(n5803), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5553) );
  INV_X1 U7321 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7895) );
  NAND2_X1 U7322 ( .A1(n5560), .A2(n7895), .ZN(n5549) );
  AND2_X1 U7323 ( .A1(n5550), .A2(n5549), .ZN(n8635) );
  NAND2_X1 U7324 ( .A1(n4402), .A2(n8635), .ZN(n5552) );
  NAND2_X1 U7325 ( .A1(n5763), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5551) );
  XNOR2_X1 U7326 ( .A(n5556), .B(n5555), .ZN(n7428) );
  NAND2_X1 U7327 ( .A1(n7428), .A2(n5800), .ZN(n5558) );
  AOI22_X1 U7328 ( .A1(n5845), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5655), .B2(
        n7659), .ZN(n5557) );
  NAND2_X2 U7329 ( .A1(n5558), .A2(n5557), .ZN(n10196) );
  NAND2_X1 U7330 ( .A1(n5762), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U7331 ( .A1(n5803), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5563) );
  NAND2_X1 U7332 ( .A1(n5577), .A2(n7658), .ZN(n5559) );
  AND2_X1 U7333 ( .A1(n5560), .A2(n5559), .ZN(n8566) );
  NAND2_X1 U7334 ( .A1(n4402), .A2(n8566), .ZN(n5562) );
  NAND2_X1 U7335 ( .A1(n5763), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5561) );
  NAND4_X1 U7336 ( .A1(n5564), .A2(n5563), .A3(n5562), .A4(n5561), .ZN(n9796)
         );
  OR2_X1 U7337 ( .A1(n10196), .A2(n8510), .ZN(n8623) );
  AND2_X1 U7338 ( .A1(n5861), .A2(n8623), .ZN(n7022) );
  NAND2_X1 U7339 ( .A1(n10065), .A2(n5854), .ZN(n5565) );
  OR2_X1 U7340 ( .A1(n10061), .A2(n9645), .ZN(n5910) );
  OAI21_X1 U7341 ( .B1(n7022), .B2(n5565), .A(n5910), .ZN(n5566) );
  INV_X1 U7342 ( .A(n5566), .ZN(n5567) );
  OR2_X1 U7343 ( .A1(n5925), .A2(n5567), .ZN(n5570) );
  NAND2_X1 U7344 ( .A1(n5925), .A2(n7089), .ZN(n5569) );
  OR2_X1 U7345 ( .A1(n10181), .A2(n10039), .ZN(n7024) );
  NAND2_X1 U7346 ( .A1(n10196), .A2(n8510), .ZN(n7021) );
  NAND2_X1 U7347 ( .A1(n10065), .A2(n7021), .ZN(n5920) );
  NAND3_X1 U7348 ( .A1(n5920), .A2(n7089), .A3(n5861), .ZN(n5568) );
  NAND4_X1 U7349 ( .A1(n5570), .A2(n5569), .A3(n7024), .A4(n5568), .ZN(n5599)
         );
  INV_X1 U7350 ( .A(n5599), .ZN(n5582) );
  NAND2_X1 U7351 ( .A1(n7419), .A2(n5800), .ZN(n5573) );
  AOI22_X1 U7352 ( .A1(n5845), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5655), .B2(
        n7425), .ZN(n5572) );
  NAND2_X1 U7353 ( .A1(n5573), .A2(n5572), .ZN(n8641) );
  NAND2_X1 U7354 ( .A1(n5803), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5581) );
  NAND2_X1 U7355 ( .A1(n5762), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5580) );
  INV_X1 U7356 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5574) );
  NAND2_X1 U7357 ( .A1(n5575), .A2(n5574), .ZN(n5576) );
  AND2_X1 U7358 ( .A1(n5577), .A2(n5576), .ZN(n8640) );
  NAND2_X1 U7359 ( .A1(n4402), .A2(n8640), .ZN(n5579) );
  NAND2_X1 U7360 ( .A1(n5763), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U7361 ( .A1(n8641), .A2(n8533), .ZN(n5862) );
  NAND2_X1 U7362 ( .A1(n8535), .A2(n8511), .ZN(n5866) );
  AND2_X1 U7363 ( .A1(n5862), .A2(n5866), .ZN(n5922) );
  NAND3_X1 U7364 ( .A1(n5582), .A2(n7089), .A3(n5922), .ZN(n5602) );
  NAND3_X1 U7365 ( .A1(n5861), .A2(n7089), .A3(n7019), .ZN(n5585) );
  NAND2_X1 U7366 ( .A1(n5862), .A2(n5854), .ZN(n5584) );
  NAND2_X1 U7367 ( .A1(n5585), .A2(n5584), .ZN(n5586) );
  XNOR2_X1 U7368 ( .A(n10196), .B(n9796), .ZN(n8558) );
  NAND3_X1 U7369 ( .A1(n5586), .A2(n10065), .A3(n8558), .ZN(n5587) );
  NOR2_X1 U7370 ( .A1(n5925), .A2(n5587), .ZN(n5598) );
  XNOR2_X1 U7371 ( .A(n5588), .B(n5589), .ZN(n7679) );
  NAND2_X1 U7372 ( .A1(n7679), .A2(n5844), .ZN(n7122) );
  AOI22_X1 U7373 ( .A1(n10316), .A2(n5655), .B1(n5815), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n7120) );
  INV_X1 U7374 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10218) );
  INV_X1 U7375 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5590) );
  NAND2_X1 U7376 ( .A1(n5591), .A2(n5590), .ZN(n5592) );
  NAND2_X1 U7377 ( .A1(n5606), .A2(n5592), .ZN(n10050) );
  OR2_X1 U7378 ( .A1(n10050), .A2(n5821), .ZN(n5594) );
  AOI22_X1 U7379 ( .A1(n5762), .A2(P1_REG1_REG_15__SCAN_IN), .B1(n5803), .B2(
        P1_REG2_REG_15__SCAN_IN), .ZN(n5593) );
  OAI211_X1 U7380 ( .C1(n5367), .C2(n10218), .A(n5594), .B(n5593), .ZN(n10012)
         );
  INV_X1 U7381 ( .A(n10012), .ZN(n9698) );
  OR2_X1 U7382 ( .A1(n10170), .A2(n9698), .ZN(n7026) );
  NAND2_X1 U7383 ( .A1(n10170), .A2(n9698), .ZN(n7025) );
  AND2_X2 U7384 ( .A1(n7026), .A2(n7025), .ZN(n10037) );
  NAND2_X1 U7385 ( .A1(n7024), .A2(n5910), .ZN(n5596) );
  NAND3_X1 U7386 ( .A1(n5596), .A2(n7089), .A3(n5595), .ZN(n5597) );
  OAI211_X1 U7387 ( .C1(n5599), .C2(n5598), .A(n10037), .B(n5597), .ZN(n5600)
         );
  INV_X1 U7388 ( .A(n5600), .ZN(n5601) );
  NAND2_X1 U7389 ( .A1(n7704), .A2(n5844), .ZN(n5605) );
  AOI22_X1 U7390 ( .A1(n5815), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7705), .B2(
        n5655), .ZN(n5604) );
  NAND2_X1 U7391 ( .A1(n5606), .A2(n4819), .ZN(n5607) );
  NAND2_X1 U7392 ( .A1(n5624), .A2(n5607), .ZN(n10018) );
  OR2_X1 U7393 ( .A1(n10018), .A2(n5821), .ZN(n5610) );
  AOI22_X1 U7394 ( .A1(n5803), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n5763), .B2(
        P1_REG0_REG_16__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U7395 ( .A1(n5762), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5608) );
  MUX2_X1 U7396 ( .A(n7026), .B(n7025), .S(n7089), .Z(n5613) );
  NAND2_X1 U7397 ( .A1(n5617), .A2(n5616), .ZN(n5619) );
  NAND2_X1 U7398 ( .A1(n7832), .A2(n5844), .ZN(n5623) );
  OAI22_X1 U7399 ( .A1(n10338), .A2(n5620), .B1(n5535), .B2(n7835), .ZN(n5621)
         );
  INV_X1 U7400 ( .A(n5621), .ZN(n5622) );
  NAND2_X1 U7401 ( .A1(n5624), .A2(n9714), .ZN(n5625) );
  AND2_X1 U7402 ( .A1(n5640), .A2(n5625), .ZN(n9997) );
  NAND2_X1 U7403 ( .A1(n9997), .A2(n4402), .ZN(n5631) );
  NAND2_X1 U7404 ( .A1(n5763), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5627) );
  NAND2_X1 U7405 ( .A1(n5803), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5626) );
  OAI211_X1 U7406 ( .C1(n5824), .C2(n5628), .A(n5627), .B(n5626), .ZN(n5629)
         );
  INV_X1 U7407 ( .A(n5629), .ZN(n5630) );
  NAND2_X1 U7408 ( .A1(n5631), .A2(n5630), .ZN(n10013) );
  INV_X1 U7409 ( .A(n10013), .ZN(n9983) );
  AND2_X1 U7410 ( .A1(n10159), .A2(n9983), .ZN(n9977) );
  INV_X1 U7411 ( .A(n9977), .ZN(n5904) );
  OR2_X1 U7412 ( .A1(n10159), .A2(n9983), .ZN(n9978) );
  NAND2_X1 U7413 ( .A1(n7879), .A2(n5844), .ZN(n5639) );
  AOI22_X1 U7414 ( .A1(n5637), .A2(n5655), .B1(n5815), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n5638) );
  NAND2_X2 U7415 ( .A1(n5639), .A2(n5638), .ZN(n10156) );
  NAND2_X1 U7416 ( .A1(n5640), .A2(n4812), .ZN(n5641) );
  NAND2_X1 U7417 ( .A1(n5659), .A2(n5641), .ZN(n9989) );
  OR2_X1 U7418 ( .A1(n9989), .A2(n5821), .ZN(n5647) );
  NAND2_X1 U7419 ( .A1(n5763), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5643) );
  NAND2_X1 U7420 ( .A1(n5803), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5642) );
  OAI211_X1 U7421 ( .C1(n5824), .C2(n5644), .A(n5643), .B(n5642), .ZN(n5645)
         );
  INV_X1 U7422 ( .A(n5645), .ZN(n5646) );
  NOR2_X1 U7423 ( .A1(n8789), .A2(n5854), .ZN(n5682) );
  AND2_X1 U7424 ( .A1(n8789), .A2(n5854), .ZN(n5674) );
  INV_X1 U7425 ( .A(n5674), .ZN(n5677) );
  NAND2_X1 U7426 ( .A1(n10156), .A2(n5677), .ZN(n5648) );
  OAI21_X1 U7427 ( .B1(n10156), .B2(n5682), .A(n5648), .ZN(n5673) );
  NAND2_X1 U7428 ( .A1(n5650), .A2(n5649), .ZN(n5652) );
  AND2_X1 U7429 ( .A1(n5652), .A2(n5651), .ZN(n5654) );
  NAND2_X1 U7430 ( .A1(n7883), .A2(n5844), .ZN(n5657) );
  AOI22_X1 U7431 ( .A1(n5845), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9990), .B2(
        n5655), .ZN(n5656) );
  NAND2_X2 U7432 ( .A1(n5657), .A2(n5656), .ZN(n10150) );
  NAND2_X1 U7433 ( .A1(n5659), .A2(n5658), .ZN(n5660) );
  AND2_X1 U7434 ( .A1(n5694), .A2(n5660), .ZN(n9960) );
  NAND2_X1 U7435 ( .A1(n9960), .A2(n4402), .ZN(n5666) );
  INV_X1 U7436 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U7437 ( .A1(n5762), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5662) );
  NAND2_X1 U7438 ( .A1(n5803), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5661) );
  OAI211_X1 U7439 ( .C1(n5663), .C2(n5367), .A(n5662), .B(n5661), .ZN(n5664)
         );
  INV_X1 U7440 ( .A(n5664), .ZN(n5665) );
  NAND2_X1 U7441 ( .A1(n5666), .A2(n5665), .ZN(n9793) );
  NAND2_X1 U7442 ( .A1(n9793), .A2(n7089), .ZN(n5683) );
  OR2_X1 U7443 ( .A1(n9793), .A2(n7089), .ZN(n5675) );
  INV_X1 U7444 ( .A(n5675), .ZN(n5667) );
  NAND2_X1 U7445 ( .A1(n10150), .A2(n5667), .ZN(n5668) );
  OAI21_X1 U7446 ( .B1(n10150), .B2(n5683), .A(n5668), .ZN(n5671) );
  MUX2_X1 U7447 ( .A(n7029), .B(n7028), .S(n7089), .Z(n5669) );
  INV_X1 U7448 ( .A(n5669), .ZN(n5670) );
  NOR2_X1 U7449 ( .A1(n5671), .A2(n5670), .ZN(n5672) );
  INV_X1 U7450 ( .A(n9793), .ZN(n9984) );
  OR2_X1 U7451 ( .A1(n10150), .A2(n9984), .ZN(n5896) );
  AND2_X1 U7452 ( .A1(n5860), .A2(n9978), .ZN(n7032) );
  NAND3_X1 U7453 ( .A1(n5896), .A2(n7032), .A3(n5854), .ZN(n5689) );
  NAND2_X1 U7454 ( .A1(n10150), .A2(n9984), .ZN(n5931) );
  NAND4_X1 U7455 ( .A1(n5931), .A2(n7089), .A3(n5905), .A4(n5904), .ZN(n5688)
         );
  NAND2_X1 U7456 ( .A1(n10156), .A2(n5674), .ZN(n5676) );
  NAND2_X1 U7457 ( .A1(n5676), .A2(n5675), .ZN(n5681) );
  OAI21_X1 U7458 ( .B1(n9793), .B2(n5677), .A(n10156), .ZN(n5680) );
  AND2_X1 U7459 ( .A1(n5682), .A2(n9793), .ZN(n5678) );
  OR2_X1 U7460 ( .A1(n10156), .A2(n5678), .ZN(n5679) );
  AOI22_X1 U7461 ( .A1(n10150), .A2(n5681), .B1(n5680), .B2(n5679), .ZN(n5687)
         );
  INV_X1 U7462 ( .A(n10150), .ZN(n9962) );
  INV_X1 U7463 ( .A(n5682), .ZN(n5684) );
  OAI21_X1 U7464 ( .B1(n10156), .B2(n5684), .A(n5683), .ZN(n5685) );
  NAND2_X1 U7465 ( .A1(n9962), .A2(n5685), .ZN(n5686) );
  NAND4_X1 U7466 ( .A1(n5689), .A2(n5688), .A3(n5687), .A4(n5686), .ZN(n5703)
         );
  XNOR2_X1 U7467 ( .A(n5691), .B(n5690), .ZN(n7979) );
  NAND2_X1 U7468 ( .A1(n7979), .A2(n5844), .ZN(n5693) );
  NAND2_X1 U7469 ( .A1(n5815), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5692) );
  NAND2_X1 U7470 ( .A1(n5694), .A2(n4813), .ZN(n5695) );
  NAND2_X1 U7471 ( .A1(n5711), .A2(n5695), .ZN(n9951) );
  OR2_X1 U7472 ( .A1(n9951), .A2(n5821), .ZN(n5701) );
  INV_X1 U7473 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n5698) );
  NAND2_X1 U7474 ( .A1(n5763), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5697) );
  NAND2_X1 U7475 ( .A1(n5803), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5696) );
  OAI211_X1 U7476 ( .C1(n5824), .C2(n5698), .A(n5697), .B(n5696), .ZN(n5699)
         );
  INV_X1 U7477 ( .A(n5699), .ZN(n5700) );
  NAND2_X1 U7478 ( .A1(n5701), .A2(n5700), .ZN(n9970) );
  INV_X1 U7479 ( .A(n9970), .ZN(n9929) );
  AND2_X1 U7480 ( .A1(n10146), .A2(n9929), .ZN(n7035) );
  INV_X1 U7481 ( .A(n7035), .ZN(n5771) );
  NAND2_X1 U7482 ( .A1(n5771), .A2(n7036), .ZN(n9946) );
  NAND2_X1 U7483 ( .A1(n5705), .A2(n5704), .ZN(n5773) );
  NAND2_X1 U7484 ( .A1(n7996), .A2(n5844), .ZN(n5709) );
  NAND2_X1 U7485 ( .A1(n5845), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5708) );
  NAND2_X1 U7486 ( .A1(n5711), .A2(n5710), .ZN(n5712) );
  AND2_X1 U7487 ( .A1(n5724), .A2(n5712), .ZN(n9933) );
  NAND2_X1 U7488 ( .A1(n9933), .A2(n4402), .ZN(n5718) );
  INV_X1 U7489 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n5715) );
  NAND2_X1 U7490 ( .A1(n5803), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5714) );
  NAND2_X1 U7491 ( .A1(n5763), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5713) );
  OAI211_X1 U7492 ( .C1(n5824), .C2(n5715), .A(n5714), .B(n5713), .ZN(n5716)
         );
  INV_X1 U7493 ( .A(n5716), .ZN(n5717) );
  NAND2_X1 U7494 ( .A1(n10141), .A2(n9948), .ZN(n7039) );
  INV_X1 U7495 ( .A(n7039), .ZN(n5719) );
  XNOR2_X1 U7496 ( .A(n5721), .B(n5720), .ZN(n6413) );
  INV_X1 U7497 ( .A(n6413), .ZN(n8959) );
  NAND2_X1 U7498 ( .A1(n6413), .A2(n5844), .ZN(n5723) );
  NAND2_X1 U7499 ( .A1(n5815), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5722) );
  INV_X1 U7500 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9745) );
  NAND2_X1 U7501 ( .A1(n5724), .A2(n9745), .ZN(n5725) );
  NAND2_X1 U7502 ( .A1(n5735), .A2(n5725), .ZN(n9913) );
  INV_X1 U7503 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n6815) );
  NAND2_X1 U7504 ( .A1(n5763), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5727) );
  NAND2_X1 U7505 ( .A1(n5803), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5726) );
  OAI211_X1 U7506 ( .C1(n5824), .C2(n6815), .A(n5727), .B(n5726), .ZN(n5728)
         );
  INV_X1 U7507 ( .A(n5728), .ZN(n5729) );
  OR2_X1 U7508 ( .A1(n10141), .A2(n9948), .ZN(n5859) );
  NAND2_X1 U7509 ( .A1(n7040), .A2(n5859), .ZN(n5899) );
  NAND2_X1 U7510 ( .A1(n10134), .A2(n9930), .ZN(n7041) );
  XNOR2_X1 U7511 ( .A(n5732), .B(n5731), .ZN(n8331) );
  NAND2_X1 U7512 ( .A1(n8331), .A2(n5844), .ZN(n5734) );
  NAND2_X1 U7513 ( .A1(n5845), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5733) );
  NAND2_X1 U7514 ( .A1(n5735), .A2(n4815), .ZN(n5736) );
  NAND2_X1 U7515 ( .A1(n5748), .A2(n5736), .ZN(n9897) );
  INV_X1 U7516 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n6935) );
  NAND2_X1 U7517 ( .A1(n5762), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5738) );
  NAND2_X1 U7518 ( .A1(n5803), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5737) );
  OAI211_X1 U7519 ( .C1(n6935), .C2(n5367), .A(n5738), .B(n5737), .ZN(n5739)
         );
  INV_X1 U7520 ( .A(n5739), .ZN(n5740) );
  NAND2_X1 U7521 ( .A1(n10129), .A2(n9887), .ZN(n5934) );
  NAND2_X1 U7522 ( .A1(n5743), .A2(n5742), .ZN(n5745) );
  NAND2_X1 U7523 ( .A1(n8477), .A2(n5844), .ZN(n5747) );
  NAND2_X1 U7524 ( .A1(n5815), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5746) );
  NAND2_X1 U7525 ( .A1(n5748), .A2(n9725), .ZN(n5749) );
  NAND2_X1 U7526 ( .A1(n5760), .A2(n5749), .ZN(n9889) );
  INV_X1 U7527 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n6916) );
  NAND2_X1 U7528 ( .A1(n5762), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5751) );
  NAND2_X1 U7529 ( .A1(n5763), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5750) );
  OAI211_X1 U7530 ( .C1(n5766), .C2(n6916), .A(n5751), .B(n5750), .ZN(n5752)
         );
  INV_X1 U7531 ( .A(n5752), .ZN(n5753) );
  NAND2_X1 U7532 ( .A1(n10127), .A2(n9871), .ZN(n9868) );
  NAND2_X1 U7533 ( .A1(n8573), .A2(n5844), .ZN(n5758) );
  NAND2_X1 U7534 ( .A1(n5845), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5757) );
  NAND2_X1 U7535 ( .A1(n5760), .A2(n5759), .ZN(n5761) );
  NAND2_X1 U7536 ( .A1(n9874), .A2(n4402), .ZN(n5769) );
  INV_X1 U7537 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n6811) );
  NAND2_X1 U7538 ( .A1(n5762), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5765) );
  NAND2_X1 U7539 ( .A1(n5763), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5764) );
  OAI211_X1 U7540 ( .C1(n5766), .C2(n6811), .A(n5765), .B(n5764), .ZN(n5767)
         );
  INV_X1 U7541 ( .A(n5767), .ZN(n5768) );
  NAND2_X1 U7542 ( .A1(n10123), .A2(n9888), .ZN(n5858) );
  NAND2_X1 U7543 ( .A1(n5858), .A2(n9868), .ZN(n9847) );
  OAI21_X1 U7544 ( .B1(n5770), .B2(n9847), .A(n7089), .ZN(n5777) );
  NAND2_X1 U7545 ( .A1(n5935), .A2(n9881), .ZN(n5900) );
  INV_X1 U7546 ( .A(n9849), .ZN(n5791) );
  AOI21_X1 U7547 ( .B1(n9868), .B2(n5900), .A(n5791), .ZN(n5775) );
  INV_X1 U7548 ( .A(n5859), .ZN(n5772) );
  OAI211_X1 U7549 ( .C1(n5772), .C2(n5771), .A(n7041), .B(n7039), .ZN(n5930)
         );
  NAND2_X1 U7550 ( .A1(n5930), .A2(n7040), .ZN(n5895) );
  OAI211_X1 U7551 ( .C1(n5773), .C2(n5899), .A(n5895), .B(n5934), .ZN(n5774)
         );
  INV_X1 U7552 ( .A(n5808), .ZN(n5812) );
  INV_X1 U7553 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9766) );
  NAND2_X1 U7554 ( .A1(n5778), .A2(n9766), .ZN(n5779) );
  NAND2_X1 U7555 ( .A1(n5818), .A2(n5779), .ZN(n9863) );
  INV_X1 U7556 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n5782) );
  NAND2_X1 U7557 ( .A1(n5803), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5781) );
  NAND2_X1 U7558 ( .A1(n5763), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5780) );
  OAI211_X1 U7559 ( .C1(n5824), .C2(n5782), .A(n5781), .B(n5780), .ZN(n5783)
         );
  INV_X1 U7560 ( .A(n5783), .ZN(n5784) );
  NAND2_X1 U7561 ( .A1(n9872), .A2(n7089), .ZN(n5793) );
  NAND2_X1 U7562 ( .A1(n8685), .A2(n5844), .ZN(n5789) );
  NAND2_X1 U7563 ( .A1(n5845), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5788) );
  NAND3_X1 U7564 ( .A1(n9858), .A2(n5858), .A3(n5854), .ZN(n5790) );
  OAI21_X1 U7565 ( .B1(n5791), .B2(n5793), .A(n5790), .ZN(n5811) );
  AOI21_X1 U7566 ( .B1(n9791), .B2(n5854), .A(n10116), .ZN(n5792) );
  AOI21_X1 U7567 ( .B1(n10116), .B2(n5793), .A(n5792), .ZN(n5810) );
  AND2_X1 U7568 ( .A1(n5797), .A2(n5796), .ZN(n5798) );
  NAND2_X1 U7569 ( .A1(n8691), .A2(n5800), .ZN(n5802) );
  NAND2_X1 U7570 ( .A1(n5845), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5801) );
  INV_X1 U7571 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n6837) );
  NAND2_X1 U7572 ( .A1(n5803), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5805) );
  NAND2_X1 U7573 ( .A1(n5763), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5804) );
  OAI211_X1 U7574 ( .C1(n6837), .C2(n5824), .A(n5805), .B(n5804), .ZN(n5806)
         );
  AOI21_X1 U7575 ( .B1(n5808), .B2(n7149), .A(n5807), .ZN(n5809) );
  NAND2_X1 U7576 ( .A1(n8715), .A2(n5844), .ZN(n5817) );
  NAND2_X1 U7577 ( .A1(n5815), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5816) );
  OAI21_X1 U7578 ( .B1(n5818), .B2(n9633), .A(n8880), .ZN(n5820) );
  NAND2_X1 U7579 ( .A1(n5820), .A2(n5819), .ZN(n8942) );
  INV_X1 U7580 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6894) );
  NAND2_X1 U7581 ( .A1(n5803), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5823) );
  NAND2_X1 U7582 ( .A1(n5763), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5822) );
  OAI211_X1 U7583 ( .C1(n5824), .C2(n6894), .A(n5823), .B(n5822), .ZN(n5825)
         );
  INV_X1 U7584 ( .A(n5825), .ZN(n5826) );
  NAND2_X1 U7585 ( .A1(n10107), .A2(n9634), .ZN(n7049) );
  MUX2_X1 U7586 ( .A(n5941), .B(n7048), .S(n7089), .Z(n5828) );
  NAND2_X1 U7587 ( .A1(n8948), .A2(n5828), .ZN(n5830) );
  MUX2_X1 U7588 ( .A(n5893), .B(n7049), .S(n7089), .Z(n5829) );
  OAI21_X1 U7589 ( .B1(n5831), .B2(n5830), .A(n5829), .ZN(n5853) );
  OAI21_X1 U7590 ( .B1(n5850), .B2(n5832), .A(n5853), .ZN(n5856) );
  INV_X1 U7591 ( .A(n10093), .ZN(n10095) );
  AOI21_X1 U7592 ( .B1(n5943), .B2(n10095), .A(n5854), .ZN(n5849) );
  NOR2_X1 U7593 ( .A1(n10087), .A2(n7057), .ZN(n5996) );
  INV_X1 U7594 ( .A(n9788), .ZN(n9837) );
  INV_X1 U7595 ( .A(SI_30_), .ZN(n5839) );
  NAND2_X1 U7596 ( .A1(n5834), .A2(n5833), .ZN(n5837) );
  NAND3_X1 U7597 ( .A1(n5837), .A2(n5836), .A3(n5835), .ZN(n5838) );
  MUX2_X1 U7598 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7388), .Z(n5841) );
  XNOR2_X1 U7599 ( .A(n5841), .B(SI_31_), .ZN(n5842) );
  NAND2_X1 U7600 ( .A1(n9617), .A2(n5844), .ZN(n5847) );
  NAND2_X1 U7601 ( .A1(n5845), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n5846) );
  INV_X1 U7602 ( .A(n5948), .ZN(n5848) );
  AOI211_X1 U7603 ( .C1(n10095), .C2(n5850), .A(n5849), .B(n5848), .ZN(n5855)
         );
  INV_X1 U7604 ( .A(n10092), .ZN(n5852) );
  INV_X1 U7605 ( .A(n7617), .ZN(n7055) );
  INV_X1 U7606 ( .A(n10083), .ZN(n9839) );
  NOR2_X1 U7607 ( .A1(n9839), .A2(n9788), .ZN(n5998) );
  AND2_X1 U7608 ( .A1(n10087), .A2(n7057), .ZN(n5993) );
  AND2_X1 U7609 ( .A1(n10116), .A2(n9872), .ZN(n7044) );
  INV_X1 U7610 ( .A(n7044), .ZN(n5857) );
  NAND2_X1 U7611 ( .A1(n9858), .A2(n9791), .ZN(n5938) );
  NAND2_X1 U7612 ( .A1(n5857), .A2(n5938), .ZN(n9856) );
  INV_X1 U7613 ( .A(n9856), .ZN(n5887) );
  NAND2_X1 U7614 ( .A1(n5860), .A2(n5905), .ZN(n9976) );
  INV_X1 U7615 ( .A(n9976), .ZN(n9980) );
  INV_X1 U7616 ( .A(n10037), .ZN(n5879) );
  XNOR2_X1 U7617 ( .A(n10181), .B(n10039), .ZN(n8742) );
  NAND2_X1 U7618 ( .A1(n5861), .A2(n10065), .ZN(n8625) );
  INV_X1 U7619 ( .A(n8625), .ZN(n7114) );
  NAND2_X1 U7620 ( .A1(n7019), .A2(n5862), .ZN(n8508) );
  INV_X1 U7621 ( .A(n8508), .ZN(n8505) );
  NAND2_X1 U7622 ( .A1(n8505), .A2(n8319), .ZN(n5876) );
  NAND2_X1 U7623 ( .A1(n5919), .A2(n7102), .ZN(n5863) );
  AND2_X1 U7624 ( .A1(n5863), .A2(n5867), .ZN(n7012) );
  NAND2_X1 U7625 ( .A1(n7096), .A2(n5864), .ZN(n5865) );
  NOR2_X1 U7626 ( .A1(n7012), .A2(n5865), .ZN(n5968) );
  NAND2_X1 U7627 ( .A1(n5867), .A2(n8262), .ZN(n5973) );
  INV_X1 U7628 ( .A(n5973), .ZN(n5871) );
  NAND2_X1 U7629 ( .A1(n8052), .A2(n5971), .ZN(n5869) );
  NAND2_X1 U7630 ( .A1(n5869), .A2(n5868), .ZN(n5870) );
  NAND2_X1 U7631 ( .A1(n5871), .A2(n5870), .ZN(n5918) );
  AND2_X1 U7632 ( .A1(n9808), .A2(n7972), .ZN(n5963) );
  NOR2_X1 U7633 ( .A1(n7725), .A2(n5963), .ZN(n7969) );
  NAND3_X1 U7634 ( .A1(n7969), .A2(n8090), .A3(n5872), .ZN(n5873) );
  NOR2_X1 U7635 ( .A1(n5918), .A2(n5873), .ZN(n5874) );
  NAND4_X1 U7636 ( .A1(n5968), .A2(n8384), .A3(n5874), .A4(n7101), .ZN(n5875)
         );
  NOR2_X1 U7637 ( .A1(n5876), .A2(n5875), .ZN(n5877) );
  NAND4_X1 U7638 ( .A1(n10064), .A2(n7114), .A3(n5877), .A4(n8558), .ZN(n5878)
         );
  NOR3_X1 U7639 ( .A1(n5879), .A2(n8742), .A3(n5878), .ZN(n5880) );
  AND2_X1 U7640 ( .A1(n7123), .A2(n5880), .ZN(n5881) );
  NAND4_X1 U7641 ( .A1(n9969), .A2(n9980), .A3(n10001), .A4(n5881), .ZN(n5882)
         );
  NOR2_X1 U7642 ( .A1(n9946), .A2(n5882), .ZN(n5883) );
  NAND3_X1 U7643 ( .A1(n9917), .A2(n7139), .A3(n5883), .ZN(n5884) );
  NAND2_X1 U7644 ( .A1(n9881), .A2(n5934), .ZN(n9902) );
  OR3_X1 U7645 ( .A1(n5884), .A2(n9886), .A3(n9902), .ZN(n5885) );
  NOR2_X1 U7646 ( .A1(n9869), .A2(n5885), .ZN(n5886) );
  NAND4_X1 U7647 ( .A1(n8948), .A2(n7149), .A3(n5887), .A4(n5886), .ZN(n5888)
         );
  NOR4_X1 U7648 ( .A1(n5998), .A2(n5996), .A3(n5993), .A4(n5888), .ZN(n5890)
         );
  XNOR2_X1 U7649 ( .A(n10093), .B(n10092), .ZN(n10101) );
  INV_X1 U7650 ( .A(n10101), .ZN(n10091) );
  NOR2_X1 U7651 ( .A1(n5947), .A2(n10091), .ZN(n5889) );
  AOI21_X1 U7652 ( .B1(n5890), .B2(n5889), .A(n4495), .ZN(n5951) );
  AOI21_X1 U7653 ( .B1(n5891), .B2(n7055), .A(n5951), .ZN(n5961) );
  INV_X1 U7654 ( .A(n5947), .ZN(n5995) );
  NAND4_X1 U7655 ( .A1(n5892), .A2(n4495), .A3(n8250), .A4(n5995), .ZN(n5960)
         );
  INV_X1 U7656 ( .A(n5893), .ZN(n5894) );
  AOI21_X1 U7657 ( .B1(n10095), .B2(n10092), .A(n5894), .ZN(n5992) );
  INV_X1 U7658 ( .A(n5992), .ZN(n5945) );
  INV_X1 U7659 ( .A(n5895), .ZN(n5903) );
  INV_X1 U7660 ( .A(n5896), .ZN(n5898) );
  INV_X1 U7661 ( .A(n5931), .ZN(n7034) );
  INV_X1 U7662 ( .A(n5905), .ZN(n7033) );
  NOR3_X1 U7663 ( .A1(n7034), .A2(n7032), .A3(n7033), .ZN(n5897) );
  NOR4_X1 U7664 ( .A1(n5899), .A2(n4697), .A3(n5898), .A4(n5897), .ZN(n5902)
         );
  INV_X1 U7665 ( .A(n5900), .ZN(n5901) );
  OAI21_X1 U7666 ( .B1(n5903), .B2(n5902), .A(n5901), .ZN(n5983) );
  NAND3_X1 U7667 ( .A1(n5905), .A2(n5904), .A3(n7029), .ZN(n5927) );
  INV_X1 U7668 ( .A(n5927), .ZN(n5916) );
  INV_X1 U7669 ( .A(n5925), .ZN(n5913) );
  INV_X1 U7670 ( .A(n7019), .ZN(n5906) );
  AOI21_X1 U7671 ( .B1(n5922), .B2(n5907), .A(n5906), .ZN(n5908) );
  OR2_X1 U7672 ( .A1(n5920), .A2(n5908), .ZN(n5909) );
  OAI211_X1 U7673 ( .C1(n7022), .C2(n4825), .A(n5910), .B(n5909), .ZN(n5912)
         );
  INV_X1 U7674 ( .A(n7024), .ZN(n5911) );
  AOI21_X1 U7675 ( .B1(n5913), .B2(n5912), .A(n5911), .ZN(n5914) );
  INV_X1 U7676 ( .A(n7025), .ZN(n5926) );
  OAI211_X1 U7677 ( .C1(n5914), .C2(n5926), .A(n7028), .B(n7026), .ZN(n5915)
         );
  NAND2_X1 U7678 ( .A1(n5916), .A2(n5915), .ZN(n5979) );
  INV_X1 U7679 ( .A(n5976), .ZN(n5929) );
  AOI22_X1 U7680 ( .A1(n5968), .A2(n5917), .B1(n5919), .B2(n5918), .ZN(n5928)
         );
  INV_X1 U7681 ( .A(n5920), .ZN(n5923) );
  NAND4_X1 U7682 ( .A1(n5923), .A2(n5922), .A3(n8317), .A4(n5921), .ZN(n5924)
         );
  NOR4_X1 U7683 ( .A1(n5927), .A2(n5926), .A3(n5925), .A4(n5924), .ZN(n5982)
         );
  OAI21_X1 U7684 ( .B1(n5929), .B2(n5928), .A(n5982), .ZN(n5933) );
  INV_X1 U7685 ( .A(n5930), .ZN(n5932) );
  NAND2_X1 U7686 ( .A1(n5932), .A2(n5931), .ZN(n5986) );
  AOI21_X1 U7687 ( .B1(n5979), .B2(n5933), .A(n5986), .ZN(n5937) );
  INV_X1 U7688 ( .A(n5934), .ZN(n5936) );
  AOI21_X1 U7689 ( .B1(n5936), .B2(n5935), .A(n9847), .ZN(n5988) );
  OAI21_X1 U7690 ( .B1(n5983), .B2(n5937), .A(n5988), .ZN(n5939) );
  NAND3_X1 U7691 ( .A1(n5939), .A2(n7045), .A3(n7048), .ZN(n5944) );
  NAND2_X1 U7692 ( .A1(n7048), .A2(n7044), .ZN(n5940) );
  NAND3_X1 U7693 ( .A1(n7049), .A2(n5941), .A3(n5940), .ZN(n5942) );
  AOI22_X1 U7694 ( .A1(n5992), .A2(n5942), .B1(n5852), .B2(n10093), .ZN(n5989)
         );
  OAI211_X1 U7695 ( .C1(n5945), .C2(n5944), .A(n5989), .B(n5943), .ZN(n5949)
         );
  AOI211_X1 U7696 ( .C1(n5949), .C2(n5948), .A(n5946), .B(n5947), .ZN(n5950)
         );
  NOR3_X1 U7697 ( .A1(n5951), .A2(n9990), .A3(n5950), .ZN(n5958) );
  OR2_X1 U7698 ( .A1(n7811), .A2(P1_U3084), .ZN(n8332) );
  INV_X1 U7699 ( .A(n8332), .ZN(n5957) );
  INV_X1 U7700 ( .A(P1_B_REG_SCAN_IN), .ZN(n5956) );
  AND2_X1 U7701 ( .A1(n7811), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5952) );
  INV_X1 U7702 ( .A(n7684), .ZN(n7690) );
  NAND2_X1 U7703 ( .A1(n10225), .A2(n7690), .ZN(n7820) );
  XNOR2_X2 U7704 ( .A(n5953), .B(n5954), .ZN(n7993) );
  NAND2_X1 U7705 ( .A1(n7051), .A2(n8059), .ZN(n7719) );
  OR2_X1 U7706 ( .A1(n7619), .A2(n7719), .ZN(n7966) );
  NOR3_X1 U7707 ( .A1(n7820), .A2(n7686), .A3(n7966), .ZN(n5955) );
  AOI211_X1 U7708 ( .C1(n5957), .C2(n8250), .A(n5956), .B(n5955), .ZN(n6001)
         );
  NOR3_X1 U7709 ( .A1(n5958), .A2(n6001), .A3(n7993), .ZN(n5959) );
  OAI211_X1 U7710 ( .C1(n5961), .C2(n8059), .A(n5960), .B(n5959), .ZN(n6008)
         );
  INV_X1 U7711 ( .A(n5963), .ZN(n5964) );
  OAI211_X1 U7712 ( .C1(n8087), .C2(n7153), .A(n4495), .B(n5964), .ZN(n5966)
         );
  NAND2_X1 U7713 ( .A1(n5966), .A2(n5965), .ZN(n5967) );
  OAI22_X1 U7714 ( .A1(n5962), .A2(n5967), .B1(n8925), .B2(n7873), .ZN(n5970)
         );
  INV_X1 U7715 ( .A(n5968), .ZN(n5969) );
  AOI21_X1 U7716 ( .B1(n5971), .B2(n5970), .A(n5969), .ZN(n5978) );
  INV_X1 U7717 ( .A(n7012), .ZN(n5975) );
  OR2_X1 U7718 ( .A1(n5973), .A2(n5972), .ZN(n5974) );
  NAND2_X1 U7719 ( .A1(n5975), .A2(n5974), .ZN(n8067) );
  INV_X1 U7720 ( .A(n8067), .ZN(n5977) );
  OAI21_X1 U7721 ( .B1(n5978), .B2(n5977), .A(n5976), .ZN(n5981) );
  INV_X1 U7722 ( .A(n5979), .ZN(n5980) );
  AOI21_X1 U7723 ( .B1(n5982), .B2(n5981), .A(n5980), .ZN(n5985) );
  INV_X1 U7724 ( .A(n5983), .ZN(n5984) );
  OAI21_X1 U7725 ( .B1(n5986), .B2(n5985), .A(n5984), .ZN(n5987) );
  AOI211_X1 U7726 ( .C1(n5988), .C2(n5987), .A(n7047), .B(n8892), .ZN(n5991)
         );
  INV_X1 U7727 ( .A(n5989), .ZN(n5990) );
  AOI21_X1 U7728 ( .B1(n5992), .B2(n5991), .A(n5990), .ZN(n5997) );
  INV_X1 U7729 ( .A(n5993), .ZN(n5994) );
  OAI211_X1 U7730 ( .C1(n5997), .C2(n5996), .A(n5995), .B(n5994), .ZN(n6000)
         );
  INV_X1 U7731 ( .A(n5998), .ZN(n5999) );
  INV_X1 U7732 ( .A(n6004), .ZN(n6002) );
  INV_X1 U7733 ( .A(n6001), .ZN(n6003) );
  NAND3_X1 U7734 ( .A1(n6002), .A2(n7941), .A3(n6003), .ZN(n6007) );
  NAND2_X1 U7735 ( .A1(n6003), .A2(n8332), .ZN(n6006) );
  NAND4_X1 U7736 ( .A1(n6004), .A2(n9990), .A3(n6003), .A4(n7993), .ZN(n6005)
         );
  AND2_X1 U7737 ( .A1(n6008), .A2(n5030), .ZN(P1_U3240) );
  INV_X1 U7738 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9186) );
  NOR2_X1 U7739 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n6009) );
  INV_X1 U7740 ( .A(n6085), .ZN(n6023) );
  INV_X1 U7741 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6012) );
  NAND2_X1 U7742 ( .A1(n6041), .A2(n6012), .ZN(n6025) );
  INV_X1 U7743 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6013) );
  NAND3_X1 U7744 ( .A1(n6029), .A2(n6026), .A3(n6013), .ZN(n6014) );
  INV_X1 U7745 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6015) );
  INV_X1 U7746 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6885) );
  NAND3_X1 U7747 ( .A1(n6016), .A2(n6015), .A3(n6885), .ZN(n6017) );
  NOR2_X1 U7748 ( .A1(n6048), .A2(n6017), .ZN(n6062) );
  NAND2_X1 U7749 ( .A1(n6062), .A2(n6018), .ZN(n6024) );
  INV_X1 U7750 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6068) );
  INV_X1 U7751 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6019) );
  NAND3_X1 U7752 ( .A1(n6068), .A2(n6065), .A3(n6019), .ZN(n6020) );
  OAI21_X1 U7753 ( .B1(n6024), .B2(n6020), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6021) );
  MUX2_X1 U7754 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6021), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n6022) );
  AND2_X1 U7755 ( .A1(n6023), .A2(n6022), .ZN(n6351) );
  NAND2_X1 U7756 ( .A1(n6024), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6066) );
  XNOR2_X1 U7757 ( .A(n6066), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7482) );
  OAI21_X1 U7758 ( .B1(n6048), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6051) );
  XNOR2_X1 U7759 ( .A(n6051), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7411) );
  NAND2_X1 U7760 ( .A1(n6025), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6046) );
  NAND2_X1 U7761 ( .A1(n6046), .A2(n6026), .ZN(n6027) );
  NAND2_X1 U7762 ( .A1(n6027), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U7763 ( .A1(n6030), .A2(n6029), .ZN(n6032) );
  NAND2_X1 U7764 ( .A1(n6032), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6028) );
  XNOR2_X1 U7765 ( .A(n6028), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7640) );
  OR2_X1 U7766 ( .A1(n6030), .A2(n6029), .ZN(n6031) );
  NAND2_X1 U7767 ( .A1(n6039), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7768 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6035) );
  NAND2_X1 U7769 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n7562) );
  NOR2_X1 U7770 ( .A1(n7561), .A2(n7562), .ZN(n7560) );
  AOI21_X1 U7771 ( .B1(n6132), .B2(P2_REG2_REG_1__SCAN_IN), .A(n7560), .ZN(
        n7573) );
  INV_X1 U7772 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6038) );
  MUX2_X1 U7773 ( .A(n6038), .B(P2_REG2_REG_2__SCAN_IN), .S(n6175), .Z(n7572)
         );
  NOR2_X1 U7774 ( .A1(n7573), .A2(n7572), .ZN(n7571) );
  INV_X1 U7775 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9459) );
  OAI21_X1 U7776 ( .B1(n6039), .B2(P2_IR_REG_2__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6040) );
  MUX2_X1 U7777 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6040), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n6043) );
  INV_X1 U7778 ( .A(n6041), .ZN(n6042) );
  MUX2_X1 U7779 ( .A(n9459), .B(P2_REG2_REG_3__SCAN_IN), .S(n7537), .Z(n7533)
         );
  INV_X1 U7780 ( .A(n7537), .ZN(n6044) );
  XNOR2_X1 U7781 ( .A(n6210), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n7599) );
  XNOR2_X1 U7782 ( .A(n7550), .B(P2_REG2_REG_5__SCAN_IN), .ZN(n7547) );
  NOR2_X1 U7783 ( .A1(n7548), .A2(n7547), .ZN(n7546) );
  INV_X1 U7784 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n8174) );
  MUX2_X1 U7785 ( .A(n8174), .B(P2_REG2_REG_6__SCAN_IN), .S(n7596), .Z(n7592)
         );
  XNOR2_X1 U7786 ( .A(n7640), .B(P2_REG2_REG_7__SCAN_IN), .ZN(n7638) );
  NAND2_X1 U7787 ( .A1(n6048), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6049) );
  XNOR2_X1 U7788 ( .A(n6049), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6267) );
  XNOR2_X1 U7789 ( .A(n6267), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n7858) );
  NOR2_X1 U7790 ( .A1(n7859), .A2(n7858), .ZN(n7857) );
  INV_X1 U7791 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n8550) );
  MUX2_X1 U7792 ( .A(n8550), .B(P2_REG2_REG_9__SCAN_IN), .S(n7411), .Z(n8044)
         );
  NAND2_X1 U7793 ( .A1(n6051), .A2(n6885), .ZN(n6052) );
  NAND2_X1 U7794 ( .A1(n6052), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6054) );
  INV_X1 U7795 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U7796 ( .A1(n6054), .A2(n6053), .ZN(n6057) );
  OR2_X1 U7797 ( .A1(n6054), .A2(n6053), .ZN(n6055) );
  XNOR2_X1 U7798 ( .A(n6280), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n8358) );
  INV_X1 U7799 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6059) );
  NAND2_X1 U7800 ( .A1(n6057), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6058) );
  XNOR2_X1 U7801 ( .A(n6058), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7429) );
  MUX2_X1 U7802 ( .A(n6059), .B(P2_REG2_REG_11__SCAN_IN), .S(n7429), .Z(n6060)
         );
  INV_X1 U7803 ( .A(n6060), .ZN(n8481) );
  OR2_X1 U7804 ( .A1(n7429), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6061) );
  INV_X1 U7805 ( .A(n6062), .ZN(n6063) );
  NAND2_X1 U7806 ( .A1(n6063), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6064) );
  XNOR2_X1 U7807 ( .A(n6064), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7476) );
  XNOR2_X1 U7808 ( .A(n7476), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n8709) );
  INV_X1 U7809 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6309) );
  XNOR2_X1 U7810 ( .A(n7482), .B(n6309), .ZN(n8720) );
  NAND2_X1 U7811 ( .A1(n6066), .A2(n6065), .ZN(n6067) );
  NAND2_X1 U7812 ( .A1(n6067), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7813 ( .A1(n6069), .A2(n6068), .ZN(n6071) );
  OR2_X1 U7814 ( .A1(n6069), .A2(n6068), .ZN(n6070) );
  INV_X1 U7815 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6332) );
  XNOR2_X1 U7816 ( .A(n6326), .B(n6332), .ZN(n9127) );
  INV_X1 U7817 ( .A(n6326), .ZN(n9133) );
  NAND2_X1 U7818 ( .A1(n6071), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6072) );
  XNOR2_X1 U7819 ( .A(n6072), .B(P2_IR_REG_15__SCAN_IN), .ZN(n9146) );
  INV_X1 U7820 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9140) );
  INV_X1 U7821 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n6872) );
  INV_X1 U7822 ( .A(n6351), .ZN(n9155) );
  AOI22_X1 U7823 ( .A1(n6351), .A2(n6872), .B1(P2_REG2_REG_16__SCAN_IN), .B2(
        n9155), .ZN(n9152) );
  NOR2_X1 U7824 ( .A1(n6085), .A2(n6033), .ZN(n6076) );
  MUX2_X1 U7825 ( .A(n6033), .B(n6076), .S(P2_IR_REG_17__SCAN_IN), .Z(n6077)
         );
  INV_X1 U7826 ( .A(n6077), .ZN(n6078) );
  AND2_X1 U7827 ( .A1(n6078), .A2(n6093), .ZN(n6362) );
  NAND2_X1 U7828 ( .A1(n6362), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6079) );
  OAI21_X1 U7829 ( .B1(n6362), .B2(P2_REG2_REG_17__SCAN_IN), .A(n6079), .ZN(
        n9166) );
  NOR2_X1 U7830 ( .A1(n9167), .A2(n9166), .ZN(n9165) );
  NOR2_X1 U7831 ( .A1(n9165), .A2(n6080), .ZN(n6083) );
  NAND2_X1 U7832 ( .A1(n6093), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6081) );
  XNOR2_X1 U7833 ( .A(n6081), .B(P2_IR_REG_18__SCAN_IN), .ZN(n9192) );
  XNOR2_X1 U7834 ( .A(n6083), .B(n6082), .ZN(n9187) );
  NOR2_X1 U7835 ( .A1(n9186), .A2(n9187), .ZN(n9185) );
  NOR2_X1 U7836 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n6084) );
  INV_X1 U7837 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7838 ( .A1(n6087), .A2(n6086), .ZN(n6114) );
  NAND2_X1 U7839 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), 
        .ZN(n6769) );
  NOR2_X1 U7840 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n6092) );
  NOR2_X1 U7841 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n6091) );
  NOR2_X1 U7842 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n6090) );
  NOR2_X1 U7843 ( .A1(n6093), .A2(n6099), .ZN(n6103) );
  NAND2_X1 U7844 ( .A1(n6103), .A2(n6096), .ZN(n6106) );
  NAND2_X1 U7845 ( .A1(n6106), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6094) );
  MUX2_X1 U7846 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6094), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6102) );
  NAND3_X1 U7847 ( .A1(n6097), .A2(n6096), .A3(n6095), .ZN(n6098) );
  NAND2_X1 U7848 ( .A1(n6102), .A2(n6122), .ZN(n8687) );
  INV_X1 U7849 ( .A(n6103), .ZN(n6104) );
  NAND2_X1 U7850 ( .A1(n6104), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6105) );
  MUX2_X1 U7851 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6105), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n6107) );
  NAND2_X1 U7852 ( .A1(n6107), .A2(n6106), .ZN(n8576) );
  NOR2_X1 U7853 ( .A1(n8687), .A2(n8576), .ZN(n6108) );
  NAND2_X1 U7854 ( .A1(n8493), .A2(n6108), .ZN(n6738) );
  NAND2_X1 U7855 ( .A1(n6109), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n6110) );
  NAND2_X1 U7856 ( .A1(n6111), .A2(n6110), .ZN(n6737) );
  NAND2_X1 U7857 ( .A1(n6112), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6113) );
  INV_X1 U7858 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6116) );
  INV_X1 U7860 ( .A(n6728), .ZN(n6121) );
  NOR2_X1 U7861 ( .A1(n6737), .A2(P2_U3152), .ZN(n8273) );
  INV_X1 U7862 ( .A(n8273), .ZN(n7379) );
  NAND2_X1 U7863 ( .A1(n6124), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6118) );
  INV_X1 U7864 ( .A(n6563), .ZN(n6562) );
  NAND2_X1 U7865 ( .A1(n6562), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8716) );
  OR2_X1 U7866 ( .A1(n6738), .A2(n8716), .ZN(n6120) );
  OAI211_X1 U7867 ( .C1(n10472), .C2(n6121), .A(n7379), .B(n6120), .ZN(n6126)
         );
  NAND2_X1 U7868 ( .A1(n6122), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6123) );
  NAND2_X1 U7869 ( .A1(n6126), .A2(n6197), .ZN(n6129) );
  INV_X1 U7870 ( .A(n10487), .ZN(n6127) );
  OR2_X2 U7871 ( .A1(n6738), .A2(n6127), .ZN(n9125) );
  NAND2_X1 U7872 ( .A1(n6129), .A2(n9125), .ZN(n6149) );
  NOR2_X1 U7873 ( .A1(n6563), .A2(n8695), .ZN(n6128) );
  INV_X1 U7874 ( .A(n8695), .ZN(n6749) );
  INV_X1 U7875 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n6877) );
  INV_X1 U7876 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n6369) );
  INV_X1 U7877 ( .A(n6362), .ZN(n9177) );
  XNOR2_X1 U7878 ( .A(n9177), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n9170) );
  OR2_X1 U7879 ( .A1(n6351), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6141) );
  XNOR2_X1 U7880 ( .A(n6351), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n9157) );
  INV_X1 U7881 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10524) );
  INV_X1 U7882 ( .A(n7640), .ZN(n7649) );
  NOR2_X1 U7883 ( .A1(n7649), .A2(n10524), .ZN(n6137) );
  INV_X1 U7884 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6130) );
  MUX2_X1 U7885 ( .A(n6130), .B(P2_REG1_REG_1__SCAN_IN), .S(n7568), .Z(n6131)
         );
  NAND3_X1 U7886 ( .A1(n6131), .A2(P2_REG1_REG_0__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n7576) );
  NAND2_X1 U7887 ( .A1(n6132), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7575) );
  INV_X1 U7888 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7852) );
  INV_X1 U7889 ( .A(n6175), .ZN(n7581) );
  NOR2_X1 U7890 ( .A1(n7581), .A2(n7852), .ZN(n7536) );
  INV_X1 U7891 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6133) );
  MUX2_X1 U7892 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6133), .S(n7537), .Z(n6134)
         );
  NAND2_X1 U7893 ( .A1(n7537), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7603) );
  INV_X1 U7894 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10519) );
  INV_X1 U7895 ( .A(n6210), .ZN(n7611) );
  NOR2_X1 U7896 ( .A1(n7611), .A2(n10519), .ZN(n7549) );
  INV_X1 U7897 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7866) );
  MUX2_X1 U7898 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n7866), .S(n7550), .Z(n6135)
         );
  OAI21_X1 U7899 ( .B1(n7606), .B2(n7549), .A(n6135), .ZN(n7586) );
  NAND2_X1 U7900 ( .A1(n7550), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7585) );
  INV_X1 U7901 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10521) );
  MUX2_X1 U7902 ( .A(n10521), .B(P2_REG1_REG_6__SCAN_IN), .S(n7596), .Z(n7584)
         );
  AOI21_X1 U7903 ( .B1(n7586), .B2(n7585), .A(n7584), .ZN(n7643) );
  INV_X1 U7904 ( .A(n7596), .ZN(n7407) );
  NOR2_X1 U7905 ( .A1(n7407), .A2(n10521), .ZN(n7642) );
  NOR2_X1 U7906 ( .A1(n7643), .A2(n7642), .ZN(n6136) );
  AOI211_X1 U7907 ( .C1(n10524), .C2(n7649), .A(n6137), .B(n6136), .ZN(n7645)
         );
  XNOR2_X1 U7908 ( .A(n6267), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n7853) );
  INV_X1 U7909 ( .A(n6267), .ZN(n7856) );
  INV_X1 U7910 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6828) );
  XOR2_X1 U7911 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n7411), .Z(n8039) );
  XNOR2_X1 U7912 ( .A(n6280), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n8352) );
  INV_X1 U7913 ( .A(n6280), .ZN(n8356) );
  XOR2_X1 U7914 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n7429), .Z(n8484) );
  AOI22_X1 U7915 ( .A1(n8483), .A2(n8484), .B1(n7429), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n8701) );
  NOR2_X1 U7916 ( .A1(n7476), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8722) );
  AOI21_X1 U7917 ( .B1(n7476), .B2(P2_REG1_REG_12__SCAN_IN), .A(n8722), .ZN(
        n8702) );
  OR2_X1 U7918 ( .A1(n7482), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6139) );
  NAND2_X1 U7919 ( .A1(n7482), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6138) );
  AND2_X1 U7920 ( .A1(n6139), .A2(n6138), .ZN(n8721) );
  OAI21_X1 U7921 ( .B1(n8723), .B2(n8722), .A(n8721), .ZN(n8725) );
  NAND2_X1 U7922 ( .A1(n8725), .A2(n6139), .ZN(n9129) );
  XNOR2_X1 U7923 ( .A(n9133), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n9130) );
  NAND2_X1 U7924 ( .A1(n9129), .A2(n9130), .ZN(n9128) );
  INV_X1 U7925 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n6873) );
  NOR2_X1 U7926 ( .A1(n9157), .A2(n9158), .ZN(n9156) );
  INV_X1 U7927 ( .A(n9156), .ZN(n6140) );
  NAND2_X1 U7928 ( .A1(n9170), .A2(n9171), .ZN(n9168) );
  AOI22_X1 U7929 ( .A1(n9192), .A2(n6877), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n6082), .ZN(n9182) );
  NAND2_X1 U7930 ( .A1(n6142), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6143) );
  XNOR2_X1 U7931 ( .A(n6143), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8193) );
  OAI21_X1 U7932 ( .B1(n10472), .B2(n6728), .A(n6197), .ZN(n6145) );
  NAND2_X1 U7933 ( .A1(n10472), .A2(n7379), .ZN(n6144) );
  NAND2_X1 U7934 ( .A1(n6145), .A2(n6144), .ZN(n9190) );
  NAND2_X1 U7935 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8978) );
  INV_X1 U7936 ( .A(n6148), .ZN(n6152) );
  NAND2_X1 U7937 ( .A1(n6149), .A2(n6563), .ZN(n9178) );
  OAI21_X1 U7938 ( .B1(n6150), .B2(n9196), .A(n9178), .ZN(n6151) );
  AOI21_X1 U7939 ( .B1(n6152), .B2(n9163), .A(n6151), .ZN(n6153) );
  NAND2_X1 U7940 ( .A1(n6157), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6156) );
  INV_X1 U7941 ( .A(n6159), .ZN(n9619) );
  OR2_X2 U7942 ( .A1(n6159), .A2(n6033), .ZN(n6161) );
  XNOR2_X2 U7943 ( .A(n6161), .B(n6160), .ZN(n8955) );
  NAND2_X1 U7944 ( .A1(n6555), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6168) );
  XNOR2_X1 U7945 ( .A(n6161), .B(P2_IR_REG_30__SCAN_IN), .ZN(n6162) );
  AND2_X4 U7946 ( .A1(n6163), .A2(n6162), .ZN(n6486) );
  NAND2_X1 U7947 ( .A1(n6486), .A2(n9462), .ZN(n6167) );
  AND2_X4 U7948 ( .A1(n6163), .A2(n8955), .ZN(n6257) );
  NAND2_X1 U7949 ( .A1(n6257), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6166) );
  INV_X1 U7950 ( .A(n8955), .ZN(n6164) );
  NAND4_X1 U7951 ( .A1(n6168), .A2(n6167), .A3(n6166), .A4(n6165), .ZN(n6600)
         );
  NAND2_X1 U7952 ( .A1(n6233), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6169) );
  NAND2_X1 U7953 ( .A1(n6202), .A2(n9460), .ZN(n6526) );
  INV_X1 U7954 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6170) );
  NAND2_X1 U7955 ( .A1(n6486), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U7956 ( .A1(n6257), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6172) );
  NAND2_X1 U7957 ( .A1(n4386), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6171) );
  NAND2_X1 U7958 ( .A1(n4423), .A2(n7384), .ZN(n6178) );
  NAND2_X1 U7959 ( .A1(n6233), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6177) );
  NAND2_X1 U7960 ( .A1(n6382), .A2(n6175), .ZN(n6176) );
  AND3_X2 U7961 ( .A1(n6178), .A2(n6177), .A3(n6176), .ZN(n7847) );
  NAND2_X1 U7962 ( .A1(n4389), .A2(n7847), .ZN(n7199) );
  NAND2_X2 U7963 ( .A1(n7197), .A2(n7199), .ZN(n7841) );
  INV_X1 U7964 ( .A(n7841), .ZN(n7839) );
  NAND2_X1 U7965 ( .A1(n6486), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6183) );
  INV_X1 U7966 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6179) );
  OR2_X1 U7967 ( .A1(n6258), .A2(n6179), .ZN(n6182) );
  NAND2_X1 U7968 ( .A1(n6257), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6181) );
  NAND2_X1 U7969 ( .A1(n7169), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6180) );
  INV_X1 U7970 ( .A(n6198), .ZN(n7740) );
  NAND2_X1 U7971 ( .A1(n4423), .A2(n6184), .ZN(n6187) );
  NAND2_X1 U7972 ( .A1(n6233), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6186) );
  INV_X2 U7973 ( .A(n6586), .ZN(n9468) );
  NAND2_X1 U7974 ( .A1(n6198), .A2(n6586), .ZN(n7353) );
  NAND2_X1 U7975 ( .A1(n7196), .A2(n7353), .ZN(n7668) );
  INV_X1 U7976 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6188) );
  OR2_X1 U7977 ( .A1(n6258), .A2(n6188), .ZN(n6192) );
  NAND2_X1 U7978 ( .A1(n4385), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6191) );
  NAND2_X1 U7979 ( .A1(n6486), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6190) );
  NAND2_X1 U7980 ( .A1(n6257), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6189) );
  NAND2_X1 U7981 ( .A1(n7388), .A2(SI_0_), .ZN(n6194) );
  INV_X1 U7982 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6193) );
  NAND2_X1 U7983 ( .A1(n6194), .A2(n6193), .ZN(n6196) );
  NAND2_X1 U7984 ( .A1(n6196), .A2(n6195), .ZN(n9628) );
  MUX2_X1 U7985 ( .A(n7564), .B(n9628), .S(n6197), .Z(n10463) );
  INV_X1 U7986 ( .A(n10463), .ZN(n10489) );
  NAND2_X1 U7987 ( .A1(n6592), .A2(n10489), .ZN(n7666) );
  NAND2_X1 U7988 ( .A1(n7668), .A2(n7666), .ZN(n7836) );
  NOR2_X1 U7989 ( .A1(n9124), .A2(n9468), .ZN(n7837) );
  NOR2_X1 U7990 ( .A1(n4389), .A2(n8189), .ZN(n6200) );
  NAND2_X1 U7991 ( .A1(n6525), .A2(n7776), .ZN(n7775) );
  NAND2_X1 U7992 ( .A1(n6202), .A2(n7922), .ZN(n6203) );
  NAND2_X1 U7993 ( .A1(n7775), .A2(n6203), .ZN(n9452) );
  NAND2_X1 U7994 ( .A1(n6555), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6209) );
  INV_X1 U7995 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6204) );
  XNOR2_X1 U7996 ( .A(n6204), .B(P2_REG3_REG_3__SCAN_IN), .ZN(n9449) );
  NAND2_X1 U7997 ( .A1(n6486), .A2(n9449), .ZN(n6208) );
  INV_X1 U7998 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6205) );
  OR2_X1 U7999 ( .A1(n6228), .A2(n6205), .ZN(n6207) );
  NAND2_X1 U8000 ( .A1(n6257), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6206) );
  NAND2_X1 U8001 ( .A1(n6382), .A2(n6210), .ZN(n6212) );
  NAND2_X1 U8002 ( .A1(n6233), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6211) );
  NAND2_X1 U8003 ( .A1(n9123), .A2(n10494), .ZN(n7750) );
  INV_X1 U8004 ( .A(n6528), .ZN(n9451) );
  NAND2_X1 U8005 ( .A1(n9452), .A2(n9451), .ZN(n9450) );
  NAND2_X1 U8006 ( .A1(n7923), .A2(n10494), .ZN(n6213) );
  NAND2_X1 U8007 ( .A1(n9450), .A2(n6213), .ZN(n7746) );
  NAND2_X1 U8008 ( .A1(n7401), .A2(n4423), .ZN(n6215) );
  AOI22_X1 U8009 ( .A1(n6233), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6382), .B2(
        n7550), .ZN(n6214) );
  AND2_X2 U8010 ( .A1(n6215), .A2(n6214), .ZN(n8196) );
  NAND2_X1 U8011 ( .A1(n7169), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6223) );
  NAND2_X1 U8012 ( .A1(n6257), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6222) );
  INV_X1 U8013 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U8014 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6216) );
  NAND2_X1 U8015 ( .A1(n6217), .A2(n6216), .ZN(n6218) );
  AND2_X1 U8016 ( .A1(n6226), .A2(n6218), .ZN(n8194) );
  NAND2_X1 U8017 ( .A1(n6486), .A2(n8194), .ZN(n6221) );
  INV_X1 U8018 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6219) );
  NAND2_X1 U8019 ( .A1(n7915), .A2(n8196), .ZN(n8115) );
  NAND2_X1 U8020 ( .A1(n6555), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U8021 ( .A1(n6257), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6231) );
  INV_X1 U8022 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6225) );
  NAND2_X1 U8023 ( .A1(n6226), .A2(n6225), .ZN(n6227) );
  AND2_X1 U8024 ( .A1(n6241), .A2(n6227), .ZN(n8177) );
  NAND2_X1 U8025 ( .A1(n6486), .A2(n8177), .ZN(n6230) );
  OR2_X1 U8026 ( .A1(n6228), .A2(n8174), .ZN(n6229) );
  NAND4_X1 U8027 ( .A1(n6232), .A2(n6231), .A3(n6230), .A4(n6229), .ZN(n9122)
         );
  NAND2_X1 U8028 ( .A1(n7403), .A2(n4423), .ZN(n6235) );
  AOI22_X1 U8029 ( .A1(n4388), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6382), .B2(
        n7596), .ZN(n6234) );
  OR2_X1 U8030 ( .A1(n9122), .A2(n8180), .ZN(n8117) );
  NAND2_X1 U8031 ( .A1(n6236), .A2(n7176), .ZN(n6238) );
  AOI22_X1 U8032 ( .A1(n4387), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6382), .B2(
        n7640), .ZN(n6237) );
  NAND2_X1 U8033 ( .A1(n6555), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6247) );
  INV_X1 U8034 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6240) );
  NAND2_X1 U8035 ( .A1(n6241), .A2(n6240), .ZN(n6242) );
  AND2_X1 U8036 ( .A1(n6270), .A2(n6242), .ZN(n8128) );
  NAND2_X1 U8037 ( .A1(n6486), .A2(n8128), .ZN(n6246) );
  NAND2_X1 U8038 ( .A1(n6257), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6245) );
  INV_X1 U8039 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6243) );
  OR2_X1 U8040 ( .A1(n6558), .A2(n6243), .ZN(n6244) );
  NOR2_X1 U8041 ( .A1(n8126), .A2(n9121), .ZN(n7222) );
  INV_X1 U8042 ( .A(n7222), .ZN(n6248) );
  AND2_X1 U8043 ( .A1(n8117), .A2(n6248), .ZN(n6250) );
  AND2_X1 U8044 ( .A1(n8115), .A2(n6250), .ZN(n6249) );
  INV_X1 U8045 ( .A(n6250), .ZN(n6251) );
  NAND2_X1 U8046 ( .A1(n8180), .A2(n9122), .ZN(n8116) );
  NAND2_X1 U8047 ( .A1(n7219), .A2(n6248), .ZN(n6252) );
  NAND2_X1 U8048 ( .A1(n7169), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6263) );
  NAND2_X1 U8049 ( .A1(n6272), .A2(n6255), .ZN(n6256) );
  AND2_X1 U8050 ( .A1(n6282), .A2(n6256), .ZN(n8552) );
  NAND2_X1 U8051 ( .A1(n6486), .A2(n8552), .ZN(n6262) );
  NAND2_X1 U8052 ( .A1(n6257), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6261) );
  INV_X1 U8053 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n6259) );
  OR2_X1 U8054 ( .A1(n7172), .A2(n6259), .ZN(n6260) );
  INV_X4 U8055 ( .A(n6264), .ZN(n7176) );
  NAND2_X1 U8056 ( .A1(n7410), .A2(n7176), .ZN(n6266) );
  AOI22_X1 U8057 ( .A1(n4388), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6382), .B2(
        n7411), .ZN(n6265) );
  NAND2_X1 U8058 ( .A1(n9587), .A2(n8209), .ZN(n7228) );
  NAND2_X1 U8059 ( .A1(n7421), .A2(n7176), .ZN(n6269) );
  AOI22_X1 U8060 ( .A1(n4387), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6382), .B2(
        n6267), .ZN(n6268) );
  NAND2_X1 U8061 ( .A1(n6269), .A2(n6268), .ZN(n8308) );
  NAND2_X1 U8062 ( .A1(n7169), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6277) );
  INV_X1 U8063 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7987) );
  NAND2_X1 U8064 ( .A1(n6270), .A2(n7987), .ZN(n6271) );
  AND2_X1 U8065 ( .A1(n6272), .A2(n6271), .ZN(n8307) );
  NAND2_X1 U8066 ( .A1(n6486), .A2(n8307), .ZN(n6276) );
  NAND2_X1 U8067 ( .A1(n6257), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6275) );
  INV_X1 U8068 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n6273) );
  OR2_X1 U8069 ( .A1(n7172), .A2(n6273), .ZN(n6274) );
  NAND4_X1 U8070 ( .A1(n6277), .A2(n6276), .A3(n6275), .A4(n6274), .ZN(n9120)
         );
  AND2_X1 U8071 ( .A1(n8308), .A2(n9120), .ZN(n8538) );
  INV_X1 U8072 ( .A(n9120), .ZN(n8545) );
  NAND2_X1 U8073 ( .A1(n8308), .A2(n8545), .ZN(n8541) );
  OR2_X1 U8074 ( .A1(n9587), .A2(n9119), .ZN(n6278) );
  AOI22_X1 U8075 ( .A1(n4388), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6382), .B2(
        n6280), .ZN(n6281) );
  NAND2_X1 U8076 ( .A1(n7169), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6288) );
  NAND2_X1 U8077 ( .A1(n6282), .A2(n8353), .ZN(n6283) );
  AND2_X1 U8078 ( .A1(n6297), .A2(n6283), .ZN(n8214) );
  NAND2_X1 U8079 ( .A1(n6486), .A2(n8214), .ZN(n6287) );
  NAND2_X1 U8080 ( .A1(n6257), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6286) );
  INV_X1 U8081 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n6284) );
  OR2_X1 U8082 ( .A1(n7172), .A2(n6284), .ZN(n6285) );
  NAND4_X1 U8083 ( .A1(n6288), .A2(n6287), .A3(n6286), .A4(n6285), .ZN(n9118)
         );
  INV_X1 U8084 ( .A(n9118), .ZN(n8546) );
  NAND2_X1 U8085 ( .A1(n9580), .A2(n8546), .ZN(n7232) );
  NAND2_X1 U8086 ( .A1(n7233), .A2(n7232), .ZN(n8220) );
  INV_X1 U8087 ( .A(n8220), .ZN(n8218) );
  INV_X1 U8088 ( .A(n6289), .ZN(n8217) );
  AND2_X1 U8089 ( .A1(n8217), .A2(n8220), .ZN(n6290) );
  AOI22_X1 U8090 ( .A1(n4476), .A2(n6290), .B1(n9118), .B2(n9580), .ZN(n6291)
         );
  NAND2_X1 U8091 ( .A1(n7428), .A2(n7176), .ZN(n6294) );
  AOI22_X1 U8092 ( .A1(n4387), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n7429), .B2(
        n6382), .ZN(n6293) );
  OR2_X1 U8093 ( .A1(n6558), .A2(n6059), .ZN(n6302) );
  INV_X1 U8094 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n6296) );
  NAND2_X1 U8095 ( .A1(n6297), .A2(n6296), .ZN(n6298) );
  AND2_X1 U8096 ( .A1(n6317), .A2(n6298), .ZN(n8231) );
  NAND2_X1 U8097 ( .A1(n6486), .A2(n8231), .ZN(n6301) );
  NAND2_X1 U8098 ( .A1(n6257), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6300) );
  INV_X1 U8099 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n6821) );
  OR2_X1 U8100 ( .A1(n7172), .A2(n6821), .ZN(n6299) );
  NAND4_X1 U8101 ( .A1(n6302), .A2(n6301), .A3(n6300), .A4(n6299), .ZN(n9117)
         );
  NOR2_X1 U8102 ( .A1(n9574), .A2(n8655), .ZN(n8650) );
  INV_X1 U8103 ( .A(n8650), .ZN(n7234) );
  NAND2_X1 U8104 ( .A1(n9574), .A2(n8655), .ZN(n8651) );
  NAND2_X1 U8105 ( .A1(n7234), .A2(n8651), .ZN(n8227) );
  NAND2_X1 U8106 ( .A1(n8225), .A2(n8227), .ZN(n8224) );
  NAND2_X1 U8107 ( .A1(n9574), .A2(n9117), .ZN(n6303) );
  NAND2_X1 U8108 ( .A1(n7481), .A2(n7176), .ZN(n6305) );
  AOI22_X1 U8109 ( .A1(n4387), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6382), .B2(
        n7482), .ZN(n6304) );
  NAND2_X1 U8110 ( .A1(n6555), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6313) );
  NAND2_X1 U8111 ( .A1(n6257), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6312) );
  INV_X1 U8112 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6307) );
  NAND2_X1 U8113 ( .A1(n6319), .A2(n6307), .ZN(n6308) );
  AND2_X1 U8114 ( .A1(n6330), .A2(n6308), .ZN(n9431) );
  NAND2_X1 U8115 ( .A1(n6486), .A2(n9431), .ZN(n6311) );
  OR2_X1 U8116 ( .A1(n6558), .A2(n6309), .ZN(n6310) );
  NAND4_X1 U8117 ( .A1(n6313), .A2(n6312), .A3(n6311), .A4(n6310), .ZN(n9115)
         );
  INV_X1 U8118 ( .A(n9115), .ZN(n8656) );
  OR2_X1 U8119 ( .A1(n9565), .A2(n8656), .ZN(n7243) );
  NAND2_X1 U8120 ( .A1(n9565), .A2(n8656), .ZN(n7253) );
  NAND2_X1 U8121 ( .A1(n6314), .A2(n7176), .ZN(n6316) );
  AOI22_X1 U8122 ( .A1(n4388), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6382), .B2(
        n7476), .ZN(n6315) );
  NAND2_X1 U8123 ( .A1(n7169), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6323) );
  INV_X1 U8124 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8703) );
  NAND2_X1 U8125 ( .A1(n6317), .A2(n8703), .ZN(n6318) );
  AND2_X1 U8126 ( .A1(n6319), .A2(n6318), .ZN(n8996) );
  NAND2_X1 U8127 ( .A1(n6486), .A2(n8996), .ZN(n6322) );
  NAND2_X1 U8128 ( .A1(n6257), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6321) );
  INV_X1 U8129 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n6898) );
  OR2_X1 U8130 ( .A1(n7172), .A2(n6898), .ZN(n6320) );
  NAND4_X1 U8131 ( .A1(n6323), .A2(n6322), .A3(n6321), .A4(n6320), .ZN(n9116)
         );
  INV_X1 U8132 ( .A(n9116), .ZN(n9417) );
  NAND2_X1 U8133 ( .A1(n6570), .A2(n9417), .ZN(n7241) );
  NAND2_X1 U8134 ( .A1(n6539), .A2(n7241), .ZN(n8653) );
  NOR2_X1 U8135 ( .A1(n6570), .A2(n9116), .ZN(n9421) );
  OR2_X1 U8136 ( .A1(n8653), .A2(n9421), .ZN(n6324) );
  INV_X1 U8137 ( .A(n9565), .ZN(n9433) );
  OAI22_X1 U8138 ( .A1(n9424), .A2(n6324), .B1(n8656), .B2(n9433), .ZN(n6325)
         );
  INV_X1 U8139 ( .A(n6325), .ZN(n8677) );
  NAND2_X1 U8140 ( .A1(n7512), .A2(n7176), .ZN(n6328) );
  AOI22_X1 U8141 ( .A1(n4387), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6326), .B2(
        n6382), .ZN(n6327) );
  INV_X1 U8142 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8613) );
  NAND2_X1 U8143 ( .A1(n6330), .A2(n8613), .ZN(n6331) );
  NAND2_X1 U8144 ( .A1(n6356), .A2(n6331), .ZN(n8673) );
  OR2_X1 U8145 ( .A1(n8673), .A2(n6561), .ZN(n6336) );
  INV_X1 U8146 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n6924) );
  OR2_X1 U8147 ( .A1(n7172), .A2(n6924), .ZN(n6335) );
  NAND2_X1 U8148 ( .A1(n6257), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6334) );
  OR2_X1 U8149 ( .A1(n6558), .A2(n6332), .ZN(n6333) );
  NAND4_X1 U8150 ( .A1(n6336), .A2(n6335), .A3(n6334), .A4(n6333), .ZN(n9400)
         );
  INV_X1 U8151 ( .A(n9400), .ZN(n9420) );
  NAND2_X1 U8152 ( .A1(n6337), .A2(n9420), .ZN(n7258) );
  OR2_X1 U8153 ( .A1(n9424), .A2(n9421), .ZN(n8678) );
  NAND3_X1 U8154 ( .A1(n8677), .A2(n8680), .A3(n8678), .ZN(n6339) );
  AOI22_X1 U8155 ( .A1(n9146), .A2(n6382), .B1(n4388), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n6347) );
  INV_X1 U8156 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n6823) );
  NAND2_X1 U8157 ( .A1(n7169), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6342) );
  NAND2_X1 U8158 ( .A1(n6257), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6341) );
  OAI211_X1 U8159 ( .C1(n7172), .C2(n6823), .A(n6342), .B(n6341), .ZN(n6343)
         );
  INV_X1 U8160 ( .A(n6343), .ZN(n6345) );
  XNOR2_X1 U8161 ( .A(n6356), .B(P2_REG3_REG_15__SCAN_IN), .ZN(n9406) );
  NAND2_X1 U8162 ( .A1(n9406), .A2(n6486), .ZN(n6344) );
  NAND2_X1 U8163 ( .A1(n6345), .A2(n6344), .ZN(n9381) );
  NAND2_X1 U8164 ( .A1(n6347), .A2(n9381), .ZN(n6346) );
  INV_X1 U8165 ( .A(n6347), .ZN(n6348) );
  INV_X1 U8166 ( .A(n9381), .ZN(n9019) );
  NAND2_X1 U8167 ( .A1(n9556), .A2(n9019), .ZN(n7263) );
  INV_X1 U8168 ( .A(n9409), .ZN(n7363) );
  NOR2_X1 U8169 ( .A1(n9556), .A2(n9381), .ZN(n6350) );
  AOI22_X1 U8170 ( .A1(n7177), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6382), .B2(
        n6351), .ZN(n6352) );
  INV_X1 U8171 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n6360) );
  INV_X1 U8172 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6354) );
  INV_X1 U8173 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6353) );
  OAI21_X1 U8174 ( .B1(n6356), .B2(n6354), .A(n6353), .ZN(n6357) );
  NAND2_X1 U8175 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_REG3_REG_15__SCAN_IN), 
        .ZN(n6355) );
  AND2_X1 U8176 ( .A1(n6357), .A2(n6365), .ZN(n9391) );
  NAND2_X1 U8177 ( .A1(n9391), .A2(n6486), .ZN(n6359) );
  AOI22_X1 U8178 ( .A1(n7169), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n6555), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n6358) );
  OAI211_X1 U8179 ( .C1(n6489), .C2(n6360), .A(n6359), .B(n6358), .ZN(n9401)
         );
  INV_X1 U8180 ( .A(n9401), .ZN(n9105) );
  AND2_X1 U8181 ( .A1(n9392), .A2(n9105), .ZN(n7269) );
  INV_X1 U8182 ( .A(n7269), .ZN(n6361) );
  NAND2_X1 U8183 ( .A1(n9379), .A2(n9378), .ZN(n9366) );
  NAND2_X1 U8184 ( .A1(n7832), .A2(n7176), .ZN(n6364) );
  AOI22_X1 U8185 ( .A1(n7177), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6382), .B2(
        n6362), .ZN(n6363) );
  INV_X1 U8186 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9172) );
  NAND2_X1 U8187 ( .A1(n6365), .A2(n9172), .ZN(n6366) );
  NAND2_X1 U8188 ( .A1(n6375), .A2(n6366), .ZN(n9362) );
  OR2_X1 U8189 ( .A1(n9362), .A2(n6561), .ZN(n6368) );
  AOI22_X1 U8190 ( .A1(n7169), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n6555), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n6367) );
  OAI211_X1 U8191 ( .C1(n6489), .C2(n6369), .A(n6368), .B(n6367), .ZN(n9382)
         );
  INV_X1 U8192 ( .A(n9382), .ZN(n6370) );
  NAND2_X1 U8193 ( .A1(n9545), .A2(n6370), .ZN(n7275) );
  NAND2_X1 U8194 ( .A1(n9392), .A2(n9401), .ZN(n9367) );
  OR2_X1 U8195 ( .A1(n9545), .A2(n9382), .ZN(n6371) );
  NAND2_X1 U8196 ( .A1(n7879), .A2(n7176), .ZN(n6373) );
  AOI22_X1 U8197 ( .A1(n7177), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6382), .B2(
        n9192), .ZN(n6372) );
  INV_X1 U8198 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n6374) );
  NAND2_X1 U8199 ( .A1(n6375), .A2(n6374), .ZN(n6376) );
  AND2_X1 U8200 ( .A1(n6387), .A2(n6376), .ZN(n9349) );
  NAND2_X1 U8201 ( .A1(n9349), .A2(n6486), .ZN(n6381) );
  NAND2_X1 U8202 ( .A1(n6555), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6378) );
  NAND2_X1 U8203 ( .A1(n4386), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6377) );
  OAI211_X1 U8204 ( .C1(n6877), .C2(n6489), .A(n6378), .B(n6377), .ZN(n6379)
         );
  INV_X1 U8205 ( .A(n6379), .ZN(n6380) );
  NAND2_X1 U8206 ( .A1(n6381), .A2(n6380), .ZN(n9359) );
  INV_X1 U8207 ( .A(n9359), .ZN(n9026) );
  INV_X1 U8208 ( .A(n9539), .ZN(n9351) );
  NAND2_X1 U8209 ( .A1(n7883), .A2(n7176), .ZN(n6384) );
  AOI22_X1 U8210 ( .A1(n4388), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6382), .B2(
        n8193), .ZN(n6383) );
  INV_X1 U8211 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6386) );
  NAND2_X1 U8212 ( .A1(n6387), .A2(n6386), .ZN(n6388) );
  NAND2_X1 U8213 ( .A1(n6404), .A2(n6388), .ZN(n9335) );
  OR2_X1 U8214 ( .A1(n9335), .A2(n6561), .ZN(n6394) );
  INV_X1 U8215 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n6391) );
  NAND2_X1 U8216 ( .A1(n6555), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6390) );
  NAND2_X1 U8217 ( .A1(n7169), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6389) );
  OAI211_X1 U8218 ( .C1(n6489), .C2(n6391), .A(n6390), .B(n6389), .ZN(n6392)
         );
  INV_X1 U8219 ( .A(n6392), .ZN(n6393) );
  NAND2_X1 U8220 ( .A1(n6394), .A2(n6393), .ZN(n9346) );
  NAND2_X1 U8221 ( .A1(n7979), .A2(n7176), .ZN(n6396) );
  NAND2_X1 U8222 ( .A1(n7177), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6395) );
  XNOR2_X1 U8223 ( .A(n6404), .B(P2_REG3_REG_20__SCAN_IN), .ZN(n9318) );
  INV_X1 U8224 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n6399) );
  NAND2_X1 U8225 ( .A1(n7169), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6398) );
  NAND2_X1 U8226 ( .A1(n6555), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6397) );
  OAI211_X1 U8227 ( .C1(n6399), .C2(n6489), .A(n6398), .B(n6397), .ZN(n6400)
         );
  AOI21_X1 U8228 ( .B1(n9318), .B2(n6486), .A(n6400), .ZN(n8987) );
  NAND2_X1 U8229 ( .A1(n9528), .A2(n8987), .ZN(n7281) );
  INV_X1 U8230 ( .A(n8987), .ZN(n9328) );
  NAND2_X1 U8231 ( .A1(n7996), .A2(n7176), .ZN(n6402) );
  NAND2_X1 U8232 ( .A1(n7177), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6401) );
  INV_X1 U8233 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9056) );
  INV_X1 U8234 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8985) );
  OAI21_X1 U8235 ( .B1(n6404), .B2(n9056), .A(n8985), .ZN(n6405) );
  NAND2_X1 U8236 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_REG3_REG_20__SCAN_IN), 
        .ZN(n6403) );
  AND2_X1 U8237 ( .A1(n6405), .A2(n6414), .ZN(n9303) );
  NAND2_X1 U8238 ( .A1(n9303), .A2(n6486), .ZN(n6411) );
  INV_X1 U8239 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n6408) );
  NAND2_X1 U8240 ( .A1(n6257), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6407) );
  NAND2_X1 U8241 ( .A1(n4386), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6406) );
  OAI211_X1 U8242 ( .C1(n7172), .C2(n6408), .A(n6407), .B(n6406), .ZN(n6409)
         );
  INV_X1 U8243 ( .A(n6409), .ZN(n6410) );
  NAND2_X1 U8244 ( .A1(n6411), .A2(n6410), .ZN(n9314) );
  INV_X1 U8245 ( .A(n9314), .ZN(n9071) );
  NAND2_X1 U8246 ( .A1(n6573), .A2(n9071), .ZN(n6412) );
  NAND2_X1 U8247 ( .A1(n6413), .A2(n7176), .ZN(n6424) );
  INV_X1 U8248 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9069) );
  NAND2_X1 U8249 ( .A1(n6414), .A2(n9069), .ZN(n6415) );
  NAND2_X1 U8250 ( .A1(n6428), .A2(n6415), .ZN(n9289) );
  OR2_X1 U8251 ( .A1(n9289), .A2(n6561), .ZN(n6421) );
  INV_X1 U8252 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n6418) );
  NAND2_X1 U8253 ( .A1(n6555), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6417) );
  NAND2_X1 U8254 ( .A1(n4386), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6416) );
  OAI211_X1 U8255 ( .C1(n6418), .C2(n6489), .A(n6417), .B(n6416), .ZN(n6419)
         );
  INV_X1 U8256 ( .A(n6419), .ZN(n6420) );
  NAND2_X1 U8257 ( .A1(n7177), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6423) );
  AND2_X1 U8258 ( .A1(n4390), .A2(n6423), .ZN(n6422) );
  NAND2_X1 U8259 ( .A1(n9520), .A2(n9264), .ZN(n7291) );
  INV_X1 U8260 ( .A(n9520), .ZN(n6425) );
  AOI22_X2 U8261 ( .A1(n9276), .A2(n6549), .B1(n6425), .B2(n9264), .ZN(n9259)
         );
  NAND2_X1 U8262 ( .A1(n8331), .A2(n7176), .ZN(n6427) );
  NAND2_X1 U8263 ( .A1(n4387), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6426) );
  INV_X1 U8264 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8969) );
  NAND2_X1 U8265 ( .A1(n6428), .A2(n8969), .ZN(n6429) );
  NAND2_X1 U8266 ( .A1(n6438), .A2(n6429), .ZN(n9269) );
  OR2_X1 U8267 ( .A1(n9269), .A2(n6561), .ZN(n6435) );
  INV_X1 U8268 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n6432) );
  NAND2_X1 U8269 ( .A1(n7169), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6431) );
  NAND2_X1 U8270 ( .A1(n6555), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6430) );
  OAI211_X1 U8271 ( .C1(n6432), .C2(n6489), .A(n6431), .B(n6430), .ZN(n6433)
         );
  INV_X1 U8272 ( .A(n6433), .ZN(n6434) );
  NAND2_X1 U8273 ( .A1(n6435), .A2(n6434), .ZN(n9282) );
  OR2_X1 U8274 ( .A1(n9515), .A2(n9070), .ZN(n7295) );
  NAND2_X1 U8275 ( .A1(n9515), .A2(n9070), .ZN(n7294) );
  NAND2_X1 U8276 ( .A1(n8477), .A2(n7176), .ZN(n6437) );
  NAND2_X1 U8277 ( .A1(n4388), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6436) );
  INV_X1 U8278 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9038) );
  OR2_X2 U8279 ( .A1(n6438), .A2(n9038), .ZN(n6460) );
  NAND2_X1 U8280 ( .A1(n6438), .A2(n9038), .ZN(n6439) );
  AND2_X1 U8281 ( .A1(n6460), .A2(n6439), .ZN(n9246) );
  NAND2_X1 U8282 ( .A1(n9246), .A2(n6486), .ZN(n6445) );
  INV_X1 U8283 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n6442) );
  NAND2_X1 U8284 ( .A1(n6555), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6441) );
  NAND2_X1 U8285 ( .A1(n4386), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6440) );
  OAI211_X1 U8286 ( .C1(n6489), .C2(n6442), .A(n6441), .B(n6440), .ZN(n6443)
         );
  INV_X1 U8287 ( .A(n6443), .ZN(n6444) );
  NAND2_X1 U8288 ( .A1(n8573), .A2(n7176), .ZN(n6448) );
  NAND2_X1 U8289 ( .A1(n4387), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6447) );
  XNOR2_X1 U8290 ( .A(n6460), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n9236) );
  NAND2_X1 U8291 ( .A1(n9236), .A2(n6486), .ZN(n6453) );
  INV_X1 U8292 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n6895) );
  NAND2_X1 U8293 ( .A1(n6257), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6450) );
  NAND2_X1 U8294 ( .A1(n6555), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6449) );
  OAI211_X1 U8295 ( .C1(n6558), .C2(n6895), .A(n6450), .B(n6449), .ZN(n6451)
         );
  INV_X1 U8296 ( .A(n6451), .ZN(n6452) );
  NAND2_X1 U8297 ( .A1(n9237), .A2(n9039), .ZN(n7301) );
  NAND2_X1 U8298 ( .A1(n9232), .A2(n6454), .ZN(n9215) );
  NAND2_X1 U8299 ( .A1(n8685), .A2(n7176), .ZN(n6456) );
  NAND2_X1 U8300 ( .A1(n7177), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6455) );
  AND2_X1 U8301 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG3_REG_26__SCAN_IN), 
        .ZN(n6457) );
  INV_X1 U8302 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9003) );
  INV_X1 U8303 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6459) );
  OAI21_X1 U8304 ( .B1(n6460), .B2(n9003), .A(n6459), .ZN(n6461) );
  NAND2_X1 U8305 ( .A1(n6475), .A2(n6461), .ZN(n9224) );
  INV_X1 U8306 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n6464) );
  NAND2_X1 U8307 ( .A1(n6257), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6463) );
  NAND2_X1 U8308 ( .A1(n6555), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6462) );
  OAI211_X1 U8309 ( .C1(n6558), .C2(n6464), .A(n6463), .B(n6462), .ZN(n6465)
         );
  INV_X1 U8310 ( .A(n6465), .ZN(n6466) );
  NAND2_X2 U8311 ( .A1(n6467), .A2(n6466), .ZN(n9203) );
  NAND2_X1 U8312 ( .A1(n9215), .A2(n9214), .ZN(n9213) );
  NAND2_X1 U8313 ( .A1(n6469), .A2(n6468), .ZN(n6470) );
  NAND2_X1 U8314 ( .A1(n7177), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6471) );
  INV_X1 U8315 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6474) );
  NAND2_X1 U8316 ( .A1(n6475), .A2(n6474), .ZN(n6476) );
  NAND2_X1 U8317 ( .A1(n6484), .A2(n6476), .ZN(n8964) );
  INV_X1 U8318 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n6479) );
  NAND2_X1 U8319 ( .A1(n6555), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6478) );
  NAND2_X1 U8320 ( .A1(n6257), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6477) );
  OAI211_X1 U8321 ( .C1(n6479), .C2(n6558), .A(n6478), .B(n6477), .ZN(n6480)
         );
  INV_X1 U8322 ( .A(n6480), .ZN(n6481) );
  XNOR2_X2 U8323 ( .A(n9493), .B(n7315), .ZN(n9209) );
  NAND2_X1 U8324 ( .A1(n7177), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6494) );
  INV_X1 U8325 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6483) );
  NAND2_X1 U8326 ( .A1(n6484), .A2(n6483), .ZN(n6485) );
  NAND2_X1 U8327 ( .A1(n6740), .A2(n6486), .ZN(n6493) );
  INV_X1 U8328 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6490) );
  NAND2_X1 U8329 ( .A1(n4386), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6488) );
  NAND2_X1 U8330 ( .A1(n6555), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6487) );
  OAI211_X1 U8331 ( .C1(n6490), .C2(n6489), .A(n6488), .B(n6487), .ZN(n6491)
         );
  INV_X1 U8332 ( .A(n6491), .ZN(n6492) );
  NAND2_X2 U8333 ( .A1(n6493), .A2(n6492), .ZN(n9204) );
  NAND3_X1 U8334 ( .A1(n6495), .A2(n6494), .A3(n9204), .ZN(n7317) );
  INV_X1 U8335 ( .A(n9204), .ZN(n6496) );
  NAND2_X1 U8336 ( .A1(n9488), .A2(n6496), .ZN(n7320) );
  INV_X1 U8337 ( .A(P2_B_REG_SCAN_IN), .ZN(n6498) );
  XNOR2_X1 U8338 ( .A(n8493), .B(n6498), .ZN(n6499) );
  NAND2_X1 U8339 ( .A1(n6499), .A2(n8576), .ZN(n6500) );
  INV_X1 U8340 ( .A(n8687), .ZN(n6516) );
  NOR4_X1 U8341 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6504) );
  NOR4_X1 U8342 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6503) );
  INV_X1 U8343 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n10480) );
  INV_X1 U8344 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n10478) );
  INV_X1 U8345 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n10475) );
  INV_X1 U8346 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n10476) );
  NAND4_X1 U8347 ( .A1(n10480), .A2(n10478), .A3(n10475), .A4(n10476), .ZN(
        n6501) );
  NOR2_X1 U8348 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n6501), .ZN(n6771) );
  NOR4_X1 U8349 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n6502) );
  AND4_X1 U8350 ( .A1(n6504), .A2(n6503), .A3(n6771), .A4(n6502), .ZN(n6509)
         );
  NOR4_X1 U8351 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n6507) );
  NOR4_X1 U8352 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n6506) );
  NOR4_X1 U8353 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n6505) );
  INV_X1 U8354 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n10473) );
  AND4_X1 U8355 ( .A1(n6507), .A2(n6506), .A3(n6505), .A4(n10473), .ZN(n6508)
         );
  NAND2_X1 U8356 ( .A1(n6509), .A2(n6508), .ZN(n6510) );
  NAND2_X1 U8357 ( .A1(n6511), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6513) );
  NAND2_X1 U8358 ( .A1(n7981), .A2(n4944), .ZN(n7378) );
  INV_X1 U8359 ( .A(n7378), .ZN(n6733) );
  NOR2_X1 U8360 ( .A1(n6728), .A2(n6733), .ZN(n6735) );
  INV_X1 U8361 ( .A(n6759), .ZN(n6520) );
  INV_X1 U8362 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10485) );
  NAND2_X1 U8363 ( .A1(n10471), .A2(n10485), .ZN(n6515) );
  AND2_X1 U8364 ( .A1(n8687), .A2(n8576), .ZN(n10486) );
  INV_X1 U8365 ( .A(n10486), .ZN(n6514) );
  NAND2_X1 U8366 ( .A1(n6515), .A2(n6514), .ZN(n6757) );
  INV_X1 U8367 ( .A(n6757), .ZN(n6519) );
  INV_X1 U8368 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10482) );
  NAND2_X1 U8369 ( .A1(n10471), .A2(n10482), .ZN(n6518) );
  NOR2_X1 U8370 ( .A1(n8493), .A2(n6516), .ZN(n10483) );
  INV_X1 U8371 ( .A(n10483), .ZN(n6517) );
  NAND3_X1 U8372 ( .A1(n6520), .A2(n6519), .A3(n7674), .ZN(n6577) );
  AND2_X1 U8373 ( .A1(n7981), .A2(n8193), .ZN(n6521) );
  NAND2_X1 U8374 ( .A1(n9552), .A2(n7998), .ZN(n6756) );
  XNOR2_X1 U8375 ( .A(n6553), .B(n6585), .ZN(n6522) );
  NAND2_X1 U8376 ( .A1(n6522), .A2(n4944), .ZN(n9425) );
  INV_X1 U8377 ( .A(n6585), .ZN(n6523) );
  NAND2_X1 U8378 ( .A1(n6523), .A2(n8193), .ZN(n8304) );
  AND2_X1 U8379 ( .A1(n9425), .A2(n8304), .ZN(n6524) );
  NOR2_X1 U8380 ( .A1(n9491), .A2(n9411), .ZN(n6583) );
  NAND2_X1 U8381 ( .A1(n7352), .A2(n7353), .ZN(n7842) );
  OAI21_X2 U8382 ( .B1(n7842), .B2(n7841), .A(n7197), .ZN(n7778) );
  INV_X1 U8383 ( .A(n6526), .ZN(n7192) );
  AND2_X1 U8384 ( .A1(n6530), .A2(n6528), .ZN(n6529) );
  NAND2_X1 U8385 ( .A1(n9442), .A2(n6529), .ZN(n6534) );
  INV_X1 U8386 ( .A(n6530), .ZN(n6532) );
  AND2_X1 U8387 ( .A1(n7750), .A2(n7213), .ZN(n6531) );
  NAND2_X1 U8388 ( .A1(n8180), .A2(n7218), .ZN(n7193) );
  NAND2_X1 U8389 ( .A1(n8172), .A2(n7193), .ZN(n8120) );
  INV_X1 U8390 ( .A(n9121), .ZN(n7988) );
  OR2_X1 U8391 ( .A1(n8126), .A2(n7988), .ZN(n8295) );
  NAND2_X1 U8392 ( .A1(n7225), .A2(n8295), .ZN(n8203) );
  INV_X1 U8393 ( .A(n7235), .ZN(n8206) );
  NOR2_X1 U8394 ( .A1(n8203), .A2(n8206), .ZN(n6535) );
  NAND2_X1 U8395 ( .A1(n8120), .A2(n6535), .ZN(n6538) );
  NAND3_X1 U8396 ( .A1(n7225), .A2(n7988), .A3(n8126), .ZN(n6536) );
  NAND3_X1 U8397 ( .A1(n6536), .A2(n7228), .A3(n8541), .ZN(n8204) );
  AOI21_X1 U8398 ( .B1(n8204), .B2(n7235), .A(n8220), .ZN(n6537) );
  NAND2_X1 U8399 ( .A1(n6538), .A2(n6537), .ZN(n8211) );
  NAND2_X1 U8400 ( .A1(n8211), .A2(n7233), .ZN(n8226) );
  INV_X1 U8401 ( .A(n6539), .ZN(n7252) );
  OR2_X1 U8402 ( .A1(n8650), .A2(n7252), .ZN(n6543) );
  INV_X1 U8403 ( .A(n8651), .ZN(n6540) );
  NOR2_X1 U8404 ( .A1(n6540), .A2(n8653), .ZN(n6541) );
  OR2_X1 U8405 ( .A1(n7252), .A2(n6541), .ZN(n6542) );
  OAI21_X1 U8406 ( .B1(n8226), .B2(n6543), .A(n6542), .ZN(n9416) );
  NAND2_X1 U8407 ( .A1(n9398), .A2(n9409), .ZN(n9399) );
  AND2_X1 U8408 ( .A1(n7275), .A2(n7274), .ZN(n9371) );
  INV_X1 U8409 ( .A(n7274), .ZN(n6545) );
  OR2_X1 U8410 ( .A1(n9539), .A2(n9026), .ZN(n7279) );
  NAND2_X1 U8411 ( .A1(n9539), .A2(n9026), .ZN(n7287) );
  NAND2_X1 U8412 ( .A1(n9344), .A2(n7287), .ZN(n9277) );
  INV_X1 U8413 ( .A(n9346), .ZN(n9080) );
  OR2_X1 U8414 ( .A1(n9535), .A2(n9080), .ZN(n7286) );
  AND2_X1 U8415 ( .A1(n9278), .A2(n7286), .ZN(n7283) );
  OR2_X1 U8416 ( .A1(n9523), .A2(n9071), .ZN(n7349) );
  AND2_X1 U8417 ( .A1(n7283), .A2(n7349), .ZN(n6546) );
  NAND2_X1 U8418 ( .A1(n9277), .A2(n6546), .ZN(n6551) );
  NAND2_X1 U8419 ( .A1(n9535), .A2(n9080), .ZN(n7350) );
  NAND2_X1 U8420 ( .A1(n7281), .A2(n7350), .ZN(n7289) );
  NAND3_X1 U8421 ( .A1(n7349), .A2(n9278), .A3(n7289), .ZN(n6547) );
  INV_X1 U8422 ( .A(n7294), .ZN(n6552) );
  NAND2_X1 U8423 ( .A1(n9251), .A2(n9250), .ZN(n9249) );
  NAND2_X1 U8424 ( .A1(n9248), .A2(n9114), .ZN(n7297) );
  OR2_X1 U8425 ( .A1(n9493), .A2(n7315), .ZN(n7318) );
  XNOR2_X1 U8426 ( .A(n7164), .B(n7369), .ZN(n6567) );
  INV_X1 U8427 ( .A(n7981), .ZN(n7355) );
  NAND2_X1 U8428 ( .A1(n6554), .A2(n7355), .ZN(n7184) );
  NAND2_X1 U8429 ( .A1(n6584), .A2(n7184), .ZN(n9385) );
  INV_X1 U8430 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8919) );
  NAND2_X1 U8431 ( .A1(n6257), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6557) );
  NAND2_X1 U8432 ( .A1(n6555), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6556) );
  OAI211_X1 U8433 ( .C1(n6558), .C2(n8919), .A(n6557), .B(n6556), .ZN(n6559)
         );
  INV_X1 U8434 ( .A(n6559), .ZN(n6560) );
  OAI21_X1 U8435 ( .B1(n8918), .B2(n6561), .A(n6560), .ZN(n9113) );
  OR2_X1 U8436 ( .A1(n6728), .A2(n6563), .ZN(n9418) );
  INV_X1 U8437 ( .A(n8308), .ZN(n8364) );
  INV_X1 U8438 ( .A(n8305), .ZN(n6569) );
  INV_X1 U8439 ( .A(n9574), .ZN(n8233) );
  NOR2_X2 U8440 ( .A1(n9430), .A2(n9565), .ZN(n9429) );
  INV_X1 U8441 ( .A(n6337), .ZN(n8676) );
  INV_X1 U8442 ( .A(n9556), .ZN(n9408) );
  NAND2_X1 U8443 ( .A1(n8671), .A2(n9408), .ZN(n9388) );
  INV_X1 U8444 ( .A(n9535), .ZN(n9338) );
  AND2_X2 U8445 ( .A1(n9244), .A2(n9248), .ZN(n9234) );
  NAND2_X2 U8446 ( .A1(n4384), .A2(n7998), .ZN(n7187) );
  INV_X1 U8447 ( .A(n8916), .ZN(n6576) );
  AOI211_X1 U8448 ( .C1(n9488), .C2(n6575), .A(n10508), .B(n6576), .ZN(n9487)
         );
  OR2_X1 U8449 ( .A1(n6577), .A2(n8193), .ZN(n8185) );
  INV_X1 U8450 ( .A(n8185), .ZN(n9472) );
  INV_X1 U8451 ( .A(n9488), .ZN(n6730) );
  NOR2_X1 U8452 ( .A1(n7187), .A2(n7981), .ZN(n6722) );
  INV_X1 U8453 ( .A(n6722), .ZN(n6578) );
  AOI22_X1 U8454 ( .A1(n6740), .A2(n10462), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n10470), .ZN(n6579) );
  OAI21_X1 U8455 ( .B1(n6730), .B2(n10464), .A(n6579), .ZN(n6580) );
  AOI21_X1 U8456 ( .B1(n9487), .B2(n9472), .A(n6580), .ZN(n6581) );
  OAI21_X1 U8457 ( .B1(n9490), .B2(n10470), .A(n6581), .ZN(n6582) );
  OR2_X1 U8458 ( .A1(n6583), .A2(n6582), .ZN(P2_U3268) );
  BUF_X4 U8459 ( .A(n6594), .Z(n6719) );
  NAND2_X1 U8460 ( .A1(n9401), .A2(n6670), .ZN(n6671) );
  INV_X1 U8461 ( .A(n6671), .ZN(n6676) );
  XNOR2_X1 U8462 ( .A(n9392), .B(n6719), .ZN(n6675) );
  XNOR2_X1 U8463 ( .A(n6594), .B(n6586), .ZN(n6590) );
  INV_X1 U8464 ( .A(n6590), .ZN(n6588) );
  NAND2_X1 U8465 ( .A1(n9124), .A2(n6591), .ZN(n6589) );
  INV_X1 U8466 ( .A(n6589), .ZN(n6587) );
  NAND2_X1 U8467 ( .A1(n6588), .A2(n6587), .ZN(n7766) );
  NAND2_X1 U8468 ( .A1(n6590), .A2(n6589), .ZN(n7765) );
  NAND2_X1 U8469 ( .A1(n6592), .A2(n6591), .ZN(n6593) );
  NAND3_X1 U8470 ( .A1(n7766), .A2(n7765), .A3(n7768), .ZN(n7767) );
  NAND2_X1 U8471 ( .A1(n7767), .A2(n7765), .ZN(n7737) );
  XNOR2_X1 U8472 ( .A(n6594), .B(n7847), .ZN(n6595) );
  NAND2_X1 U8473 ( .A1(n4389), .A2(n6591), .ZN(n6596) );
  XNOR2_X1 U8474 ( .A(n6595), .B(n6596), .ZN(n7738) );
  INV_X1 U8475 ( .A(n6595), .ZN(n6598) );
  INV_X1 U8476 ( .A(n6596), .ZN(n6597) );
  NAND2_X1 U8477 ( .A1(n6598), .A2(n6597), .ZN(n6599) );
  XNOR2_X1 U8478 ( .A(n6719), .B(n9460), .ZN(n6603) );
  NAND2_X1 U8479 ( .A1(n9445), .A2(n6591), .ZN(n6601) );
  XNOR2_X1 U8480 ( .A(n6603), .B(n6601), .ZN(n7920) );
  INV_X1 U8481 ( .A(n6601), .ZN(n6602) );
  AND2_X1 U8482 ( .A1(n6603), .A2(n6602), .ZN(n6604) );
  AOI21_X1 U8483 ( .B1(n7921), .B2(n7920), .A(n6604), .ZN(n9047) );
  XNOR2_X1 U8484 ( .A(n6719), .B(n10494), .ZN(n6605) );
  NAND2_X1 U8485 ( .A1(n9123), .A2(n6670), .ZN(n6606) );
  NAND2_X1 U8486 ( .A1(n6605), .A2(n6606), .ZN(n7707) );
  INV_X1 U8487 ( .A(n6605), .ZN(n6608) );
  INV_X1 U8488 ( .A(n6606), .ZN(n6607) );
  NAND2_X1 U8489 ( .A1(n6608), .A2(n6607), .ZN(n6609) );
  AND2_X1 U8490 ( .A1(n7707), .A2(n6609), .ZN(n9046) );
  XNOR2_X1 U8491 ( .A(n6719), .B(n8196), .ZN(n6612) );
  NAND2_X1 U8492 ( .A1(n9443), .A2(n6670), .ZN(n6613) );
  XNOR2_X1 U8493 ( .A(n6612), .B(n6613), .ZN(n7709) );
  INV_X1 U8494 ( .A(n7707), .ZN(n6610) );
  NOR2_X1 U8495 ( .A1(n7709), .A2(n6610), .ZN(n6611) );
  INV_X1 U8496 ( .A(n6612), .ZN(n6615) );
  INV_X1 U8497 ( .A(n6613), .ZN(n6614) );
  NAND2_X1 U8498 ( .A1(n6615), .A2(n6614), .ZN(n6616) );
  INV_X2 U8499 ( .A(n6719), .ZN(n6715) );
  XNOR2_X1 U8500 ( .A(n8180), .B(n6715), .ZN(n6617) );
  NAND2_X1 U8501 ( .A1(n9122), .A2(n6670), .ZN(n6618) );
  NAND2_X1 U8502 ( .A1(n6617), .A2(n6618), .ZN(n6623) );
  INV_X1 U8503 ( .A(n6617), .ZN(n6620) );
  INV_X1 U8504 ( .A(n6618), .ZN(n6619) );
  NAND2_X1 U8505 ( .A1(n6620), .A2(n6619), .ZN(n6621) );
  INV_X1 U8506 ( .A(n7913), .ZN(n6622) );
  NAND2_X1 U8507 ( .A1(n7910), .A2(n6623), .ZN(n7904) );
  XNOR2_X1 U8508 ( .A(n8126), .B(n6715), .ZN(n6625) );
  NAND2_X1 U8509 ( .A1(n9121), .A2(n6670), .ZN(n6624) );
  XNOR2_X1 U8510 ( .A(n6625), .B(n6624), .ZN(n7903) );
  XNOR2_X1 U8511 ( .A(n8308), .B(n6719), .ZN(n6637) );
  NAND2_X1 U8512 ( .A1(n9120), .A2(n6670), .ZN(n6635) );
  XNOR2_X1 U8513 ( .A(n6637), .B(n6635), .ZN(n8145) );
  XNOR2_X1 U8514 ( .A(n9580), .B(n6715), .ZN(n6629) );
  INV_X1 U8515 ( .A(n6629), .ZN(n6627) );
  NAND2_X1 U8516 ( .A1(n9118), .A2(n6670), .ZN(n6628) );
  INV_X1 U8517 ( .A(n6628), .ZN(n6626) );
  NAND2_X1 U8518 ( .A1(n6627), .A2(n6626), .ZN(n6644) );
  INV_X1 U8519 ( .A(n6644), .ZN(n6632) );
  XNOR2_X1 U8520 ( .A(n6629), .B(n6628), .ZN(n8159) );
  INV_X1 U8521 ( .A(n8159), .ZN(n6630) );
  XNOR2_X1 U8522 ( .A(n9587), .B(n6715), .ZN(n6638) );
  NAND2_X1 U8523 ( .A1(n9119), .A2(n6670), .ZN(n6639) );
  NAND2_X1 U8524 ( .A1(n6638), .A2(n6639), .ZN(n8157) );
  AND2_X1 U8525 ( .A1(n6630), .A2(n8157), .ZN(n6631) );
  AND2_X1 U8526 ( .A1(n8145), .A2(n6634), .ZN(n6633) );
  NAND2_X1 U8527 ( .A1(n7986), .A2(n6633), .ZN(n6648) );
  INV_X1 U8528 ( .A(n6634), .ZN(n6646) );
  INV_X1 U8529 ( .A(n6635), .ZN(n6636) );
  NAND2_X1 U8530 ( .A1(n6637), .A2(n6636), .ZN(n8146) );
  INV_X1 U8531 ( .A(n6638), .ZN(n6641) );
  INV_X1 U8532 ( .A(n6639), .ZN(n6640) );
  NAND2_X1 U8533 ( .A1(n6641), .A2(n6640), .ZN(n6642) );
  NAND2_X1 U8534 ( .A1(n8157), .A2(n6642), .ZN(n8150) );
  INV_X1 U8535 ( .A(n8150), .ZN(n6643) );
  AND2_X1 U8536 ( .A1(n8146), .A2(n6643), .ZN(n8147) );
  AND2_X1 U8537 ( .A1(n8147), .A2(n6644), .ZN(n6645) );
  OR2_X1 U8538 ( .A1(n6646), .A2(n6645), .ZN(n6647) );
  NAND2_X1 U8539 ( .A1(n6648), .A2(n6647), .ZN(n8165) );
  XNOR2_X1 U8540 ( .A(n9574), .B(n6719), .ZN(n6651) );
  NAND2_X1 U8541 ( .A1(n9117), .A2(n6670), .ZN(n6649) );
  XNOR2_X1 U8542 ( .A(n6651), .B(n6649), .ZN(n8166) );
  INV_X1 U8543 ( .A(n6649), .ZN(n6650) );
  AND2_X1 U8544 ( .A1(n6651), .A2(n6650), .ZN(n6652) );
  XNOR2_X1 U8545 ( .A(n6570), .B(n6715), .ZN(n6653) );
  NAND2_X1 U8546 ( .A1(n9116), .A2(n6670), .ZN(n6654) );
  NAND2_X1 U8547 ( .A1(n6653), .A2(n6654), .ZN(n6658) );
  INV_X1 U8548 ( .A(n6653), .ZN(n6656) );
  INV_X1 U8549 ( .A(n6654), .ZN(n6655) );
  NAND2_X1 U8550 ( .A1(n6656), .A2(n6655), .ZN(n6657) );
  AND2_X1 U8551 ( .A1(n6658), .A2(n6657), .ZN(n8993) );
  NAND2_X1 U8552 ( .A1(n8994), .A2(n8993), .ZN(n8992) );
  NAND2_X1 U8553 ( .A1(n8992), .A2(n6658), .ZN(n8373) );
  XNOR2_X1 U8554 ( .A(n9565), .B(n6715), .ZN(n6659) );
  NAND2_X1 U8555 ( .A1(n9115), .A2(n6670), .ZN(n6660) );
  XNOR2_X1 U8556 ( .A(n6659), .B(n6660), .ZN(n8372) );
  INV_X1 U8557 ( .A(n8372), .ZN(n6663) );
  INV_X1 U8558 ( .A(n6659), .ZN(n6662) );
  INV_X1 U8559 ( .A(n6660), .ZN(n6661) );
  XNOR2_X1 U8560 ( .A(n6337), .B(n6715), .ZN(n6664) );
  NAND2_X1 U8561 ( .A1(n9400), .A2(n6670), .ZN(n6665) );
  NAND2_X1 U8562 ( .A1(n6664), .A2(n6665), .ZN(n6669) );
  INV_X1 U8563 ( .A(n6664), .ZN(n6667) );
  INV_X1 U8564 ( .A(n6665), .ZN(n6666) );
  NAND2_X1 U8565 ( .A1(n6667), .A2(n6666), .ZN(n6668) );
  AND2_X1 U8566 ( .A1(n6669), .A2(n6668), .ZN(n8609) );
  XNOR2_X1 U8567 ( .A(n9556), .B(n6715), .ZN(n9009) );
  NAND2_X1 U8568 ( .A1(n9381), .A2(n6670), .ZN(n9011) );
  AND2_X1 U8569 ( .A1(n9009), .A2(n9011), .ZN(n6674) );
  XNOR2_X1 U8570 ( .A(n6675), .B(n6671), .ZN(n9013) );
  NAND2_X1 U8571 ( .A1(n9382), .A2(n6670), .ZN(n6678) );
  XNOR2_X1 U8572 ( .A(n9545), .B(n6719), .ZN(n6677) );
  XOR2_X1 U8573 ( .A(n6678), .B(n6677), .Z(n9024) );
  XNOR2_X1 U8574 ( .A(n9539), .B(n6719), .ZN(n6680) );
  NAND2_X1 U8575 ( .A1(n9359), .A2(n6670), .ZN(n6679) );
  XNOR2_X1 U8576 ( .A(n6680), .B(n6679), .ZN(n9077) );
  INV_X1 U8577 ( .A(n6679), .ZN(n6681) );
  AND2_X1 U8578 ( .A1(n9346), .A2(n6670), .ZN(n6683) );
  XNOR2_X1 U8579 ( .A(n9535), .B(n6719), .ZN(n6682) );
  NOR2_X1 U8580 ( .A1(n6682), .A2(n6683), .ZN(n6684) );
  AOI21_X1 U8581 ( .B1(n6683), .B2(n6682), .A(n6684), .ZN(n8975) );
  INV_X1 U8582 ( .A(n6684), .ZN(n6685) );
  XNOR2_X1 U8583 ( .A(n9528), .B(n6719), .ZN(n6686) );
  NOR2_X1 U8584 ( .A1(n8987), .A2(n7759), .ZN(n6687) );
  XNOR2_X1 U8585 ( .A(n6686), .B(n6687), .ZN(n9054) );
  INV_X1 U8586 ( .A(n6686), .ZN(n6689) );
  INV_X1 U8587 ( .A(n6687), .ZN(n6688) );
  XNOR2_X1 U8588 ( .A(n9523), .B(n6719), .ZN(n6693) );
  NAND2_X1 U8589 ( .A1(n9314), .A2(n6670), .ZN(n6690) );
  XNOR2_X1 U8590 ( .A(n6693), .B(n6690), .ZN(n8983) );
  NAND2_X1 U8591 ( .A1(n8984), .A2(n8983), .ZN(n9064) );
  XNOR2_X1 U8592 ( .A(n9520), .B(n6719), .ZN(n9065) );
  NOR2_X1 U8593 ( .A1(n9264), .A2(n7759), .ZN(n9066) );
  NOR2_X1 U8594 ( .A1(n9065), .A2(n9066), .ZN(n6696) );
  INV_X1 U8595 ( .A(n6690), .ZN(n6692) );
  AND2_X1 U8596 ( .A1(n6693), .A2(n6692), .ZN(n9062) );
  OAI21_X1 U8597 ( .B1(n9062), .B2(n9066), .A(n9065), .ZN(n6691) );
  OAI21_X2 U8598 ( .B1(n9064), .B2(n6696), .A(n6695), .ZN(n6702) );
  XNOR2_X1 U8599 ( .A(n9515), .B(n6719), .ZN(n6700) );
  INV_X1 U8600 ( .A(n9035), .ZN(n6698) );
  INV_X1 U8601 ( .A(n9034), .ZN(n6697) );
  XNOR2_X2 U8602 ( .A(n6702), .B(n6701), .ZN(n9033) );
  AND2_X1 U8603 ( .A1(n9282), .A2(n6670), .ZN(n9032) );
  XNOR2_X1 U8604 ( .A(n9498), .B(n6715), .ZN(n6708) );
  NAND2_X1 U8605 ( .A1(n9203), .A2(n6670), .ZN(n6709) );
  NAND2_X1 U8606 ( .A1(n6708), .A2(n6709), .ZN(n9089) );
  NAND2_X1 U8607 ( .A1(n9084), .A2(n5047), .ZN(n6714) );
  NAND3_X1 U8608 ( .A1(n9089), .A2(n9001), .A3(n9087), .ZN(n6712) );
  INV_X1 U8609 ( .A(n6708), .ZN(n6711) );
  INV_X1 U8610 ( .A(n6709), .ZN(n6710) );
  NAND2_X1 U8611 ( .A1(n6711), .A2(n6710), .ZN(n9088) );
  XNOR2_X1 U8612 ( .A(n9493), .B(n6715), .ZN(n6717) );
  NAND2_X1 U8613 ( .A1(n9220), .A2(n6670), .ZN(n6716) );
  NOR2_X1 U8614 ( .A1(n6717), .A2(n6716), .ZN(n6718) );
  AOI21_X1 U8615 ( .B1(n6717), .B2(n6716), .A(n6718), .ZN(n8962) );
  NAND2_X1 U8616 ( .A1(n9204), .A2(n6670), .ZN(n6720) );
  XNOR2_X1 U8617 ( .A(n6720), .B(n6719), .ZN(n6726) );
  NAND2_X1 U8618 ( .A1(n6734), .A2(n6722), .ZN(n6723) );
  NOR3_X1 U8619 ( .A1(n6730), .A2(n9108), .A3(n6726), .ZN(n6724) );
  AOI21_X1 U8620 ( .B1(n6730), .B2(n6726), .A(n6724), .ZN(n6732) );
  NAND3_X1 U8621 ( .A1(n9488), .A2(n9023), .A3(n6726), .ZN(n6725) );
  OAI21_X1 U8622 ( .B1(n9488), .B2(n6726), .A(n6725), .ZN(n6727) );
  AND2_X1 U8623 ( .A1(n10507), .A2(n6728), .ZN(n6729) );
  OAI21_X1 U8624 ( .B1(n6730), .B2(n9023), .A(n9110), .ZN(n6731) );
  AOI21_X1 U8625 ( .B1(n6736), .B2(n6756), .A(n6735), .ZN(n7742) );
  NAND3_X1 U8626 ( .A1(n7742), .A2(n6738), .A3(n6737), .ZN(n6739) );
  AOI22_X1 U8627 ( .A1(n9113), .A2(n9092), .B1(n6740), .B2(n9102), .ZN(n6742)
         );
  AOI22_X1 U8628 ( .A1(n9220), .A2(n9103), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n6741) );
  NAND2_X1 U8629 ( .A1(n6743), .A2(n5028), .ZN(P2_U3222) );
  NAND2_X1 U8630 ( .A1(n9623), .A2(n7176), .ZN(n6745) );
  NAND2_X1 U8631 ( .A1(n7177), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6744) );
  NAND2_X1 U8632 ( .A1(n8953), .A2(n7176), .ZN(n6747) );
  NAND2_X1 U8633 ( .A1(n7177), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6746) );
  NAND2_X1 U8634 ( .A1(n8915), .A2(n8900), .ZN(n9198) );
  NAND2_X1 U8635 ( .A1(n6749), .A2(P2_B_REG_SCAN_IN), .ZN(n6750) );
  AND2_X1 U8636 ( .A1(n9444), .A2(n6750), .ZN(n8911) );
  NAND2_X1 U8637 ( .A1(n6257), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6754) );
  NAND2_X1 U8638 ( .A1(n7169), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6753) );
  INV_X1 U8639 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n6751) );
  OR2_X1 U8640 ( .A1(n7172), .A2(n6751), .ZN(n6752) );
  AND3_X1 U8641 ( .A1(n6754), .A2(n6753), .A3(n6752), .ZN(n7180) );
  INV_X1 U8642 ( .A(n7180), .ZN(n7431) );
  NAND2_X1 U8643 ( .A1(n8911), .A2(n7431), .ZN(n9480) );
  NAND2_X1 U8644 ( .A1(n7182), .A2(n9588), .ZN(n6755) );
  NAND2_X1 U8645 ( .A1(n6757), .A2(n6756), .ZN(n6758) );
  NAND2_X1 U8646 ( .A1(n9482), .A2(n10516), .ZN(n6762) );
  OR2_X1 U8647 ( .A1(n10516), .A2(n6760), .ZN(n6761) );
  NAND2_X1 U8648 ( .A1(n6762), .A2(n6761), .ZN(n7011) );
  NOR4_X1 U8649 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n7073) );
  INV_X1 U8650 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10357) );
  INV_X1 U8651 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10356) );
  INV_X1 U8652 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10358) );
  INV_X1 U8653 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10360) );
  NAND4_X1 U8654 ( .A1(n10357), .A2(n10356), .A3(n10358), .A4(n10360), .ZN(
        n7069) );
  INV_X1 U8655 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n6849) );
  INV_X1 U8656 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6989) );
  NOR4_X1 U8657 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_18__SCAN_IN), 
        .A3(n6849), .A4(n6989), .ZN(n6767) );
  NOR4_X1 U8658 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(P1_REG3_REG_9__SCAN_IN), 
        .A3(P1_REG2_REG_22__SCAN_IN), .A4(n8174), .ZN(n6764) );
  NOR4_X1 U8659 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(P1_DATAO_REG_15__SCAN_IN), 
        .A3(SI_13_), .A4(n6898), .ZN(n6763) );
  NAND4_X1 U8660 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_DATAO_REG_0__SCAN_IN), 
        .A3(n6764), .A4(n6763), .ZN(n6765) );
  NOR3_X1 U8661 ( .A1(n6765), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n6766) );
  NAND2_X1 U8662 ( .A1(n6767), .A2(n6766), .ZN(n6768) );
  NOR4_X1 U8663 ( .A1(n7069), .A2(n6769), .A3(n7562), .A4(n6768), .ZN(n6770)
         );
  NAND4_X1 U8664 ( .A1(n7073), .A2(P2_DATAO_REG_9__SCAN_IN), .A3(
        P1_REG0_REG_16__SCAN_IN), .A4(n6770), .ZN(n6797) );
  NAND4_X1 U8665 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_REG0_REG_23__SCAN_IN), 
        .A3(n6771), .A4(P2_REG0_REG_10__SCAN_IN), .ZN(n6796) );
  NOR4_X1 U8666 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(P1_REG2_REG_18__SCAN_IN), 
        .A3(P2_REG2_REG_16__SCAN_IN), .A4(P2_REG1_REG_15__SCAN_IN), .ZN(n6772)
         );
  NAND3_X1 U8667 ( .A1(SI_10_), .A2(P1_REG1_REG_27__SCAN_IN), .A3(n6772), .ZN(
        n6795) );
  NAND4_X1 U8668 ( .A1(n8575), .A2(n4539), .A3(SI_7_), .A4(
        P2_REG3_REG_14__SCAN_IN), .ZN(n6774) );
  NAND2_X1 U8669 ( .A1(P2_REG2_REG_24__SCAN_IN), .A2(P1_DATAO_REG_5__SCAN_IN), 
        .ZN(n6773) );
  NOR4_X1 U8670 ( .A1(n6774), .A2(n8718), .A3(n6773), .A4(
        P2_REG0_REG_11__SCAN_IN), .ZN(n6788) );
  NAND4_X1 U8671 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(P1_REG1_REG_12__SCAN_IN), 
        .A3(P2_REG0_REG_14__SCAN_IN), .A4(n6923), .ZN(n6776) );
  NAND4_X1 U8672 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), 
        .A3(P1_REG1_REG_13__SCAN_IN), .A4(n10237), .ZN(n6775) );
  NOR2_X1 U8673 ( .A1(n6776), .A2(n6775), .ZN(n6783) );
  INV_X1 U8674 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9462) );
  NAND4_X1 U8675 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(P2_REG0_REG_15__SCAN_IN), 
        .A3(n6831), .A4(n9462), .ZN(n6778) );
  NAND4_X1 U8676 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(P2_DATAO_REG_28__SCAN_IN), 
        .A3(P1_REG1_REG_0__SCAN_IN), .A4(n6916), .ZN(n6777) );
  NOR2_X1 U8677 ( .A1(n6778), .A2(n6777), .ZN(n6782) );
  NAND4_X1 U8678 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), 
        .A3(n6483), .A4(n6828), .ZN(n6779) );
  INV_X1 U8679 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7974) );
  NOR2_X1 U8680 ( .A1(n6779), .A2(n7974), .ZN(n6781) );
  INV_X1 U8681 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10177) );
  NOR4_X1 U8682 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_REG0_REG_21__SCAN_IN), 
        .A3(n10177), .A4(n4812), .ZN(n6780) );
  NAND4_X1 U8683 ( .A1(n6783), .A2(n6782), .A3(n6781), .A4(n6780), .ZN(n6784)
         );
  NOR2_X1 U8684 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(n6784), .ZN(n6787) );
  NOR4_X1 U8685 ( .A1(P2_U3152), .A2(n6785), .A3(P2_IR_REG_11__SCAN_IN), .A4(
        P2_IR_REG_25__SCAN_IN), .ZN(n6786) );
  NAND4_X1 U8686 ( .A1(n6788), .A2(P1_D_REG_6__SCAN_IN), .A3(n6787), .A4(n6786), .ZN(n6793) );
  NAND4_X1 U8687 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_REG1_REG_18__SCAN_IN), 
        .A3(P2_REG3_REG_2__SCAN_IN), .A4(n6852), .ZN(n6792) );
  NAND4_X1 U8688 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), 
        .A3(P1_D_REG_2__SCAN_IN), .A4(P2_REG2_REG_26__SCAN_IN), .ZN(n6791) );
  NAND4_X1 U8689 ( .A1(n10289), .A2(n10440), .A3(n6789), .A4(
        P2_D_REG_27__SCAN_IN), .ZN(n6790) );
  OR4_X1 U8690 ( .A1(n6793), .A2(n6792), .A3(n6791), .A4(n6790), .ZN(n6794) );
  NOR4_X1 U8691 ( .A1(n6797), .A2(n6796), .A3(n6795), .A4(n6794), .ZN(n6809)
         );
  INV_X1 U8692 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8954) );
  NOR4_X1 U8693 ( .A1(P2_REG2_REG_9__SCAN_IN), .A2(P2_REG2_REG_27__SCAN_IN), 
        .A3(n6811), .A4(n8954), .ZN(n6798) );
  NAND3_X1 U8694 ( .A1(P1_REG0_REG_8__SCAN_IN), .A2(P2_REG2_REG_29__SCAN_IN), 
        .A3(n6798), .ZN(n6807) );
  NAND4_X1 U8695 ( .A1(P1_REG0_REG_19__SCAN_IN), .A2(P1_REG0_REG_12__SCAN_IN), 
        .A3(P1_REG0_REG_7__SCAN_IN), .A4(P2_REG1_REG_5__SCAN_IN), .ZN(n6799)
         );
  NOR3_X1 U8696 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(n6799), .ZN(n6805) );
  NAND4_X1 U8697 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(P2_DATAO_REG_30__SCAN_IN), 
        .A3(n7483), .A4(n7895), .ZN(n6802) );
  NAND4_X1 U8698 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .A3(
        P2_REG2_REG_25__SCAN_IN), .A4(n6894), .ZN(n6801) );
  INV_X1 U8699 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n6912) );
  NAND4_X1 U8700 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P2_REG1_REG_14__SCAN_IN), 
        .A3(n6912), .A4(n9459), .ZN(n6800) );
  NOR4_X1 U8701 ( .A1(SI_5_), .A2(n6802), .A3(n6801), .A4(n6800), .ZN(n6803)
         );
  AND4_X1 U8702 ( .A1(n6803), .A2(P2_REG2_REG_18__SCAN_IN), .A3(
        P1_REG0_REG_3__SCAN_IN), .A4(n9069), .ZN(n6804) );
  NAND4_X1 U8703 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(P2_REG0_REG_5__SCAN_IN), 
        .A3(n6805), .A4(n6804), .ZN(n6806) );
  NOR4_X1 U8704 ( .A1(P1_REG1_REG_22__SCAN_IN), .A2(n7682), .A3(n6807), .A4(
        n6806), .ZN(n6808) );
  AOI21_X1 U8705 ( .B1(n6809), .B2(n6808), .A(n8478), .ZN(n7009) );
  INV_X1 U8706 ( .A(keyinput97), .ZN(n7008) );
  AOI22_X1 U8707 ( .A1(n7658), .A2(keyinput25), .B1(keyinput63), .B2(n6811), 
        .ZN(n6810) );
  OAI221_X1 U8708 ( .B1(n7658), .B2(keyinput25), .C1(n6811), .C2(keyinput63), 
        .A(n6810), .ZN(n6819) );
  AOI22_X1 U8709 ( .A1(n6479), .A2(keyinput59), .B1(keyinput20), .B2(n8954), 
        .ZN(n6812) );
  OAI221_X1 U8710 ( .B1(n6479), .B2(keyinput59), .C1(n8954), .C2(keyinput20), 
        .A(n6812), .ZN(n6818) );
  INV_X1 U8711 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10359) );
  AOI22_X1 U8712 ( .A1(n8550), .A2(keyinput41), .B1(n10359), .B2(keyinput119), 
        .ZN(n6813) );
  OAI221_X1 U8713 ( .B1(n8550), .B2(keyinput41), .C1(n10359), .C2(keyinput119), 
        .A(n6813), .ZN(n6817) );
  AOI22_X1 U8714 ( .A1(n6815), .A2(keyinput28), .B1(n7682), .B2(keyinput11), 
        .ZN(n6814) );
  OAI221_X1 U8715 ( .B1(n6815), .B2(keyinput28), .C1(n7682), .C2(keyinput11), 
        .A(n6814), .ZN(n6816) );
  NOR4_X1 U8716 ( .A1(n6819), .A2(n6818), .A3(n6817), .A4(n6816), .ZN(n7007)
         );
  AOI22_X1 U8717 ( .A1(n7974), .A2(keyinput37), .B1(keyinput53), .B2(n6821), 
        .ZN(n6820) );
  OAI221_X1 U8718 ( .B1(n7974), .B2(keyinput37), .C1(n6821), .C2(keyinput53), 
        .A(n6820), .ZN(n6826) );
  AOI22_X1 U8719 ( .A1(n10476), .A2(keyinput116), .B1(keyinput56), .B2(n6823), 
        .ZN(n6822) );
  OAI221_X1 U8720 ( .B1(n10476), .B2(keyinput116), .C1(n6823), .C2(keyinput56), 
        .A(n6822), .ZN(n6825) );
  INV_X1 U8721 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n10479) );
  XNOR2_X1 U8722 ( .A(n10479), .B(keyinput10), .ZN(n6824) );
  OR3_X1 U8723 ( .A1(n6826), .A2(n6825), .A3(n6824), .ZN(n6835) );
  AOI22_X1 U8724 ( .A1(n6829), .A2(keyinput121), .B1(keyinput45), .B2(n6828), 
        .ZN(n6827) );
  OAI221_X1 U8725 ( .B1(n6829), .B2(keyinput121), .C1(n6828), .C2(keyinput45), 
        .A(n6827), .ZN(n6834) );
  AOI22_X1 U8726 ( .A1(n9462), .A2(keyinput46), .B1(n6831), .B2(keyinput55), 
        .ZN(n6830) );
  OAI221_X1 U8727 ( .B1(n9462), .B2(keyinput46), .C1(n6831), .C2(keyinput55), 
        .A(n6830), .ZN(n6833) );
  INV_X1 U8728 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10366) );
  XNOR2_X1 U8729 ( .A(n10366), .B(keyinput34), .ZN(n6832) );
  OR4_X1 U8730 ( .A1(n6835), .A2(n6834), .A3(n6833), .A4(n6832), .ZN(n6862) );
  AOI22_X1 U8731 ( .A1(n10360), .A2(keyinput105), .B1(keyinput57), .B2(n6837), 
        .ZN(n6836) );
  OAI221_X1 U8732 ( .B1(n10360), .B2(keyinput105), .C1(n6837), .C2(keyinput57), 
        .A(n6836), .ZN(n6838) );
  INV_X1 U8733 ( .A(n6838), .ZN(n6858) );
  XNOR2_X1 U8734 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput15), .ZN(n6842) );
  XNOR2_X1 U8735 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput69), .ZN(n6841) );
  XNOR2_X1 U8736 ( .A(P2_IR_REG_28__SCAN_IN), .B(keyinput1), .ZN(n6840) );
  XNOR2_X1 U8737 ( .A(keyinput125), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n6839) );
  NAND4_X1 U8738 ( .A1(n6842), .A2(n6841), .A3(n6840), .A4(n6839), .ZN(n6848)
         );
  XNOR2_X1 U8739 ( .A(keyinput113), .B(P2_IR_REG_24__SCAN_IN), .ZN(n6846) );
  XNOR2_X1 U8740 ( .A(keyinput87), .B(P2_REG2_REG_3__SCAN_IN), .ZN(n6845) );
  XNOR2_X1 U8741 ( .A(keyinput91), .B(P1_D_REG_6__SCAN_IN), .ZN(n6844) );
  XNOR2_X1 U8742 ( .A(keyinput85), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n6843) );
  NAND4_X1 U8743 ( .A1(n6846), .A2(n6845), .A3(n6844), .A4(n6843), .ZN(n6847)
         );
  NOR2_X1 U8744 ( .A1(n6848), .A2(n6847), .ZN(n6857) );
  XNOR2_X1 U8745 ( .A(keyinput77), .B(n6849), .ZN(n6851) );
  INV_X1 U8746 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10385) );
  XNOR2_X1 U8747 ( .A(keyinput51), .B(n10385), .ZN(n6850) );
  NOR2_X1 U8748 ( .A1(n6851), .A2(n6850), .ZN(n6856) );
  XNOR2_X1 U8749 ( .A(keyinput64), .B(n6852), .ZN(n6854) );
  XNOR2_X1 U8750 ( .A(keyinput6), .B(n6483), .ZN(n6853) );
  NOR2_X1 U8751 ( .A1(n6854), .A2(n6853), .ZN(n6855) );
  NAND4_X1 U8752 ( .A1(n6858), .A2(n6857), .A3(n6856), .A4(n6855), .ZN(n6861)
         );
  XNOR2_X1 U8753 ( .A(n10357), .B(keyinput65), .ZN(n6860) );
  XNOR2_X1 U8754 ( .A(n10480), .B(keyinput29), .ZN(n6859) );
  NOR4_X1 U8755 ( .A1(n6862), .A2(n6861), .A3(n6860), .A4(n6859), .ZN(n6870)
         );
  INV_X1 U8756 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n6864) );
  OAI22_X1 U8757 ( .A1(n7895), .A2(keyinput79), .B1(n6864), .B2(keyinput8), 
        .ZN(n6863) );
  AOI221_X1 U8758 ( .B1(n7895), .B2(keyinput79), .C1(keyinput8), .C2(n6864), 
        .A(n6863), .ZN(n6869) );
  INV_X1 U8759 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n10474) );
  OAI22_X1 U8760 ( .A1(P2_U3152), .A2(keyinput61), .B1(n10474), .B2(
        keyinput100), .ZN(n6865) );
  AOI221_X1 U8761 ( .B1(P2_U3152), .B2(keyinput61), .C1(keyinput100), .C2(
        n10474), .A(n6865), .ZN(n6868) );
  OAI22_X1 U8762 ( .A1(n7483), .A2(keyinput88), .B1(n9186), .B2(keyinput52), 
        .ZN(n6866) );
  AOI221_X1 U8763 ( .B1(n7483), .B2(keyinput88), .C1(keyinput52), .C2(n9186), 
        .A(n6866), .ZN(n6867) );
  NAND4_X1 U8764 ( .A1(n6870), .A2(n6869), .A3(n6868), .A4(n6867), .ZN(n7005)
         );
  AOI22_X1 U8765 ( .A1(n6873), .A2(keyinput19), .B1(n6872), .B2(keyinput38), 
        .ZN(n6871) );
  OAI221_X1 U8766 ( .B1(n6873), .B2(keyinput19), .C1(n6872), .C2(keyinput38), 
        .A(n6871), .ZN(n6881) );
  AOI22_X1 U8767 ( .A1(n10237), .A2(keyinput112), .B1(n10358), .B2(keyinput54), 
        .ZN(n6874) );
  OAI221_X1 U8768 ( .B1(n10237), .B2(keyinput112), .C1(n10358), .C2(keyinput54), .A(n6874), .ZN(n6880) );
  AOI22_X1 U8769 ( .A1(n8174), .A2(keyinput84), .B1(n10475), .B2(keyinput27), 
        .ZN(n6875) );
  OAI221_X1 U8770 ( .B1(n8174), .B2(keyinput84), .C1(n10475), .C2(keyinput27), 
        .A(n6875), .ZN(n6879) );
  INV_X1 U8771 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n10477) );
  AOI22_X1 U8772 ( .A1(n6877), .A2(keyinput21), .B1(n10477), .B2(keyinput108), 
        .ZN(n6876) );
  OAI221_X1 U8773 ( .B1(n6877), .B2(keyinput21), .C1(n10477), .C2(keyinput108), 
        .A(n6876), .ZN(n6878) );
  NOR4_X1 U8774 ( .A1(n6881), .A2(n6880), .A3(n6879), .A4(n6878), .ZN(n6932)
         );
  INV_X1 U8775 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10361) );
  AOI22_X1 U8776 ( .A1(n7866), .A2(keyinput17), .B1(n10361), .B2(keyinput86), 
        .ZN(n6882) );
  OAI221_X1 U8777 ( .B1(n7866), .B2(keyinput17), .C1(n10361), .C2(keyinput86), 
        .A(n6882), .ZN(n6890) );
  INV_X1 U8778 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10426) );
  AOI22_X1 U8779 ( .A1(n8919), .A2(keyinput44), .B1(n10426), .B2(keyinput111), 
        .ZN(n6883) );
  OAI221_X1 U8780 ( .B1(n8919), .B2(keyinput44), .C1(n10426), .C2(keyinput111), 
        .A(n6883), .ZN(n6889) );
  INV_X1 U8781 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10362) );
  AOI22_X1 U8782 ( .A1(n6885), .A2(keyinput3), .B1(n10362), .B2(keyinput4), 
        .ZN(n6884) );
  OAI221_X1 U8783 ( .B1(n6885), .B2(keyinput3), .C1(n10362), .C2(keyinput4), 
        .A(n6884), .ZN(n6888) );
  AOI22_X1 U8784 ( .A1(n5124), .A2(keyinput0), .B1(n8718), .B2(keyinput22), 
        .ZN(n6886) );
  OAI221_X1 U8785 ( .B1(n5124), .B2(keyinput0), .C1(n8718), .C2(keyinput22), 
        .A(n6886), .ZN(n6887) );
  NOR4_X1 U8786 ( .A1(n6890), .A2(n6889), .A3(n6888), .A4(n6887), .ZN(n6931)
         );
  AOI22_X1 U8787 ( .A1(n6892), .A2(keyinput99), .B1(n4539), .B2(keyinput30), 
        .ZN(n6891) );
  OAI221_X1 U8788 ( .B1(n6892), .B2(keyinput99), .C1(n4539), .C2(keyinput30), 
        .A(n6891), .ZN(n6902) );
  AOI22_X1 U8789 ( .A1(n6895), .A2(keyinput2), .B1(n6894), .B2(keyinput13), 
        .ZN(n6893) );
  OAI221_X1 U8790 ( .B1(n6895), .B2(keyinput2), .C1(n6894), .C2(keyinput13), 
        .A(n6893), .ZN(n6901) );
  AOI22_X1 U8791 ( .A1(n7526), .A2(keyinput36), .B1(n8496), .B2(keyinput60), 
        .ZN(n6896) );
  OAI221_X1 U8792 ( .B1(n7526), .B2(keyinput36), .C1(n8496), .C2(keyinput60), 
        .A(n6896), .ZN(n6900) );
  AOI22_X1 U8793 ( .A1(n6898), .A2(keyinput58), .B1(n7680), .B2(keyinput122), 
        .ZN(n6897) );
  OAI221_X1 U8794 ( .B1(n6898), .B2(keyinput58), .C1(n7680), .C2(keyinput122), 
        .A(n6897), .ZN(n6899) );
  OR4_X1 U8795 ( .A1(n6902), .A2(n6901), .A3(n6900), .A4(n6899), .ZN(n6908) );
  INV_X1 U8796 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10365) );
  AOI22_X1 U8797 ( .A1(n10365), .A2(keyinput76), .B1(keyinput106), .B2(n6464), 
        .ZN(n6903) );
  OAI221_X1 U8798 ( .B1(n10365), .B2(keyinput76), .C1(n6464), .C2(keyinput106), 
        .A(n6903), .ZN(n6907) );
  INV_X1 U8799 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n6905) );
  AOI22_X1 U8800 ( .A1(n8334), .A2(keyinput98), .B1(keyinput127), .B2(n6905), 
        .ZN(n6904) );
  OAI221_X1 U8801 ( .B1(n8334), .B2(keyinput98), .C1(n6905), .C2(keyinput127), 
        .A(n6904), .ZN(n6906) );
  NOR3_X1 U8802 ( .A1(n6908), .A2(n6907), .A3(n6906), .ZN(n6930) );
  AOI22_X1 U8803 ( .A1(n4812), .A2(keyinput18), .B1(keyinput124), .B2(n10177), 
        .ZN(n6909) );
  OAI221_X1 U8804 ( .B1(n4812), .B2(keyinput18), .C1(n10177), .C2(keyinput124), 
        .A(n6909), .ZN(n6921) );
  INV_X1 U8805 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6911) );
  AOI22_X1 U8806 ( .A1(n6912), .A2(keyinput42), .B1(keyinput70), .B2(n6911), 
        .ZN(n6910) );
  OAI221_X1 U8807 ( .B1(n6912), .B2(keyinput42), .C1(n6911), .C2(keyinput70), 
        .A(n6910), .ZN(n6920) );
  AOI22_X1 U8808 ( .A1(n6914), .A2(keyinput9), .B1(keyinput114), .B2(n8575), 
        .ZN(n6913) );
  OAI221_X1 U8809 ( .B1(n6914), .B2(keyinput9), .C1(n8575), .C2(keyinput114), 
        .A(n6913), .ZN(n6919) );
  AOI22_X1 U8810 ( .A1(n6917), .A2(keyinput67), .B1(keyinput103), .B2(n6916), 
        .ZN(n6915) );
  OAI221_X1 U8811 ( .B1(n6917), .B2(keyinput67), .C1(n6916), .C2(keyinput103), 
        .A(n6915), .ZN(n6918) );
  OR4_X1 U8812 ( .A1(n6921), .A2(n6920), .A3(n6919), .A4(n6918), .ZN(n6928) );
  AOI22_X1 U8813 ( .A1(n6924), .A2(keyinput16), .B1(n6923), .B2(keyinput81), 
        .ZN(n6922) );
  OAI221_X1 U8814 ( .B1(n6924), .B2(keyinput16), .C1(n6923), .C2(keyinput81), 
        .A(n6922), .ZN(n6927) );
  INV_X1 U8815 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10436) );
  AOI22_X1 U8816 ( .A1(n10356), .A2(keyinput68), .B1(keyinput95), .B2(n10436), 
        .ZN(n6925) );
  OAI221_X1 U8817 ( .B1(n10356), .B2(keyinput68), .C1(n10436), .C2(keyinput95), 
        .A(n6925), .ZN(n6926) );
  NOR3_X1 U8818 ( .A1(n6928), .A2(n6927), .A3(n6926), .ZN(n6929) );
  NAND4_X1 U8819 ( .A1(n6932), .A2(n6931), .A3(n6930), .A4(n6929), .ZN(n7004)
         );
  INV_X1 U8820 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10568) );
  AOI22_X1 U8821 ( .A1(n6219), .A2(keyinput7), .B1(keyinput50), .B2(n10568), 
        .ZN(n6933) );
  OAI221_X1 U8822 ( .B1(n6219), .B2(keyinput7), .C1(n10568), .C2(keyinput50), 
        .A(n6933), .ZN(n6999) );
  AOI22_X1 U8823 ( .A1(n6935), .A2(keyinput126), .B1(keyinput5), .B2(n10245), 
        .ZN(n6934) );
  OAI221_X1 U8824 ( .B1(n6935), .B2(keyinput126), .C1(n10245), .C2(keyinput5), 
        .A(n6934), .ZN(n6943) );
  INV_X1 U8825 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6937) );
  AOI22_X1 U8826 ( .A1(n6937), .A2(keyinput123), .B1(n8613), .B2(keyinput40), 
        .ZN(n6936) );
  OAI221_X1 U8827 ( .B1(n6937), .B2(keyinput123), .C1(n8613), .C2(keyinput40), 
        .A(n6936), .ZN(n6942) );
  INV_X1 U8828 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6939) );
  AOI22_X1 U8829 ( .A1(n6940), .A2(keyinput107), .B1(keyinput66), .B2(n6939), 
        .ZN(n6938) );
  OAI221_X1 U8830 ( .B1(n6940), .B2(keyinput107), .C1(n6939), .C2(keyinput66), 
        .A(n6938), .ZN(n6941) );
  OR3_X1 U8831 ( .A1(n6943), .A2(n6942), .A3(n6941), .ZN(n6998) );
  XNOR2_X1 U8832 ( .A(SI_5_), .B(keyinput117), .ZN(n6947) );
  XNOR2_X1 U8833 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput82), .ZN(n6946) );
  XNOR2_X1 U8834 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput96), .ZN(n6945) );
  XNOR2_X1 U8835 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(keyinput110), .ZN(n6944)
         );
  NAND4_X1 U8836 ( .A1(n6947), .A2(n6946), .A3(n6945), .A4(n6944), .ZN(n6953)
         );
  XNOR2_X1 U8837 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput14), .ZN(n6951) );
  XNOR2_X1 U8838 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput89), .ZN(n6950) );
  XNOR2_X1 U8839 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput90), .ZN(n6949) );
  XNOR2_X1 U8840 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput93), .ZN(n6948) );
  NAND4_X1 U8841 ( .A1(n6951), .A2(n6950), .A3(n6949), .A4(n6948), .ZN(n6952)
         );
  NOR2_X1 U8842 ( .A1(n6953), .A2(n6952), .ZN(n6987) );
  XNOR2_X1 U8843 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput71), .ZN(n6957) );
  XNOR2_X1 U8844 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput48), .ZN(n6956) );
  XNOR2_X1 U8845 ( .A(P1_REG0_REG_12__SCAN_IN), .B(keyinput32), .ZN(n6955) );
  XNOR2_X1 U8846 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput35), .ZN(n6954) );
  NAND4_X1 U8847 ( .A1(n6957), .A2(n6956), .A3(n6955), .A4(n6954), .ZN(n6963)
         );
  XNOR2_X1 U8848 ( .A(P1_REG0_REG_16__SCAN_IN), .B(keyinput94), .ZN(n6961) );
  XNOR2_X1 U8849 ( .A(P1_REG1_REG_12__SCAN_IN), .B(keyinput23), .ZN(n6960) );
  XNOR2_X1 U8850 ( .A(P1_REG0_REG_19__SCAN_IN), .B(keyinput39), .ZN(n6959) );
  XNOR2_X1 U8851 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput72), .ZN(n6958) );
  NAND4_X1 U8852 ( .A1(n6961), .A2(n6960), .A3(n6959), .A4(n6958), .ZN(n6962)
         );
  NOR2_X1 U8853 ( .A1(n6963), .A2(n6962), .ZN(n6986) );
  XNOR2_X1 U8854 ( .A(P1_REG3_REG_8__SCAN_IN), .B(keyinput62), .ZN(n6967) );
  XNOR2_X1 U8855 ( .A(P1_REG3_REG_4__SCAN_IN), .B(keyinput47), .ZN(n6966) );
  XNOR2_X1 U8856 ( .A(P2_IR_REG_0__SCAN_IN), .B(keyinput104), .ZN(n6965) );
  XNOR2_X1 U8857 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput74), .ZN(n6964) );
  NAND4_X1 U8858 ( .A1(n6967), .A2(n6966), .A3(n6965), .A4(n6964), .ZN(n6973)
         );
  XNOR2_X1 U8859 ( .A(P2_IR_REG_12__SCAN_IN), .B(keyinput12), .ZN(n6971) );
  XNOR2_X1 U8860 ( .A(P2_REG0_REG_10__SCAN_IN), .B(keyinput24), .ZN(n6970) );
  XNOR2_X1 U8861 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput78), .ZN(n6969) );
  XNOR2_X1 U8862 ( .A(P2_REG0_REG_21__SCAN_IN), .B(keyinput115), .ZN(n6968) );
  NAND4_X1 U8863 ( .A1(n6971), .A2(n6970), .A3(n6969), .A4(n6968), .ZN(n6972)
         );
  NOR2_X1 U8864 ( .A1(n6973), .A2(n6972), .ZN(n6985) );
  XNOR2_X1 U8865 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(keyinput33), .ZN(n6977) );
  XNOR2_X1 U8866 ( .A(P2_REG2_REG_0__SCAN_IN), .B(keyinput73), .ZN(n6976) );
  XNOR2_X1 U8867 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput80), .ZN(n6975) );
  XNOR2_X1 U8868 ( .A(SI_7_), .B(keyinput109), .ZN(n6974) );
  NAND4_X1 U8869 ( .A1(n6977), .A2(n6976), .A3(n6975), .A4(n6974), .ZN(n6983)
         );
  XNOR2_X1 U8870 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput120), .ZN(n6981) );
  XNOR2_X1 U8871 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(keyinput101), .ZN(n6980) );
  XNOR2_X1 U8872 ( .A(P1_REG3_REG_3__SCAN_IN), .B(keyinput75), .ZN(n6979) );
  XNOR2_X1 U8873 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput83), .ZN(n6978) );
  NAND4_X1 U8874 ( .A1(n6981), .A2(n6980), .A3(n6979), .A4(n6978), .ZN(n6982)
         );
  NOR2_X1 U8875 ( .A1(n6983), .A2(n6982), .ZN(n6984) );
  NAND4_X1 U8876 ( .A1(n6987), .A2(n6986), .A3(n6985), .A4(n6984), .ZN(n6997)
         );
  AOI22_X1 U8877 ( .A1(n6989), .A2(keyinput102), .B1(n7987), .B2(keyinput43), 
        .ZN(n6988) );
  OAI221_X1 U8878 ( .B1(n6989), .B2(keyinput102), .C1(n7987), .C2(keyinput43), 
        .A(n6988), .ZN(n6995) );
  XNOR2_X1 U8879 ( .A(n6990), .B(keyinput118), .ZN(n6994) );
  XNOR2_X1 U8880 ( .A(n9069), .B(keyinput26), .ZN(n6993) );
  XNOR2_X1 U8881 ( .A(SI_10_), .B(keyinput49), .ZN(n6991) );
  OAI21_X1 U8882 ( .B1(keyinput97), .B2(n8478), .A(n6991), .ZN(n6992) );
  OR4_X1 U8883 ( .A1(n6995), .A2(n6994), .A3(n6993), .A4(n6992), .ZN(n6996) );
  NOR4_X1 U8884 ( .A1(n6999), .A2(n6998), .A3(n6997), .A4(n6996), .ZN(n7002)
         );
  INV_X1 U8885 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10232) );
  OAI22_X1 U8886 ( .A1(n10478), .A2(keyinput92), .B1(n10232), .B2(keyinput31), 
        .ZN(n7000) );
  AOI221_X1 U8887 ( .B1(n10478), .B2(keyinput92), .C1(keyinput31), .C2(n10232), 
        .A(n7000), .ZN(n7001) );
  NAND2_X1 U8888 ( .A1(n7002), .A2(n7001), .ZN(n7003) );
  NOR3_X1 U8889 ( .A1(n7005), .A2(n7004), .A3(n7003), .ZN(n7006) );
  OAI211_X1 U8890 ( .C1(n7009), .C2(n7008), .A(n7007), .B(n7006), .ZN(n7010)
         );
  XNOR2_X1 U8891 ( .A(n7011), .B(n7010), .ZN(P2_U3518) );
  INV_X1 U8892 ( .A(n8319), .ZN(n8315) );
  INV_X1 U8893 ( .A(n8317), .ZN(n7013) );
  NOR2_X1 U8894 ( .A1(n8315), .A2(n7013), .ZN(n7014) );
  NAND2_X1 U8895 ( .A1(n8318), .A2(n7014), .ZN(n7016) );
  NAND2_X1 U8896 ( .A1(n7016), .A2(n7015), .ZN(n8383) );
  NAND2_X1 U8897 ( .A1(n8383), .A2(n8384), .ZN(n7018) );
  NAND2_X1 U8898 ( .A1(n8509), .A2(n8505), .ZN(n7020) );
  OAI21_X2 U8899 ( .B1(n8741), .B2(n8742), .A(n7024), .ZN(n10038) );
  NAND2_X1 U8900 ( .A1(n10038), .A2(n7025), .ZN(n7027) );
  INV_X1 U8901 ( .A(n7028), .ZN(n7030) );
  OR2_X1 U8902 ( .A1(n9977), .A2(n7033), .ZN(n9963) );
  OR2_X1 U8903 ( .A1(n9963), .A2(n7034), .ZN(n9943) );
  NOR2_X1 U8904 ( .A1(n5045), .A2(n4697), .ZN(n7037) );
  INV_X1 U8905 ( .A(n9927), .ZN(n7038) );
  INV_X1 U8906 ( .A(n9881), .ZN(n7042) );
  NOR2_X1 U8907 ( .A1(n9886), .A2(n7042), .ZN(n7043) );
  AOI21_X1 U8908 ( .B1(n7045), .B2(n9847), .A(n7044), .ZN(n7046) );
  XNOR2_X1 U8909 ( .A(n7050), .B(n10101), .ZN(n7059) );
  NAND2_X1 U8910 ( .A1(n7051), .A2(n9990), .ZN(n7053) );
  INV_X1 U8911 ( .A(n7993), .ZN(n7155) );
  NAND2_X1 U8912 ( .A1(n4495), .A2(n7155), .ZN(n7052) );
  NAND2_X1 U8913 ( .A1(n10288), .A2(P1_B_REG_SCAN_IN), .ZN(n7054) );
  NAND2_X1 U8914 ( .A1(n10068), .A2(n7054), .ZN(n9836) );
  NAND2_X1 U8915 ( .A1(n9790), .A2(n10011), .ZN(n7056) );
  OAI21_X1 U8916 ( .B1(n7057), .B2(n9836), .A(n7056), .ZN(n7058) );
  NAND2_X1 U8917 ( .A1(n4509), .A2(n4757), .ZN(n7063) );
  NAND2_X1 U8918 ( .A1(n7061), .A2(n7063), .ZN(n8479) );
  OAI21_X1 U8919 ( .B1(n8479), .B2(P1_B_REG_SCAN_IN), .A(n7082), .ZN(n7062) );
  INV_X1 U8920 ( .A(n7062), .ZN(n7068) );
  NAND2_X1 U8921 ( .A1(n7063), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7064) );
  MUX2_X1 U8922 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7064), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n7066) );
  NAND2_X1 U8923 ( .A1(n7066), .A2(n7065), .ZN(n8574) );
  NAND3_X1 U8924 ( .A1(n8574), .A2(P1_B_REG_SCAN_IN), .A3(n8479), .ZN(n7067)
         );
  NOR2_X1 U8925 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .ZN(
        n7072) );
  NOR4_X1 U8926 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n7071) );
  INV_X1 U8927 ( .A(n7069), .ZN(n7070) );
  AND4_X1 U8928 ( .A1(n7073), .A2(n7072), .A3(n7071), .A4(n7070), .ZN(n7079)
         );
  NOR4_X1 U8929 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n7077) );
  NOR4_X1 U8930 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n7076) );
  NOR4_X1 U8931 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_27__SCAN_IN), .ZN(n7075) );
  NOR4_X1 U8932 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n7074) );
  AND4_X1 U8933 ( .A1(n7077), .A2(n7076), .A3(n7075), .A4(n7074), .ZN(n7078)
         );
  NAND2_X1 U8934 ( .A1(n7079), .A2(n7078), .ZN(n7080) );
  NAND2_X1 U8935 ( .A1(n10355), .A2(n7080), .ZN(n7612) );
  OR2_X1 U8936 ( .A1(n7617), .A2(n7941), .ZN(n7813) );
  NAND2_X1 U8937 ( .A1(n7612), .A2(n7615), .ZN(n7964) );
  INV_X1 U8938 ( .A(n7964), .ZN(n7088) );
  INV_X1 U8939 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n7081) );
  NAND2_X1 U8940 ( .A1(n10355), .A2(n7081), .ZN(n7084) );
  INV_X1 U8941 ( .A(n7082), .ZN(n8690) );
  NAND2_X1 U8942 ( .A1(n8574), .A2(n8690), .ZN(n7083) );
  NAND2_X1 U8943 ( .A1(n7084), .A2(n7083), .ZN(n7963) );
  INV_X1 U8944 ( .A(n7963), .ZN(n10224) );
  INV_X1 U8945 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n7085) );
  NAND2_X1 U8946 ( .A1(n10355), .A2(n7085), .ZN(n7087) );
  NAND2_X1 U8947 ( .A1(n8479), .A2(n8690), .ZN(n7086) );
  NAND3_X1 U8948 ( .A1(n7088), .A2(n10224), .A3(n7975), .ZN(n7156) );
  NAND2_X1 U8949 ( .A1(n7090), .A2(n8092), .ZN(n7932) );
  INV_X1 U8950 ( .A(n7932), .ZN(n7093) );
  AOI22_X1 U8951 ( .A1(n7932), .A2(n7929), .B1(n9805), .B2(n7873), .ZN(n7092)
         );
  NAND2_X1 U8952 ( .A1(n7094), .A2(n10380), .ZN(n7095) );
  NAND2_X1 U8953 ( .A1(n7934), .A2(n7095), .ZN(n8105) );
  NAND2_X1 U8954 ( .A1(n8052), .A2(n7096), .ZN(n8106) );
  NAND2_X1 U8955 ( .A1(n8105), .A2(n8106), .ZN(n7099) );
  NAND2_X1 U8956 ( .A1(n7097), .A2(n10388), .ZN(n7098) );
  NAND2_X1 U8957 ( .A1(n7099), .A2(n7098), .ZN(n8060) );
  NAND2_X1 U8958 ( .A1(n9802), .A2(n8246), .ZN(n8252) );
  AND2_X1 U8959 ( .A1(n8255), .A2(n8252), .ZN(n7100) );
  NAND2_X1 U8960 ( .A1(n8060), .A2(n7100), .ZN(n8075) );
  NAND3_X1 U8961 ( .A1(n8255), .A2(n8061), .A3(n8252), .ZN(n7104) );
  NAND2_X1 U8962 ( .A1(n8346), .A2(n8011), .ZN(n7103) );
  NAND2_X1 U8963 ( .A1(n7104), .A2(n7103), .ZN(n8073) );
  NAND2_X1 U8964 ( .A1(n8073), .A2(n8076), .ZN(n7106) );
  INV_X1 U8965 ( .A(n8286), .ZN(n9800) );
  NAND2_X1 U8966 ( .A1(n8286), .A2(n5491), .ZN(n7105) );
  INV_X1 U8967 ( .A(n8386), .ZN(n9799) );
  NAND2_X1 U8968 ( .A1(n10427), .A2(n9799), .ZN(n7109) );
  AND2_X1 U8969 ( .A1(n8535), .A2(n9798), .ZN(n7111) );
  OR2_X1 U8970 ( .A1(n8535), .A2(n9798), .ZN(n7110) );
  NAND2_X1 U8971 ( .A1(n8504), .A2(n8508), .ZN(n7113) );
  INV_X1 U8972 ( .A(n8533), .ZN(n9797) );
  OR2_X1 U8973 ( .A1(n8641), .A2(n9797), .ZN(n7112) );
  NAND2_X1 U8974 ( .A1(n7113), .A2(n7112), .ZN(n8619) );
  NOR2_X1 U8975 ( .A1(n10196), .A2(n9796), .ZN(n8618) );
  OR2_X1 U8976 ( .A1(n8618), .A2(n7114), .ZN(n7118) );
  NAND2_X1 U8977 ( .A1(n10196), .A2(n9796), .ZN(n8620) );
  INV_X1 U8978 ( .A(n10072), .ZN(n9795) );
  NAND2_X1 U8979 ( .A1(n10193), .A2(n9795), .ZN(n7115) );
  AND2_X1 U8980 ( .A1(n7116), .A2(n7115), .ZN(n7117) );
  AND2_X1 U8981 ( .A1(n10061), .A2(n9794), .ZN(n7119) );
  NOR2_X1 U8982 ( .A1(n10181), .A2(n10069), .ZN(n10033) );
  INV_X1 U8983 ( .A(n7120), .ZN(n7121) );
  AND2_X1 U8984 ( .A1(n4465), .A2(n7122), .ZN(n7126) );
  OR2_X1 U8985 ( .A1(n10033), .A2(n7126), .ZN(n10026) );
  NAND2_X1 U8986 ( .A1(n10170), .A2(n10012), .ZN(n7124) );
  NAND2_X1 U8987 ( .A1(n10181), .A2(n10069), .ZN(n10034) );
  AND2_X1 U8988 ( .A1(n7124), .A2(n10034), .ZN(n7125) );
  NOR2_X1 U8989 ( .A1(n7126), .A2(n7125), .ZN(n10027) );
  NAND2_X1 U8990 ( .A1(n10165), .A2(n5611), .ZN(n7128) );
  OR2_X1 U8991 ( .A1(n10159), .A2(n10013), .ZN(n7129) );
  NAND2_X1 U8992 ( .A1(n9995), .A2(n7129), .ZN(n7131) );
  NAND2_X1 U8993 ( .A1(n10159), .A2(n10013), .ZN(n7130) );
  NAND2_X1 U8994 ( .A1(n7131), .A2(n7130), .ZN(n9975) );
  NAND2_X1 U8995 ( .A1(n9975), .A2(n9976), .ZN(n7133) );
  NAND2_X1 U8996 ( .A1(n10156), .A2(n10003), .ZN(n7132) );
  NAND2_X1 U8997 ( .A1(n7133), .A2(n7132), .ZN(n9957) );
  OR2_X1 U8998 ( .A1(n10150), .A2(n9793), .ZN(n7134) );
  NAND2_X1 U8999 ( .A1(n9957), .A2(n7134), .ZN(n7136) );
  NAND2_X1 U9000 ( .A1(n10150), .A2(n9793), .ZN(n7135) );
  AND2_X1 U9001 ( .A1(n10146), .A2(n9970), .ZN(n7138) );
  INV_X1 U9002 ( .A(n9948), .ZN(n9921) );
  OR2_X1 U9003 ( .A1(n10134), .A2(n9903), .ZN(n7140) );
  NAND2_X1 U9004 ( .A1(n9909), .A2(n7140), .ZN(n7142) );
  NAND2_X1 U9005 ( .A1(n10134), .A2(n9903), .ZN(n7141) );
  OR2_X1 U9006 ( .A1(n10129), .A2(n9919), .ZN(n7143) );
  AND2_X1 U9007 ( .A1(n10127), .A2(n9905), .ZN(n7144) );
  NAND2_X1 U9008 ( .A1(n9867), .A2(n9869), .ZN(n7146) );
  OR2_X1 U9009 ( .A1(n10123), .A2(n9792), .ZN(n7145) );
  NAND2_X1 U9010 ( .A1(n7146), .A2(n7145), .ZN(n9855) );
  NOR2_X1 U9011 ( .A1(n10116), .A2(n9791), .ZN(n7148) );
  NAND2_X1 U9012 ( .A1(n10116), .A2(n9791), .ZN(n7147) );
  NAND2_X1 U9013 ( .A1(n10107), .A2(n9790), .ZN(n10097) );
  NAND2_X1 U9014 ( .A1(n10103), .A2(n10097), .ZN(n7151) );
  NAND2_X2 U9015 ( .A1(n7619), .A2(n7719), .ZN(n8836) );
  AND2_X1 U9016 ( .A1(n7966), .A2(n8836), .ZN(n7152) );
  NOR2_X4 U9017 ( .A1(n8379), .A2(n8535), .ZN(n8506) );
  INV_X1 U9018 ( .A(n8641), .ZN(n8507) );
  INV_X1 U9019 ( .A(n10181), .ZN(n8737) );
  NAND2_X1 U9020 ( .A1(n10057), .A2(n8737), .ZN(n8734) );
  OR2_X2 U9021 ( .A1(n8734), .A2(n10170), .ZN(n10048) );
  NOR2_X4 U9022 ( .A1(n10048), .A2(n10165), .ZN(n10017) );
  INV_X1 U9023 ( .A(n10159), .ZN(n10000) );
  INV_X1 U9024 ( .A(n10141), .ZN(n9936) );
  AND2_X2 U9025 ( .A1(n9950), .A2(n9936), .ZN(n9931) );
  INV_X1 U9026 ( .A(n10134), .ZN(n9916) );
  INV_X1 U9027 ( .A(n10123), .ZN(n9877) );
  AND2_X2 U9028 ( .A1(n9857), .A2(n9858), .ZN(n9859) );
  INV_X1 U9029 ( .A(n10107), .ZN(n8945) );
  NAND2_X1 U9030 ( .A1(n8250), .A2(n5946), .ZN(n7971) );
  OR2_X1 U9031 ( .A1(n7156), .A2(n9990), .ZN(n8643) );
  INV_X1 U9032 ( .A(n8643), .ZN(n10024) );
  NOR2_X1 U9033 ( .A1(n7971), .A2(n7993), .ZN(n7613) );
  INV_X1 U9034 ( .A(n10049), .ZN(n10059) );
  AOI22_X1 U9035 ( .A1(n7157), .A2(n10059), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n10020), .ZN(n7158) );
  OAI21_X1 U9036 ( .B1(n10095), .B2(n9999), .A(n7158), .ZN(n7159) );
  AOI21_X1 U9037 ( .B1(n10098), .B2(n10024), .A(n7159), .ZN(n7160) );
  NAND3_X1 U9038 ( .A1(n5044), .A2(n7161), .A3(n7160), .ZN(P1_U3355) );
  INV_X1 U9039 ( .A(n7317), .ZN(n7162) );
  INV_X1 U9040 ( .A(n9113), .ZN(n7165) );
  NAND2_X1 U9041 ( .A1(n7180), .A2(n6554), .ZN(n7173) );
  INV_X1 U9042 ( .A(n7166), .ZN(n7332) );
  INV_X1 U9043 ( .A(n7167), .ZN(n7168) );
  NAND2_X1 U9044 ( .A1(n4386), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n7171) );
  NAND2_X1 U9045 ( .A1(n6257), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n7170) );
  OAI211_X1 U9046 ( .C1(n7172), .C2(n6760), .A(n7171), .B(n7170), .ZN(n9112)
         );
  NAND2_X1 U9047 ( .A1(n8900), .A2(n9112), .ZN(n7371) );
  NAND2_X1 U9048 ( .A1(n7174), .A2(n7173), .ZN(n7175) );
  NAND2_X1 U9049 ( .A1(n9617), .A2(n7176), .ZN(n7179) );
  NAND2_X1 U9050 ( .A1(n7177), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n7178) );
  NOR2_X1 U9051 ( .A1(n9478), .A2(n7180), .ZN(n7337) );
  INV_X1 U9052 ( .A(n9112), .ZN(n7181) );
  AND2_X1 U9053 ( .A1(n7182), .A2(n7181), .ZN(n7331) );
  NOR2_X1 U9054 ( .A1(n7337), .A2(n7331), .ZN(n7374) );
  INV_X1 U9055 ( .A(n9478), .ZN(n9199) );
  XNOR2_X1 U9056 ( .A(n7183), .B(n4944), .ZN(n7186) );
  INV_X1 U9057 ( .A(n7184), .ZN(n7185) );
  INV_X1 U9058 ( .A(n7187), .ZN(n10488) );
  INV_X1 U9059 ( .A(n6584), .ZN(n7346) );
  INV_X1 U9060 ( .A(n7188), .ZN(n7191) );
  NAND2_X1 U9061 ( .A1(n7194), .A2(n7188), .ZN(n7356) );
  NAND2_X1 U9062 ( .A1(n7213), .A2(n7750), .ZN(n7357) );
  INV_X1 U9063 ( .A(n7214), .ZN(n7190) );
  OAI21_X1 U9064 ( .B1(n7192), .B2(n7191), .A(n7190), .ZN(n7195) );
  NAND3_X1 U9065 ( .A1(n7195), .A2(n7194), .A3(n7193), .ZN(n7210) );
  NAND2_X1 U9066 ( .A1(n6592), .A2(n10463), .ZN(n10456) );
  INV_X1 U9067 ( .A(n7196), .ZN(n7198) );
  INV_X1 U9068 ( .A(n7197), .ZN(n7204) );
  AOI211_X1 U9069 ( .C1(n7353), .C2(n10456), .A(n7198), .B(n7204), .ZN(n7200)
         );
  INV_X1 U9070 ( .A(n7199), .ZN(n7202) );
  NOR2_X1 U9071 ( .A1(n7200), .A2(n7202), .ZN(n7207) );
  AOI21_X1 U9072 ( .B1(n6554), .B2(n10456), .A(n7352), .ZN(n7203) );
  INV_X1 U9073 ( .A(n7353), .ZN(n7201) );
  NOR3_X1 U9074 ( .A1(n7203), .A2(n7202), .A3(n7201), .ZN(n7205) );
  NOR2_X1 U9075 ( .A1(n7205), .A2(n7204), .ZN(n7206) );
  NOR2_X1 U9076 ( .A1(n8180), .A2(n7218), .ZN(n7217) );
  INV_X1 U9077 ( .A(n7357), .ZN(n7212) );
  AOI22_X1 U9078 ( .A1(n7214), .A2(n7213), .B1(n7212), .B2(n7211), .ZN(n7215)
         );
  NOR2_X1 U9079 ( .A1(n7215), .A2(n7217), .ZN(n7216) );
  NAND3_X1 U9080 ( .A1(n8180), .A2(n7218), .A3(n7340), .ZN(n7220) );
  AND2_X1 U9081 ( .A1(n7220), .A2(n7219), .ZN(n7221) );
  MUX2_X1 U9082 ( .A(n8126), .B(n9121), .S(n7339), .Z(n7223) );
  MUX2_X1 U9083 ( .A(n8541), .B(n7225), .S(n7339), .Z(n7226) );
  NAND2_X1 U9084 ( .A1(n7233), .A2(n7235), .ZN(n7230) );
  INV_X1 U9085 ( .A(n7228), .ZN(n7229) );
  MUX2_X1 U9086 ( .A(n7230), .B(n7229), .S(n7339), .Z(n7231) );
  INV_X1 U9087 ( .A(n7232), .ZN(n7236) );
  NOR2_X1 U9088 ( .A1(n7231), .A2(n7236), .ZN(n7240) );
  NAND2_X1 U9089 ( .A1(n8651), .A2(n7232), .ZN(n7238) );
  OAI211_X1 U9090 ( .C1(n7236), .C2(n7235), .A(n7234), .B(n7233), .ZN(n7237)
         );
  MUX2_X1 U9091 ( .A(n7238), .B(n7237), .S(n7339), .Z(n7239) );
  INV_X1 U9092 ( .A(n7241), .ZN(n7247) );
  INV_X1 U9093 ( .A(n7243), .ZN(n7251) );
  NOR2_X1 U9094 ( .A1(n7247), .A2(n7339), .ZN(n7248) );
  OAI211_X1 U9095 ( .C1(n7249), .C2(n8650), .A(n7248), .B(n7253), .ZN(n7256)
         );
  NOR2_X1 U9096 ( .A1(n7253), .A2(n7340), .ZN(n7250) );
  AOI21_X1 U9097 ( .B1(n7340), .B2(n7251), .A(n7250), .ZN(n7255) );
  NAND3_X1 U9098 ( .A1(n7253), .A2(n7252), .A3(n7340), .ZN(n7254) );
  NAND4_X1 U9099 ( .A1(n7256), .A2(n6544), .A3(n7255), .A4(n7254), .ZN(n7260)
         );
  MUX2_X1 U9100 ( .A(n7258), .B(n7257), .S(n7339), .Z(n7259) );
  OAI21_X1 U9101 ( .B1(n7261), .B2(n7260), .A(n7259), .ZN(n7262) );
  INV_X1 U9102 ( .A(n7263), .ZN(n7266) );
  INV_X1 U9103 ( .A(n7264), .ZN(n7265) );
  MUX2_X1 U9104 ( .A(n7266), .B(n7265), .S(n7339), .Z(n7267) );
  INV_X1 U9105 ( .A(n7268), .ZN(n7270) );
  MUX2_X1 U9106 ( .A(n7270), .B(n7269), .S(n7339), .Z(n7271) );
  NAND2_X1 U9107 ( .A1(n7279), .A2(n7274), .ZN(n7277) );
  INV_X1 U9108 ( .A(n7275), .ZN(n7276) );
  MUX2_X1 U9109 ( .A(n7277), .B(n7276), .S(n7340), .Z(n7278) );
  INV_X1 U9110 ( .A(n7279), .ZN(n7280) );
  OAI211_X1 U9111 ( .C1(n7285), .C2(n7280), .A(n7287), .B(n7350), .ZN(n7284)
         );
  INV_X1 U9112 ( .A(n7281), .ZN(n7282) );
  INV_X1 U9113 ( .A(n7348), .ZN(n9279) );
  INV_X1 U9114 ( .A(n7286), .ZN(n7351) );
  AOI21_X1 U9115 ( .B1(n7288), .B2(n7287), .A(n7351), .ZN(n7290) );
  OAI211_X1 U9116 ( .C1(n7290), .C2(n7289), .A(n7349), .B(n9278), .ZN(n7292)
         );
  MUX2_X1 U9117 ( .A(n7295), .B(n7294), .S(n7339), .Z(n7296) );
  INV_X1 U9118 ( .A(n9114), .ZN(n9265) );
  NAND2_X1 U9119 ( .A1(n9508), .A2(n9265), .ZN(n7298) );
  MUX2_X1 U9120 ( .A(n7298), .B(n7297), .S(n7339), .Z(n7299) );
  NAND3_X1 U9121 ( .A1(n7300), .A2(n9228), .A3(n7299), .ZN(n7306) );
  INV_X1 U9122 ( .A(n7311), .ZN(n7303) );
  INV_X1 U9123 ( .A(n7301), .ZN(n7302) );
  OAI21_X1 U9124 ( .B1(n7303), .B2(n7302), .A(n7339), .ZN(n7305) );
  INV_X1 U9125 ( .A(n7309), .ZN(n7304) );
  AOI21_X1 U9126 ( .B1(n7306), .B2(n7305), .A(n7304), .ZN(n7307) );
  INV_X1 U9127 ( .A(n7307), .ZN(n7314) );
  AOI21_X1 U9128 ( .B1(n7309), .B2(n7308), .A(n7339), .ZN(n7310) );
  INV_X1 U9129 ( .A(n7310), .ZN(n7313) );
  NAND3_X1 U9130 ( .A1(n9493), .A2(n7315), .A3(n7339), .ZN(n7316) );
  OAI211_X1 U9131 ( .C1(n7318), .C2(n7339), .A(n7317), .B(n7316), .ZN(n7319)
         );
  NOR2_X1 U9132 ( .A1(n9488), .A2(n7340), .ZN(n7322) );
  OAI211_X1 U9133 ( .C1(n7324), .C2(n9204), .A(n7332), .B(n7336), .ZN(n7329)
         );
  NOR4_X1 U9134 ( .A1(n7325), .A2(n7330), .A3(n7174), .A4(n7340), .ZN(n7328)
         );
  INV_X1 U9135 ( .A(n7325), .ZN(n7372) );
  NOR2_X1 U9136 ( .A1(n7372), .A2(n7339), .ZN(n7327) );
  NOR4_X1 U9137 ( .A1(n7325), .A2(n8900), .A3(n7340), .A4(n9112), .ZN(n7326)
         );
  INV_X1 U9138 ( .A(n7330), .ZN(n7335) );
  INV_X1 U9139 ( .A(n7331), .ZN(n7333) );
  NAND3_X1 U9140 ( .A1(n7333), .A2(n7340), .A3(n7332), .ZN(n7334) );
  INV_X1 U9141 ( .A(n7337), .ZN(n7341) );
  NAND2_X1 U9142 ( .A1(n7338), .A2(n7341), .ZN(n7344) );
  NAND3_X1 U9143 ( .A1(n9199), .A2(n7431), .A3(n7339), .ZN(n7343) );
  NAND4_X1 U9144 ( .A1(n7341), .A2(n8900), .A3(n7340), .A4(n9112), .ZN(n7342)
         );
  NAND4_X1 U9145 ( .A1(n7345), .A2(n7344), .A3(n7343), .A4(n7342), .ZN(n7347)
         );
  OAI21_X1 U9146 ( .B1(n7347), .B2(n7346), .A(n7981), .ZN(n7377) );
  INV_X1 U9147 ( .A(n8908), .ZN(n7370) );
  NAND2_X1 U9148 ( .A1(n7349), .A2(n4518), .ZN(n9306) );
  INV_X1 U9149 ( .A(n8653), .ZN(n8663) );
  INV_X1 U9150 ( .A(n7352), .ZN(n7354) );
  AND2_X1 U9151 ( .A1(n7354), .A2(n7353), .ZN(n7667) );
  NAND4_X1 U9152 ( .A1(n7667), .A2(n7839), .A3(n7355), .A4(n10456), .ZN(n7358)
         );
  NOR4_X1 U9153 ( .A1(n7358), .A2(n6525), .A3(n7357), .A4(n7356), .ZN(n7359)
         );
  NAND4_X1 U9154 ( .A1(n7359), .A2(n8218), .A3(n8544), .A4(n4422), .ZN(n7360)
         );
  INV_X1 U9155 ( .A(n8299), .ZN(n8293) );
  NOR4_X1 U9156 ( .A1(n7360), .A2(n8227), .A3(n8121), .A4(n8293), .ZN(n7361)
         );
  NAND4_X1 U9157 ( .A1(n6544), .A2(n9424), .A3(n8663), .A4(n7361), .ZN(n7362)
         );
  NOR4_X1 U9158 ( .A1(n9357), .A2(n9378), .A3(n7363), .A4(n7362), .ZN(n7364)
         );
  NAND4_X1 U9159 ( .A1(n7365), .A2(n9352), .A3(n9340), .A4(n7364), .ZN(n7366)
         );
  NOR4_X1 U9160 ( .A1(n9261), .A2(n6549), .A3(n9306), .A4(n7366), .ZN(n7367)
         );
  NAND4_X1 U9161 ( .A1(n9219), .A2(n9228), .A3(n7367), .A4(n9250), .ZN(n7368)
         );
  NOR4_X1 U9162 ( .A1(n7370), .A2(n7369), .A3(n9209), .A4(n7368), .ZN(n7373)
         );
  NAND4_X1 U9163 ( .A1(n7374), .A2(n7373), .A3(n7372), .A4(n7371), .ZN(n7375)
         );
  NOR4_X1 U9164 ( .A1(n10472), .A2(n9418), .A3(n8695), .A4(n7378), .ZN(n7381)
         );
  OAI21_X1 U9165 ( .B1(n7379), .B2(n6553), .A(P2_B_REG_SCAN_IN), .ZN(n7380) );
  OR2_X1 U9166 ( .A1(n7381), .A2(n7380), .ZN(n7382) );
  INV_X1 U9167 ( .A(n9125), .ZN(P2_U3966) );
  OR2_X2 U9168 ( .A1(n7383), .A2(P1_U3084), .ZN(n9807) );
  INV_X1 U9169 ( .A(n9807), .ZN(P1_U4006) );
  NOR2_X1 U9170 ( .A1(n7388), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9621) );
  NAND2_X1 U9171 ( .A1(n7388), .A2(P2_U3152), .ZN(n9627) );
  OAI222_X1 U9172 ( .A1(n9624), .A2(n7385), .B1(n9627), .B2(n4676), .C1(
        P2_U3152), .C2(n7581), .ZN(P2_U3356) );
  INV_X1 U9173 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n7386) );
  OAI222_X1 U9174 ( .A1(n9624), .A2(n7386), .B1(n9627), .B2(n7398), .C1(
        P2_U3152), .C2(n7568), .ZN(P2_U3357) );
  OAI222_X1 U9175 ( .A1(n9624), .A2(n7387), .B1(n9627), .B2(n7391), .C1(
        P2_U3152), .C2(n6044), .ZN(P2_U3355) );
  AND2_X1 U9176 ( .A1(n5398), .A2(P1_U3084), .ZN(n8330) );
  INV_X1 U9177 ( .A(n7390), .ZN(n10274) );
  OAI222_X1 U9178 ( .A1(n10238), .A2(n7392), .B1(n4391), .B2(n7391), .C1(
        P1_U3084), .C2(n10274), .ZN(P1_U3350) );
  INV_X1 U9179 ( .A(n7393), .ZN(n7394) );
  OAI222_X1 U9180 ( .A1(n9624), .A2(n5219), .B1(n9627), .B2(n7394), .C1(
        P2_U3152), .C2(n7611), .ZN(P2_U3354) );
  INV_X1 U9181 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7395) );
  OAI222_X1 U9182 ( .A1(n10238), .A2(n7395), .B1(n4391), .B2(n7394), .C1(
        P1_U3084), .C2(n7701), .ZN(P1_U3349) );
  INV_X1 U9183 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7397) );
  OAI222_X1 U9184 ( .A1(n5010), .A2(P1_U3084), .B1(n4391), .B2(n7398), .C1(
        n7397), .C2(n10238), .ZN(P1_U3352) );
  INV_X1 U9185 ( .A(n7399), .ZN(n10298) );
  OAI222_X1 U9186 ( .A1(n10298), .A2(P1_U3084), .B1(n4391), .B2(n4676), .C1(
        n7400), .C2(n10238), .ZN(P1_U3351) );
  INV_X1 U9187 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7402) );
  INV_X1 U9188 ( .A(n7401), .ZN(n7405) );
  INV_X1 U9189 ( .A(n7550), .ZN(n7557) );
  OAI222_X1 U9190 ( .A1(n9624), .A2(n7402), .B1(n9627), .B2(n7405), .C1(
        P2_U3152), .C2(n7557), .ZN(P2_U3353) );
  INV_X1 U9191 ( .A(n7403), .ZN(n7408) );
  INV_X1 U9192 ( .A(n10238), .ZN(n10229) );
  AOI22_X1 U9193 ( .A1(n9818), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n10229), .ZN(n7404) );
  OAI21_X1 U9194 ( .B1(n7408), .B2(n4391), .A(n7404), .ZN(P1_U3347) );
  INV_X1 U9195 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7406) );
  OAI222_X1 U9196 ( .A1(n10238), .A2(n7406), .B1(n4391), .B2(n7405), .C1(
        P1_U3084), .C2(n7451), .ZN(P1_U3348) );
  INV_X1 U9197 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7409) );
  OAI222_X1 U9198 ( .A1(n9624), .A2(n7409), .B1(n9627), .B2(n7408), .C1(
        P2_U3152), .C2(n7407), .ZN(P2_U3352) );
  INV_X1 U9199 ( .A(n9627), .ZN(n8714) );
  INV_X1 U9200 ( .A(n8714), .ZN(n8956) );
  INV_X1 U9201 ( .A(n7410), .ZN(n7414) );
  INV_X1 U9202 ( .A(n7411), .ZN(n8042) );
  OAI222_X1 U9203 ( .A1(n8956), .A2(n7414), .B1(n8042), .B2(P2_U3152), .C1(
        n7412), .C2(n9624), .ZN(P2_U3349) );
  OAI222_X1 U9204 ( .A1(n10238), .A2(n7415), .B1(n4391), .B2(n7414), .C1(n7413), .C2(P1_U3084), .ZN(P1_U3344) );
  INV_X1 U9205 ( .A(n6236), .ZN(n7417) );
  OAI222_X1 U9206 ( .A1(n9624), .A2(n4539), .B1(n9627), .B2(n7417), .C1(
        P2_U3152), .C2(n7649), .ZN(P2_U3351) );
  INV_X1 U9207 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7418) );
  INV_X1 U9208 ( .A(n7488), .ZN(n7416) );
  OAI222_X1 U9209 ( .A1(n10238), .A2(n7418), .B1(n4391), .B2(n7417), .C1(
        P1_U3084), .C2(n7416), .ZN(P1_U3346) );
  INV_X1 U9210 ( .A(n7419), .ZN(n7426) );
  OAI222_X1 U9211 ( .A1(n8956), .A2(n7426), .B1(n8356), .B2(P2_U3152), .C1(
        n7420), .C2(n9624), .ZN(P2_U3348) );
  INV_X1 U9212 ( .A(n7421), .ZN(n7423) );
  INV_X1 U9213 ( .A(n7462), .ZN(n7461) );
  OAI222_X1 U9214 ( .A1(n10238), .A2(n7422), .B1(n4391), .B2(n7423), .C1(
        P1_U3084), .C2(n7461), .ZN(P1_U3345) );
  OAI222_X1 U9215 ( .A1(n9624), .A2(n7424), .B1(n8956), .B2(n7423), .C1(
        P2_U3152), .C2(n7856), .ZN(P2_U3350) );
  NOR2_X1 U9216 ( .A1(n9174), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U9217 ( .A(n7425), .ZN(n7502) );
  OAI222_X1 U9218 ( .A1(n10238), .A2(n7427), .B1(n4391), .B2(n7426), .C1(n7502), .C2(P1_U3084), .ZN(P1_U3343) );
  INV_X1 U9219 ( .A(n7428), .ZN(n7435) );
  INV_X1 U9220 ( .A(n7429), .ZN(n8489) );
  OAI222_X1 U9221 ( .A1(n8956), .A2(n7435), .B1(n8489), .B2(P2_U3152), .C1(
        n7430), .C2(n9624), .ZN(P2_U3347) );
  INV_X1 U9222 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n7433) );
  NAND2_X1 U9223 ( .A1(P2_U3966), .A2(n7431), .ZN(n7432) );
  OAI21_X1 U9224 ( .B1(P2_U3966), .B2(n7433), .A(n7432), .ZN(P2_U3583) );
  OAI222_X1 U9225 ( .A1(n10238), .A2(n7436), .B1(n4391), .B2(n7435), .C1(n7434), .C2(P1_U3084), .ZN(P1_U3342) );
  INV_X1 U9226 ( .A(n10342), .ZN(n7900) );
  INV_X1 U9227 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7447) );
  INV_X1 U9228 ( .A(n7437), .ZN(n7439) );
  NAND2_X1 U9229 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n7683) );
  AOI211_X1 U9230 ( .C1(n7439), .C2(n7683), .A(n7438), .B(n10305), .ZN(n7445)
         );
  NAND2_X1 U9231 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n7441) );
  AOI211_X1 U9232 ( .C1(n7442), .C2(n7441), .A(n7440), .B(n10300), .ZN(n7444)
         );
  INV_X1 U9233 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7729) );
  OAI22_X1 U9234 ( .A1(n10339), .A2(n5010), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7729), .ZN(n7443) );
  NOR3_X1 U9235 ( .A1(n7445), .A2(n7444), .A3(n7443), .ZN(n7446) );
  OAI21_X1 U9236 ( .B1(n7900), .B2(n7447), .A(n7446), .ZN(P1_U3242) );
  INV_X1 U9237 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7460) );
  AOI211_X1 U9238 ( .C1(n7450), .C2(n7449), .A(n10300), .B(n7448), .ZN(n7458)
         );
  AND2_X1 U9239 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n8243) );
  NOR2_X1 U9240 ( .A1(n10339), .A2(n7451), .ZN(n7457) );
  OR3_X1 U9241 ( .A1(n7692), .A2(n7453), .A3(n7452), .ZN(n7454) );
  AOI21_X1 U9242 ( .B1(n7455), .B2(n7454), .A(n10305), .ZN(n7456) );
  NOR4_X1 U9243 ( .A1(n7458), .A2(n8243), .A3(n7457), .A4(n7456), .ZN(n7459)
         );
  OAI21_X1 U9244 ( .B1(n7900), .B2(n7460), .A(n7459), .ZN(P1_U3246) );
  NAND2_X1 U9245 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8284) );
  OAI21_X1 U9246 ( .B1(n10339), .B2(n7461), .A(n8284), .ZN(n7468) );
  INV_X1 U9247 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10453) );
  MUX2_X1 U9248 ( .A(n10453), .B(P1_REG1_REG_8__SCAN_IN), .S(n7462), .Z(n7466)
         );
  NAND2_X1 U9249 ( .A1(n7489), .A2(n7463), .ZN(n7465) );
  INV_X1 U9250 ( .A(n7523), .ZN(n7464) );
  AOI211_X1 U9251 ( .C1(n7466), .C2(n7465), .A(n10300), .B(n7464), .ZN(n7467)
         );
  AOI211_X1 U9252 ( .C1(n10342), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n7468), .B(
        n7467), .ZN(n7475) );
  INV_X1 U9253 ( .A(n7469), .ZN(n7473) );
  NOR3_X1 U9254 ( .A1(n7485), .A2(n7471), .A3(n7470), .ZN(n7472) );
  OAI21_X1 U9255 ( .B1(n7473), .B2(n7472), .A(n10348), .ZN(n7474) );
  NAND2_X1 U9256 ( .A1(n7475), .A2(n7474), .ZN(P1_U3249) );
  INV_X1 U9257 ( .A(n6314), .ZN(n7479) );
  INV_X1 U9258 ( .A(n7476), .ZN(n8706) );
  OAI222_X1 U9259 ( .A1(n9624), .A2(n7477), .B1(n8956), .B2(n7479), .C1(
        P2_U3152), .C2(n8706), .ZN(P2_U3346) );
  OAI222_X1 U9260 ( .A1(n10238), .A2(n7480), .B1(n4391), .B2(n7479), .C1(
        P1_U3084), .C2(n7478), .ZN(P1_U3341) );
  INV_X1 U9261 ( .A(n7481), .ZN(n7497) );
  INV_X1 U9262 ( .A(n7482), .ZN(n8728) );
  OAI222_X1 U9263 ( .A1(n8956), .A2(n7497), .B1(n8728), .B2(P2_U3152), .C1(
        n7483), .C2(n9624), .ZN(P2_U3345) );
  INV_X1 U9264 ( .A(n7484), .ZN(n7486) );
  AOI21_X1 U9265 ( .B1(n4493), .B2(n7486), .A(n7485), .ZN(n7496) );
  INV_X1 U9266 ( .A(n10339), .ZN(n10317) );
  AND2_X1 U9267 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n8032) );
  INV_X1 U9268 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10259) );
  NOR2_X1 U9269 ( .A1(n7900), .A2(n10259), .ZN(n7487) );
  AOI211_X1 U9270 ( .C1(n10317), .C2(n7488), .A(n8032), .B(n7487), .ZN(n7495)
         );
  INV_X1 U9271 ( .A(n7489), .ZN(n7493) );
  NOR3_X1 U9272 ( .A1(n9809), .A2(n7491), .A3(n7490), .ZN(n7492) );
  OAI21_X1 U9273 ( .B1(n7493), .B2(n7492), .A(n10344), .ZN(n7494) );
  OAI211_X1 U9274 ( .C1(n7496), .C2(n10305), .A(n7495), .B(n7494), .ZN(
        P1_U3248) );
  OAI222_X1 U9275 ( .A1(n10238), .A2(n7498), .B1(n4391), .B2(n7497), .C1(n8140), .C2(P1_U3084), .ZN(P1_U3340) );
  NAND3_X1 U9276 ( .A1(n7516), .A2(n7500), .A3(n7499), .ZN(n7501) );
  NAND2_X1 U9277 ( .A1(n7501), .A2(n10348), .ZN(n7510) );
  NAND2_X1 U9278 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8417) );
  OAI21_X1 U9279 ( .B1(n10339), .B2(n7502), .A(n8417), .ZN(n7508) );
  INV_X1 U9280 ( .A(n7655), .ZN(n7506) );
  NAND3_X1 U9281 ( .A1(n7520), .A2(n7504), .A3(n7503), .ZN(n7505) );
  AOI21_X1 U9282 ( .B1(n7506), .B2(n7505), .A(n10300), .ZN(n7507) );
  AOI211_X1 U9283 ( .C1(n10342), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n7508), .B(
        n7507), .ZN(n7509) );
  OAI21_X1 U9284 ( .B1(n7511), .B2(n7510), .A(n7509), .ZN(P1_U3251) );
  INV_X1 U9285 ( .A(n7512), .ZN(n7514) );
  OAI222_X1 U9286 ( .A1(n8956), .A2(n7514), .B1(n9133), .B2(P2_U3152), .C1(
        n7513), .C2(n9624), .ZN(P2_U3344) );
  OAI222_X1 U9287 ( .A1(n10238), .A2(n7515), .B1(n4391), .B2(n7514), .C1(n8425), .C2(P1_U3084), .ZN(P1_U3339) );
  INV_X1 U9288 ( .A(n7516), .ZN(n7517) );
  AOI211_X1 U9289 ( .C1(n7519), .C2(n7518), .A(n10305), .B(n7517), .ZN(n7531)
         );
  INV_X1 U9290 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10565) );
  INV_X1 U9291 ( .A(n7520), .ZN(n7525) );
  AOI21_X1 U9292 ( .B1(n7523), .B2(n7522), .A(n7521), .ZN(n7524) );
  OAI21_X1 U9293 ( .B1(n7525), .B2(n7524), .A(n10344), .ZN(n7529) );
  NOR2_X1 U9294 ( .A1(n7526), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8530) );
  AOI21_X1 U9295 ( .B1(n10317), .B2(n7527), .A(n8530), .ZN(n7528) );
  OAI211_X1 U9296 ( .C1(n10565), .C2(n7900), .A(n7529), .B(n7528), .ZN(n7530)
         );
  OR2_X1 U9297 ( .A1(n7531), .A2(n7530), .ZN(P1_U3250) );
  AOI211_X1 U9298 ( .C1(n7534), .C2(n7533), .A(n7532), .B(n9184), .ZN(n7545)
         );
  INV_X1 U9299 ( .A(n7535), .ZN(n7578) );
  INV_X1 U9300 ( .A(n7536), .ZN(n7539) );
  MUX2_X1 U9301 ( .A(n6133), .B(P2_REG1_REG_3__SCAN_IN), .S(n7537), .Z(n7538)
         );
  NAND3_X1 U9302 ( .A1(n7578), .A2(n7539), .A3(n7538), .ZN(n7540) );
  NAND3_X1 U9303 ( .A1(n9169), .A2(n7604), .A3(n7540), .ZN(n7543) );
  NOR2_X1 U9304 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9462), .ZN(n7541) );
  AOI21_X1 U9305 ( .B1(n9174), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n7541), .ZN(
        n7542) );
  OAI211_X1 U9306 ( .C1(n9178), .C2(n6044), .A(n7543), .B(n7542), .ZN(n7544)
         );
  OR2_X1 U9307 ( .A1(n7545), .A2(n7544), .ZN(P2_U3248) );
  AOI211_X1 U9308 ( .C1(n7548), .C2(n7547), .A(n9184), .B(n7546), .ZN(n7559)
         );
  INV_X1 U9309 ( .A(n7549), .ZN(n7552) );
  MUX2_X1 U9310 ( .A(n7866), .B(P2_REG1_REG_5__SCAN_IN), .S(n7550), .Z(n7551)
         );
  NAND2_X1 U9311 ( .A1(n7552), .A2(n7551), .ZN(n7553) );
  OAI211_X1 U9312 ( .C1(n7606), .C2(n7553), .A(n9169), .B(n7586), .ZN(n7556)
         );
  AND2_X1 U9313 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7554) );
  AOI21_X1 U9314 ( .B1(n9174), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n7554), .ZN(
        n7555) );
  OAI211_X1 U9315 ( .C1(n9178), .C2(n7557), .A(n7556), .B(n7555), .ZN(n7558)
         );
  OR2_X1 U9316 ( .A1(n7559), .A2(n7558), .ZN(P2_U3250) );
  AOI211_X1 U9317 ( .C1(n7562), .C2(n7561), .A(n7560), .B(n9184), .ZN(n7570)
         );
  INV_X1 U9318 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10517) );
  MUX2_X1 U9319 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6130), .S(n7568), .Z(n7563)
         );
  OAI21_X1 U9320 ( .B1(n10517), .B2(n7564), .A(n7563), .ZN(n7565) );
  NAND3_X1 U9321 ( .A1(n9169), .A2(n7576), .A3(n7565), .ZN(n7567) );
  AOI22_X1 U9322 ( .A1(n9174), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n7566) );
  OAI211_X1 U9323 ( .C1(n9178), .C2(n7568), .A(n7567), .B(n7566), .ZN(n7569)
         );
  OR2_X1 U9324 ( .A1(n7570), .A2(n7569), .ZN(P2_U3246) );
  AOI211_X1 U9325 ( .C1(n7573), .C2(n7572), .A(n7571), .B(n9184), .ZN(n7583)
         );
  NAND3_X1 U9326 ( .A1(n7576), .A2(n7575), .A3(n7574), .ZN(n7577) );
  NAND3_X1 U9327 ( .A1(n9169), .A2(n7578), .A3(n7577), .ZN(n7580) );
  AOI22_X1 U9328 ( .A1(n9174), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n7579) );
  OAI211_X1 U9329 ( .C1(n9178), .C2(n7581), .A(n7580), .B(n7579), .ZN(n7582)
         );
  OR2_X1 U9330 ( .A1(n7583), .A2(n7582), .ZN(P2_U3247) );
  INV_X1 U9331 ( .A(n9178), .ZN(n9193) );
  INV_X1 U9332 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7590) );
  INV_X1 U9333 ( .A(n7643), .ZN(n7588) );
  NAND3_X1 U9334 ( .A1(n7586), .A2(n7585), .A3(n7584), .ZN(n7587) );
  NAND3_X1 U9335 ( .A1(n9169), .A2(n7588), .A3(n7587), .ZN(n7589) );
  NAND2_X1 U9336 ( .A1(P2_U3152), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7914) );
  OAI211_X1 U9337 ( .C1(n9190), .C2(n7590), .A(n7589), .B(n7914), .ZN(n7595)
         );
  AOI211_X1 U9338 ( .C1(n7593), .C2(n7592), .A(n9184), .B(n7591), .ZN(n7594)
         );
  AOI211_X1 U9339 ( .C1(n9193), .C2(n7596), .A(n7595), .B(n7594), .ZN(n7597)
         );
  INV_X1 U9340 ( .A(n7597), .ZN(P2_U3251) );
  AOI211_X1 U9341 ( .C1(n7600), .C2(n7599), .A(n7598), .B(n9184), .ZN(n7601)
         );
  INV_X1 U9342 ( .A(n7601), .ZN(n7610) );
  AND2_X1 U9343 ( .A1(P2_U3152), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7608) );
  AND3_X1 U9344 ( .A1(n7604), .A2(n7603), .A3(n7602), .ZN(n7605) );
  NOR3_X1 U9345 ( .A1(n9196), .A2(n7606), .A3(n7605), .ZN(n7607) );
  AOI211_X1 U9346 ( .C1(n9174), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n7608), .B(
        n7607), .ZN(n7609) );
  OAI211_X1 U9347 ( .C1(n9178), .C2(n7611), .A(n7610), .B(n7609), .ZN(P2_U3249) );
  NAND3_X1 U9348 ( .A1(n10226), .A2(n10224), .A3(n7612), .ZN(n7628) );
  INV_X1 U9349 ( .A(n7613), .ZN(n7728) );
  INV_X1 U9350 ( .A(n10225), .ZN(n10354) );
  NOR2_X1 U9351 ( .A1(n7728), .A2(n10354), .ZN(n7614) );
  NAND2_X1 U9352 ( .A1(n7628), .A2(n7614), .ZN(n7817) );
  OR2_X1 U9353 ( .A1(n7628), .A2(n7966), .ZN(n7819) );
  NAND2_X1 U9354 ( .A1(n10225), .A2(n7684), .ZN(n7616) );
  NAND3_X1 U9355 ( .A1(n10225), .A2(n7617), .A3(n10400), .ZN(n7618) );
  INV_X1 U9356 ( .A(n8865), .ZN(n7621) );
  NAND2_X1 U9357 ( .A1(n7621), .A2(n9808), .ZN(n7623) );
  NAND2_X1 U9358 ( .A1(n9808), .A2(n8004), .ZN(n7626) );
  AOI22_X1 U9359 ( .A1(n8439), .A2(n7982), .B1(n7624), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n7625) );
  NAND2_X1 U9360 ( .A1(n7626), .A2(n7625), .ZN(n7790) );
  NAND2_X1 U9361 ( .A1(n7627), .A2(n7790), .ZN(n7792) );
  OAI21_X1 U9362 ( .B1(n7627), .B2(n7790), .A(n7792), .ZN(n7685) );
  AOI22_X1 U9363 ( .A1(n9780), .A2(n9806), .B1(n9772), .B2(n7685), .ZN(n7630)
         );
  NAND2_X1 U9364 ( .A1(n7628), .A2(n10400), .ZN(n7814) );
  AND2_X1 U9365 ( .A1(n8347), .A2(n7814), .ZN(n7878) );
  INV_X1 U9366 ( .A(n7878), .ZN(n8927) );
  NAND2_X1 U9367 ( .A1(n8927), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n7629) );
  OAI211_X1 U9368 ( .C1(n9771), .C2(n7972), .A(n7630), .B(n7629), .ZN(P1_U3230) );
  INV_X1 U9369 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7631) );
  OAI211_X1 U9370 ( .C1(n9196), .C2(P2_REG1_REG_0__SCAN_IN), .A(
        P2_IR_REG_0__SCAN_IN), .B(n9178), .ZN(n7632) );
  AOI21_X1 U9371 ( .B1(n9163), .B2(n7631), .A(n7632), .ZN(n7636) );
  AOI21_X1 U9372 ( .B1(n9169), .B2(P2_REG1_REG_0__SCAN_IN), .A(
        P2_IR_REG_0__SCAN_IN), .ZN(n7635) );
  AOI22_X1 U9373 ( .A1(n9174), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n7634) );
  NAND3_X1 U9374 ( .A1(n7632), .A2(n9163), .A3(P2_REG2_REG_0__SCAN_IN), .ZN(
        n7633) );
  OAI211_X1 U9375 ( .C1(n7636), .C2(n7635), .A(n7634), .B(n7633), .ZN(P2_U3245) );
  AOI211_X1 U9376 ( .C1(n4492), .C2(n7638), .A(n9184), .B(n7637), .ZN(n7639)
         );
  INV_X1 U9377 ( .A(n7639), .ZN(n7648) );
  AND2_X1 U9378 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7906) );
  MUX2_X1 U9379 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10524), .S(n7640), .Z(n7641)
         );
  NOR3_X1 U9380 ( .A1(n7643), .A2(n7642), .A3(n7641), .ZN(n7644) );
  NOR3_X1 U9381 ( .A1(n7645), .A2(n7644), .A3(n9196), .ZN(n7646) );
  AOI211_X1 U9382 ( .C1(n9174), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n7906), .B(
        n7646), .ZN(n7647) );
  OAI211_X1 U9383 ( .C1(n9178), .C2(n7649), .A(n7648), .B(n7647), .ZN(P2_U3252) );
  OAI21_X1 U9384 ( .B1(n7652), .B2(n7651), .A(n7650), .ZN(n7664) );
  INV_X1 U9385 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7662) );
  INV_X1 U9386 ( .A(n7892), .ZN(n7657) );
  NOR3_X1 U9387 ( .A1(n7655), .A2(n7654), .A3(n7653), .ZN(n7656) );
  OAI21_X1 U9388 ( .B1(n7657), .B2(n7656), .A(n10344), .ZN(n7661) );
  NOR2_X1 U9389 ( .A1(n7658), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8451) );
  AOI21_X1 U9390 ( .B1(n10317), .B2(n7659), .A(n8451), .ZN(n7660) );
  OAI211_X1 U9391 ( .C1(n7662), .C2(n7900), .A(n7661), .B(n7660), .ZN(n7663)
         );
  AOI21_X1 U9392 ( .B1(n7664), .B2(n10348), .A(n7663), .ZN(n7665) );
  INV_X1 U9393 ( .A(n7665), .ZN(P1_U3252) );
  INV_X1 U9394 ( .A(n9552), .ZN(n9594) );
  OAI21_X1 U9395 ( .B1(n7668), .B2(n7666), .A(n7836), .ZN(n9470) );
  INV_X1 U9396 ( .A(n9470), .ZN(n7672) );
  INV_X1 U9397 ( .A(n10457), .ZN(n7762) );
  AOI211_X1 U9398 ( .C1(n7762), .C2(n7668), .A(n9263), .B(n7667), .ZN(n7670)
         );
  OAI22_X1 U9399 ( .A1(n7924), .A2(n9419), .B1(n9418), .B2(n7774), .ZN(n7669)
         );
  NOR2_X1 U9400 ( .A1(n7670), .A2(n7669), .ZN(n9473) );
  AOI211_X1 U9401 ( .C1(n10489), .C2(n9468), .A(n10508), .B(n7846), .ZN(n9471)
         );
  AOI21_X1 U9402 ( .B1(n9588), .B2(n9468), .A(n9471), .ZN(n7671) );
  OAI211_X1 U9403 ( .C1(n9579), .C2(n7672), .A(n9473), .B(n7671), .ZN(n7677)
         );
  NAND2_X1 U9404 ( .A1(n7677), .A2(n10516), .ZN(n7673) );
  OAI21_X1 U9405 ( .B1(n10516), .B2(n6179), .A(n7673), .ZN(P2_U3454) );
  INV_X1 U9406 ( .A(n7674), .ZN(n7675) );
  NAND2_X1 U9407 ( .A1(n7677), .A2(n10526), .ZN(n7678) );
  OAI21_X1 U9408 ( .B1(n10526), .B2(n6130), .A(n7678), .ZN(P2_U3521) );
  INV_X1 U9409 ( .A(n7679), .ZN(n7681) );
  OAI222_X1 U9410 ( .A1(n9624), .A2(n7680), .B1(n8956), .B2(n7681), .C1(
        P2_U3152), .C2(n6073), .ZN(P2_U3343) );
  OAI222_X1 U9411 ( .A1(n10238), .A2(n7682), .B1(n4391), .B2(n7681), .C1(
        P1_U3084), .C2(n5173), .ZN(P1_U3338) );
  NOR2_X1 U9412 ( .A1(n7684), .A2(n7683), .ZN(n10291) );
  NOR2_X1 U9413 ( .A1(n7685), .A2(n7684), .ZN(n7687) );
  MUX2_X1 U9414 ( .A(n10291), .B(n7687), .S(n7686), .Z(n7691) );
  INV_X1 U9415 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7688) );
  NAND2_X1 U9416 ( .A1(n10288), .A2(n7688), .ZN(n7689) );
  AOI21_X1 U9417 ( .B1(n7690), .B2(n7689), .A(P1_IR_REG_0__SCAN_IN), .ZN(
        n10292) );
  OR3_X1 U9418 ( .A1(n7691), .A2(n10292), .A3(n9807), .ZN(n10312) );
  INV_X1 U9419 ( .A(n7692), .ZN(n7693) );
  OAI21_X1 U9420 ( .B1(n4489), .B2(n7694), .A(n7693), .ZN(n7699) );
  OAI21_X1 U9421 ( .B1(n7697), .B2(n7696), .A(n7695), .ZN(n7698) );
  AOI22_X1 U9422 ( .A1(n7699), .A2(n10348), .B1(n10344), .B2(n7698), .ZN(n7700) );
  NAND2_X1 U9423 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7823) );
  OAI211_X1 U9424 ( .C1(n10339), .C2(n7701), .A(n7700), .B(n7823), .ZN(n7702)
         );
  INV_X1 U9425 ( .A(n7702), .ZN(n7703) );
  OAI211_X1 U9426 ( .C1(n10245), .C2(n7900), .A(n10312), .B(n7703), .ZN(
        P1_U3245) );
  INV_X1 U9427 ( .A(n7704), .ZN(n7718) );
  AOI22_X1 U9428 ( .A1(n7705), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n10229), .ZN(n7706) );
  OAI21_X1 U9429 ( .B1(n7718), .B2(n4391), .A(n7706), .ZN(P1_U3337) );
  NAND2_X1 U9430 ( .A1(n9045), .A2(n7707), .ZN(n7708) );
  XOR2_X1 U9431 ( .A(n7709), .B(n7708), .Z(n7715) );
  NAND2_X1 U9432 ( .A1(n9444), .A2(n9122), .ZN(n7711) );
  NAND2_X1 U9433 ( .A1(n9446), .A2(n9123), .ZN(n7710) );
  NAND2_X1 U9434 ( .A1(n7711), .A2(n7710), .ZN(n7754) );
  AOI22_X1 U9435 ( .A1(n8615), .A2(n7754), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n7713) );
  NAND2_X1 U9436 ( .A1(n9102), .A2(n8194), .ZN(n7712) );
  OAI211_X1 U9437 ( .C1(n8196), .C2(n9023), .A(n7713), .B(n7712), .ZN(n7714)
         );
  AOI21_X1 U9438 ( .B1(n7715), .B2(n9048), .A(n7714), .ZN(n7716) );
  INV_X1 U9439 ( .A(n7716), .ZN(P2_U3229) );
  OAI222_X1 U9440 ( .A1(n8956), .A2(n7718), .B1(n9155), .B2(P2_U3152), .C1(
        n7717), .C2(n9624), .ZN(P2_U3342) );
  OR2_X1 U9441 ( .A1(n7719), .A2(n7723), .ZN(n7722) );
  NAND3_X1 U9442 ( .A1(n8250), .A2(n4495), .A3(n7941), .ZN(n7721) );
  NAND2_X1 U9443 ( .A1(n7723), .A2(n9990), .ZN(n8256) );
  OAI21_X1 U9444 ( .B1(n7726), .B2(n7724), .A(n7931), .ZN(n10370) );
  AOI21_X1 U9445 ( .B1(n10090), .B2(n8256), .A(n10370), .ZN(n7731) );
  XNOR2_X1 U9446 ( .A(n7726), .B(n7725), .ZN(n7727) );
  INV_X1 U9447 ( .A(n9808), .ZN(n8924) );
  OAI222_X1 U9448 ( .A1(n7727), .A2(n10044), .B1(n10040), .B2(n8925), .C1(
        n10071), .C2(n8924), .ZN(n10372) );
  OAI22_X1 U9449 ( .A1(n10049), .A2(n7729), .B1(n7728), .B2(n8934), .ZN(n7730)
         );
  NOR3_X1 U9450 ( .A1(n7731), .A2(n10372), .A3(n7730), .ZN(n7736) );
  NAND2_X1 U9451 ( .A1(n7153), .A2(n7982), .ZN(n7733) );
  NAND2_X1 U9452 ( .A1(n10429), .A2(n7733), .ZN(n7734) );
  NOR2_X1 U9453 ( .A1(n7732), .A2(n7734), .ZN(n10368) );
  AOI22_X1 U9454 ( .A1(n10024), .A2(n10368), .B1(P1_REG2_REG_1__SCAN_IN), .B2(
        n10020), .ZN(n7735) );
  OAI21_X1 U9455 ( .B1(n7736), .B2(n10020), .A(n7735), .ZN(P1_U3290) );
  XOR2_X1 U9456 ( .A(n7737), .B(n7738), .Z(n7739) );
  AOI22_X1 U9457 ( .A1(n9108), .A2(n8189), .B1(n9048), .B2(n7739), .ZN(n7744)
         );
  OAI22_X1 U9458 ( .A1(n6202), .A2(n9419), .B1(n9418), .B2(n7740), .ZN(n7843)
         );
  INV_X1 U9459 ( .A(n10472), .ZN(n7741) );
  NAND2_X1 U9460 ( .A1(n7742), .A2(n7741), .ZN(n7770) );
  AOI22_X1 U9461 ( .A1(n8615), .A2(n7843), .B1(n7770), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n7743) );
  NAND2_X1 U9462 ( .A1(n7744), .A2(n7743), .ZN(P2_U3239) );
  OAI21_X1 U9463 ( .B1(n7746), .B2(n6527), .A(n7745), .ZN(n8199) );
  AOI21_X1 U9464 ( .B1(n9438), .B2(n7747), .A(n10508), .ZN(n7749) );
  NAND2_X1 U9465 ( .A1(n7749), .A2(n7748), .ZN(n8202) );
  OAI21_X1 U9466 ( .B1(n8196), .B2(n10507), .A(n8202), .ZN(n7757) );
  NAND2_X1 U9467 ( .A1(n9442), .A2(n6528), .ZN(n9441) );
  NAND2_X1 U9468 ( .A1(n9441), .A2(n7750), .ZN(n7753) );
  NAND2_X1 U9469 ( .A1(n7753), .A2(n7752), .ZN(n7751) );
  OAI211_X1 U9470 ( .C1(n7753), .C2(n7752), .A(n7751), .B(n10460), .ZN(n7756)
         );
  INV_X1 U9471 ( .A(n7754), .ZN(n7755) );
  NAND2_X1 U9472 ( .A1(n7756), .A2(n7755), .ZN(n8198) );
  AOI211_X1 U9473 ( .C1(n10512), .C2(n8199), .A(n7757), .B(n8198), .ZN(n7864)
         );
  NAND2_X1 U9474 ( .A1(n10514), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n7758) );
  OAI21_X1 U9475 ( .B1(n7864), .B2(n10514), .A(n7758), .ZN(P2_U3466) );
  NAND2_X1 U9476 ( .A1(n9444), .A2(n9124), .ZN(n10458) );
  INV_X1 U9477 ( .A(n8615), .ZN(n9004) );
  AOI22_X1 U9478 ( .A1(n9108), .A2(n10489), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n7770), .ZN(n7764) );
  INV_X1 U9479 ( .A(n10456), .ZN(n7760) );
  MUX2_X1 U9480 ( .A(n7760), .B(n10489), .S(n7759), .Z(n7761) );
  OAI21_X1 U9481 ( .B1(n7762), .B2(n7761), .A(n9048), .ZN(n7763) );
  OAI211_X1 U9482 ( .C1(n10458), .C2(n9004), .A(n7764), .B(n7763), .ZN(
        P2_U3234) );
  AOI22_X1 U9483 ( .A1(n9468), .A2(n9108), .B1(n9092), .B2(n4389), .ZN(n7773)
         );
  AND2_X1 U9484 ( .A1(n7766), .A2(n7765), .ZN(n7769) );
  OAI21_X1 U9485 ( .B1(n7769), .B2(n7768), .A(n7767), .ZN(n7771) );
  AOI22_X1 U9486 ( .A1(n9048), .A2(n7771), .B1(n7770), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n7772) );
  OAI211_X1 U9487 ( .C1(n7774), .C2(n9072), .A(n7773), .B(n7772), .ZN(P2_U3224) );
  INV_X1 U9488 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7784) );
  OAI21_X1 U9489 ( .B1(n7776), .B2(n6525), .A(n7775), .ZN(n9461) );
  INV_X1 U9490 ( .A(n9461), .ZN(n7782) );
  XNOR2_X1 U9491 ( .A(n7778), .B(n7777), .ZN(n7779) );
  AOI222_X1 U9492 ( .A1(n4389), .A2(n9446), .B1(n9123), .B2(n9444), .C1(n10460), .C2(n7779), .ZN(n9458) );
  AOI21_X1 U9493 ( .B1(n9460), .B2(n7845), .A(n7780), .ZN(n9463) );
  AOI22_X1 U9494 ( .A1(n9463), .A2(n9589), .B1(n9588), .B2(n9460), .ZN(n7781)
         );
  OAI211_X1 U9495 ( .C1(n9579), .C2(n7782), .A(n9458), .B(n7781), .ZN(n7785)
         );
  NAND2_X1 U9496 ( .A1(n7785), .A2(n10516), .ZN(n7783) );
  OAI21_X1 U9497 ( .B1(n10516), .B2(n7784), .A(n7783), .ZN(P2_U3460) );
  NAND2_X1 U9498 ( .A1(n7785), .A2(n10526), .ZN(n7786) );
  OAI21_X1 U9499 ( .B1(n10526), .B2(n6133), .A(n7786), .ZN(P2_U3523) );
  OAI22_X1 U9500 ( .A1(n7097), .A2(n4401), .B1(n10388), .B2(n8012), .ZN(n7787)
         );
  XNOR2_X1 U9501 ( .A(n7787), .B(n8872), .ZN(n7999) );
  OAI22_X1 U9502 ( .A1(n7097), .A2(n8865), .B1(n10388), .B2(n4401), .ZN(n8000)
         );
  XNOR2_X1 U9503 ( .A(n7999), .B(n8000), .ZN(n7810) );
  XNOR2_X1 U9504 ( .A(n7788), .B(n8836), .ZN(n7799) );
  OAI22_X1 U9505 ( .A1(n8925), .A2(n8865), .B1(n8092), .B2(n4401), .ZN(n7800)
         );
  NAND2_X1 U9506 ( .A1(n7799), .A2(n7800), .ZN(n7869) );
  AND2_X1 U9507 ( .A1(n8869), .A2(n7153), .ZN(n7789) );
  INV_X1 U9508 ( .A(n7790), .ZN(n7791) );
  NAND2_X1 U9509 ( .A1(n7791), .A2(n8836), .ZN(n7793) );
  NAND2_X1 U9510 ( .A1(n9806), .A2(n8004), .ZN(n7795) );
  NAND2_X1 U9511 ( .A1(n8785), .A2(n7153), .ZN(n7794) );
  NAND2_X1 U9512 ( .A1(n7795), .A2(n7794), .ZN(n7796) );
  XNOR2_X1 U9513 ( .A(n7796), .B(n8836), .ZN(n7797) );
  INV_X1 U9514 ( .A(n7799), .ZN(n7802) );
  INV_X1 U9515 ( .A(n7800), .ZN(n7801) );
  NAND2_X1 U9516 ( .A1(n7802), .A2(n7801), .ZN(n7950) );
  OAI22_X1 U9517 ( .A1(n7094), .A2(n4401), .B1(n10380), .B2(n8012), .ZN(n7804)
         );
  XNOR2_X1 U9518 ( .A(n7804), .B(n8836), .ZN(n7806) );
  OAI22_X1 U9519 ( .A1(n7094), .A2(n8865), .B1(n10380), .B2(n4401), .ZN(n7805)
         );
  OR2_X1 U9520 ( .A1(n7806), .A2(n7805), .ZN(n7808) );
  NAND2_X1 U9521 ( .A1(n7806), .A2(n7805), .ZN(n7807) );
  AND2_X1 U9522 ( .A1(n7808), .A2(n7807), .ZN(n7951) );
  NAND2_X1 U9523 ( .A1(n7954), .A2(n7808), .ZN(n7809) );
  OAI21_X1 U9524 ( .B1(n7810), .B2(n7809), .A(n8003), .ZN(n7830) );
  AND3_X1 U9525 ( .A1(n7813), .A2(n7812), .A3(n7811), .ZN(n7815) );
  NAND2_X1 U9526 ( .A1(n7815), .A2(n7814), .ZN(n7816) );
  NAND2_X1 U9527 ( .A1(n7816), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7818) );
  INV_X1 U9528 ( .A(n8110), .ZN(n7828) );
  INV_X1 U9529 ( .A(n7819), .ZN(n7822) );
  INV_X1 U9530 ( .A(n7820), .ZN(n7821) );
  NAND2_X1 U9531 ( .A1(n9780), .A2(n9802), .ZN(n7824) );
  OAI211_X1 U9532 ( .C1(n9778), .C2(n7094), .A(n7824), .B(n7823), .ZN(n7825)
         );
  INV_X1 U9533 ( .A(n7825), .ZN(n7827) );
  NAND2_X1 U9534 ( .A1(n9784), .A2(n8109), .ZN(n7826) );
  OAI211_X1 U9535 ( .C1(n9782), .C2(n7828), .A(n7827), .B(n7826), .ZN(n7829)
         );
  AOI21_X1 U9536 ( .B1(n7830), .B2(n9772), .A(n7829), .ZN(n7831) );
  INV_X1 U9537 ( .A(n7831), .ZN(P1_U3228) );
  INV_X1 U9538 ( .A(n7832), .ZN(n7834) );
  OAI222_X1 U9539 ( .A1(n8956), .A2(n7834), .B1(n9177), .B2(P2_U3152), .C1(
        n7833), .C2(n9624), .ZN(P2_U3341) );
  OAI222_X1 U9540 ( .A1(n10238), .A2(n7835), .B1(n4391), .B2(n7834), .C1(
        n10338), .C2(P1_U3084), .ZN(P1_U3336) );
  INV_X1 U9541 ( .A(n7836), .ZN(n7838) );
  NOR2_X1 U9542 ( .A1(n7838), .A2(n7837), .ZN(n7840) );
  XNOR2_X1 U9543 ( .A(n7839), .B(n7840), .ZN(n8190) );
  XNOR2_X1 U9544 ( .A(n7841), .B(n7842), .ZN(n7844) );
  AOI21_X1 U9545 ( .B1(n7844), .B2(n10460), .A(n7843), .ZN(n8186) );
  OAI211_X1 U9546 ( .C1(n7846), .C2(n7847), .A(n9589), .B(n7845), .ZN(n8184)
         );
  OAI211_X1 U9547 ( .C1(n7847), .C2(n10507), .A(n8186), .B(n8184), .ZN(n7848)
         );
  AOI21_X1 U9548 ( .B1(n10512), .B2(n8190), .A(n7848), .ZN(n7850) );
  OR2_X1 U9549 ( .A1(n10514), .A2(n7850), .ZN(n7849) );
  OAI21_X1 U9550 ( .B1(n10516), .B2(n6170), .A(n7849), .ZN(P2_U3457) );
  OR2_X1 U9551 ( .A1(n10523), .A2(n7850), .ZN(n7851) );
  OAI21_X1 U9552 ( .B1(n10526), .B2(n7852), .A(n7851), .ZN(P2_U3522) );
  XOR2_X1 U9553 ( .A(n7853), .B(n4488), .Z(n7862) );
  NOR2_X1 U9554 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7987), .ZN(n7854) );
  AOI21_X1 U9555 ( .B1(n9174), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n7854), .ZN(
        n7855) );
  OAI21_X1 U9556 ( .B1(n9178), .B2(n7856), .A(n7855), .ZN(n7861) );
  AOI211_X1 U9557 ( .C1(n7859), .C2(n7858), .A(n9184), .B(n7857), .ZN(n7860)
         );
  AOI211_X1 U9558 ( .C1(n9169), .C2(n7862), .A(n7861), .B(n7860), .ZN(n7863)
         );
  INV_X1 U9559 ( .A(n7863), .ZN(P2_U3253) );
  OR2_X1 U9560 ( .A1(n7864), .A2(n10523), .ZN(n7865) );
  OAI21_X1 U9561 ( .B1(n10526), .B2(n7866), .A(n7865), .ZN(P2_U3525) );
  INV_X1 U9562 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7877) );
  NOR2_X1 U9563 ( .A1(n7867), .A2(n7868), .ZN(n8929) );
  NAND2_X1 U9564 ( .A1(n8929), .A2(n8930), .ZN(n8928) );
  INV_X1 U9565 ( .A(n7868), .ZN(n7871) );
  NAND2_X1 U9566 ( .A1(n7869), .A2(n7950), .ZN(n7870) );
  AOI21_X1 U9567 ( .B1(n8928), .B2(n7871), .A(n7870), .ZN(n7953) );
  AND3_X1 U9568 ( .A1(n8928), .A2(n7871), .A3(n7870), .ZN(n7872) );
  OAI21_X1 U9569 ( .B1(n7953), .B2(n7872), .A(n9772), .ZN(n7876) );
  INV_X1 U9570 ( .A(n8347), .ZN(n8031) );
  NAND2_X1 U9571 ( .A1(n7873), .A2(n10428), .ZN(n10374) );
  OAI22_X1 U9572 ( .A1(n8031), .A2(n10374), .B1(n9778), .B2(n8087), .ZN(n7874)
         );
  AOI21_X1 U9573 ( .B1(n9780), .B2(n9804), .A(n7874), .ZN(n7875) );
  OAI211_X1 U9574 ( .C1(n7878), .C2(n7877), .A(n7876), .B(n7875), .ZN(P1_U3235) );
  INV_X1 U9575 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7880) );
  INV_X1 U9576 ( .A(n7879), .ZN(n7881) );
  OAI222_X1 U9577 ( .A1(n9624), .A2(n7880), .B1(n9627), .B2(n7881), .C1(
        P2_U3152), .C2(n6082), .ZN(P2_U3340) );
  INV_X1 U9578 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7882) );
  OAI222_X1 U9579 ( .A1(n10238), .A2(n7882), .B1(n4391), .B2(n7881), .C1(
        P1_U3084), .C2(n9827), .ZN(P1_U3335) );
  INV_X1 U9580 ( .A(n7883), .ZN(n7885) );
  OAI222_X1 U9581 ( .A1(n10238), .A2(n7884), .B1(n4391), .B2(n7885), .C1(
        P1_U3084), .C2(n8059), .ZN(P1_U3334) );
  OAI222_X1 U9582 ( .A1(n9624), .A2(n7886), .B1(n9627), .B2(n7885), .C1(
        P2_U3152), .C2(n4944), .ZN(P2_U3339) );
  AOI211_X1 U9583 ( .C1(n7889), .C2(n7888), .A(n10305), .B(n7887), .ZN(n7902)
         );
  INV_X1 U9584 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7899) );
  AND3_X1 U9585 ( .A1(n7892), .A2(n7891), .A3(n7890), .ZN(n7893) );
  OAI21_X1 U9586 ( .B1(n7894), .B2(n7893), .A(n10344), .ZN(n7898) );
  NOR2_X1 U9587 ( .A1(n7895), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8471) );
  AOI21_X1 U9588 ( .B1(n10317), .B2(n7896), .A(n8471), .ZN(n7897) );
  OAI211_X1 U9589 ( .C1(n7900), .C2(n7899), .A(n7898), .B(n7897), .ZN(n7901)
         );
  OR2_X1 U9590 ( .A1(n7902), .A2(n7901), .ZN(P1_U3253) );
  XNOR2_X1 U9591 ( .A(n7904), .B(n7903), .ZN(n7909) );
  AOI22_X1 U9592 ( .A1(n9092), .A2(n9120), .B1(n9103), .B2(n9122), .ZN(n7908)
         );
  NOR2_X1 U9593 ( .A1(n9023), .A2(n4845), .ZN(n7905) );
  AOI211_X1 U9594 ( .C1(n9102), .C2(n8128), .A(n7906), .B(n7905), .ZN(n7907)
         );
  OAI211_X1 U9595 ( .C1(n7909), .C2(n9110), .A(n7908), .B(n7907), .ZN(P2_U3215) );
  INV_X1 U9596 ( .A(n7910), .ZN(n7911) );
  AOI21_X1 U9597 ( .B1(n7913), .B2(n7912), .A(n7911), .ZN(n7919) );
  OAI21_X1 U9598 ( .B1(n9023), .B2(n4847), .A(n7914), .ZN(n7917) );
  OAI22_X1 U9599 ( .A1(n7988), .A2(n9106), .B1(n9072), .B2(n7915), .ZN(n7916)
         );
  AOI211_X1 U9600 ( .C1(n8177), .C2(n9102), .A(n7917), .B(n7916), .ZN(n7918)
         );
  OAI21_X1 U9601 ( .B1(n7919), .B2(n9110), .A(n7918), .ZN(P2_U3241) );
  XNOR2_X1 U9602 ( .A(n4394), .B(n7920), .ZN(n7928) );
  OAI22_X1 U9603 ( .A1(n9023), .A2(n7922), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9462), .ZN(n7926) );
  OAI22_X1 U9604 ( .A1(n7924), .A2(n9072), .B1(n9106), .B2(n7923), .ZN(n7925)
         );
  AOI211_X1 U9605 ( .C1(n9102), .C2(n9462), .A(n7926), .B(n7925), .ZN(n7927)
         );
  OAI21_X1 U9606 ( .B1(n9110), .B2(n7928), .A(n7927), .ZN(P2_U3220) );
  INV_X1 U9607 ( .A(n7929), .ZN(n7930) );
  NAND2_X1 U9608 ( .A1(n7931), .A2(n7930), .ZN(n8089) );
  NOR2_X1 U9609 ( .A1(n8089), .A2(n8090), .ZN(n8088) );
  NAND2_X1 U9610 ( .A1(n7933), .A2(n7932), .ZN(n7935) );
  OAI21_X1 U9611 ( .B1(n8088), .B2(n7935), .A(n7934), .ZN(n10384) );
  INV_X1 U9612 ( .A(n10384), .ZN(n7949) );
  INV_X1 U9613 ( .A(n5917), .ZN(n7939) );
  INV_X1 U9614 ( .A(n7936), .ZN(n7937) );
  AOI21_X1 U9615 ( .B1(n7939), .B2(n7938), .A(n7937), .ZN(n7940) );
  OAI222_X1 U9616 ( .A1(n10040), .A2(n7097), .B1(n10071), .B2(n8925), .C1(
        n7940), .C2(n10044), .ZN(n10382) );
  NAND2_X1 U9617 ( .A1(n10382), .A2(n10078), .ZN(n7948) );
  INV_X1 U9618 ( .A(n7941), .ZN(n7942) );
  OR2_X1 U9619 ( .A1(n7971), .A2(n7942), .ZN(n7943) );
  OAI21_X1 U9620 ( .B1(n7154), .B2(n10380), .A(n8107), .ZN(n10381) );
  NOR2_X1 U9621 ( .A1(n10063), .A2(n10381), .ZN(n7946) );
  OAI22_X1 U9622 ( .A1(n10078), .A2(n7944), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10049), .ZN(n7945) );
  AOI211_X1 U9623 ( .C1(n10060), .C2(n7959), .A(n7946), .B(n7945), .ZN(n7947)
         );
  OAI211_X1 U9624 ( .C1(n10009), .C2(n7949), .A(n7948), .B(n7947), .ZN(
        P1_U3288) );
  INV_X1 U9625 ( .A(n7950), .ZN(n7952) );
  NOR3_X1 U9626 ( .A1(n7953), .A2(n7952), .A3(n7951), .ZN(n7956) );
  INV_X1 U9627 ( .A(n7954), .ZN(n7955) );
  OAI21_X1 U9628 ( .B1(n7956), .B2(n7955), .A(n9772), .ZN(n7961) );
  NAND2_X1 U9629 ( .A1(n9780), .A2(n9803), .ZN(n7957) );
  NAND2_X1 U9630 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n10273) );
  OAI211_X1 U9631 ( .C1(n9778), .C2(n8925), .A(n7957), .B(n10273), .ZN(n7958)
         );
  AOI21_X1 U9632 ( .B1(n9784), .B2(n7959), .A(n7958), .ZN(n7960) );
  OAI211_X1 U9633 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9782), .A(n7961), .B(
        n7960), .ZN(P1_U3216) );
  NAND2_X1 U9634 ( .A1(n10184), .A2(n5946), .ZN(n7962) );
  NAND2_X1 U9635 ( .A1(n7963), .A2(n7962), .ZN(n7965) );
  NOR2_X4 U9636 ( .A1(n7976), .A2(n10226), .ZN(n10437) );
  INV_X1 U9637 ( .A(n7971), .ZN(n7968) );
  INV_X1 U9638 ( .A(n7966), .ZN(n7967) );
  NOR3_X1 U9639 ( .A1(n7969), .A2(n7968), .A3(n7967), .ZN(n7970) );
  AOI21_X1 U9640 ( .B1(n10068), .B2(n9806), .A(n7970), .ZN(n7985) );
  OAI21_X1 U9641 ( .B1(n7972), .B2(n7971), .A(n7985), .ZN(n7977) );
  NAND2_X1 U9642 ( .A1(n7977), .A2(n10437), .ZN(n7973) );
  OAI21_X1 U9643 ( .B1(n10437), .B2(n7974), .A(n7973), .ZN(P1_U3454) );
  NOR2_X4 U9644 ( .A1(n7976), .A2(n7975), .ZN(n10455) );
  NAND2_X1 U9645 ( .A1(n7977), .A2(n10455), .ZN(n7978) );
  OAI21_X1 U9646 ( .B1(n10455), .B2(n5124), .A(n7978), .ZN(P1_U3523) );
  INV_X1 U9647 ( .A(n7979), .ZN(n7994) );
  OAI222_X1 U9648 ( .A1(n8956), .A2(n7994), .B1(n7981), .B2(P2_U3152), .C1(
        n7980), .C2(n9624), .ZN(P2_U3338) );
  AOI22_X1 U9649 ( .A1(n10020), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n10059), .ZN(n7984) );
  OAI21_X1 U9650 ( .B1(n10007), .B2(n10060), .A(n7982), .ZN(n7983) );
  OAI211_X1 U9651 ( .C1(n7985), .C2(n10020), .A(n7984), .B(n7983), .ZN(
        P1_U3291) );
  XNOR2_X1 U9652 ( .A(n7986), .B(n8145), .ZN(n7992) );
  OAI22_X1 U9653 ( .A1(n9023), .A2(n8364), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7987), .ZN(n7990) );
  OAI22_X1 U9654 ( .A1(n7988), .A2(n9072), .B1(n9106), .B2(n8209), .ZN(n7989)
         );
  AOI211_X1 U9655 ( .C1(n8307), .C2(n9102), .A(n7990), .B(n7989), .ZN(n7991)
         );
  OAI21_X1 U9656 ( .B1(n7992), .B2(n9110), .A(n7991), .ZN(P2_U3223) );
  OAI222_X1 U9657 ( .A1(n10238), .A2(n7995), .B1(n4391), .B2(n7994), .C1(n7993), .C2(P1_U3084), .ZN(P1_U3333) );
  INV_X1 U9658 ( .A(n7996), .ZN(n8957) );
  OAI222_X1 U9659 ( .A1(n8956), .A2(n8957), .B1(n7998), .B2(P2_U3152), .C1(
        n7997), .C2(n9624), .ZN(P2_U3337) );
  INV_X1 U9660 ( .A(n7999), .ZN(n8001) );
  OR2_X1 U9661 ( .A1(n8001), .A2(n8000), .ZN(n8002) );
  NAND2_X1 U9662 ( .A1(n9802), .A2(n8869), .ZN(n8006) );
  NAND2_X1 U9663 ( .A1(n8246), .A2(n8785), .ZN(n8005) );
  NAND2_X1 U9664 ( .A1(n8006), .A2(n8005), .ZN(n8007) );
  XNOR2_X1 U9665 ( .A(n8007), .B(n8836), .ZN(n8238) );
  INV_X1 U9666 ( .A(n8238), .ZN(n8010) );
  NAND2_X1 U9667 ( .A1(n9802), .A2(n8874), .ZN(n8009) );
  NAND2_X1 U9668 ( .A1(n8246), .A2(n8869), .ZN(n8008) );
  NAND2_X1 U9669 ( .A1(n8009), .A2(n8008), .ZN(n8016) );
  INV_X1 U9670 ( .A(n8016), .ZN(n8241) );
  AND2_X1 U9671 ( .A1(n8010), .A2(n8241), .ZN(n8019) );
  OAI22_X1 U9672 ( .A1(n8346), .A2(n8012), .B1(n8011), .B2(n4401), .ZN(n8013)
         );
  XNOR2_X1 U9673 ( .A(n8013), .B(n8836), .ZN(n8020) );
  OR2_X1 U9674 ( .A1(n8346), .A2(n4401), .ZN(n8015) );
  NAND2_X1 U9675 ( .A1(n9801), .A2(n8874), .ZN(n8014) );
  NAND2_X1 U9676 ( .A1(n8015), .A2(n8014), .ZN(n8021) );
  NAND2_X1 U9677 ( .A1(n8020), .A2(n8021), .ZN(n8339) );
  NAND2_X1 U9678 ( .A1(n8238), .A2(n8016), .ZN(n8017) );
  AND2_X1 U9679 ( .A1(n8339), .A2(n8017), .ZN(n8018) );
  INV_X1 U9680 ( .A(n8020), .ZN(n8023) );
  INV_X1 U9681 ( .A(n8021), .ZN(n8022) );
  NAND2_X1 U9682 ( .A1(n8023), .A2(n8022), .ZN(n8338) );
  NAND2_X1 U9683 ( .A1(n8080), .A2(n8869), .ZN(n8026) );
  OR2_X1 U9684 ( .A1(n8286), .A2(n8865), .ZN(n8025) );
  AND2_X1 U9685 ( .A1(n8026), .A2(n8025), .ZN(n8277) );
  NAND2_X1 U9686 ( .A1(n8080), .A2(n8785), .ZN(n8028) );
  OR2_X1 U9687 ( .A1(n8286), .A2(n4401), .ZN(n8027) );
  NAND2_X1 U9688 ( .A1(n8028), .A2(n8027), .ZN(n8029) );
  XNOR2_X1 U9689 ( .A(n8029), .B(n8836), .ZN(n8276) );
  XOR2_X1 U9690 ( .A(n8277), .B(n8276), .Z(n8030) );
  XNOR2_X1 U9691 ( .A(n8278), .B(n8030), .ZN(n8037) );
  NAND2_X1 U9692 ( .A1(n8080), .A2(n10428), .ZN(n10421) );
  NOR2_X1 U9693 ( .A1(n8031), .A2(n10421), .ZN(n8035) );
  INV_X1 U9694 ( .A(n9778), .ZN(n9735) );
  AOI21_X1 U9695 ( .B1(n9735), .B2(n9801), .A(n8032), .ZN(n8033) );
  OAI21_X1 U9696 ( .B1(n8386), .B2(n9683), .A(n8033), .ZN(n8034) );
  AOI211_X1 U9697 ( .C1(n8079), .C2(n9713), .A(n8035), .B(n8034), .ZN(n8036)
         );
  OAI21_X1 U9698 ( .B1(n8037), .B2(n9760), .A(n8036), .ZN(P1_U3211) );
  XOR2_X1 U9699 ( .A(n8039), .B(n8038), .Z(n8048) );
  NAND2_X1 U9700 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n8152) );
  INV_X1 U9701 ( .A(n8152), .ZN(n8040) );
  AOI21_X1 U9702 ( .B1(n9174), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8040), .ZN(
        n8041) );
  OAI21_X1 U9703 ( .B1(n9178), .B2(n8042), .A(n8041), .ZN(n8047) );
  AOI211_X1 U9704 ( .C1(n8045), .C2(n8044), .A(n9184), .B(n8043), .ZN(n8046)
         );
  AOI211_X1 U9705 ( .C1(n9169), .C2(n8048), .A(n8047), .B(n8046), .ZN(n8049)
         );
  INV_X1 U9706 ( .A(n8049), .ZN(P2_U3254) );
  OAI21_X1 U9707 ( .B1(n5015), .B2(n10401), .A(n10429), .ZN(n8050) );
  NOR2_X1 U9708 ( .A1(n8050), .A2(n8257), .ZN(n10403) );
  INV_X1 U9709 ( .A(n8051), .ZN(n8249) );
  NAND2_X1 U9710 ( .A1(n9801), .A2(n10068), .ZN(n10399) );
  OAI21_X1 U9711 ( .B1(n10049), .B2(n8249), .A(n10399), .ZN(n8058) );
  NAND2_X1 U9712 ( .A1(n8053), .A2(n8052), .ZN(n8054) );
  NAND2_X1 U9713 ( .A1(n8054), .A2(n8061), .ZN(n8263) );
  OAI21_X1 U9714 ( .B1(n8061), .B2(n8054), .A(n8263), .ZN(n8055) );
  NAND2_X1 U9715 ( .A1(n8055), .A2(n10074), .ZN(n8057) );
  OR2_X1 U9716 ( .A1(n7097), .A2(n10071), .ZN(n8056) );
  NAND2_X1 U9717 ( .A1(n8057), .A2(n8056), .ZN(n10407) );
  AOI211_X1 U9718 ( .C1(n10403), .C2(n8059), .A(n8058), .B(n10407), .ZN(n8066)
         );
  OR2_X1 U9719 ( .A1(n8060), .A2(n8061), .ZN(n8253) );
  NAND2_X1 U9720 ( .A1(n8060), .A2(n8061), .ZN(n8062) );
  AND2_X1 U9721 ( .A1(n8253), .A2(n8062), .ZN(n10398) );
  INV_X1 U9722 ( .A(n10009), .ZN(n10030) );
  OAI22_X1 U9723 ( .A1(n10078), .A2(n8063), .B1(n9999), .B2(n10401), .ZN(n8064) );
  AOI21_X1 U9724 ( .B1(n10398), .B2(n10030), .A(n8064), .ZN(n8065) );
  OAI21_X1 U9725 ( .B1(n8066), .B2(n10020), .A(n8065), .ZN(P1_U3286) );
  NAND3_X1 U9726 ( .A1(n8068), .A2(n8076), .A3(n8067), .ZN(n8069) );
  NAND2_X1 U9727 ( .A1(n8318), .A2(n8069), .ZN(n8070) );
  NAND2_X1 U9728 ( .A1(n8070), .A2(n10074), .ZN(n8072) );
  AOI22_X1 U9729 ( .A1(n9799), .A2(n10068), .B1(n10011), .B2(n9801), .ZN(n8071) );
  NAND2_X1 U9730 ( .A1(n8072), .A2(n8071), .ZN(n10425) );
  INV_X1 U9731 ( .A(n10425), .ZN(n8085) );
  INV_X1 U9732 ( .A(n8073), .ZN(n8074) );
  NAND2_X1 U9733 ( .A1(n8075), .A2(n8074), .ZN(n8077) );
  XNOR2_X1 U9734 ( .A(n8077), .B(n8076), .ZN(n10420) );
  AOI21_X1 U9735 ( .B1(n8259), .B2(n8080), .A(n10413), .ZN(n8078) );
  NAND2_X1 U9736 ( .A1(n8078), .A2(n8323), .ZN(n10422) );
  AOI22_X1 U9737 ( .A1(n10020), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n8079), .B2(
        n10059), .ZN(n8082) );
  NAND2_X1 U9738 ( .A1(n10060), .A2(n8080), .ZN(n8081) );
  OAI211_X1 U9739 ( .C1(n10422), .C2(n8643), .A(n8082), .B(n8081), .ZN(n8083)
         );
  AOI21_X1 U9740 ( .B1(n10420), .B2(n10030), .A(n8083), .ZN(n8084) );
  OAI21_X1 U9741 ( .B1(n8085), .B2(n10020), .A(n8084), .ZN(P1_U3284) );
  XOR2_X1 U9742 ( .A(n5962), .B(n8090), .Z(n8086) );
  OAI222_X1 U9743 ( .A1(n10040), .A2(n7094), .B1(n10071), .B2(n8087), .C1(
        n8086), .C2(n10044), .ZN(n10376) );
  INV_X1 U9744 ( .A(n10376), .ZN(n8099) );
  AOI21_X1 U9745 ( .B1(n8090), .B2(n8089), .A(n8088), .ZN(n8091) );
  INV_X1 U9746 ( .A(n8091), .ZN(n10378) );
  NOR2_X1 U9747 ( .A1(n9999), .A2(n8092), .ZN(n8097) );
  OR2_X1 U9748 ( .A1(n7732), .A2(n8092), .ZN(n8093) );
  NOR2_X1 U9749 ( .A1(n10049), .A2(n7877), .ZN(n8094) );
  AOI21_X1 U9750 ( .B1(n10020), .B2(P1_REG2_REG_2__SCAN_IN), .A(n8094), .ZN(
        n8095) );
  OAI21_X1 U9751 ( .B1(n10063), .B2(n10375), .A(n8095), .ZN(n8096) );
  AOI211_X1 U9752 ( .C1(n10378), .C2(n10030), .A(n8097), .B(n8096), .ZN(n8098)
         );
  OAI21_X1 U9753 ( .B1(n8099), .B2(n10020), .A(n8098), .ZN(P1_U3289) );
  INV_X1 U9754 ( .A(n8106), .ZN(n8100) );
  XNOR2_X1 U9755 ( .A(n8101), .B(n8100), .ZN(n8104) );
  NAND2_X1 U9756 ( .A1(n9802), .A2(n10068), .ZN(n8102) );
  OAI21_X1 U9757 ( .B1(n7094), .B2(n10071), .A(n8102), .ZN(n8103) );
  AOI21_X1 U9758 ( .B1(n8104), .B2(n10074), .A(n8103), .ZN(n10395) );
  XNOR2_X1 U9759 ( .A(n8106), .B(n8105), .ZN(n10387) );
  AND2_X1 U9760 ( .A1(n8107), .A2(n8109), .ZN(n8108) );
  OR2_X1 U9761 ( .A1(n8108), .A2(n5015), .ZN(n10389) );
  NAND2_X1 U9762 ( .A1(n10060), .A2(n8109), .ZN(n8112) );
  AOI22_X1 U9763 ( .A1(n10020), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n8110), .B2(
        n10059), .ZN(n8111) );
  OAI211_X1 U9764 ( .C1(n10389), .C2(n10063), .A(n8112), .B(n8111), .ZN(n8113)
         );
  AOI21_X1 U9765 ( .B1(n10387), .B2(n10030), .A(n8113), .ZN(n8114) );
  OAI21_X1 U9766 ( .B1(n10395), .B2(n10020), .A(n8114), .ZN(P1_U3287) );
  NAND2_X1 U9767 ( .A1(n7745), .A2(n8115), .ZN(n8171) );
  NAND2_X1 U9768 ( .A1(n8171), .A2(n8116), .ZN(n8118) );
  NAND2_X1 U9769 ( .A1(n8118), .A2(n8117), .ZN(n8119) );
  XNOR2_X1 U9770 ( .A(n8119), .B(n8121), .ZN(n10513) );
  INV_X1 U9771 ( .A(n10513), .ZN(n8133) );
  NOR2_X1 U9772 ( .A1(n8120), .A2(n8121), .ZN(n8297) );
  NAND2_X1 U9773 ( .A1(n8120), .A2(n8121), .ZN(n8122) );
  NAND2_X1 U9774 ( .A1(n8122), .A2(n9385), .ZN(n8123) );
  OR2_X1 U9775 ( .A1(n8297), .A2(n8123), .ZN(n8125) );
  AOI22_X1 U9776 ( .A1(n9446), .A2(n9122), .B1(n9444), .B2(n9120), .ZN(n8124)
         );
  NAND2_X1 U9777 ( .A1(n8125), .A2(n8124), .ZN(n10510) );
  NOR2_X2 U9778 ( .A1(n8185), .A2(n10508), .ZN(n9464) );
  XNOR2_X1 U9779 ( .A(n8176), .B(n8126), .ZN(n10509) );
  INV_X1 U9780 ( .A(n10509), .ZN(n8127) );
  NAND2_X1 U9781 ( .A1(n9464), .A2(n8127), .ZN(n8130) );
  AOI22_X1 U9782 ( .A1(n10461), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n8128), .B2(
        n10462), .ZN(n8129) );
  OAI211_X1 U9783 ( .C1(n4845), .C2(n10464), .A(n8130), .B(n8129), .ZN(n8131)
         );
  AOI21_X1 U9784 ( .B1(n10510), .B2(n9457), .A(n8131), .ZN(n8132) );
  OAI21_X1 U9785 ( .B1(n9411), .B2(n8133), .A(n8132), .ZN(P2_U3289) );
  AOI21_X1 U9786 ( .B1(n4483), .B2(n8135), .A(n8134), .ZN(n8144) );
  XOR2_X1 U9787 ( .A(n8137), .B(n8136), .Z(n8138) );
  NAND2_X1 U9788 ( .A1(n8138), .A2(n10348), .ZN(n8143) );
  NOR2_X1 U9789 ( .A1(n8139), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8602) );
  NOR2_X1 U9790 ( .A1(n10339), .A2(n8140), .ZN(n8141) );
  AOI211_X1 U9791 ( .C1(n10342), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n8602), .B(
        n8141), .ZN(n8142) );
  OAI211_X1 U9792 ( .C1(n8144), .C2(n10300), .A(n8143), .B(n8142), .ZN(
        P1_U3254) );
  NAND2_X1 U9793 ( .A1(n7986), .A2(n8145), .ZN(n8148) );
  NAND2_X1 U9794 ( .A1(n8148), .A2(n8146), .ZN(n8151) );
  NAND2_X1 U9795 ( .A1(n8148), .A2(n8147), .ZN(n8158) );
  INV_X1 U9796 ( .A(n8158), .ZN(n8149) );
  AOI21_X1 U9797 ( .B1(n8151), .B2(n8150), .A(n8149), .ZN(n8156) );
  INV_X1 U9798 ( .A(n9587), .ZN(n8554) );
  OAI21_X1 U9799 ( .B1(n9023), .B2(n8554), .A(n8152), .ZN(n8154) );
  OAI22_X1 U9800 ( .A1(n8545), .A2(n9072), .B1(n9106), .B2(n8546), .ZN(n8153)
         );
  AOI211_X1 U9801 ( .C1(n8552), .C2(n9102), .A(n8154), .B(n8153), .ZN(n8155)
         );
  OAI21_X1 U9802 ( .B1(n8156), .B2(n9110), .A(n8155), .ZN(P2_U3233) );
  NAND2_X1 U9803 ( .A1(n8158), .A2(n8157), .ZN(n8160) );
  XNOR2_X1 U9804 ( .A(n8159), .B(n8160), .ZN(n8164) );
  OAI22_X1 U9805 ( .A1(n9023), .A2(n4543), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8353), .ZN(n8162) );
  OAI22_X1 U9806 ( .A1(n8209), .A2(n9072), .B1(n9106), .B2(n8655), .ZN(n8161)
         );
  AOI211_X1 U9807 ( .C1(n8214), .C2(n9102), .A(n8162), .B(n8161), .ZN(n8163)
         );
  OAI21_X1 U9808 ( .B1(n8164), .B2(n9110), .A(n8163), .ZN(P2_U3219) );
  XNOR2_X1 U9809 ( .A(n8165), .B(n8166), .ZN(n8170) );
  OAI22_X1 U9810 ( .A1(n9072), .A2(n8546), .B1(n8233), .B2(n9023), .ZN(n8168)
         );
  OAI22_X1 U9811 ( .A1(n9106), .A2(n9417), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6296), .ZN(n8167) );
  AOI211_X1 U9812 ( .C1(n8231), .C2(n9102), .A(n8168), .B(n8167), .ZN(n8169)
         );
  OAI21_X1 U9813 ( .B1(n8170), .B2(n9110), .A(n8169), .ZN(P2_U3238) );
  XNOR2_X1 U9814 ( .A(n8171), .B(n4422), .ZN(n10500) );
  AOI222_X1 U9815 ( .A1(n10460), .A2(n8173), .B1(n9121), .B2(n9444), .C1(n9443), .C2(n9446), .ZN(n10502) );
  MUX2_X1 U9816 ( .A(n8174), .B(n10502), .S(n9457), .Z(n8182) );
  INV_X1 U9817 ( .A(n9464), .ZN(n10465) );
  NAND2_X1 U9818 ( .A1(n7748), .A2(n8180), .ZN(n8175) );
  NAND2_X1 U9819 ( .A1(n8176), .A2(n8175), .ZN(n10501) );
  INV_X1 U9820 ( .A(n8177), .ZN(n8178) );
  OAI22_X1 U9821 ( .A1(n10465), .A2(n10501), .B1(n8178), .B2(n9290), .ZN(n8179) );
  AOI21_X1 U9822 ( .B1(n9469), .B2(n8180), .A(n8179), .ZN(n8181) );
  OAI211_X1 U9823 ( .C1(n9411), .C2(n10500), .A(n8182), .B(n8181), .ZN(
        P2_U3290) );
  INV_X1 U9824 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n8183) );
  OAI22_X1 U9825 ( .A1(n8185), .A2(n8184), .B1(n8183), .B2(n9290), .ZN(n8188)
         );
  NOR2_X1 U9826 ( .A1(n10461), .A2(n8186), .ZN(n8187) );
  AOI211_X1 U9827 ( .C1(n10461), .C2(P2_REG2_REG_2__SCAN_IN), .A(n8188), .B(
        n8187), .ZN(n8192) );
  AOI22_X1 U9828 ( .A1(n10467), .A2(n8190), .B1(n9469), .B2(n8189), .ZN(n8191)
         );
  NAND2_X1 U9829 ( .A1(n8192), .A2(n8191), .ZN(P2_U3294) );
  OR2_X1 U9830 ( .A1(n10461), .A2(n8193), .ZN(n9334) );
  AOI22_X1 U9831 ( .A1(n10461), .A2(P2_REG2_REG_5__SCAN_IN), .B1(n8194), .B2(
        n10462), .ZN(n8195) );
  OAI21_X1 U9832 ( .B1(n10464), .B2(n8196), .A(n8195), .ZN(n8197) );
  AOI21_X1 U9833 ( .B1(n9457), .B2(n8198), .A(n8197), .ZN(n8201) );
  NAND2_X1 U9834 ( .A1(n10467), .A2(n8199), .ZN(n8200) );
  OAI211_X1 U9835 ( .C1(n8202), .C2(n9334), .A(n8201), .B(n8200), .ZN(P2_U3291) );
  INV_X1 U9836 ( .A(n8203), .ZN(n8205) );
  AOI21_X1 U9837 ( .B1(n8120), .B2(n8205), .A(n8204), .ZN(n8207) );
  NOR3_X1 U9838 ( .A1(n8207), .A2(n8206), .A3(n8218), .ZN(n8208) );
  NOR2_X1 U9839 ( .A1(n8208), .A2(n9263), .ZN(n8212) );
  OAI22_X1 U9840 ( .A1(n8655), .A2(n9419), .B1(n9418), .B2(n8209), .ZN(n8210)
         );
  AOI21_X1 U9841 ( .B1(n8212), .B2(n8211), .A(n8210), .ZN(n9586) );
  AOI21_X1 U9842 ( .B1(n9580), .B2(n8213), .A(n8229), .ZN(n9581) );
  AOI22_X1 U9843 ( .A1(n10461), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n8214), .B2(
        n10462), .ZN(n8215) );
  OAI21_X1 U9844 ( .B1(n10464), .B2(n4543), .A(n8215), .ZN(n8216) );
  AOI21_X1 U9845 ( .B1(n9581), .B2(n9464), .A(n8216), .ZN(n8223) );
  INV_X1 U9846 ( .A(n8291), .ZN(n8294) );
  OAI21_X1 U9847 ( .B1(n8294), .B2(n8217), .A(n4476), .ZN(n8219) );
  NAND2_X1 U9848 ( .A1(n8219), .A2(n8218), .ZN(n9583) );
  INV_X1 U9849 ( .A(n8219), .ZN(n8221) );
  NAND2_X1 U9850 ( .A1(n8221), .A2(n8220), .ZN(n9582) );
  NAND3_X1 U9851 ( .A1(n9583), .A2(n10467), .A3(n9582), .ZN(n8222) );
  OAI211_X1 U9852 ( .C1(n9586), .C2(n10461), .A(n8223), .B(n8222), .ZN(
        P2_U3286) );
  OAI21_X1 U9853 ( .B1(n8225), .B2(n8227), .A(n8224), .ZN(n9578) );
  XNOR2_X1 U9854 ( .A(n8226), .B(n8227), .ZN(n8228) );
  AOI222_X1 U9855 ( .A1(n9385), .A2(n8228), .B1(n9116), .B2(n9444), .C1(n9118), 
        .C2(n9446), .ZN(n9577) );
  MUX2_X1 U9856 ( .A(n6059), .B(n9577), .S(n9457), .Z(n8236) );
  INV_X1 U9857 ( .A(n8229), .ZN(n8230) );
  AOI21_X1 U9858 ( .B1(n9574), .B2(n8230), .A(n6572), .ZN(n9575) );
  INV_X1 U9859 ( .A(n8231), .ZN(n8232) );
  OAI22_X1 U9860 ( .A1(n10464), .A2(n8233), .B1(n9290), .B2(n8232), .ZN(n8234)
         );
  AOI21_X1 U9861 ( .B1(n9575), .B2(n9464), .A(n8234), .ZN(n8235) );
  OAI211_X1 U9862 ( .C1(n9411), .C2(n9578), .A(n8236), .B(n8235), .ZN(P2_U3285) );
  INV_X1 U9863 ( .A(n8237), .ZN(n8239) );
  NOR2_X1 U9864 ( .A1(n8239), .A2(n8238), .ZN(n8335) );
  AOI21_X1 U9865 ( .B1(n8239), .B2(n8238), .A(n8335), .ZN(n8240) );
  NAND2_X1 U9866 ( .A1(n8240), .A2(n8241), .ZN(n8337) );
  OAI21_X1 U9867 ( .B1(n8241), .B2(n8240), .A(n8337), .ZN(n8242) );
  NAND2_X1 U9868 ( .A1(n8242), .A2(n9772), .ZN(n8248) );
  AOI21_X1 U9869 ( .B1(n9780), .B2(n9801), .A(n8243), .ZN(n8244) );
  OAI21_X1 U9870 ( .B1(n7097), .B2(n9778), .A(n8244), .ZN(n8245) );
  AOI21_X1 U9871 ( .B1(n9784), .B2(n8246), .A(n8245), .ZN(n8247) );
  OAI211_X1 U9872 ( .C1(n9782), .C2(n8249), .A(n8248), .B(n8247), .ZN(P1_U3225) );
  OAI222_X1 U9873 ( .A1(n10238), .A2(n8251), .B1(n4391), .B2(n8959), .C1(
        P1_U3084), .C2(n8250), .ZN(P1_U3331) );
  NAND2_X1 U9874 ( .A1(n8253), .A2(n8252), .ZN(n8254) );
  XNOR2_X1 U9875 ( .A(n8255), .B(n8254), .ZN(n10410) );
  INV_X1 U9876 ( .A(n10410), .ZN(n8271) );
  NOR2_X1 U9877 ( .A1(n10020), .A2(n8256), .ZN(n10081) );
  OR2_X1 U9878 ( .A1(n8257), .A2(n8346), .ZN(n8258) );
  NAND2_X1 U9879 ( .A1(n8259), .A2(n8258), .ZN(n10414) );
  AOI22_X1 U9880 ( .A1(n10060), .A2(n8260), .B1(n10059), .B2(n8345), .ZN(n8261) );
  OAI21_X1 U9881 ( .B1(n10063), .B2(n10414), .A(n8261), .ZN(n8270) );
  NAND2_X1 U9882 ( .A1(n8263), .A2(n8262), .ZN(n8265) );
  XNOR2_X1 U9883 ( .A(n8265), .B(n8264), .ZN(n8266) );
  NAND2_X1 U9884 ( .A1(n8266), .A2(n10074), .ZN(n8268) );
  AOI22_X1 U9885 ( .A1(n9800), .A2(n10068), .B1(n10011), .B2(n9802), .ZN(n8267) );
  OAI211_X1 U9886 ( .C1(n10410), .C2(n10090), .A(n8268), .B(n8267), .ZN(n10417) );
  MUX2_X1 U9887 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10417), .S(n10078), .Z(n8269) );
  AOI211_X1 U9888 ( .C1(n8271), .C2(n10081), .A(n8270), .B(n8269), .ZN(n8272)
         );
  INV_X1 U9889 ( .A(n8272), .ZN(P1_U3285) );
  INV_X1 U9890 ( .A(n8331), .ZN(n8275) );
  AOI21_X1 U9891 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n9621), .A(n8273), .ZN(
        n8274) );
  OAI21_X1 U9892 ( .B1(n8275), .B2(n9627), .A(n8274), .ZN(P2_U3335) );
  NOR2_X1 U9893 ( .A1(n8386), .A2(n8865), .ZN(n8282) );
  AOI21_X1 U9894 ( .B1(n10427), .B2(n8869), .A(n8282), .ZN(n8523) );
  INV_X1 U9895 ( .A(n8523), .ZN(n8522) );
  XNOR2_X1 U9896 ( .A(n8525), .B(n8522), .ZN(n8283) );
  XNOR2_X1 U9897 ( .A(n8462), .B(n8283), .ZN(n8290) );
  NAND2_X1 U9898 ( .A1(n9780), .A2(n9798), .ZN(n8285) );
  OAI211_X1 U9899 ( .C1(n9778), .C2(n8286), .A(n8285), .B(n8284), .ZN(n8287)
         );
  AOI21_X1 U9900 ( .B1(n9713), .B2(n8324), .A(n8287), .ZN(n8289) );
  NAND2_X1 U9901 ( .A1(n9784), .A2(n10427), .ZN(n8288) );
  OAI211_X1 U9902 ( .C1(n8290), .C2(n9760), .A(n8289), .B(n8288), .ZN(P1_U3219) );
  NOR2_X1 U9903 ( .A1(n8291), .A2(n8299), .ZN(n8539) );
  INV_X1 U9904 ( .A(n8539), .ZN(n8292) );
  OAI21_X1 U9905 ( .B1(n8294), .B2(n8293), .A(n8292), .ZN(n8303) );
  INV_X1 U9906 ( .A(n8295), .ZN(n8296) );
  NOR2_X1 U9907 ( .A1(n8297), .A2(n8296), .ZN(n8298) );
  NAND2_X1 U9908 ( .A1(n8298), .A2(n8299), .ZN(n8542) );
  OAI21_X1 U9909 ( .B1(n8299), .B2(n8298), .A(n8542), .ZN(n8300) );
  NAND2_X1 U9910 ( .A1(n8300), .A2(n9385), .ZN(n8302) );
  AOI22_X1 U9911 ( .A1(n9446), .A2(n9121), .B1(n9444), .B2(n9119), .ZN(n8301)
         );
  OAI211_X1 U9912 ( .C1(n9425), .C2(n8303), .A(n8302), .B(n8301), .ZN(n8366)
         );
  INV_X1 U9913 ( .A(n8366), .ZN(n8313) );
  INV_X1 U9914 ( .A(n8303), .ZN(n8368) );
  NOR2_X1 U9915 ( .A1(n10461), .A2(n8304), .ZN(n9396) );
  OAI21_X1 U9916 ( .B1(n8306), .B2(n8364), .A(n8305), .ZN(n8365) );
  AOI22_X1 U9917 ( .A1(n10461), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n8307), .B2(
        n10462), .ZN(n8310) );
  NAND2_X1 U9918 ( .A1(n9469), .A2(n8308), .ZN(n8309) );
  OAI211_X1 U9919 ( .C1(n10465), .C2(n8365), .A(n8310), .B(n8309), .ZN(n8311)
         );
  AOI21_X1 U9920 ( .B1(n8368), .B2(n9396), .A(n8311), .ZN(n8312) );
  OAI21_X1 U9921 ( .B1(n8313), .B2(n10470), .A(n8312), .ZN(P2_U3288) );
  OAI21_X1 U9922 ( .B1(n8316), .B2(n8315), .A(n8314), .ZN(n10433) );
  NAND2_X1 U9923 ( .A1(n8318), .A2(n8317), .ZN(n8320) );
  XNOR2_X1 U9924 ( .A(n8320), .B(n8319), .ZN(n8321) );
  AOI222_X1 U9925 ( .A1(n9800), .A2(n10011), .B1(n10074), .B2(n8321), .C1(
        n9798), .C2(n10068), .ZN(n10432) );
  MUX2_X1 U9926 ( .A(n5167), .B(n10432), .S(n10078), .Z(n8329) );
  INV_X1 U9927 ( .A(n8379), .ZN(n8322) );
  AOI21_X1 U9928 ( .B1(n10427), .B2(n8323), .A(n8322), .ZN(n10430) );
  INV_X1 U9929 ( .A(n10427), .ZN(n8326) );
  INV_X1 U9930 ( .A(n8324), .ZN(n8325) );
  OAI22_X1 U9931 ( .A1(n9999), .A2(n8326), .B1(n10049), .B2(n8325), .ZN(n8327)
         );
  AOI21_X1 U9932 ( .B1(n10430), .B2(n10007), .A(n8327), .ZN(n8328) );
  OAI211_X1 U9933 ( .C1(n10009), .C2(n10433), .A(n8329), .B(n8328), .ZN(
        P1_U3283) );
  NAND2_X1 U9934 ( .A1(n8331), .A2(n8330), .ZN(n8333) );
  OAI211_X1 U9935 ( .C1(n8334), .C2(n10238), .A(n8333), .B(n8332), .ZN(
        P1_U3330) );
  INV_X1 U9936 ( .A(n8335), .ZN(n8336) );
  NAND2_X1 U9937 ( .A1(n8337), .A2(n8336), .ZN(n8341) );
  NAND2_X1 U9938 ( .A1(n8339), .A2(n8338), .ZN(n8340) );
  XNOR2_X1 U9939 ( .A(n8341), .B(n8340), .ZN(n8350) );
  NAND2_X1 U9940 ( .A1(n9780), .A2(n9800), .ZN(n8342) );
  NAND2_X1 U9941 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9821) );
  OAI211_X1 U9942 ( .C1(n9778), .C2(n8343), .A(n8342), .B(n9821), .ZN(n8344)
         );
  AOI21_X1 U9943 ( .B1(n9713), .B2(n8345), .A(n8344), .ZN(n8349) );
  NOR2_X1 U9944 ( .A1(n8346), .A2(n10400), .ZN(n10411) );
  NAND2_X1 U9945 ( .A1(n8347), .A2(n10411), .ZN(n8348) );
  OAI211_X1 U9946 ( .C1(n8350), .C2(n9760), .A(n8349), .B(n8348), .ZN(P1_U3237) );
  XOR2_X1 U9947 ( .A(n8352), .B(n8351), .Z(n8362) );
  NOR2_X1 U9948 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8353), .ZN(n8354) );
  AOI21_X1 U9949 ( .B1(n9174), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n8354), .ZN(
        n8355) );
  OAI21_X1 U9950 ( .B1(n9178), .B2(n8356), .A(n8355), .ZN(n8361) );
  AOI211_X1 U9951 ( .C1(n8359), .C2(n8358), .A(n9184), .B(n8357), .ZN(n8360)
         );
  AOI211_X1 U9952 ( .C1(n9169), .C2(n8362), .A(n8361), .B(n8360), .ZN(n8363)
         );
  INV_X1 U9953 ( .A(n8363), .ZN(P2_U3255) );
  OAI22_X1 U9954 ( .A1(n8365), .A2(n10508), .B1(n8364), .B2(n10507), .ZN(n8367) );
  AOI211_X1 U9955 ( .C1(n9552), .C2(n8368), .A(n8367), .B(n8366), .ZN(n8371)
         );
  NAND2_X1 U9956 ( .A1(n10514), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8369) );
  OAI21_X1 U9957 ( .B1(n8371), .B2(n10514), .A(n8369), .ZN(P2_U3475) );
  NAND2_X1 U9958 ( .A1(n10523), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8370) );
  OAI21_X1 U9959 ( .B1(n8371), .B2(n10523), .A(n8370), .ZN(P2_U3528) );
  XNOR2_X1 U9960 ( .A(n8373), .B(n8372), .ZN(n8377) );
  AOI22_X1 U9961 ( .A1(n9103), .A2(n9116), .B1(n9102), .B2(n9431), .ZN(n8374)
         );
  NAND2_X1 U9962 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8727) );
  OAI211_X1 U9963 ( .C1(n9106), .C2(n9420), .A(n8374), .B(n8727), .ZN(n8375)
         );
  AOI21_X1 U9964 ( .B1(n9565), .B2(n9108), .A(n8375), .ZN(n8376) );
  OAI21_X1 U9965 ( .B1(n8377), .B2(n9110), .A(n8376), .ZN(P2_U3236) );
  XNOR2_X1 U9966 ( .A(n8378), .B(n8384), .ZN(n8502) );
  INV_X1 U9967 ( .A(n8506), .ZN(n8381) );
  NAND2_X1 U9968 ( .A1(n8379), .A2(n8535), .ZN(n8380) );
  NAND2_X1 U9969 ( .A1(n8381), .A2(n8380), .ZN(n8498) );
  INV_X1 U9970 ( .A(n8535), .ZN(n8382) );
  OAI22_X1 U9971 ( .A1(n8498), .A2(n10413), .B1(n8382), .B2(n10400), .ZN(n8391) );
  INV_X1 U9972 ( .A(n10090), .ZN(n10386) );
  NAND2_X1 U9973 ( .A1(n8502), .A2(n10386), .ZN(n8390) );
  INV_X1 U9974 ( .A(n8384), .ZN(n8385) );
  XNOR2_X1 U9975 ( .A(n8383), .B(n8385), .ZN(n8388) );
  OAI22_X1 U9976 ( .A1(n8386), .A2(n10071), .B1(n8533), .B2(n10040), .ZN(n8387) );
  AOI21_X1 U9977 ( .B1(n8388), .B2(n10074), .A(n8387), .ZN(n8389) );
  NAND2_X1 U9978 ( .A1(n8390), .A2(n8389), .ZN(n8499) );
  AOI211_X1 U9979 ( .C1(n10184), .C2(n8502), .A(n8391), .B(n8499), .ZN(n8394)
         );
  NAND2_X1 U9980 ( .A1(n10452), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n8392) );
  OAI21_X1 U9981 ( .B1(n8394), .B2(n10452), .A(n8392), .ZN(P1_U3532) );
  NAND2_X1 U9982 ( .A1(n10435), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8393) );
  OAI21_X1 U9983 ( .B1(n8394), .B2(n10435), .A(n8393), .ZN(P1_U3481) );
  NAND2_X1 U9984 ( .A1(n8535), .A2(n8785), .ZN(n8396) );
  NAND2_X1 U9985 ( .A1(n9798), .A2(n8004), .ZN(n8395) );
  NAND2_X1 U9986 ( .A1(n8396), .A2(n8395), .ZN(n8397) );
  XNOR2_X1 U9987 ( .A(n8397), .B(n8836), .ZN(n8400) );
  NAND2_X1 U9988 ( .A1(n8535), .A2(n8869), .ZN(n8399) );
  NAND2_X1 U9989 ( .A1(n9798), .A2(n8874), .ZN(n8398) );
  NAND2_X1 U9990 ( .A1(n8399), .A2(n8398), .ZN(n8401) );
  OAI21_X1 U9991 ( .B1(n8525), .B2(n8523), .A(n8521), .ZN(n8435) );
  OR2_X1 U9992 ( .A1(n8462), .A2(n8435), .ZN(n8405) );
  NAND3_X1 U9993 ( .A1(n8525), .A2(n8523), .A3(n8521), .ZN(n8404) );
  INV_X1 U9994 ( .A(n8400), .ZN(n8403) );
  INV_X1 U9995 ( .A(n8401), .ZN(n8402) );
  NAND2_X1 U9996 ( .A1(n8403), .A2(n8402), .ZN(n8520) );
  AND2_X1 U9997 ( .A1(n8404), .A2(n8520), .ZN(n8437) );
  NAND2_X1 U9998 ( .A1(n8405), .A2(n8437), .ZN(n8416) );
  NAND2_X1 U9999 ( .A1(n8641), .A2(n8785), .ZN(n8407) );
  OR2_X1 U10000 ( .A1(n8533), .A2(n4401), .ZN(n8406) );
  NAND2_X1 U10001 ( .A1(n8407), .A2(n8406), .ZN(n8408) );
  XNOR2_X1 U10002 ( .A(n8408), .B(n8836), .ZN(n8411) );
  NAND2_X1 U10003 ( .A1(n8641), .A2(n8869), .ZN(n8410) );
  OR2_X1 U10004 ( .A1(n8533), .A2(n8865), .ZN(n8409) );
  NAND2_X1 U10005 ( .A1(n8410), .A2(n8409), .ZN(n8412) );
  NAND2_X1 U10006 ( .A1(n8411), .A2(n8412), .ZN(n8434) );
  INV_X1 U10007 ( .A(n8411), .ZN(n8414) );
  INV_X1 U10008 ( .A(n8412), .ZN(n8413) );
  NAND2_X1 U10009 ( .A1(n8414), .A2(n8413), .ZN(n8436) );
  NAND2_X1 U10010 ( .A1(n8434), .A2(n8436), .ZN(n8415) );
  XNOR2_X1 U10011 ( .A(n8416), .B(n8415), .ZN(n8422) );
  NAND2_X1 U10012 ( .A1(n9780), .A2(n9796), .ZN(n8418) );
  OAI211_X1 U10013 ( .C1(n9778), .C2(n8511), .A(n8418), .B(n8417), .ZN(n8420)
         );
  NOR2_X1 U10014 ( .A1(n9771), .A2(n8507), .ZN(n8419) );
  AOI211_X1 U10015 ( .C1(n8640), .C2(n9713), .A(n8420), .B(n8419), .ZN(n8421)
         );
  OAI21_X1 U10016 ( .B1(n8422), .B2(n9760), .A(n8421), .ZN(P1_U3215) );
  AOI21_X1 U10017 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n8424), .A(n8423), .ZN(
        n8433) );
  NAND2_X1 U10018 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9644) );
  OAI21_X1 U10019 ( .B1(n10339), .B2(n8425), .A(n9644), .ZN(n8431) );
  AOI21_X1 U10020 ( .B1(n8428), .B2(n8427), .A(n8426), .ZN(n8429) );
  NOR2_X1 U10021 ( .A1(n8429), .A2(n10300), .ZN(n8430) );
  AOI211_X1 U10022 ( .C1(n10342), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n8431), .B(
        n8430), .ZN(n8432) );
  OAI21_X1 U10023 ( .B1(n8433), .B2(n10305), .A(n8432), .ZN(P1_U3255) );
  INV_X1 U10024 ( .A(n10196), .ZN(n8568) );
  INV_X1 U10025 ( .A(n8434), .ZN(n8438) );
  OR2_X1 U10026 ( .A1(n8435), .A2(n8438), .ZN(n8460) );
  OR2_X1 U10027 ( .A1(n8462), .A2(n8460), .ZN(n8448) );
  NAND2_X1 U10028 ( .A1(n8448), .A2(n8446), .ZN(n8444) );
  NAND2_X1 U10029 ( .A1(n10196), .A2(n8785), .ZN(n8441) );
  NAND2_X1 U10030 ( .A1(n9796), .A2(n8869), .ZN(n8440) );
  NAND2_X1 U10031 ( .A1(n8441), .A2(n8440), .ZN(n8442) );
  XNOR2_X1 U10032 ( .A(n8442), .B(n8872), .ZN(n8456) );
  AND2_X1 U10033 ( .A1(n9796), .A2(n8874), .ZN(n8443) );
  AOI21_X1 U10034 ( .B1(n10196), .B2(n8869), .A(n8443), .ZN(n8457) );
  XNOR2_X1 U10035 ( .A(n8456), .B(n8457), .ZN(n8445) );
  AOI21_X1 U10036 ( .B1(n8444), .B2(n8445), .A(n9760), .ZN(n8450) );
  INV_X1 U10037 ( .A(n8445), .ZN(n8447) );
  NAND2_X1 U10038 ( .A1(n8448), .A2(n8463), .ZN(n8449) );
  NAND2_X1 U10039 ( .A1(n8450), .A2(n8449), .ZN(n8455) );
  AOI21_X1 U10040 ( .B1(n9780), .B2(n9795), .A(n8451), .ZN(n8452) );
  OAI21_X1 U10041 ( .B1(n8533), .B2(n9778), .A(n8452), .ZN(n8453) );
  AOI21_X1 U10042 ( .B1(n8566), .B2(n9713), .A(n8453), .ZN(n8454) );
  OAI211_X1 U10043 ( .C1(n8568), .C2(n9771), .A(n8455), .B(n8454), .ZN(
        P1_U3234) );
  INV_X1 U10044 ( .A(n8456), .ZN(n8459) );
  INV_X1 U10045 ( .A(n8457), .ZN(n8458) );
  AND2_X1 U10046 ( .A1(n8459), .A2(n8458), .ZN(n8464) );
  OR2_X1 U10047 ( .A1(n8460), .A2(n8464), .ZN(n8461) );
  OR2_X2 U10048 ( .A1(n8462), .A2(n8461), .ZN(n8583) );
  AND2_X1 U10049 ( .A1(n8583), .A2(n8580), .ZN(n8470) );
  NAND2_X1 U10050 ( .A1(n10193), .A2(n8785), .ZN(n8466) );
  OR2_X1 U10051 ( .A1(n10072), .A2(n4401), .ZN(n8465) );
  NAND2_X1 U10052 ( .A1(n8466), .A2(n8465), .ZN(n8467) );
  XNOR2_X1 U10053 ( .A(n8467), .B(n8872), .ZN(n8584) );
  NOR2_X1 U10054 ( .A1(n10072), .A2(n8865), .ZN(n8468) );
  AOI21_X1 U10055 ( .B1(n10193), .B2(n8869), .A(n8468), .ZN(n8579) );
  INV_X1 U10056 ( .A(n8579), .ZN(n8585) );
  XNOR2_X1 U10057 ( .A(n8584), .B(n8585), .ZN(n8469) );
  XNOR2_X1 U10058 ( .A(n8470), .B(n8469), .ZN(n8476) );
  NAND2_X1 U10059 ( .A1(n9713), .A2(n8635), .ZN(n8473) );
  AOI21_X1 U10060 ( .B1(n9780), .B2(n9794), .A(n8471), .ZN(n8472) );
  OAI211_X1 U10061 ( .C1(n8510), .C2(n9778), .A(n8473), .B(n8472), .ZN(n8474)
         );
  AOI21_X1 U10062 ( .B1(n9784), .B2(n10193), .A(n8474), .ZN(n8475) );
  OAI21_X1 U10063 ( .B1(n8476), .B2(n9760), .A(n8475), .ZN(P1_U3222) );
  INV_X1 U10064 ( .A(n8477), .ZN(n8494) );
  OAI222_X1 U10065 ( .A1(P1_U3084), .A2(n8479), .B1(n4391), .B2(n8494), .C1(
        n8478), .C2(n10238), .ZN(P1_U3329) );
  OAI21_X1 U10066 ( .B1(n8482), .B2(n8481), .A(n8480), .ZN(n8491) );
  XOR2_X1 U10067 ( .A(n8484), .B(n8483), .Z(n8485) );
  NAND2_X1 U10068 ( .A1(n8485), .A2(n9169), .ZN(n8488) );
  NOR2_X1 U10069 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6296), .ZN(n8486) );
  AOI21_X1 U10070 ( .B1(n9174), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n8486), .ZN(
        n8487) );
  OAI211_X1 U10071 ( .C1(n9178), .C2(n8489), .A(n8488), .B(n8487), .ZN(n8490)
         );
  AOI21_X1 U10072 ( .B1(n8491), .B2(n9163), .A(n8490), .ZN(n8492) );
  INV_X1 U10073 ( .A(n8492), .ZN(P2_U3256) );
  INV_X1 U10074 ( .A(n8493), .ZN(n8495) );
  OAI222_X1 U10075 ( .A1(n9624), .A2(n8496), .B1(P2_U3152), .B2(n8495), .C1(
        n9627), .C2(n8494), .ZN(P2_U3334) );
  AOI22_X1 U10076 ( .A1(n10060), .A2(n8535), .B1(n10059), .B2(n8529), .ZN(
        n8497) );
  OAI21_X1 U10077 ( .B1(n8498), .B2(n10063), .A(n8497), .ZN(n8501) );
  MUX2_X1 U10078 ( .A(n8499), .B(P1_REG2_REG_9__SCAN_IN), .S(n10020), .Z(n8500) );
  AOI211_X1 U10079 ( .C1(n8502), .C2(n10081), .A(n8501), .B(n8500), .ZN(n8503)
         );
  INV_X1 U10080 ( .A(n8503), .ZN(P1_U3282) );
  XNOR2_X1 U10081 ( .A(n8504), .B(n8505), .ZN(n8515) );
  INV_X1 U10082 ( .A(n8515), .ZN(n8648) );
  OAI211_X1 U10083 ( .C1(n8506), .C2(n8507), .A(n8565), .B(n10429), .ZN(n8644)
         );
  OAI21_X1 U10084 ( .B1(n8507), .B2(n10400), .A(n8644), .ZN(n8516) );
  XNOR2_X1 U10085 ( .A(n8509), .B(n8508), .ZN(n8513) );
  OAI22_X1 U10086 ( .A1(n8511), .A2(n10071), .B1(n8510), .B2(n10040), .ZN(
        n8512) );
  AOI21_X1 U10087 ( .B1(n8513), .B2(n10074), .A(n8512), .ZN(n8514) );
  OAI21_X1 U10088 ( .B1(n8515), .B2(n10090), .A(n8514), .ZN(n8645) );
  AOI211_X1 U10089 ( .C1(n10184), .C2(n8648), .A(n8516), .B(n8645), .ZN(n8519)
         );
  NAND2_X1 U10090 ( .A1(n10435), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n8517) );
  OAI21_X1 U10091 ( .B1(n8519), .B2(n10435), .A(n8517), .ZN(P1_U3484) );
  NAND2_X1 U10092 ( .A1(n10452), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8518) );
  OAI21_X1 U10093 ( .B1(n8519), .B2(n10452), .A(n8518), .ZN(P1_U3533) );
  NAND2_X1 U10094 ( .A1(n8521), .A2(n8520), .ZN(n8528) );
  NOR2_X1 U10095 ( .A1(n8462), .A2(n8522), .ZN(n8526) );
  INV_X1 U10096 ( .A(n8462), .ZN(n8524) );
  OAI22_X1 U10097 ( .A1(n8526), .A2(n8525), .B1(n8524), .B2(n8523), .ZN(n8527)
         );
  XOR2_X1 U10098 ( .A(n8528), .B(n8527), .Z(n8537) );
  NAND2_X1 U10099 ( .A1(n9713), .A2(n8529), .ZN(n8532) );
  AOI21_X1 U10100 ( .B1(n9735), .B2(n9799), .A(n8530), .ZN(n8531) );
  OAI211_X1 U10101 ( .C1(n8533), .C2(n9683), .A(n8532), .B(n8531), .ZN(n8534)
         );
  AOI21_X1 U10102 ( .B1(n9784), .B2(n8535), .A(n8534), .ZN(n8536) );
  OAI21_X1 U10103 ( .B1(n8537), .B2(n9760), .A(n8536), .ZN(P1_U3229) );
  NOR2_X1 U10104 ( .A1(n8539), .A2(n8538), .ZN(n8540) );
  XNOR2_X1 U10105 ( .A(n8540), .B(n8544), .ZN(n9593) );
  INV_X1 U10106 ( .A(n9396), .ZN(n9434) );
  NAND2_X1 U10107 ( .A1(n8542), .A2(n8541), .ZN(n8543) );
  XNOR2_X1 U10108 ( .A(n8544), .B(n8543), .ZN(n8549) );
  OAI22_X1 U10109 ( .A1(n8546), .A2(n9419), .B1(n9418), .B2(n8545), .ZN(n8548)
         );
  NOR2_X1 U10110 ( .A1(n9593), .A2(n9425), .ZN(n8547) );
  AOI211_X1 U10111 ( .C1(n8549), .C2(n9385), .A(n8548), .B(n8547), .ZN(n9592)
         );
  MUX2_X1 U10112 ( .A(n8550), .B(n9592), .S(n9457), .Z(n8557) );
  NAND2_X1 U10113 ( .A1(n8305), .A2(n9587), .ZN(n8551) );
  AND2_X1 U10114 ( .A1(n8213), .A2(n8551), .ZN(n9590) );
  INV_X1 U10115 ( .A(n8552), .ZN(n8553) );
  OAI22_X1 U10116 ( .A1(n10464), .A2(n8554), .B1(n8553), .B2(n9290), .ZN(n8555) );
  AOI21_X1 U10117 ( .B1(n9464), .B2(n9590), .A(n8555), .ZN(n8556) );
  OAI211_X1 U10118 ( .C1(n9593), .C2(n9434), .A(n8557), .B(n8556), .ZN(
        P2_U3287) );
  XOR2_X1 U10119 ( .A(n8619), .B(n8558), .Z(n8563) );
  INV_X1 U10120 ( .A(n8563), .ZN(n10200) );
  INV_X1 U10121 ( .A(n10081), .ZN(n8572) );
  XNOR2_X1 U10122 ( .A(n8559), .B(n8558), .ZN(n8561) );
  AOI22_X1 U10123 ( .A1(n10011), .A2(n9797), .B1(n9795), .B2(n10068), .ZN(
        n8560) );
  OAI21_X1 U10124 ( .B1(n8561), .B2(n10044), .A(n8560), .ZN(n8562) );
  AOI21_X1 U10125 ( .B1(n8563), .B2(n10386), .A(n8562), .ZN(n10199) );
  MUX2_X1 U10126 ( .A(n5169), .B(n10199), .S(n10078), .Z(n8571) );
  INV_X1 U10127 ( .A(n8632), .ZN(n8564) );
  AOI21_X1 U10128 ( .B1(n10196), .B2(n8565), .A(n8564), .ZN(n10197) );
  INV_X1 U10129 ( .A(n8566), .ZN(n8567) );
  OAI22_X1 U10130 ( .A1(n8568), .A2(n9999), .B1(n8567), .B2(n10049), .ZN(n8569) );
  AOI21_X1 U10131 ( .B1(n10197), .B2(n10007), .A(n8569), .ZN(n8570) );
  OAI211_X1 U10132 ( .C1(n10200), .C2(n8572), .A(n8571), .B(n8570), .ZN(
        P1_U3280) );
  INV_X1 U10133 ( .A(n8573), .ZN(n8577) );
  OAI222_X1 U10134 ( .A1(n10238), .A2(n8575), .B1(n4391), .B2(n8577), .C1(
        P1_U3084), .C2(n8574), .ZN(P1_U3328) );
  OAI222_X1 U10135 ( .A1(n9624), .A2(n8578), .B1(n9627), .B2(n8577), .C1(n8576), .C2(P2_U3152), .ZN(P2_U3333) );
  NAND2_X1 U10136 ( .A1(n8584), .A2(n8579), .ZN(n8581) );
  INV_X1 U10137 ( .A(n8584), .ZN(n8586) );
  NAND2_X1 U10138 ( .A1(n8586), .A2(n8585), .ZN(n8587) );
  NAND2_X1 U10139 ( .A1(n10061), .A2(n8785), .ZN(n8589) );
  NAND2_X1 U10140 ( .A1(n9794), .A2(n8869), .ZN(n8588) );
  NAND2_X1 U10141 ( .A1(n8589), .A2(n8588), .ZN(n8590) );
  XNOR2_X1 U10142 ( .A(n8590), .B(n8836), .ZN(n8593) );
  NAND2_X1 U10143 ( .A1(n10061), .A2(n8869), .ZN(n8592) );
  NAND2_X1 U10144 ( .A1(n9794), .A2(n8874), .ZN(n8591) );
  NAND2_X1 U10145 ( .A1(n8592), .A2(n8591), .ZN(n8594) );
  AND2_X1 U10146 ( .A1(n8593), .A2(n8594), .ZN(n8598) );
  INV_X1 U10147 ( .A(n8593), .ZN(n8596) );
  INV_X1 U10148 ( .A(n8594), .ZN(n8595) );
  NAND2_X1 U10149 ( .A1(n8596), .A2(n8595), .ZN(n8746) );
  INV_X1 U10150 ( .A(n8746), .ZN(n8600) );
  OAI21_X1 U10151 ( .B1(n8600), .B2(n8598), .A(n8597), .ZN(n8599) );
  OAI21_X1 U10152 ( .B1(n8747), .B2(n8600), .A(n8599), .ZN(n8601) );
  NAND2_X1 U10153 ( .A1(n8601), .A2(n9772), .ZN(n8606) );
  AOI21_X1 U10154 ( .B1(n9780), .B2(n10069), .A(n8602), .ZN(n8603) );
  OAI21_X1 U10155 ( .B1(n10072), .B2(n9778), .A(n8603), .ZN(n8604) );
  AOI21_X1 U10156 ( .B1(n10058), .B2(n9713), .A(n8604), .ZN(n8605) );
  OAI211_X1 U10157 ( .C1(n10186), .C2(n9771), .A(n8606), .B(n8605), .ZN(
        P1_U3232) );
  OAI21_X1 U10158 ( .B1(n8609), .B2(n8608), .A(n8607), .ZN(n8610) );
  NAND2_X1 U10159 ( .A1(n8610), .A2(n9048), .ZN(n8617) );
  NAND2_X1 U10160 ( .A1(n9444), .A2(n9381), .ZN(n8612) );
  NAND2_X1 U10161 ( .A1(n9446), .A2(n9115), .ZN(n8611) );
  NAND2_X1 U10162 ( .A1(n8612), .A2(n8611), .ZN(n8668) );
  NOR2_X1 U10163 ( .A1(n8613), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9131) );
  NOR2_X1 U10164 ( .A1(n9095), .A2(n8673), .ZN(n8614) );
  AOI211_X1 U10165 ( .C1(n8615), .C2(n8668), .A(n9131), .B(n8614), .ZN(n8616)
         );
  OAI211_X1 U10166 ( .C1(n8676), .C2(n9023), .A(n8617), .B(n8616), .ZN(
        P2_U3217) );
  OR2_X1 U10167 ( .A1(n8619), .A2(n8618), .ZN(n8621) );
  NAND2_X1 U10168 ( .A1(n8621), .A2(n8620), .ZN(n8622) );
  XNOR2_X1 U10169 ( .A(n8622), .B(n8625), .ZN(n10195) );
  NAND2_X1 U10170 ( .A1(n8624), .A2(n8623), .ZN(n8626) );
  XNOR2_X1 U10171 ( .A(n8625), .B(n8626), .ZN(n8627) );
  NAND2_X1 U10172 ( .A1(n8627), .A2(n10074), .ZN(n8629) );
  AOI22_X1 U10173 ( .A1(n10011), .A2(n9796), .B1(n9794), .B2(n10068), .ZN(
        n8628) );
  NAND2_X1 U10174 ( .A1(n8629), .A2(n8628), .ZN(n10191) );
  INV_X1 U10175 ( .A(n10191), .ZN(n8630) );
  MUX2_X1 U10176 ( .A(n5170), .B(n8630), .S(n10078), .Z(n8639) );
  NAND2_X1 U10177 ( .A1(n8632), .A2(n10193), .ZN(n8633) );
  NAND2_X1 U10178 ( .A1(n8633), .A2(n10429), .ZN(n8634) );
  NOR2_X1 U10179 ( .A1(n8631), .A2(n8634), .ZN(n10192) );
  INV_X1 U10180 ( .A(n8635), .ZN(n8636) );
  OAI22_X1 U10181 ( .A1(n5017), .A2(n9999), .B1(n10049), .B2(n8636), .ZN(n8637) );
  AOI21_X1 U10182 ( .B1(n10192), .B2(n10024), .A(n8637), .ZN(n8638) );
  OAI211_X1 U10183 ( .C1(n10009), .C2(n10195), .A(n8639), .B(n8638), .ZN(
        P1_U3279) );
  AOI22_X1 U10184 ( .A1(n10060), .A2(n8641), .B1(n8640), .B2(n10059), .ZN(
        n8642) );
  OAI21_X1 U10185 ( .B1(n8644), .B2(n8643), .A(n8642), .ZN(n8647) );
  MUX2_X1 U10186 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n8645), .S(n10078), .Z(
        n8646) );
  AOI211_X1 U10187 ( .C1(n10081), .C2(n8648), .A(n8647), .B(n8646), .ZN(n8649)
         );
  INV_X1 U10188 ( .A(n8649), .ZN(P1_U3281) );
  OR2_X1 U10189 ( .A1(n8226), .A2(n8650), .ZN(n8652) );
  NAND2_X1 U10190 ( .A1(n8652), .A2(n8651), .ZN(n8654) );
  AOI21_X1 U10191 ( .B1(n8654), .B2(n8653), .A(n9263), .ZN(n8659) );
  OR2_X1 U10192 ( .A1(n8654), .A2(n8653), .ZN(n8658) );
  OAI22_X1 U10193 ( .A1(n8656), .A2(n9419), .B1(n9418), .B2(n8655), .ZN(n8657)
         );
  AOI21_X1 U10194 ( .B1(n8659), .B2(n8658), .A(n8657), .ZN(n9572) );
  XOR2_X1 U10195 ( .A(n8660), .B(n6570), .Z(n9570) );
  AOI22_X1 U10196 ( .A1(n10470), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n8996), 
        .B2(n10462), .ZN(n8661) );
  OAI21_X1 U10197 ( .B1(n10464), .B2(n6571), .A(n8661), .ZN(n8665) );
  NOR2_X1 U10198 ( .A1(n8662), .A2(n8663), .ZN(n9422) );
  AOI21_X1 U10199 ( .B1(n8663), .B2(n8662), .A(n9422), .ZN(n9573) );
  NOR2_X1 U10200 ( .A1(n9573), .A2(n9411), .ZN(n8664) );
  AOI211_X1 U10201 ( .C1(n9570), .C2(n9464), .A(n8665), .B(n8664), .ZN(n8666)
         );
  OAI21_X1 U10202 ( .B1(n10461), .B2(n9572), .A(n8666), .ZN(P2_U3284) );
  AOI21_X1 U10203 ( .B1(n8667), .B2(n8680), .A(n9263), .ZN(n8670) );
  AOI21_X1 U10204 ( .B1(n8670), .B2(n8669), .A(n8668), .ZN(n9563) );
  INV_X1 U10205 ( .A(n9429), .ZN(n8672) );
  AOI211_X1 U10206 ( .C1(n6337), .C2(n8672), .A(n10508), .B(n8671), .ZN(n9561)
         );
  INV_X1 U10207 ( .A(n8673), .ZN(n8674) );
  AOI22_X1 U10208 ( .A1(n10470), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8674), 
        .B2(n10462), .ZN(n8675) );
  OAI21_X1 U10209 ( .B1(n8676), .B2(n10464), .A(n8675), .ZN(n8683) );
  INV_X1 U10210 ( .A(n8662), .ZN(n8679) );
  OAI21_X1 U10211 ( .B1(n8679), .B2(n8678), .A(n8677), .ZN(n8681) );
  XNOR2_X1 U10212 ( .A(n8681), .B(n8680), .ZN(n9564) );
  NOR2_X1 U10213 ( .A1(n9564), .A2(n9411), .ZN(n8682) );
  AOI211_X1 U10214 ( .C1(n9561), .C2(n9472), .A(n8683), .B(n8682), .ZN(n8684)
         );
  OAI21_X1 U10215 ( .B1(n10461), .B2(n9563), .A(n8684), .ZN(P2_U3282) );
  INV_X1 U10216 ( .A(n8685), .ZN(n8689) );
  OAI222_X1 U10217 ( .A1(n8956), .A2(n8689), .B1(P2_U3152), .B2(n8687), .C1(
        n8686), .C2(n9624), .ZN(P2_U3332) );
  OAI222_X1 U10218 ( .A1(P1_U3084), .A2(n8690), .B1(n4391), .B2(n8689), .C1(
        n8688), .C2(n10238), .ZN(P1_U3327) );
  INV_X1 U10219 ( .A(n8691), .ZN(n8696) );
  AOI21_X1 U10220 ( .B1(n10229), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n8692), 
        .ZN(n8693) );
  OAI21_X1 U10221 ( .B1(n8696), .B2(n4391), .A(n8693), .ZN(P1_U3326) );
  OAI222_X1 U10222 ( .A1(n8956), .A2(n8696), .B1(n8695), .B2(P2_U3152), .C1(
        n8694), .C2(n9624), .ZN(P2_U3331) );
  INV_X1 U10223 ( .A(n8715), .ZN(n8699) );
  AOI21_X1 U10224 ( .B1(n10229), .B2(P2_DATAO_REG_28__SCAN_IN), .A(n8697), 
        .ZN(n8698) );
  OAI21_X1 U10225 ( .B1(n8699), .B2(n4391), .A(n8698), .ZN(P1_U3325) );
  INV_X1 U10226 ( .A(n8723), .ZN(n8700) );
  OAI21_X1 U10227 ( .B1(n8702), .B2(n8701), .A(n8700), .ZN(n8712) );
  NOR2_X1 U10228 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8703), .ZN(n8704) );
  AOI21_X1 U10229 ( .B1(n9174), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n8704), .ZN(
        n8705) );
  OAI21_X1 U10230 ( .B1(n9178), .B2(n8706), .A(n8705), .ZN(n8711) );
  AOI211_X1 U10231 ( .C1(n8709), .C2(n8708), .A(n9184), .B(n8707), .ZN(n8710)
         );
  AOI211_X1 U10232 ( .C1(n9169), .C2(n8712), .A(n8711), .B(n8710), .ZN(n8713)
         );
  INV_X1 U10233 ( .A(n8713), .ZN(P2_U3257) );
  NAND2_X1 U10234 ( .A1(n8715), .A2(n8714), .ZN(n8717) );
  OAI211_X1 U10235 ( .C1(n9624), .C2(n8718), .A(n8717), .B(n8716), .ZN(
        P2_U3330) );
  OAI21_X1 U10236 ( .B1(n8720), .B2(n4487), .A(n8719), .ZN(n8731) );
  OR3_X1 U10237 ( .A1(n8723), .A2(n8722), .A3(n8721), .ZN(n8724) );
  AOI21_X1 U10238 ( .B1(n8725), .B2(n8724), .A(n9196), .ZN(n8730) );
  NAND2_X1 U10239 ( .A1(n9174), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n8726) );
  OAI211_X1 U10240 ( .C1(n9178), .C2(n8728), .A(n8727), .B(n8726), .ZN(n8729)
         );
  AOI211_X1 U10241 ( .C1(n8731), .C2(n9163), .A(n8730), .B(n8729), .ZN(n8732)
         );
  INV_X1 U10242 ( .A(n8732), .ZN(P2_U3258) );
  XOR2_X1 U10243 ( .A(n8742), .B(n8733), .Z(n10183) );
  INV_X1 U10244 ( .A(n10057), .ZN(n8736) );
  INV_X1 U10245 ( .A(n8734), .ZN(n8735) );
  AOI211_X1 U10246 ( .C1(n10181), .C2(n8736), .A(n10413), .B(n8735), .ZN(
        n10180) );
  NOR2_X1 U10247 ( .A1(n8737), .A2(n9999), .ZN(n8740) );
  INV_X1 U10248 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n8738) );
  OAI22_X1 U10249 ( .A1(n10078), .A2(n8738), .B1(n9648), .B2(n10049), .ZN(
        n8739) );
  AOI211_X1 U10250 ( .C1(n10180), .C2(n10024), .A(n8740), .B(n8739), .ZN(n8745) );
  XNOR2_X1 U10251 ( .A(n8741), .B(n8742), .ZN(n8743) );
  OAI222_X1 U10252 ( .A1(n10040), .A2(n9698), .B1(n10071), .B2(n9645), .C1(
        n8743), .C2(n10044), .ZN(n10179) );
  NAND2_X1 U10253 ( .A1(n10179), .A2(n10078), .ZN(n8744) );
  OAI211_X1 U10254 ( .C1(n10183), .C2(n10009), .A(n8745), .B(n8744), .ZN(
        P1_U3277) );
  NAND2_X1 U10255 ( .A1(n10181), .A2(n8785), .ZN(n8749) );
  NAND2_X1 U10256 ( .A1(n10069), .A2(n8869), .ZN(n8748) );
  NAND2_X1 U10257 ( .A1(n8749), .A2(n8748), .ZN(n8750) );
  XNOR2_X1 U10258 ( .A(n8750), .B(n8872), .ZN(n8757) );
  NAND2_X1 U10259 ( .A1(n10181), .A2(n8869), .ZN(n8752) );
  NAND2_X1 U10260 ( .A1(n10069), .A2(n8874), .ZN(n8751) );
  NAND2_X1 U10261 ( .A1(n8752), .A2(n8751), .ZN(n9643) );
  NAND2_X1 U10262 ( .A1(n10170), .A2(n8785), .ZN(n8754) );
  NAND2_X1 U10263 ( .A1(n10012), .A2(n8869), .ZN(n8753) );
  NAND2_X1 U10264 ( .A1(n8754), .A2(n8753), .ZN(n8755) );
  XNOR2_X1 U10265 ( .A(n8755), .B(n8872), .ZN(n8762) );
  INV_X1 U10266 ( .A(n8756), .ZN(n8759) );
  INV_X1 U10267 ( .A(n8757), .ZN(n8758) );
  NAND2_X1 U10268 ( .A1(n10170), .A2(n8869), .ZN(n8761) );
  NAND2_X1 U10269 ( .A1(n10012), .A2(n8874), .ZN(n8760) );
  NAND2_X1 U10270 ( .A1(n8761), .A2(n8760), .ZN(n9775) );
  INV_X1 U10271 ( .A(n8762), .ZN(n8763) );
  NAND2_X1 U10272 ( .A1(n10159), .A2(n8785), .ZN(n8765) );
  NAND2_X1 U10273 ( .A1(n10013), .A2(n8869), .ZN(n8764) );
  NAND2_X1 U10274 ( .A1(n8765), .A2(n8764), .ZN(n8766) );
  XNOR2_X1 U10275 ( .A(n8766), .B(n8872), .ZN(n9710) );
  NAND2_X1 U10276 ( .A1(n10159), .A2(n8869), .ZN(n8768) );
  NAND2_X1 U10277 ( .A1(n10013), .A2(n8874), .ZN(n8767) );
  AND2_X1 U10278 ( .A1(n8768), .A2(n8767), .ZN(n8776) );
  NOR2_X1 U10279 ( .A1(n10041), .A2(n8865), .ZN(n8769) );
  AOI21_X1 U10280 ( .B1(n10165), .B2(n8869), .A(n8769), .ZN(n8775) );
  NAND2_X1 U10281 ( .A1(n10165), .A2(n8785), .ZN(n8771) );
  OR2_X1 U10282 ( .A1(n10041), .A2(n4401), .ZN(n8770) );
  NAND2_X1 U10283 ( .A1(n8771), .A2(n8770), .ZN(n8772) );
  XNOR2_X1 U10284 ( .A(n8772), .B(n8872), .ZN(n9707) );
  OAI22_X1 U10285 ( .A1(n9710), .A2(n8776), .B1(n8775), .B2(n9707), .ZN(n8773)
         );
  INV_X1 U10286 ( .A(n8773), .ZN(n8774) );
  INV_X1 U10287 ( .A(n9707), .ZN(n9705) );
  INV_X1 U10288 ( .A(n8775), .ZN(n9704) );
  INV_X1 U10289 ( .A(n8776), .ZN(n9709) );
  OAI21_X1 U10290 ( .B1(n9705), .B2(n9704), .A(n9709), .ZN(n8778) );
  NOR2_X1 U10291 ( .A1(n9709), .A2(n9704), .ZN(n8777) );
  AOI22_X1 U10292 ( .A1(n8778), .A2(n9710), .B1(n9707), .B2(n8777), .ZN(n8779)
         );
  NAND2_X1 U10293 ( .A1(n10150), .A2(n8785), .ZN(n8782) );
  NAND2_X1 U10294 ( .A1(n9793), .A2(n8869), .ZN(n8781) );
  NAND2_X1 U10295 ( .A1(n8782), .A2(n8781), .ZN(n8783) );
  XNOR2_X1 U10296 ( .A(n8783), .B(n8836), .ZN(n8795) );
  INV_X1 U10297 ( .A(n8795), .ZN(n9670) );
  AND2_X1 U10298 ( .A1(n9793), .A2(n8874), .ZN(n8784) );
  AOI21_X1 U10299 ( .B1(n10150), .B2(n8869), .A(n8784), .ZN(n9669) );
  NAND2_X1 U10300 ( .A1(n9670), .A2(n9669), .ZN(n9668) );
  NAND2_X1 U10301 ( .A1(n10156), .A2(n8785), .ZN(n8787) );
  NAND2_X1 U10302 ( .A1(n10003), .A2(n8869), .ZN(n8786) );
  NAND2_X1 U10303 ( .A1(n8787), .A2(n8786), .ZN(n8788) );
  XNOR2_X1 U10304 ( .A(n8788), .B(n8872), .ZN(n9665) );
  NOR2_X1 U10305 ( .A1(n8789), .A2(n8865), .ZN(n8790) );
  AOI21_X1 U10306 ( .B1(n10156), .B2(n8869), .A(n8790), .ZN(n9754) );
  NAND2_X1 U10307 ( .A1(n9665), .A2(n9754), .ZN(n8791) );
  NAND2_X1 U10308 ( .A1(n9668), .A2(n8791), .ZN(n8798) );
  OAI21_X1 U10309 ( .B1(n9665), .B2(n9754), .A(n9669), .ZN(n8796) );
  INV_X1 U10310 ( .A(n9669), .ZN(n8792) );
  INV_X1 U10311 ( .A(n9754), .ZN(n9667) );
  AND2_X1 U10312 ( .A1(n8792), .A2(n9667), .ZN(n8794) );
  INV_X1 U10313 ( .A(n9665), .ZN(n8793) );
  AOI22_X1 U10314 ( .A1(n8796), .A2(n8795), .B1(n8794), .B2(n8793), .ZN(n8797)
         );
  NAND2_X1 U10315 ( .A1(n10146), .A2(n8785), .ZN(n8800) );
  NAND2_X1 U10316 ( .A1(n9970), .A2(n8869), .ZN(n8799) );
  NAND2_X1 U10317 ( .A1(n8800), .A2(n8799), .ZN(n8801) );
  XNOR2_X1 U10318 ( .A(n8801), .B(n8836), .ZN(n8805) );
  NAND2_X1 U10319 ( .A1(n10146), .A2(n8869), .ZN(n8803) );
  NAND2_X1 U10320 ( .A1(n9970), .A2(n8874), .ZN(n8802) );
  NAND2_X1 U10321 ( .A1(n8803), .A2(n8802), .ZN(n8806) );
  AND2_X1 U10322 ( .A1(n8805), .A2(n8806), .ZN(n9731) );
  INV_X1 U10323 ( .A(n9731), .ZN(n8804) );
  INV_X1 U10324 ( .A(n8805), .ZN(n8808) );
  INV_X1 U10325 ( .A(n8806), .ZN(n8807) );
  NAND2_X1 U10326 ( .A1(n8808), .A2(n8807), .ZN(n9730) );
  NAND2_X1 U10327 ( .A1(n10141), .A2(n8785), .ZN(n8811) );
  OR2_X1 U10328 ( .A1(n9948), .A2(n4401), .ZN(n8810) );
  NAND2_X1 U10329 ( .A1(n8811), .A2(n8810), .ZN(n8812) );
  XNOR2_X1 U10330 ( .A(n8812), .B(n8836), .ZN(n8814) );
  NOR2_X1 U10331 ( .A1(n9948), .A2(n8865), .ZN(n8813) );
  AOI21_X1 U10332 ( .B1(n10141), .B2(n8869), .A(n8813), .ZN(n8815) );
  XNOR2_X1 U10333 ( .A(n8814), .B(n8815), .ZN(n9679) );
  INV_X1 U10334 ( .A(n8814), .ZN(n8816) );
  NAND2_X1 U10335 ( .A1(n8816), .A2(n8815), .ZN(n8817) );
  AND2_X1 U10336 ( .A1(n9903), .A2(n8874), .ZN(n8818) );
  AOI21_X1 U10337 ( .B1(n10134), .B2(n8869), .A(n8818), .ZN(n8822) );
  NAND2_X1 U10338 ( .A1(n10134), .A2(n8439), .ZN(n8820) );
  NAND2_X1 U10339 ( .A1(n9903), .A2(n8869), .ZN(n8819) );
  NAND2_X1 U10340 ( .A1(n8820), .A2(n8819), .ZN(n8821) );
  XNOR2_X1 U10341 ( .A(n8821), .B(n8872), .ZN(n9743) );
  NAND2_X1 U10342 ( .A1(n9742), .A2(n9743), .ZN(n8824) );
  NAND2_X1 U10343 ( .A1(n8823), .A2(n8822), .ZN(n9741) );
  NAND2_X1 U10344 ( .A1(n10123), .A2(n8439), .ZN(n8826) );
  NAND2_X1 U10345 ( .A1(n9792), .A2(n8869), .ZN(n8825) );
  NAND2_X1 U10346 ( .A1(n8826), .A2(n8825), .ZN(n8827) );
  XNOR2_X1 U10347 ( .A(n8827), .B(n8836), .ZN(n8852) );
  NOR2_X1 U10348 ( .A1(n9888), .A2(n8865), .ZN(n8828) );
  AOI21_X1 U10349 ( .B1(n10123), .B2(n8869), .A(n8828), .ZN(n8850) );
  XNOR2_X1 U10350 ( .A(n8852), .B(n8850), .ZN(n9689) );
  NAND2_X1 U10351 ( .A1(n10127), .A2(n8785), .ZN(n8830) );
  NAND2_X1 U10352 ( .A1(n9905), .A2(n8869), .ZN(n8829) );
  NAND2_X1 U10353 ( .A1(n8830), .A2(n8829), .ZN(n8831) );
  XNOR2_X1 U10354 ( .A(n8831), .B(n8836), .ZN(n8842) );
  NAND2_X1 U10355 ( .A1(n10127), .A2(n8869), .ZN(n8833) );
  NAND2_X1 U10356 ( .A1(n9905), .A2(n8874), .ZN(n8832) );
  NAND2_X1 U10357 ( .A1(n8833), .A2(n8832), .ZN(n8843) );
  NAND2_X1 U10358 ( .A1(n8842), .A2(n8843), .ZN(n9687) );
  NAND2_X1 U10359 ( .A1(n10129), .A2(n8439), .ZN(n8835) );
  NAND2_X1 U10360 ( .A1(n9919), .A2(n8869), .ZN(n8834) );
  NAND2_X1 U10361 ( .A1(n8835), .A2(n8834), .ZN(n8837) );
  XNOR2_X1 U10362 ( .A(n8837), .B(n8836), .ZN(n9652) );
  NAND2_X1 U10363 ( .A1(n10129), .A2(n8869), .ZN(n8839) );
  NAND2_X1 U10364 ( .A1(n9919), .A2(n8874), .ZN(n8838) );
  NAND2_X1 U10365 ( .A1(n8839), .A2(n8838), .ZN(n8841) );
  NAND2_X1 U10366 ( .A1(n9652), .A2(n8841), .ZN(n8840) );
  NAND4_X1 U10367 ( .A1(n9655), .A2(n9689), .A3(n9687), .A4(n8840), .ZN(n8849)
         );
  INV_X1 U10368 ( .A(n9652), .ZN(n9654) );
  INV_X1 U10369 ( .A(n8841), .ZN(n9656) );
  NAND3_X1 U10370 ( .A1(n9687), .A2(n9654), .A3(n9656), .ZN(n8846) );
  INV_X1 U10371 ( .A(n8842), .ZN(n8845) );
  INV_X1 U10372 ( .A(n8843), .ZN(n8844) );
  NAND2_X1 U10373 ( .A1(n8845), .A2(n8844), .ZN(n9688) );
  NAND2_X1 U10374 ( .A1(n8846), .A2(n9688), .ZN(n8847) );
  NAND2_X1 U10375 ( .A1(n9689), .A2(n8847), .ZN(n8848) );
  INV_X1 U10376 ( .A(n8850), .ZN(n8851) );
  NOR2_X1 U10377 ( .A1(n8852), .A2(n8851), .ZN(n9763) );
  NAND2_X1 U10378 ( .A1(n10116), .A2(n8439), .ZN(n8854) );
  NAND2_X1 U10379 ( .A1(n9791), .A2(n8869), .ZN(n8853) );
  NAND2_X1 U10380 ( .A1(n8854), .A2(n8853), .ZN(n8855) );
  XNOR2_X1 U10381 ( .A(n8855), .B(n8872), .ZN(n8857) );
  AND2_X1 U10382 ( .A1(n9791), .A2(n8874), .ZN(n8856) );
  AOI21_X1 U10383 ( .B1(n10116), .B2(n8869), .A(n8856), .ZN(n8858) );
  XNOR2_X1 U10384 ( .A(n8857), .B(n8858), .ZN(n9762) );
  INV_X1 U10385 ( .A(n8857), .ZN(n8860) );
  INV_X1 U10386 ( .A(n8858), .ZN(n8859) );
  AND2_X1 U10387 ( .A1(n8860), .A2(n8859), .ZN(n9631) );
  NAND2_X1 U10388 ( .A1(n7150), .A2(n8439), .ZN(n8863) );
  OR2_X1 U10389 ( .A1(n9852), .A2(n4401), .ZN(n8862) );
  NAND2_X1 U10390 ( .A1(n8863), .A2(n8862), .ZN(n8864) );
  XNOR2_X1 U10391 ( .A(n8864), .B(n8872), .ZN(n8868) );
  NOR2_X1 U10392 ( .A1(n9852), .A2(n8865), .ZN(n8866) );
  AOI21_X1 U10393 ( .B1(n7150), .B2(n8869), .A(n8866), .ZN(n8867) );
  NAND2_X1 U10394 ( .A1(n8868), .A2(n8867), .ZN(n8883) );
  OAI21_X1 U10395 ( .B1(n8868), .B2(n8867), .A(n8883), .ZN(n9630) );
  NAND2_X1 U10396 ( .A1(n10107), .A2(n8439), .ZN(n8871) );
  NAND2_X1 U10397 ( .A1(n9790), .A2(n8869), .ZN(n8870) );
  NAND2_X1 U10398 ( .A1(n8871), .A2(n8870), .ZN(n8873) );
  XNOR2_X1 U10399 ( .A(n8873), .B(n8872), .ZN(n8876) );
  AOI22_X1 U10400 ( .A1(n10107), .A2(n8869), .B1(n8874), .B2(n9790), .ZN(n8875) );
  XNOR2_X1 U10401 ( .A(n8876), .B(n8875), .ZN(n8884) );
  INV_X1 U10402 ( .A(n8884), .ZN(n8877) );
  NAND2_X1 U10403 ( .A1(n8877), .A2(n9772), .ZN(n8878) );
  OAI21_X1 U10404 ( .B1(n9632), .B2(n5048), .A(n8879), .ZN(n8888) );
  OAI22_X1 U10405 ( .A1(n8942), .A2(n9782), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8880), .ZN(n8881) );
  AOI21_X1 U10406 ( .B1(n9780), .B2(n10092), .A(n8881), .ZN(n8882) );
  OAI21_X1 U10407 ( .B1(n9852), .B2(n9778), .A(n8882), .ZN(n8886) );
  NOR3_X1 U10408 ( .A1(n8884), .A2(n8883), .A3(n9760), .ZN(n8885) );
  AOI211_X1 U10409 ( .C1(n9784), .C2(n10107), .A(n8886), .B(n8885), .ZN(n8887)
         );
  NAND2_X1 U10410 ( .A1(n8888), .A2(n8887), .ZN(P1_U3218) );
  XNOR2_X1 U10411 ( .A(n8889), .B(n8892), .ZN(n10115) );
  INV_X1 U10412 ( .A(n9859), .ZN(n8890) );
  AOI21_X1 U10413 ( .B1(n7150), .B2(n8890), .A(n8938), .ZN(n10112) );
  AOI22_X1 U10414 ( .A1(n9637), .A2(n10059), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10020), .ZN(n8891) );
  OAI21_X1 U10415 ( .B1(n9639), .B2(n9999), .A(n8891), .ZN(n8898) );
  AOI21_X1 U10416 ( .B1(n8893), .B2(n8892), .A(n10044), .ZN(n8896) );
  OAI22_X1 U10417 ( .A1(n9634), .A2(n10040), .B1(n9872), .B2(n10071), .ZN(
        n8894) );
  AOI21_X1 U10418 ( .B1(n8896), .B2(n8895), .A(n8894), .ZN(n10114) );
  NOR2_X1 U10419 ( .A1(n10114), .A2(n10020), .ZN(n8897) );
  AOI211_X1 U10420 ( .C1(n10112), .C2(n10007), .A(n8898), .B(n8897), .ZN(n8899) );
  OAI21_X1 U10421 ( .B1(n10115), .B2(n10009), .A(n8899), .ZN(P1_U3264) );
  NOR2_X1 U10422 ( .A1(n10461), .A2(n9480), .ZN(n9201) );
  NOR2_X1 U10423 ( .A1(n8900), .A2(n10464), .ZN(n8901) );
  AOI211_X1 U10424 ( .C1(n10461), .C2(P2_REG2_REG_30__SCAN_IN), .A(n9201), .B(
        n8901), .ZN(n8902) );
  OAI21_X1 U10425 ( .B1(n8903), .B2(n10465), .A(n8902), .ZN(P2_U3266) );
  NAND2_X1 U10426 ( .A1(n8905), .A2(n8904), .ZN(n8906) );
  NAND2_X1 U10427 ( .A1(n4988), .A2(n7370), .ZN(n8909) );
  NAND2_X1 U10428 ( .A1(n8910), .A2(n8909), .ZN(n8914) );
  OR2_X1 U10429 ( .A1(n9485), .A2(n10461), .ZN(n8923) );
  AOI21_X1 U10430 ( .B1(n9483), .B2(n8916), .A(n8915), .ZN(n9484) );
  INV_X1 U10431 ( .A(n9483), .ZN(n8917) );
  NOR2_X1 U10432 ( .A1(n8917), .A2(n10464), .ZN(n8921) );
  OAI22_X1 U10433 ( .A1(n9457), .A2(n8919), .B1(n8918), .B2(n9290), .ZN(n8920)
         );
  AOI211_X1 U10434 ( .C1(n9484), .C2(n9464), .A(n8921), .B(n8920), .ZN(n8922)
         );
  OAI211_X1 U10435 ( .C1(n9486), .C2(n9411), .A(n8923), .B(n8922), .ZN(
        P2_U3267) );
  OAI22_X1 U10436 ( .A1(n9683), .A2(n8925), .B1(n8924), .B2(n9778), .ZN(n8926)
         );
  AOI21_X1 U10437 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n8927), .A(n8926), .ZN(
        n8933) );
  OAI21_X1 U10438 ( .B1(n8930), .B2(n8929), .A(n8928), .ZN(n8931) );
  NAND2_X1 U10439 ( .A1(n8931), .A2(n9772), .ZN(n8932) );
  OAI211_X1 U10440 ( .C1(n8934), .C2(n9771), .A(n8933), .B(n8932), .ZN(
        P1_U3220) );
  INV_X1 U10441 ( .A(n8938), .ZN(n8941) );
  INV_X1 U10442 ( .A(n8939), .ZN(n8940) );
  AOI21_X1 U10443 ( .B1(n10107), .B2(n8941), .A(n8940), .ZN(n10108) );
  INV_X1 U10444 ( .A(n8942), .ZN(n8943) );
  AOI22_X1 U10445 ( .A1(n8943), .A2(n10059), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n10020), .ZN(n8944) );
  OAI21_X1 U10446 ( .B1(n8945), .B2(n9999), .A(n8944), .ZN(n8951) );
  OAI21_X1 U10447 ( .B1(n8948), .B2(n8947), .A(n8946), .ZN(n8949) );
  OAI21_X1 U10448 ( .B1(n10111), .B2(n10009), .A(n8952), .ZN(P1_U3263) );
  INV_X1 U10449 ( .A(n8953), .ZN(n10233) );
  OAI222_X1 U10450 ( .A1(n8956), .A2(n10233), .B1(n8955), .B2(P2_U3152), .C1(
        n8954), .C2(n9624), .ZN(P2_U3328) );
  OAI222_X1 U10451 ( .A1(n10238), .A2(n8958), .B1(n4391), .B2(n8957), .C1(
        n5946), .C2(P1_U3084), .ZN(P1_U3332) );
  OAI222_X1 U10452 ( .A1(n9624), .A2(n8960), .B1(n9627), .B2(n8959), .C1(
        P2_U3152), .C2(n4384), .ZN(P2_U3336) );
  OAI211_X1 U10453 ( .C1(n8963), .C2(n8962), .A(n8961), .B(n9048), .ZN(n8968)
         );
  AOI22_X1 U10454 ( .A1(n9204), .A2(n9092), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n8967) );
  INV_X1 U10455 ( .A(n8964), .ZN(n9205) );
  AOI22_X1 U10456 ( .A1(n9103), .A2(n9203), .B1(n9205), .B2(n9102), .ZN(n8966)
         );
  NAND2_X1 U10457 ( .A1(n9493), .A2(n9108), .ZN(n8965) );
  NAND4_X1 U10458 ( .A1(n8968), .A2(n8967), .A3(n8966), .A4(n8965), .ZN(
        P2_U3216) );
  XNOR2_X1 U10459 ( .A(n9033), .B(n9032), .ZN(n8973) );
  OAI22_X1 U10460 ( .A1(n9106), .A2(n9265), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8969), .ZN(n8971) );
  OAI22_X1 U10461 ( .A1(n9072), .A2(n9264), .B1(n9095), .B2(n9269), .ZN(n8970)
         );
  AOI211_X1 U10462 ( .C1(n9515), .C2(n9108), .A(n8971), .B(n8970), .ZN(n8972)
         );
  OAI21_X1 U10463 ( .B1(n8973), .B2(n9110), .A(n8972), .ZN(P2_U3218) );
  OAI21_X1 U10464 ( .B1(n8976), .B2(n8975), .A(n8974), .ZN(n8977) );
  NAND2_X1 U10465 ( .A1(n8977), .A2(n9048), .ZN(n8982) );
  INV_X1 U10466 ( .A(n8978), .ZN(n8980) );
  OAI22_X1 U10467 ( .A1(n9072), .A2(n9026), .B1(n9095), .B2(n9335), .ZN(n8979)
         );
  AOI211_X1 U10468 ( .C1(n9092), .C2(n9328), .A(n8980), .B(n8979), .ZN(n8981)
         );
  OAI211_X1 U10469 ( .C1(n9338), .C2(n9023), .A(n8982), .B(n8981), .ZN(
        P2_U3221) );
  XNOR2_X1 U10470 ( .A(n8984), .B(n8983), .ZN(n8991) );
  OAI22_X1 U10471 ( .A1(n9106), .A2(n9264), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8985), .ZN(n8989) );
  INV_X1 U10472 ( .A(n9303), .ZN(n8986) );
  OAI22_X1 U10473 ( .A1(n9072), .A2(n8987), .B1(n9095), .B2(n8986), .ZN(n8988)
         );
  AOI211_X1 U10474 ( .C1(n9523), .C2(n9108), .A(n8989), .B(n8988), .ZN(n8990)
         );
  OAI21_X1 U10475 ( .B1(n8991), .B2(n9110), .A(n8990), .ZN(P2_U3225) );
  OAI21_X1 U10476 ( .B1(n8994), .B2(n8993), .A(n8992), .ZN(n8995) );
  NAND2_X1 U10477 ( .A1(n8995), .A2(n9048), .ZN(n9000) );
  AOI22_X1 U10478 ( .A1(n9092), .A2(n9115), .B1(P2_REG3_REG_12__SCAN_IN), .B2(
        P2_U3152), .ZN(n8999) );
  AOI22_X1 U10479 ( .A1(n9103), .A2(n9117), .B1(n9102), .B2(n8996), .ZN(n8998)
         );
  NAND2_X1 U10480 ( .A1(n9108), .A2(n6570), .ZN(n8997) );
  NAND4_X1 U10481 ( .A1(n9000), .A2(n8999), .A3(n8998), .A4(n8997), .ZN(
        P2_U3226) );
  INV_X1 U10482 ( .A(n9001), .ZN(n9085) );
  XNOR2_X1 U10483 ( .A(n9087), .B(n9085), .ZN(n9002) );
  XNOR2_X1 U10484 ( .A(n9084), .B(n9002), .ZN(n9008) );
  AOI22_X1 U10485 ( .A1(n9203), .A2(n9444), .B1(n9446), .B2(n9114), .ZN(n9230)
         );
  OAI22_X1 U10486 ( .A1(n9230), .A2(n9004), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9003), .ZN(n9005) );
  AOI21_X1 U10487 ( .B1(n9236), .B2(n9102), .A(n9005), .ZN(n9007) );
  NAND2_X1 U10488 ( .A1(n9237), .A2(n9108), .ZN(n9006) );
  OAI211_X1 U10489 ( .C1(n9008), .C2(n9110), .A(n9007), .B(n9006), .ZN(
        P2_U3227) );
  INV_X1 U10490 ( .A(n9392), .ZN(n9549) );
  NAND2_X1 U10491 ( .A1(n9010), .A2(n9009), .ZN(n9012) );
  OAI21_X1 U10492 ( .B1(n9010), .B2(n9009), .A(n9012), .ZN(n9100) );
  INV_X1 U10493 ( .A(n9011), .ZN(n9101) );
  NOR2_X1 U10494 ( .A1(n9100), .A2(n9101), .ZN(n9099) );
  INV_X1 U10495 ( .A(n9012), .ZN(n9014) );
  NOR3_X1 U10496 ( .A1(n9099), .A2(n9014), .A3(n9013), .ZN(n9017) );
  INV_X1 U10497 ( .A(n4392), .ZN(n9016) );
  OAI21_X1 U10498 ( .B1(n9017), .B2(n9016), .A(n9048), .ZN(n9022) );
  AND2_X1 U10499 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n9153) );
  INV_X1 U10500 ( .A(n9391), .ZN(n9018) );
  OAI22_X1 U10501 ( .A1(n9072), .A2(n9019), .B1(n9095), .B2(n9018), .ZN(n9020)
         );
  AOI211_X1 U10502 ( .C1(n9092), .C2(n9382), .A(n9153), .B(n9020), .ZN(n9021)
         );
  OAI211_X1 U10503 ( .C1(n9549), .C2(n9023), .A(n9022), .B(n9021), .ZN(
        P2_U3228) );
  XNOR2_X1 U10504 ( .A(n4511), .B(n9024), .ZN(n9030) );
  OAI22_X1 U10505 ( .A1(n9106), .A2(n9026), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9172), .ZN(n9028) );
  OAI22_X1 U10506 ( .A1(n9072), .A2(n9105), .B1(n9095), .B2(n9362), .ZN(n9027)
         );
  AOI211_X1 U10507 ( .C1(n9545), .C2(n9108), .A(n9028), .B(n9027), .ZN(n9029)
         );
  OAI21_X1 U10508 ( .B1(n9030), .B2(n9110), .A(n9029), .ZN(P2_U3230) );
  AOI21_X1 U10509 ( .B1(n9033), .B2(n9032), .A(n9031), .ZN(n9037) );
  XNOR2_X1 U10510 ( .A(n9035), .B(n9034), .ZN(n9036) );
  XNOR2_X1 U10511 ( .A(n9037), .B(n9036), .ZN(n9044) );
  OAI22_X1 U10512 ( .A1(n9106), .A2(n9039), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9038), .ZN(n9042) );
  INV_X1 U10513 ( .A(n9246), .ZN(n9040) );
  OAI22_X1 U10514 ( .A1(n9072), .A2(n9070), .B1(n9095), .B2(n9040), .ZN(n9041)
         );
  AOI211_X1 U10515 ( .C1(n9508), .C2(n9108), .A(n9042), .B(n9041), .ZN(n9043)
         );
  OAI21_X1 U10516 ( .B1(n9044), .B2(n9110), .A(n9043), .ZN(P2_U3231) );
  AOI22_X1 U10517 ( .A1(n9103), .A2(n9445), .B1(n9092), .B2(n9443), .ZN(n9053)
         );
  AOI22_X1 U10518 ( .A1(n9108), .A2(n9440), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3152), .ZN(n9052) );
  OAI21_X1 U10519 ( .B1(n9047), .B2(n9046), .A(n9045), .ZN(n9049) );
  NAND2_X1 U10520 ( .A1(n9049), .A2(n9048), .ZN(n9051) );
  NAND2_X1 U10521 ( .A1(n9102), .A2(n9449), .ZN(n9050) );
  NAND4_X1 U10522 ( .A1(n9053), .A2(n9052), .A3(n9051), .A4(n9050), .ZN(
        P2_U3232) );
  XNOR2_X1 U10523 ( .A(n9055), .B(n9054), .ZN(n9061) );
  OAI22_X1 U10524 ( .A1(n9106), .A2(n9071), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9056), .ZN(n9059) );
  INV_X1 U10525 ( .A(n9318), .ZN(n9057) );
  OAI22_X1 U10526 ( .A1(n9072), .A2(n9080), .B1(n9095), .B2(n9057), .ZN(n9058)
         );
  AOI211_X1 U10527 ( .C1(n9528), .C2(n9108), .A(n9059), .B(n9058), .ZN(n9060)
         );
  OAI21_X1 U10528 ( .B1(n9061), .B2(n9110), .A(n9060), .ZN(P2_U3235) );
  INV_X1 U10529 ( .A(n9062), .ZN(n9063) );
  NAND2_X1 U10530 ( .A1(n9064), .A2(n9063), .ZN(n9068) );
  XOR2_X1 U10531 ( .A(n9066), .B(n9065), .Z(n9067) );
  XNOR2_X1 U10532 ( .A(n9068), .B(n9067), .ZN(n9076) );
  OAI22_X1 U10533 ( .A1(n9106), .A2(n9070), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9069), .ZN(n9074) );
  OAI22_X1 U10534 ( .A1(n9072), .A2(n9071), .B1(n9095), .B2(n9289), .ZN(n9073)
         );
  AOI211_X1 U10535 ( .C1(n9520), .C2(n9108), .A(n9074), .B(n9073), .ZN(n9075)
         );
  OAI21_X1 U10536 ( .B1(n9076), .B2(n9110), .A(n9075), .ZN(P2_U3237) );
  XNOR2_X1 U10537 ( .A(n9078), .B(n9077), .ZN(n9083) );
  AOI22_X1 U10538 ( .A1(n9103), .A2(n9382), .B1(n9102), .B2(n9349), .ZN(n9079)
         );
  NAND2_X1 U10539 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9189) );
  OAI211_X1 U10540 ( .C1(n9106), .C2(n9080), .A(n9079), .B(n9189), .ZN(n9081)
         );
  AOI21_X1 U10541 ( .B1(n9539), .B2(n9108), .A(n9081), .ZN(n9082) );
  OAI21_X1 U10542 ( .B1(n9083), .B2(n9110), .A(n9082), .ZN(P2_U3240) );
  OAI21_X1 U10543 ( .B1(n9087), .B2(n9084), .A(n9086), .ZN(n9091) );
  NAND2_X1 U10544 ( .A1(n9089), .A2(n9088), .ZN(n9090) );
  XNOR2_X1 U10545 ( .A(n9091), .B(n9090), .ZN(n9098) );
  AOI22_X1 U10546 ( .A1(n9220), .A2(n9092), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n9094) );
  NAND2_X1 U10547 ( .A1(n9103), .A2(n9252), .ZN(n9093) );
  OAI211_X1 U10548 ( .C1(n9224), .C2(n9095), .A(n9094), .B(n9093), .ZN(n9096)
         );
  AOI21_X1 U10549 ( .B1(n9498), .B2(n9108), .A(n9096), .ZN(n9097) );
  OAI21_X1 U10550 ( .B1(n9098), .B2(n9110), .A(n9097), .ZN(P2_U3242) );
  AOI21_X1 U10551 ( .B1(n9101), .B2(n9100), .A(n9099), .ZN(n9111) );
  AOI22_X1 U10552 ( .A1(n9103), .A2(n9400), .B1(n9102), .B2(n9406), .ZN(n9104)
         );
  NAND2_X1 U10553 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9143) );
  OAI211_X1 U10554 ( .C1(n9106), .C2(n9105), .A(n9104), .B(n9143), .ZN(n9107)
         );
  AOI21_X1 U10555 ( .B1(n9556), .B2(n9108), .A(n9107), .ZN(n9109) );
  OAI21_X1 U10556 ( .B1(n9111), .B2(n9110), .A(n9109), .ZN(P2_U3243) );
  MUX2_X1 U10557 ( .A(n9112), .B(P2_DATAO_REG_30__SCAN_IN), .S(n9125), .Z(
        P2_U3582) );
  MUX2_X1 U10558 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n9113), .S(P2_U3966), .Z(
        P2_U3581) );
  MUX2_X1 U10559 ( .A(n9204), .B(P2_DATAO_REG_28__SCAN_IN), .S(n9125), .Z(
        P2_U3580) );
  MUX2_X1 U10560 ( .A(n9220), .B(P2_DATAO_REG_27__SCAN_IN), .S(n9125), .Z(
        P2_U3579) );
  MUX2_X1 U10561 ( .A(n9203), .B(P2_DATAO_REG_26__SCAN_IN), .S(n9125), .Z(
        P2_U3578) );
  MUX2_X1 U10562 ( .A(n9252), .B(P2_DATAO_REG_25__SCAN_IN), .S(n9125), .Z(
        P2_U3577) );
  MUX2_X1 U10563 ( .A(n9114), .B(P2_DATAO_REG_24__SCAN_IN), .S(n9125), .Z(
        P2_U3576) );
  MUX2_X1 U10564 ( .A(n9282), .B(P2_DATAO_REG_23__SCAN_IN), .S(n9125), .Z(
        P2_U3575) );
  MUX2_X1 U10565 ( .A(n4390), .B(P2_DATAO_REG_22__SCAN_IN), .S(n9125), .Z(
        P2_U3574) );
  MUX2_X1 U10566 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n9314), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U10567 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n9328), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U10568 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n9346), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U10569 ( .A(n9359), .B(P2_DATAO_REG_18__SCAN_IN), .S(n9125), .Z(
        P2_U3570) );
  MUX2_X1 U10570 ( .A(n9382), .B(P2_DATAO_REG_17__SCAN_IN), .S(n9125), .Z(
        P2_U3569) );
  MUX2_X1 U10571 ( .A(n9401), .B(P2_DATAO_REG_16__SCAN_IN), .S(n9125), .Z(
        P2_U3568) );
  MUX2_X1 U10572 ( .A(n9381), .B(P2_DATAO_REG_15__SCAN_IN), .S(n9125), .Z(
        P2_U3567) );
  MUX2_X1 U10573 ( .A(n9400), .B(P2_DATAO_REG_14__SCAN_IN), .S(n9125), .Z(
        P2_U3566) );
  MUX2_X1 U10574 ( .A(n9115), .B(P2_DATAO_REG_13__SCAN_IN), .S(n9125), .Z(
        P2_U3565) );
  MUX2_X1 U10575 ( .A(n9116), .B(P2_DATAO_REG_12__SCAN_IN), .S(n9125), .Z(
        P2_U3564) );
  MUX2_X1 U10576 ( .A(n9117), .B(P2_DATAO_REG_11__SCAN_IN), .S(n9125), .Z(
        P2_U3563) );
  MUX2_X1 U10577 ( .A(n9118), .B(P2_DATAO_REG_10__SCAN_IN), .S(n9125), .Z(
        P2_U3562) );
  MUX2_X1 U10578 ( .A(n9119), .B(P2_DATAO_REG_9__SCAN_IN), .S(n9125), .Z(
        P2_U3561) );
  MUX2_X1 U10579 ( .A(n9120), .B(P2_DATAO_REG_8__SCAN_IN), .S(n9125), .Z(
        P2_U3560) );
  MUX2_X1 U10580 ( .A(n9121), .B(P2_DATAO_REG_7__SCAN_IN), .S(n9125), .Z(
        P2_U3559) );
  MUX2_X1 U10581 ( .A(n9122), .B(P2_DATAO_REG_6__SCAN_IN), .S(n9125), .Z(
        P2_U3558) );
  MUX2_X1 U10582 ( .A(n9443), .B(P2_DATAO_REG_5__SCAN_IN), .S(n9125), .Z(
        P2_U3557) );
  MUX2_X1 U10583 ( .A(n9123), .B(P2_DATAO_REG_4__SCAN_IN), .S(n9125), .Z(
        P2_U3556) );
  MUX2_X1 U10584 ( .A(n9445), .B(P2_DATAO_REG_3__SCAN_IN), .S(n9125), .Z(
        P2_U3555) );
  MUX2_X1 U10585 ( .A(n4389), .B(P2_DATAO_REG_2__SCAN_IN), .S(n9125), .Z(
        P2_U3554) );
  MUX2_X1 U10586 ( .A(n9124), .B(P2_DATAO_REG_1__SCAN_IN), .S(n9125), .Z(
        P2_U3553) );
  MUX2_X1 U10587 ( .A(n6592), .B(P2_DATAO_REG_0__SCAN_IN), .S(n9125), .Z(
        P2_U3552) );
  XOR2_X1 U10588 ( .A(n9127), .B(n9126), .Z(n9137) );
  OAI21_X1 U10589 ( .B1(n9130), .B2(n9129), .A(n9128), .ZN(n9135) );
  AOI21_X1 U10590 ( .B1(n9174), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n9131), .ZN(
        n9132) );
  OAI21_X1 U10591 ( .B1(n9178), .B2(n9133), .A(n9132), .ZN(n9134) );
  AOI21_X1 U10592 ( .B1(n9135), .B2(n9169), .A(n9134), .ZN(n9136) );
  OAI21_X1 U10593 ( .B1(n9137), .B2(n9184), .A(n9136), .ZN(P2_U3259) );
  XNOR2_X1 U10594 ( .A(n9138), .B(P2_REG1_REG_15__SCAN_IN), .ZN(n9149) );
  OAI21_X1 U10595 ( .B1(n9141), .B2(n9140), .A(n9139), .ZN(n9142) );
  NAND2_X1 U10596 ( .A1(n9142), .A2(n9163), .ZN(n9148) );
  INV_X1 U10597 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n9144) );
  OAI21_X1 U10598 ( .B1(n9190), .B2(n9144), .A(n9143), .ZN(n9145) );
  AOI21_X1 U10599 ( .B1(n9193), .B2(n9146), .A(n9145), .ZN(n9147) );
  OAI211_X1 U10600 ( .C1(n9196), .C2(n9149), .A(n9148), .B(n9147), .ZN(
        P2_U3260) );
  AOI21_X1 U10601 ( .B1(n9152), .B2(n9151), .A(n9150), .ZN(n9162) );
  AOI21_X1 U10602 ( .B1(n9174), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n9153), .ZN(
        n9154) );
  OAI21_X1 U10603 ( .B1(n9178), .B2(n9155), .A(n9154), .ZN(n9161) );
  AOI21_X1 U10604 ( .B1(n9158), .B2(n9157), .A(n9156), .ZN(n9159) );
  NOR2_X1 U10605 ( .A1(n9159), .A2(n9196), .ZN(n9160) );
  AOI211_X1 U10606 ( .C1(n9163), .C2(n9162), .A(n9161), .B(n9160), .ZN(n9164)
         );
  INV_X1 U10607 ( .A(n9164), .ZN(P2_U3261) );
  AOI211_X1 U10608 ( .C1(n9167), .C2(n9166), .A(n9165), .B(n9184), .ZN(n9180)
         );
  OAI211_X1 U10609 ( .C1(n9171), .C2(n9170), .A(n9169), .B(n9168), .ZN(n9176)
         );
  NOR2_X1 U10610 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9172), .ZN(n9173) );
  AOI21_X1 U10611 ( .B1(n9174), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n9173), .ZN(
        n9175) );
  OAI211_X1 U10612 ( .C1(n9178), .C2(n9177), .A(n9176), .B(n9175), .ZN(n9179)
         );
  OR2_X1 U10613 ( .A1(n9180), .A2(n9179), .ZN(P2_U3262) );
  AOI21_X1 U10614 ( .B1(n9183), .B2(n9182), .A(n9181), .ZN(n9197) );
  AOI211_X1 U10615 ( .C1(n9187), .C2(n9186), .A(n9185), .B(n9184), .ZN(n9188)
         );
  INV_X1 U10616 ( .A(n9188), .ZN(n9195) );
  OAI21_X1 U10617 ( .B1(n9190), .B2(n10568), .A(n9189), .ZN(n9191) );
  AOI21_X1 U10618 ( .B1(n9193), .B2(n9192), .A(n9191), .ZN(n9194) );
  OAI211_X1 U10619 ( .C1(n9197), .C2(n9196), .A(n9195), .B(n9194), .ZN(
        P2_U3263) );
  XNOR2_X1 U10620 ( .A(n9198), .B(n9478), .ZN(n9481) );
  NOR2_X1 U10621 ( .A1(n9199), .A2(n10464), .ZN(n9200) );
  AOI211_X1 U10622 ( .C1(n10461), .C2(P2_REG2_REG_31__SCAN_IN), .A(n9201), .B(
        n9200), .ZN(n9202) );
  OAI21_X1 U10623 ( .B1(n9481), .B2(n10465), .A(n9202), .ZN(P2_U3265) );
  AOI211_X1 U10624 ( .C1(n9493), .C2(n4409), .A(n10508), .B(n4859), .ZN(n9492)
         );
  AOI22_X1 U10625 ( .A1(n9205), .A2(n10462), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n10470), .ZN(n9206) );
  OAI21_X1 U10626 ( .B1(n9207), .B2(n10464), .A(n9206), .ZN(n9212) );
  OAI21_X1 U10627 ( .B1(n9210), .B2(n9209), .A(n9208), .ZN(n9211) );
  OAI21_X1 U10628 ( .B1(n9215), .B2(n9214), .A(n9213), .ZN(n9216) );
  INV_X1 U10629 ( .A(n9216), .ZN(n9501) );
  OAI21_X1 U10630 ( .B1(n9219), .B2(n9218), .A(n9217), .ZN(n9221) );
  AOI222_X1 U10631 ( .A1(n9385), .A2(n9221), .B1(n9220), .B2(n9444), .C1(n9252), .C2(n9446), .ZN(n9500) );
  AOI21_X1 U10632 ( .B1(n9235), .B2(n9498), .A(n10508), .ZN(n9222) );
  AND2_X1 U10633 ( .A1(n9222), .A2(n4409), .ZN(n9497) );
  NAND2_X1 U10634 ( .A1(n9497), .A2(n4944), .ZN(n9223) );
  OAI211_X1 U10635 ( .C1(n9290), .C2(n9224), .A(n4400), .B(n9223), .ZN(n9225)
         );
  NAND2_X1 U10636 ( .A1(n9225), .A2(n9457), .ZN(n9227) );
  AOI22_X1 U10637 ( .A1(n9498), .A2(n9469), .B1(n10461), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n9226) );
  OAI211_X1 U10638 ( .C1(n9501), .C2(n9411), .A(n9227), .B(n9226), .ZN(
        P2_U3270) );
  XNOR2_X1 U10639 ( .A(n9229), .B(n9228), .ZN(n9231) );
  OAI21_X1 U10640 ( .B1(n9231), .B2(n9263), .A(n9230), .ZN(n9504) );
  INV_X1 U10641 ( .A(n9504), .ZN(n9242) );
  OAI21_X1 U10642 ( .B1(n9233), .B2(n4994), .A(n9232), .ZN(n9506) );
  OAI211_X1 U10643 ( .C1(n9503), .C2(n9234), .A(n9235), .B(n9589), .ZN(n9502)
         );
  AOI22_X1 U10644 ( .A1(n10470), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n9236), 
        .B2(n10462), .ZN(n9239) );
  NAND2_X1 U10645 ( .A1(n9237), .A2(n9469), .ZN(n9238) );
  OAI211_X1 U10646 ( .C1(n9502), .C2(n9334), .A(n9239), .B(n9238), .ZN(n9240)
         );
  AOI21_X1 U10647 ( .B1(n9506), .B2(n10467), .A(n9240), .ZN(n9241) );
  OAI21_X1 U10648 ( .B1(n9242), .B2(n10470), .A(n9241), .ZN(P2_U3271) );
  XOR2_X1 U10649 ( .A(n9243), .B(n9250), .Z(n9512) );
  INV_X1 U10650 ( .A(n9244), .ZN(n9245) );
  AOI21_X1 U10651 ( .B1(n9508), .B2(n9245), .A(n9234), .ZN(n9509) );
  AOI22_X1 U10652 ( .A1(n10470), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n9246), 
        .B2(n10462), .ZN(n9247) );
  OAI21_X1 U10653 ( .B1(n9248), .B2(n10464), .A(n9247), .ZN(n9256) );
  OAI211_X1 U10654 ( .C1(n9251), .C2(n9250), .A(n9249), .B(n10460), .ZN(n9254)
         );
  AOI22_X1 U10655 ( .A1(n9252), .A2(n9444), .B1(n9446), .B2(n9282), .ZN(n9253)
         );
  AND2_X1 U10656 ( .A1(n9254), .A2(n9253), .ZN(n9511) );
  NOR2_X1 U10657 ( .A1(n9511), .A2(n10470), .ZN(n9255) );
  AOI211_X1 U10658 ( .C1(n9509), .C2(n9464), .A(n9256), .B(n9255), .ZN(n9257)
         );
  OAI21_X1 U10659 ( .B1(n9512), .B2(n9411), .A(n9257), .ZN(P2_U3272) );
  OAI21_X1 U10660 ( .B1(n9259), .B2(n9261), .A(n9258), .ZN(n9517) );
  AOI21_X1 U10661 ( .B1(n9261), .B2(n9260), .A(n4475), .ZN(n9262) );
  OAI222_X1 U10662 ( .A1(n9419), .A2(n9265), .B1(n9418), .B2(n9264), .C1(n9263), .C2(n9262), .ZN(n9513) );
  OAI21_X1 U10663 ( .B1(n9287), .B2(n9266), .A(n9589), .ZN(n9267) );
  NOR2_X1 U10664 ( .A1(n9267), .A2(n9244), .ZN(n9514) );
  NAND2_X1 U10665 ( .A1(n9514), .A2(n9472), .ZN(n9272) );
  NAND2_X1 U10666 ( .A1(n10470), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n9268) );
  OAI21_X1 U10667 ( .B1(n9290), .B2(n9269), .A(n9268), .ZN(n9270) );
  AOI21_X1 U10668 ( .B1(n9515), .B2(n9469), .A(n9270), .ZN(n9271) );
  NAND2_X1 U10669 ( .A1(n9272), .A2(n9271), .ZN(n9273) );
  AOI21_X1 U10670 ( .B1(n9513), .B2(n9457), .A(n9273), .ZN(n9274) );
  OAI21_X1 U10671 ( .B1(n9411), .B2(n9517), .A(n9274), .ZN(P2_U3273) );
  XNOR2_X1 U10672 ( .A(n9276), .B(n9275), .ZN(n9522) );
  INV_X1 U10673 ( .A(n9278), .ZN(n9297) );
  NOR3_X1 U10674 ( .A1(n9310), .A2(n9297), .A3(n9306), .ZN(n9296) );
  OAI21_X1 U10675 ( .B1(n9296), .B2(n9279), .A(n6549), .ZN(n9281) );
  NAND3_X1 U10676 ( .A1(n9281), .A2(n9280), .A3(n10460), .ZN(n9284) );
  AOI22_X1 U10677 ( .A1(n9282), .A2(n9444), .B1(n9446), .B2(n9314), .ZN(n9283)
         );
  NAND2_X1 U10678 ( .A1(n9284), .A2(n9283), .ZN(n9518) );
  NAND2_X1 U10679 ( .A1(n9302), .A2(n9520), .ZN(n9285) );
  NAND2_X1 U10680 ( .A1(n9285), .A2(n9589), .ZN(n9286) );
  NOR2_X1 U10681 ( .A1(n9287), .A2(n9286), .ZN(n9519) );
  NAND2_X1 U10682 ( .A1(n9519), .A2(n9472), .ZN(n9293) );
  NAND2_X1 U10683 ( .A1(n10470), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n9288) );
  OAI21_X1 U10684 ( .B1(n9290), .B2(n9289), .A(n9288), .ZN(n9291) );
  AOI21_X1 U10685 ( .B1(n9520), .B2(n9469), .A(n9291), .ZN(n9292) );
  NAND2_X1 U10686 ( .A1(n9293), .A2(n9292), .ZN(n9294) );
  AOI21_X1 U10687 ( .B1(n9518), .B2(n9457), .A(n9294), .ZN(n9295) );
  OAI21_X1 U10688 ( .B1(n9411), .B2(n9522), .A(n9295), .ZN(P2_U3274) );
  INV_X1 U10689 ( .A(n9296), .ZN(n9299) );
  OAI21_X1 U10690 ( .B1(n9310), .B2(n9297), .A(n9306), .ZN(n9298) );
  NAND2_X1 U10691 ( .A1(n9299), .A2(n9298), .ZN(n9300) );
  AOI222_X1 U10692 ( .A1(n9385), .A2(n9300), .B1(n4390), .B2(n9444), .C1(n9328), .C2(n9446), .ZN(n9526) );
  AOI21_X1 U10693 ( .B1(n9523), .B2(n9317), .A(n4854), .ZN(n9524) );
  AOI22_X1 U10694 ( .A1(n10470), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9303), 
        .B2(n10462), .ZN(n9304) );
  OAI21_X1 U10695 ( .B1(n6573), .B2(n10464), .A(n9304), .ZN(n9308) );
  XNOR2_X1 U10696 ( .A(n9305), .B(n9306), .ZN(n9527) );
  NOR2_X1 U10697 ( .A1(n9527), .A2(n9411), .ZN(n9307) );
  AOI211_X1 U10698 ( .C1(n9524), .C2(n9464), .A(n9308), .B(n9307), .ZN(n9309)
         );
  OAI21_X1 U10699 ( .B1(n9526), .B2(n10470), .A(n9309), .ZN(P2_U3275) );
  INV_X1 U10700 ( .A(n9310), .ZN(n9313) );
  OAI21_X1 U10701 ( .B1(n9326), .B2(n9311), .A(n9321), .ZN(n9312) );
  NAND3_X1 U10702 ( .A1(n9313), .A2(n10460), .A3(n9312), .ZN(n9316) );
  AOI22_X1 U10703 ( .A1(n9314), .A2(n9444), .B1(n9446), .B2(n9346), .ZN(n9315)
         );
  AOI21_X1 U10704 ( .B1(n9528), .B2(n9331), .A(n9301), .ZN(n9529) );
  AOI22_X1 U10705 ( .A1(n10461), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9318), 
        .B2(n10462), .ZN(n9319) );
  OAI21_X1 U10706 ( .B1(n4856), .B2(n10464), .A(n9319), .ZN(n9320) );
  AOI21_X1 U10707 ( .B1(n9529), .B2(n9464), .A(n9320), .ZN(n9325) );
  OR2_X1 U10708 ( .A1(n9322), .A2(n9321), .ZN(n9530) );
  NAND3_X1 U10709 ( .A1(n9530), .A2(n10467), .A3(n9323), .ZN(n9324) );
  OAI211_X1 U10710 ( .C1(n9533), .C2(n10461), .A(n9325), .B(n9324), .ZN(
        P2_U3276) );
  INV_X1 U10711 ( .A(n9326), .ZN(n9327) );
  OAI21_X1 U10712 ( .B1(n9340), .B2(n9277), .A(n9327), .ZN(n9329) );
  AOI222_X1 U10713 ( .A1(n9385), .A2(n9329), .B1(n9328), .B2(n9444), .C1(n9359), .C2(n9446), .ZN(n9537) );
  INV_X1 U10714 ( .A(n9330), .ZN(n9333) );
  INV_X1 U10715 ( .A(n9331), .ZN(n9332) );
  AOI211_X1 U10716 ( .C1(n9535), .C2(n9333), .A(n10508), .B(n9332), .ZN(n9534)
         );
  INV_X1 U10717 ( .A(n9334), .ZN(n9374) );
  INV_X1 U10718 ( .A(n9335), .ZN(n9336) );
  AOI22_X1 U10719 ( .A1(n10470), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n9336), 
        .B2(n10462), .ZN(n9337) );
  OAI21_X1 U10720 ( .B1(n9338), .B2(n10464), .A(n9337), .ZN(n9342) );
  XOR2_X1 U10721 ( .A(n9339), .B(n9340), .Z(n9538) );
  NOR2_X1 U10722 ( .A1(n9538), .A2(n9411), .ZN(n9341) );
  AOI211_X1 U10723 ( .C1(n9534), .C2(n9374), .A(n9342), .B(n9341), .ZN(n9343)
         );
  OAI21_X1 U10724 ( .B1(n9537), .B2(n10470), .A(n9343), .ZN(P2_U3277) );
  OAI21_X1 U10725 ( .B1(n9352), .B2(n9345), .A(n9344), .ZN(n9347) );
  AOI222_X1 U10726 ( .A1(n9385), .A2(n9347), .B1(n9346), .B2(n9444), .C1(n9382), .C2(n9446), .ZN(n9542) );
  INV_X1 U10727 ( .A(n9361), .ZN(n9348) );
  AOI21_X1 U10728 ( .B1(n9539), .B2(n9348), .A(n9330), .ZN(n9540) );
  AOI22_X1 U10729 ( .A1(n10470), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9349), 
        .B2(n10462), .ZN(n9350) );
  OAI21_X1 U10730 ( .B1(n9351), .B2(n10464), .A(n9350), .ZN(n9355) );
  XNOR2_X1 U10731 ( .A(n9353), .B(n9352), .ZN(n9543) );
  NOR2_X1 U10732 ( .A1(n9543), .A2(n9411), .ZN(n9354) );
  AOI211_X1 U10733 ( .C1(n9540), .C2(n9464), .A(n9355), .B(n9354), .ZN(n9356)
         );
  OAI21_X1 U10734 ( .B1(n9542), .B2(n10470), .A(n9356), .ZN(P2_U3278) );
  XNOR2_X1 U10735 ( .A(n9358), .B(n9357), .ZN(n9360) );
  AOI222_X1 U10736 ( .A1(n9385), .A2(n9360), .B1(n9359), .B2(n9444), .C1(n9401), .C2(n9446), .ZN(n9547) );
  AOI211_X1 U10737 ( .C1(n9545), .C2(n9390), .A(n10508), .B(n9361), .ZN(n9544)
         );
  INV_X1 U10738 ( .A(n9545), .ZN(n9365) );
  INV_X1 U10739 ( .A(n9362), .ZN(n9363) );
  AOI22_X1 U10740 ( .A1(n10470), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n9363), 
        .B2(n10462), .ZN(n9364) );
  OAI21_X1 U10741 ( .B1(n9365), .B2(n10464), .A(n9364), .ZN(n9373) );
  NAND2_X1 U10742 ( .A1(n9366), .A2(n9367), .ZN(n9370) );
  INV_X1 U10743 ( .A(n9368), .ZN(n9369) );
  AOI21_X1 U10744 ( .B1(n9371), .B2(n9370), .A(n9369), .ZN(n9548) );
  NOR2_X1 U10745 ( .A1(n9548), .A2(n9411), .ZN(n9372) );
  AOI211_X1 U10746 ( .C1(n9544), .C2(n9374), .A(n9373), .B(n9372), .ZN(n9375)
         );
  OAI21_X1 U10747 ( .B1(n9547), .B2(n10470), .A(n9375), .ZN(P2_U3279) );
  INV_X1 U10748 ( .A(n9378), .ZN(n9377) );
  XNOR2_X1 U10749 ( .A(n9376), .B(n9377), .ZN(n9386) );
  OR2_X1 U10750 ( .A1(n9379), .A2(n9378), .ZN(n9380) );
  NAND2_X1 U10751 ( .A1(n9366), .A2(n9380), .ZN(n9387) );
  AOI22_X1 U10752 ( .A1(n9382), .A2(n9444), .B1(n9446), .B2(n9381), .ZN(n9383)
         );
  OAI21_X1 U10753 ( .B1(n9387), .B2(n9425), .A(n9383), .ZN(n9384) );
  AOI21_X1 U10754 ( .B1(n9386), .B2(n9385), .A(n9384), .ZN(n9555) );
  INV_X1 U10755 ( .A(n9387), .ZN(n9553) );
  NAND2_X1 U10756 ( .A1(n9388), .A2(n9392), .ZN(n9389) );
  NAND2_X1 U10757 ( .A1(n9390), .A2(n9389), .ZN(n9550) );
  AOI22_X1 U10758 ( .A1(n10461), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n9391), 
        .B2(n10462), .ZN(n9394) );
  NAND2_X1 U10759 ( .A1(n9392), .A2(n9469), .ZN(n9393) );
  OAI211_X1 U10760 ( .C1(n9550), .C2(n10465), .A(n9394), .B(n9393), .ZN(n9395)
         );
  AOI21_X1 U10761 ( .B1(n9553), .B2(n9396), .A(n9395), .ZN(n9397) );
  OAI21_X1 U10762 ( .B1(n9555), .B2(n10470), .A(n9397), .ZN(P2_U3280) );
  OAI211_X1 U10763 ( .C1(n9409), .C2(n9398), .A(n9399), .B(n10460), .ZN(n9403)
         );
  AOI22_X1 U10764 ( .A1(n9401), .A2(n9444), .B1(n9446), .B2(n9400), .ZN(n9402)
         );
  AND2_X1 U10765 ( .A1(n9403), .A2(n9402), .ZN(n9559) );
  INV_X1 U10766 ( .A(n8671), .ZN(n9405) );
  INV_X1 U10767 ( .A(n9388), .ZN(n9404) );
  AOI21_X1 U10768 ( .B1(n9556), .B2(n9405), .A(n9404), .ZN(n9557) );
  AOI22_X1 U10769 ( .A1(n10461), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n9406), 
        .B2(n10462), .ZN(n9407) );
  OAI21_X1 U10770 ( .B1(n9408), .B2(n10464), .A(n9407), .ZN(n9413) );
  XNOR2_X1 U10771 ( .A(n9410), .B(n9409), .ZN(n9560) );
  NOR2_X1 U10772 ( .A1(n9560), .A2(n9411), .ZN(n9412) );
  AOI211_X1 U10773 ( .C1(n9557), .C2(n9464), .A(n9413), .B(n9412), .ZN(n9414)
         );
  OAI21_X1 U10774 ( .B1(n9559), .B2(n10470), .A(n9414), .ZN(P2_U3281) );
  OAI21_X1 U10775 ( .B1(n9424), .B2(n9416), .A(n9415), .ZN(n9428) );
  OAI22_X1 U10776 ( .A1(n9420), .A2(n9419), .B1(n9418), .B2(n9417), .ZN(n9427)
         );
  NOR2_X1 U10777 ( .A1(n9422), .A2(n9421), .ZN(n9423) );
  XOR2_X1 U10778 ( .A(n9424), .B(n9423), .Z(n9569) );
  NOR2_X1 U10779 ( .A1(n9569), .A2(n9425), .ZN(n9426) );
  AOI211_X1 U10780 ( .C1(n10460), .C2(n9428), .A(n9427), .B(n9426), .ZN(n9568)
         );
  AOI21_X1 U10781 ( .B1(n9565), .B2(n9430), .A(n9429), .ZN(n9566) );
  AOI22_X1 U10782 ( .A1(n10461), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n9431), 
        .B2(n10462), .ZN(n9432) );
  OAI21_X1 U10783 ( .B1(n10464), .B2(n9433), .A(n9432), .ZN(n9436) );
  NOR2_X1 U10784 ( .A1(n9569), .A2(n9434), .ZN(n9435) );
  AOI211_X1 U10785 ( .C1(n9566), .C2(n9464), .A(n9436), .B(n9435), .ZN(n9437)
         );
  OAI21_X1 U10786 ( .B1(n9568), .B2(n10461), .A(n9437), .ZN(P2_U3283) );
  INV_X1 U10787 ( .A(n7780), .ZN(n9439) );
  AOI21_X1 U10788 ( .B1(n9440), .B2(n9439), .A(n6568), .ZN(n10493) );
  AOI22_X1 U10789 ( .A1(n9469), .A2(n9440), .B1(n9464), .B2(n10493), .ZN(n9456) );
  OAI211_X1 U10790 ( .C1(n9442), .C2(n6528), .A(n9441), .B(n10460), .ZN(n9448)
         );
  AOI22_X1 U10791 ( .A1(n9446), .A2(n9445), .B1(n9444), .B2(n9443), .ZN(n9447)
         );
  NAND2_X1 U10792 ( .A1(n9448), .A2(n9447), .ZN(n10496) );
  AOI22_X1 U10793 ( .A1(n9457), .A2(n10496), .B1(n9449), .B2(n10462), .ZN(
        n9455) );
  NAND2_X1 U10794 ( .A1(n10470), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9454) );
  OAI21_X1 U10795 ( .B1(n9452), .B2(n9451), .A(n9450), .ZN(n10498) );
  NAND2_X1 U10796 ( .A1(n10467), .A2(n10498), .ZN(n9453) );
  NAND4_X1 U10797 ( .A1(n9456), .A2(n9455), .A3(n9454), .A4(n9453), .ZN(
        P2_U3292) );
  MUX2_X1 U10798 ( .A(n9459), .B(n9458), .S(n9457), .Z(n9467) );
  AOI22_X1 U10799 ( .A1(n10467), .A2(n9461), .B1(n9469), .B2(n9460), .ZN(n9466) );
  AOI22_X1 U10800 ( .A1(n9464), .A2(n9463), .B1(n10462), .B2(n9462), .ZN(n9465) );
  NAND3_X1 U10801 ( .A1(n9467), .A2(n9466), .A3(n9465), .ZN(P2_U3293) );
  AOI22_X1 U10802 ( .A1(n10467), .A2(n9470), .B1(n9469), .B2(n9468), .ZN(n9477) );
  AOI22_X1 U10803 ( .A1(n9472), .A2(n9471), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n10462), .ZN(n9476) );
  NOR2_X1 U10804 ( .A1(n9473), .A2(n10461), .ZN(n9474) );
  AOI21_X1 U10805 ( .B1(n10461), .B2(P2_REG2_REG_1__SCAN_IN), .A(n9474), .ZN(
        n9475) );
  NAND3_X1 U10806 ( .A1(n9477), .A2(n9476), .A3(n9475), .ZN(P2_U3295) );
  NAND2_X1 U10807 ( .A1(n9478), .A2(n9588), .ZN(n9479) );
  OAI211_X1 U10808 ( .C1(n9481), .C2(n10508), .A(n9480), .B(n9479), .ZN(n9595)
         );
  MUX2_X1 U10809 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9595), .S(n10526), .Z(
        P2_U3551) );
  MUX2_X1 U10810 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9482), .S(n10526), .Z(
        P2_U3550) );
  AOI21_X1 U10811 ( .B1(n9588), .B2(n9488), .A(n9487), .ZN(n9489) );
  OAI211_X1 U10812 ( .C1(n9579), .C2(n9491), .A(n9490), .B(n9489), .ZN(n9597)
         );
  MUX2_X1 U10813 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9597), .S(n10526), .Z(
        P2_U3548) );
  AOI21_X1 U10814 ( .B1(n9588), .B2(n9493), .A(n9492), .ZN(n9494) );
  OAI211_X1 U10815 ( .C1(n9579), .C2(n9496), .A(n9495), .B(n9494), .ZN(n9598)
         );
  MUX2_X1 U10816 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9598), .S(n10526), .Z(
        P2_U3547) );
  AOI21_X1 U10817 ( .B1(n9588), .B2(n9498), .A(n9497), .ZN(n9499) );
  OAI211_X1 U10818 ( .C1(n9579), .C2(n9501), .A(n4400), .B(n9499), .ZN(n9599)
         );
  MUX2_X1 U10819 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9599), .S(n10526), .Z(
        P2_U3546) );
  OAI21_X1 U10820 ( .B1(n9503), .B2(n10507), .A(n9502), .ZN(n9505) );
  AOI211_X1 U10821 ( .C1(n10512), .C2(n9506), .A(n9505), .B(n9504), .ZN(n9507)
         );
  INV_X1 U10822 ( .A(n9507), .ZN(n9600) );
  MUX2_X1 U10823 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9600), .S(n10526), .Z(
        P2_U3545) );
  AOI22_X1 U10824 ( .A1(n9509), .A2(n9589), .B1(n9588), .B2(n9508), .ZN(n9510)
         );
  OAI211_X1 U10825 ( .C1(n9512), .C2(n9579), .A(n9511), .B(n9510), .ZN(n9601)
         );
  MUX2_X1 U10826 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9601), .S(n10526), .Z(
        P2_U3544) );
  AOI211_X1 U10827 ( .C1(n9588), .C2(n9515), .A(n9514), .B(n9513), .ZN(n9516)
         );
  OAI21_X1 U10828 ( .B1(n9579), .B2(n9517), .A(n9516), .ZN(n9602) );
  MUX2_X1 U10829 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9602), .S(n10526), .Z(
        P2_U3543) );
  AOI211_X1 U10830 ( .C1(n9588), .C2(n9520), .A(n9519), .B(n9518), .ZN(n9521)
         );
  OAI21_X1 U10831 ( .B1(n9579), .B2(n9522), .A(n9521), .ZN(n9603) );
  MUX2_X1 U10832 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9603), .S(n10526), .Z(
        P2_U3542) );
  AOI22_X1 U10833 ( .A1(n9524), .A2(n9589), .B1(n9588), .B2(n9523), .ZN(n9525)
         );
  OAI211_X1 U10834 ( .C1(n9579), .C2(n9527), .A(n9526), .B(n9525), .ZN(n9604)
         );
  MUX2_X1 U10835 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9604), .S(n10526), .Z(
        P2_U3541) );
  AOI22_X1 U10836 ( .A1(n9529), .A2(n9589), .B1(n9588), .B2(n9528), .ZN(n9532)
         );
  NAND3_X1 U10837 ( .A1(n9530), .A2(n10512), .A3(n9323), .ZN(n9531) );
  NAND3_X1 U10838 ( .A1(n9533), .A2(n9532), .A3(n9531), .ZN(n9605) );
  MUX2_X1 U10839 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9605), .S(n10526), .Z(
        P2_U3540) );
  AOI21_X1 U10840 ( .B1(n9588), .B2(n9535), .A(n9534), .ZN(n9536) );
  OAI211_X1 U10841 ( .C1(n9579), .C2(n9538), .A(n9537), .B(n9536), .ZN(n9606)
         );
  MUX2_X1 U10842 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9606), .S(n10526), .Z(
        P2_U3539) );
  AOI22_X1 U10843 ( .A1(n9540), .A2(n9589), .B1(n9588), .B2(n9539), .ZN(n9541)
         );
  OAI211_X1 U10844 ( .C1(n9579), .C2(n9543), .A(n9542), .B(n9541), .ZN(n9607)
         );
  MUX2_X1 U10845 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9607), .S(n10526), .Z(
        P2_U3538) );
  AOI21_X1 U10846 ( .B1(n9588), .B2(n9545), .A(n9544), .ZN(n9546) );
  OAI211_X1 U10847 ( .C1(n9579), .C2(n9548), .A(n9547), .B(n9546), .ZN(n9608)
         );
  MUX2_X1 U10848 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9608), .S(n10526), .Z(
        P2_U3537) );
  OAI22_X1 U10849 ( .A1(n9550), .A2(n10508), .B1(n9549), .B2(n10507), .ZN(
        n9551) );
  AOI21_X1 U10850 ( .B1(n9553), .B2(n9552), .A(n9551), .ZN(n9554) );
  NAND2_X1 U10851 ( .A1(n9555), .A2(n9554), .ZN(n9609) );
  MUX2_X1 U10852 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9609), .S(n10526), .Z(
        P2_U3536) );
  AOI22_X1 U10853 ( .A1(n9557), .A2(n9589), .B1(n9588), .B2(n9556), .ZN(n9558)
         );
  OAI211_X1 U10854 ( .C1(n9579), .C2(n9560), .A(n9559), .B(n9558), .ZN(n9610)
         );
  MUX2_X1 U10855 ( .A(n9610), .B(P2_REG1_REG_15__SCAN_IN), .S(n10523), .Z(
        P2_U3535) );
  AOI21_X1 U10856 ( .B1(n9588), .B2(n6337), .A(n9561), .ZN(n9562) );
  OAI211_X1 U10857 ( .C1(n9579), .C2(n9564), .A(n9563), .B(n9562), .ZN(n9611)
         );
  MUX2_X1 U10858 ( .A(n9611), .B(P2_REG1_REG_14__SCAN_IN), .S(n10523), .Z(
        P2_U3534) );
  AOI22_X1 U10859 ( .A1(n9566), .A2(n9589), .B1(n9588), .B2(n9565), .ZN(n9567)
         );
  OAI211_X1 U10860 ( .C1(n9569), .C2(n9594), .A(n9568), .B(n9567), .ZN(n9612)
         );
  MUX2_X1 U10861 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n9612), .S(n10526), .Z(
        P2_U3533) );
  AOI22_X1 U10862 ( .A1(n9570), .A2(n9589), .B1(n9588), .B2(n6570), .ZN(n9571)
         );
  OAI211_X1 U10863 ( .C1(n9573), .C2(n9579), .A(n9572), .B(n9571), .ZN(n9613)
         );
  MUX2_X1 U10864 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n9613), .S(n10526), .Z(
        P2_U3532) );
  AOI22_X1 U10865 ( .A1(n9575), .A2(n9589), .B1(n9588), .B2(n9574), .ZN(n9576)
         );
  OAI211_X1 U10866 ( .C1(n9579), .C2(n9578), .A(n9577), .B(n9576), .ZN(n9614)
         );
  MUX2_X1 U10867 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n9614), .S(n10526), .Z(
        P2_U3531) );
  AOI22_X1 U10868 ( .A1(n9581), .A2(n9589), .B1(n9588), .B2(n9580), .ZN(n9585)
         );
  NAND3_X1 U10869 ( .A1(n9583), .A2(n10512), .A3(n9582), .ZN(n9584) );
  NAND3_X1 U10870 ( .A1(n9586), .A2(n9585), .A3(n9584), .ZN(n9615) );
  MUX2_X1 U10871 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n9615), .S(n10526), .Z(
        P2_U3530) );
  AOI22_X1 U10872 ( .A1(n9590), .A2(n9589), .B1(n9588), .B2(n9587), .ZN(n9591)
         );
  OAI211_X1 U10873 ( .C1(n9594), .C2(n9593), .A(n9592), .B(n9591), .ZN(n9616)
         );
  MUX2_X1 U10874 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n9616), .S(n10526), .Z(
        P2_U3529) );
  MUX2_X1 U10875 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9595), .S(n10516), .Z(
        P2_U3519) );
  MUX2_X1 U10876 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9597), .S(n10516), .Z(
        P2_U3516) );
  MUX2_X1 U10877 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9598), .S(n10516), .Z(
        P2_U3515) );
  MUX2_X1 U10878 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9599), .S(n10516), .Z(
        P2_U3514) );
  MUX2_X1 U10879 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9600), .S(n10516), .Z(
        P2_U3513) );
  MUX2_X1 U10880 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9601), .S(n10516), .Z(
        P2_U3512) );
  MUX2_X1 U10881 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9602), .S(n10516), .Z(
        P2_U3511) );
  MUX2_X1 U10882 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9603), .S(n10516), .Z(
        P2_U3510) );
  MUX2_X1 U10883 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9604), .S(n10516), .Z(
        P2_U3509) );
  MUX2_X1 U10884 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9605), .S(n10516), .Z(
        P2_U3508) );
  MUX2_X1 U10885 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9606), .S(n10516), .Z(
        P2_U3507) );
  MUX2_X1 U10886 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9607), .S(n10516), .Z(
        P2_U3505) );
  MUX2_X1 U10887 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9608), .S(n10516), .Z(
        P2_U3502) );
  MUX2_X1 U10888 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9609), .S(n10516), .Z(
        P2_U3499) );
  MUX2_X1 U10889 ( .A(n9610), .B(P2_REG0_REG_15__SCAN_IN), .S(n10514), .Z(
        P2_U3496) );
  MUX2_X1 U10890 ( .A(n9611), .B(P2_REG0_REG_14__SCAN_IN), .S(n10514), .Z(
        P2_U3493) );
  MUX2_X1 U10891 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n9612), .S(n10516), .Z(
        P2_U3490) );
  MUX2_X1 U10892 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n9613), .S(n10516), .Z(
        P2_U3487) );
  MUX2_X1 U10893 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n9614), .S(n10516), .Z(
        P2_U3484) );
  MUX2_X1 U10894 ( .A(P2_REG0_REG_10__SCAN_IN), .B(n9615), .S(n10516), .Z(
        P2_U3481) );
  MUX2_X1 U10895 ( .A(P2_REG0_REG_9__SCAN_IN), .B(n9616), .S(n10516), .Z(
        P2_U3478) );
  INV_X1 U10896 ( .A(n9617), .ZN(n10231) );
  NOR4_X1 U10897 ( .A1(n9619), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3152), .A4(
        n6033), .ZN(n9620) );
  AOI21_X1 U10898 ( .B1(n9621), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9620), .ZN(
        n9622) );
  OAI21_X1 U10899 ( .B1(n10231), .B2(n9627), .A(n9622), .ZN(P2_U3327) );
  INV_X1 U10900 ( .A(n9623), .ZN(n10236) );
  OAI222_X1 U10901 ( .A1(n9627), .A2(n10236), .B1(n9626), .B2(P2_U3152), .C1(
        n9625), .C2(n9624), .ZN(P2_U3329) );
  INV_X1 U10902 ( .A(n9628), .ZN(n9629) );
  MUX2_X1 U10903 ( .A(n9629), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  OAI22_X1 U10904 ( .A1(n9872), .A2(n9778), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9633), .ZN(n9636) );
  NOR2_X1 U10905 ( .A1(n9634), .A2(n9683), .ZN(n9635) );
  AOI211_X1 U10906 ( .C1(n9637), .C2(n9713), .A(n9636), .B(n9635), .ZN(n9638)
         );
  NAND2_X1 U10907 ( .A1(n9641), .A2(n9640), .ZN(n9642) );
  XOR2_X1 U10908 ( .A(n9643), .B(n9642), .Z(n9651) );
  OAI21_X1 U10909 ( .B1(n9778), .B2(n9645), .A(n9644), .ZN(n9646) );
  AOI21_X1 U10910 ( .B1(n9780), .B2(n10012), .A(n9646), .ZN(n9647) );
  OAI21_X1 U10911 ( .B1(n9782), .B2(n9648), .A(n9647), .ZN(n9649) );
  AOI21_X1 U10912 ( .B1(n9784), .B2(n10181), .A(n9649), .ZN(n9650) );
  OAI21_X1 U10913 ( .B1(n9651), .B2(n9760), .A(n9650), .ZN(P1_U3213) );
  INV_X1 U10914 ( .A(n9655), .ZN(n9653) );
  NAND2_X1 U10915 ( .A1(n9653), .A2(n9652), .ZN(n9657) );
  NAND2_X1 U10916 ( .A1(n9657), .A2(n9656), .ZN(n9722) );
  INV_X1 U10917 ( .A(n9722), .ZN(n9659) );
  NAND2_X1 U10918 ( .A1(n9655), .A2(n9654), .ZN(n9721) );
  AOI21_X1 U10919 ( .B1(n9657), .B2(n9721), .A(n9656), .ZN(n9658) );
  AOI21_X1 U10920 ( .B1(n9659), .B2(n9721), .A(n9658), .ZN(n9664) );
  NAND2_X1 U10921 ( .A1(n9905), .A2(n9780), .ZN(n9661) );
  AOI22_X1 U10922 ( .A1(n9903), .A2(n9735), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n9660) );
  OAI211_X1 U10923 ( .C1(n9782), .C2(n9897), .A(n9661), .B(n9660), .ZN(n9662)
         );
  AOI21_X1 U10924 ( .B1(n10129), .B2(n9784), .A(n9662), .ZN(n9663) );
  OAI21_X1 U10925 ( .B1(n9664), .B2(n9760), .A(n9663), .ZN(P1_U3214) );
  NOR2_X1 U10926 ( .A1(n9666), .A2(n9665), .ZN(n9751) );
  NAND2_X1 U10927 ( .A1(n9666), .A2(n9665), .ZN(n9752) );
  OAI21_X1 U10928 ( .B1(n9751), .B2(n9667), .A(n9752), .ZN(n9672) );
  OAI21_X1 U10929 ( .B1(n9670), .B2(n9669), .A(n9668), .ZN(n9671) );
  XNOR2_X1 U10930 ( .A(n9672), .B(n9671), .ZN(n9678) );
  NAND2_X1 U10931 ( .A1(n9713), .A2(n9960), .ZN(n9675) );
  AOI21_X1 U10932 ( .B1(n9735), .B2(n10003), .A(n9673), .ZN(n9674) );
  OAI211_X1 U10933 ( .C1(n9929), .C2(n9683), .A(n9675), .B(n9674), .ZN(n9676)
         );
  AOI21_X1 U10934 ( .B1(n10150), .B2(n9784), .A(n9676), .ZN(n9677) );
  OAI21_X1 U10935 ( .B1(n9678), .B2(n9760), .A(n9677), .ZN(P1_U3217) );
  XOR2_X1 U10936 ( .A(n9680), .B(n9679), .Z(n9686) );
  AOI22_X1 U10937 ( .A1(n9970), .A2(n9735), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n9682) );
  NAND2_X1 U10938 ( .A1(n9713), .A2(n9933), .ZN(n9681) );
  OAI211_X1 U10939 ( .C1(n9930), .C2(n9683), .A(n9682), .B(n9681), .ZN(n9684)
         );
  AOI21_X1 U10940 ( .B1(n10141), .B2(n9784), .A(n9684), .ZN(n9685) );
  OAI21_X1 U10941 ( .B1(n9686), .B2(n9760), .A(n9685), .ZN(P1_U3221) );
  NAND2_X1 U10942 ( .A1(n9688), .A2(n9687), .ZN(n9720) );
  INV_X1 U10943 ( .A(n9688), .ZN(n9690) );
  NOR3_X1 U10944 ( .A1(n9724), .A2(n9690), .A3(n9689), .ZN(n9691) );
  AOI22_X1 U10945 ( .A1(n9874), .A2(n9713), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9692) );
  OAI21_X1 U10946 ( .B1(n9871), .B2(n9778), .A(n9692), .ZN(n9693) );
  AOI21_X1 U10947 ( .B1(n9780), .B2(n9791), .A(n9693), .ZN(n9694) );
  OAI211_X1 U10948 ( .C1(n9877), .C2(n9771), .A(n9695), .B(n9694), .ZN(
        P1_U3223) );
  XNOR2_X1 U10949 ( .A(n9707), .B(n9704), .ZN(n9697) );
  XNOR2_X1 U10950 ( .A(n9696), .B(n9697), .ZN(n9703) );
  AND2_X1 U10951 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10328) );
  NOR2_X1 U10952 ( .A1(n9778), .A2(n9698), .ZN(n9699) );
  AOI211_X1 U10953 ( .C1(n9780), .C2(n10013), .A(n10328), .B(n9699), .ZN(n9700) );
  OAI21_X1 U10954 ( .B1(n9782), .B2(n10018), .A(n9700), .ZN(n9701) );
  AOI21_X1 U10955 ( .B1(n10165), .B2(n9784), .A(n9701), .ZN(n9702) );
  OAI21_X1 U10956 ( .B1(n9703), .B2(n9760), .A(n9702), .ZN(P1_U3224) );
  INV_X1 U10957 ( .A(n9696), .ZN(n9708) );
  OAI21_X1 U10958 ( .B1(n9696), .B2(n9705), .A(n9704), .ZN(n9706) );
  OAI21_X1 U10959 ( .B1(n9708), .B2(n9707), .A(n9706), .ZN(n9712) );
  XNOR2_X1 U10960 ( .A(n9710), .B(n9709), .ZN(n9711) );
  XNOR2_X1 U10961 ( .A(n9712), .B(n9711), .ZN(n9719) );
  NAND2_X1 U10962 ( .A1(n9713), .A2(n9997), .ZN(n9716) );
  NOR2_X1 U10963 ( .A1(n9714), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10341) );
  AOI21_X1 U10964 ( .B1(n10003), .B2(n9780), .A(n10341), .ZN(n9715) );
  OAI211_X1 U10965 ( .C1(n10041), .C2(n9778), .A(n9716), .B(n9715), .ZN(n9717)
         );
  AOI21_X1 U10966 ( .B1(n10159), .B2(n9784), .A(n9717), .ZN(n9718) );
  OAI21_X1 U10967 ( .B1(n9719), .B2(n9760), .A(n9718), .ZN(P1_U3226) );
  AND3_X1 U10968 ( .A1(n9722), .A2(n9721), .A3(n9720), .ZN(n9723) );
  OAI21_X1 U10969 ( .B1(n9724), .B2(n9723), .A(n9772), .ZN(n9729) );
  NOR2_X1 U10970 ( .A1(n9889), .A2(n9782), .ZN(n9727) );
  OAI22_X1 U10971 ( .A1(n9887), .A2(n9778), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9725), .ZN(n9726) );
  AOI211_X1 U10972 ( .C1(n9792), .C2(n9780), .A(n9727), .B(n9726), .ZN(n9728)
         );
  OAI211_X1 U10973 ( .C1(n5025), .C2(n9771), .A(n9729), .B(n9728), .ZN(
        P1_U3227) );
  INV_X1 U10974 ( .A(n9730), .ZN(n9732) );
  NOR2_X1 U10975 ( .A1(n9732), .A2(n9731), .ZN(n9733) );
  XNOR2_X1 U10976 ( .A(n9734), .B(n9733), .ZN(n9740) );
  NAND2_X1 U10977 ( .A1(n9921), .A2(n9780), .ZN(n9737) );
  AOI22_X1 U10978 ( .A1(n9735), .A2(n9793), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9736) );
  OAI211_X1 U10979 ( .C1(n9782), .C2(n9951), .A(n9737), .B(n9736), .ZN(n9738)
         );
  AOI21_X1 U10980 ( .B1(n10146), .B2(n9784), .A(n9738), .ZN(n9739) );
  OAI21_X1 U10981 ( .B1(n9740), .B2(n9760), .A(n9739), .ZN(P1_U3231) );
  NAND2_X1 U10982 ( .A1(n9742), .A2(n9741), .ZN(n9744) );
  XNOR2_X1 U10983 ( .A(n9744), .B(n9743), .ZN(n9750) );
  OAI22_X1 U10984 ( .A1(n9948), .A2(n9778), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9745), .ZN(n9746) );
  AOI21_X1 U10985 ( .B1(n9919), .B2(n9780), .A(n9746), .ZN(n9747) );
  OAI21_X1 U10986 ( .B1(n9782), .B2(n9913), .A(n9747), .ZN(n9748) );
  AOI21_X1 U10987 ( .B1(n10134), .B2(n9784), .A(n9748), .ZN(n9749) );
  OAI21_X1 U10988 ( .B1(n9750), .B2(n9760), .A(n9749), .ZN(P1_U3233) );
  INV_X1 U10989 ( .A(n9751), .ZN(n9753) );
  NAND2_X1 U10990 ( .A1(n9753), .A2(n9752), .ZN(n9755) );
  XNOR2_X1 U10991 ( .A(n9755), .B(n9754), .ZN(n9761) );
  NAND2_X1 U10992 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9826) );
  OAI21_X1 U10993 ( .B1(n9778), .B2(n9983), .A(n9826), .ZN(n9756) );
  AOI21_X1 U10994 ( .B1(n9780), .B2(n9793), .A(n9756), .ZN(n9757) );
  OAI21_X1 U10995 ( .B1(n9782), .B2(n9989), .A(n9757), .ZN(n9758) );
  AOI21_X1 U10996 ( .B1(n10156), .B2(n9784), .A(n9758), .ZN(n9759) );
  OAI21_X1 U10997 ( .B1(n9761), .B2(n9760), .A(n9759), .ZN(P1_U3236) );
  OAI21_X1 U10998 ( .B1(n9764), .B2(n9763), .A(n9762), .ZN(n9765) );
  NAND3_X1 U10999 ( .A1(n4898), .A2(n9772), .A3(n9765), .ZN(n9770) );
  NOR2_X1 U11000 ( .A1(n9888), .A2(n9778), .ZN(n9768) );
  OAI22_X1 U11001 ( .A1(n9863), .A2(n9782), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9766), .ZN(n9767) );
  AOI211_X1 U11002 ( .C1(n4807), .C2(n9780), .A(n9768), .B(n9767), .ZN(n9769)
         );
  OAI211_X1 U11003 ( .C1(n9858), .C2(n9771), .A(n9770), .B(n9769), .ZN(
        P1_U3238) );
  INV_X1 U11004 ( .A(n9777), .ZN(n9774) );
  OAI21_X1 U11005 ( .B1(n9774), .B2(n9773), .A(n9772), .ZN(n9787) );
  AOI21_X1 U11006 ( .B1(n9777), .B2(n9776), .A(n9775), .ZN(n9786) );
  NAND2_X1 U11007 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10314)
         );
  OAI21_X1 U11008 ( .B1(n9778), .B2(n10039), .A(n10314), .ZN(n9779) );
  AOI21_X1 U11009 ( .B1(n9780), .B2(n5611), .A(n9779), .ZN(n9781) );
  OAI21_X1 U11010 ( .B1(n9782), .B2(n10050), .A(n9781), .ZN(n9783) );
  AOI21_X1 U11011 ( .B1(n10170), .B2(n9784), .A(n9783), .ZN(n9785) );
  OAI21_X1 U11012 ( .B1(n9787), .B2(n9786), .A(n9785), .ZN(P1_U3239) );
  MUX2_X1 U11013 ( .A(n9788), .B(P1_DATAO_REG_31__SCAN_IN), .S(n9807), .Z(
        P1_U3586) );
  MUX2_X1 U11014 ( .A(n9789), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9807), .Z(
        P1_U3585) );
  MUX2_X1 U11015 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n10092), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U11016 ( .A(n9790), .B(P1_DATAO_REG_28__SCAN_IN), .S(n9807), .Z(
        P1_U3583) );
  MUX2_X1 U11017 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n4807), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U11018 ( .A(n9791), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9807), .Z(
        P1_U3581) );
  MUX2_X1 U11019 ( .A(n9792), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9807), .Z(
        P1_U3580) );
  MUX2_X1 U11020 ( .A(n9905), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9807), .Z(
        P1_U3579) );
  MUX2_X1 U11021 ( .A(n9919), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9807), .Z(
        P1_U3578) );
  MUX2_X1 U11022 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9903), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U11023 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9921), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U11024 ( .A(n9970), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9807), .Z(
        P1_U3575) );
  MUX2_X1 U11025 ( .A(n9793), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9807), .Z(
        P1_U3574) );
  MUX2_X1 U11026 ( .A(n10003), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9807), .Z(
        P1_U3573) );
  MUX2_X1 U11027 ( .A(n10013), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9807), .Z(
        P1_U3572) );
  MUX2_X1 U11028 ( .A(n5611), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9807), .Z(
        P1_U3571) );
  MUX2_X1 U11029 ( .A(n10012), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9807), .Z(
        P1_U3570) );
  MUX2_X1 U11030 ( .A(n10069), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9807), .Z(
        P1_U3569) );
  MUX2_X1 U11031 ( .A(n9794), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9807), .Z(
        P1_U3568) );
  MUX2_X1 U11032 ( .A(n9795), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9807), .Z(
        P1_U3567) );
  MUX2_X1 U11033 ( .A(n9796), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9807), .Z(
        P1_U3566) );
  MUX2_X1 U11034 ( .A(n9797), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9807), .Z(
        P1_U3565) );
  MUX2_X1 U11035 ( .A(n9798), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9807), .Z(
        P1_U3564) );
  MUX2_X1 U11036 ( .A(n9799), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9807), .Z(
        P1_U3563) );
  MUX2_X1 U11037 ( .A(n9800), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9807), .Z(
        P1_U3562) );
  MUX2_X1 U11038 ( .A(n9801), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9807), .Z(
        P1_U3561) );
  MUX2_X1 U11039 ( .A(n9802), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9807), .Z(
        P1_U3560) );
  MUX2_X1 U11040 ( .A(n9803), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9807), .Z(
        P1_U3559) );
  MUX2_X1 U11041 ( .A(n9804), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9807), .Z(
        P1_U3558) );
  MUX2_X1 U11042 ( .A(n9805), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9807), .Z(
        P1_U3557) );
  MUX2_X1 U11043 ( .A(n9806), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9807), .Z(
        P1_U3556) );
  MUX2_X1 U11044 ( .A(n9808), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9807), .Z(
        P1_U3555) );
  INV_X1 U11045 ( .A(n9809), .ZN(n9810) );
  OAI21_X1 U11046 ( .B1(n9812), .B2(n9811), .A(n9810), .ZN(n9817) );
  AOI211_X1 U11047 ( .C1(n9815), .C2(n9814), .A(n10305), .B(n9813), .ZN(n9816)
         );
  AOI21_X1 U11048 ( .B1(n10344), .B2(n9817), .A(n9816), .ZN(n9822) );
  NAND2_X1 U11049 ( .A1(n10342), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9820) );
  NAND2_X1 U11050 ( .A1(n10317), .A2(n9818), .ZN(n9819) );
  NAND4_X1 U11051 ( .A1(n9822), .A2(n9821), .A3(n9820), .A4(n9819), .ZN(
        P1_U3247) );
  AOI21_X1 U11052 ( .B1(n9825), .B2(n9824), .A(n9823), .ZN(n9834) );
  OAI21_X1 U11053 ( .B1(n10339), .B2(n9827), .A(n9826), .ZN(n9828) );
  AOI21_X1 U11054 ( .B1(n10342), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n9828), .ZN(
        n9833) );
  OAI211_X1 U11055 ( .C1(n9831), .C2(n9830), .A(n10348), .B(n9829), .ZN(n9832)
         );
  OAI211_X1 U11056 ( .C1(n9834), .C2(n10300), .A(n9833), .B(n9832), .ZN(
        P1_U3259) );
  NAND2_X1 U11057 ( .A1(n9843), .A2(n9842), .ZN(n9835) );
  XNOR2_X1 U11058 ( .A(n9835), .B(n10083), .ZN(n10085) );
  NOR2_X1 U11059 ( .A1(n9837), .A2(n9836), .ZN(n10086) );
  INV_X1 U11060 ( .A(n10086), .ZN(n9838) );
  NOR2_X1 U11061 ( .A1(n10020), .A2(n9838), .ZN(n9845) );
  NOR2_X1 U11062 ( .A1(n9839), .A2(n9999), .ZN(n9840) );
  AOI211_X1 U11063 ( .C1(n10020), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9845), .B(
        n9840), .ZN(n9841) );
  OAI21_X1 U11064 ( .B1(n10085), .B2(n10063), .A(n9841), .ZN(P1_U3261) );
  XNOR2_X1 U11065 ( .A(n9843), .B(n9842), .ZN(n10089) );
  NOR2_X1 U11066 ( .A1(n9843), .A2(n9999), .ZN(n9844) );
  AOI211_X1 U11067 ( .C1(n10020), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9845), .B(
        n9844), .ZN(n9846) );
  OAI21_X1 U11068 ( .B1(n10089), .B2(n10063), .A(n9846), .ZN(P1_U3262) );
  INV_X1 U11069 ( .A(n9847), .ZN(n9848) );
  NAND2_X1 U11070 ( .A1(n9883), .A2(n9848), .ZN(n9850) );
  NAND2_X1 U11071 ( .A1(n9850), .A2(n9849), .ZN(n9851) );
  XNOR2_X1 U11072 ( .A(n9851), .B(n9856), .ZN(n9854) );
  OAI22_X1 U11073 ( .A1(n9852), .A2(n10040), .B1(n9888), .B2(n10071), .ZN(
        n9853) );
  AOI21_X1 U11074 ( .B1(n9854), .B2(n10074), .A(n9853), .ZN(n10119) );
  XOR2_X1 U11075 ( .A(n9856), .B(n9855), .Z(n10120) );
  OR2_X1 U11076 ( .A1(n10120), .A2(n10009), .ZN(n9866) );
  NOR2_X1 U11077 ( .A1(n9858), .A2(n9857), .ZN(n9860) );
  NOR2_X1 U11078 ( .A1(n9860), .A2(n9859), .ZN(n10117) );
  NAND2_X1 U11079 ( .A1(n10116), .A2(n10060), .ZN(n9862) );
  NAND2_X1 U11080 ( .A1(n10020), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n9861) );
  OAI211_X1 U11081 ( .C1(n10049), .C2(n9863), .A(n9862), .B(n9861), .ZN(n9864)
         );
  AOI21_X1 U11082 ( .B1(n10117), .B2(n10007), .A(n9864), .ZN(n9865) );
  OAI211_X1 U11083 ( .C1(n10020), .C2(n10119), .A(n9866), .B(n9865), .ZN(
        P1_U3265) );
  XOR2_X1 U11084 ( .A(n9869), .B(n9867), .Z(n10124) );
  NAND2_X1 U11085 ( .A1(n9883), .A2(n9868), .ZN(n9870) );
  INV_X1 U11086 ( .A(n4424), .ZN(n9873) );
  AOI211_X1 U11087 ( .C1(n10123), .C2(n9873), .A(n10413), .B(n9857), .ZN(
        n10122) );
  NAND2_X1 U11088 ( .A1(n10122), .A2(n10024), .ZN(n9876) );
  AOI22_X1 U11089 ( .A1(n9874), .A2(n10059), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10020), .ZN(n9875) );
  OAI211_X1 U11090 ( .C1(n9877), .C2(n9999), .A(n9876), .B(n9875), .ZN(n9878)
         );
  AOI21_X1 U11091 ( .B1(n10121), .B2(n10078), .A(n9878), .ZN(n9879) );
  OAI21_X1 U11092 ( .B1(n10124), .B2(n10009), .A(n9879), .ZN(P1_U3266) );
  XNOR2_X1 U11093 ( .A(n9880), .B(n9886), .ZN(n10128) );
  NAND2_X1 U11094 ( .A1(n9882), .A2(n9881), .ZN(n9885) );
  INV_X1 U11095 ( .A(n9883), .ZN(n9884) );
  AOI211_X1 U11096 ( .C1(n10127), .C2(n9895), .A(n10413), .B(n4424), .ZN(
        n10126) );
  INV_X1 U11097 ( .A(n10126), .ZN(n9890) );
  OAI22_X1 U11098 ( .A1(n9890), .A2(n9990), .B1(n10049), .B2(n9889), .ZN(n9891) );
  OAI21_X1 U11099 ( .B1(n10125), .B2(n9891), .A(n10078), .ZN(n9893) );
  AOI22_X1 U11100 ( .A1(n10127), .A2(n10060), .B1(n10020), .B2(
        P1_REG2_REG_24__SCAN_IN), .ZN(n9892) );
  OAI211_X1 U11101 ( .C1(n10128), .C2(n10009), .A(n9893), .B(n9892), .ZN(
        P1_U3267) );
  XNOR2_X1 U11102 ( .A(n9894), .B(n9902), .ZN(n10133) );
  INV_X1 U11103 ( .A(n9895), .ZN(n9896) );
  AOI21_X1 U11104 ( .B1(n10129), .B2(n9910), .A(n9896), .ZN(n10130) );
  INV_X1 U11105 ( .A(n10129), .ZN(n9900) );
  INV_X1 U11106 ( .A(n9897), .ZN(n9898) );
  AOI22_X1 U11107 ( .A1(n9898), .A2(n10059), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n10020), .ZN(n9899) );
  OAI21_X1 U11108 ( .B1(n9900), .B2(n9999), .A(n9899), .ZN(n9907) );
  XOR2_X1 U11109 ( .A(n9902), .B(n9901), .Z(n9904) );
  AOI211_X1 U11110 ( .C1(n10130), .C2(n10007), .A(n9907), .B(n9906), .ZN(n9908) );
  OAI21_X1 U11111 ( .B1(n10009), .B2(n10133), .A(n9908), .ZN(P1_U3268) );
  XOR2_X1 U11112 ( .A(n9909), .B(n9917), .Z(n10138) );
  INV_X1 U11113 ( .A(n9931), .ZN(n9912) );
  INV_X1 U11114 ( .A(n9910), .ZN(n9911) );
  AOI21_X1 U11115 ( .B1(n10134), .B2(n9912), .A(n9911), .ZN(n10135) );
  INV_X1 U11116 ( .A(n9913), .ZN(n9914) );
  AOI22_X1 U11117 ( .A1(n9914), .A2(n10059), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n10020), .ZN(n9915) );
  OAI21_X1 U11118 ( .B1(n9916), .B2(n9999), .A(n9915), .ZN(n9923) );
  XNOR2_X1 U11119 ( .A(n9918), .B(n9917), .ZN(n9920) );
  AOI222_X1 U11120 ( .A1(n9921), .A2(n10011), .B1(n10074), .B2(n9920), .C1(
        n9919), .C2(n10068), .ZN(n10137) );
  NOR2_X1 U11121 ( .A1(n10137), .A2(n10020), .ZN(n9922) );
  AOI211_X1 U11122 ( .C1(n10135), .C2(n10007), .A(n9923), .B(n9922), .ZN(n9924) );
  OAI21_X1 U11123 ( .B1(n10009), .B2(n10138), .A(n9924), .ZN(P1_U3269) );
  INV_X1 U11124 ( .A(n9925), .ZN(n9926) );
  AOI21_X1 U11125 ( .B1(n9938), .B2(n9927), .A(n9926), .ZN(n9928) );
  OAI222_X1 U11126 ( .A1(n10040), .A2(n9930), .B1(n10071), .B2(n9929), .C1(
        n9928), .C2(n10044), .ZN(n10139) );
  OAI21_X1 U11127 ( .B1(n9950), .B2(n9936), .A(n10429), .ZN(n9932) );
  NOR2_X1 U11128 ( .A1(n9932), .A2(n9931), .ZN(n10140) );
  NAND2_X1 U11129 ( .A1(n10140), .A2(n10024), .ZN(n9935) );
  AOI22_X1 U11130 ( .A1(n9933), .A2(n10059), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n10020), .ZN(n9934) );
  OAI211_X1 U11131 ( .C1(n9936), .C2(n9999), .A(n9935), .B(n9934), .ZN(n9940)
         );
  OAI21_X1 U11132 ( .B1(n4447), .B2(n9938), .A(n9937), .ZN(n10143) );
  NOR2_X1 U11133 ( .A1(n10143), .A2(n10009), .ZN(n9939) );
  AOI211_X1 U11134 ( .C1(n10078), .C2(n10139), .A(n9940), .B(n9939), .ZN(n9941) );
  INV_X1 U11135 ( .A(n9941), .ZN(P1_U3270) );
  XNOR2_X1 U11136 ( .A(n9942), .B(n9946), .ZN(n10148) );
  OR2_X1 U11137 ( .A1(n10002), .A2(n9943), .ZN(n9945) );
  AND2_X1 U11138 ( .A1(n9945), .A2(n9944), .ZN(n9947) );
  XNOR2_X1 U11139 ( .A(n9947), .B(n9946), .ZN(n9949) );
  OAI222_X1 U11140 ( .A1(n9949), .A2(n10044), .B1(n10040), .B2(n9948), .C1(
        n10071), .C2(n9984), .ZN(n10144) );
  AOI211_X1 U11141 ( .C1(n10146), .C2(n9958), .A(n10413), .B(n9950), .ZN(
        n10145) );
  NAND2_X1 U11142 ( .A1(n10145), .A2(n10024), .ZN(n9954) );
  INV_X1 U11143 ( .A(n9951), .ZN(n9952) );
  AOI22_X1 U11144 ( .A1(n9952), .A2(n10059), .B1(P1_REG2_REG_20__SCAN_IN), 
        .B2(n10020), .ZN(n9953) );
  OAI211_X1 U11145 ( .C1(n5022), .C2(n9999), .A(n9954), .B(n9953), .ZN(n9955)
         );
  AOI21_X1 U11146 ( .B1(n10144), .B2(n10078), .A(n9955), .ZN(n9956) );
  OAI21_X1 U11147 ( .B1(n10148), .B2(n10009), .A(n9956), .ZN(P1_U3271) );
  XOR2_X1 U11148 ( .A(n9957), .B(n9969), .Z(n10153) );
  INV_X1 U11149 ( .A(n9958), .ZN(n9959) );
  AOI211_X1 U11150 ( .C1(n10150), .C2(n9986), .A(n10413), .B(n9959), .ZN(
        n10149) );
  AOI22_X1 U11151 ( .A1(n9960), .A2(n10059), .B1(n10020), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n9961) );
  OAI21_X1 U11152 ( .B1(n9962), .B2(n9999), .A(n9961), .ZN(n9973) );
  OR2_X1 U11153 ( .A1(n10002), .A2(n9963), .ZN(n9966) );
  AND2_X1 U11154 ( .A1(n9964), .A2(n9966), .ZN(n9968) );
  NAND2_X1 U11155 ( .A1(n9966), .A2(n9965), .ZN(n9967) );
  OAI21_X1 U11156 ( .B1(n9969), .B2(n9968), .A(n9967), .ZN(n9971) );
  AOI222_X1 U11157 ( .A1(n9971), .A2(n10074), .B1(n9970), .B2(n10068), .C1(
        n10003), .C2(n10011), .ZN(n10152) );
  NOR2_X1 U11158 ( .A1(n10152), .A2(n10020), .ZN(n9972) );
  AOI211_X1 U11159 ( .C1(n10149), .C2(n10024), .A(n9973), .B(n9972), .ZN(n9974) );
  OAI21_X1 U11160 ( .B1(n10009), .B2(n10153), .A(n9974), .ZN(P1_U3272) );
  XNOR2_X1 U11161 ( .A(n9975), .B(n9976), .ZN(n10158) );
  OR2_X1 U11162 ( .A1(n10002), .A2(n9977), .ZN(n9979) );
  NAND2_X1 U11163 ( .A1(n9979), .A2(n9978), .ZN(n9981) );
  XNOR2_X1 U11164 ( .A(n9981), .B(n9980), .ZN(n9982) );
  OAI222_X1 U11165 ( .A1(n10040), .A2(n9984), .B1(n10071), .B2(n9983), .C1(
        n9982), .C2(n10044), .ZN(n10154) );
  INV_X1 U11166 ( .A(n9985), .ZN(n9988) );
  INV_X1 U11167 ( .A(n9986), .ZN(n9987) );
  AOI211_X1 U11168 ( .C1(n10156), .C2(n9988), .A(n10413), .B(n9987), .ZN(
        n10155) );
  INV_X1 U11169 ( .A(n10155), .ZN(n9991) );
  OAI22_X1 U11170 ( .A1(n9991), .A2(n9990), .B1(n10049), .B2(n9989), .ZN(n9992) );
  OAI21_X1 U11171 ( .B1(n10154), .B2(n9992), .A(n10078), .ZN(n9994) );
  AOI22_X1 U11172 ( .A1(n10156), .A2(n10060), .B1(P1_REG2_REG_18__SCAN_IN), 
        .B2(n10020), .ZN(n9993) );
  OAI211_X1 U11173 ( .C1(n10158), .C2(n10009), .A(n9994), .B(n9993), .ZN(
        P1_U3273) );
  XOR2_X1 U11174 ( .A(n9995), .B(n10001), .Z(n10163) );
  INV_X1 U11175 ( .A(n10017), .ZN(n9996) );
  AOI21_X1 U11176 ( .B1(n10159), .B2(n9996), .A(n9985), .ZN(n10160) );
  AOI22_X1 U11177 ( .A1(n10020), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9997), 
        .B2(n10059), .ZN(n9998) );
  OAI21_X1 U11178 ( .B1(n10000), .B2(n9999), .A(n9998), .ZN(n10006) );
  XNOR2_X1 U11179 ( .A(n10002), .B(n10001), .ZN(n10004) );
  AOI222_X1 U11180 ( .A1(n5611), .A2(n10011), .B1(n10074), .B2(n10004), .C1(
        n10003), .C2(n10068), .ZN(n10162) );
  NOR2_X1 U11181 ( .A1(n10162), .A2(n10020), .ZN(n10005) );
  AOI211_X1 U11182 ( .C1(n10160), .C2(n10007), .A(n10006), .B(n10005), .ZN(
        n10008) );
  OAI21_X1 U11183 ( .B1(n10009), .B2(n10163), .A(n10008), .ZN(P1_U3274) );
  XOR2_X1 U11184 ( .A(n7123), .B(n10010), .Z(n10014) );
  AOI222_X1 U11185 ( .A1(n10014), .A2(n10074), .B1(n10013), .B2(n10068), .C1(
        n10012), .C2(n10011), .ZN(n10169) );
  NAND2_X1 U11186 ( .A1(n10048), .A2(n10165), .ZN(n10015) );
  NAND2_X1 U11187 ( .A1(n10015), .A2(n10429), .ZN(n10016) );
  NOR2_X1 U11188 ( .A1(n10017), .A2(n10016), .ZN(n10164) );
  NAND2_X1 U11189 ( .A1(n10165), .A2(n10060), .ZN(n10022) );
  NOR2_X1 U11190 ( .A1(n10018), .A2(n10049), .ZN(n10019) );
  AOI21_X1 U11191 ( .B1(n10020), .B2(P1_REG2_REG_16__SCAN_IN), .A(n10019), 
        .ZN(n10021) );
  NAND2_X1 U11192 ( .A1(n10022), .A2(n10021), .ZN(n10023) );
  AOI21_X1 U11193 ( .B1(n10164), .B2(n10024), .A(n10023), .ZN(n10032) );
  NOR2_X1 U11194 ( .A1(n8733), .A2(n10026), .ZN(n10028) );
  NOR2_X1 U11195 ( .A1(n10028), .A2(n10027), .ZN(n10029) );
  NAND2_X1 U11196 ( .A1(n10029), .A2(n7123), .ZN(n10166) );
  NAND3_X1 U11197 ( .A1(n10025), .A2(n10166), .A3(n10030), .ZN(n10031) );
  OAI211_X1 U11198 ( .C1(n10169), .C2(n10020), .A(n10032), .B(n10031), .ZN(
        P1_U3275) );
  OR2_X1 U11199 ( .A1(n8733), .A2(n10033), .ZN(n10035) );
  NAND2_X1 U11200 ( .A1(n10035), .A2(n10034), .ZN(n10036) );
  XNOR2_X1 U11201 ( .A(n10036), .B(n10037), .ZN(n10174) );
  XNOR2_X1 U11202 ( .A(n10038), .B(n10037), .ZN(n10045) );
  OAI22_X1 U11203 ( .A1(n10041), .A2(n10040), .B1(n10039), .B2(n10071), .ZN(
        n10042) );
  INV_X1 U11204 ( .A(n10042), .ZN(n10043) );
  OAI21_X1 U11205 ( .B1(n10045), .B2(n10044), .A(n10043), .ZN(n10046) );
  AOI21_X1 U11206 ( .B1(n10174), .B2(n10386), .A(n10046), .ZN(n10176) );
  NAND2_X1 U11207 ( .A1(n8734), .A2(n10170), .ZN(n10047) );
  NAND2_X1 U11208 ( .A1(n10048), .A2(n10047), .ZN(n10172) );
  OAI22_X1 U11209 ( .A1(n10078), .A2(n6864), .B1(n10050), .B2(n10049), .ZN(
        n10051) );
  AOI21_X1 U11210 ( .B1(n10170), .B2(n10060), .A(n10051), .ZN(n10052) );
  OAI21_X1 U11211 ( .B1(n10172), .B2(n10063), .A(n10052), .ZN(n10053) );
  AOI21_X1 U11212 ( .B1(n10174), .B2(n10081), .A(n10053), .ZN(n10054) );
  OAI21_X1 U11213 ( .B1(n10176), .B2(n10020), .A(n10054), .ZN(P1_U3276) );
  XNOR2_X1 U11214 ( .A(n10055), .B(n10064), .ZN(n10185) );
  NOR2_X1 U11215 ( .A1(n8631), .A2(n10186), .ZN(n10056) );
  OR2_X1 U11216 ( .A1(n10057), .A2(n10056), .ZN(n10187) );
  AOI22_X1 U11217 ( .A1(n10061), .A2(n10060), .B1(n10059), .B2(n10058), .ZN(
        n10062) );
  OAI21_X1 U11218 ( .B1(n10187), .B2(n10063), .A(n10062), .ZN(n10080) );
  NAND2_X1 U11219 ( .A1(n10185), .A2(n10386), .ZN(n10077) );
  NAND3_X1 U11220 ( .A1(n10066), .A2(n4822), .A3(n10065), .ZN(n10067) );
  NAND2_X1 U11221 ( .A1(n4399), .A2(n10067), .ZN(n10075) );
  NAND2_X1 U11222 ( .A1(n10069), .A2(n10068), .ZN(n10070) );
  OAI21_X1 U11223 ( .B1(n10072), .B2(n10071), .A(n10070), .ZN(n10073) );
  AOI21_X1 U11224 ( .B1(n10075), .B2(n10074), .A(n10073), .ZN(n10076) );
  NAND2_X1 U11225 ( .A1(n10077), .A2(n10076), .ZN(n10189) );
  MUX2_X1 U11226 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n10189), .S(n10078), .Z(
        n10079) );
  AOI211_X1 U11227 ( .C1(n10185), .C2(n10081), .A(n10080), .B(n10079), .ZN(
        n10082) );
  INV_X1 U11228 ( .A(n10082), .ZN(P1_U3278) );
  AOI21_X1 U11229 ( .B1(n10083), .B2(n10428), .A(n10086), .ZN(n10084) );
  OAI21_X1 U11230 ( .B1(n10085), .B2(n10413), .A(n10084), .ZN(n10201) );
  MUX2_X1 U11231 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n10201), .S(n10455), .Z(
        P1_U3554) );
  AOI21_X1 U11232 ( .B1(n10087), .B2(n10428), .A(n10086), .ZN(n10088) );
  OAI21_X1 U11233 ( .B1(n10089), .B2(n10413), .A(n10088), .ZN(n10202) );
  MUX2_X1 U11234 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n10202), .S(n10455), .Z(
        P1_U3553) );
  INV_X1 U11235 ( .A(n10184), .ZN(n10409) );
  NAND2_X1 U11236 ( .A1(n10090), .A2(n10409), .ZN(n10419) );
  NAND4_X1 U11237 ( .A1(n10103), .A2(n10091), .A3(n10419), .A4(n10097), .ZN(
        n10105) );
  NAND2_X1 U11238 ( .A1(n10092), .A2(n10419), .ZN(n10094) );
  OAI211_X1 U11239 ( .C1(n10097), .C2(n10094), .A(n10093), .B(n10400), .ZN(
        n10100) );
  NAND2_X1 U11240 ( .A1(n5852), .A2(n10419), .ZN(n10096) );
  OAI21_X1 U11241 ( .B1(n10097), .B2(n10096), .A(n10095), .ZN(n10099) );
  INV_X1 U11242 ( .A(n10419), .ZN(n10102) );
  MUX2_X1 U11243 ( .A(n10203), .B(P1_REG1_REG_29__SCAN_IN), .S(n10452), .Z(
        P1_U3552) );
  AOI22_X1 U11244 ( .A1(n10108), .A2(n10429), .B1(n10428), .B2(n10107), .ZN(
        n10109) );
  MUX2_X1 U11245 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n10204), .S(n10455), .Z(
        P1_U3551) );
  AOI22_X1 U11246 ( .A1(n10112), .A2(n10429), .B1(n10428), .B2(n7150), .ZN(
        n10113) );
  OAI211_X1 U11247 ( .C1(n10115), .C2(n10102), .A(n10114), .B(n10113), .ZN(
        n10205) );
  MUX2_X1 U11248 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10205), .S(n10455), .Z(
        P1_U3550) );
  AOI22_X1 U11249 ( .A1(n10117), .A2(n10429), .B1(n10428), .B2(n10116), .ZN(
        n10118) );
  OAI211_X1 U11250 ( .C1(n10120), .C2(n10102), .A(n10119), .B(n10118), .ZN(
        n10206) );
  MUX2_X1 U11251 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10206), .S(n10455), .Z(
        P1_U3549) );
  MUX2_X1 U11252 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10207), .S(n10455), .Z(
        P1_U3548) );
  MUX2_X1 U11253 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10208), .S(n10455), .Z(
        P1_U3547) );
  AOI22_X1 U11254 ( .A1(n10130), .A2(n10429), .B1(n10428), .B2(n10129), .ZN(
        n10131) );
  OAI211_X1 U11255 ( .C1(n10102), .C2(n10133), .A(n10132), .B(n10131), .ZN(
        n10209) );
  MUX2_X1 U11256 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10209), .S(n10455), .Z(
        P1_U3546) );
  AOI22_X1 U11257 ( .A1(n10135), .A2(n10429), .B1(n10428), .B2(n10134), .ZN(
        n10136) );
  OAI211_X1 U11258 ( .C1(n10138), .C2(n10102), .A(n10137), .B(n10136), .ZN(
        n10210) );
  MUX2_X1 U11259 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10210), .S(n10455), .Z(
        P1_U3545) );
  AOI211_X1 U11260 ( .C1(n10428), .C2(n10141), .A(n10140), .B(n10139), .ZN(
        n10142) );
  OAI21_X1 U11261 ( .B1(n10102), .B2(n10143), .A(n10142), .ZN(n10211) );
  MUX2_X1 U11262 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10211), .S(n10455), .Z(
        P1_U3544) );
  AOI211_X1 U11263 ( .C1(n10428), .C2(n10146), .A(n10145), .B(n10144), .ZN(
        n10147) );
  OAI21_X1 U11264 ( .B1(n10102), .B2(n10148), .A(n10147), .ZN(n10212) );
  MUX2_X1 U11265 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10212), .S(n10455), .Z(
        P1_U3543) );
  AOI21_X1 U11266 ( .B1(n10428), .B2(n10150), .A(n10149), .ZN(n10151) );
  OAI211_X1 U11267 ( .C1(n10153), .C2(n10102), .A(n10152), .B(n10151), .ZN(
        n10213) );
  MUX2_X1 U11268 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10213), .S(n10455), .Z(
        P1_U3542) );
  AOI211_X1 U11269 ( .C1(n10428), .C2(n10156), .A(n10155), .B(n10154), .ZN(
        n10157) );
  OAI21_X1 U11270 ( .B1(n10102), .B2(n10158), .A(n10157), .ZN(n10214) );
  MUX2_X1 U11271 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10214), .S(n10455), .Z(
        P1_U3541) );
  AOI22_X1 U11272 ( .A1(n10160), .A2(n10429), .B1(n10428), .B2(n10159), .ZN(
        n10161) );
  OAI211_X1 U11273 ( .C1(n10102), .C2(n10163), .A(n10162), .B(n10161), .ZN(
        n10215) );
  MUX2_X1 U11274 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10215), .S(n10455), .Z(
        P1_U3540) );
  AOI21_X1 U11275 ( .B1(n10428), .B2(n10165), .A(n10164), .ZN(n10168) );
  NAND3_X1 U11276 ( .A1(n10025), .A2(n10419), .A3(n10166), .ZN(n10167) );
  NAND3_X1 U11277 ( .A1(n10169), .A2(n10168), .A3(n10167), .ZN(n10216) );
  MUX2_X1 U11278 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10216), .S(n10455), .Z(
        P1_U3539) );
  INV_X1 U11279 ( .A(n10170), .ZN(n10171) );
  OAI22_X1 U11280 ( .A1(n10172), .A2(n10413), .B1(n10171), .B2(n10400), .ZN(
        n10173) );
  AOI21_X1 U11281 ( .B1(n10174), .B2(n10184), .A(n10173), .ZN(n10175) );
  AND2_X1 U11282 ( .A1(n10176), .A2(n10175), .ZN(n10217) );
  MUX2_X1 U11283 ( .A(n10177), .B(n10217), .S(n10455), .Z(n10178) );
  INV_X1 U11284 ( .A(n10178), .ZN(P1_U3538) );
  AOI211_X1 U11285 ( .C1(n10428), .C2(n10181), .A(n10180), .B(n10179), .ZN(
        n10182) );
  OAI21_X1 U11286 ( .B1(n10102), .B2(n10183), .A(n10182), .ZN(n10220) );
  MUX2_X1 U11287 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10220), .S(n10455), .Z(
        P1_U3537) );
  AND2_X1 U11288 ( .A1(n10185), .A2(n10184), .ZN(n10190) );
  OAI22_X1 U11289 ( .A1(n10187), .A2(n10413), .B1(n10186), .B2(n10400), .ZN(
        n10188) );
  MUX2_X1 U11290 ( .A(n10221), .B(P1_REG1_REG_13__SCAN_IN), .S(n10452), .Z(
        P1_U3536) );
  AOI211_X1 U11291 ( .C1(n10428), .C2(n10193), .A(n10192), .B(n10191), .ZN(
        n10194) );
  OAI21_X1 U11292 ( .B1(n10102), .B2(n10195), .A(n10194), .ZN(n10222) );
  MUX2_X1 U11293 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10222), .S(n10455), .Z(
        P1_U3535) );
  AOI22_X1 U11294 ( .A1(n10197), .A2(n10429), .B1(n10428), .B2(n10196), .ZN(
        n10198) );
  OAI211_X1 U11295 ( .C1(n10409), .C2(n10200), .A(n10199), .B(n10198), .ZN(
        n10223) );
  MUX2_X1 U11296 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10223), .S(n10455), .Z(
        P1_U3534) );
  MUX2_X1 U11297 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n10201), .S(n10437), .Z(
        P1_U3522) );
  MUX2_X1 U11298 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10202), .S(n10437), .Z(
        P1_U3521) );
  MUX2_X1 U11299 ( .A(n10203), .B(P1_REG0_REG_29__SCAN_IN), .S(n10435), .Z(
        P1_U3520) );
  MUX2_X1 U11300 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n10204), .S(n10437), .Z(
        P1_U3519) );
  MUX2_X1 U11301 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10205), .S(n10437), .Z(
        P1_U3518) );
  MUX2_X1 U11302 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10206), .S(n10437), .Z(
        P1_U3517) );
  MUX2_X1 U11303 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10207), .S(n10437), .Z(
        P1_U3516) );
  MUX2_X1 U11304 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10208), .S(n10437), .Z(
        P1_U3515) );
  MUX2_X1 U11305 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10209), .S(n10437), .Z(
        P1_U3514) );
  MUX2_X1 U11306 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10210), .S(n10437), .Z(
        P1_U3513) );
  MUX2_X1 U11307 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10211), .S(n10437), .Z(
        P1_U3512) );
  MUX2_X1 U11308 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10212), .S(n10437), .Z(
        P1_U3511) );
  MUX2_X1 U11309 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10213), .S(n10437), .Z(
        P1_U3510) );
  MUX2_X1 U11310 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10214), .S(n10437), .Z(
        P1_U3508) );
  MUX2_X1 U11311 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10215), .S(n10437), .Z(
        P1_U3505) );
  MUX2_X1 U11312 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10216), .S(n10437), .Z(
        P1_U3502) );
  MUX2_X1 U11313 ( .A(n10218), .B(n10217), .S(n10437), .Z(n10219) );
  INV_X1 U11314 ( .A(n10219), .ZN(P1_U3499) );
  MUX2_X1 U11315 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10220), .S(n10437), .Z(
        P1_U3496) );
  MUX2_X1 U11316 ( .A(n10221), .B(P1_REG0_REG_13__SCAN_IN), .S(n10435), .Z(
        P1_U3493) );
  MUX2_X1 U11317 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n10222), .S(n10437), .Z(
        P1_U3490) );
  MUX2_X1 U11318 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n10223), .S(n10437), .Z(
        P1_U3487) );
  MUX2_X1 U11319 ( .A(P1_D_REG_1__SCAN_IN), .B(n10224), .S(n10225), .Z(
        P1_U3441) );
  MUX2_X1 U11320 ( .A(P1_D_REG_0__SCAN_IN), .B(n10226), .S(n10225), .Z(
        P1_U3440) );
  NOR4_X1 U11321 ( .A1(n10227), .A2(P1_IR_REG_30__SCAN_IN), .A3(n5143), .A4(
        P1_U3084), .ZN(n10228) );
  AOI21_X1 U11322 ( .B1(n10229), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10228), 
        .ZN(n10230) );
  OAI21_X1 U11323 ( .B1(n10231), .B2(n4391), .A(n10230), .ZN(P1_U3322) );
  OAI222_X1 U11324 ( .A1(n10234), .A2(P1_U3084), .B1(n4391), .B2(n10233), .C1(
        n10232), .C2(n10238), .ZN(P1_U3323) );
  OAI222_X1 U11325 ( .A1(n10238), .A2(n10237), .B1(n4391), .B2(n10236), .C1(
        n10235), .C2(P1_U3084), .ZN(P1_U3324) );
  MUX2_X1 U11326 ( .A(n10239), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  NOR2_X1 U11327 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10240) );
  AOI21_X1 U11328 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n10240), .ZN(n10534) );
  NOR2_X1 U11329 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10241) );
  AOI21_X1 U11330 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n10241), .ZN(n10537) );
  NOR2_X1 U11331 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10242) );
  AOI21_X1 U11332 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10242), .ZN(n10540) );
  NOR2_X1 U11333 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10243) );
  AOI21_X1 U11334 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n10243), .ZN(n10543) );
  NOR2_X1 U11335 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10244) );
  AOI21_X1 U11336 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10244), .ZN(n10546) );
  NOR2_X1 U11337 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10252) );
  INV_X1 U11338 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10246) );
  AOI22_X1 U11339 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n10246), .B1(
        P2_ADDR_REG_4__SCAN_IN), .B2(n10245), .ZN(n10576) );
  NAND2_X1 U11340 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n10250) );
  XOR2_X1 U11341 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10574) );
  NAND2_X1 U11342 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n10248) );
  XOR2_X1 U11343 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10571) );
  AOI21_X1 U11344 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10527) );
  INV_X1 U11345 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10531) );
  NAND3_X1 U11346 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10529) );
  OAI21_X1 U11347 ( .B1(n10527), .B2(n10531), .A(n10529), .ZN(n10570) );
  NAND2_X1 U11348 ( .A1(n10571), .A2(n10570), .ZN(n10247) );
  NAND2_X1 U11349 ( .A1(n10248), .A2(n10247), .ZN(n10573) );
  NAND2_X1 U11350 ( .A1(n10574), .A2(n10573), .ZN(n10249) );
  NAND2_X1 U11351 ( .A1(n10250), .A2(n10249), .ZN(n10575) );
  NOR2_X1 U11352 ( .A1(n10576), .A2(n10575), .ZN(n10251) );
  NOR2_X1 U11353 ( .A1(n10252), .A2(n10251), .ZN(n10253) );
  NOR2_X1 U11354 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10253), .ZN(n10559) );
  NAND2_X1 U11355 ( .A1(n10255), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n10257) );
  XOR2_X1 U11356 ( .A(n10255), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10557) );
  NAND2_X1 U11357 ( .A1(n10557), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n10256) );
  NAND2_X1 U11358 ( .A1(n10257), .A2(n10256), .ZN(n10258) );
  NAND2_X1 U11359 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n10258), .ZN(n10261) );
  XNOR2_X1 U11360 ( .A(n10259), .B(n10258), .ZN(n10572) );
  NAND2_X1 U11361 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10572), .ZN(n10260) );
  NAND2_X1 U11362 ( .A1(n10261), .A2(n10260), .ZN(n10262) );
  NAND2_X1 U11363 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n10262), .ZN(n10264) );
  XOR2_X1 U11364 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n10262), .Z(n10556) );
  NAND2_X1 U11365 ( .A1(n10556), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n10263) );
  NAND2_X1 U11366 ( .A1(n10264), .A2(n10263), .ZN(n10265) );
  NAND2_X1 U11367 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10265), .ZN(n10561) );
  NAND2_X1 U11368 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n10266) );
  OAI21_X1 U11369 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10266), .ZN(n10554) );
  NAND2_X1 U11370 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n10267) );
  OAI21_X1 U11371 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n10267), .ZN(n10551) );
  NOR2_X1 U11372 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10268) );
  AOI21_X1 U11373 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n10268), .ZN(n10548) );
  NAND2_X1 U11374 ( .A1(n10549), .A2(n10548), .ZN(n10547) );
  NAND2_X1 U11375 ( .A1(n10546), .A2(n10545), .ZN(n10544) );
  NAND2_X1 U11376 ( .A1(n10543), .A2(n10542), .ZN(n10541) );
  OAI21_X1 U11377 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10541), .ZN(n10539) );
  NAND2_X1 U11378 ( .A1(n10539), .A2(n10540), .ZN(n10538) );
  OAI21_X1 U11379 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10538), .ZN(n10536) );
  NAND2_X1 U11380 ( .A1(n10537), .A2(n10536), .ZN(n10535) );
  OAI21_X1 U11381 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10535), .ZN(n10533) );
  NAND2_X1 U11382 ( .A1(n10534), .A2(n10533), .ZN(n10532) );
  NOR2_X1 U11383 ( .A1(n10568), .A2(n10567), .ZN(n10269) );
  NAND2_X1 U11384 ( .A1(n10568), .A2(n10567), .ZN(n10566) );
  OAI21_X1 U11385 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n10269), .A(n10566), 
        .ZN(n10272) );
  XNOR2_X1 U11386 ( .A(n10270), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n10271) );
  XNOR2_X1 U11387 ( .A(n10272), .B(n10271), .ZN(ADD_1071_U4) );
  OAI21_X1 U11388 ( .B1(n10339), .B2(n10274), .A(n10273), .ZN(n10275) );
  AOI21_X1 U11389 ( .B1(n10342), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n10275), .ZN(
        n10286) );
  AOI211_X1 U11390 ( .C1(n10278), .C2(n10277), .A(n10276), .B(n10305), .ZN(
        n10279) );
  INV_X1 U11391 ( .A(n10279), .ZN(n10285) );
  AOI211_X1 U11392 ( .C1(n10282), .C2(n10281), .A(n10300), .B(n10280), .ZN(
        n10283) );
  INV_X1 U11393 ( .A(n10283), .ZN(n10284) );
  NAND3_X1 U11394 ( .A1(n10286), .A2(n10285), .A3(n10284), .ZN(P1_U3244) );
  XNOR2_X1 U11395 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11396 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AOI22_X1 U11397 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n10342), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .ZN(n10297) );
  AOI21_X1 U11398 ( .B1(n10289), .B2(P1_REG1_REG_0__SCAN_IN), .A(n10288), .ZN(
        n10290) );
  NOR4_X1 U11399 ( .A1(n10292), .A2(n10291), .A3(n10290), .A4(P1_U3084), .ZN(
        n10293) );
  NAND2_X1 U11400 ( .A1(P1_U3083), .A2(n10293), .ZN(n10296) );
  NAND3_X1 U11401 ( .A1(n10344), .A2(P1_IR_REG_0__SCAN_IN), .A3(n5124), .ZN(
        n10295) );
  NAND3_X1 U11402 ( .A1(n10297), .A2(n10296), .A3(n10295), .ZN(P1_U3241) );
  OAI22_X1 U11403 ( .A1(n10339), .A2(n10298), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7877), .ZN(n10299) );
  AOI21_X1 U11404 ( .B1(n10342), .B2(P1_ADDR_REG_2__SCAN_IN), .A(n10299), .ZN(
        n10313) );
  AOI211_X1 U11405 ( .C1(n10303), .C2(n10302), .A(n10301), .B(n10300), .ZN(
        n10304) );
  INV_X1 U11406 ( .A(n10304), .ZN(n10311) );
  AOI211_X1 U11407 ( .C1(n10308), .C2(n10307), .A(n10306), .B(n10305), .ZN(
        n10309) );
  INV_X1 U11408 ( .A(n10309), .ZN(n10310) );
  NAND4_X1 U11409 ( .A1(n10313), .A2(n10312), .A3(n10311), .A4(n10310), .ZN(
        P1_U3243) );
  INV_X1 U11410 ( .A(n10314), .ZN(n10315) );
  AOI21_X1 U11411 ( .B1(n10317), .B2(n10316), .A(n10315), .ZN(n10325) );
  OAI211_X1 U11412 ( .C1(n10319), .C2(P1_REG1_REG_15__SCAN_IN), .A(n10344), 
        .B(n10318), .ZN(n10324) );
  NAND2_X1 U11413 ( .A1(n10342), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n10323) );
  OAI211_X1 U11414 ( .C1(n10321), .C2(P1_REG2_REG_15__SCAN_IN), .A(n10348), 
        .B(n10320), .ZN(n10322) );
  NAND4_X1 U11415 ( .A1(n10325), .A2(n10324), .A3(n10323), .A4(n10322), .ZN(
        P1_U3256) );
  NOR2_X1 U11416 ( .A1(n10339), .A2(n10326), .ZN(n10327) );
  AOI211_X1 U11417 ( .C1(n10342), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n10328), 
        .B(n10327), .ZN(n10337) );
  OAI211_X1 U11418 ( .C1(n10331), .C2(n10330), .A(n10344), .B(n10329), .ZN(
        n10336) );
  OAI211_X1 U11419 ( .C1(n10334), .C2(n10333), .A(n10348), .B(n10332), .ZN(
        n10335) );
  NAND3_X1 U11420 ( .A1(n10337), .A2(n10336), .A3(n10335), .ZN(P1_U3257) );
  NOR2_X1 U11421 ( .A1(n10339), .A2(n10338), .ZN(n10340) );
  AOI211_X1 U11422 ( .C1(n10342), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n10341), 
        .B(n10340), .ZN(n10353) );
  OAI211_X1 U11423 ( .C1(n10346), .C2(n10345), .A(n10344), .B(n10343), .ZN(
        n10352) );
  OAI211_X1 U11424 ( .C1(n10350), .C2(n10349), .A(n10348), .B(n10347), .ZN(
        n10351) );
  NAND3_X1 U11425 ( .A1(n10353), .A2(n10352), .A3(n10351), .ZN(P1_U3258) );
  AND2_X1 U11426 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10364), .ZN(P1_U3292) );
  NOR2_X1 U11427 ( .A1(n10367), .A2(n10356), .ZN(P1_U3293) );
  AND2_X1 U11428 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10364), .ZN(P1_U3294) );
  AND2_X1 U11429 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10364), .ZN(P1_U3295) );
  AND2_X1 U11430 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10364), .ZN(P1_U3296) );
  AND2_X1 U11431 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10364), .ZN(P1_U3297) );
  AND2_X1 U11432 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10364), .ZN(P1_U3298) );
  NOR2_X1 U11433 ( .A1(n10367), .A2(n10357), .ZN(P1_U3299) );
  NOR2_X1 U11434 ( .A1(n10367), .A2(n10358), .ZN(P1_U3300) );
  AND2_X1 U11435 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10364), .ZN(P1_U3301) );
  AND2_X1 U11436 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10364), .ZN(P1_U3302) );
  AND2_X1 U11437 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10364), .ZN(P1_U3303) );
  AND2_X1 U11438 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10364), .ZN(P1_U3304) );
  AND2_X1 U11439 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10364), .ZN(P1_U3305) );
  NOR2_X1 U11440 ( .A1(n10367), .A2(n10359), .ZN(P1_U3306) );
  NOR2_X1 U11441 ( .A1(n10367), .A2(n10360), .ZN(P1_U3307) );
  AND2_X1 U11442 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10364), .ZN(P1_U3308) );
  AND2_X1 U11443 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10364), .ZN(P1_U3309) );
  AND2_X1 U11444 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10364), .ZN(P1_U3310) );
  NOR2_X1 U11445 ( .A1(n10367), .A2(n10361), .ZN(P1_U3311) );
  AND2_X1 U11446 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10364), .ZN(P1_U3312) );
  NOR2_X1 U11447 ( .A1(n10367), .A2(n10362), .ZN(P1_U3313) );
  AND2_X1 U11448 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10364), .ZN(P1_U3314) );
  AND2_X1 U11449 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10364), .ZN(P1_U3315) );
  AND2_X1 U11450 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10364), .ZN(P1_U3316) );
  INV_X1 U11451 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10363) );
  NOR2_X1 U11452 ( .A1(n10367), .A2(n10363), .ZN(P1_U3317) );
  AND2_X1 U11453 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10364), .ZN(P1_U3318) );
  AND2_X1 U11454 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10364), .ZN(P1_U3319) );
  NOR2_X1 U11455 ( .A1(n10367), .A2(n10365), .ZN(P1_U3320) );
  NOR2_X1 U11456 ( .A1(n10367), .A2(n10366), .ZN(P1_U3321) );
  AOI21_X1 U11457 ( .B1(n10428), .B2(n7153), .A(n10368), .ZN(n10369) );
  OAI21_X1 U11458 ( .B1(n10370), .B2(n10102), .A(n10369), .ZN(n10371) );
  NOR2_X1 U11459 ( .A1(n10372), .A2(n10371), .ZN(n10439) );
  INV_X1 U11460 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10373) );
  AOI22_X1 U11461 ( .A1(n10437), .A2(n10439), .B1(n10373), .B2(n10435), .ZN(
        P1_U3457) );
  OAI21_X1 U11462 ( .B1(n10375), .B2(n10413), .A(n10374), .ZN(n10377) );
  AOI211_X1 U11463 ( .C1(n10419), .C2(n10378), .A(n10377), .B(n10376), .ZN(
        n10441) );
  INV_X1 U11464 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10379) );
  AOI22_X1 U11465 ( .A1(n10437), .A2(n10441), .B1(n10379), .B2(n10435), .ZN(
        P1_U3460) );
  OAI22_X1 U11466 ( .A1(n10381), .A2(n10413), .B1(n10380), .B2(n10400), .ZN(
        n10383) );
  AOI211_X1 U11467 ( .C1(n10419), .C2(n10384), .A(n10383), .B(n10382), .ZN(
        n10443) );
  AOI22_X1 U11468 ( .A1(n10437), .A2(n10443), .B1(n10385), .B2(n10435), .ZN(
        P1_U3463) );
  INV_X1 U11469 ( .A(n10387), .ZN(n10393) );
  NAND2_X1 U11470 ( .A1(n10387), .A2(n10386), .ZN(n10392) );
  OAI22_X1 U11471 ( .A1(n10389), .A2(n10413), .B1(n10388), .B2(n10400), .ZN(
        n10390) );
  INV_X1 U11472 ( .A(n10390), .ZN(n10391) );
  OAI211_X1 U11473 ( .C1(n10393), .C2(n10409), .A(n10392), .B(n10391), .ZN(
        n10394) );
  INV_X1 U11474 ( .A(n10394), .ZN(n10396) );
  AND2_X1 U11475 ( .A1(n10396), .A2(n10395), .ZN(n10445) );
  INV_X1 U11476 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10397) );
  AOI22_X1 U11477 ( .A1(n10437), .A2(n10445), .B1(n10397), .B2(n10435), .ZN(
        P1_U3466) );
  NAND2_X1 U11478 ( .A1(n10398), .A2(n10419), .ZN(n10405) );
  OAI21_X1 U11479 ( .B1(n10401), .B2(n10400), .A(n10399), .ZN(n10402) );
  NOR2_X1 U11480 ( .A1(n10403), .A2(n10402), .ZN(n10404) );
  NAND2_X1 U11481 ( .A1(n10405), .A2(n10404), .ZN(n10406) );
  NOR2_X1 U11482 ( .A1(n10407), .A2(n10406), .ZN(n10447) );
  INV_X1 U11483 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10408) );
  AOI22_X1 U11484 ( .A1(n10437), .A2(n10447), .B1(n10408), .B2(n10435), .ZN(
        P1_U3469) );
  NOR2_X1 U11485 ( .A1(n10410), .A2(n10409), .ZN(n10416) );
  INV_X1 U11486 ( .A(n10411), .ZN(n10412) );
  OAI21_X1 U11487 ( .B1(n10414), .B2(n10413), .A(n10412), .ZN(n10415) );
  NOR3_X1 U11488 ( .A1(n10417), .A2(n10416), .A3(n10415), .ZN(n10449) );
  INV_X1 U11489 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10418) );
  AOI22_X1 U11490 ( .A1(n10437), .A2(n10449), .B1(n10418), .B2(n10435), .ZN(
        P1_U3472) );
  AND2_X1 U11491 ( .A1(n10420), .A2(n10419), .ZN(n10424) );
  NAND2_X1 U11492 ( .A1(n10422), .A2(n10421), .ZN(n10423) );
  NOR3_X1 U11493 ( .A1(n10425), .A2(n10424), .A3(n10423), .ZN(n10451) );
  AOI22_X1 U11494 ( .A1(n10437), .A2(n10451), .B1(n10426), .B2(n10435), .ZN(
        P1_U3475) );
  AOI22_X1 U11495 ( .A1(n10430), .A2(n10429), .B1(n10428), .B2(n10427), .ZN(
        n10431) );
  OAI211_X1 U11496 ( .C1(n10102), .C2(n10433), .A(n10432), .B(n10431), .ZN(
        n10434) );
  INV_X1 U11497 ( .A(n10434), .ZN(n10454) );
  AOI22_X1 U11498 ( .A1(n10437), .A2(n10454), .B1(n10436), .B2(n10435), .ZN(
        P1_U3478) );
  AOI22_X1 U11499 ( .A1(n10455), .A2(n10439), .B1(n10438), .B2(n10452), .ZN(
        P1_U3524) );
  AOI22_X1 U11500 ( .A1(n10455), .A2(n10441), .B1(n10440), .B2(n10452), .ZN(
        P1_U3525) );
  AOI22_X1 U11501 ( .A1(n10455), .A2(n10443), .B1(n10442), .B2(n10452), .ZN(
        P1_U3526) );
  AOI22_X1 U11502 ( .A1(n10455), .A2(n10445), .B1(n10444), .B2(n10452), .ZN(
        P1_U3527) );
  AOI22_X1 U11503 ( .A1(n10455), .A2(n10447), .B1(n10446), .B2(n10452), .ZN(
        P1_U3528) );
  AOI22_X1 U11504 ( .A1(n10455), .A2(n10449), .B1(n10448), .B2(n10452), .ZN(
        P1_U3529) );
  AOI22_X1 U11505 ( .A1(n10455), .A2(n10451), .B1(n10450), .B2(n10452), .ZN(
        P1_U3530) );
  AOI22_X1 U11506 ( .A1(n10455), .A2(n10454), .B1(n10453), .B2(n10452), .ZN(
        P1_U3531) );
  NAND2_X1 U11507 ( .A1(n10457), .A2(n10456), .ZN(n10490) );
  INV_X1 U11508 ( .A(n10458), .ZN(n10459) );
  AOI21_X1 U11509 ( .B1(n10460), .B2(n10490), .A(n10459), .ZN(n10492) );
  AOI22_X1 U11510 ( .A1(n10462), .A2(P2_REG3_REG_0__SCAN_IN), .B1(
        P2_REG2_REG_0__SCAN_IN), .B2(n10461), .ZN(n10469) );
  AOI21_X1 U11511 ( .B1(n10465), .B2(n10464), .A(n10463), .ZN(n10466) );
  AOI21_X1 U11512 ( .B1(n10467), .B2(n10490), .A(n10466), .ZN(n10468) );
  OAI211_X1 U11513 ( .C1(n10470), .C2(n10492), .A(n10469), .B(n10468), .ZN(
        P2_U3296) );
  AND2_X1 U11514 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10484), .ZN(P2_U3297) );
  AND2_X1 U11515 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10484), .ZN(P2_U3298) );
  AND2_X1 U11516 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10484), .ZN(P2_U3299) );
  NOR2_X1 U11517 ( .A1(n10481), .A2(n10473), .ZN(P2_U3300) );
  NOR2_X1 U11518 ( .A1(n10481), .A2(n10474), .ZN(P2_U3301) );
  NOR2_X1 U11519 ( .A1(n10481), .A2(n10475), .ZN(P2_U3302) );
  NOR2_X1 U11520 ( .A1(n10481), .A2(n10476), .ZN(P2_U3303) );
  AND2_X1 U11521 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10484), .ZN(P2_U3304) );
  AND2_X1 U11522 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10484), .ZN(P2_U3305) );
  AND2_X1 U11523 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10484), .ZN(P2_U3306) );
  AND2_X1 U11524 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10484), .ZN(P2_U3307) );
  AND2_X1 U11525 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10484), .ZN(P2_U3308) );
  AND2_X1 U11526 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10484), .ZN(P2_U3309) );
  NOR2_X1 U11527 ( .A1(n10481), .A2(n10477), .ZN(P2_U3310) );
  AND2_X1 U11528 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10484), .ZN(P2_U3311) );
  AND2_X1 U11529 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10484), .ZN(P2_U3312) );
  AND2_X1 U11530 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10484), .ZN(P2_U3313) );
  AND2_X1 U11531 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10484), .ZN(P2_U3314) );
  AND2_X1 U11532 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10484), .ZN(P2_U3315) );
  AND2_X1 U11533 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10484), .ZN(P2_U3316) );
  NOR2_X1 U11534 ( .A1(n10481), .A2(n10478), .ZN(P2_U3317) );
  AND2_X1 U11535 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10484), .ZN(P2_U3318) );
  AND2_X1 U11536 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10484), .ZN(P2_U3319) );
  AND2_X1 U11537 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10484), .ZN(P2_U3320) );
  AND2_X1 U11538 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10484), .ZN(P2_U3321) );
  AND2_X1 U11539 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10484), .ZN(P2_U3322) );
  NOR2_X1 U11540 ( .A1(n10481), .A2(n10479), .ZN(P2_U3323) );
  NOR2_X1 U11541 ( .A1(n10481), .A2(n10480), .ZN(P2_U3324) );
  AND2_X1 U11542 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10484), .ZN(P2_U3325) );
  AND2_X1 U11543 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10484), .ZN(P2_U3326) );
  AOI22_X1 U11544 ( .A1(n10487), .A2(n10483), .B1(n10482), .B2(n10484), .ZN(
        P2_U3437) );
  AOI22_X1 U11545 ( .A1(n10487), .A2(n10486), .B1(n10485), .B2(n10484), .ZN(
        P2_U3438) );
  AOI22_X1 U11546 ( .A1(n10512), .A2(n10490), .B1(n10489), .B2(n10488), .ZN(
        n10491) );
  AND2_X1 U11547 ( .A1(n10492), .A2(n10491), .ZN(n10518) );
  AOI22_X1 U11548 ( .A1(n10516), .A2(n10518), .B1(n6188), .B2(n10514), .ZN(
        P2_U3451) );
  INV_X1 U11549 ( .A(n10493), .ZN(n10495) );
  OAI22_X1 U11550 ( .A1(n10495), .A2(n10508), .B1(n10494), .B2(n10507), .ZN(
        n10497) );
  AOI211_X1 U11551 ( .C1(n10512), .C2(n10498), .A(n10497), .B(n10496), .ZN(
        n10520) );
  INV_X1 U11552 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10499) );
  AOI22_X1 U11553 ( .A1(n10516), .A2(n10520), .B1(n10499), .B2(n10514), .ZN(
        P2_U3463) );
  INV_X1 U11554 ( .A(n10500), .ZN(n10505) );
  OAI22_X1 U11555 ( .A1(n10501), .A2(n10508), .B1(n4847), .B2(n10507), .ZN(
        n10504) );
  INV_X1 U11556 ( .A(n10502), .ZN(n10503) );
  AOI211_X1 U11557 ( .C1(n10505), .C2(n10512), .A(n10504), .B(n10503), .ZN(
        n10522) );
  INV_X1 U11558 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10506) );
  AOI22_X1 U11559 ( .A1(n10516), .A2(n10522), .B1(n10506), .B2(n10514), .ZN(
        P2_U3469) );
  OAI22_X1 U11560 ( .A1(n10509), .A2(n10508), .B1(n4845), .B2(n10507), .ZN(
        n10511) );
  AOI211_X1 U11561 ( .C1(n10513), .C2(n10512), .A(n10511), .B(n10510), .ZN(
        n10525) );
  INV_X1 U11562 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10515) );
  AOI22_X1 U11563 ( .A1(n10516), .A2(n10525), .B1(n10515), .B2(n10514), .ZN(
        P2_U3472) );
  AOI22_X1 U11564 ( .A1(n10526), .A2(n10518), .B1(n10517), .B2(n10523), .ZN(
        P2_U3520) );
  AOI22_X1 U11565 ( .A1(n10526), .A2(n10520), .B1(n10519), .B2(n10523), .ZN(
        P2_U3524) );
  AOI22_X1 U11566 ( .A1(n10526), .A2(n10522), .B1(n10521), .B2(n10523), .ZN(
        P2_U3526) );
  AOI22_X1 U11567 ( .A1(n10526), .A2(n10525), .B1(n10524), .B2(n10523), .ZN(
        P2_U3527) );
  INV_X1 U11568 ( .A(n10527), .ZN(n10528) );
  NAND2_X1 U11569 ( .A1(n10529), .A2(n10528), .ZN(n10530) );
  XOR2_X1 U11570 ( .A(n10531), .B(n10530), .Z(ADD_1071_U5) );
  XOR2_X1 U11571 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11572 ( .B1(n10534), .B2(n10533), .A(n10532), .ZN(ADD_1071_U56) );
  OAI21_X1 U11573 ( .B1(n10537), .B2(n10536), .A(n10535), .ZN(ADD_1071_U57) );
  OAI21_X1 U11574 ( .B1(n10540), .B2(n10539), .A(n10538), .ZN(ADD_1071_U58) );
  OAI21_X1 U11575 ( .B1(n10543), .B2(n10542), .A(n10541), .ZN(ADD_1071_U59) );
  OAI21_X1 U11576 ( .B1(n10546), .B2(n10545), .A(n10544), .ZN(ADD_1071_U60) );
  OAI21_X1 U11577 ( .B1(n10549), .B2(n10548), .A(n10547), .ZN(ADD_1071_U61) );
  AOI21_X1 U11578 ( .B1(n10552), .B2(n10551), .A(n10550), .ZN(ADD_1071_U62) );
  AOI21_X1 U11579 ( .B1(n10555), .B2(n10554), .A(n10553), .ZN(ADD_1071_U63) );
  XOR2_X1 U11580 ( .A(n10556), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  XOR2_X1 U11581 ( .A(n10557), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11582 ( .A1(n10559), .A2(n10558), .ZN(n10560) );
  XOR2_X1 U11583 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10560), .Z(ADD_1071_U51) );
  AOI222_X1 U11584 ( .A1(n10565), .A2(n10564), .B1(n10565), .B2(n10563), .C1(
        n10562), .C2(n10561), .ZN(ADD_1071_U47) );
  OAI21_X1 U11585 ( .B1(n10568), .B2(n10567), .A(n10566), .ZN(n10569) );
  XNOR2_X1 U11586 ( .A(n10569), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U11587 ( .A(n10571), .B(n10570), .Z(ADD_1071_U54) );
  XOR2_X1 U11588 ( .A(n10572), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  XOR2_X1 U11589 ( .A(n10574), .B(n10573), .Z(ADD_1071_U53) );
  XNOR2_X1 U11590 ( .A(n10576), .B(n10575), .ZN(ADD_1071_U52) );
  XNOR2_X1 U7859 ( .A(n6117), .B(n6116), .ZN(n6574) );
  INV_X1 U4919 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6914) );
  CLKBUF_X1 U4938 ( .A(n9025), .Z(n4511) );
  CLKBUF_X1 U5384 ( .A(n6258), .Z(n7172) );
  CLKBUF_X1 U5913 ( .A(n6198), .Z(n9124) );
endmodule

