

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4264, n4265, n4266, n4267, n4268, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10007;

  INV_X1 U4766 ( .A(P2_STATE_REG_SCAN_IN), .ZN(n10007) );
  OR2_X1 U4767 ( .A1(n9693), .A2(n6934), .ZN(n9683) );
  AND3_X1 U4768 ( .A1(n4953), .A2(n4952), .A3(n4951), .ZN(n9920) );
  CLKBUF_X2 U4769 ( .A(n4940), .Z(n4266) );
  CLKBUF_X2 U4770 ( .A(n4940), .Z(n8231) );
  OAI21_X1 U4771 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        n4868), .ZN(n4656) );
  INV_X1 U4774 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U4775 ( .A(n8393), .ZN(n8385) );
  INV_X1 U4776 ( .A(n8999), .ZN(n5709) );
  INV_X1 U4777 ( .A(n4869), .ZN(n4940) );
  NAND2_X1 U4778 ( .A1(n4478), .A2(n4477), .ZN(n8363) );
  NAND2_X1 U4780 ( .A1(n6167), .A2(n5561), .ZN(n5665) );
  NAND2_X1 U4781 ( .A1(n7344), .A2(n5147), .ZN(n7352) );
  INV_X1 U4782 ( .A(n8239), .ZN(n5481) );
  AND2_X1 U4783 ( .A1(n8609), .A2(n8608), .ZN(n8611) );
  AND3_X1 U4784 ( .A1(n4930), .A2(n4929), .A3(n4928), .ZN(n6915) );
  NAND2_X1 U4785 ( .A1(n8285), .A2(n8279), .ZN(n8408) );
  INV_X1 U4786 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8964) );
  AND2_X1 U4787 ( .A1(n4716), .A2(n4318), .ZN(n9074) );
  AND2_X1 U4788 ( .A1(n7941), .A2(n7940), .ZN(n4640) );
  OAI21_X1 U4789 ( .B1(n5195), .B2(n5194), .A(n5198), .ZN(n5222) );
  NAND3_X1 U4790 ( .A1(n4517), .A2(n7159), .A3(n4516), .ZN(n7344) );
  XNOR2_X1 U4791 ( .A(n4363), .B(n5029), .ZN(n6315) );
  INV_X1 U4792 ( .A(n8583), .ZN(n8569) );
  INV_X2 U4793 ( .A(n8688), .ZN(n7135) );
  NAND2_X1 U4794 ( .A1(n4543), .A2(n4540), .ZN(n8441) );
  XNOR2_X1 U4795 ( .A(n5573), .B(n5572), .ZN(n7939) );
  AND4_X2 U4796 ( .A1(n4353), .A2(n5547), .A3(n5546), .A4(n5785), .ZN(n4264)
         );
  NOR2_X2 U4797 ( .A1(n8557), .A2(n8079), .ZN(n8547) );
  NAND2_X2 U4798 ( .A1(n5175), .A2(n4840), .ZN(n5177) );
  OR2_X2 U4799 ( .A1(n6726), .A2(n9725), .ZN(n9722) );
  OAI21_X2 U4800 ( .B1(n5153), .B2(n5152), .A(n5154), .ZN(n5175) );
  NAND2_X2 U4801 ( .A1(n4500), .A2(n4503), .ZN(n5153) );
  INV_X2 U4802 ( .A(n8283), .ZN(n4267) );
  OAI211_X2 U4803 ( .C1(n6167), .C2(n6364), .A(n5706), .B(n5705), .ZN(n6934)
         );
  INV_X4 U4805 ( .A(n6055), .ZN(n9001) );
  INV_X1 U4806 ( .A(n8444), .ZN(n8241) );
  OAI21_X2 U4807 ( .B1(n7520), .B2(n7522), .A(n7519), .ZN(n7521) );
  NAND2_X2 U4808 ( .A1(n7440), .A2(n7439), .ZN(n7520) );
  OAI21_X2 U4809 ( .B1(n7521), .B2(n4779), .A(n4776), .ZN(n7641) );
  OR2_X1 U4810 ( .A1(n6112), .A2(n6113), .ZN(n4362) );
  NAND2_X1 U4811 ( .A1(n8520), .A2(n8527), .ZN(n8519) );
  NAND2_X1 U4812 ( .A1(n5933), .A2(n5932), .ZN(n7661) );
  NAND2_X1 U4813 ( .A1(n5922), .A2(n5923), .ZN(n7619) );
  OAI21_X1 U4814 ( .B1(n5868), .B2(n4731), .A(n4730), .ZN(n5922) );
  NAND2_X1 U4815 ( .A1(n5383), .A2(n5382), .ZN(n5413) );
  CLKBUF_X2 U4816 ( .A(n5709), .Z(n6105) );
  NAND4_X1 U4817 ( .A1(n5740), .A2(n5739), .A3(n5738), .A4(n5737), .ZN(n9676)
         );
  NAND2_X1 U4818 ( .A1(n8274), .A2(n8275), .ZN(n8402) );
  NAND2_X1 U4819 ( .A1(n8464), .A2(n9916), .ZN(n8275) );
  AND2_X1 U4821 ( .A1(n4414), .A2(n5636), .ZN(n6714) );
  NAND2_X2 U4822 ( .A1(n8241), .A2(n8436), .ZN(n8399) );
  INV_X4 U4823 ( .A(n6167), .ZN(n5635) );
  XNOR2_X1 U4824 ( .A(n5487), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8444) );
  AOI21_X1 U4825 ( .B1(n8087), .B2(n8659), .A(n8086), .ZN(n8723) );
  OAI21_X1 U4826 ( .B1(n4474), .B2(n4283), .A(n4471), .ZN(n8094) );
  NOR2_X1 U4827 ( .A1(n8066), .A2(n4330), .ZN(n4766) );
  NAND2_X1 U4828 ( .A1(n8066), .A2(n4330), .ZN(n4767) );
  INV_X1 U4829 ( .A(n9459), .ZN(n5868) );
  NAND2_X1 U4830 ( .A1(n8363), .A2(n8364), .ZN(n8594) );
  NOR2_X1 U4831 ( .A1(n8324), .A2(n8325), .ZN(n4432) );
  OAI21_X1 U4832 ( .B1(n5371), .B2(n5370), .A(n5372), .ZN(n5381) );
  MUX2_X1 U4833 ( .A(n8323), .B(n8322), .S(n8393), .Z(n8324) );
  NAND2_X1 U4834 ( .A1(n7798), .A2(n7909), .ZN(n7794) );
  NAND2_X1 U4835 ( .A1(n5897), .A2(n5896), .ZN(n9421) );
  NAND2_X1 U4836 ( .A1(n5162), .A2(n5161), .ZN(n7438) );
  NAND2_X1 U4837 ( .A1(n5177), .A2(n5176), .ZN(n5195) );
  INV_X2 U4838 ( .A(n9737), .ZN(n9739) );
  NAND2_X1 U4839 ( .A1(n5016), .A2(n5015), .ZN(n6767) );
  OAI211_X1 U4840 ( .C1(n6167), .C2(n6394), .A(n5764), .B(n5763), .ZN(n7179)
         );
  NAND2_X1 U4841 ( .A1(n5789), .A2(n5788), .ZN(n7315) );
  INV_X1 U4842 ( .A(n7130), .ZN(n9926) );
  NAND2_X1 U4843 ( .A1(n4602), .A2(n4600), .ZN(n7130) );
  OR2_X1 U4844 ( .A1(n5297), .A2(n8117), .ZN(n5316) );
  OAI21_X1 U4845 ( .B1(n5056), .B2(n5055), .A(n5057), .ZN(n5079) );
  AND2_X2 U4846 ( .A1(n5625), .A2(n5592), .ZN(n8996) );
  INV_X1 U4847 ( .A(n5643), .ZN(n6055) );
  INV_X2 U4848 ( .A(n6715), .ZN(n6713) );
  NAND4_X1 U4849 ( .A1(n5779), .A2(n5778), .A3(n5777), .A4(n5776), .ZN(n9122)
         );
  NAND4_X1 U4850 ( .A1(n5680), .A2(n5679), .A3(n5678), .A4(n5677), .ZN(n9125)
         );
  AND2_X2 U4851 ( .A1(n6371), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  CLKBUF_X1 U4852 ( .A(n6133), .Z(n8041) );
  CLKBUF_X1 U4853 ( .A(n6132), .Z(n8043) );
  INV_X1 U4854 ( .A(n6132), .ZN(n6134) );
  NAND4_X1 U4855 ( .A1(n4914), .A2(n4913), .A3(n4912), .A4(n4911), .ZN(n8464)
         );
  AND2_X2 U4856 ( .A1(n4610), .A2(n4609), .ZN(n5482) );
  NAND4_X1 U4857 ( .A1(n4886), .A2(n4885), .A3(n4884), .A4(n4883), .ZN(n8465)
         );
  NAND4_X1 U4858 ( .A1(n4890), .A2(n4889), .A3(n4888), .A4(n4887), .ZN(n8467)
         );
  BUF_X2 U4859 ( .A(n4954), .Z(n6328) );
  BUF_X2 U4860 ( .A(n4972), .Z(n6329) );
  INV_X1 U4861 ( .A(n5602), .ZN(n7701) );
  AND2_X2 U4862 ( .A1(n4882), .A2(n8973), .ZN(n4954) );
  NAND2_X1 U4863 ( .A1(n4900), .A2(n4899), .ZN(n4920) );
  NAND2_X1 U4864 ( .A1(n5581), .A2(n5582), .ZN(n7358) );
  XNOR2_X1 U4865 ( .A(n5558), .B(P1_IR_REG_28__SCAN_IN), .ZN(n6140) );
  OAI21_X1 U4866 ( .B1(n4851), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5487) );
  INV_X1 U4867 ( .A(n5597), .ZN(n5598) );
  NAND2_X1 U4868 ( .A1(n9443), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U4869 ( .A1(n5589), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5591) );
  OAI21_X1 U4870 ( .B1(n5951), .B2(n4271), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5573) );
  NOR2_X1 U4871 ( .A1(n4542), .A2(n4541), .ZN(n4540) );
  AND2_X1 U4872 ( .A1(n5110), .A2(n5109), .ZN(n5140) );
  NAND2_X1 U4873 ( .A1(n4867), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4865) );
  NAND2_X1 U4874 ( .A1(n4866), .A2(n4376), .ZN(n4543) );
  NOR2_X1 U4875 ( .A1(n5067), .A2(n5066), .ZN(n5110) );
  OR2_X1 U4876 ( .A1(n5002), .A2(n5001), .ZN(n5044) );
  AND2_X1 U4877 ( .A1(n4264), .A2(n5556), .ZN(n4551) );
  NAND2_X1 U4878 ( .A1(n4658), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4657) );
  INV_X1 U4879 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5724) );
  INV_X1 U4880 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4868) );
  CLKBUF_X1 U4881 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n9556) );
  INV_X1 U4882 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5545) );
  NOR2_X2 U4883 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5660) );
  NOR2_X1 U4884 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5565) );
  INV_X1 U4885 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5547) );
  NOR2_X1 U4886 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4541) );
  NOR2_X1 U4887 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n4740) );
  NOR2_X1 U4888 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4739) );
  NOR2_X1 U4889 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4842) );
  NOR2_X2 U4890 ( .A1(n5554), .A2(n5553), .ZN(n5555) );
  AND2_X1 U4891 ( .A1(n5625), .A2(n5592), .ZN(n4268) );
  AND2_X1 U4892 ( .A1(n5410), .A2(n4475), .ZN(n4474) );
  AND2_X2 U4893 ( .A1(n8047), .A2(n7701), .ZN(n5676) );
  XNOR2_X1 U4894 ( .A(n9727), .B(n6718), .ZN(n6922) );
  INV_X2 U4895 ( .A(n6936), .ZN(n6718) );
  OAI222_X1 U4896 ( .A1(n8048), .A2(n8092), .B1(P1_U3084), .B2(n8047), .C1(
        n8046), .C2(n8045), .ZN(P1_U3323) );
  AND2_X4 U4897 ( .A1(n8047), .A2(n5602), .ZN(n5675) );
  INV_X1 U4899 ( .A(n5663), .ZN(n4270) );
  NAND2_X4 U4900 ( .A1(n6167), .A2(n7715), .ZN(n5663) );
  XNOR2_X2 U4901 ( .A(n4874), .B(P2_IR_REG_1__SCAN_IN), .ZN(n6212) );
  AOI21_X1 U4902 ( .B1(n9310), .B2(n4683), .A(n8003), .ZN(n4395) );
  INV_X1 U4903 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n4844) );
  NAND2_X1 U4904 ( .A1(n5246), .A2(n4859), .ZN(n4849) );
  NAND2_X1 U4905 ( .A1(n5935), .A2(n5566), .ZN(n5951) );
  NAND2_X1 U4906 ( .A1(n8375), .A2(n8385), .ZN(n4465) );
  AOI21_X1 U4907 ( .B1(n8732), .B2(n8563), .A(n8385), .ZN(n4466) );
  OR2_X1 U4908 ( .A1(n8759), .A2(n8104), .ZN(n8076) );
  NOR2_X1 U4909 ( .A1(n9032), .A2(n4297), .ZN(n4718) );
  INV_X1 U4910 ( .A(n9063), .ZN(n4719) );
  INV_X1 U4911 ( .A(n4628), .ZN(n4627) );
  OAI21_X1 U4912 ( .B1(n5516), .B2(n4629), .A(n7694), .ZN(n4628) );
  NOR2_X1 U4913 ( .A1(n4505), .A2(n4502), .ZN(n4501) );
  INV_X1 U4914 ( .A(n5080), .ZN(n4502) );
  INV_X1 U4915 ( .A(n4506), .ZN(n4505) );
  AND2_X1 U4916 ( .A1(n5024), .A2(n5028), .ZN(n5030) );
  OAI21_X1 U4917 ( .B1(n5561), .B2(n4361), .A(n4360), .ZN(n5023) );
  NAND2_X1 U4918 ( .A1(n5561), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n4360) );
  OR2_X1 U4919 ( .A1(n5475), .A2(n5474), .ZN(n5526) );
  NAND2_X1 U4920 ( .A1(n4287), .A2(n8363), .ZN(n4593) );
  NAND2_X1 U4921 ( .A1(n8594), .A2(n4760), .ZN(n4759) );
  INV_X1 U4922 ( .A(n4761), .ZN(n4760) );
  OR2_X1 U4923 ( .A1(n8783), .A2(n8155), .ZN(n8339) );
  OR2_X1 U4924 ( .A1(n8465), .A2(n6884), .ZN(n6585) );
  INV_X1 U4925 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4859) );
  NOR2_X2 U4926 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4903) );
  AND2_X1 U4927 ( .A1(n7727), .A2(n7930), .ZN(n7898) );
  INV_X1 U4928 ( .A(n8027), .ZN(n4832) );
  OR2_X1 U4929 ( .A1(n9351), .A2(n9009), .ZN(n8028) );
  OR2_X1 U4930 ( .A1(n9360), .A2(n9105), .ZN(n8024) );
  NOR2_X1 U4931 ( .A1(n9235), .A2(n4794), .ZN(n4793) );
  OR2_X1 U4932 ( .A1(n9377), .A2(n9382), .ZN(n4567) );
  AND2_X1 U4933 ( .A1(n5746), .A2(n4678), .ZN(n7089) );
  AND2_X1 U4934 ( .A1(n5745), .A2(n4679), .ZN(n4678) );
  NAND2_X1 U4935 ( .A1(n5635), .A2(n6383), .ZN(n4679) );
  OR2_X2 U4936 ( .A1(n6133), .A2(n7940), .ZN(n6723) );
  NOR2_X1 U4937 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n4812) );
  INV_X1 U4938 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5556) );
  OAI21_X1 U4939 ( .B1(n5308), .B2(n5307), .A(n5309), .ZN(n5326) );
  AND2_X1 U4940 ( .A1(n5327), .A2(n5313), .ZN(n5325) );
  AND2_X1 U4941 ( .A1(n5244), .A2(n5227), .ZN(n5242) );
  NAND2_X1 U4942 ( .A1(n6837), .A2(n4617), .ZN(n6761) );
  AND2_X1 U4943 ( .A1(n5021), .A2(n4999), .ZN(n4617) );
  NAND2_X1 U4944 ( .A1(n9472), .A2(n5211), .ZN(n7543) );
  INV_X1 U4945 ( .A(n5532), .ZN(n5463) );
  AND4_X1 U4946 ( .A1(n5168), .A2(n5167), .A3(n5166), .A4(n5165), .ZN(n7434)
         );
  AND4_X1 U4947 ( .A1(n5095), .A2(n5094), .A3(n5093), .A4(n5092), .ZN(n8180)
         );
  AND2_X1 U4949 ( .A1(n8091), .A2(n8973), .ZN(n4972) );
  AND2_X1 U4950 ( .A1(n8091), .A2(n4881), .ZN(n4973) );
  AND2_X1 U4951 ( .A1(n4882), .A2(n4881), .ZN(n5443) );
  NOR2_X1 U4952 ( .A1(n8473), .A2(n8480), .ZN(n8492) );
  NAND2_X1 U4953 ( .A1(n8535), .A2(n8060), .ZN(n8520) );
  OR2_X1 U4954 ( .A1(n8732), .A2(n8530), .ZN(n8060) );
  OR2_X1 U4955 ( .A1(n8747), .A2(n4477), .ZN(n8058) );
  AOI21_X1 U4956 ( .B1(n4778), .B2(n4777), .A(n4304), .ZN(n4776) );
  INV_X1 U4957 ( .A(n8422), .ZN(n4777) );
  NOR2_X1 U4958 ( .A1(n8422), .A2(n4596), .ZN(n4595) );
  INV_X1 U4959 ( .A(n7523), .ZN(n4596) );
  INV_X1 U4960 ( .A(n4573), .ZN(n4572) );
  AND2_X1 U4961 ( .A1(n8301), .A2(n4570), .ZN(n4569) );
  INV_X2 U4962 ( .A(n6195), .ZN(n5294) );
  AND2_X1 U4963 ( .A1(n4863), .A2(n4327), .ZN(n4780) );
  INV_X1 U4964 ( .A(n4783), .ZN(n4782) );
  INV_X1 U4965 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4877) );
  NAND2_X1 U4966 ( .A1(n5488), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5513) );
  INV_X1 U4967 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4860) );
  AND2_X1 U4968 ( .A1(n5178), .A2(n4323), .ZN(n5246) );
  NAND2_X1 U4969 ( .A1(n5838), .A2(n5837), .ZN(n7388) );
  AND2_X1 U4970 ( .A1(n7939), .A2(n9137), .ZN(n7977) );
  NAND2_X1 U4971 ( .A1(n7970), .A2(n7890), .ZN(n8030) );
  NAND2_X1 U4972 ( .A1(n4785), .A2(n4787), .ZN(n9218) );
  AOI21_X1 U4973 ( .B1(n4789), .B2(n4792), .A(n4788), .ZN(n4787) );
  AOI21_X1 U4974 ( .B1(n4392), .B2(n4394), .A(n4308), .ZN(n4391) );
  NAND2_X1 U4975 ( .A1(n9397), .A2(n9114), .ZN(n4683) );
  INV_X2 U4976 ( .A(n5665), .ZN(n7777) );
  NAND2_X1 U4977 ( .A1(n6730), .A2(n6729), .ZN(n9704) );
  AND2_X1 U4978 ( .A1(n4736), .A2(n4837), .ZN(n5935) );
  NOR2_X1 U4979 ( .A1(n4738), .A2(n4306), .ZN(n4736) );
  NAND2_X1 U4980 ( .A1(n5525), .A2(n5524), .ZN(n8725) );
  NAND2_X1 U4981 ( .A1(n4450), .A2(n4447), .ZN(n8265) );
  NAND2_X1 U4982 ( .A1(n8251), .A2(n8393), .ZN(n4450) );
  NAND2_X1 U4983 ( .A1(n8267), .A2(n4302), .ZN(n4447) );
  OR2_X1 U4984 ( .A1(n4441), .A2(n4437), .ZN(n4436) );
  NOR2_X1 U4985 ( .A1(n8324), .A2(n4442), .ZN(n4440) );
  INV_X1 U4986 ( .A(n8321), .ZN(n4437) );
  NOR2_X1 U4987 ( .A1(n4349), .A2(n4305), .ZN(n4348) );
  INV_X1 U4988 ( .A(n7829), .ZN(n4349) );
  NOR2_X1 U4989 ( .A1(n8355), .A2(n4457), .ZN(n4456) );
  AND2_X1 U4990 ( .A1(n8343), .A2(n8393), .ZN(n4457) );
  AND2_X1 U4991 ( .A1(n4452), .A2(n4451), .ZN(n8361) );
  NAND2_X1 U4992 ( .A1(n4467), .A2(n8374), .ZN(n8377) );
  NAND2_X1 U4993 ( .A1(n7920), .A2(n7745), .ZN(n4817) );
  INV_X1 U4994 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n5155) );
  NAND2_X1 U4995 ( .A1(n8747), .A2(n8165), .ZN(n8364) );
  NOR3_X1 U4996 ( .A1(n8676), .A2(n8618), .A3(n4417), .ZN(n4550) );
  NOR2_X1 U4997 ( .A1(n8764), .A2(n8771), .ZN(n4418) );
  NOR2_X1 U4998 ( .A1(n8072), .A2(n4585), .ZN(n4584) );
  INV_X1 U4999 ( .A(n8331), .ZN(n4585) );
  OR2_X1 U5000 ( .A1(n8795), .A2(n7552), .ZN(n4421) );
  NAND2_X1 U5001 ( .A1(n5212), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5232) );
  INV_X1 U5002 ( .A(n7238), .ZN(n4753) );
  AND2_X1 U5003 ( .A1(n4267), .A2(n8285), .ZN(n4576) );
  NAND2_X1 U5004 ( .A1(n8461), .A2(n6995), .ZN(n8249) );
  OR2_X1 U5005 ( .A1(n6995), .A2(n8461), .ZN(n8267) );
  NAND2_X1 U5006 ( .A1(n8675), .A2(n8052), .ZN(n4775) );
  INV_X1 U5007 ( .A(n9096), .ZN(n4705) );
  OR2_X1 U5008 ( .A1(n6001), .A2(n6000), .ZN(n6002) );
  AOI21_X1 U5009 ( .B1(n4718), .B2(n4720), .A(n4337), .ZN(n4717) );
  INV_X1 U5010 ( .A(n9065), .ZN(n4720) );
  OAI21_X1 U5011 ( .B1(n7686), .B2(n4724), .A(n4721), .ZN(n4729) );
  AOI21_X1 U5012 ( .B1(n4723), .B2(n4722), .A(n4316), .ZN(n4721) );
  INV_X1 U5013 ( .A(n4728), .ZN(n4722) );
  NAND2_X1 U5014 ( .A1(n4293), .A2(n7895), .ZN(n4370) );
  NOR2_X1 U5015 ( .A1(n7966), .A2(n8030), .ZN(n4654) );
  OR2_X1 U5016 ( .A1(n9337), .A2(n7788), .ZN(n7890) );
  NOR2_X1 U5017 ( .A1(n9177), .A2(n4829), .ZN(n4828) );
  INV_X1 U5018 ( .A(n8026), .ZN(n4829) );
  INV_X1 U5019 ( .A(n4807), .ZN(n4801) );
  OR2_X1 U5020 ( .A1(n9382), .A2(n9250), .ZN(n7903) );
  NOR2_X1 U5021 ( .A1(n9283), .A2(n4808), .ZN(n4807) );
  INV_X1 U5022 ( .A(n4674), .ZN(n4672) );
  OR2_X1 U5023 ( .A1(n7669), .A2(n7690), .ZN(n7761) );
  OR2_X1 U5024 ( .A1(n7560), .A2(n9512), .ZN(n7827) );
  AND2_X1 U5025 ( .A1(n7055), .A2(n7738), .ZN(n7744) );
  NAND2_X1 U5026 ( .A1(n4559), .A2(n5561), .ZN(n4413) );
  INV_X1 U5027 ( .A(n6292), .ZN(n4559) );
  NAND2_X1 U5028 ( .A1(n7715), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4412) );
  OR2_X1 U5029 ( .A1(n9345), .A2(n9179), .ZN(n7900) );
  OR3_X1 U5030 ( .A1(n4562), .A2(n9421), .A3(n9410), .ZN(n4561) );
  NOR3_X1 U5031 ( .A1(n7569), .A2(n9421), .A3(n9499), .ZN(n7584) );
  XNOR2_X1 U5032 ( .A(n7709), .B(n7710), .ZN(n7720) );
  NAND2_X1 U5033 ( .A1(n4625), .A2(n4623), .ZN(n7705) );
  AOI21_X1 U5034 ( .B1(n4627), .B2(n4629), .A(n4624), .ZN(n4623) );
  INV_X1 U5035 ( .A(n7696), .ZN(n4624) );
  INV_X1 U5036 ( .A(n5450), .ZN(n4632) );
  NAND2_X1 U5037 ( .A1(n5290), .A2(n5289), .ZN(n5308) );
  NAND2_X1 U5038 ( .A1(n5287), .A2(n5286), .ZN(n5290) );
  INV_X1 U5039 ( .A(n5285), .ZN(n5286) );
  INV_X1 U5040 ( .A(n4738), .ZN(n4737) );
  AOI21_X1 U5041 ( .B1(n4504), .B2(n4506), .A(n4311), .ZN(n4503) );
  AOI21_X1 U5042 ( .B1(n5027), .B2(n5026), .A(n4313), .ZN(n5056) );
  NAND2_X1 U5043 ( .A1(n5028), .A2(n5029), .ZN(n5034) );
  NAND2_X1 U5044 ( .A1(n4986), .A2(n4985), .ZN(n5027) );
  INV_X1 U5045 ( .A(n4945), .ZN(n4498) );
  OAI21_X1 U5046 ( .B1(n5561), .B2(P1_DATAO_REG_4__SCAN_IN), .A(n4366), .ZN(
        n4965) );
  NAND2_X1 U5047 ( .A1(n5561), .A2(n6298), .ZN(n4366) );
  NOR2_X2 U5048 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5544) );
  NAND2_X1 U5049 ( .A1(n5617), .A2(n4872), .ZN(n4898) );
  INV_X1 U5050 ( .A(n8215), .ZN(n4472) );
  INV_X1 U5051 ( .A(n5409), .ZN(n4470) );
  NAND2_X1 U5052 ( .A1(n5356), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5400) );
  NAND2_X1 U5053 ( .A1(n9471), .A2(n5189), .ZN(n9472) );
  AND2_X1 U5054 ( .A1(n5100), .A2(n5078), .ZN(n4619) );
  AOI21_X1 U5055 ( .B1(n4619), .B2(n4520), .A(n4519), .ZN(n4518) );
  INV_X1 U5056 ( .A(n5101), .ZN(n4519) );
  INV_X1 U5057 ( .A(n5074), .ZN(n4520) );
  XNOR2_X1 U5058 ( .A(n5482), .B(n6884), .ZN(n6842) );
  INV_X1 U5059 ( .A(n5264), .ZN(n4511) );
  AOI21_X1 U5060 ( .B1(n8397), .B2(n8398), .A(n8396), .ZN(n8435) );
  AOI21_X1 U5061 ( .B1(n8435), .B2(n8434), .A(n5535), .ZN(n4446) );
  AND4_X1 U5062 ( .A1(n5007), .A2(n5006), .A3(n5005), .A4(n5004), .ZN(n6825)
         );
  AND4_X1 U5063 ( .A1(n4994), .A2(n4993), .A3(n4992), .A4(n4991), .ZN(n6751)
         );
  NOR2_X1 U5064 ( .A1(n6204), .A2(n4292), .ZN(n6239) );
  OR2_X1 U5065 ( .A1(n6239), .A2(n6238), .ZN(n4537) );
  OR2_X1 U5066 ( .A1(n6278), .A2(n6277), .ZN(n4530) );
  AND2_X1 U5067 ( .A1(n4530), .A2(n4529), .ZN(n6210) );
  NAND2_X1 U5068 ( .A1(n6216), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4529) );
  OR2_X1 U5069 ( .A1(n6210), .A2(n6209), .ZN(n4528) );
  NOR2_X1 U5070 ( .A1(n7211), .A2(n7210), .ZN(n4525) );
  AOI21_X1 U5071 ( .B1(n7206), .B2(n7207), .A(n7205), .ZN(n7211) );
  NOR2_X1 U5072 ( .A1(n8522), .A2(n8720), .ZN(n8513) );
  NAND2_X1 U5073 ( .A1(n8582), .A2(n8067), .ZN(n8565) );
  NOR2_X1 U5074 ( .A1(n8565), .A2(n8732), .ZN(n8539) );
  AND2_X1 U5075 ( .A1(n5468), .A2(n5467), .ZN(n8563) );
  OR2_X1 U5076 ( .A1(n8542), .A2(n5463), .ZN(n5468) );
  AOI21_X1 U5077 ( .B1(n4591), .B2(n8078), .A(n4590), .ZN(n4589) );
  INV_X1 U5078 ( .A(n8371), .ZN(n4590) );
  OR2_X1 U5079 ( .A1(n8611), .A2(n4592), .ZN(n4588) );
  AND2_X1 U5080 ( .A1(n4588), .A2(n4586), .ZN(n8557) );
  AND2_X1 U5081 ( .A1(n4589), .A2(n4587), .ZN(n4586) );
  INV_X1 U5082 ( .A(n8558), .ZN(n4587) );
  NAND2_X1 U5083 ( .A1(n4759), .A2(n8058), .ZN(n4757) );
  AND2_X1 U5084 ( .A1(n8618), .A2(n8634), .ZN(n4761) );
  OR2_X1 U5085 ( .A1(n8607), .A2(n4759), .ZN(n8593) );
  OR2_X1 U5086 ( .A1(n8611), .A2(n4287), .ZN(n4594) );
  NAND2_X1 U5087 ( .A1(n8077), .A2(n8075), .ZN(n4606) );
  AOI21_X1 U5088 ( .B1(n8077), .B2(n4605), .A(n8246), .ZN(n4604) );
  OR2_X1 U5089 ( .A1(n8771), .A2(n8126), .ZN(n8352) );
  AOI21_X1 U5090 ( .B1(n4772), .B2(n4771), .A(n4332), .ZN(n4770) );
  INV_X1 U5091 ( .A(n8052), .ZN(n4771) );
  NOR2_X1 U5092 ( .A1(n8676), .A2(n8771), .ZN(n8668) );
  AND2_X1 U5093 ( .A1(n8352), .A2(n8075), .ZN(n8660) );
  INV_X1 U5094 ( .A(n4584), .ZN(n4583) );
  INV_X1 U5095 ( .A(n7634), .ZN(n7635) );
  AOI21_X1 U5096 ( .B1(n4584), .B2(n4582), .A(n4581), .ZN(n4580) );
  INV_X1 U5097 ( .A(n8345), .ZN(n4581) );
  OR2_X1 U5098 ( .A1(n8695), .A2(n8778), .ZN(n8676) );
  AND2_X1 U5099 ( .A1(n8348), .A2(n8346), .ZN(n8674) );
  OR2_X1 U5100 ( .A1(n8787), .A2(n8203), .ZN(n8331) );
  NAND2_X1 U5101 ( .A1(n7635), .A2(n7640), .ZN(n8071) );
  NOR2_X1 U5102 ( .A1(n8421), .A2(n4599), .ZN(n4598) );
  INV_X1 U5103 ( .A(n8315), .ZN(n4599) );
  AOI21_X1 U5104 ( .B1(n4752), .B2(n4751), .A(n4756), .ZN(n4750) );
  NOR2_X1 U5105 ( .A1(n7361), .A2(n8456), .ZN(n4756) );
  INV_X1 U5106 ( .A(n8414), .ZN(n4751) );
  AND2_X1 U5107 ( .A1(n8416), .A2(n8417), .ZN(n7365) );
  NOR2_X1 U5108 ( .A1(n4575), .A2(n7239), .ZN(n4573) );
  NAND2_X1 U5109 ( .A1(n7073), .A2(n8411), .ZN(n4574) );
  CLKBUF_X1 U5110 ( .A(n7247), .Z(n4371) );
  AND2_X1 U5111 ( .A1(n8298), .A2(n8300), .ZN(n8413) );
  AND2_X1 U5112 ( .A1(n8296), .A2(n8294), .ZN(n8411) );
  NOR2_X1 U5113 ( .A1(n4267), .A2(n4372), .ZN(n4746) );
  NOR2_X1 U5114 ( .A1(n8408), .A2(n4747), .ZN(n4372) );
  INV_X1 U5115 ( .A(n6744), .ZN(n4747) );
  OR2_X1 U5116 ( .A1(n6308), .A2(n4869), .ZN(n4602) );
  NAND2_X1 U5117 ( .A1(n6743), .A2(n6742), .ZN(n7124) );
  NAND2_X1 U5118 ( .A1(n7124), .A2(n8408), .ZN(n7123) );
  AND2_X1 U5119 ( .A1(n6583), .A2(n6995), .ZN(n7126) );
  NAND2_X1 U5120 ( .A1(n6588), .A2(n8405), .ZN(n7013) );
  AOI21_X1 U5121 ( .B1(n6585), .B2(n6889), .A(n4375), .ZN(n7005) );
  INV_X1 U5122 ( .A(n8564), .ZN(n8654) );
  NAND2_X1 U5123 ( .A1(n8240), .A2(n8434), .ZN(n8659) );
  NAND2_X1 U5124 ( .A1(n8233), .A2(n8232), .ZN(n8712) );
  NAND2_X1 U5125 ( .A1(n5272), .A2(n5271), .ZN(n8783) );
  NAND2_X1 U5126 ( .A1(n5500), .A2(n5499), .ZN(n9885) );
  XNOR2_X1 U5127 ( .A(n4878), .B(P2_IR_REG_30__SCAN_IN), .ZN(n4882) );
  NAND2_X1 U5128 ( .A1(n8965), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4878) );
  XNOR2_X1 U5129 ( .A(n4880), .B(P2_IR_REG_29__SCAN_IN), .ZN(n4881) );
  NAND2_X1 U5130 ( .A1(n4460), .A2(n4780), .ZN(n4879) );
  INV_X1 U5131 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5512) );
  XNOR2_X1 U5132 ( .A(n4850), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8255) );
  NAND2_X1 U5133 ( .A1(n5178), .A2(n4522), .ZN(n5228) );
  NOR2_X1 U5134 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n4741) );
  AOI21_X1 U5135 ( .B1(n4409), .B2(P1_IR_REG_31__SCAN_IN), .A(n4314), .ZN(
        n4408) );
  XNOR2_X1 U5136 ( .A(n5733), .B(n5731), .ZN(n6703) );
  INV_X1 U5137 ( .A(n9675), .ZN(n9702) );
  AOI21_X1 U5138 ( .B1(n9728), .B2(n4268), .A(n5624), .ZN(n6433) );
  INV_X1 U5139 ( .A(n7136), .ZN(n4700) );
  AOI21_X1 U5140 ( .B1(n9130), .B2(n9129), .A(n9128), .ZN(n9132) );
  INV_X1 U5141 ( .A(n4828), .ZN(n4827) );
  NAND2_X1 U5142 ( .A1(n4272), .A2(n4832), .ZN(n4824) );
  INV_X1 U5143 ( .A(n9111), .ZN(n9179) );
  NAND2_X1 U5144 ( .A1(n4823), .A2(n4832), .ZN(n4831) );
  INV_X1 U5145 ( .A(n4830), .ZN(n9175) );
  AND2_X1 U5146 ( .A1(n6151), .A2(n6096), .ZN(n9172) );
  NAND2_X1 U5147 ( .A1(n8028), .A2(n7901), .ZN(n9177) );
  INV_X1 U5148 ( .A(n4793), .ZN(n4790) );
  NAND2_X1 U5149 ( .A1(n4278), .A2(n4796), .ZN(n4795) );
  NOR2_X1 U5150 ( .A1(n9243), .A2(n9258), .ZN(n8007) );
  AOI21_X1 U5151 ( .B1(n4395), .B2(n4393), .A(n4309), .ZN(n4392) );
  INV_X1 U5152 ( .A(n4683), .ZN(n4393) );
  INV_X1 U5153 ( .A(n4395), .ZN(n4394) );
  NAND2_X1 U5154 ( .A1(n4806), .A2(n4809), .ZN(n4805) );
  INV_X1 U5155 ( .A(n9283), .ZN(n4806) );
  NAND2_X1 U5156 ( .A1(n9297), .A2(n4807), .ZN(n4804) );
  INV_X1 U5157 ( .A(n8013), .ZN(n4809) );
  AND2_X1 U5158 ( .A1(n7905), .A2(n8013), .ZN(n9310) );
  AOI21_X1 U5159 ( .B1(n7999), .B2(n7998), .A(n4387), .ZN(n9315) );
  AND2_X1 U5160 ( .A1(n9410), .A2(n9115), .ZN(n4387) );
  INV_X1 U5161 ( .A(n4669), .ZN(n4668) );
  OAI21_X1 U5162 ( .B1(n4670), .B2(n4675), .A(n4676), .ZN(n4669) );
  NAND2_X1 U5163 ( .A1(n4677), .A2(n9496), .ZN(n4676) );
  NAND2_X1 U5164 ( .A1(n9499), .A2(n9118), .ZN(n4674) );
  OR2_X1 U5165 ( .A1(n9499), .A2(n9118), .ZN(n4675) );
  NAND2_X1 U5166 ( .A1(n7562), .A2(n7561), .ZN(n9490) );
  OAI22_X1 U5167 ( .A1(n7319), .A2(n4659), .B1(n7382), .B2(n4660), .ZN(n7384)
         );
  NAND2_X1 U5168 ( .A1(n4663), .A2(n7380), .ZN(n4659) );
  INV_X1 U5169 ( .A(n4661), .ZN(n4660) );
  AND2_X1 U5170 ( .A1(n7563), .A2(n7825), .ZN(n9511) );
  OR2_X1 U5171 ( .A1(n7899), .A2(n6141), .ZN(n9699) );
  NAND2_X1 U5172 ( .A1(n7196), .A2(n7195), .ZN(n7314) );
  INV_X1 U5173 ( .A(n7091), .ZN(n4682) );
  NAND2_X1 U5174 ( .A1(n4835), .A2(n4833), .ZN(n7948) );
  AOI21_X1 U5175 ( .B1(n4276), .B2(n7058), .A(n4834), .ZN(n4833) );
  NAND2_X1 U5176 ( .A1(n7046), .A2(n7047), .ZN(n7092) );
  INV_X1 U5177 ( .A(n9701), .ZN(n9726) );
  OR2_X1 U5178 ( .A1(n7899), .A2(n6423), .ZN(n9701) );
  NAND2_X1 U5179 ( .A1(n8030), .A2(n4331), .ZN(n4689) );
  INV_X1 U5180 ( .A(n8030), .ZN(n4690) );
  NAND2_X1 U5181 ( .A1(n6092), .A2(n6091), .ZN(n9351) );
  NAND2_X1 U5182 ( .A1(n5972), .A2(n5971), .ZN(n9397) );
  INV_X1 U5183 ( .A(n7669), .ZN(n9414) );
  NAND2_X1 U5184 ( .A1(n5453), .A2(n5452), .ZN(n5517) );
  OAI21_X1 U5185 ( .B1(n5413), .B2(n4633), .A(n4631), .ZN(n5453) );
  INV_X1 U5186 ( .A(n4634), .ZN(n4633) );
  AOI21_X1 U5187 ( .B1(n4634), .B2(n4636), .A(n4632), .ZN(n4631) );
  XNOR2_X1 U5188 ( .A(n5517), .B(n5516), .ZN(n7592) );
  XNOR2_X1 U5189 ( .A(n5451), .B(n5450), .ZN(n7540) );
  NAND2_X1 U5190 ( .A1(n4630), .A2(n4634), .ZN(n5451) );
  NAND2_X1 U5191 ( .A1(n5413), .A2(n4637), .ZN(n4630) );
  AND2_X1 U5192 ( .A1(n5382), .A2(n5377), .ZN(n5380) );
  NAND2_X1 U5193 ( .A1(n4524), .A2(n5327), .ZN(n5345) );
  NAND2_X1 U5194 ( .A1(n4486), .A2(n5244), .ZN(n5269) );
  NAND2_X1 U5195 ( .A1(n4490), .A2(n4646), .ZN(n4486) );
  NAND2_X1 U5196 ( .A1(n5177), .A2(n4491), .ZN(n4490) );
  NAND2_X1 U5197 ( .A1(n4645), .A2(n4650), .ZN(n5243) );
  NAND2_X1 U5198 ( .A1(n5195), .A2(n4652), .ZN(n4645) );
  OR2_X1 U5199 ( .A1(n5660), .A2(n5934), .ZN(n5662) );
  NAND2_X1 U5200 ( .A1(n4481), .A2(n4336), .ZN(n4480) );
  NAND2_X1 U5201 ( .A1(n8725), .A2(n9854), .ZN(n4481) );
  NAND2_X1 U5202 ( .A1(n5219), .A2(n7544), .ZN(n4513) );
  AND4_X1 U5203 ( .A1(n5237), .A2(n5236), .A3(n5235), .A4(n5234), .ZN(n8154)
         );
  AND4_X1 U5204 ( .A1(n5145), .A2(n5144), .A3(n5143), .A4(n5142), .ZN(n7328)
         );
  NAND2_X1 U5205 ( .A1(n4995), .A2(n6831), .ZN(n6837) );
  NAND2_X1 U5206 ( .A1(n5538), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9860) );
  INV_X1 U5207 ( .A(n9835), .ZN(n9845) );
  NAND2_X1 U5208 ( .A1(n6329), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8084) );
  NAND2_X1 U5209 ( .A1(n6695), .A2(n6696), .ZN(n6789) );
  OR2_X1 U5210 ( .A1(n4295), .A2(n8492), .ZN(n8474) );
  AND2_X1 U5211 ( .A1(n6187), .A2(n6186), .ZN(n9879) );
  OAI21_X1 U5212 ( .B1(n8506), .B2(n8507), .A(n8505), .ZN(n4532) );
  INV_X1 U5213 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8507) );
  NAND2_X1 U5214 ( .A1(n9886), .A2(n6879), .ZN(n8679) );
  OR2_X1 U5215 ( .A1(n4852), .A2(n4860), .ZN(n4853) );
  OAI21_X1 U5216 ( .B1(n4849), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n4852) );
  NAND2_X1 U5217 ( .A1(n9053), .A2(n4714), .ZN(n4365) );
  INV_X1 U5218 ( .A(n9038), .ZN(n4364) );
  NAND2_X1 U5219 ( .A1(n6061), .A2(n6060), .ZN(n9360) );
  NAND2_X1 U5220 ( .A1(n6031), .A2(n6030), .ZN(n9377) );
  OR2_X1 U5221 ( .A1(n9026), .A2(n9799), .ZN(n9095) );
  AND3_X1 U5222 ( .A1(n6145), .A2(n9799), .A3(n7899), .ZN(n9086) );
  INV_X1 U5223 ( .A(n9095), .ZN(n9107) );
  OAI21_X1 U5224 ( .B1(n9632), .B2(n4868), .A(n9140), .ZN(n4357) );
  AOI21_X1 U5225 ( .B1(n9448), .B2(n7777), .A(n7719), .ZN(n9145) );
  INV_X1 U5226 ( .A(n9351), .ZN(n9174) );
  NAND2_X1 U5227 ( .A1(n9343), .A2(n4403), .ZN(n4401) );
  NAND2_X1 U5228 ( .A1(n4404), .A2(n4690), .ZN(n4403) );
  NOR2_X1 U5229 ( .A1(n4400), .A2(n9823), .ZN(n4398) );
  NOR2_X1 U5230 ( .A1(n9342), .A2(n4335), .ZN(n4400) );
  INV_X1 U5231 ( .A(n4688), .ZN(n4402) );
  NAND2_X1 U5232 ( .A1(n9807), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n4691) );
  OR2_X1 U5233 ( .A1(n5951), .A2(n4275), .ZN(n5589) );
  INV_X1 U5234 ( .A(n8265), .ZN(n8269) );
  NOR2_X1 U5235 ( .A1(n8325), .A2(n4442), .ZN(n4441) );
  AOI21_X1 U5236 ( .B1(n4435), .B2(n4438), .A(n8423), .ZN(n4434) );
  NOR2_X1 U5237 ( .A1(n4439), .A2(n8321), .ZN(n4438) );
  AOI21_X1 U5238 ( .B1(n4434), .B2(n4429), .A(n8338), .ZN(n4430) );
  NOR2_X1 U5239 ( .A1(n8354), .A2(n8385), .ZN(n4455) );
  OR2_X1 U5240 ( .A1(n8244), .A2(n8594), .ZN(n8358) );
  NAND2_X1 U5241 ( .A1(n8358), .A2(n8385), .ZN(n4451) );
  INV_X1 U5242 ( .A(n4815), .ZN(n4813) );
  INV_X1 U5243 ( .A(SI_15_), .ZN(n8815) );
  INV_X1 U5244 ( .A(n4727), .ZN(n4725) );
  INV_X1 U5245 ( .A(n5871), .ZN(n4733) );
  NAND2_X1 U5246 ( .A1(n6714), .A2(n6715), .ZN(n4377) );
  NAND2_X1 U5247 ( .A1(n9414), .A2(n4563), .ZN(n4562) );
  INV_X1 U5248 ( .A(n5518), .ZN(n4629) );
  NAND2_X1 U5249 ( .A1(n5265), .A2(n5244), .ZN(n4489) );
  AND2_X1 U5250 ( .A1(n4491), .A2(n4485), .ZN(n4484) );
  INV_X1 U5251 ( .A(n4489), .ZN(n4485) );
  INV_X1 U5252 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5223) );
  INV_X1 U5253 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n5199) );
  NAND2_X1 U5254 ( .A1(n5157), .A2(n5156), .ZN(n5176) );
  INV_X1 U5255 ( .A(n4839), .ZN(n4504) );
  NOR2_X1 U5256 ( .A1(n5123), .A2(n4507), .ZN(n4506) );
  INV_X1 U5257 ( .A(n5103), .ZN(n4507) );
  NAND2_X1 U5258 ( .A1(n5126), .A2(n5125), .ZN(n5154) );
  OR2_X1 U5259 ( .A1(n5032), .A2(n5031), .ZN(n5033) );
  INV_X1 U5260 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4622) );
  OR2_X1 U5261 ( .A1(n6875), .A2(n5511), .ZN(n5536) );
  INV_X1 U5262 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n4974) );
  OR2_X1 U5263 ( .A1(n8725), .A2(n8096), .ZN(n8380) );
  NAND2_X1 U5264 ( .A1(n6329), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5423) );
  NAND2_X1 U5265 ( .A1(n6329), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5465) );
  INV_X1 U5266 ( .A(n4607), .ZN(n4605) );
  NAND2_X1 U5267 ( .A1(n4418), .A2(n8629), .ZN(n4417) );
  AND2_X1 U5268 ( .A1(n8646), .A2(n8352), .ZN(n4607) );
  INV_X1 U5269 ( .A(n8660), .ZN(n4774) );
  NAND2_X1 U5270 ( .A1(n4580), .A2(n4583), .ZN(n4579) );
  NAND2_X1 U5271 ( .A1(n8300), .A2(n4571), .ZN(n4570) );
  NOR2_X1 U5272 ( .A1(n8411), .A2(n4575), .ZN(n4571) );
  INV_X1 U5273 ( .A(n8413), .ZN(n7070) );
  NOR2_X1 U5274 ( .A1(n4423), .A2(n9853), .ZN(n4422) );
  INV_X1 U5275 ( .A(n4424), .ZN(n4423) );
  AND2_X1 U5276 ( .A1(n4425), .A2(n9926), .ZN(n4424) );
  AND2_X1 U5277 ( .A1(n8249), .A2(n6747), .ZN(n8251) );
  NAND2_X1 U5278 ( .A1(n4449), .A2(n4448), .ZN(n8248) );
  NOR2_X1 U5279 ( .A1(n8595), .A2(n8742), .ZN(n8582) );
  INV_X1 U5280 ( .A(SI_21_), .ZN(n8906) );
  NAND2_X1 U5281 ( .A1(n4780), .A2(n5178), .ZN(n4867) );
  NAND2_X1 U5282 ( .A1(n4864), .A2(n4784), .ZN(n4783) );
  INV_X1 U5283 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4864) );
  INV_X1 U5284 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4784) );
  INV_X1 U5285 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5486) );
  NAND2_X1 U5286 ( .A1(n4621), .A2(n4620), .ZN(n4851) );
  NOR2_X1 U5287 ( .A1(n4848), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n4620) );
  INV_X1 U5288 ( .A(n4849), .ZN(n4621) );
  AND2_X1 U5289 ( .A1(n4855), .A2(n4523), .ZN(n4522) );
  INV_X1 U5290 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n4523) );
  OR2_X1 U5291 ( .A1(n5063), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5129) );
  INV_X1 U5292 ( .A(n9055), .ZN(n4712) );
  INV_X1 U5293 ( .A(n4732), .ZN(n4731) );
  AOI21_X1 U5294 ( .B1(n4732), .B2(n9458), .A(n4310), .ZN(n4730) );
  NOR2_X1 U5295 ( .A1(n4291), .A2(n4733), .ZN(n4732) );
  INV_X1 U5296 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5755) );
  INV_X1 U5297 ( .A(n8047), .ZN(n5603) );
  NAND2_X1 U5298 ( .A1(n4554), .A2(n4553), .ZN(n4552) );
  INV_X1 U5299 ( .A(n4556), .ZN(n4554) );
  NAND2_X1 U5300 ( .A1(n9174), .A2(n4557), .ZN(n4556) );
  INV_X1 U5301 ( .A(n4386), .ZN(n4382) );
  NAND2_X1 U5302 ( .A1(n9233), .A2(n4566), .ZN(n4565) );
  INV_X1 U5303 ( .A(n4567), .ZN(n4566) );
  NAND2_X1 U5304 ( .A1(n5939), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5954) );
  INV_X1 U5305 ( .A(n7670), .ZN(n4667) );
  NOR2_X1 U5306 ( .A1(n4671), .A2(n7670), .ZN(n4666) );
  OAI21_X1 U5307 ( .B1(n9493), .B2(n4315), .A(n4816), .ZN(n7672) );
  NAND2_X1 U5308 ( .A1(n4817), .A2(n4818), .ZN(n4816) );
  INV_X1 U5309 ( .A(n7843), .ZN(n4818) );
  OAI21_X1 U5310 ( .B1(n7318), .B2(n4662), .A(n7383), .ZN(n4661) );
  INV_X1 U5311 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5790) );
  OR2_X1 U5312 ( .A1(n5791), .A2(n5790), .ZN(n5821) );
  NOR2_X1 U5313 ( .A1(n7197), .A2(n7315), .ZN(n7308) );
  NAND2_X1 U5314 ( .A1(n9676), .A2(n7089), .ZN(n7796) );
  NAND2_X1 U5315 ( .A1(n6134), .A2(n9137), .ZN(n6724) );
  NAND2_X1 U5316 ( .A1(n6938), .A2(n6937), .ZN(n4815) );
  INV_X1 U5317 ( .A(n9698), .ZN(n4814) );
  AND2_X1 U5318 ( .A1(n7706), .A2(n7700), .ZN(n7704) );
  NAND2_X1 U5319 ( .A1(n4812), .A2(n4410), .ZN(n4409) );
  INV_X1 U5320 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4410) );
  AND2_X1 U5321 ( .A1(n5452), .A2(n5437), .ZN(n5450) );
  INV_X1 U5322 ( .A(n5416), .ZN(n4638) );
  AOI21_X1 U5323 ( .B1(n5412), .B2(n4637), .A(n4635), .ZN(n4634) );
  INV_X1 U5324 ( .A(n5431), .ZN(n4635) );
  NAND2_X1 U5325 ( .A1(n5567), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5570) );
  AOI21_X1 U5326 ( .B1(n4271), .B2(P1_IR_REG_31__SCAN_IN), .A(
        P1_IR_REG_20__SCAN_IN), .ZN(n4735) );
  NAND2_X1 U5327 ( .A1(n5570), .A2(n5569), .ZN(n5586) );
  INV_X1 U5328 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5569) );
  NAND2_X1 U5329 ( .A1(n4483), .A2(n4487), .ZN(n5287) );
  INV_X1 U5330 ( .A(n4488), .ZN(n4487) );
  NAND2_X1 U5331 ( .A1(n5177), .A2(n4484), .ZN(n4483) );
  OAI21_X1 U5332 ( .B1(n4646), .B2(n4489), .A(n5268), .ZN(n4488) );
  AOI21_X1 U5333 ( .B1(n4650), .B2(n4648), .A(n4647), .ZN(n4646) );
  INV_X1 U5334 ( .A(n5242), .ZN(n4647) );
  INV_X1 U5335 ( .A(n4652), .ZN(n4648) );
  NOR2_X1 U5336 ( .A1(n4649), .A2(n4492), .ZN(n4491) );
  INV_X1 U5337 ( .A(n5176), .ZN(n4492) );
  INV_X1 U5338 ( .A(n4650), .ZN(n4649) );
  NOR2_X1 U5339 ( .A1(n5221), .A2(n4653), .ZN(n4652) );
  INV_X1 U5340 ( .A(n5198), .ZN(n4653) );
  AOI21_X1 U5341 ( .B1(n4652), .B2(n5194), .A(n4651), .ZN(n4650) );
  INV_X1 U5342 ( .A(n5220), .ZN(n4651) );
  NAND2_X1 U5343 ( .A1(n5331), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5358) );
  INV_X1 U5344 ( .A(n5333), .ZN(n5331) );
  NAND2_X1 U5345 ( .A1(n4468), .A2(n8123), .ZN(n8128) );
  NAND2_X1 U5346 ( .A1(n8125), .A2(n5324), .ZN(n4468) );
  INV_X1 U5347 ( .A(n5253), .ZN(n5251) );
  AND2_X1 U5348 ( .A1(n6858), .A2(n4959), .ZN(n4960) );
  NAND2_X1 U5349 ( .A1(n9855), .A2(n5074), .ZN(n8175) );
  OR2_X1 U5350 ( .A1(n6171), .A2(n6172), .ZN(n8125) );
  NAND2_X1 U5351 ( .A1(n8175), .A2(n4619), .ZN(n9833) );
  INV_X1 U5352 ( .A(n6657), .ZN(n4613) );
  OAI21_X1 U5353 ( .B1(n4960), .B2(n4284), .A(n7991), .ZN(n4515) );
  AND2_X1 U5354 ( .A1(n8392), .A2(n8389), .ZN(n8400) );
  NAND2_X1 U5355 ( .A1(n6329), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5527) );
  AND2_X1 U5356 ( .A1(n5408), .A2(n5407), .ZN(n8057) );
  AND2_X1 U5357 ( .A1(n5365), .A2(n5364), .ZN(n8104) );
  INV_X1 U5358 ( .A(n6328), .ZN(n5530) );
  AND4_X1 U5359 ( .A1(n5049), .A2(n5048), .A3(n5047), .A4(n5046), .ZN(n6954)
         );
  NAND2_X1 U5360 ( .A1(n6240), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4536) );
  AND2_X1 U5361 ( .A1(n4535), .A2(n4534), .ZN(n6250) );
  INV_X1 U5362 ( .A(n6251), .ZN(n4534) );
  OR2_X1 U5363 ( .A1(n5039), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5063) );
  AOI21_X1 U5364 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n6791), .A(n6790), .ZN(
        n6793) );
  AOI211_X1 U5365 ( .C1(n7219), .C2(P2_REG1_REG_14__SCAN_IN), .A(n7215), .B(
        n7217), .ZN(n7415) );
  NOR2_X1 U5366 ( .A1(n4525), .A2(n4345), .ZN(n7508) );
  NOR2_X1 U5367 ( .A1(n8479), .A2(n8478), .ZN(n9874) );
  NAND2_X1 U5368 ( .A1(n8226), .A2(n8225), .ZN(n8515) );
  NAND2_X1 U5369 ( .A1(n8380), .A2(n8381), .ZN(n8527) );
  NAND2_X1 U5370 ( .A1(n5386), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5441) );
  NAND2_X1 U5371 ( .A1(n4550), .A2(n4478), .ZN(n8595) );
  INV_X1 U5372 ( .A(n4550), .ZN(n8616) );
  INV_X1 U5373 ( .A(n8356), .ZN(n8632) );
  OR2_X1 U5374 ( .A1(n8653), .A2(n8343), .ZN(n4608) );
  NAND2_X1 U5375 ( .A1(n4608), .A2(n4607), .ZN(n8645) );
  NOR2_X1 U5376 ( .A1(n8676), .A2(n4416), .ZN(n8640) );
  INV_X1 U5377 ( .A(n4418), .ZN(n4416) );
  NAND2_X1 U5378 ( .A1(n8160), .A2(n8701), .ZN(n4420) );
  NOR3_X1 U5379 ( .A1(n7528), .A2(n4421), .A3(n8787), .ZN(n8694) );
  NOR2_X1 U5380 ( .A1(n7528), .A2(n4421), .ZN(n7643) );
  NAND2_X1 U5381 ( .A1(n7599), .A2(n4778), .ZN(n7638) );
  NAND2_X1 U5382 ( .A1(n7442), .A2(n8319), .ZN(n7528) );
  NAND2_X1 U5383 ( .A1(n7521), .A2(n8422), .ZN(n7599) );
  NAND2_X1 U5384 ( .A1(n5163), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5182) );
  NOR2_X1 U5385 ( .A1(n7438), .A2(n7373), .ZN(n7442) );
  NAND2_X1 U5386 ( .A1(n4549), .A2(n4548), .ZN(n7373) );
  AND4_X1 U5387 ( .A1(n5115), .A2(n5114), .A3(n5113), .A4(n5112), .ZN(n7345)
         );
  AND3_X1 U5388 ( .A1(n7126), .A2(n4422), .A3(n7111), .ZN(n7078) );
  AOI21_X1 U5389 ( .B1(n4746), .B2(n4747), .A(n4307), .ZN(n4744) );
  NAND2_X1 U5390 ( .A1(n7126), .A2(n4424), .ZN(n6783) );
  NAND2_X1 U5391 ( .A1(n7126), .A2(n9926), .ZN(n7125) );
  OR2_X1 U5392 ( .A1(n9936), .A2(n8583), .ZN(n6878) );
  NAND2_X1 U5393 ( .A1(n6585), .A2(n6584), .ZN(n8403) );
  NAND2_X1 U5394 ( .A1(n8260), .A2(n8403), .ZN(n7000) );
  NAND2_X1 U5395 ( .A1(n8064), .A2(n8063), .ZN(n8720) );
  NAND2_X1 U5396 ( .A1(n4775), .A2(n8053), .ZN(n8661) );
  NAND2_X1 U5397 ( .A1(n4775), .A2(n4772), .ZN(n8770) );
  OR2_X1 U5398 ( .A1(n8399), .A2(n5535), .ZN(n9936) );
  AND2_X1 U5399 ( .A1(n8442), .A2(n9899), .ZN(n9475) );
  INV_X1 U5400 ( .A(n9936), .ZN(n9912) );
  INV_X1 U5401 ( .A(n6884), .ZN(n9907) );
  INV_X1 U5402 ( .A(n9475), .ZN(n9934) );
  AND2_X1 U5403 ( .A1(n6181), .A2(n9893), .ZN(n9886) );
  NOR2_X1 U5404 ( .A1(n4781), .A2(n8964), .ZN(n4376) );
  INV_X1 U5405 ( .A(n4867), .ZN(n4542) );
  OR2_X1 U5406 ( .A1(n5494), .A2(n4783), .ZN(n4866) );
  NAND2_X1 U5407 ( .A1(n5178), .A2(n4863), .ZN(n5494) );
  AOI21_X1 U5408 ( .B1(n4849), .B2(P2_IR_REG_31__SCAN_IN), .A(n4494), .ZN(
        n4493) );
  NAND2_X1 U5409 ( .A1(n4495), .A2(n4860), .ZN(n4494) );
  NAND2_X1 U5410 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), 
        .ZN(n4495) );
  NAND2_X1 U5411 ( .A1(n5178), .A2(n4855), .ZN(n5203) );
  NAND2_X1 U5412 ( .A1(n4903), .A2(n4842), .ZN(n4947) );
  AOI21_X1 U5413 ( .B1(n4277), .B2(n4709), .A(n4333), .ZN(n4704) );
  INV_X1 U5414 ( .A(n9191), .ZN(n9009) );
  NOR2_X1 U5415 ( .A1(n5756), .A2(n5755), .ZN(n5774) );
  NAND2_X1 U5416 ( .A1(n7683), .A2(n7684), .ZN(n4727) );
  OR2_X1 U5417 ( .A1(n7683), .A2(n7684), .ZN(n4728) );
  INV_X1 U5418 ( .A(n6682), .ZN(n5711) );
  AND2_X1 U5419 ( .A1(n6005), .A2(n5599), .ZN(n6020) );
  CLKBUF_X1 U5420 ( .A(n9062), .Z(n4354) );
  NAND2_X1 U5421 ( .A1(n4354), .A2(n9063), .ZN(n9061) );
  NAND2_X1 U5422 ( .A1(n5868), .A2(n5867), .ZN(n9462) );
  INV_X1 U5423 ( .A(n6040), .ZN(n4715) );
  OR2_X1 U5424 ( .A1(n5821), .A2(n6445), .ZN(n5840) );
  INV_X1 U5425 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5839) );
  INV_X1 U5426 ( .A(n9125), .ZN(n6928) );
  AND3_X1 U5427 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5735) );
  OR2_X1 U5428 ( .A1(n4710), .A2(n4708), .ZN(n4707) );
  INV_X1 U5429 ( .A(n4713), .ZN(n4708) );
  AND2_X1 U5430 ( .A1(n9038), .A2(n4711), .ZN(n4710) );
  NAND2_X1 U5431 ( .A1(n4712), .A2(n4714), .ZN(n4711) );
  NAND2_X1 U5432 ( .A1(n4713), .A2(n4714), .ZN(n4709) );
  INV_X1 U5433 ( .A(n4369), .ZN(n4368) );
  OAI21_X1 U5434 ( .B1(n7898), .B2(n7897), .A(n4370), .ZN(n4369) );
  NAND2_X1 U5435 ( .A1(n4644), .A2(n9721), .ZN(n4643) );
  INV_X1 U5436 ( .A(n7935), .ZN(n4644) );
  NAND2_X1 U5437 ( .A1(n7934), .A2(n9137), .ZN(n4642) );
  INV_X1 U5438 ( .A(n5675), .ZN(n6049) );
  INV_X2 U5439 ( .A(n5991), .ZN(n7723) );
  INV_X1 U5440 ( .A(n5676), .ZN(n5991) );
  NAND2_X1 U5441 ( .A1(n6153), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5677) );
  NOR2_X1 U5442 ( .A1(n6462), .A2(n6461), .ZN(n6460) );
  CLKBUF_X1 U5443 ( .A(n5741), .Z(n5743) );
  AOI21_X1 U5444 ( .B1(n6366), .B2(n9818), .A(n6378), .ZN(n6367) );
  AOI21_X1 U5445 ( .B1(n9528), .B2(n7448), .A(n7447), .ZN(n9620) );
  AOI21_X1 U5446 ( .B1(n7450), .B2(n7449), .A(n9618), .ZN(n7451) );
  NOR3_X1 U5447 ( .A1(n9197), .A2(n9337), .A3(n4552), .ZN(n9148) );
  NOR2_X1 U5448 ( .A1(n9197), .A2(n4552), .ZN(n9157) );
  NOR2_X1 U5449 ( .A1(n9197), .A2(n9355), .ZN(n9186) );
  NAND2_X1 U5450 ( .A1(n4693), .A2(n4692), .ZN(n9196) );
  OR2_X1 U5451 ( .A1(n9366), .A2(n9206), .ZN(n4692) );
  NAND2_X1 U5452 ( .A1(n9212), .A2(n4298), .ZN(n4693) );
  NOR3_X1 U5453 ( .A1(n9269), .A2(n9366), .A3(n4565), .ZN(n9213) );
  NAND2_X1 U5454 ( .A1(n4380), .A2(n4379), .ZN(n9212) );
  OR2_X1 U5455 ( .A1(n4381), .A2(n4694), .ZN(n4379) );
  NAND2_X1 U5456 ( .A1(n8006), .A2(n4303), .ZN(n4380) );
  NOR2_X1 U5457 ( .A1(n4296), .A2(n4382), .ZN(n4381) );
  NOR2_X1 U5458 ( .A1(n9269), .A2(n4565), .ZN(n9229) );
  AND2_X1 U5459 ( .A1(n6020), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6032) );
  NOR2_X1 U5460 ( .A1(n9269), .A2(n4567), .ZN(n9242) );
  NAND2_X1 U5461 ( .A1(n4799), .A2(n4797), .ZN(n9256) );
  AOI21_X1 U5462 ( .B1(n4800), .B2(n4803), .A(n4798), .ZN(n4797) );
  AOI21_X1 U5463 ( .B1(n4802), .B2(n4801), .A(n8017), .ZN(n4800) );
  NOR2_X1 U5464 ( .A1(n5974), .A2(n5973), .ZN(n6005) );
  AND2_X1 U5465 ( .A1(n9321), .A2(n9305), .ZN(n9303) );
  AND2_X1 U5466 ( .A1(n9296), .A2(n8012), .ZN(n9316) );
  NAND2_X1 U5467 ( .A1(n4388), .A2(n4664), .ZN(n7999) );
  AOI21_X1 U5468 ( .B1(n4666), .B2(n4668), .A(n4665), .ZN(n4664) );
  NAND2_X1 U5469 ( .A1(n9490), .A2(n4300), .ZN(n4388) );
  NOR2_X1 U5470 ( .A1(n9414), .A2(n7690), .ZN(n4665) );
  NOR2_X1 U5471 ( .A1(n5898), .A2(n7625), .ZN(n5912) );
  NAND2_X1 U5472 ( .A1(n4819), .A2(n7567), .ZN(n9491) );
  INV_X1 U5473 ( .A(n9493), .ZN(n4819) );
  NAND2_X1 U5474 ( .A1(n5855), .A2(n5854), .ZN(n7560) );
  AOI21_X1 U5475 ( .B1(n7757), .B2(n7813), .A(n4822), .ZN(n4821) );
  INV_X1 U5476 ( .A(n7746), .ZN(n4822) );
  NAND2_X1 U5477 ( .A1(n7381), .A2(n7380), .ZN(n9505) );
  AND2_X1 U5478 ( .A1(n7308), .A2(n7312), .ZN(n9507) );
  NAND2_X1 U5479 ( .A1(n7314), .A2(n7313), .ZN(n7319) );
  NAND2_X1 U5480 ( .A1(n7319), .A2(n7318), .ZN(n7381) );
  OR2_X1 U5481 ( .A1(n7188), .A2(n7813), .ZN(n7386) );
  AND2_X1 U5482 ( .A1(n7821), .A2(n7808), .ZN(n7915) );
  NAND2_X1 U5483 ( .A1(n4560), .A2(n7094), .ZN(n7197) );
  INV_X1 U5484 ( .A(n7172), .ZN(n4560) );
  NAND2_X1 U5485 ( .A1(n7097), .A2(n7096), .ZN(n7196) );
  AND2_X1 U5486 ( .A1(n7803), .A2(n7804), .ZN(n7911) );
  NAND2_X1 U5487 ( .A1(n7174), .A2(n7173), .ZN(n7172) );
  AND2_X1 U5488 ( .A1(n7795), .A2(n7796), .ZN(n7909) );
  NOR2_X1 U5489 ( .A1(n9684), .A2(n7053), .ZN(n7174) );
  INV_X1 U5490 ( .A(n7089), .ZN(n7053) );
  NAND2_X1 U5491 ( .A1(n7057), .A2(n7736), .ZN(n9673) );
  AND2_X1 U5492 ( .A1(n7741), .A2(n7743), .ZN(n9680) );
  NAND2_X1 U5493 ( .A1(n4411), .A2(n6167), .ZN(n4414) );
  NAND2_X1 U5494 ( .A1(n5635), .A2(n5634), .ZN(n5636) );
  NAND2_X1 U5495 ( .A1(n4413), .A2(n4412), .ZN(n4411) );
  NAND2_X1 U5496 ( .A1(n6714), .A2(n4558), .ZN(n9716) );
  NOR2_X1 U5497 ( .A1(n9425), .A2(n4405), .ZN(n4404) );
  INV_X1 U5498 ( .A(n4689), .ZN(n4405) );
  NOR2_X1 U5499 ( .A1(n8030), .A2(n4331), .ZN(n4688) );
  NAND2_X1 U5500 ( .A1(n5988), .A2(n5987), .ZN(n9391) );
  OR2_X1 U5501 ( .A1(n6736), .A2(n7977), .ZN(n9799) );
  NAND2_X1 U5502 ( .A1(n8043), .A2(n8041), .ZN(n6736) );
  INV_X1 U5503 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4811) );
  XNOR2_X1 U5504 ( .A(n7720), .B(SI_30_), .ZN(n8224) );
  XNOR2_X1 U5505 ( .A(n7705), .B(n7704), .ZN(n8062) );
  AND2_X1 U5506 ( .A1(n7696), .A2(n5523), .ZN(n7694) );
  AND2_X1 U5507 ( .A1(n5518), .A2(n5456), .ZN(n5516) );
  CLKBUF_X1 U5508 ( .A(n6140), .Z(n6141) );
  XNOR2_X1 U5509 ( .A(n5433), .B(n5432), .ZN(n7535) );
  NAND2_X1 U5510 ( .A1(n4639), .A2(n5416), .ZN(n5433) );
  OR2_X1 U5511 ( .A1(n5413), .A2(n5412), .ZN(n4639) );
  XNOR2_X1 U5512 ( .A(n5588), .B(n5587), .ZN(n6132) );
  INV_X1 U5513 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U5514 ( .A1(n5586), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U5515 ( .A1(n4264), .A2(n4837), .ZN(n5835) );
  NAND2_X1 U5516 ( .A1(n4508), .A2(n5103), .ZN(n5124) );
  NAND2_X1 U5517 ( .A1(n5102), .A2(n4839), .ZN(n4508) );
  NAND2_X1 U5518 ( .A1(n5011), .A2(n5024), .ZN(n4363) );
  NAND2_X1 U5519 ( .A1(n5027), .A2(n5025), .ZN(n5008) );
  NAND2_X1 U5520 ( .A1(n4496), .A2(n4497), .ZN(n4986) );
  AOI21_X1 U5521 ( .B1(n4963), .B2(n4498), .A(n4312), .ZN(n4497) );
  AND3_X1 U5522 ( .A1(n5660), .A2(n5544), .A3(n5545), .ZN(n5723) );
  AND2_X1 U5523 ( .A1(n5660), .A2(n5544), .ZN(n5700) );
  XNOR2_X1 U5524 ( .A(n4898), .B(n4873), .ZN(n4897) );
  AOI21_X1 U5525 ( .B1(n8103), .B2(n4469), .A(n4334), .ZN(n4471) );
  NOR2_X1 U5526 ( .A1(n4283), .A2(n4470), .ZN(n4469) );
  NAND2_X1 U5527 ( .A1(n5458), .A2(n5457), .ZN(n8732) );
  NAND2_X1 U5528 ( .A1(n8175), .A2(n5078), .ZN(n9836) );
  AND4_X1 U5529 ( .A1(n5072), .A2(n5071), .A3(n5070), .A4(n5069), .ZN(n9832)
         );
  AND2_X1 U5530 ( .A1(n6838), .A2(n4918), .ZN(n6656) );
  NAND2_X1 U5531 ( .A1(n6656), .A2(n6657), .ZN(n6850) );
  NAND2_X1 U5532 ( .A1(n5296), .A2(n5295), .ZN(n8778) );
  INV_X1 U5533 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8840) );
  AND4_X1 U5534 ( .A1(n5279), .A2(n5278), .A3(n5277), .A4(n5276), .ZN(n8155)
         );
  NAND2_X1 U5535 ( .A1(n7491), .A2(n4618), .ZN(n8201) );
  NAND2_X1 U5536 ( .A1(n7491), .A2(n5241), .ZN(n8152) );
  NAND2_X1 U5537 ( .A1(n9845), .A2(n8239), .ZN(n8202) );
  OR2_X1 U5538 ( .A1(n8209), .A2(n8562), .ZN(n9831) );
  NAND2_X1 U5539 ( .A1(n7352), .A2(n4301), .ZN(n9471) );
  NAND2_X1 U5540 ( .A1(n7352), .A2(n5151), .ZN(n7326) );
  NAND2_X1 U5541 ( .A1(n5355), .A2(n5354), .ZN(n8759) );
  NAND2_X1 U5542 ( .A1(n4518), .A2(n4521), .ZN(n4516) );
  INV_X1 U5543 ( .A(n4619), .ZN(n4521) );
  NAND2_X1 U5544 ( .A1(n4616), .A2(n4893), .ZN(n6846) );
  INV_X1 U5545 ( .A(n6618), .ZN(n4616) );
  AOI21_X1 U5546 ( .B1(n4618), .B2(n4512), .A(n4511), .ZN(n4510) );
  NAND2_X1 U5547 ( .A1(n4611), .A2(n4514), .ZN(n7997) );
  NAND2_X1 U5548 ( .A1(n6656), .A2(n4612), .ZN(n4611) );
  INV_X1 U5549 ( .A(n4515), .ZN(n4514) );
  NOR2_X1 U5550 ( .A1(n4613), .A2(n4284), .ZN(n4612) );
  NAND2_X1 U5551 ( .A1(n4473), .A2(n8139), .ZN(n8216) );
  NAND2_X1 U5552 ( .A1(n4474), .A2(n4476), .ZN(n4473) );
  NOR2_X1 U5553 ( .A1(n4446), .A2(n4445), .ZN(n4444) );
  AND2_X1 U5554 ( .A1(n8437), .A2(n8436), .ZN(n4445) );
  NAND2_X1 U5555 ( .A1(n7088), .A2(n8583), .ZN(n8442) );
  INV_X1 U5556 ( .A(n8104), .ZN(n8648) );
  NAND2_X1 U5557 ( .A1(n6329), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n4980) );
  NAND2_X1 U5558 ( .A1(n4972), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n4911) );
  NAND2_X1 U5559 ( .A1(n4972), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n4883) );
  INV_X2 U5560 ( .A(P2_U3966), .ZN(n8466) );
  AOI21_X1 U5561 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n6253), .A(n6254), .ZN(
        n6231) );
  AOI21_X1 U5562 ( .B1(n6266), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6267), .ZN(
        n6281) );
  INV_X1 U5563 ( .A(n4530), .ZN(n6276) );
  INV_X1 U5564 ( .A(n4528), .ZN(n6630) );
  AND2_X1 U5565 ( .A1(n4528), .A2(n4527), .ZN(n6633) );
  NAND2_X1 U5566 ( .A1(n6631), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4527) );
  NOR2_X1 U5567 ( .A1(n6662), .A2(n6663), .ZN(n6693) );
  NOR2_X1 U5568 ( .A1(n6660), .A2(n4539), .ZN(n6663) );
  AND2_X1 U5569 ( .A1(n6666), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4539) );
  AOI21_X1 U5570 ( .B1(n6666), .B2(P2_REG1_REG_9__SCAN_IN), .A(n6665), .ZN(
        n6669) );
  NOR2_X1 U5571 ( .A1(n6693), .A2(n4538), .ZN(n6695) );
  AND2_X1 U5572 ( .A1(n6694), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4538) );
  OAI21_X1 U5573 ( .B1(n6970), .B2(n6969), .A(n4526), .ZN(n7206) );
  OR2_X1 U5574 ( .A1(n6968), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4526) );
  INV_X1 U5575 ( .A(n4525), .ZN(n7411) );
  NOR2_X1 U5576 ( .A1(n8474), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8493) );
  INV_X1 U5577 ( .A(n8515), .ZN(n8719) );
  INV_X1 U5578 ( .A(n8085), .ZN(n8086) );
  AOI22_X1 U5579 ( .A1(n8549), .A2(n8656), .B1(n8509), .B2(n8449), .ZN(n8085)
         );
  NAND2_X1 U5580 ( .A1(n5439), .A2(n5438), .ZN(n8737) );
  NAND2_X1 U5581 ( .A1(n4588), .A2(n4589), .ZN(n8559) );
  NAND2_X1 U5582 ( .A1(n8593), .A2(n8058), .ZN(n8576) );
  INV_X1 U5583 ( .A(n4594), .ZN(n8588) );
  NAND2_X1 U5584 ( .A1(n5379), .A2(n5378), .ZN(n8618) );
  CLKBUF_X1 U5585 ( .A(n8603), .Z(n8605) );
  NAND2_X1 U5586 ( .A1(n5315), .A2(n5314), .ZN(n8771) );
  OAI21_X1 U5587 ( .B1(n7635), .B2(n4583), .A(n4580), .ZN(n8685) );
  NAND2_X1 U5588 ( .A1(n8071), .A2(n8331), .ZN(n8705) );
  NAND2_X1 U5589 ( .A1(n5231), .A2(n5230), .ZN(n8795) );
  NAND2_X1 U5590 ( .A1(n4597), .A2(n7523), .ZN(n7526) );
  NAND2_X1 U5591 ( .A1(n7433), .A2(n8315), .ZN(n7524) );
  NAND2_X1 U5592 ( .A1(n5181), .A2(n5180), .ZN(n9476) );
  NAND2_X1 U5593 ( .A1(n4748), .A2(n4750), .ZN(n7363) );
  NAND2_X1 U5594 ( .A1(n4754), .A2(n7238), .ZN(n7362) );
  NAND2_X1 U5595 ( .A1(n4371), .A2(n8414), .ZN(n4754) );
  NAND2_X1 U5596 ( .A1(n4574), .A2(n4573), .ZN(n7248) );
  NAND2_X1 U5597 ( .A1(n4762), .A2(n7069), .ZN(n7071) );
  NAND2_X1 U5598 ( .A1(n4577), .A2(n8285), .ZN(n6750) );
  NAND2_X1 U5599 ( .A1(n7123), .A2(n6744), .ZN(n6745) );
  OAI21_X1 U5600 ( .B1(n7124), .B2(n4747), .A(n4746), .ZN(n6773) );
  AND3_X1 U5601 ( .A1(n4971), .A2(n4970), .A3(n4969), .ZN(n6995) );
  NAND2_X1 U5602 ( .A1(n8688), .A2(n6887), .ZN(n8700) );
  NAND2_X1 U5603 ( .A1(n8688), .A2(n6888), .ZN(n8711) );
  INV_X1 U5604 ( .A(n8700), .ZN(n8666) );
  AND2_X1 U5605 ( .A1(n8723), .A2(n8722), .ZN(n4373) );
  INV_X1 U5606 ( .A(n4428), .ZN(n4427) );
  OAI21_X1 U5607 ( .B1(n8723), .B2(n9942), .A(n4769), .ZN(n4428) );
  NAND2_X1 U5608 ( .A1(n9942), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n4769) );
  AOI21_X1 U5609 ( .B1(n8721), .B2(n9912), .A(n4547), .ZN(n8722) );
  AND2_X1 U5610 ( .A1(n8720), .A2(n9475), .ZN(n4547) );
  AND2_X1 U5611 ( .A1(n6180), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9893) );
  AND2_X1 U5612 ( .A1(n5178), .A2(n4461), .ZN(n4459) );
  AND2_X1 U5613 ( .A1(n4877), .A2(n4462), .ZN(n4461) );
  INV_X1 U5614 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8907) );
  NAND2_X1 U5615 ( .A1(n5489), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5491) );
  INV_X1 U5616 ( .A(n8255), .ZN(n8436) );
  INV_X1 U5617 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7087) );
  XNOR2_X1 U5618 ( .A(n4845), .B(n4847), .ZN(n7088) );
  NAND2_X1 U5619 ( .A1(n4854), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4845) );
  INV_X1 U5620 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6808) );
  NAND2_X1 U5621 ( .A1(n4849), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5270) );
  INV_X1 U5622 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n8831) );
  INV_X1 U5623 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n8891) );
  INV_X1 U5624 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6421) );
  INV_X1 U5625 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6338) );
  INV_X1 U5626 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6319) );
  INV_X1 U5627 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6307) );
  INV_X1 U5628 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6305) );
  INV_X1 U5629 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n8933) );
  AND2_X1 U5630 ( .A1(n4701), .A2(n4698), .ZN(n7138) );
  INV_X1 U5631 ( .A(n5816), .ZN(n4698) );
  NAND2_X1 U5632 ( .A1(n4702), .A2(n4274), .ZN(n4701) );
  INV_X1 U5633 ( .A(n7146), .ZN(n4702) );
  NAND2_X1 U5634 ( .A1(n5820), .A2(n5819), .ZN(n7402) );
  AND2_X1 U5635 ( .A1(n9015), .A2(n9086), .ZN(n9005) );
  AND2_X1 U5636 ( .A1(n6109), .A2(n6108), .ZN(n9014) );
  AND2_X1 U5637 ( .A1(n9061), .A2(n9065), .ZN(n9031) );
  NAND2_X1 U5639 ( .A1(n4726), .A2(n4727), .ZN(n9045) );
  NAND2_X1 U5640 ( .A1(n4355), .A2(n4728), .ZN(n4726) );
  INV_X1 U5641 ( .A(n9222), .ZN(n9251) );
  INV_X1 U5642 ( .A(n6934), .ZN(n9764) );
  NAND2_X1 U5643 ( .A1(n6004), .A2(n6003), .ZN(n9385) );
  INV_X1 U5644 ( .A(n9119), .ZN(n9512) );
  AND2_X1 U5645 ( .A1(n9462), .A2(n5871), .ZN(n7425) );
  OAI22_X1 U5646 ( .A1(n6863), .A2(n4279), .B1(n4697), .B2(n4699), .ZN(n7230)
         );
  INV_X1 U5647 ( .A(n4346), .ZN(n4697) );
  INV_X1 U5648 ( .A(n9468), .ZN(n9099) );
  INV_X1 U5649 ( .A(n9221), .ZN(n9105) );
  NAND2_X1 U5650 ( .A1(n4706), .A2(n4707), .ZN(n9098) );
  OR2_X1 U5651 ( .A1(n9054), .A2(n4709), .ZN(n4706) );
  INV_X1 U5652 ( .A(n7986), .ZN(n4351) );
  NOR2_X1 U5653 ( .A1(n6442), .A2(n9604), .ZN(n6444) );
  AOI21_X1 U5654 ( .B1(n6493), .B2(n6517), .A(n6513), .ZN(n6515) );
  AND2_X1 U5655 ( .A1(n9551), .A2(n6355), .ZN(n9663) );
  INV_X1 U5656 ( .A(n9334), .ZN(n9149) );
  OAI21_X1 U5657 ( .B1(n9189), .B2(n4824), .A(n4825), .ZN(n8031) );
  AOI21_X1 U5658 ( .B1(n4272), .B2(n4827), .A(n4826), .ZN(n4825) );
  NAND2_X1 U5659 ( .A1(n4830), .A2(n4272), .ZN(n9161) );
  NAND2_X1 U5660 ( .A1(n4831), .A2(n8026), .ZN(n9176) );
  NAND2_X1 U5661 ( .A1(n4786), .A2(n4789), .ZN(n9220) );
  NAND2_X1 U5662 ( .A1(n4796), .A2(n4791), .ZN(n4786) );
  NAND2_X1 U5663 ( .A1(n4795), .A2(n8021), .ZN(n9234) );
  NAND2_X1 U5664 ( .A1(n4383), .A2(n4386), .ZN(n9228) );
  NAND2_X1 U5665 ( .A1(n8006), .A2(n4285), .ZN(n4383) );
  NAND2_X1 U5666 ( .A1(n6019), .A2(n6018), .ZN(n9382) );
  NAND2_X1 U5667 ( .A1(n4390), .A2(n4392), .ZN(n9268) );
  OR2_X1 U5668 ( .A1(n9311), .A2(n4394), .ZN(n4390) );
  AOI21_X1 U5669 ( .B1(n9297), .B2(n8014), .A(n4809), .ZN(n9284) );
  NAND2_X1 U5670 ( .A1(n4804), .A2(n4805), .ZN(n9282) );
  AND2_X1 U5671 ( .A1(n4684), .A2(n4683), .ZN(n9281) );
  NAND2_X1 U5672 ( .A1(n5953), .A2(n5952), .ZN(n9405) );
  NAND2_X1 U5673 ( .A1(n5938), .A2(n5937), .ZN(n9410) );
  NAND2_X1 U5674 ( .A1(n5911), .A2(n5910), .ZN(n7669) );
  OAI21_X1 U5675 ( .B1(n9490), .B2(n4670), .A(n4668), .ZN(n7671) );
  NAND2_X1 U5676 ( .A1(n4673), .A2(n4674), .ZN(n7575) );
  NAND2_X1 U5677 ( .A1(n9490), .A2(n4675), .ZN(n4673) );
  NAND2_X1 U5678 ( .A1(n5876), .A2(n5875), .ZN(n9499) );
  OR3_X1 U5679 ( .A1(n6736), .A2(n6722), .A3(n7980), .ZN(n9709) );
  NAND2_X1 U5680 ( .A1(n7092), .A2(n7091), .ZN(n7171) );
  INV_X1 U5681 ( .A(n9556), .ZN(n5620) );
  AND2_X1 U5682 ( .A1(n9260), .A2(n9717), .ZN(n9696) );
  INV_X1 U5683 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5594) );
  XNOR2_X1 U5684 ( .A(n7718), .B(n7717), .ZN(n9448) );
  XNOR2_X1 U5685 ( .A(n7695), .B(n7694), .ZN(n7772) );
  NAND2_X1 U5686 ( .A1(n4626), .A2(n5518), .ZN(n7695) );
  NAND2_X1 U5687 ( .A1(n5517), .A2(n5516), .ZN(n4626) );
  XNOR2_X1 U5688 ( .A(n5576), .B(n5575), .ZN(n7559) );
  XNOR2_X1 U5689 ( .A(n5381), .B(n5380), .ZN(n7261) );
  INV_X1 U5690 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8948) );
  INV_X1 U5691 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7703) );
  INV_X1 U5692 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6810) );
  INV_X1 U5693 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6569) );
  INV_X1 U5694 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6510) );
  INV_X1 U5695 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n8934) );
  INV_X1 U5696 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6339) );
  INV_X1 U5697 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n8890) );
  INV_X1 U5698 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6321) );
  INV_X1 U5699 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6309) );
  XNOR2_X1 U5700 ( .A(n5008), .B(n5031), .ZN(n6308) );
  INV_X1 U5701 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6302) );
  INV_X1 U5702 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6298) );
  XNOR2_X1 U5703 ( .A(n4964), .B(n4963), .ZN(n6300) );
  NAND2_X1 U5704 ( .A1(n4499), .A2(n4945), .ZN(n4964) );
  INV_X1 U5705 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6297) );
  XNOR2_X1 U5706 ( .A(n5683), .B(n5682), .ZN(n6412) );
  NOR2_X1 U5707 ( .A1(n7298), .A2(n9994), .ZN(n9982) );
  AOI21_X1 U5708 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9980), .ZN(n9979) );
  NOR2_X1 U5709 ( .A1(n9979), .A2(n9978), .ZN(n9977) );
  NAND2_X1 U5710 ( .A1(n6837), .A2(n4999), .ZN(n6763) );
  AND2_X1 U5711 ( .A1(n8725), .A2(n9845), .ZN(n4482) );
  AOI21_X1 U5712 ( .B1(n4533), .B2(n8569), .A(n4532), .ZN(n4531) );
  OAI21_X1 U5713 ( .B1(n8724), .B2(n4768), .A(n4763), .ZN(P2_U3517) );
  NAND2_X1 U5714 ( .A1(n9944), .A2(n9931), .ZN(n4768) );
  INV_X1 U5715 ( .A(n4764), .ZN(n4763) );
  OAI21_X1 U5716 ( .B1(n8722), .B2(n9942), .A(n4427), .ZN(n4764) );
  OAI21_X1 U5717 ( .B1(n9174), .B2(n9095), .A(n6160), .ZN(n6161) );
  XNOR2_X1 U5718 ( .A(n4365), .B(n4364), .ZN(n9044) );
  NAND2_X1 U5719 ( .A1(n4358), .A2(n4356), .ZN(P1_U3260) );
  NAND2_X1 U5720 ( .A1(n9139), .A2(n9721), .ZN(n4358) );
  AOI21_X1 U5721 ( .B1(n9138), .B2(n9137), .A(n4357), .ZN(n4356) );
  NAND2_X1 U5722 ( .A1(n9823), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n4406) );
  NAND2_X1 U5723 ( .A1(n4401), .A2(n9826), .ZN(n4399) );
  NAND2_X1 U5724 ( .A1(n9809), .A2(n9805), .ZN(n4687) );
  INV_X1 U5725 ( .A(n4686), .ZN(n4685) );
  OAI21_X1 U5726 ( .B1(n9343), .B2(n9807), .A(n4691), .ZN(n4686) );
  OR2_X1 U5727 ( .A1(n4275), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n4271) );
  AND2_X1 U5728 ( .A1(n9162), .A2(n8028), .ZN(n4272) );
  INV_X1 U5729 ( .A(n8462), .ZN(n4448) );
  INV_X1 U5730 ( .A(n9219), .ZN(n4788) );
  AND2_X1 U5731 ( .A1(n4745), .A2(n4744), .ZN(n4273) );
  NOR2_X1 U5732 ( .A1(n7145), .A2(n5815), .ZN(n4274) );
  OR2_X1 U5733 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n4275) );
  AND2_X1 U5734 ( .A1(n7796), .A2(n7743), .ZN(n4276) );
  AND2_X1 U5735 ( .A1(n4707), .A2(n4705), .ZN(n4277) );
  AND2_X1 U5736 ( .A1(n7902), .A2(n8021), .ZN(n4278) );
  INV_X1 U5737 ( .A(n8016), .ZN(n4798) );
  XNOR2_X1 U5738 ( .A(n8742), .B(n8561), .ZN(n8575) );
  INV_X1 U5739 ( .A(n8575), .ZN(n4359) );
  OAI21_X1 U5740 ( .B1(n4440), .B2(n4432), .A(n4436), .ZN(n4429) );
  AND2_X1 U5741 ( .A1(n5392), .A2(n5391), .ZN(n8165) );
  INV_X1 U5742 ( .A(n8165), .ZN(n4477) );
  NAND2_X1 U5743 ( .A1(n4274), .A2(n4346), .ZN(n4279) );
  AND2_X1 U5744 ( .A1(n4750), .A2(n4755), .ZN(n4280) );
  OAI21_X2 U5745 ( .B1(n6167), .B2(n5620), .A(n5619), .ZN(n6800) );
  INV_X1 U5746 ( .A(n6800), .ZN(n4558) );
  OR3_X1 U5747 ( .A1(n7569), .A2(n4562), .A3(n9421), .ZN(n4281) );
  INV_X1 U5748 ( .A(n9421), .ZN(n4677) );
  INV_X1 U5749 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4846) );
  INV_X1 U5750 ( .A(n9366), .ZN(n9217) );
  NAND2_X1 U5751 ( .A1(n5563), .A2(n5562), .ZN(n9366) );
  NAND2_X1 U5752 ( .A1(n8103), .A2(n5409), .ZN(n4476) );
  OR2_X1 U5753 ( .A1(n6167), .A2(n9576), .ZN(n4282) );
  INV_X1 U5754 ( .A(n6926), .ZN(n6927) );
  NAND2_X1 U5755 ( .A1(n5250), .A2(n5249), .ZN(n8787) );
  NAND2_X1 U5756 ( .A1(n8139), .A2(n4472), .ZN(n4283) );
  AND2_X1 U5757 ( .A1(n4962), .A2(n4961), .ZN(n4284) );
  NOR2_X1 U5758 ( .A1(n8007), .A2(n4384), .ZN(n4285) );
  AND2_X1 U5759 ( .A1(n4804), .A2(n4802), .ZN(n4286) );
  INV_X1 U5760 ( .A(n8021), .ZN(n4794) );
  OR2_X1 U5761 ( .A1(n8594), .A2(n8589), .ZN(n4287) );
  AND2_X1 U5762 ( .A1(n8006), .A2(n8005), .ZN(n4288) );
  AND2_X1 U5763 ( .A1(n4594), .A2(n8363), .ZN(n4289) );
  AND2_X1 U5764 ( .A1(n4963), .A2(n4941), .ZN(n4290) );
  NAND2_X1 U5765 ( .A1(n5773), .A2(n5772), .ZN(n7194) );
  INV_X1 U5766 ( .A(n8029), .ZN(n4826) );
  AND2_X1 U5767 ( .A1(n7423), .A2(n5888), .ZN(n4291) );
  AND2_X1 U5768 ( .A1(n6212), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4292) );
  AND2_X1 U5769 ( .A1(n7930), .A2(n7897), .ZN(n4293) );
  INV_X1 U5770 ( .A(n8317), .ZN(n4442) );
  NOR2_X1 U5771 ( .A1(n8607), .A2(n4761), .ZN(n4294) );
  AND2_X1 U5772 ( .A1(n8331), .A2(n8329), .ZN(n7640) );
  INV_X1 U5773 ( .A(n7640), .ZN(n4582) );
  AND2_X1 U5774 ( .A1(n8473), .A2(n8480), .ZN(n4295) );
  AND2_X1 U5775 ( .A1(n9233), .A2(n9251), .ZN(n4296) );
  AND2_X1 U5776 ( .A1(n9065), .A2(n4719), .ZN(n4297) );
  NAND2_X1 U5777 ( .A1(n5330), .A2(n5329), .ZN(n8764) );
  OR2_X1 U5778 ( .A1(n9217), .A2(n9236), .ZN(n4298) );
  AND2_X1 U5779 ( .A1(n4795), .A2(n4793), .ZN(n4299) );
  INV_X1 U5780 ( .A(n4803), .ZN(n4802) );
  NAND2_X1 U5781 ( .A1(n4805), .A2(n8015), .ZN(n4803) );
  NAND2_X1 U5782 ( .A1(n7781), .A2(n7780), .ZN(n9337) );
  INV_X1 U5783 ( .A(n7380), .ZN(n4662) );
  AND2_X1 U5784 ( .A1(n4668), .A2(n4667), .ZN(n4300) );
  INV_X1 U5785 ( .A(n4555), .ZN(n9170) );
  NOR2_X1 U5786 ( .A1(n9197), .A2(n4556), .ZN(n4555) );
  INV_X1 U5787 ( .A(n4568), .ZN(n9259) );
  NOR2_X1 U5788 ( .A1(n9269), .A2(n9382), .ZN(n4568) );
  INV_X1 U5789 ( .A(n4792), .ZN(n4791) );
  NAND2_X1 U5790 ( .A1(n7872), .A2(n4278), .ZN(n4792) );
  AND2_X1 U5791 ( .A1(n5174), .A2(n5151), .ZN(n4301) );
  INV_X1 U5792 ( .A(n4671), .ZN(n4670) );
  NOR2_X1 U5793 ( .A1(n7574), .A2(n4672), .ZN(n4671) );
  AND2_X1 U5794 ( .A1(n8248), .A2(n8385), .ZN(n4302) );
  AND2_X1 U5795 ( .A1(n4285), .A2(n4385), .ZN(n4303) );
  AND2_X1 U5796 ( .A1(n8795), .A2(n8453), .ZN(n4304) );
  INV_X1 U5797 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8924) );
  NAND2_X1 U5798 ( .A1(n7090), .A2(n7053), .ZN(n7795) );
  INV_X1 U5799 ( .A(n7795), .ZN(n4834) );
  INV_X1 U5800 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4781) );
  AND2_X1 U5801 ( .A1(n7828), .A2(n7827), .ZN(n4305) );
  NAND2_X1 U5802 ( .A1(n5565), .A2(n5564), .ZN(n4306) );
  INV_X1 U5803 ( .A(n6617), .ZN(n4893) );
  INV_X1 U5804 ( .A(n9920), .ZN(n4449) );
  AND2_X1 U5805 ( .A1(n6825), .A2(n4425), .ZN(n4307) );
  NOR2_X1 U5806 ( .A1(n9385), .A2(n9113), .ZN(n4308) );
  INV_X1 U5807 ( .A(n8423), .ZN(n4443) );
  INV_X1 U5808 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5590) );
  INV_X1 U5809 ( .A(n4773), .ZN(n4772) );
  NAND2_X1 U5810 ( .A1(n4774), .A2(n8053), .ZN(n4773) );
  NOR2_X1 U5811 ( .A1(n9293), .A2(n9090), .ZN(n4309) );
  AND2_X1 U5812 ( .A1(n5889), .A2(n7422), .ZN(n4310) );
  AND2_X1 U5813 ( .A1(n5122), .A2(SI_11_), .ZN(n4311) );
  AND2_X1 U5814 ( .A1(n4966), .A2(SI_4_), .ZN(n4312) );
  NAND2_X1 U5815 ( .A1(n5034), .A2(n5033), .ZN(n4313) );
  AND2_X1 U5816 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n4314) );
  INV_X1 U5817 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6301) );
  INV_X1 U5818 ( .A(n4724), .ZN(n4723) );
  OR2_X1 U5819 ( .A1(n9046), .A2(n4725), .ZN(n4724) );
  NAND2_X1 U5820 ( .A1(n6043), .A2(n6042), .ZN(n9370) );
  NAND2_X1 U5821 ( .A1(n4818), .A2(n7567), .ZN(n4315) );
  AND2_X1 U5822 ( .A1(n5966), .A2(n5965), .ZN(n4316) );
  INV_X1 U5823 ( .A(n6767), .ZN(n4425) );
  AND2_X1 U5824 ( .A1(n5328), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n4317) );
  AND2_X1 U5825 ( .A1(n4717), .A2(n4715), .ZN(n4318) );
  AND2_X1 U5826 ( .A1(n4812), .A2(n4811), .ZN(n4319) );
  AND2_X1 U5827 ( .A1(n7093), .A2(n7173), .ZN(n4320) );
  AND2_X1 U5828 ( .A1(n4757), .A2(n8575), .ZN(n4321) );
  AND2_X1 U5829 ( .A1(n7737), .A2(n6937), .ZN(n4322) );
  AND2_X1 U5830 ( .A1(n8290), .A2(n8291), .ZN(n8410) );
  NOR2_X1 U5831 ( .A1(n7365), .A2(n4753), .ZN(n4752) );
  AND2_X1 U5832 ( .A1(n4522), .A2(n8924), .ZN(n4323) );
  AND2_X1 U5833 ( .A1(n7942), .A2(n4642), .ZN(n4324) );
  AND2_X1 U5834 ( .A1(n7070), .A2(n7069), .ZN(n4325) );
  AND2_X1 U5835 ( .A1(n8674), .A2(n4579), .ZN(n4326) );
  AND2_X1 U5836 ( .A1(n4782), .A2(n4781), .ZN(n4327) );
  AND2_X1 U5837 ( .A1(n4608), .A2(n8352), .ZN(n4328) );
  NAND2_X1 U5838 ( .A1(n4790), .A2(n7872), .ZN(n4789) );
  AND2_X1 U5839 ( .A1(n5263), .A2(n5241), .ZN(n4618) );
  INV_X1 U5840 ( .A(n4592), .ZN(n4591) );
  NAND2_X1 U5841 ( .A1(n4593), .A2(n4359), .ZN(n4592) );
  INV_X1 U5842 ( .A(n4694), .ZN(n4385) );
  AND2_X1 U5843 ( .A1(n9370), .A2(n9222), .ZN(n4694) );
  INV_X1 U5844 ( .A(n4779), .ZN(n4778) );
  NAND2_X1 U5845 ( .A1(n8423), .A2(n7598), .ZN(n4779) );
  INV_X1 U5846 ( .A(n7088), .ZN(n5535) );
  NAND2_X1 U5847 ( .A1(n6075), .A2(n6074), .ZN(n9355) );
  INV_X1 U5848 ( .A(n9355), .ZN(n4557) );
  NAND2_X1 U5849 ( .A1(n7775), .A2(n7774), .ZN(n9345) );
  INV_X1 U5850 ( .A(n9345), .ZN(n4553) );
  OR2_X1 U5851 ( .A1(n7569), .A2(n9499), .ZN(n4329) );
  AND2_X1 U5852 ( .A1(n8061), .A2(n8096), .ZN(n4330) );
  INV_X1 U5853 ( .A(n8017), .ZN(n4810) );
  NOR2_X1 U5854 ( .A1(n4553), .A2(n9179), .ZN(n4331) );
  NAND2_X1 U5855 ( .A1(n5385), .A2(n5384), .ZN(n8747) );
  INV_X1 U5856 ( .A(n8747), .ZN(n4478) );
  AND2_X1 U5857 ( .A1(n8771), .A2(n8647), .ZN(n4332) );
  AND2_X1 U5858 ( .A1(n6089), .A2(n6088), .ZN(n4333) );
  NAND2_X1 U5859 ( .A1(n4513), .A2(n7492), .ZN(n7491) );
  NOR3_X1 U5860 ( .A1(n7528), .A2(n4421), .A3(n4420), .ZN(n4419) );
  AND2_X1 U5861 ( .A1(n5449), .A2(n5448), .ZN(n4334) );
  INV_X1 U5862 ( .A(n8014), .ZN(n4808) );
  NOR2_X1 U5863 ( .A1(n7569), .A2(n4561), .ZN(n4564) );
  AND2_X1 U5864 ( .A1(n4404), .A2(n4402), .ZN(n4335) );
  NAND2_X1 U5865 ( .A1(n6058), .A2(n6059), .ZN(n4714) );
  INV_X1 U5866 ( .A(n4415), .ZN(n8625) );
  NOR2_X1 U5867 ( .A1(n8676), .A2(n4417), .ZN(n4415) );
  AND2_X1 U5868 ( .A1(n5540), .A2(n5539), .ZN(n4336) );
  NOR2_X1 U5869 ( .A1(n6029), .A2(n6028), .ZN(n4337) );
  INV_X1 U5870 ( .A(n4684), .ZN(n9402) );
  OR2_X1 U5871 ( .A1(n9311), .A2(n9310), .ZN(n4684) );
  OR2_X1 U5872 ( .A1(n7528), .A2(n7552), .ZN(n4338) );
  AND2_X1 U5873 ( .A1(n5346), .A2(n5327), .ZN(n4339) );
  AND2_X1 U5874 ( .A1(n9491), .A2(n7745), .ZN(n7576) );
  AND2_X1 U5875 ( .A1(n7599), .A2(n7598), .ZN(n4340) );
  AND2_X1 U5876 ( .A1(n4837), .A2(n4737), .ZN(n4341) );
  NOR2_X1 U5877 ( .A1(n6736), .A2(n7939), .ZN(n4342) );
  INV_X2 U5878 ( .A(n9942), .ZN(n9944) );
  INV_X1 U5879 ( .A(n9499), .ZN(n4563) );
  INV_X1 U5880 ( .A(n7492), .ZN(n4512) );
  AND2_X1 U5881 ( .A1(n6850), .A2(n4960), .ZN(n4343) );
  INV_X2 U5882 ( .A(n9952), .ZN(n9954) );
  OR2_X1 U5883 ( .A1(n5494), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4344) );
  NAND2_X1 U5884 ( .A1(n4378), .A2(n7042), .ZN(n9679) );
  AND2_X1 U5885 ( .A1(n8316), .A2(n8315), .ZN(n8419) );
  INV_X1 U5886 ( .A(n8419), .ZN(n4755) );
  INV_X1 U5887 ( .A(n4973), .ZN(n5000) );
  AND2_X1 U5888 ( .A1(n9478), .A2(n9475), .ZN(n9854) );
  INV_X1 U5889 ( .A(n4637), .ZN(n4636) );
  NOR2_X1 U5890 ( .A1(n5432), .A2(n4638), .ZN(n4637) );
  AND2_X1 U5891 ( .A1(n7416), .A2(n7441), .ZN(n4345) );
  NAND2_X1 U5892 ( .A1(n7126), .A2(n4422), .ZN(n4426) );
  INV_X1 U5893 ( .A(n4549), .ZN(n7251) );
  NOR2_X1 U5894 ( .A1(n7252), .A2(n7265), .ZN(n4549) );
  NAND2_X1 U5895 ( .A1(n5834), .A2(n5833), .ZN(n4346) );
  NAND2_X1 U5896 ( .A1(n4574), .A2(n8294), .ZN(n4347) );
  NOR2_X1 U5897 ( .A1(n5815), .A2(n7148), .ZN(n5816) );
  XNOR2_X1 U5898 ( .A(n4865), .B(n4877), .ZN(n5534) );
  AND2_X1 U5899 ( .A1(n9707), .A2(n9748), .ZN(n9425) );
  NAND2_X1 U5900 ( .A1(n5139), .A2(n5138), .ZN(n7361) );
  INV_X1 U5901 ( .A(n7361), .ZN(n4548) );
  INV_X1 U5902 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4462) );
  INV_X1 U5903 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5575) );
  NAND2_X1 U5904 ( .A1(n4854), .A2(n4853), .ZN(n8583) );
  INV_X1 U5905 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4847) );
  INV_X1 U5906 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n4361) );
  MUX2_X1 U5907 ( .A(n7863), .B(n7862), .S(n7897), .Z(n7866) );
  MUX2_X1 U5908 ( .A(n7871), .B(n7870), .S(n7897), .Z(n7879) );
  NAND2_X1 U5909 ( .A1(n7856), .A2(n7855), .ZN(n7861) );
  NAND2_X1 U5910 ( .A1(n6727), .A2(n4377), .ZN(n6726) );
  NAND2_X1 U5911 ( .A1(n7908), .A2(n6728), .ZN(n6938) );
  NOR3_X1 U5912 ( .A1(n7938), .A2(n7974), .A3(n7899), .ZN(n7933) );
  AOI21_X1 U5913 ( .B1(n4655), .B2(n4654), .A(n7891), .ZN(n7892) );
  NAND2_X1 U5914 ( .A1(n7845), .A2(n4348), .ZN(n4374) );
  NAND2_X1 U5915 ( .A1(n7824), .A2(n7823), .ZN(n7845) );
  NAND2_X1 U5916 ( .A1(n4350), .A2(n7985), .ZN(P1_U3240) );
  NAND2_X1 U5917 ( .A1(n4352), .A2(n4351), .ZN(n4350) );
  NAND2_X1 U5918 ( .A1(n4641), .A2(n4640), .ZN(n4352) );
  MUX2_X1 U5919 ( .A(n7888), .B(n7900), .S(n7897), .Z(n7894) );
  AOI21_X1 U5920 ( .B1(n9072), .B2(n9075), .A(n9074), .ZN(n6057) );
  AOI21_X2 U5921 ( .B1(n8978), .B2(n8980), .A(n8977), .ZN(n9054) );
  NAND2_X1 U5922 ( .A1(n6112), .A2(n6113), .ZN(n9013) );
  NAND2_X1 U5923 ( .A1(n6703), .A2(n6702), .ZN(n6701) );
  NAND2_X1 U5924 ( .A1(n9062), .A2(n4718), .ZN(n4716) );
  NOR2_X2 U5925 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n4353) );
  NAND2_X1 U5926 ( .A1(n7620), .A2(n7618), .ZN(n7623) );
  NAND2_X1 U5927 ( .A1(n8987), .A2(n6002), .ZN(n9062) );
  NAND2_X1 U5928 ( .A1(n4703), .A2(n4704), .ZN(n6112) );
  NAND2_X1 U5929 ( .A1(n5649), .A2(n5650), .ZN(n9020) );
  NAND2_X1 U5930 ( .A1(n5631), .A2(n6432), .ZN(n5649) );
  NAND2_X1 U5931 ( .A1(n4362), .A2(n9013), .ZN(n6135) );
  NAND2_X1 U5932 ( .A1(n5925), .A2(n5924), .ZN(n7620) );
  NAND2_X1 U5933 ( .A1(n7657), .A2(n7661), .ZN(n7686) );
  INV_X1 U5934 ( .A(n4729), .ZN(n5984) );
  NOR2_X1 U5935 ( .A1(n6057), .A2(n6056), .ZN(n8977) );
  NAND2_X1 U5936 ( .A1(n6680), .A2(n5717), .ZN(n5733) );
  NAND2_X1 U5937 ( .A1(n6525), .A2(n5674), .ZN(n6532) );
  OAI21_X2 U5938 ( .B1(n5578), .B2(n4409), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5560) );
  NAND2_X1 U5939 ( .A1(n7660), .A2(n7659), .ZN(n7657) );
  NAND3_X1 U5940 ( .A1(n5585), .A2(n6127), .A3(n5584), .ZN(n6165) );
  NAND2_X1 U5941 ( .A1(n5326), .A2(n5325), .ZN(n4524) );
  NAND2_X1 U5942 ( .A1(n5381), .A2(n5380), .ZN(n5383) );
  NAND2_X1 U5943 ( .A1(n5349), .A2(n5348), .ZN(n5371) );
  NAND2_X1 U5944 ( .A1(n5079), .A2(n4838), .ZN(n5081) );
  NAND2_X1 U5945 ( .A1(n8081), .A2(n8066), .ZN(n8227) );
  NAND2_X1 U5946 ( .A1(n8988), .A2(n8989), .ZN(n8987) );
  NAND2_X1 U5947 ( .A1(n5652), .A2(n5651), .ZN(n9021) );
  NAND2_X1 U5948 ( .A1(n8692), .A2(n8704), .ZN(n8691) );
  NAND2_X1 U5949 ( .A1(n6579), .A2(n8407), .ZN(n6743) );
  NAND2_X1 U5950 ( .A1(n7068), .A2(n7067), .ZN(n4762) );
  NAND2_X1 U5951 ( .A1(n6956), .A2(n6955), .ZN(n7066) );
  INV_X1 U5952 ( .A(n6584), .ZN(n4375) );
  AOI21_X2 U5953 ( .B1(n8639), .B2(n8055), .A(n8054), .ZN(n8624) );
  OAI21_X2 U5954 ( .B1(n8724), .B2(n8785), .A(n4373), .ZN(n4546) );
  NAND2_X1 U5955 ( .A1(n7433), .A2(n4598), .ZN(n4597) );
  NAND2_X1 U5956 ( .A1(n7601), .A2(n8330), .ZN(n7632) );
  NAND2_X1 U5957 ( .A1(n4273), .A2(n6776), .ZN(n6956) );
  NAND2_X1 U5958 ( .A1(n4748), .A2(n4280), .ZN(n7440) );
  NAND2_X1 U5959 ( .A1(n4576), .A2(n4577), .ZN(n6778) );
  INV_X1 U5960 ( .A(n4603), .ZN(n8609) );
  NAND2_X1 U5961 ( .A1(n4749), .A2(n4752), .ZN(n4748) );
  NAND2_X1 U5962 ( .A1(n7237), .A2(n7236), .ZN(n7247) );
  NAND2_X1 U5963 ( .A1(n4758), .A2(n4321), .ZN(n8574) );
  NAND2_X2 U5964 ( .A1(n4924), .A2(n4923), .ZN(n4942) );
  NAND2_X1 U5965 ( .A1(n8377), .A2(n8546), .ZN(n4464) );
  NAND2_X1 U5966 ( .A1(n8370), .A2(n8372), .ZN(n4467) );
  INV_X1 U5967 ( .A(n4429), .ZN(n4435) );
  INV_X1 U5968 ( .A(n4434), .ZN(n4431) );
  OAI21_X1 U5969 ( .B1(n4454), .B2(n4453), .A(n8608), .ZN(n4452) );
  NAND2_X1 U5970 ( .A1(n8344), .A2(n8075), .ZN(n4458) );
  NAND2_X1 U5971 ( .A1(n4433), .A2(n8337), .ZN(n8347) );
  NOR2_X1 U5972 ( .A1(n8438), .A2(n4444), .ZN(n8439) );
  NAND2_X1 U5973 ( .A1(n4367), .A2(n7797), .ZN(n7802) );
  NAND3_X1 U5974 ( .A1(n7794), .A2(n7795), .A3(n7799), .ZN(n4367) );
  NOR3_X2 U5975 ( .A1(n7889), .A2(n7886), .A3(n9160), .ZN(n7887) );
  MUX2_X1 U5976 ( .A(n7852), .B(n7851), .S(n7897), .Z(n7853) );
  OAI21_X2 U5977 ( .B1(n7896), .B2(n7895), .A(n4368), .ZN(n7938) );
  NAND3_X2 U5978 ( .A1(n5667), .A2(n5666), .A3(n4282), .ZN(n6936) );
  OAI21_X1 U5979 ( .B1(n7933), .B2(n4643), .A(n4324), .ZN(n4641) );
  NAND2_X1 U5980 ( .A1(n4716), .A2(n4717), .ZN(n6041) );
  NOR2_X1 U5981 ( .A1(n5816), .A2(n4700), .ZN(n4699) );
  NAND2_X1 U5982 ( .A1(n5580), .A2(n5557), .ZN(n5574) );
  NAND2_X1 U5983 ( .A1(n7230), .A2(n7229), .ZN(n7228) );
  NAND2_X1 U5984 ( .A1(n8574), .A2(n8059), .ZN(n8555) );
  NAND2_X2 U5985 ( .A1(n8691), .A2(n8051), .ZN(n8675) );
  NAND2_X1 U5986 ( .A1(n8537), .A2(n8536), .ZN(n8535) );
  NAND2_X1 U5987 ( .A1(n4546), .A2(n9954), .ZN(n4545) );
  OAI21_X1 U5988 ( .B1(n8504), .B2(n8569), .A(n4531), .ZN(P2_U3264) );
  OAI21_X1 U5989 ( .B1(n8503), .B2(n8500), .A(n8499), .ZN(n4533) );
  NAND2_X1 U5990 ( .A1(n4374), .A2(n7846), .ZN(n7839) );
  MUX2_X2 U5991 ( .A(n7802), .B(n7801), .S(n7881), .Z(n7814) );
  NAND2_X1 U5992 ( .A1(n7889), .A2(n8028), .ZN(n4655) );
  AND2_X4 U5993 ( .A1(n5136), .A2(n4844), .ZN(n5178) );
  NAND2_X1 U5994 ( .A1(n8519), .A2(n4766), .ZN(n4765) );
  AND2_X2 U5995 ( .A1(n8603), .A2(n8604), .ZN(n8607) );
  NAND2_X1 U5996 ( .A1(n4545), .A2(n4544), .ZN(P2_U3549) );
  NAND3_X1 U5997 ( .A1(n7946), .A2(n7945), .A3(n4377), .ZN(n7951) );
  OAI21_X1 U5998 ( .B1(n9679), .B2(n9680), .A(n7045), .ZN(n7048) );
  NAND2_X1 U5999 ( .A1(n7041), .A2(n7907), .ZN(n4378) );
  NAND2_X1 U6000 ( .A1(n6930), .A2(n6929), .ZN(n7041) );
  INV_X1 U6001 ( .A(n8005), .ZN(n4384) );
  OR2_X1 U6002 ( .A1(n9377), .A2(n9112), .ZN(n4386) );
  NAND2_X1 U6003 ( .A1(n9311), .A2(n4392), .ZN(n4389) );
  NAND2_X1 U6004 ( .A1(n4389), .A2(n4391), .ZN(n8004) );
  NAND2_X1 U6005 ( .A1(n9154), .A2(n4398), .ZN(n4396) );
  NAND2_X1 U6006 ( .A1(n9154), .A2(n4688), .ZN(n4397) );
  OAI211_X1 U6007 ( .C1(n9154), .C2(n4399), .A(n4396), .B(n4406), .ZN(P1_U3552) );
  OAI211_X1 U6008 ( .C1(n9154), .C2(n4690), .A(n4689), .B(n4397), .ZN(n9344)
         );
  INV_X1 U6009 ( .A(n5578), .ZN(n4407) );
  OAI21_X1 U6010 ( .B1(n4407), .B2(n5934), .A(n4408), .ZN(n5558) );
  NOR2_X2 U6011 ( .A1(n5577), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n5580) );
  INV_X1 U6012 ( .A(n4419), .ZN(n8695) );
  INV_X1 U6013 ( .A(n4426), .ZN(n6959) );
  OAI21_X1 U6014 ( .B1(n8318), .B2(n4431), .A(n4430), .ZN(n4433) );
  INV_X1 U6015 ( .A(n4432), .ZN(n4439) );
  NAND2_X1 U6016 ( .A1(n8632), .A2(n8357), .ZN(n4453) );
  AOI21_X1 U6017 ( .B1(n4458), .B2(n4456), .A(n4455), .ZN(n4454) );
  AND2_X1 U6018 ( .A1(n5178), .A2(n4877), .ZN(n4460) );
  NAND2_X1 U6019 ( .A1(n4459), .A2(n4780), .ZN(n8965) );
  NAND2_X1 U6020 ( .A1(n4463), .A2(n4465), .ZN(n8379) );
  NAND2_X1 U6021 ( .A1(n4464), .A2(n4466), .ZN(n4463) );
  NAND2_X1 U6022 ( .A1(n5410), .A2(n4476), .ZN(n8140) );
  INV_X1 U6023 ( .A(n8135), .ZN(n4475) );
  OAI21_X1 U6024 ( .B1(n5543), .B2(n8725), .A(n4479), .ZN(P2_U3222) );
  AOI21_X1 U6025 ( .B1(n5542), .B2(n4482), .A(n4480), .ZN(n4479) );
  INV_X1 U6026 ( .A(n4493), .ZN(n4854) );
  NAND2_X1 U6027 ( .A1(n4942), .A2(n4941), .ZN(n4499) );
  NAND2_X1 U6028 ( .A1(n4942), .A2(n4290), .ZN(n4496) );
  NAND2_X1 U6029 ( .A1(n5081), .A2(n4501), .ZN(n4500) );
  NAND2_X1 U6030 ( .A1(n5081), .A2(n5080), .ZN(n5102) );
  NAND2_X1 U6031 ( .A1(n4509), .A2(n4510), .ZN(n5284) );
  NAND3_X1 U6032 ( .A1(n5219), .A2(n7544), .A3(n4618), .ZN(n4509) );
  NAND2_X1 U6033 ( .A1(n9855), .A2(n4518), .ZN(n4517) );
  NAND2_X1 U6034 ( .A1(n4524), .A2(n4339), .ZN(n5349) );
  INV_X1 U6035 ( .A(n4537), .ZN(n6237) );
  INV_X1 U6036 ( .A(n4535), .ZN(n6252) );
  NAND2_X1 U6037 ( .A1(n4537), .A2(n4536), .ZN(n4535) );
  AND2_X2 U6038 ( .A1(n6195), .A2(n5561), .ZN(n4902) );
  NAND2_X2 U6039 ( .A1(n8441), .A2(n5534), .ZN(n6195) );
  NAND2_X1 U6040 ( .A1(n9952), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n4544) );
  NAND3_X1 U6041 ( .A1(n5555), .A2(n4551), .A3(n4837), .ZN(n5577) );
  INV_X2 U6042 ( .A(n5741), .ZN(n4837) );
  NAND3_X1 U6043 ( .A1(n5555), .A2(n4837), .A3(n4264), .ZN(n6128) );
  INV_X2 U6044 ( .A(n6714), .ZN(n9719) );
  INV_X1 U6045 ( .A(n4564), .ZN(n9322) );
  OAI21_X1 U6046 ( .B1(n7073), .B2(n4572), .A(n4569), .ZN(n7240) );
  INV_X1 U6047 ( .A(n8294), .ZN(n4575) );
  NAND2_X1 U6048 ( .A1(n6778), .A2(n6777), .ZN(n6957) );
  NAND2_X1 U6049 ( .A1(n7119), .A2(n7118), .ZN(n4577) );
  NAND2_X1 U6050 ( .A1(n4578), .A2(n4326), .ZN(n8074) );
  NAND2_X1 U6051 ( .A1(n7635), .A2(n4580), .ZN(n4578) );
  NAND2_X1 U6052 ( .A1(n4597), .A2(n4595), .ZN(n7601) );
  NOR2_X1 U6053 ( .A1(n4317), .A2(n4601), .ZN(n4600) );
  NOR2_X1 U6054 ( .A1(n6195), .A2(n6306), .ZN(n4601) );
  OAI21_X1 U6055 ( .B1(n8653), .B2(n4606), .A(n4604), .ZN(n4603) );
  OR2_X1 U6056 ( .A1(n8436), .A2(n7088), .ZN(n8240) );
  NAND2_X1 U6057 ( .A1(n8444), .A2(n8583), .ZN(n6580) );
  NAND2_X1 U6058 ( .A1(n7088), .A2(n8255), .ZN(n4609) );
  NAND3_X1 U6059 ( .A1(n8436), .A2(n8444), .A3(n8583), .ZN(n4610) );
  NAND2_X1 U6060 ( .A1(n6618), .A2(n4895), .ZN(n4614) );
  NAND3_X1 U6061 ( .A1(n4615), .A2(n4614), .A3(n6844), .ZN(n6838) );
  NAND2_X1 U6062 ( .A1(n6617), .A2(n4895), .ZN(n4615) );
  AOI21_X1 U6063 ( .B1(n8528), .B2(n8428), .A(n8080), .ZN(n8081) );
  INV_X1 U6064 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4742) );
  OAI21_X1 U6065 ( .B1(n8230), .B2(n8229), .A(n8228), .ZN(n8236) );
  BUF_X4 U6066 ( .A(n4870), .Z(n7715) );
  NOR2_X1 U6067 ( .A1(n8723), .A2(n7135), .ZN(n8088) );
  NAND2_X1 U6068 ( .A1(n4622), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4658) );
  NAND2_X1 U6069 ( .A1(n5517), .A2(n4627), .ZN(n4625) );
  NAND2_X2 U6070 ( .A1(n4657), .A2(n4656), .ZN(n4870) );
  NAND2_X1 U6071 ( .A1(n7384), .A2(n7917), .ZN(n7562) );
  INV_X1 U6072 ( .A(n7382), .ZN(n4663) );
  NAND2_X1 U6073 ( .A1(n4681), .A2(n4680), .ZN(n7098) );
  AOI21_X1 U6074 ( .B1(n7912), .B2(n4682), .A(n4320), .ZN(n4680) );
  NAND3_X1 U6075 ( .A1(n7046), .A2(n7912), .A3(n7047), .ZN(n4681) );
  OAI21_X1 U6076 ( .B1(n9344), .B2(n4687), .A(n4685), .ZN(P1_U3520) );
  NAND2_X1 U6077 ( .A1(n4695), .A2(n9084), .ZN(n8988) );
  NAND2_X1 U6078 ( .A1(n9085), .A2(n9083), .ZN(n4695) );
  NOR2_X1 U6079 ( .A1(n9082), .A2(n4695), .ZN(n9088) );
  OAI21_X1 U6080 ( .B1(n6526), .B2(n4696), .A(n6525), .ZN(n6527) );
  NAND2_X1 U6081 ( .A1(n4696), .A2(n6526), .ZN(n6525) );
  AND2_X1 U6082 ( .A1(n5653), .A2(n9021), .ZN(n4696) );
  NAND4_X1 U6083 ( .A1(n5660), .A2(n5544), .A3(n5545), .A4(n5724), .ZN(n5741)
         );
  NAND2_X1 U6084 ( .A1(n9054), .A2(n4277), .ZN(n4703) );
  NAND2_X1 U6085 ( .A1(n9054), .A2(n9055), .ZN(n9053) );
  NAND2_X1 U6086 ( .A1(n6073), .A2(n6072), .ZN(n4713) );
  INV_X1 U6087 ( .A(n5951), .ZN(n4734) );
  OAI21_X1 U6088 ( .B1(n4734), .B2(n5934), .A(n4735), .ZN(n5567) );
  NAND2_X1 U6089 ( .A1(n4264), .A2(n5548), .ZN(n4738) );
  NAND4_X1 U6090 ( .A1(n4843), .A2(n4741), .A3(n4740), .A4(n4739), .ZN(n4743)
         );
  NAND3_X1 U6091 ( .A1(n4842), .A2(n4903), .A3(n4742), .ZN(n4949) );
  NOR2_X2 U6092 ( .A1(n4949), .A2(n4743), .ZN(n5136) );
  NAND2_X1 U6093 ( .A1(n7124), .A2(n4746), .ZN(n4745) );
  INV_X1 U6094 ( .A(n7247), .ZN(n4749) );
  NAND2_X1 U6095 ( .A1(n8607), .A2(n8058), .ZN(n4758) );
  NAND2_X1 U6096 ( .A1(n4762), .A2(n4325), .ZN(n7237) );
  OAI211_X2 U6097 ( .C1(n8519), .C2(n8430), .A(n4767), .B(n4765), .ZN(n8724)
         );
  OAI21_X2 U6098 ( .B1(n8675), .B2(n4773), .A(n4770), .ZN(n8639) );
  INV_X1 U6099 ( .A(n9248), .ZN(n4796) );
  NAND2_X1 U6100 ( .A1(n9248), .A2(n4789), .ZN(n4785) );
  NAND2_X1 U6101 ( .A1(n9297), .A2(n4800), .ZN(n4799) );
  AND2_X2 U6102 ( .A1(n5580), .A2(n4319), .ZN(n5596) );
  NAND2_X1 U6103 ( .A1(n6938), .A2(n4322), .ZN(n7056) );
  NOR2_X1 U6104 ( .A1(n7952), .A2(n4813), .ZN(n7751) );
  XNOR2_X1 U6105 ( .A(n4815), .B(n4814), .ZN(n9705) );
  NAND2_X1 U6106 ( .A1(n7188), .A2(n7757), .ZN(n4820) );
  NAND2_X1 U6107 ( .A1(n4820), .A2(n4821), .ZN(n9510) );
  INV_X1 U6108 ( .A(n9189), .ZN(n4823) );
  NAND2_X1 U6109 ( .A1(n4831), .A2(n4828), .ZN(n4830) );
  NAND2_X1 U6110 ( .A1(n9673), .A2(n4276), .ZN(n4835) );
  OR2_X2 U6111 ( .A1(n9673), .A2(n7058), .ZN(n4836) );
  AND2_X2 U6112 ( .A1(n4836), .A2(n7743), .ZN(n7798) );
  INV_X8 U6113 ( .A(n4870), .ZN(n5561) );
  XNOR2_X2 U6114 ( .A(n5399), .B(n5398), .ZN(n8103) );
  NAND2_X1 U6115 ( .A1(n5571), .A2(n5586), .ZN(n6133) );
  CLKBUF_X1 U6116 ( .A(n6863), .Z(n7146) );
  INV_X1 U6117 ( .A(n5649), .ZN(n5652) );
  CLKBUF_X1 U6118 ( .A(n6726), .Z(n9724) );
  OAI21_X1 U6119 ( .B1(n9274), .B2(n9286), .A(n8004), .ZN(n9254) );
  BUF_X4 U6120 ( .A(n4902), .Z(n5328) );
  NAND2_X2 U6121 ( .A1(n6882), .A2(n8679), .ZN(n8688) );
  INV_X1 U6122 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5559) );
  NAND2_X2 U6123 ( .A1(n7175), .A2(n9709), .ZN(n9737) );
  INV_X1 U6124 ( .A(n7939), .ZN(n7940) );
  AND2_X1 U6125 ( .A1(n5080), .A2(n5062), .ZN(n4838) );
  AND2_X1 U6126 ( .A1(n5103), .A2(n5086), .ZN(n4839) );
  AND2_X1 U6127 ( .A1(n5176), .A2(n5159), .ZN(n4840) );
  INV_X1 U6128 ( .A(n9560), .ZN(n5634) );
  INV_X1 U6129 ( .A(n8725), .ZN(n8061) );
  INV_X1 U6130 ( .A(n8430), .ZN(n8066) );
  NOR2_X1 U6131 ( .A1(n5163), .A2(n5141), .ZN(n4841) );
  AOI21_X1 U6132 ( .B1(n8525), .B2(n5532), .A(n5480), .ZN(n8096) );
  INV_X1 U6133 ( .A(n7911), .ZN(n7096) );
  NAND2_X1 U6134 ( .A1(n5284), .A2(n8199), .ZN(n8111) );
  INV_X1 U6135 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5548) );
  INV_X1 U6136 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5546) );
  XNOR2_X1 U6137 ( .A(n5709), .B(n5646), .ZN(n5650) );
  INV_X1 U6138 ( .A(n9494), .ZN(n7567) );
  NAND2_X1 U6139 ( .A1(n6713), .A2(n9719), .ZN(n6727) );
  INV_X1 U6140 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5082) );
  INV_X1 U6141 ( .A(n5358), .ZN(n5356) );
  INV_X1 U6142 ( .A(n5274), .ZN(n5273) );
  INV_X1 U6143 ( .A(n5213), .ZN(n5212) );
  INV_X1 U6144 ( .A(n5402), .ZN(n5386) );
  INV_X1 U6145 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n4855) );
  INV_X1 U6146 ( .A(n5625), .ZN(n5637) );
  INV_X1 U6147 ( .A(n5627), .ZN(n5628) );
  INV_X1 U6148 ( .A(n5650), .ZN(n5651) );
  INV_X1 U6149 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5566) );
  INV_X1 U6150 ( .A(SI_12_), .ZN(n5125) );
  INV_X1 U6151 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5785) );
  INV_X1 U6152 ( .A(n6762), .ZN(n5021) );
  INV_X1 U6153 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5001) );
  OR2_X1 U6154 ( .A1(n5232), .A2(n8840), .ZN(n5253) );
  AND2_X1 U6155 ( .A1(n5140), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5163) );
  NAND2_X1 U6156 ( .A1(n5273), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5297) );
  AOI21_X1 U6157 ( .B1(n8236), .B2(n8400), .A(n8395), .ZN(n8237) );
  OR2_X1 U6158 ( .A1(n5441), .A2(n5440), .ZN(n5461) );
  NOR2_X1 U6159 ( .A1(n4975), .A2(n4974), .ZN(n4989) );
  OR2_X1 U6160 ( .A1(n8742), .A2(n8450), .ZN(n8059) );
  AND2_X1 U6161 ( .A1(n9886), .A2(n6619), .ZN(n6877) );
  INV_X1 U6162 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7625) );
  INV_X1 U6163 ( .A(n5923), .ZN(n5924) );
  NAND2_X1 U6164 ( .A1(n5623), .A2(n5622), .ZN(n5624) );
  INV_X1 U6165 ( .A(n9458), .ZN(n5867) );
  NAND2_X1 U6166 ( .A1(n4270), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5667) );
  INV_X1 U6167 ( .A(n8041), .ZN(n7931) );
  OR2_X1 U6168 ( .A1(n5954), .A2(n9047), .ZN(n5974) );
  AND2_X1 U6169 ( .A1(n5912), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5939) );
  OR2_X1 U6170 ( .A1(n9683), .A2(n9687), .ZN(n9684) );
  INV_X1 U6171 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5557) );
  OR2_X1 U6172 ( .A1(n5400), .A2(n8106), .ZN(n5402) );
  INV_X1 U6173 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5066) );
  INV_X1 U6174 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5043) );
  NAND2_X1 U6175 ( .A1(n5251), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5274) );
  AND2_X1 U6176 ( .A1(n8467), .A2(n9898), .ZN(n6889) );
  INV_X1 U6177 ( .A(n7325), .ZN(n5174) );
  AND2_X1 U6178 ( .A1(n5526), .A2(n5476), .ZN(n8525) );
  OR2_X1 U6179 ( .A1(n5316), .A2(n6174), .ZN(n5333) );
  INV_X1 U6180 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8820) );
  NAND2_X1 U6181 ( .A1(n6877), .A2(n6876), .ZN(n6882) );
  INV_X1 U6182 ( .A(n8659), .ZN(n8707) );
  NAND2_X1 U6183 ( .A1(n5513), .A2(n5512), .ZN(n5489) );
  AND2_X1 U6184 ( .A1(n5600), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6062) );
  NOR2_X1 U6185 ( .A1(n5840), .A2(n5839), .ZN(n5856) );
  OR2_X1 U6186 ( .A1(n5733), .A2(n5732), .ZN(n5734) );
  NAND2_X1 U6187 ( .A1(n6134), .A2(n7931), .ZN(n7899) );
  AND2_X1 U6188 ( .A1(n7782), .A2(n6152), .ZN(n9158) );
  AND2_X1 U6189 ( .A1(n6032), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6044) );
  INV_X1 U6190 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6445) );
  OR2_X1 U6191 ( .A1(n9553), .A2(n6423), .ZN(n9658) );
  INV_X1 U6192 ( .A(n9370), .ZN(n9233) );
  INV_X1 U6193 ( .A(n9115), .ZN(n9319) );
  INV_X1 U6194 ( .A(n9116), .ZN(n7690) );
  OR2_X1 U6195 ( .A1(n5878), .A2(n5877), .ZN(n5898) );
  INV_X1 U6196 ( .A(n9137), .ZN(n9721) );
  NAND2_X1 U6197 ( .A1(n9737), .A2(n4342), .ZN(n9710) );
  INV_X1 U6198 ( .A(n9801), .ZN(n9717) );
  INV_X1 U6199 ( .A(n9799), .ZN(n9422) );
  INV_X1 U6200 ( .A(n9704), .ZN(n9733) );
  NAND2_X1 U6201 ( .A1(n6167), .A2(n9450), .ZN(n5619) );
  INV_X1 U6202 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5934) );
  OR3_X1 U6203 ( .A1(n7335), .A2(n7536), .A3(n7542), .ZN(n6181) );
  OR2_X1 U6204 ( .A1(n5182), .A2(n8820), .ZN(n5213) );
  OR2_X1 U6205 ( .A1(n5044), .A2(n5043), .ZN(n5067) );
  XNOR2_X1 U6206 ( .A(n6842), .B(n4894), .ZN(n6618) );
  OR2_X1 U6207 ( .A1(n6179), .A2(n6186), .ZN(n8564) );
  AND2_X1 U6208 ( .A1(n8444), .A2(n8255), .ZN(n6581) );
  INV_X1 U6209 ( .A(n8656), .ZN(n8562) );
  AND2_X1 U6210 ( .A1(n5427), .A2(n5426), .ZN(n8561) );
  AND4_X1 U6211 ( .A1(n5258), .A2(n5257), .A3(n5256), .A4(n5255), .ZN(n8203)
         );
  INV_X1 U6212 ( .A(n6974), .ZN(n6968) );
  AND2_X1 U6213 ( .A1(n6192), .A2(n8441), .ZN(n9871) );
  AND2_X1 U6214 ( .A1(n6190), .A2(n5534), .ZN(n9876) );
  INV_X1 U6215 ( .A(n8711), .ZN(n8662) );
  AND2_X1 U6216 ( .A1(n6581), .A2(n6186), .ZN(n8656) );
  OR2_X1 U6217 ( .A1(n9892), .A2(n5501), .ZN(n6875) );
  AND2_X1 U6218 ( .A1(n7600), .A2(n7480), .ZN(n8785) );
  INV_X1 U6219 ( .A(n8785), .ZN(n9931) );
  OR2_X1 U6220 ( .A1(n6572), .A2(n6571), .ZN(n6609) );
  INV_X1 U6221 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5012) );
  INV_X1 U6222 ( .A(n7783), .ZN(n6038) );
  OR2_X1 U6223 ( .A1(n5991), .A2(n5695), .ZN(n5696) );
  INV_X1 U6224 ( .A(n9658), .ZN(n9636) );
  INV_X1 U6225 ( .A(n9632), .ZN(n9661) );
  INV_X1 U6226 ( .A(n9145), .ZN(n9330) );
  NAND2_X1 U6227 ( .A1(n8024), .A2(n8023), .ZN(n9205) );
  AND2_X1 U6228 ( .A1(n9737), .A2(n9137), .ZN(n9260) );
  INV_X1 U6229 ( .A(n9709), .ZN(n9718) );
  INV_X1 U6230 ( .A(n9699), .ZN(n9729) );
  AND2_X1 U6231 ( .A1(n6136), .A2(n6311), .ZN(n6479) );
  OR2_X1 U6232 ( .A1(n6736), .A2(n7940), .ZN(n9801) );
  INV_X1 U6233 ( .A(n9425), .ZN(n9805) );
  AND2_X1 U6234 ( .A1(n6479), .A2(n6478), .ZN(n6721) );
  NAND2_X1 U6235 ( .A1(n6165), .A2(n6131), .ZN(n6722) );
  INV_X1 U6236 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5572) );
  AND2_X1 U6237 ( .A1(n5908), .A2(n5895), .ZN(n9624) );
  INV_X1 U6238 ( .A(n8506), .ZN(n9870) );
  OR2_X1 U6239 ( .A1(n8209), .A2(n8564), .ZN(n8219) );
  INV_X1 U6240 ( .A(n8563), .ZN(n8530) );
  INV_X1 U6241 ( .A(n8057), .ZN(n8634) );
  AND4_X1 U6242 ( .A1(n5218), .A2(n5217), .A3(n5216), .A4(n5215), .ZN(n7602)
         );
  INV_X1 U6243 ( .A(n9876), .ZN(n9861) );
  INV_X1 U6244 ( .A(n9871), .ZN(n9862) );
  AND2_X1 U6245 ( .A1(n7606), .A2(n7605), .ZN(n8800) );
  OR2_X1 U6246 ( .A1(n6609), .A2(n6875), .ZN(n9952) );
  OR2_X1 U6247 ( .A1(n6609), .A2(n6573), .ZN(n9942) );
  NAND2_X1 U6248 ( .A1(n9886), .A2(n9885), .ZN(n9890) );
  INV_X1 U6249 ( .A(n4881), .ZN(n8973) );
  XNOR2_X1 U6250 ( .A(n5491), .B(n5490), .ZN(n7335) );
  INV_X1 U6251 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6544) );
  INV_X1 U6252 ( .A(n8967), .ZN(n8971) );
  INV_X1 U6253 ( .A(n9391), .ZN(n9293) );
  NAND2_X1 U6254 ( .A1(n6139), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9468) );
  INV_X1 U6255 ( .A(n7388), .ZN(n9535) );
  INV_X1 U6256 ( .A(n9086), .ZN(n9460) );
  OR2_X1 U6257 ( .A1(n9553), .A2(n6141), .ZN(n9627) );
  INV_X1 U6258 ( .A(n9663), .ZN(n9621) );
  INV_X1 U6259 ( .A(n9696), .ZN(n9153) );
  NAND2_X1 U6260 ( .A1(n9737), .A2(n9682), .ZN(n9329) );
  AND2_X2 U6261 ( .A1(n6429), .A2(n6479), .ZN(n9826) );
  OR3_X1 U6262 ( .A1(n9418), .A2(n9417), .A3(n9416), .ZN(n9441) );
  AND2_X2 U6263 ( .A1(n6721), .A2(n6481), .ZN(n9809) );
  INV_X1 U6264 ( .A(n6722), .ZN(n6311) );
  NAND2_X1 U6265 ( .A1(n6311), .A2(n6475), .ZN(n9744) );
  INV_X1 U6266 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n8935) );
  INV_X1 U6267 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6336) );
  NOR2_X1 U6268 ( .A1(n9996), .A2(n9995), .ZN(n9994) );
  NOR2_X1 U6269 ( .A1(n9982), .A2(n9981), .ZN(n9980) );
  AND2_X1 U6270 ( .A1(n6169), .A2(n9893), .ZN(P2_U3966) );
  NOR2_X1 U6271 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n4843) );
  NAND2_X1 U6272 ( .A1(n4847), .A2(n4846), .ZN(n4848) );
  NAND2_X1 U6273 ( .A1(n4851), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4850) );
  NOR2_X1 U6274 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n4858) );
  NOR2_X1 U6275 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n4857) );
  NOR2_X1 U6276 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n4856) );
  NAND4_X1 U6277 ( .A1(n4858), .A2(n4857), .A3(n4856), .A4(n4855), .ZN(n4862)
         );
  NAND4_X1 U6278 ( .A1(n4860), .A2(n4859), .A3(n8924), .A4(n5486), .ZN(n4861)
         );
  NOR2_X1 U6279 ( .A1(n4862), .A2(n4861), .ZN(n4863) );
  NAND2_X1 U6280 ( .A1(n6195), .A2(n7715), .ZN(n4869) );
  AND2_X1 U6281 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4871) );
  NAND2_X1 U6282 ( .A1(n5561), .A2(n4871), .ZN(n5617) );
  NAND3_X1 U6283 ( .A1(n7715), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n4872) );
  INV_X1 U6284 ( .A(SI_1_), .ZN(n4873) );
  MUX2_X1 U6285 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5561), .Z(n4896) );
  XNOR2_X1 U6286 ( .A(n4897), .B(n4896), .ZN(n6292) );
  NAND2_X1 U6287 ( .A1(n4902), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4876) );
  NAND2_X1 U6288 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4874) );
  NAND2_X1 U6289 ( .A1(n5294), .A2(n6212), .ZN(n4875) );
  OAI211_X2 U6290 ( .C1(n4869), .C2(n6292), .A(n4876), .B(n4875), .ZN(n6884)
         );
  NAND2_X1 U6291 ( .A1(n4879), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4880) );
  NAND2_X1 U6292 ( .A1(n5443), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n4886) );
  INV_X1 U6293 ( .A(n4882), .ZN(n8091) );
  NAND2_X1 U6294 ( .A1(n4973), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4885) );
  NAND2_X1 U6295 ( .A1(n4954), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4884) );
  OR2_X4 U6296 ( .A1(n8442), .A2(n8399), .ZN(n8239) );
  NAND2_X1 U6297 ( .A1(n8465), .A2(n8239), .ZN(n4894) );
  NAND2_X1 U6298 ( .A1(n5443), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n4890) );
  NAND2_X1 U6299 ( .A1(n4973), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4889) );
  NAND2_X1 U6300 ( .A1(n4954), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n4888) );
  NAND2_X1 U6301 ( .A1(n4972), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n4887) );
  NAND2_X1 U6302 ( .A1(n7715), .A2(SI_0_), .ZN(n4891) );
  XNOR2_X1 U6303 ( .A(n4891), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8976) );
  MUX2_X1 U6304 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8976), .S(n6195), .Z(n9898) );
  NAND2_X1 U6305 ( .A1(n6889), .A2(n8239), .ZN(n6821) );
  INV_X1 U6306 ( .A(n9898), .ZN(n6947) );
  NAND2_X1 U6307 ( .A1(n5482), .A2(n6947), .ZN(n4892) );
  NAND2_X1 U6308 ( .A1(n6821), .A2(n4892), .ZN(n6617) );
  NAND2_X1 U6309 ( .A1(n6842), .A2(n4894), .ZN(n4895) );
  NAND2_X1 U6310 ( .A1(n4897), .A2(n4896), .ZN(n4900) );
  NAND2_X1 U6311 ( .A1(n4898), .A2(SI_1_), .ZN(n4899) );
  INV_X1 U6312 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6290) );
  INV_X1 U6313 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6295) );
  MUX2_X1 U6314 ( .A(n6290), .B(n6295), .S(n5561), .Z(n4921) );
  XNOR2_X1 U6315 ( .A(n4921), .B(SI_2_), .ZN(n4919) );
  XNOR2_X1 U6316 ( .A(n4920), .B(n4919), .ZN(n6294) );
  INV_X1 U6317 ( .A(n6294), .ZN(n4901) );
  NAND2_X1 U6318 ( .A1(n4940), .A2(n4901), .ZN(n4910) );
  NAND2_X1 U6319 ( .A1(n4902), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n4909) );
  NOR2_X1 U6320 ( .A1(n4903), .A2(n8964), .ZN(n4904) );
  NAND2_X1 U6321 ( .A1(n4904), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n4907) );
  INV_X1 U6322 ( .A(n4904), .ZN(n4906) );
  INV_X1 U6323 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4905) );
  NAND2_X1 U6324 ( .A1(n4906), .A2(n4905), .ZN(n4926) );
  AND2_X1 U6325 ( .A1(n4907), .A2(n4926), .ZN(n6240) );
  NAND2_X1 U6326 ( .A1(n5294), .A2(n6240), .ZN(n4908) );
  AND3_X2 U6327 ( .A1(n4910), .A2(n4909), .A3(n4908), .ZN(n9916) );
  XNOR2_X1 U6328 ( .A(n9916), .B(n5482), .ZN(n4915) );
  NAND2_X1 U6329 ( .A1(n5443), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n4914) );
  NAND2_X1 U6330 ( .A1(n4973), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4913) );
  NAND2_X1 U6331 ( .A1(n4954), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4912) );
  NAND2_X1 U6332 ( .A1(n8464), .A2(n8239), .ZN(n4916) );
  XNOR2_X1 U6333 ( .A(n4915), .B(n4916), .ZN(n6844) );
  INV_X1 U6334 ( .A(n4915), .ZN(n4917) );
  NAND2_X1 U6335 ( .A1(n4917), .A2(n4916), .ZN(n4918) );
  NAND2_X1 U6336 ( .A1(n4920), .A2(n4919), .ZN(n4924) );
  INV_X1 U6337 ( .A(n4921), .ZN(n4922) );
  NAND2_X1 U6338 ( .A1(n4922), .A2(SI_2_), .ZN(n4923) );
  MUX2_X1 U6339 ( .A(n8933), .B(n6297), .S(n5561), .Z(n4943) );
  XNOR2_X1 U6340 ( .A(n4943), .B(SI_3_), .ZN(n4941) );
  XNOR2_X1 U6341 ( .A(n4942), .B(n4941), .ZN(n6296) );
  INV_X1 U6342 ( .A(n6296), .ZN(n4925) );
  NAND2_X1 U6343 ( .A1(n4266), .A2(n4925), .ZN(n4930) );
  NAND2_X1 U6344 ( .A1(n5328), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n4929) );
  NAND2_X1 U6345 ( .A1(n4926), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4927) );
  XNOR2_X1 U6346 ( .A(n4927), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6253) );
  NAND2_X1 U6347 ( .A1(n5294), .A2(n6253), .ZN(n4928) );
  XNOR2_X1 U6348 ( .A(n6915), .B(n5482), .ZN(n4936) );
  INV_X1 U6349 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n4931) );
  NAND2_X1 U6350 ( .A1(n5443), .A2(n4931), .ZN(n4935) );
  NAND2_X1 U6351 ( .A1(n4973), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4934) );
  NAND2_X1 U6352 ( .A1(n6328), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4933) );
  NAND2_X1 U6353 ( .A1(n4972), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n4932) );
  NAND4_X1 U6354 ( .A1(n4935), .A2(n4934), .A3(n4933), .A4(n4932), .ZN(n8463)
         );
  AND2_X1 U6355 ( .A1(n8463), .A2(n8239), .ZN(n4937) );
  NAND2_X1 U6356 ( .A1(n4936), .A2(n4937), .ZN(n4959) );
  INV_X1 U6357 ( .A(n4936), .ZN(n6857) );
  INV_X1 U6358 ( .A(n4937), .ZN(n4938) );
  NAND2_X1 U6359 ( .A1(n6857), .A2(n4938), .ZN(n4939) );
  AND2_X1 U6360 ( .A1(n4959), .A2(n4939), .ZN(n6657) );
  INV_X1 U6361 ( .A(n4943), .ZN(n4944) );
  NAND2_X1 U6362 ( .A1(n4944), .A2(SI_3_), .ZN(n4945) );
  XNOR2_X1 U6363 ( .A(n4965), .B(SI_4_), .ZN(n4963) );
  INV_X1 U6364 ( .A(n6300), .ZN(n4946) );
  NAND2_X1 U6365 ( .A1(n8231), .A2(n4946), .ZN(n4953) );
  NAND2_X1 U6366 ( .A1(n5328), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n4952) );
  NAND2_X1 U6367 ( .A1(n4947), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4948) );
  MUX2_X1 U6368 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4948), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n4950) );
  AND2_X1 U6369 ( .A1(n4950), .A2(n4949), .ZN(n6228) );
  NAND2_X1 U6370 ( .A1(n5294), .A2(n6228), .ZN(n4951) );
  XNOR2_X1 U6371 ( .A(n9920), .B(n5482), .ZN(n7990) );
  NAND2_X1 U6372 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n4975) );
  OAI21_X1 U6373 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n4975), .ZN(n7018) );
  INV_X1 U6374 ( .A(n7018), .ZN(n6856) );
  NAND2_X1 U6375 ( .A1(n5443), .A2(n6856), .ZN(n4958) );
  NAND2_X1 U6376 ( .A1(n4973), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4957) );
  NAND2_X1 U6377 ( .A1(n6328), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4956) );
  NAND2_X1 U6378 ( .A1(n4972), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n4955) );
  NAND4_X1 U6379 ( .A1(n4958), .A2(n4957), .A3(n4956), .A4(n4955), .ZN(n8462)
         );
  NAND2_X1 U6380 ( .A1(n8462), .A2(n8239), .ZN(n4961) );
  XNOR2_X1 U6381 ( .A(n7990), .B(n4961), .ZN(n6858) );
  INV_X1 U6382 ( .A(n7990), .ZN(n4962) );
  INV_X1 U6383 ( .A(n4965), .ZN(n4966) );
  MUX2_X1 U6384 ( .A(n6305), .B(n6302), .S(n5561), .Z(n4987) );
  XNOR2_X1 U6385 ( .A(n4987), .B(SI_5_), .ZN(n4985) );
  XNOR2_X1 U6386 ( .A(n4986), .B(n4985), .ZN(n6304) );
  INV_X1 U6387 ( .A(n6304), .ZN(n4967) );
  NAND2_X1 U6388 ( .A1(n8231), .A2(n4967), .ZN(n4971) );
  NAND2_X1 U6389 ( .A1(n5328), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n4970) );
  NAND2_X1 U6390 ( .A1(n4949), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4968) );
  XNOR2_X1 U6391 ( .A(n4968), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6266) );
  NAND2_X1 U6392 ( .A1(n5294), .A2(n6266), .ZN(n4969) );
  XNOR2_X1 U6393 ( .A(n6995), .B(n5482), .ZN(n4981) );
  INV_X2 U6394 ( .A(n5000), .ZN(n6327) );
  NAND2_X1 U6395 ( .A1(n6327), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4979) );
  AND2_X1 U6396 ( .A1(n4975), .A2(n4974), .ZN(n4976) );
  NOR2_X1 U6397 ( .A1(n4989), .A2(n4976), .ZN(n6990) );
  NAND2_X1 U6398 ( .A1(n5532), .A2(n6990), .ZN(n4978) );
  NAND2_X1 U6399 ( .A1(n6328), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4977) );
  NAND4_X1 U6400 ( .A1(n4980), .A2(n4979), .A3(n4978), .A4(n4977), .ZN(n8461)
         );
  NAND2_X1 U6401 ( .A1(n8461), .A2(n8239), .ZN(n4982) );
  XNOR2_X1 U6402 ( .A(n4981), .B(n4982), .ZN(n7991) );
  INV_X1 U6403 ( .A(n4981), .ZN(n6832) );
  NAND2_X1 U6404 ( .A1(n6832), .A2(n4982), .ZN(n4983) );
  NAND2_X1 U6405 ( .A1(n7997), .A2(n4983), .ZN(n4995) );
  INV_X2 U6406 ( .A(n5482), .ZN(n5459) );
  NOR2_X1 U6407 ( .A1(n4949), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5013) );
  OR2_X1 U6408 ( .A1(n5013), .A2(n8964), .ZN(n4984) );
  XNOR2_X1 U6409 ( .A(n4984), .B(n5012), .ZN(n6306) );
  INV_X1 U6410 ( .A(n4987), .ZN(n4988) );
  NAND2_X1 U6411 ( .A1(n4988), .A2(SI_5_), .ZN(n5025) );
  MUX2_X1 U6412 ( .A(n6307), .B(n6309), .S(n5561), .Z(n5009) );
  XNOR2_X1 U6413 ( .A(n5009), .B(SI_6_), .ZN(n5031) );
  XNOR2_X1 U6414 ( .A(n5459), .B(n7130), .ZN(n4996) );
  NAND2_X1 U6415 ( .A1(n6329), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n4994) );
  NAND2_X1 U6416 ( .A1(n6327), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4993) );
  NAND2_X1 U6417 ( .A1(n4989), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5002) );
  OR2_X1 U6418 ( .A1(n4989), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n4990) );
  AND2_X1 U6419 ( .A1(n5002), .A2(n4990), .ZN(n7127) );
  NAND2_X1 U6420 ( .A1(n5532), .A2(n7127), .ZN(n4992) );
  NAND2_X1 U6421 ( .A1(n6328), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4991) );
  OR2_X1 U6422 ( .A1(n6751), .A2(n5481), .ZN(n4998) );
  XNOR2_X1 U6423 ( .A(n4996), .B(n4998), .ZN(n6831) );
  INV_X1 U6424 ( .A(n4996), .ZN(n4997) );
  NAND2_X1 U6425 ( .A1(n4998), .A2(n4997), .ZN(n4999) );
  NAND2_X1 U6426 ( .A1(n6329), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5007) );
  NAND2_X1 U6427 ( .A1(n6327), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5006) );
  NAND2_X1 U6428 ( .A1(n5002), .A2(n5001), .ZN(n5003) );
  AND2_X1 U6429 ( .A1(n5044), .A2(n5003), .ZN(n6894) );
  NAND2_X1 U6430 ( .A1(n5443), .A2(n6894), .ZN(n5005) );
  NAND2_X1 U6431 ( .A1(n6328), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5004) );
  NOR2_X1 U6432 ( .A1(n6825), .A2(n5481), .ZN(n5017) );
  NAND2_X1 U6433 ( .A1(n5008), .A2(n5031), .ZN(n5011) );
  INV_X1 U6434 ( .A(n5009), .ZN(n5010) );
  NAND2_X1 U6435 ( .A1(n5010), .A2(SI_6_), .ZN(n5024) );
  XNOR2_X1 U6436 ( .A(n5023), .B(SI_7_), .ZN(n5029) );
  NAND2_X1 U6437 ( .A1(n6315), .A2(n8231), .ZN(n5016) );
  NAND2_X1 U6438 ( .A1(n5013), .A2(n5012), .ZN(n5039) );
  NAND2_X1 U6439 ( .A1(n5039), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5014) );
  XNOR2_X1 U6440 ( .A(n5014), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6631) );
  AOI22_X1 U6441 ( .A1(n5328), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5294), .B2(
        n6631), .ZN(n5015) );
  XNOR2_X1 U6442 ( .A(n6767), .B(n5459), .ZN(n9849) );
  NAND2_X1 U6443 ( .A1(n5017), .A2(n9849), .ZN(n5022) );
  INV_X1 U6444 ( .A(n9849), .ZN(n5019) );
  INV_X1 U6445 ( .A(n5017), .ZN(n5018) );
  NAND2_X1 U6446 ( .A1(n5019), .A2(n5018), .ZN(n5020) );
  NAND2_X1 U6447 ( .A1(n5022), .A2(n5020), .ZN(n6762) );
  NAND2_X1 U6448 ( .A1(n6761), .A2(n5022), .ZN(n5054) );
  NAND2_X1 U6449 ( .A1(n5023), .A2(SI_7_), .ZN(n5028) );
  AND2_X1 U6450 ( .A1(n5025), .A2(n5030), .ZN(n5026) );
  INV_X1 U6451 ( .A(n5030), .ZN(n5032) );
  MUX2_X1 U6452 ( .A(n6319), .B(n6321), .S(n5561), .Z(n5036) );
  INV_X1 U6453 ( .A(SI_8_), .ZN(n5035) );
  NAND2_X1 U6454 ( .A1(n5036), .A2(n5035), .ZN(n5057) );
  INV_X1 U6455 ( .A(n5036), .ZN(n5037) );
  NAND2_X1 U6456 ( .A1(n5037), .A2(SI_8_), .ZN(n5038) );
  NAND2_X1 U6457 ( .A1(n5057), .A2(n5038), .ZN(n5055) );
  XNOR2_X1 U6458 ( .A(n5056), .B(n5055), .ZN(n6318) );
  NAND2_X1 U6459 ( .A1(n6318), .A2(n8231), .ZN(n5042) );
  NAND2_X1 U6460 ( .A1(n5063), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5040) );
  XNOR2_X1 U6461 ( .A(n5040), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6645) );
  AOI22_X1 U6462 ( .A1(n5328), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5294), .B2(
        n6645), .ZN(n5041) );
  NAND2_X1 U6463 ( .A1(n5042), .A2(n5041), .ZN(n9853) );
  XNOR2_X1 U6464 ( .A(n9853), .B(n5459), .ZN(n5050) );
  NAND2_X1 U6465 ( .A1(n5044), .A2(n5043), .ZN(n5045) );
  NAND2_X1 U6466 ( .A1(n5067), .A2(n5045), .ZN(n9859) );
  INV_X1 U6467 ( .A(n9859), .ZN(n6902) );
  NAND2_X1 U6468 ( .A1(n5532), .A2(n6902), .ZN(n5049) );
  NAND2_X1 U6469 ( .A1(n6327), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5048) );
  NAND2_X1 U6470 ( .A1(n4954), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5047) );
  NAND2_X1 U6471 ( .A1(n6329), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5046) );
  NOR2_X1 U6472 ( .A1(n6954), .A2(n5481), .ZN(n5051) );
  NAND2_X1 U6473 ( .A1(n5050), .A2(n5051), .ZN(n5073) );
  INV_X1 U6474 ( .A(n5050), .ZN(n8183) );
  INV_X1 U6475 ( .A(n5051), .ZN(n5052) );
  NAND2_X1 U6476 ( .A1(n8183), .A2(n5052), .ZN(n5053) );
  AND2_X1 U6477 ( .A1(n5073), .A2(n5053), .ZN(n9846) );
  NAND2_X1 U6478 ( .A1(n5054), .A2(n9846), .ZN(n9855) );
  INV_X1 U6479 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5058) );
  MUX2_X1 U6480 ( .A(n5058), .B(n8890), .S(n5561), .Z(n5060) );
  INV_X1 U6481 ( .A(SI_9_), .ZN(n5059) );
  NAND2_X1 U6482 ( .A1(n5060), .A2(n5059), .ZN(n5080) );
  INV_X1 U6483 ( .A(n5060), .ZN(n5061) );
  NAND2_X1 U6484 ( .A1(n5061), .A2(SI_9_), .ZN(n5062) );
  XNOR2_X1 U6485 ( .A(n5079), .B(n4838), .ZN(n6322) );
  NAND2_X1 U6486 ( .A1(n6322), .A2(n8231), .ZN(n5065) );
  NAND2_X1 U6487 ( .A1(n5129), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5087) );
  XNOR2_X1 U6488 ( .A(n5087), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6666) );
  AOI22_X1 U6489 ( .A1(n5328), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5294), .B2(
        n6666), .ZN(n5064) );
  NAND2_X1 U6490 ( .A1(n5065), .A2(n5064), .ZN(n8182) );
  XNOR2_X1 U6491 ( .A(n8182), .B(n5482), .ZN(n5077) );
  NAND2_X1 U6492 ( .A1(n6329), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5072) );
  NAND2_X1 U6493 ( .A1(n6327), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5071) );
  AND2_X1 U6494 ( .A1(n5067), .A2(n5066), .ZN(n5068) );
  NOR2_X1 U6495 ( .A1(n5110), .A2(n5068), .ZN(n8177) );
  NAND2_X1 U6496 ( .A1(n5532), .A2(n8177), .ZN(n5070) );
  NAND2_X1 U6497 ( .A1(n6328), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5069) );
  NOR2_X1 U6498 ( .A1(n9832), .A2(n5481), .ZN(n5075) );
  XNOR2_X1 U6499 ( .A(n5077), .B(n5075), .ZN(n8184) );
  AND2_X1 U6500 ( .A1(n8184), .A2(n5073), .ZN(n5074) );
  INV_X1 U6501 ( .A(n5075), .ZN(n5076) );
  NAND2_X1 U6502 ( .A1(n5077), .A2(n5076), .ZN(n5078) );
  MUX2_X1 U6503 ( .A(n5082), .B(n6336), .S(n5561), .Z(n5084) );
  INV_X1 U6504 ( .A(SI_10_), .ZN(n5083) );
  NAND2_X1 U6505 ( .A1(n5084), .A2(n5083), .ZN(n5103) );
  INV_X1 U6506 ( .A(n5084), .ZN(n5085) );
  NAND2_X1 U6507 ( .A1(n5085), .A2(SI_10_), .ZN(n5086) );
  XNOR2_X1 U6508 ( .A(n5102), .B(n4839), .ZN(n6325) );
  NAND2_X1 U6509 ( .A1(n6325), .A2(n4266), .ZN(n5090) );
  INV_X1 U6510 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5131) );
  NAND2_X1 U6511 ( .A1(n5087), .A2(n5131), .ZN(n5088) );
  NAND2_X1 U6512 ( .A1(n5088), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5104) );
  XNOR2_X1 U6513 ( .A(n5104), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6694) );
  AOI22_X1 U6514 ( .A1(n5328), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5294), .B2(
        n6694), .ZN(n5089) );
  NAND2_X1 U6515 ( .A1(n5090), .A2(n5089), .ZN(n9840) );
  XNOR2_X1 U6516 ( .A(n9840), .B(n5459), .ZN(n5096) );
  XNOR2_X1 U6517 ( .A(n5110), .B(P2_REG3_REG_10__SCAN_IN), .ZN(n9842) );
  INV_X1 U6518 ( .A(n9842), .ZN(n5091) );
  NAND2_X1 U6519 ( .A1(n5443), .A2(n5091), .ZN(n5095) );
  NAND2_X1 U6520 ( .A1(n6327), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5094) );
  NAND2_X1 U6521 ( .A1(n4954), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5093) );
  NAND2_X1 U6522 ( .A1(n6329), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5092) );
  NOR2_X1 U6523 ( .A1(n8180), .A2(n5481), .ZN(n5097) );
  NAND2_X1 U6524 ( .A1(n5096), .A2(n5097), .ZN(n5101) );
  INV_X1 U6525 ( .A(n5096), .ZN(n7161) );
  INV_X1 U6526 ( .A(n5097), .ZN(n5098) );
  NAND2_X1 U6527 ( .A1(n7161), .A2(n5098), .ZN(n5099) );
  NAND2_X1 U6528 ( .A1(n5101), .A2(n5099), .ZN(n9837) );
  INV_X1 U6529 ( .A(n9837), .ZN(n5100) );
  MUX2_X1 U6530 ( .A(n6338), .B(n6339), .S(n5561), .Z(n5121) );
  XNOR2_X1 U6531 ( .A(n5121), .B(SI_11_), .ZN(n5120) );
  XNOR2_X1 U6532 ( .A(n5124), .B(n5120), .ZN(n6337) );
  NAND2_X1 U6533 ( .A1(n6337), .A2(n4266), .ZN(n5108) );
  INV_X1 U6534 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5132) );
  NAND2_X1 U6535 ( .A1(n5104), .A2(n5132), .ZN(n5105) );
  NAND2_X1 U6536 ( .A1(n5105), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5106) );
  XNOR2_X1 U6537 ( .A(n5106), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6791) );
  AOI22_X1 U6538 ( .A1(n5328), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5294), .B2(
        n6791), .ZN(n5107) );
  NAND2_X1 U6539 ( .A1(n5108), .A2(n5107), .ZN(n7265) );
  XNOR2_X1 U6540 ( .A(n7265), .B(n5459), .ZN(n5116) );
  NAND2_X1 U6541 ( .A1(n6329), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5115) );
  NAND2_X1 U6542 ( .A1(n6327), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5114) );
  AND2_X1 U6543 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n5109) );
  AOI21_X1 U6544 ( .B1(n5110), .B2(P2_REG3_REG_10__SCAN_IN), .A(
        P2_REG3_REG_11__SCAN_IN), .ZN(n5111) );
  OR2_X1 U6545 ( .A1(n5140), .A2(n5111), .ZN(n7165) );
  INV_X1 U6546 ( .A(n7165), .ZN(n7266) );
  NAND2_X1 U6547 ( .A1(n5532), .A2(n7266), .ZN(n5113) );
  NAND2_X1 U6548 ( .A1(n6328), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5112) );
  NOR2_X1 U6549 ( .A1(n7345), .A2(n5481), .ZN(n5117) );
  NAND2_X1 U6550 ( .A1(n5116), .A2(n5117), .ZN(n5146) );
  INV_X1 U6551 ( .A(n5116), .ZN(n7346) );
  INV_X1 U6552 ( .A(n5117), .ZN(n5118) );
  NAND2_X1 U6553 ( .A1(n7346), .A2(n5118), .ZN(n5119) );
  AND2_X1 U6554 ( .A1(n5146), .A2(n5119), .ZN(n7159) );
  INV_X1 U6555 ( .A(n5120), .ZN(n5123) );
  INV_X1 U6556 ( .A(n5121), .ZN(n5122) );
  MUX2_X1 U6557 ( .A(n6421), .B(n8934), .S(n5561), .Z(n5126) );
  INV_X1 U6558 ( .A(n5126), .ZN(n5127) );
  NAND2_X1 U6559 ( .A1(n5127), .A2(SI_12_), .ZN(n5128) );
  NAND2_X1 U6560 ( .A1(n5154), .A2(n5128), .ZN(n5152) );
  XNOR2_X1 U6561 ( .A(n5153), .B(n5152), .ZN(n6420) );
  NAND2_X1 U6562 ( .A1(n6420), .A2(n8231), .ZN(n5139) );
  INV_X1 U6563 ( .A(n5129), .ZN(n5134) );
  INV_X1 U6564 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5130) );
  AND3_X1 U6565 ( .A1(n5132), .A2(n5131), .A3(n5130), .ZN(n5133) );
  AOI21_X1 U6566 ( .B1(n5134), .B2(n5133), .A(n8964), .ZN(n5135) );
  MUX2_X1 U6567 ( .A(n8964), .B(n5135), .S(P2_IR_REG_12__SCAN_IN), .Z(n5137)
         );
  OR2_X1 U6568 ( .A1(n5137), .A2(n5136), .ZN(n6974) );
  AOI22_X1 U6569 ( .A1(n5328), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5294), .B2(
        n6968), .ZN(n5138) );
  XNOR2_X1 U6570 ( .A(n7361), .B(n5482), .ZN(n5150) );
  NAND2_X1 U6571 ( .A1(n6329), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5145) );
  NAND2_X1 U6572 ( .A1(n6327), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5144) );
  NOR2_X1 U6573 ( .A1(n5140), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5141) );
  NAND2_X1 U6574 ( .A1(n5532), .A2(n4841), .ZN(n5143) );
  NAND2_X1 U6575 ( .A1(n6328), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5142) );
  NOR2_X1 U6576 ( .A1(n7328), .A2(n5481), .ZN(n5148) );
  XNOR2_X1 U6577 ( .A(n5150), .B(n5148), .ZN(n7357) );
  AND2_X1 U6578 ( .A1(n7357), .A2(n5146), .ZN(n5147) );
  INV_X1 U6579 ( .A(n5148), .ZN(n5149) );
  NAND2_X1 U6580 ( .A1(n5150), .A2(n5149), .ZN(n5151) );
  MUX2_X1 U6581 ( .A(n5155), .B(n6510), .S(n5561), .Z(n5157) );
  INV_X1 U6582 ( .A(SI_13_), .ZN(n5156) );
  INV_X1 U6583 ( .A(n5157), .ZN(n5158) );
  NAND2_X1 U6584 ( .A1(n5158), .A2(SI_13_), .ZN(n5159) );
  XNOR2_X1 U6585 ( .A(n5175), .B(n4840), .ZN(n6507) );
  NAND2_X1 U6586 ( .A1(n6507), .A2(n8231), .ZN(n5162) );
  OR2_X1 U6587 ( .A1(n5136), .A2(n8964), .ZN(n5160) );
  XNOR2_X1 U6588 ( .A(n5160), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6985) );
  AOI22_X1 U6589 ( .A1(n5328), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5294), .B2(
        n6985), .ZN(n5161) );
  XNOR2_X1 U6590 ( .A(n7438), .B(n5459), .ZN(n5169) );
  NAND2_X1 U6591 ( .A1(n6329), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5168) );
  NAND2_X1 U6592 ( .A1(n6327), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5167) );
  OR2_X1 U6593 ( .A1(n5163), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5164) );
  AND2_X1 U6594 ( .A1(n5164), .A2(n5182), .ZN(n7375) );
  NAND2_X1 U6595 ( .A1(n5532), .A2(n7375), .ZN(n5166) );
  NAND2_X1 U6596 ( .A1(n6328), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5165) );
  NOR2_X1 U6597 ( .A1(n7434), .A2(n5481), .ZN(n5170) );
  NAND2_X1 U6598 ( .A1(n5169), .A2(n5170), .ZN(n9470) );
  INV_X1 U6599 ( .A(n5169), .ZN(n5172) );
  INV_X1 U6600 ( .A(n5170), .ZN(n5171) );
  NAND2_X1 U6601 ( .A1(n5172), .A2(n5171), .ZN(n5173) );
  NAND2_X1 U6602 ( .A1(n9470), .A2(n5173), .ZN(n7325) );
  MUX2_X1 U6603 ( .A(n8891), .B(n8935), .S(n5561), .Z(n5196) );
  XNOR2_X1 U6604 ( .A(n5196), .B(SI_14_), .ZN(n5193) );
  XNOR2_X1 U6605 ( .A(n5195), .B(n5193), .ZN(n6511) );
  NAND2_X1 U6606 ( .A1(n6511), .A2(n8231), .ZN(n5181) );
  OR2_X1 U6607 ( .A1(n5178), .A2(n8964), .ZN(n5179) );
  XNOR2_X1 U6608 ( .A(n5179), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7219) );
  AOI22_X1 U6609 ( .A1(n5328), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5294), .B2(
        n7219), .ZN(n5180) );
  XNOR2_X1 U6610 ( .A(n9476), .B(n5459), .ZN(n5190) );
  NAND2_X1 U6611 ( .A1(n5182), .A2(n8820), .ZN(n5183) );
  NAND2_X1 U6612 ( .A1(n5213), .A2(n5183), .ZN(n9482) );
  INV_X1 U6613 ( .A(n9482), .ZN(n5184) );
  NAND2_X1 U6614 ( .A1(n5443), .A2(n5184), .ZN(n5188) );
  NAND2_X1 U6615 ( .A1(n6327), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5187) );
  NAND2_X1 U6616 ( .A1(n6328), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U6617 ( .A1(n6329), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5185) );
  NAND4_X1 U6618 ( .A1(n5188), .A2(n5187), .A3(n5186), .A4(n5185), .ZN(n8454)
         );
  NAND2_X1 U6619 ( .A1(n8454), .A2(n8239), .ZN(n5191) );
  XNOR2_X1 U6620 ( .A(n5190), .B(n5191), .ZN(n9473) );
  AND2_X1 U6621 ( .A1(n9473), .A2(n9470), .ZN(n5189) );
  INV_X1 U6622 ( .A(n5190), .ZN(n5192) );
  NAND2_X1 U6623 ( .A1(n5192), .A2(n5191), .ZN(n5209) );
  NAND2_X1 U6624 ( .A1(n9472), .A2(n5209), .ZN(n5207) );
  INV_X1 U6625 ( .A(n5193), .ZN(n5194) );
  INV_X1 U6626 ( .A(n5196), .ZN(n5197) );
  NAND2_X1 U6627 ( .A1(n5197), .A2(SI_14_), .ZN(n5198) );
  MUX2_X1 U6628 ( .A(n6544), .B(n5199), .S(n5561), .Z(n5200) );
  NAND2_X1 U6629 ( .A1(n5200), .A2(n8815), .ZN(n5220) );
  INV_X1 U6630 ( .A(n5200), .ZN(n5201) );
  NAND2_X1 U6631 ( .A1(n5201), .A2(SI_15_), .ZN(n5202) );
  NAND2_X1 U6632 ( .A1(n5220), .A2(n5202), .ZN(n5221) );
  XNOR2_X1 U6633 ( .A(n5222), .B(n5221), .ZN(n6539) );
  NAND2_X1 U6634 ( .A1(n6539), .A2(n4266), .ZN(n5206) );
  NAND2_X1 U6635 ( .A1(n5203), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5204) );
  XNOR2_X1 U6636 ( .A(n5204), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7509) );
  AOI22_X1 U6637 ( .A1(n5328), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5294), .B2(
        n7509), .ZN(n5205) );
  NAND2_X2 U6638 ( .A1(n5206), .A2(n5205), .ZN(n7552) );
  XNOR2_X1 U6639 ( .A(n7552), .B(n5482), .ZN(n5208) );
  NAND2_X2 U6640 ( .A1(n5207), .A2(n5208), .ZN(n7544) );
  INV_X1 U6641 ( .A(n5208), .ZN(n5210) );
  AND2_X1 U6642 ( .A1(n5210), .A2(n5209), .ZN(n5211) );
  INV_X1 U6643 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7548) );
  NAND2_X1 U6644 ( .A1(n5213), .A2(n7548), .ZN(n5214) );
  AND2_X1 U6645 ( .A1(n5232), .A2(n5214), .ZN(n7547) );
  NAND2_X1 U6646 ( .A1(n5443), .A2(n7547), .ZN(n5218) );
  NAND2_X1 U6647 ( .A1(n6327), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5217) );
  NAND2_X1 U6648 ( .A1(n6328), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5216) );
  NAND2_X1 U6649 ( .A1(n6329), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5215) );
  OR2_X1 U6650 ( .A1(n7602), .A2(n5481), .ZN(n7546) );
  NAND2_X1 U6651 ( .A1(n7543), .A2(n7546), .ZN(n5219) );
  MUX2_X1 U6652 ( .A(n8831), .B(n5223), .S(n5561), .Z(n5225) );
  INV_X1 U6653 ( .A(SI_16_), .ZN(n5224) );
  NAND2_X1 U6654 ( .A1(n5225), .A2(n5224), .ZN(n5244) );
  INV_X1 U6655 ( .A(n5225), .ZN(n5226) );
  NAND2_X1 U6656 ( .A1(n5226), .A2(SI_16_), .ZN(n5227) );
  XNOR2_X1 U6657 ( .A(n5243), .B(n5242), .ZN(n6541) );
  NAND2_X1 U6658 ( .A1(n6541), .A2(n8231), .ZN(n5231) );
  NAND2_X1 U6659 ( .A1(n5228), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5229) );
  XNOR2_X1 U6660 ( .A(n5229), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8477) );
  AOI22_X1 U6661 ( .A1(n5328), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5294), .B2(
        n8477), .ZN(n5230) );
  XNOR2_X1 U6662 ( .A(n8795), .B(n5482), .ZN(n5240) );
  NAND2_X1 U6663 ( .A1(n6329), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5237) );
  NAND2_X1 U6664 ( .A1(n6327), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5236) );
  NAND2_X1 U6665 ( .A1(n5232), .A2(n8840), .ZN(n5233) );
  AND2_X1 U6666 ( .A1(n5253), .A2(n5233), .ZN(n7609) );
  NAND2_X1 U6667 ( .A1(n5532), .A2(n7609), .ZN(n5235) );
  NAND2_X1 U6668 ( .A1(n6328), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5234) );
  NOR2_X1 U6669 ( .A1(n8154), .A2(n5481), .ZN(n5238) );
  XNOR2_X1 U6670 ( .A(n5240), .B(n5238), .ZN(n7492) );
  INV_X1 U6671 ( .A(n5238), .ZN(n5239) );
  NAND2_X1 U6672 ( .A1(n5240), .A2(n5239), .ZN(n5241) );
  INV_X1 U6673 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n5245) );
  MUX2_X1 U6674 ( .A(n5245), .B(n6569), .S(n5561), .Z(n5266) );
  XNOR2_X1 U6675 ( .A(n5266), .B(SI_17_), .ZN(n5265) );
  XNOR2_X1 U6676 ( .A(n5269), .B(n5265), .ZN(n6566) );
  NAND2_X1 U6677 ( .A1(n6566), .A2(n4266), .ZN(n5250) );
  INV_X1 U6678 ( .A(n5246), .ZN(n5247) );
  NAND2_X1 U6679 ( .A1(n5247), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5248) );
  XNOR2_X1 U6680 ( .A(n5248), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9875) );
  AOI22_X1 U6681 ( .A1(n5328), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5294), .B2(
        n9875), .ZN(n5249) );
  XNOR2_X1 U6682 ( .A(n8787), .B(n5459), .ZN(n5259) );
  NAND2_X1 U6683 ( .A1(n6329), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5258) );
  INV_X1 U6684 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5252) );
  NAND2_X1 U6685 ( .A1(n5253), .A2(n5252), .ZN(n5254) );
  AND2_X1 U6686 ( .A1(n5274), .A2(n5254), .ZN(n8157) );
  NAND2_X1 U6687 ( .A1(n5532), .A2(n8157), .ZN(n5257) );
  NAND2_X1 U6688 ( .A1(n6327), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5256) );
  NAND2_X1 U6689 ( .A1(n6328), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5255) );
  NOR2_X1 U6690 ( .A1(n8203), .A2(n5481), .ZN(n5260) );
  NAND2_X1 U6691 ( .A1(n5259), .A2(n5260), .ZN(n5264) );
  INV_X1 U6692 ( .A(n5259), .ZN(n8204) );
  INV_X1 U6693 ( .A(n5260), .ZN(n5261) );
  NAND2_X1 U6694 ( .A1(n8204), .A2(n5261), .ZN(n5262) );
  NAND2_X1 U6695 ( .A1(n5264), .A2(n5262), .ZN(n8151) );
  INV_X1 U6696 ( .A(n8151), .ZN(n5263) );
  INV_X1 U6697 ( .A(n5266), .ZN(n5267) );
  NAND2_X1 U6698 ( .A1(n5267), .A2(SI_17_), .ZN(n5268) );
  MUX2_X1 U6699 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5561), .Z(n5288) );
  XNOR2_X1 U6700 ( .A(n5288), .B(SI_18_), .ZN(n5285) );
  XNOR2_X1 U6701 ( .A(n5287), .B(n5285), .ZN(n6674) );
  NAND2_X1 U6702 ( .A1(n6674), .A2(n8231), .ZN(n5272) );
  XNOR2_X1 U6703 ( .A(n5270), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8480) );
  AOI22_X1 U6704 ( .A1(n5328), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5294), .B2(
        n8480), .ZN(n5271) );
  XNOR2_X1 U6705 ( .A(n8783), .B(n5459), .ZN(n8112) );
  INV_X1 U6706 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8208) );
  NAND2_X1 U6707 ( .A1(n5274), .A2(n8208), .ZN(n5275) );
  NAND2_X1 U6708 ( .A1(n5297), .A2(n5275), .ZN(n8207) );
  OR2_X1 U6709 ( .A1(n8207), .A2(n5463), .ZN(n5279) );
  NAND2_X1 U6710 ( .A1(n6329), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U6711 ( .A1(n6327), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5277) );
  NAND2_X1 U6712 ( .A1(n4954), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5276) );
  NOR2_X1 U6713 ( .A1(n8155), .A2(n5481), .ZN(n5280) );
  NAND2_X1 U6714 ( .A1(n8112), .A2(n5280), .ZN(n5301) );
  INV_X1 U6715 ( .A(n8112), .ZN(n5282) );
  INV_X1 U6716 ( .A(n5280), .ZN(n5281) );
  NAND2_X1 U6717 ( .A1(n5282), .A2(n5281), .ZN(n5283) );
  AND2_X1 U6718 ( .A1(n5301), .A2(n5283), .ZN(n8199) );
  NAND2_X1 U6719 ( .A1(n5288), .A2(SI_18_), .ZN(n5289) );
  MUX2_X1 U6720 ( .A(n6808), .B(n6810), .S(n5561), .Z(n5291) );
  INV_X1 U6721 ( .A(SI_19_), .ZN(n8916) );
  NAND2_X1 U6722 ( .A1(n5291), .A2(n8916), .ZN(n5309) );
  INV_X1 U6723 ( .A(n5291), .ZN(n5292) );
  NAND2_X1 U6724 ( .A1(n5292), .A2(SI_19_), .ZN(n5293) );
  NAND2_X1 U6725 ( .A1(n5309), .A2(n5293), .ZN(n5307) );
  XNOR2_X1 U6726 ( .A(n5308), .B(n5307), .ZN(n6807) );
  NAND2_X1 U6727 ( .A1(n6807), .A2(n8231), .ZN(n5296) );
  AOI22_X1 U6728 ( .A1(n5328), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8569), .B2(
        n5294), .ZN(n5295) );
  XNOR2_X1 U6729 ( .A(n8778), .B(n5459), .ZN(n5303) );
  INV_X1 U6730 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8681) );
  INV_X1 U6731 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8117) );
  NAND2_X1 U6732 ( .A1(n5297), .A2(n8117), .ZN(n5298) );
  NAND2_X1 U6733 ( .A1(n5316), .A2(n5298), .ZN(n8680) );
  OR2_X1 U6734 ( .A1(n8680), .A2(n5463), .ZN(n5300) );
  AOI22_X1 U6735 ( .A1(n6329), .A2(P2_REG0_REG_19__SCAN_IN), .B1(n6327), .B2(
        P2_REG1_REG_19__SCAN_IN), .ZN(n5299) );
  OAI211_X1 U6736 ( .C1(n5530), .C2(n8681), .A(n5300), .B(n5299), .ZN(n8657)
         );
  NAND2_X1 U6737 ( .A1(n8657), .A2(n8239), .ZN(n5304) );
  XNOR2_X1 U6738 ( .A(n5303), .B(n5304), .ZN(n8114) );
  AND2_X1 U6739 ( .A1(n8114), .A2(n5301), .ZN(n5302) );
  NAND2_X1 U6740 ( .A1(n8111), .A2(n5302), .ZN(n8122) );
  INV_X1 U6741 ( .A(n5303), .ZN(n5305) );
  NAND2_X1 U6742 ( .A1(n5305), .A2(n5304), .ZN(n5306) );
  NAND2_X1 U6743 ( .A1(n8122), .A2(n5306), .ZN(n6171) );
  MUX2_X1 U6744 ( .A(n7087), .B(n7703), .S(n5561), .Z(n5311) );
  INV_X1 U6745 ( .A(SI_20_), .ZN(n5310) );
  NAND2_X1 U6746 ( .A1(n5311), .A2(n5310), .ZN(n5327) );
  INV_X1 U6747 ( .A(n5311), .ZN(n5312) );
  NAND2_X1 U6748 ( .A1(n5312), .A2(SI_20_), .ZN(n5313) );
  XNOR2_X1 U6749 ( .A(n5326), .B(n5325), .ZN(n7086) );
  NAND2_X1 U6750 ( .A1(n7086), .A2(n4266), .ZN(n5315) );
  NAND2_X1 U6751 ( .A1(n5328), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5314) );
  XNOR2_X1 U6752 ( .A(n8771), .B(n5459), .ZN(n5320) );
  INV_X1 U6753 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n6174) );
  NAND2_X1 U6754 ( .A1(n5316), .A2(n6174), .ZN(n5317) );
  NAND2_X1 U6755 ( .A1(n5333), .A2(n5317), .ZN(n8663) );
  AOI22_X1 U6756 ( .A1(n6329), .A2(P2_REG0_REG_20__SCAN_IN), .B1(n6327), .B2(
        P2_REG1_REG_20__SCAN_IN), .ZN(n5319) );
  NAND2_X1 U6757 ( .A1(n6328), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5318) );
  OAI211_X1 U6758 ( .C1(n8663), .C2(n5463), .A(n5319), .B(n5318), .ZN(n8647)
         );
  AND2_X1 U6759 ( .A1(n8647), .A2(n8239), .ZN(n5321) );
  NAND2_X1 U6760 ( .A1(n5320), .A2(n5321), .ZN(n5324) );
  INV_X1 U6761 ( .A(n5320), .ZN(n8127) );
  INV_X1 U6762 ( .A(n5321), .ZN(n5322) );
  NAND2_X1 U6763 ( .A1(n8127), .A2(n5322), .ZN(n5323) );
  NAND2_X1 U6764 ( .A1(n5324), .A2(n5323), .ZN(n6172) );
  MUX2_X1 U6765 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n5561), .Z(n5347) );
  XNOR2_X1 U6766 ( .A(n5347), .B(n8906), .ZN(n5346) );
  XNOR2_X1 U6767 ( .A(n5345), .B(n5346), .ZN(n7084) );
  NAND2_X1 U6768 ( .A1(n7084), .A2(n4266), .ZN(n5330) );
  NAND2_X1 U6769 ( .A1(n5328), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5329) );
  XNOR2_X1 U6770 ( .A(n8764), .B(n5459), .ZN(n5343) );
  INV_X1 U6771 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5332) );
  NAND2_X1 U6772 ( .A1(n5333), .A2(n5332), .ZN(n5334) );
  AND2_X1 U6773 ( .A1(n5358), .A2(n5334), .ZN(n8642) );
  NAND2_X1 U6774 ( .A1(n8642), .A2(n5443), .ZN(n5340) );
  INV_X1 U6775 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n5337) );
  NAND2_X1 U6776 ( .A1(n6329), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5336) );
  NAND2_X1 U6777 ( .A1(n6327), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5335) );
  OAI211_X1 U6778 ( .C1(n5337), .C2(n5530), .A(n5336), .B(n5335), .ZN(n5338)
         );
  INV_X1 U6779 ( .A(n5338), .ZN(n5339) );
  NAND2_X1 U6780 ( .A1(n5340), .A2(n5339), .ZN(n8655) );
  NAND2_X1 U6781 ( .A1(n8655), .A2(n8239), .ZN(n5341) );
  XNOR2_X1 U6782 ( .A(n5343), .B(n5341), .ZN(n8123) );
  INV_X1 U6783 ( .A(n5341), .ZN(n5342) );
  NAND2_X1 U6784 ( .A1(n5343), .A2(n5342), .ZN(n5344) );
  NAND2_X1 U6785 ( .A1(n8128), .A2(n5344), .ZN(n5368) );
  NAND2_X1 U6786 ( .A1(n5347), .A2(SI_21_), .ZN(n5348) );
  INV_X1 U6787 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7227) );
  MUX2_X1 U6788 ( .A(n7227), .B(n8948), .S(n5561), .Z(n5351) );
  INV_X1 U6789 ( .A(SI_22_), .ZN(n5350) );
  NAND2_X1 U6790 ( .A1(n5351), .A2(n5350), .ZN(n5372) );
  INV_X1 U6791 ( .A(n5351), .ZN(n5352) );
  NAND2_X1 U6792 ( .A1(n5352), .A2(SI_22_), .ZN(n5353) );
  NAND2_X1 U6793 ( .A1(n5372), .A2(n5353), .ZN(n5370) );
  XNOR2_X1 U6794 ( .A(n5371), .B(n5370), .ZN(n7226) );
  NAND2_X1 U6795 ( .A1(n7226), .A2(n8231), .ZN(n5355) );
  NAND2_X1 U6796 ( .A1(n5328), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5354) );
  XNOR2_X1 U6797 ( .A(n8759), .B(n5482), .ZN(n5366) );
  XNOR2_X1 U6798 ( .A(n5368), .B(n5366), .ZN(n8190) );
  INV_X1 U6799 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n5357) );
  NAND2_X1 U6800 ( .A1(n5358), .A2(n5357), .ZN(n5359) );
  NAND2_X1 U6801 ( .A1(n5400), .A2(n5359), .ZN(n8193) );
  OR2_X1 U6802 ( .A1(n8193), .A2(n5463), .ZN(n5365) );
  INV_X1 U6803 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U6804 ( .A1(n6329), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6805 ( .A1(n6327), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5360) );
  OAI211_X1 U6806 ( .C1(n5362), .C2(n5530), .A(n5361), .B(n5360), .ZN(n5363)
         );
  INV_X1 U6807 ( .A(n5363), .ZN(n5364) );
  NAND2_X1 U6808 ( .A1(n8648), .A2(n8239), .ZN(n8189) );
  INV_X1 U6809 ( .A(n5366), .ZN(n5367) );
  NOR2_X1 U6810 ( .A1(n5368), .A2(n5367), .ZN(n5369) );
  AOI21_X1 U6811 ( .B1(n8190), .B2(n8189), .A(n5369), .ZN(n5397) );
  INV_X1 U6812 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5373) );
  INV_X1 U6813 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7264) );
  MUX2_X1 U6814 ( .A(n5373), .B(n7264), .S(n5561), .Z(n5375) );
  INV_X1 U6815 ( .A(SI_23_), .ZN(n5374) );
  NAND2_X1 U6816 ( .A1(n5375), .A2(n5374), .ZN(n5382) );
  INV_X1 U6817 ( .A(n5375), .ZN(n5376) );
  NAND2_X1 U6818 ( .A1(n5376), .A2(SI_23_), .ZN(n5377) );
  NAND2_X1 U6819 ( .A1(n7261), .A2(n8231), .ZN(n5379) );
  NAND2_X1 U6820 ( .A1(n5328), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5378) );
  XNOR2_X1 U6821 ( .A(n8618), .B(n5459), .ZN(n5398) );
  AND2_X1 U6822 ( .A1(n5397), .A2(n5398), .ZN(n8161) );
  INV_X1 U6823 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7334) );
  INV_X1 U6824 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7360) );
  MUX2_X1 U6825 ( .A(n7334), .B(n7360), .S(n5561), .Z(n5414) );
  XNOR2_X1 U6826 ( .A(n5414), .B(SI_24_), .ZN(n5411) );
  XNOR2_X1 U6827 ( .A(n5413), .B(n5411), .ZN(n7333) );
  NAND2_X1 U6828 ( .A1(n7333), .A2(n4266), .ZN(n5385) );
  NAND2_X1 U6829 ( .A1(n4902), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5384) );
  XNOR2_X1 U6830 ( .A(n8747), .B(n5459), .ZN(n5394) );
  INV_X1 U6831 ( .A(n5394), .ZN(n8163) );
  INV_X1 U6832 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8106) );
  INV_X1 U6833 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8171) );
  NAND2_X1 U6834 ( .A1(n5402), .A2(n8171), .ZN(n5387) );
  NAND2_X1 U6835 ( .A1(n5441), .A2(n5387), .ZN(n8598) );
  OR2_X1 U6836 ( .A1(n8598), .A2(n5463), .ZN(n5392) );
  INV_X1 U6837 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8597) );
  NAND2_X1 U6838 ( .A1(n6329), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5389) );
  NAND2_X1 U6839 ( .A1(n6327), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5388) );
  OAI211_X1 U6840 ( .C1(n8597), .C2(n5530), .A(n5389), .B(n5388), .ZN(n5390)
         );
  INV_X1 U6841 ( .A(n5390), .ZN(n5391) );
  NOR2_X1 U6842 ( .A1(n8165), .A2(n5481), .ZN(n5393) );
  INV_X1 U6843 ( .A(n5393), .ZN(n8167) );
  NAND2_X1 U6844 ( .A1(n8163), .A2(n8167), .ZN(n5396) );
  AND2_X1 U6845 ( .A1(n5394), .A2(n5393), .ZN(n5395) );
  AOI21_X1 U6846 ( .B1(n8161), .B2(n5396), .A(n5395), .ZN(n5410) );
  INV_X1 U6847 ( .A(n5397), .ZN(n5399) );
  NAND2_X1 U6848 ( .A1(n5400), .A2(n8106), .ZN(n5401) );
  AND2_X1 U6849 ( .A1(n5402), .A2(n5401), .ZN(n8617) );
  NAND2_X1 U6850 ( .A1(n8617), .A2(n5532), .ZN(n5408) );
  INV_X1 U6851 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U6852 ( .A1(n6329), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5404) );
  NAND2_X1 U6853 ( .A1(n6327), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5403) );
  OAI211_X1 U6854 ( .C1(n5405), .C2(n5530), .A(n5404), .B(n5403), .ZN(n5406)
         );
  INV_X1 U6855 ( .A(n5406), .ZN(n5407) );
  NAND2_X1 U6856 ( .A1(n8634), .A2(n8239), .ZN(n8101) );
  AOI21_X1 U6857 ( .B1(n8163), .B2(n8165), .A(n8101), .ZN(n5409) );
  INV_X1 U6858 ( .A(n5411), .ZN(n5412) );
  INV_X1 U6859 ( .A(n5414), .ZN(n5415) );
  NAND2_X1 U6860 ( .A1(n5415), .A2(SI_24_), .ZN(n5416) );
  INV_X1 U6861 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7539) );
  MUX2_X1 U6862 ( .A(n8907), .B(n7539), .S(n5561), .Z(n5418) );
  INV_X1 U6863 ( .A(SI_25_), .ZN(n5417) );
  NAND2_X1 U6864 ( .A1(n5418), .A2(n5417), .ZN(n5431) );
  INV_X1 U6865 ( .A(n5418), .ZN(n5419) );
  NAND2_X1 U6866 ( .A1(n5419), .A2(SI_25_), .ZN(n5420) );
  NAND2_X1 U6867 ( .A1(n5431), .A2(n5420), .ZN(n5432) );
  NAND2_X1 U6868 ( .A1(n7535), .A2(n4266), .ZN(n5422) );
  NAND2_X1 U6869 ( .A1(n5328), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5421) );
  NAND2_X2 U6870 ( .A1(n5422), .A2(n5421), .ZN(n8742) );
  XNOR2_X1 U6871 ( .A(n8742), .B(n5459), .ZN(n8137) );
  XNOR2_X1 U6872 ( .A(n5441), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n8145) );
  NAND2_X1 U6873 ( .A1(n8145), .A2(n5532), .ZN(n5427) );
  NAND2_X1 U6874 ( .A1(n6327), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5424) );
  OAI211_X1 U6875 ( .C1(n5530), .C2(n8882), .A(n5424), .B(n5423), .ZN(n5425)
         );
  INV_X1 U6876 ( .A(n5425), .ZN(n5426) );
  NOR2_X1 U6877 ( .A1(n8561), .A2(n5481), .ZN(n5428) );
  AND2_X1 U6878 ( .A1(n8137), .A2(n5428), .ZN(n8135) );
  INV_X1 U6879 ( .A(n8137), .ZN(n5430) );
  INV_X1 U6880 ( .A(n5428), .ZN(n5429) );
  NAND2_X1 U6881 ( .A1(n5430), .A2(n5429), .ZN(n8139) );
  INV_X1 U6882 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7541) );
  INV_X1 U6883 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7557) );
  MUX2_X1 U6884 ( .A(n7541), .B(n7557), .S(n5561), .Z(n5435) );
  INV_X1 U6885 ( .A(SI_26_), .ZN(n5434) );
  NAND2_X1 U6886 ( .A1(n5435), .A2(n5434), .ZN(n5452) );
  INV_X1 U6887 ( .A(n5435), .ZN(n5436) );
  NAND2_X1 U6888 ( .A1(n5436), .A2(SI_26_), .ZN(n5437) );
  NAND2_X1 U6889 ( .A1(n7540), .A2(n8231), .ZN(n5439) );
  NAND2_X1 U6890 ( .A1(n5328), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5438) );
  XNOR2_X1 U6891 ( .A(n8737), .B(n5459), .ZN(n5449) );
  INV_X1 U6892 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8146) );
  INV_X1 U6893 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8218) );
  OAI21_X1 U6894 ( .B1(n5441), .B2(n8146), .A(n8218), .ZN(n5442) );
  NAND2_X1 U6895 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG3_REG_26__SCAN_IN), 
        .ZN(n5440) );
  AND2_X1 U6896 ( .A1(n5442), .A2(n5461), .ZN(n8217) );
  INV_X1 U6897 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n5446) );
  NAND2_X1 U6898 ( .A1(n6329), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5445) );
  NAND2_X1 U6899 ( .A1(n6327), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5444) );
  OAI211_X1 U6900 ( .C1(n5446), .C2(n5530), .A(n5445), .B(n5444), .ZN(n5447)
         );
  AOI21_X1 U6901 ( .B1(n8217), .B2(n5532), .A(n5447), .ZN(n8144) );
  NOR2_X1 U6902 ( .A1(n8144), .A2(n5481), .ZN(n5448) );
  XNOR2_X1 U6903 ( .A(n5449), .B(n5448), .ZN(n8215) );
  INV_X1 U6904 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7596) );
  INV_X1 U6905 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n6090) );
  MUX2_X1 U6906 ( .A(n7596), .B(n6090), .S(n5561), .Z(n5454) );
  INV_X1 U6907 ( .A(SI_27_), .ZN(n8888) );
  NAND2_X1 U6908 ( .A1(n5454), .A2(n8888), .ZN(n5518) );
  INV_X1 U6909 ( .A(n5454), .ZN(n5455) );
  NAND2_X1 U6910 ( .A1(n5455), .A2(SI_27_), .ZN(n5456) );
  NAND2_X1 U6911 ( .A1(n7592), .A2(n4266), .ZN(n5458) );
  NAND2_X1 U6912 ( .A1(n5328), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5457) );
  XNOR2_X1 U6913 ( .A(n8732), .B(n5459), .ZN(n5471) );
  INV_X1 U6914 ( .A(n5461), .ZN(n5460) );
  NAND2_X1 U6915 ( .A1(n5460), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5475) );
  INV_X1 U6916 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8095) );
  NAND2_X1 U6917 ( .A1(n5461), .A2(n8095), .ZN(n5462) );
  NAND2_X1 U6918 ( .A1(n5475), .A2(n5462), .ZN(n8542) );
  INV_X1 U6919 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8541) );
  NAND2_X1 U6920 ( .A1(n6327), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5464) );
  OAI211_X1 U6921 ( .C1(n8541), .C2(n5530), .A(n5465), .B(n5464), .ZN(n5466)
         );
  INV_X1 U6922 ( .A(n5466), .ZN(n5467) );
  NAND2_X1 U6923 ( .A1(n8530), .A2(n8239), .ZN(n5469) );
  XNOR2_X1 U6924 ( .A(n5471), .B(n5469), .ZN(n8093) );
  NAND2_X1 U6925 ( .A1(n8094), .A2(n8093), .ZN(n5473) );
  INV_X1 U6926 ( .A(n5469), .ZN(n5470) );
  NAND2_X1 U6927 ( .A1(n5471), .A2(n5470), .ZN(n5472) );
  NAND2_X1 U6928 ( .A1(n5473), .A2(n5472), .ZN(n5485) );
  INV_X1 U6929 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U6930 ( .A1(n5475), .A2(n5474), .ZN(n5476) );
  INV_X1 U6931 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n5479) );
  NAND2_X1 U6932 ( .A1(n6329), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5478) );
  NAND2_X1 U6933 ( .A1(n6327), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5477) );
  OAI211_X1 U6934 ( .C1(n5479), .C2(n5530), .A(n5478), .B(n5477), .ZN(n5480)
         );
  OR2_X1 U6935 ( .A1(n8096), .A2(n5481), .ZN(n5483) );
  XNOR2_X1 U6936 ( .A(n5483), .B(n5482), .ZN(n5484) );
  XNOR2_X1 U6937 ( .A(n5485), .B(n5484), .ZN(n5542) );
  INV_X1 U6938 ( .A(n5542), .ZN(n5515) );
  NAND2_X1 U6939 ( .A1(n5487), .A2(n5486), .ZN(n5488) );
  INV_X1 U6940 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5490) );
  NAND2_X1 U6941 ( .A1(n4344), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5492) );
  MUX2_X1 U6942 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5492), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5493) );
  NAND2_X1 U6943 ( .A1(n5493), .A2(n4866), .ZN(n7542) );
  AND2_X1 U6944 ( .A1(n7335), .A2(n7542), .ZN(n9892) );
  INV_X1 U6945 ( .A(n7542), .ZN(n5500) );
  NAND2_X1 U6946 ( .A1(n5494), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5495) );
  MUX2_X1 U6947 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5495), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5496) );
  NAND2_X1 U6948 ( .A1(n5496), .A2(n4344), .ZN(n7536) );
  INV_X1 U6949 ( .A(P2_B_REG_SCAN_IN), .ZN(n5497) );
  XOR2_X1 U6950 ( .A(n7335), .B(n5497), .Z(n5498) );
  NAND2_X1 U6951 ( .A1(n7536), .A2(n5498), .ZN(n5499) );
  NOR2_X1 U6952 ( .A1(n9885), .A2(P2_D_REG_0__SCAN_IN), .ZN(n5501) );
  NOR4_X1 U6953 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n5505) );
  NOR4_X1 U6954 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5504) );
  NOR4_X1 U6955 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n5503) );
  NOR4_X1 U6956 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n5502) );
  AND4_X1 U6957 ( .A1(n5505), .A2(n5504), .A3(n5503), .A4(n5502), .ZN(n5510)
         );
  NOR2_X1 U6958 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .ZN(
        n8928) );
  NOR4_X1 U6959 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5508) );
  NOR4_X1 U6960 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n5507) );
  NOR4_X1 U6961 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n5506) );
  AND4_X1 U6962 ( .A1(n8928), .A2(n5508), .A3(n5507), .A4(n5506), .ZN(n5509)
         );
  AOI21_X1 U6963 ( .B1(n5510), .B2(n5509), .A(n9885), .ZN(n6571) );
  NAND2_X1 U6964 ( .A1(n7542), .A2(n7536), .ZN(n9895) );
  OAI21_X1 U6965 ( .B1(P2_D_REG_1__SCAN_IN), .B2(n9885), .A(n9895), .ZN(n6570)
         );
  NOR2_X1 U6966 ( .A1(n6571), .A2(n6570), .ZN(n6874) );
  INV_X1 U6967 ( .A(n6874), .ZN(n5511) );
  INV_X1 U6968 ( .A(n5536), .ZN(n5514) );
  XNOR2_X1 U6969 ( .A(n5513), .B(n5512), .ZN(n6180) );
  NAND2_X1 U6970 ( .A1(n5514), .A2(n9886), .ZN(n5533) );
  INV_X1 U6971 ( .A(n8399), .ZN(n9899) );
  OR3_X2 U6972 ( .A1(n5533), .A2(n9475), .A3(n6581), .ZN(n9835) );
  NAND2_X1 U6973 ( .A1(n5515), .A2(n9845), .ZN(n5543) );
  INV_X1 U6974 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7773) );
  INV_X1 U6975 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5519) );
  MUX2_X1 U6976 ( .A(n7773), .B(n5519), .S(n7715), .Z(n5521) );
  INV_X1 U6977 ( .A(SI_28_), .ZN(n5520) );
  NAND2_X1 U6978 ( .A1(n5521), .A2(n5520), .ZN(n7696) );
  INV_X1 U6979 ( .A(n5521), .ZN(n5522) );
  NAND2_X1 U6980 ( .A1(n5522), .A2(SI_28_), .ZN(n5523) );
  NAND2_X1 U6981 ( .A1(n7772), .A2(n4266), .ZN(n5525) );
  NAND2_X1 U6982 ( .A1(n5328), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5524) );
  INV_X1 U6983 ( .A(n5526), .ZN(n8068) );
  INV_X1 U6984 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n5529) );
  NAND2_X1 U6985 ( .A1(n6327), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5528) );
  OAI211_X1 U6986 ( .C1(n5530), .C2(n5529), .A(n5528), .B(n5527), .ZN(n5531)
         );
  AOI21_X1 U6987 ( .B1(n8068), .B2(n5532), .A(n5531), .ZN(n8065) );
  INV_X1 U6988 ( .A(n8065), .ZN(n8529) );
  OR2_X1 U6989 ( .A1(n5533), .A2(n8442), .ZN(n8209) );
  INV_X1 U6990 ( .A(n6581), .ZN(n6179) );
  INV_X1 U6991 ( .A(n5534), .ZN(n6186) );
  INV_X1 U6992 ( .A(n8219), .ZN(n9828) );
  INV_X1 U6993 ( .A(n9831), .ZN(n8194) );
  AOI22_X1 U6994 ( .A1(n8529), .A2(n9828), .B1(n8530), .B2(n8194), .ZN(n5540)
         );
  NAND2_X1 U6995 ( .A1(n5536), .A2(n6878), .ZN(n5541) );
  NAND2_X1 U6996 ( .A1(n8442), .A2(n6581), .ZN(n6619) );
  AND3_X1 U6997 ( .A1(n6181), .A2(n6180), .A3(n6619), .ZN(n5537) );
  NAND2_X1 U6998 ( .A1(n5541), .A2(n5537), .ZN(n5538) );
  INV_X1 U6999 ( .A(n9860), .ZN(n8211) );
  AOI22_X1 U7000 ( .A1(n8525), .A2(n8211), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n5539) );
  AND2_X1 U7001 ( .A1(n5541), .A2(n9886), .ZN(n9478) );
  NAND3_X1 U7002 ( .A1(n5565), .A2(n5566), .A3(n5548), .ZN(n5554) );
  NOR2_X1 U7003 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5552) );
  NOR2_X1 U7004 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5551) );
  NOR2_X1 U7005 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5550) );
  NOR2_X1 U7006 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5549) );
  NAND4_X1 U7007 ( .A1(n5552), .A2(n5551), .A3(n5550), .A4(n5549), .ZN(n5553)
         );
  XNOR2_X2 U7008 ( .A(n5560), .B(n5559), .ZN(n9546) );
  NAND2_X4 U7009 ( .A1(n6140), .A2(n9546), .ZN(n6167) );
  NAND2_X1 U7010 ( .A1(n7333), .A2(n7777), .ZN(n5563) );
  OR2_X1 U7011 ( .A1(n5663), .A2(n7360), .ZN(n5562) );
  NOR2_X1 U7012 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5564) );
  INV_X1 U7013 ( .A(n5570), .ZN(n5568) );
  NAND2_X1 U7014 ( .A1(n5568), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n5571) );
  NAND2_X1 U7015 ( .A1(n5574), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5576) );
  INV_X1 U7016 ( .A(n7559), .ZN(n5585) );
  BUF_X1 U7017 ( .A(n5577), .Z(n5578) );
  NAND2_X1 U7018 ( .A1(n5578), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5579) );
  MUX2_X1 U7019 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5579), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5581) );
  INV_X1 U7020 ( .A(n5580), .ZN(n5582) );
  INV_X1 U7021 ( .A(n7358), .ZN(n5584) );
  NAND2_X1 U7022 ( .A1(n5582), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5583) );
  XNOR2_X1 U7023 ( .A(n5583), .B(P1_IR_REG_25__SCAN_IN), .ZN(n6127) );
  INV_X1 U7024 ( .A(n6165), .ZN(n5621) );
  NOR2_X2 U7025 ( .A1(n6723), .A2(n5621), .ZN(n5643) );
  INV_X4 U7026 ( .A(n6055), .ZN(n8995) );
  AND2_X2 U7027 ( .A1(n6723), .A2(n6165), .ZN(n5625) );
  XNOR2_X2 U7028 ( .A(n5591), .B(n5590), .ZN(n9137) );
  NAND2_X1 U7029 ( .A1(n6132), .A2(n7977), .ZN(n5592) );
  NOR2_X1 U7030 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n5593) );
  NAND2_X1 U7031 ( .A1(n5596), .A2(n5593), .ZN(n9443) );
  XNOR2_X2 U7032 ( .A(n5595), .B(n5594), .ZN(n8047) );
  AOI21_X1 U7033 ( .B1(n5596), .B2(n5559), .A(n5934), .ZN(n5597) );
  XNOR2_X2 U7034 ( .A(n5598), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5602) );
  NAND2_X1 U7035 ( .A1(n5675), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5608) );
  AND2_X4 U7036 ( .A1(n5602), .A2(n5603), .ZN(n7783) );
  INV_X1 U7037 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5601) );
  NAND2_X1 U7038 ( .A1(n5735), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U7039 ( .A1(n5774), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5791) );
  NAND2_X1 U7040 ( .A1(n5856), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5878) );
  INV_X1 U7041 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5877) );
  INV_X1 U7042 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9047) );
  INV_X1 U7043 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5973) );
  AND2_X1 U7044 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n5599) );
  NAND2_X1 U7045 ( .A1(n6044), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6045) );
  INV_X1 U7046 ( .A(n6045), .ZN(n5600) );
  AOI21_X1 U7047 ( .B1(n5601), .B2(n6045), .A(n6062), .ZN(n9215) );
  NAND2_X1 U7048 ( .A1(n7783), .A2(n9215), .ZN(n5607) );
  AND2_X2 U7049 ( .A1(n5603), .A2(n7701), .ZN(n5654) );
  BUF_X2 U7050 ( .A(n5654), .Z(n6153) );
  INV_X1 U7051 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n5604) );
  OR2_X1 U7052 ( .A1(n6098), .A2(n5604), .ZN(n5606) );
  NAND2_X1 U7053 ( .A1(n7723), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5605) );
  NAND4_X1 U7054 ( .A1(n5608), .A2(n5607), .A3(n5606), .A4(n5605), .ZN(n9206)
         );
  AOI22_X1 U7055 ( .A1(n9366), .A2(n8995), .B1(n8996), .B2(n9206), .ZN(n6059)
         );
  INV_X2 U7056 ( .A(n5637), .ZN(n9002) );
  AOI22_X1 U7057 ( .A1(n9366), .A2(n9002), .B1(n8995), .B2(n9206), .ZN(n5609)
         );
  NAND2_X2 U7058 ( .A1(n6724), .A2(n6723), .ZN(n8999) );
  XNOR2_X1 U7059 ( .A(n5609), .B(n8999), .ZN(n6058) );
  NAND2_X1 U7060 ( .A1(n7783), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5614) );
  NAND2_X1 U7061 ( .A1(n5676), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5612) );
  NAND2_X1 U7062 ( .A1(n5654), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U7063 ( .A1(n5675), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5610) );
  AND3_X1 U7064 ( .A1(n5612), .A2(n5611), .A3(n5610), .ZN(n5613) );
  NAND2_X2 U7065 ( .A1(n5614), .A2(n5613), .ZN(n9728) );
  INV_X1 U7066 ( .A(SI_0_), .ZN(n5616) );
  INV_X1 U7067 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5615) );
  OAI21_X1 U7068 ( .B1(n7715), .B2(n5616), .A(n5615), .ZN(n5618) );
  AND2_X1 U7069 ( .A1(n5617), .A2(n5618), .ZN(n9450) );
  NAND2_X1 U7070 ( .A1(n6800), .A2(n5643), .ZN(n5623) );
  NAND2_X1 U7071 ( .A1(n5621), .A2(n9556), .ZN(n5622) );
  NAND2_X1 U7072 ( .A1(n9728), .A2(n5643), .ZN(n5629) );
  INV_X1 U7073 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9555) );
  NAND2_X1 U7074 ( .A1(n6800), .A2(n5625), .ZN(n5626) );
  OAI21_X1 U7075 ( .B1(n6165), .B2(n9555), .A(n5626), .ZN(n5627) );
  NAND2_X1 U7076 ( .A1(n5629), .A2(n5628), .ZN(n5630) );
  NAND2_X1 U7077 ( .A1(n6433), .A2(n5630), .ZN(n6432) );
  INV_X1 U7078 ( .A(n5630), .ZN(n6431) );
  NAND2_X1 U7079 ( .A1(n6431), .A2(n8999), .ZN(n5631) );
  INV_X1 U7080 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6293) );
  INV_X1 U7081 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5633) );
  NAND2_X1 U7082 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n9556), .ZN(n5632) );
  XNOR2_X1 U7083 ( .A(n5633), .B(n5632), .ZN(n9560) );
  NAND2_X1 U7084 ( .A1(n9719), .A2(n5625), .ZN(n5645) );
  NAND2_X1 U7085 ( .A1(n7783), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5642) );
  NAND2_X1 U7086 ( .A1(n5676), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5640) );
  NAND2_X1 U7087 ( .A1(n5654), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5639) );
  NAND2_X1 U7088 ( .A1(n5675), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5638) );
  AND3_X1 U7089 ( .A1(n5640), .A2(n5639), .A3(n5638), .ZN(n5641) );
  NAND2_X2 U7090 ( .A1(n5642), .A2(n5641), .ZN(n6715) );
  NAND2_X1 U7091 ( .A1(n6715), .A2(n5643), .ZN(n5644) );
  NAND2_X1 U7092 ( .A1(n5645), .A2(n5644), .ZN(n5646) );
  NAND2_X1 U7093 ( .A1(n6715), .A2(n8996), .ZN(n5648) );
  NAND2_X1 U7094 ( .A1(n9719), .A2(n9001), .ZN(n5647) );
  NAND2_X1 U7095 ( .A1(n5648), .A2(n5647), .ZN(n9022) );
  NAND2_X1 U7096 ( .A1(n9020), .A2(n9022), .ZN(n5653) );
  NAND2_X1 U7097 ( .A1(n5675), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5659) );
  NAND2_X1 U7098 ( .A1(n7783), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5658) );
  NAND2_X1 U7099 ( .A1(n5676), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5657) );
  INV_X1 U7100 ( .A(n5654), .ZN(n5655) );
  INV_X1 U7101 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6341) );
  OR2_X1 U7102 ( .A1(n5655), .A2(n6341), .ZN(n5656) );
  NAND4_X2 U7103 ( .A1(n5659), .A2(n5658), .A3(n5657), .A4(n5656), .ZN(n9727)
         );
  NAND2_X1 U7104 ( .A1(n9727), .A2(n5643), .ZN(n5669) );
  INV_X1 U7105 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U7106 ( .A1(n5662), .A2(n5661), .ZN(n5681) );
  OAI21_X1 U7107 ( .B1(n5662), .B2(n5661), .A(n5681), .ZN(n9576) );
  INV_X1 U7108 ( .A(n5663), .ZN(n5664) );
  OR2_X1 U7109 ( .A1(n5665), .A2(n6294), .ZN(n5666) );
  NAND2_X1 U7110 ( .A1(n6936), .A2(n5625), .ZN(n5668) );
  NAND2_X1 U7111 ( .A1(n5669), .A2(n5668), .ZN(n5670) );
  XNOR2_X1 U7112 ( .A(n5670), .B(n8999), .ZN(n5671) );
  AOI22_X1 U7113 ( .A1(n9727), .A2(n8996), .B1(n9001), .B2(n6936), .ZN(n5672)
         );
  XNOR2_X1 U7114 ( .A(n5671), .B(n5672), .ZN(n6526) );
  INV_X1 U7115 ( .A(n5671), .ZN(n5673) );
  NAND2_X1 U7116 ( .A1(n5673), .A2(n5672), .ZN(n5674) );
  INV_X1 U7117 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n8917) );
  NAND2_X1 U7118 ( .A1(n7783), .A2(n8917), .ZN(n5680) );
  NAND2_X1 U7119 ( .A1(n5675), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U7120 ( .A1(n5676), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U7121 ( .A1(n9125), .A2(n9001), .ZN(n5687) );
  NAND2_X1 U7122 ( .A1(n5681), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5683) );
  INV_X1 U7123 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5682) );
  OR2_X1 U7124 ( .A1(n5663), .A2(n6297), .ZN(n5685) );
  OR2_X1 U7125 ( .A1(n5665), .A2(n6296), .ZN(n5684) );
  OAI211_X1 U7126 ( .C1(n6167), .C2(n6412), .A(n5685), .B(n5684), .ZN(n6926)
         );
  NAND2_X1 U7127 ( .A1(n6926), .A2(n9002), .ZN(n5686) );
  NAND2_X1 U7128 ( .A1(n5687), .A2(n5686), .ZN(n5688) );
  XNOR2_X1 U7129 ( .A(n5688), .B(n8999), .ZN(n5689) );
  AOI22_X1 U7130 ( .A1(n9125), .A2(n8996), .B1(n8995), .B2(n6926), .ZN(n5690)
         );
  XNOR2_X1 U7131 ( .A(n5689), .B(n5690), .ZN(n6531) );
  NAND2_X1 U7132 ( .A1(n6532), .A2(n6531), .ZN(n5693) );
  INV_X1 U7133 ( .A(n5689), .ZN(n5691) );
  NAND2_X1 U7134 ( .A1(n5691), .A2(n5690), .ZN(n5692) );
  NAND2_X1 U7135 ( .A1(n5693), .A2(n5692), .ZN(n6679) );
  INV_X1 U7136 ( .A(n6679), .ZN(n5712) );
  NAND2_X1 U7137 ( .A1(n6148), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5699) );
  INV_X1 U7138 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5694) );
  XNOR2_X1 U7139 ( .A(n5694), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n6933) );
  NAND2_X1 U7140 ( .A1(n7783), .A2(n6933), .ZN(n5698) );
  NAND2_X1 U7141 ( .A1(n6153), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5697) );
  INV_X1 U7142 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5695) );
  NAND4_X1 U7143 ( .A1(n5699), .A2(n5698), .A3(n5697), .A4(n5696), .ZN(n9675)
         );
  NAND2_X1 U7144 ( .A1(n9675), .A2(n8995), .ZN(n5708) );
  NOR2_X1 U7145 ( .A1(n5700), .A2(n5934), .ZN(n5701) );
  MUX2_X1 U7146 ( .A(n5934), .B(n5701), .S(P1_IR_REG_4__SCAN_IN), .Z(n5702) );
  INV_X1 U7147 ( .A(n5702), .ZN(n5704) );
  INV_X1 U7148 ( .A(n5723), .ZN(n5703) );
  NAND2_X1 U7149 ( .A1(n5704), .A2(n5703), .ZN(n6364) );
  OR2_X1 U7150 ( .A1(n7779), .A2(n6298), .ZN(n5706) );
  OR2_X1 U7151 ( .A1(n5665), .A2(n6300), .ZN(n5705) );
  NAND2_X1 U7152 ( .A1(n6934), .A2(n9002), .ZN(n5707) );
  NAND2_X1 U7153 ( .A1(n5708), .A2(n5707), .ZN(n5710) );
  XNOR2_X1 U7154 ( .A(n5710), .B(n6105), .ZN(n5713) );
  AOI22_X1 U7155 ( .A1(n9675), .A2(n8996), .B1(n8995), .B2(n6934), .ZN(n5714)
         );
  XNOR2_X1 U7156 ( .A(n5713), .B(n5714), .ZN(n6682) );
  NAND2_X1 U7157 ( .A1(n5712), .A2(n5711), .ZN(n6680) );
  INV_X1 U7158 ( .A(n5713), .ZN(n5716) );
  INV_X1 U7159 ( .A(n5714), .ZN(n5715) );
  NAND2_X1 U7160 ( .A1(n5716), .A2(n5715), .ZN(n5717) );
  NAND2_X1 U7161 ( .A1(n6148), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5722) );
  AOI21_X1 U7162 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5718) );
  NOR2_X1 U7163 ( .A1(n5718), .A2(n5735), .ZN(n9686) );
  NAND2_X1 U7164 ( .A1(n7783), .A2(n9686), .ZN(n5721) );
  NAND2_X1 U7165 ( .A1(n6153), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5720) );
  NAND2_X1 U7166 ( .A1(n7723), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5719) );
  NAND4_X1 U7167 ( .A1(n5722), .A2(n5721), .A3(n5720), .A4(n5719), .ZN(n9124)
         );
  NAND2_X1 U7168 ( .A1(n9124), .A2(n8995), .ZN(n5729) );
  OR2_X1 U7169 ( .A1(n5723), .A2(n5934), .ZN(n5725) );
  XNOR2_X1 U7170 ( .A(n5725), .B(n5724), .ZN(n6459) );
  OR2_X1 U7171 ( .A1(n7779), .A2(n6302), .ZN(n5727) );
  OR2_X1 U7172 ( .A1(n5665), .A2(n6304), .ZN(n5726) );
  OAI211_X1 U7173 ( .C1(n6167), .C2(n6459), .A(n5727), .B(n5726), .ZN(n9687)
         );
  NAND2_X1 U7174 ( .A1(n9687), .A2(n9002), .ZN(n5728) );
  NAND2_X1 U7175 ( .A1(n5729), .A2(n5728), .ZN(n5730) );
  XNOR2_X1 U7176 ( .A(n5730), .B(n6105), .ZN(n5731) );
  AOI22_X1 U7177 ( .A1(n9124), .A2(n8996), .B1(n8995), .B2(n9687), .ZN(n6702)
         );
  INV_X1 U7178 ( .A(n5731), .ZN(n5732) );
  NAND2_X1 U7179 ( .A1(n6701), .A2(n5734), .ZN(n6812) );
  INV_X2 U7180 ( .A(n6049), .ZN(n6148) );
  NAND2_X1 U7181 ( .A1(n6148), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5740) );
  OAI21_X1 U7182 ( .B1(n5735), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5756), .ZN(
        n6816) );
  INV_X1 U7183 ( .A(n6816), .ZN(n7052) );
  NAND2_X1 U7184 ( .A1(n7783), .A2(n7052), .ZN(n5739) );
  INV_X1 U7185 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5736) );
  OR2_X1 U7186 ( .A1(n6098), .A2(n5736), .ZN(n5738) );
  NAND2_X1 U7187 ( .A1(n7723), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5737) );
  NAND2_X1 U7188 ( .A1(n9676), .A2(n8995), .ZN(n5748) );
  NAND2_X1 U7189 ( .A1(n5743), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5742) );
  MUX2_X1 U7190 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5742), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n5744) );
  OR2_X1 U7191 ( .A1(n5743), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5770) );
  AND2_X1 U7192 ( .A1(n5744), .A2(n5770), .ZN(n6383) );
  INV_X1 U7193 ( .A(n6383), .ZN(n6366) );
  OR2_X1 U7194 ( .A1(n5665), .A2(n6308), .ZN(n5746) );
  OR2_X1 U7195 ( .A1(n7779), .A2(n6309), .ZN(n5745) );
  NAND2_X1 U7196 ( .A1(n7053), .A2(n9002), .ZN(n5747) );
  NAND2_X1 U7197 ( .A1(n5748), .A2(n5747), .ZN(n5749) );
  XNOR2_X1 U7198 ( .A(n5749), .B(n8999), .ZN(n5750) );
  AOI22_X1 U7199 ( .A1(n9676), .A2(n8996), .B1(n8995), .B2(n7053), .ZN(n5751)
         );
  XNOR2_X1 U7200 ( .A(n5750), .B(n5751), .ZN(n6811) );
  NAND2_X1 U7201 ( .A1(n6812), .A2(n6811), .ZN(n5754) );
  INV_X1 U7202 ( .A(n5750), .ZN(n5752) );
  NAND2_X1 U7203 ( .A1(n5752), .A2(n5751), .ZN(n5753) );
  NAND2_X1 U7204 ( .A1(n5754), .A2(n5753), .ZN(n6863) );
  NAND2_X1 U7205 ( .A1(n6148), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5761) );
  AND2_X1 U7206 ( .A1(n5756), .A2(n5755), .ZN(n5757) );
  NOR2_X1 U7207 ( .A1(n5774), .A2(n5757), .ZN(n6867) );
  NAND2_X1 U7208 ( .A1(n7783), .A2(n6867), .ZN(n5760) );
  INV_X1 U7209 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7177) );
  OR2_X1 U7210 ( .A1(n6098), .A2(n7177), .ZN(n5759) );
  NAND2_X1 U7211 ( .A1(n7723), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5758) );
  NAND4_X1 U7212 ( .A1(n5761), .A2(n5760), .A3(n5759), .A4(n5758), .ZN(n9123)
         );
  NAND2_X1 U7213 ( .A1(n9123), .A2(n8995), .ZN(n5766) );
  NAND2_X1 U7214 ( .A1(n5770), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5762) );
  XNOR2_X1 U7215 ( .A(n5762), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6387) );
  INV_X1 U7216 ( .A(n6387), .ZN(n6394) );
  NAND2_X1 U7217 ( .A1(n6315), .A2(n7777), .ZN(n5764) );
  INV_X1 U7218 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6317) );
  OR2_X1 U7219 ( .A1(n7779), .A2(n6317), .ZN(n5763) );
  NAND2_X1 U7220 ( .A1(n7179), .A2(n9002), .ZN(n5765) );
  NAND2_X1 U7221 ( .A1(n5766), .A2(n5765), .ZN(n5767) );
  XNOR2_X1 U7222 ( .A(n5767), .B(n6105), .ZN(n6865) );
  NAND2_X1 U7223 ( .A1(n9123), .A2(n8996), .ZN(n5769) );
  NAND2_X1 U7224 ( .A1(n7179), .A2(n8995), .ZN(n5768) );
  AND2_X1 U7225 ( .A1(n5769), .A2(n5768), .ZN(n6864) );
  AND2_X1 U7226 ( .A1(n6865), .A2(n6864), .ZN(n7028) );
  NAND2_X1 U7227 ( .A1(n6318), .A2(n7777), .ZN(n5773) );
  NOR2_X1 U7228 ( .A1(n5770), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5786) );
  OR2_X1 U7229 ( .A1(n5786), .A2(n5934), .ZN(n5771) );
  XNOR2_X1 U7230 ( .A(n5771), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6447) );
  AOI22_X1 U7231 ( .A1(n4270), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5635), .B2(
        n6447), .ZN(n5772) );
  NAND2_X1 U7232 ( .A1(n7194), .A2(n9002), .ZN(n5781) );
  NAND2_X1 U7233 ( .A1(n6148), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5779) );
  OR2_X1 U7234 ( .A1(n5774), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5775) );
  AND2_X1 U7235 ( .A1(n5791), .A2(n5775), .ZN(n7103) );
  NAND2_X1 U7236 ( .A1(n7783), .A2(n7103), .ZN(n5778) );
  INV_X1 U7237 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n8918) );
  OR2_X1 U7238 ( .A1(n6098), .A2(n8918), .ZN(n5777) );
  NAND2_X1 U7239 ( .A1(n7723), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5776) );
  NAND2_X1 U7240 ( .A1(n9122), .A2(n8995), .ZN(n5780) );
  NAND2_X1 U7241 ( .A1(n5781), .A2(n5780), .ZN(n5782) );
  XNOR2_X1 U7242 ( .A(n5782), .B(n6105), .ZN(n7032) );
  NAND2_X1 U7243 ( .A1(n7194), .A2(n8995), .ZN(n5784) );
  NAND2_X1 U7244 ( .A1(n9122), .A2(n8996), .ZN(n5783) );
  AND2_X1 U7245 ( .A1(n5784), .A2(n5783), .ZN(n5809) );
  AND2_X1 U7246 ( .A1(n7032), .A2(n5809), .ZN(n5813) );
  OR2_X1 U7247 ( .A1(n7028), .A2(n5813), .ZN(n7145) );
  NAND2_X1 U7248 ( .A1(n6322), .A2(n7777), .ZN(n5789) );
  NAND2_X1 U7249 ( .A1(n5786), .A2(n5785), .ZN(n5817) );
  NAND2_X1 U7250 ( .A1(n5817), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5787) );
  XNOR2_X1 U7251 ( .A(n5787), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9610) );
  AOI22_X1 U7252 ( .A1(n5664), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5635), .B2(
        n9610), .ZN(n5788) );
  NAND2_X1 U7253 ( .A1(n7315), .A2(n9002), .ZN(n5798) );
  NAND2_X1 U7254 ( .A1(n6148), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5796) );
  NAND2_X1 U7255 ( .A1(n5791), .A2(n5790), .ZN(n5792) );
  AND2_X1 U7256 ( .A1(n5821), .A2(n5792), .ZN(n7199) );
  NAND2_X1 U7257 ( .A1(n7783), .A2(n7199), .ZN(n5795) );
  NAND2_X1 U7258 ( .A1(n7723), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5794) );
  NAND2_X1 U7259 ( .A1(n6153), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5793) );
  NAND4_X1 U7260 ( .A1(n5796), .A2(n5795), .A3(n5794), .A4(n5793), .ZN(n9121)
         );
  NAND2_X1 U7261 ( .A1(n9121), .A2(n8995), .ZN(n5797) );
  NAND2_X1 U7262 ( .A1(n5798), .A2(n5797), .ZN(n5799) );
  XNOR2_X1 U7263 ( .A(n5799), .B(n6105), .ZN(n5801) );
  AND2_X1 U7264 ( .A1(n9121), .A2(n8996), .ZN(n5800) );
  AOI21_X1 U7265 ( .B1(n7315), .B2(n8995), .A(n5800), .ZN(n5802) );
  NAND2_X1 U7266 ( .A1(n5801), .A2(n5802), .ZN(n5806) );
  INV_X1 U7267 ( .A(n5806), .ZN(n5815) );
  INV_X1 U7268 ( .A(n5801), .ZN(n5804) );
  INV_X1 U7269 ( .A(n5802), .ZN(n5803) );
  NAND2_X1 U7270 ( .A1(n5804), .A2(n5803), .ZN(n5805) );
  NAND2_X1 U7271 ( .A1(n5806), .A2(n5805), .ZN(n7152) );
  INV_X1 U7272 ( .A(n7152), .ZN(n5814) );
  INV_X1 U7273 ( .A(n6865), .ZN(n5808) );
  INV_X1 U7274 ( .A(n6864), .ZN(n5807) );
  NAND2_X1 U7275 ( .A1(n5808), .A2(n5807), .ZN(n7029) );
  INV_X1 U7276 ( .A(n7032), .ZN(n5810) );
  INV_X1 U7277 ( .A(n5809), .ZN(n7031) );
  NAND2_X1 U7278 ( .A1(n5810), .A2(n7031), .ZN(n5811) );
  AND2_X1 U7279 ( .A1(n5811), .A2(n7029), .ZN(n5812) );
  OR2_X1 U7280 ( .A1(n5813), .A2(n5812), .ZN(n7147) );
  AND2_X1 U7281 ( .A1(n5814), .A2(n7147), .ZN(n7148) );
  NAND2_X1 U7282 ( .A1(n6325), .A2(n7777), .ZN(n5820) );
  OAI21_X1 U7283 ( .B1(n5817), .B2(P1_IR_REG_9__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5818) );
  XNOR2_X1 U7284 ( .A(n5818), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6485) );
  AOI22_X1 U7285 ( .A1(n5664), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5635), .B2(
        n6485), .ZN(n5819) );
  NAND2_X1 U7286 ( .A1(n7402), .A2(n9002), .ZN(n5828) );
  NAND2_X1 U7287 ( .A1(n6148), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5826) );
  NAND2_X1 U7288 ( .A1(n5821), .A2(n6445), .ZN(n5822) );
  AND2_X1 U7289 ( .A1(n5840), .A2(n5822), .ZN(n7310) );
  NAND2_X1 U7290 ( .A1(n7783), .A2(n7310), .ZN(n5825) );
  INV_X1 U7291 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6453) );
  OR2_X1 U7292 ( .A1(n6098), .A2(n6453), .ZN(n5824) );
  NAND2_X1 U7293 ( .A1(n7723), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5823) );
  NAND4_X1 U7294 ( .A1(n5826), .A2(n5825), .A3(n5824), .A4(n5823), .ZN(n9120)
         );
  NAND2_X1 U7295 ( .A1(n9120), .A2(n8995), .ZN(n5827) );
  NAND2_X1 U7296 ( .A1(n5828), .A2(n5827), .ZN(n5829) );
  XNOR2_X1 U7297 ( .A(n5829), .B(n6105), .ZN(n5834) );
  INV_X1 U7298 ( .A(n5834), .ZN(n5832) );
  AND2_X1 U7299 ( .A1(n9120), .A2(n8996), .ZN(n5830) );
  AOI21_X1 U7300 ( .B1(n7402), .B2(n9001), .A(n5830), .ZN(n5833) );
  INV_X1 U7301 ( .A(n5833), .ZN(n5831) );
  NAND2_X1 U7302 ( .A1(n5832), .A2(n5831), .ZN(n7136) );
  NAND2_X1 U7303 ( .A1(n6337), .A2(n7777), .ZN(n5838) );
  NAND2_X1 U7304 ( .A1(n5835), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5836) );
  XNOR2_X1 U7305 ( .A(n5836), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6492) );
  AOI22_X1 U7306 ( .A1(n5664), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5635), .B2(
        n6492), .ZN(n5837) );
  NAND2_X1 U7307 ( .A1(n7388), .A2(n9002), .ZN(n5847) );
  NAND2_X1 U7308 ( .A1(n6148), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5845) );
  AND2_X1 U7309 ( .A1(n5840), .A2(n5839), .ZN(n5841) );
  NOR2_X1 U7310 ( .A1(n5856), .A2(n5841), .ZN(n9518) );
  NAND2_X1 U7311 ( .A1(n7783), .A2(n9518), .ZN(n5844) );
  NAND2_X1 U7312 ( .A1(n7723), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5843) );
  OR2_X1 U7313 ( .A1(n6098), .A2(n6518), .ZN(n5842) );
  NAND4_X1 U7314 ( .A1(n5845), .A2(n5844), .A3(n5843), .A4(n5842), .ZN(n9455)
         );
  NAND2_X1 U7315 ( .A1(n9455), .A2(n8995), .ZN(n5846) );
  NAND2_X1 U7316 ( .A1(n5847), .A2(n5846), .ZN(n5848) );
  XNOR2_X1 U7317 ( .A(n5848), .B(n8999), .ZN(n5852) );
  AND2_X1 U7318 ( .A1(n9455), .A2(n8996), .ZN(n5849) );
  AOI21_X1 U7319 ( .B1(n7388), .B2(n8995), .A(n5849), .ZN(n5850) );
  XNOR2_X1 U7320 ( .A(n5852), .B(n5850), .ZN(n7229) );
  INV_X1 U7321 ( .A(n5850), .ZN(n5851) );
  NAND2_X1 U7322 ( .A1(n5852), .A2(n5851), .ZN(n5853) );
  NAND2_X1 U7323 ( .A1(n7228), .A2(n5853), .ZN(n9459) );
  NAND2_X1 U7324 ( .A1(n6420), .A2(n7777), .ZN(n5855) );
  OR2_X1 U7325 ( .A1(n4341), .A2(n5934), .ZN(n5891) );
  XNOR2_X1 U7326 ( .A(n5891), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6550) );
  AOI22_X1 U7327 ( .A1(n5664), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5635), .B2(
        n6550), .ZN(n5854) );
  NAND2_X1 U7328 ( .A1(n7560), .A2(n9002), .ZN(n5864) );
  OR2_X1 U7329 ( .A1(n5856), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5857) );
  NAND2_X1 U7330 ( .A1(n5878), .A2(n5857), .ZN(n9467) );
  INV_X1 U7331 ( .A(n9467), .ZN(n7395) );
  NAND2_X1 U7332 ( .A1(n7783), .A2(n7395), .ZN(n5862) );
  NAND2_X1 U7333 ( .A1(n6148), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5861) );
  NAND2_X1 U7334 ( .A1(n7723), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5860) );
  INV_X1 U7335 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n5858) );
  OR2_X1 U7336 ( .A1(n6098), .A2(n5858), .ZN(n5859) );
  NAND4_X1 U7337 ( .A1(n5862), .A2(n5861), .A3(n5860), .A4(n5859), .ZN(n9119)
         );
  NAND2_X1 U7338 ( .A1(n9119), .A2(n8995), .ZN(n5863) );
  NAND2_X1 U7339 ( .A1(n5864), .A2(n5863), .ZN(n5865) );
  XNOR2_X1 U7340 ( .A(n5865), .B(n6105), .ZN(n5870) );
  AND2_X1 U7341 ( .A1(n9119), .A2(n8996), .ZN(n5866) );
  AOI21_X1 U7342 ( .B1(n7560), .B2(n9001), .A(n5866), .ZN(n5869) );
  XNOR2_X1 U7343 ( .A(n5870), .B(n5869), .ZN(n9458) );
  NAND2_X1 U7344 ( .A1(n5870), .A2(n5869), .ZN(n5871) );
  NAND2_X1 U7345 ( .A1(n6507), .A2(n7777), .ZN(n5876) );
  INV_X1 U7346 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5872) );
  NAND2_X1 U7347 ( .A1(n5891), .A2(n5872), .ZN(n5873) );
  NAND2_X1 U7348 ( .A1(n5873), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5874) );
  XNOR2_X1 U7349 ( .A(n5874), .B(P1_IR_REG_13__SCAN_IN), .ZN(n6559) );
  AOI22_X1 U7350 ( .A1(n5664), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5635), .B2(
        n6559), .ZN(n5875) );
  NAND2_X1 U7351 ( .A1(n9499), .A2(n9002), .ZN(n5885) );
  NAND2_X1 U7352 ( .A1(n6148), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5883) );
  NAND2_X1 U7353 ( .A1(n5878), .A2(n5877), .ZN(n5879) );
  AND2_X1 U7354 ( .A1(n5898), .A2(n5879), .ZN(n9497) );
  NAND2_X1 U7355 ( .A1(n7783), .A2(n9497), .ZN(n5882) );
  NAND2_X1 U7356 ( .A1(n6153), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5881) );
  NAND2_X1 U7357 ( .A1(n7723), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5880) );
  NAND4_X1 U7358 ( .A1(n5883), .A2(n5882), .A3(n5881), .A4(n5880), .ZN(n9118)
         );
  NAND2_X1 U7359 ( .A1(n9118), .A2(n8995), .ZN(n5884) );
  NAND2_X1 U7360 ( .A1(n5885), .A2(n5884), .ZN(n5886) );
  XNOR2_X1 U7361 ( .A(n5886), .B(n6105), .ZN(n7423) );
  AND2_X1 U7362 ( .A1(n9118), .A2(n8996), .ZN(n5887) );
  AOI21_X1 U7363 ( .B1(n9499), .B2(n8995), .A(n5887), .ZN(n5888) );
  INV_X1 U7364 ( .A(n7423), .ZN(n5889) );
  INV_X1 U7365 ( .A(n5888), .ZN(n7422) );
  NAND2_X1 U7366 ( .A1(n6511), .A2(n7777), .ZN(n5897) );
  OAI21_X1 U7367 ( .B1(P1_IR_REG_13__SCAN_IN), .B2(P1_IR_REG_12__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5890) );
  AND2_X1 U7368 ( .A1(n5891), .A2(n5890), .ZN(n5893) );
  INV_X1 U7369 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U7370 ( .A1(n5893), .A2(n5892), .ZN(n5908) );
  INV_X1 U7371 ( .A(n5893), .ZN(n5894) );
  NAND2_X1 U7372 ( .A1(n5894), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5895) );
  AOI22_X1 U7373 ( .A1(n5664), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5635), .B2(
        n9624), .ZN(n5896) );
  NAND2_X1 U7374 ( .A1(n9421), .A2(n9002), .ZN(n5906) );
  NAND2_X1 U7375 ( .A1(n6148), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5904) );
  AND2_X1 U7376 ( .A1(n5898), .A2(n7625), .ZN(n5899) );
  NOR2_X1 U7377 ( .A1(n5912), .A2(n5899), .ZN(n7628) );
  NAND2_X1 U7378 ( .A1(n7783), .A2(n7628), .ZN(n5903) );
  INV_X1 U7379 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n5900) );
  OR2_X1 U7380 ( .A1(n6098), .A2(n5900), .ZN(n5902) );
  NAND2_X1 U7381 ( .A1(n7723), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5901) );
  NAND4_X1 U7382 ( .A1(n5904), .A2(n5903), .A3(n5902), .A4(n5901), .ZN(n9117)
         );
  NAND2_X1 U7383 ( .A1(n9117), .A2(n8995), .ZN(n5905) );
  NAND2_X1 U7384 ( .A1(n5906), .A2(n5905), .ZN(n5907) );
  XNOR2_X1 U7385 ( .A(n5907), .B(n8999), .ZN(n5923) );
  NAND2_X1 U7386 ( .A1(n6539), .A2(n7777), .ZN(n5911) );
  NAND2_X1 U7387 ( .A1(n5908), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5909) );
  XNOR2_X1 U7388 ( .A(n5909), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9635) );
  AOI22_X1 U7389 ( .A1(n5664), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5635), .B2(
        n9635), .ZN(n5910) );
  NAND2_X1 U7390 ( .A1(n7669), .A2(n9002), .ZN(n5920) );
  NAND2_X1 U7391 ( .A1(n6148), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5918) );
  NOR2_X1 U7392 ( .A1(n5912), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5913) );
  OR2_X1 U7393 ( .A1(n5939), .A2(n5913), .ZN(n7664) );
  INV_X1 U7394 ( .A(n7664), .ZN(n5914) );
  NAND2_X1 U7395 ( .A1(n7783), .A2(n5914), .ZN(n5917) );
  INV_X1 U7396 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7583) );
  OR2_X1 U7397 ( .A1(n6098), .A2(n7583), .ZN(n5916) );
  NAND2_X1 U7398 ( .A1(n7723), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5915) );
  NAND4_X1 U7399 ( .A1(n5918), .A2(n5917), .A3(n5916), .A4(n5915), .ZN(n9116)
         );
  NAND2_X1 U7400 ( .A1(n9116), .A2(n9001), .ZN(n5919) );
  NAND2_X1 U7401 ( .A1(n5920), .A2(n5919), .ZN(n5921) );
  XNOR2_X1 U7402 ( .A(n5921), .B(n6105), .ZN(n5931) );
  AND2_X1 U7403 ( .A1(n7619), .A2(n5931), .ZN(n5928) );
  INV_X1 U7404 ( .A(n5922), .ZN(n5925) );
  NAND2_X1 U7405 ( .A1(n9421), .A2(n8995), .ZN(n5927) );
  NAND2_X1 U7406 ( .A1(n9117), .A2(n8996), .ZN(n5926) );
  NAND2_X1 U7407 ( .A1(n5927), .A2(n5926), .ZN(n7618) );
  NAND2_X1 U7408 ( .A1(n5928), .A2(n7623), .ZN(n7660) );
  NAND2_X1 U7409 ( .A1(n7669), .A2(n8995), .ZN(n5930) );
  NAND2_X1 U7410 ( .A1(n9116), .A2(n8996), .ZN(n5929) );
  NAND2_X1 U7411 ( .A1(n5930), .A2(n5929), .ZN(n7659) );
  NAND2_X1 U7412 ( .A1(n7623), .A2(n7619), .ZN(n5933) );
  INV_X1 U7413 ( .A(n5931), .ZN(n5932) );
  NAND2_X1 U7414 ( .A1(n6541), .A2(n7777), .ZN(n5938) );
  OR2_X1 U7415 ( .A1(n5935), .A2(n5934), .ZN(n5936) );
  XNOR2_X1 U7416 ( .A(n5936), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7462) );
  AOI22_X1 U7417 ( .A1(n5664), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5635), .B2(
        n7462), .ZN(n5937) );
  NAND2_X1 U7418 ( .A1(n9410), .A2(n9002), .ZN(n5947) );
  NAND2_X1 U7419 ( .A1(n6148), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5945) );
  OR2_X1 U7420 ( .A1(n5939), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5940) );
  AND2_X1 U7421 ( .A1(n5954), .A2(n5940), .ZN(n7687) );
  NAND2_X1 U7422 ( .A1(n7783), .A2(n7687), .ZN(n5944) );
  NAND2_X1 U7423 ( .A1(n7723), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5943) );
  INV_X1 U7424 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n5941) );
  OR2_X1 U7425 ( .A1(n6098), .A2(n5941), .ZN(n5942) );
  NAND4_X1 U7426 ( .A1(n5945), .A2(n5944), .A3(n5943), .A4(n5942), .ZN(n9115)
         );
  NAND2_X1 U7427 ( .A1(n9115), .A2(n8995), .ZN(n5946) );
  NAND2_X1 U7428 ( .A1(n5947), .A2(n5946), .ZN(n5948) );
  XNOR2_X1 U7429 ( .A(n5948), .B(n8999), .ZN(n7683) );
  NAND2_X1 U7430 ( .A1(n9410), .A2(n8995), .ZN(n5950) );
  NAND2_X1 U7431 ( .A1(n9115), .A2(n8996), .ZN(n5949) );
  NAND2_X1 U7432 ( .A1(n5950), .A2(n5949), .ZN(n7684) );
  NAND2_X1 U7433 ( .A1(n6566), .A2(n7777), .ZN(n5953) );
  NAND2_X1 U7434 ( .A1(n5951), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5968) );
  XNOR2_X1 U7435 ( .A(n5968), .B(P1_IR_REG_17__SCAN_IN), .ZN(n7460) );
  AOI22_X1 U7436 ( .A1(n5664), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5635), .B2(
        n7460), .ZN(n5952) );
  NAND2_X1 U7437 ( .A1(n9405), .A2(n9002), .ZN(n5962) );
  NAND2_X1 U7438 ( .A1(n6148), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5960) );
  NAND2_X1 U7439 ( .A1(n5954), .A2(n9047), .ZN(n5955) );
  AND2_X1 U7440 ( .A1(n5974), .A2(n5955), .ZN(n9323) );
  NAND2_X1 U7441 ( .A1(n7783), .A2(n9323), .ZN(n5959) );
  INV_X1 U7442 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n5956) );
  OR2_X1 U7443 ( .A1(n6098), .A2(n5956), .ZN(n5958) );
  NAND2_X1 U7444 ( .A1(n7723), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5957) );
  NAND4_X1 U7445 ( .A1(n5960), .A2(n5959), .A3(n5958), .A4(n5957), .ZN(n9301)
         );
  NAND2_X1 U7446 ( .A1(n9301), .A2(n9001), .ZN(n5961) );
  NAND2_X1 U7447 ( .A1(n5962), .A2(n5961), .ZN(n5963) );
  XNOR2_X1 U7448 ( .A(n5963), .B(n6105), .ZN(n5966) );
  AND2_X1 U7449 ( .A1(n9301), .A2(n8996), .ZN(n5964) );
  AOI21_X1 U7450 ( .B1(n9405), .B2(n9001), .A(n5964), .ZN(n5965) );
  XNOR2_X1 U7451 ( .A(n5966), .B(n5965), .ZN(n9046) );
  NAND2_X1 U7452 ( .A1(n6674), .A2(n7777), .ZN(n5972) );
  INV_X1 U7453 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5967) );
  NAND2_X1 U7454 ( .A1(n5968), .A2(n5967), .ZN(n5969) );
  NAND2_X1 U7455 ( .A1(n5969), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5970) );
  XNOR2_X1 U7456 ( .A(n5970), .B(P1_IR_REG_18__SCAN_IN), .ZN(n7472) );
  AOI22_X1 U7457 ( .A1(n5664), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5635), .B2(
        n7472), .ZN(n5971) );
  NAND2_X1 U7458 ( .A1(n9397), .A2(n9002), .ZN(n5981) );
  AND2_X1 U7459 ( .A1(n5974), .A2(n5973), .ZN(n5975) );
  OR2_X1 U7460 ( .A1(n5975), .A2(n6005), .ZN(n9306) );
  INV_X1 U7461 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9129) );
  INV_X1 U7462 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9307) );
  OR2_X1 U7463 ( .A1(n6098), .A2(n9307), .ZN(n5976) );
  OAI21_X1 U7464 ( .B1(n6049), .B2(n9129), .A(n5976), .ZN(n5977) );
  INV_X1 U7465 ( .A(n5977), .ZN(n5979) );
  NAND2_X1 U7466 ( .A1(n7723), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5978) );
  OAI211_X1 U7467 ( .C1(n6038), .C2(n9306), .A(n5979), .B(n5978), .ZN(n9114)
         );
  NAND2_X1 U7468 ( .A1(n9114), .A2(n8995), .ZN(n5980) );
  NAND2_X1 U7469 ( .A1(n5981), .A2(n5980), .ZN(n5982) );
  XNOR2_X1 U7470 ( .A(n5982), .B(n8999), .ZN(n5985) );
  NAND2_X1 U7471 ( .A1(n5984), .A2(n5985), .ZN(n9085) );
  AND2_X1 U7472 ( .A1(n9114), .A2(n8996), .ZN(n5983) );
  AOI21_X1 U7473 ( .B1(n9397), .B2(n8995), .A(n5983), .ZN(n9083) );
  INV_X1 U7474 ( .A(n5985), .ZN(n5986) );
  NAND2_X1 U7475 ( .A1(n4729), .A2(n5986), .ZN(n9084) );
  NAND2_X1 U7476 ( .A1(n6807), .A2(n7777), .ZN(n5988) );
  AOI22_X1 U7477 ( .A1(n5664), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9721), .B2(
        n5635), .ZN(n5987) );
  NAND2_X1 U7478 ( .A1(n9391), .A2(n9002), .ZN(n5997) );
  INV_X1 U7479 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n8817) );
  NAND2_X1 U7480 ( .A1(n6148), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7481 ( .A1(n6153), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5989) );
  OAI211_X1 U7482 ( .C1(n5991), .C2(n8817), .A(n5990), .B(n5989), .ZN(n5992)
         );
  INV_X1 U7483 ( .A(n5992), .ZN(n5995) );
  INV_X1 U7484 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5993) );
  XNOR2_X1 U7485 ( .A(n6005), .B(n5993), .ZN(n9290) );
  NAND2_X1 U7486 ( .A1(n9290), .A2(n7783), .ZN(n5994) );
  NAND2_X1 U7487 ( .A1(n5995), .A2(n5994), .ZN(n9300) );
  NAND2_X1 U7488 ( .A1(n9300), .A2(n9001), .ZN(n5996) );
  NAND2_X1 U7489 ( .A1(n5997), .A2(n5996), .ZN(n5998) );
  XNOR2_X1 U7490 ( .A(n5998), .B(n8999), .ZN(n6001) );
  AOI22_X1 U7491 ( .A1(n9391), .A2(n8995), .B1(n8996), .B2(n9300), .ZN(n5999)
         );
  XNOR2_X1 U7492 ( .A(n6001), .B(n5999), .ZN(n8989) );
  INV_X1 U7493 ( .A(n5999), .ZN(n6000) );
  NAND2_X1 U7494 ( .A1(n7086), .A2(n7777), .ZN(n6004) );
  OR2_X1 U7495 ( .A1(n7779), .A2(n7703), .ZN(n6003) );
  NAND2_X1 U7496 ( .A1(n9385), .A2(n9002), .ZN(n6010) );
  AOI21_X1 U7497 ( .B1(n6005), .B2(P1_REG3_REG_19__SCAN_IN), .A(
        P1_REG3_REG_20__SCAN_IN), .ZN(n6006) );
  OR2_X1 U7498 ( .A1(n6020), .A2(n6006), .ZN(n9271) );
  AOI22_X1 U7499 ( .A1(n6148), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n6153), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n6008) );
  NAND2_X1 U7500 ( .A1(n7723), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6007) );
  OAI211_X1 U7501 ( .C1(n9271), .C2(n6038), .A(n6008), .B(n6007), .ZN(n9113)
         );
  NAND2_X1 U7502 ( .A1(n9113), .A2(n9001), .ZN(n6009) );
  NAND2_X1 U7503 ( .A1(n6010), .A2(n6009), .ZN(n6011) );
  XNOR2_X1 U7504 ( .A(n6011), .B(n8999), .ZN(n6014) );
  NAND2_X1 U7505 ( .A1(n9385), .A2(n9001), .ZN(n6013) );
  NAND2_X1 U7506 ( .A1(n9113), .A2(n8996), .ZN(n6012) );
  NAND2_X1 U7507 ( .A1(n6013), .A2(n6012), .ZN(n6015) );
  NAND2_X1 U7508 ( .A1(n6014), .A2(n6015), .ZN(n9063) );
  INV_X1 U7509 ( .A(n6014), .ZN(n6017) );
  INV_X1 U7510 ( .A(n6015), .ZN(n6016) );
  NAND2_X1 U7511 ( .A1(n6017), .A2(n6016), .ZN(n9065) );
  NAND2_X1 U7512 ( .A1(n7084), .A2(n7777), .ZN(n6019) );
  INV_X1 U7513 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8943) );
  OR2_X1 U7514 ( .A1(n5663), .A2(n8943), .ZN(n6018) );
  NOR2_X1 U7515 ( .A1(n6020), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6021) );
  OR2_X1 U7516 ( .A1(n6032), .A2(n6021), .ZN(n9261) );
  AOI22_X1 U7517 ( .A1(n6148), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n7723), .B2(
        P1_REG0_REG_21__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U7518 ( .A1(n6153), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6022) );
  OAI211_X1 U7519 ( .C1(n9261), .C2(n6038), .A(n6023), .B(n6022), .ZN(n9276)
         );
  AOI22_X1 U7520 ( .A1(n9382), .A2(n8995), .B1(n8996), .B2(n9276), .ZN(n6027)
         );
  NAND2_X1 U7521 ( .A1(n9382), .A2(n9002), .ZN(n6025) );
  NAND2_X1 U7522 ( .A1(n9276), .A2(n9001), .ZN(n6024) );
  NAND2_X1 U7523 ( .A1(n6025), .A2(n6024), .ZN(n6026) );
  XNOR2_X1 U7524 ( .A(n6026), .B(n8999), .ZN(n6029) );
  XOR2_X1 U7525 ( .A(n6027), .B(n6029), .Z(n9032) );
  INV_X1 U7526 ( .A(n6027), .ZN(n6028) );
  NAND2_X1 U7527 ( .A1(n7226), .A2(n7777), .ZN(n6031) );
  OR2_X1 U7528 ( .A1(n5663), .A2(n8948), .ZN(n6030) );
  NOR2_X1 U7529 ( .A1(n6032), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6033) );
  OR2_X1 U7530 ( .A1(n6044), .A2(n6033), .ZN(n9244) );
  INV_X1 U7531 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9245) );
  NAND2_X1 U7532 ( .A1(n6148), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U7533 ( .A1(n7723), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6034) );
  OAI211_X1 U7534 ( .C1(n6098), .C2(n9245), .A(n6035), .B(n6034), .ZN(n6036)
         );
  INV_X1 U7535 ( .A(n6036), .ZN(n6037) );
  OAI21_X1 U7536 ( .B1(n9244), .B2(n6038), .A(n6037), .ZN(n9112) );
  AOI22_X1 U7537 ( .A1(n9377), .A2(n9001), .B1(n8996), .B2(n9112), .ZN(n6040)
         );
  NAND2_X1 U7538 ( .A1(n6041), .A2(n6040), .ZN(n9072) );
  INV_X1 U7539 ( .A(n9377), .ZN(n9243) );
  INV_X1 U7540 ( .A(n9112), .ZN(n9258) );
  OAI22_X1 U7541 ( .A1(n9243), .A2(n5637), .B1(n9258), .B2(n6055), .ZN(n6039)
         );
  XNOR2_X1 U7542 ( .A(n6039), .B(n8999), .ZN(n9075) );
  NAND2_X1 U7543 ( .A1(n7261), .A2(n7777), .ZN(n6043) );
  OR2_X1 U7544 ( .A1(n5663), .A2(n7264), .ZN(n6042) );
  OR2_X1 U7545 ( .A1(n6044), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6046) );
  AND2_X1 U7546 ( .A1(n6046), .A2(n6045), .ZN(n9231) );
  NAND2_X1 U7547 ( .A1(n9231), .A2(n7783), .ZN(n6052) );
  INV_X1 U7548 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n8944) );
  NAND2_X1 U7549 ( .A1(n7723), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6048) );
  NAND2_X1 U7550 ( .A1(n6153), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6047) );
  OAI211_X1 U7551 ( .C1(n6049), .C2(n8944), .A(n6048), .B(n6047), .ZN(n6050)
         );
  INV_X1 U7552 ( .A(n6050), .ZN(n6051) );
  NAND2_X1 U7553 ( .A1(n6052), .A2(n6051), .ZN(n9222) );
  AOI22_X1 U7554 ( .A1(n9370), .A2(n9002), .B1(n8995), .B2(n9222), .ZN(n6053)
         );
  XNOR2_X1 U7555 ( .A(n6053), .B(n8999), .ZN(n6056) );
  NAND2_X1 U7556 ( .A1(n6057), .A2(n6056), .ZN(n8978) );
  INV_X1 U7557 ( .A(n8996), .ZN(n6054) );
  OAI22_X1 U7558 ( .A1(n9233), .A2(n6055), .B1(n9251), .B2(n6054), .ZN(n8980)
         );
  XOR2_X1 U7559 ( .A(n6059), .B(n6058), .Z(n9055) );
  NAND2_X1 U7560 ( .A1(n7535), .A2(n7777), .ZN(n6061) );
  OR2_X1 U7561 ( .A1(n5663), .A2(n7539), .ZN(n6060) );
  NAND2_X1 U7562 ( .A1(n9360), .A2(n9002), .ZN(n6069) );
  NAND2_X1 U7563 ( .A1(n5675), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6067) );
  NAND2_X1 U7564 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n6062), .ZN(n6078) );
  OAI21_X1 U7565 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n6062), .A(n6078), .ZN(
        n9041) );
  INV_X1 U7566 ( .A(n9041), .ZN(n9200) );
  NAND2_X1 U7567 ( .A1(n7783), .A2(n9200), .ZN(n6066) );
  INV_X1 U7568 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n6063) );
  OR2_X1 U7569 ( .A1(n6098), .A2(n6063), .ZN(n6065) );
  NAND2_X1 U7570 ( .A1(n7723), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6064) );
  NAND4_X1 U7571 ( .A1(n6067), .A2(n6066), .A3(n6065), .A4(n6064), .ZN(n9221)
         );
  NAND2_X1 U7572 ( .A1(n9221), .A2(n9001), .ZN(n6068) );
  NAND2_X1 U7573 ( .A1(n6069), .A2(n6068), .ZN(n6070) );
  XNOR2_X1 U7574 ( .A(n6070), .B(n8999), .ZN(n6071) );
  AOI22_X1 U7575 ( .A1(n9360), .A2(n8995), .B1(n8996), .B2(n9221), .ZN(n6072)
         );
  XNOR2_X1 U7576 ( .A(n6071), .B(n6072), .ZN(n9038) );
  INV_X1 U7577 ( .A(n6071), .ZN(n6073) );
  NAND2_X1 U7578 ( .A1(n7540), .A2(n7777), .ZN(n6075) );
  OR2_X1 U7579 ( .A1(n5663), .A2(n7557), .ZN(n6074) );
  NAND2_X1 U7580 ( .A1(n9355), .A2(n9002), .ZN(n6085) );
  NAND2_X1 U7581 ( .A1(n6148), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6083) );
  INV_X1 U7582 ( .A(n6078), .ZN(n6076) );
  NAND2_X1 U7583 ( .A1(n6076), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6095) );
  INV_X1 U7584 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6077) );
  NAND2_X1 U7585 ( .A1(n6078), .A2(n6077), .ZN(n6079) );
  AND2_X1 U7586 ( .A1(n6095), .A2(n6079), .ZN(n9187) );
  NAND2_X1 U7587 ( .A1(n7783), .A2(n9187), .ZN(n6082) );
  NAND2_X1 U7588 ( .A1(n6153), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6081) );
  NAND2_X1 U7589 ( .A1(n7723), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6080) );
  NAND4_X1 U7590 ( .A1(n6083), .A2(n6082), .A3(n6081), .A4(n6080), .ZN(n9207)
         );
  NAND2_X1 U7591 ( .A1(n9207), .A2(n9001), .ZN(n6084) );
  NAND2_X1 U7592 ( .A1(n6085), .A2(n6084), .ZN(n6086) );
  XNOR2_X1 U7593 ( .A(n6086), .B(n6105), .ZN(n6089) );
  AND2_X1 U7594 ( .A1(n9207), .A2(n8996), .ZN(n6087) );
  AOI21_X1 U7595 ( .B1(n9355), .B2(n8995), .A(n6087), .ZN(n6088) );
  NOR2_X1 U7596 ( .A1(n6089), .A2(n6088), .ZN(n9096) );
  NAND2_X1 U7597 ( .A1(n7592), .A2(n7777), .ZN(n6092) );
  OR2_X1 U7598 ( .A1(n5663), .A2(n6090), .ZN(n6091) );
  NAND2_X1 U7599 ( .A1(n9351), .A2(n9002), .ZN(n6104) );
  NAND2_X1 U7600 ( .A1(n5675), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6102) );
  INV_X1 U7601 ( .A(n6095), .ZN(n6093) );
  NAND2_X1 U7602 ( .A1(n6093), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6151) );
  INV_X1 U7603 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6094) );
  NAND2_X1 U7604 ( .A1(n6095), .A2(n6094), .ZN(n6096) );
  NAND2_X1 U7605 ( .A1(n7783), .A2(n9172), .ZN(n6101) );
  NAND2_X1 U7606 ( .A1(n7723), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6100) );
  INV_X1 U7607 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n6097) );
  OR2_X1 U7608 ( .A1(n6098), .A2(n6097), .ZN(n6099) );
  NAND4_X1 U7609 ( .A1(n6102), .A2(n6101), .A3(n6100), .A4(n6099), .ZN(n9191)
         );
  NAND2_X1 U7610 ( .A1(n9191), .A2(n8995), .ZN(n6103) );
  NAND2_X1 U7611 ( .A1(n6104), .A2(n6103), .ZN(n6106) );
  XNOR2_X1 U7612 ( .A(n6106), .B(n6105), .ZN(n6109) );
  INV_X1 U7613 ( .A(n6109), .ZN(n6111) );
  AND2_X1 U7614 ( .A1(n9191), .A2(n8996), .ZN(n6107) );
  AOI21_X1 U7615 ( .B1(n9351), .B2(n9001), .A(n6107), .ZN(n6108) );
  INV_X1 U7616 ( .A(n6108), .ZN(n6110) );
  AOI21_X1 U7617 ( .B1(n6111), .B2(n6110), .A(n9014), .ZN(n6113) );
  NAND2_X1 U7618 ( .A1(n7358), .A2(P1_B_REG_SCAN_IN), .ZN(n6114) );
  OAI22_X1 U7619 ( .A1(n6127), .A2(n6114), .B1(P1_B_REG_SCAN_IN), .B2(n7358), 
        .ZN(n6115) );
  OR2_X1 U7620 ( .A1(n6115), .A2(n7559), .ZN(n6475) );
  NOR4_X1 U7621 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6119) );
  NOR4_X1 U7622 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6118) );
  NOR4_X1 U7623 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6117) );
  NOR4_X1 U7624 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6116) );
  AND4_X1 U7625 ( .A1(n6119), .A2(n6118), .A3(n6117), .A4(n6116), .ZN(n6125)
         );
  NOR2_X1 U7626 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .ZN(
        n6123) );
  NOR4_X1 U7627 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6122) );
  NOR4_X1 U7628 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n6121) );
  NOR4_X1 U7629 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n6120) );
  AND4_X1 U7630 ( .A1(n6123), .A2(n6122), .A3(n6121), .A4(n6120), .ZN(n6124)
         );
  NAND2_X1 U7631 ( .A1(n6125), .A2(n6124), .ZN(n6472) );
  INV_X1 U7632 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6312) );
  NOR2_X1 U7633 ( .A1(n6472), .A2(n6312), .ZN(n6126) );
  NAND2_X1 U7634 ( .A1(n7559), .A2(n7358), .ZN(n6474) );
  OAI21_X1 U7635 ( .B1(n6475), .B2(n6126), .A(n6474), .ZN(n6428) );
  INV_X1 U7636 ( .A(n6127), .ZN(n7537) );
  NAND2_X1 U7637 ( .A1(n7559), .A2(n7537), .ZN(n6313) );
  OAI21_X1 U7638 ( .B1(n6475), .B2(P1_D_REG_1__SCAN_IN), .A(n6313), .ZN(n6719)
         );
  OR2_X1 U7639 ( .A1(n6428), .A2(n6719), .ZN(n6143) );
  NAND2_X1 U7640 ( .A1(n6128), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6129) );
  MUX2_X1 U7641 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6129), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n6130) );
  NAND2_X1 U7642 ( .A1(n6130), .A2(n5578), .ZN(n7262) );
  AND2_X1 U7643 ( .A1(n7262), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6131) );
  NOR2_X1 U7644 ( .A1(n6143), .A2(n6722), .ZN(n6145) );
  NAND2_X1 U7645 ( .A1(n6135), .A2(n9086), .ZN(n6163) );
  NAND2_X1 U7646 ( .A1(n4342), .A2(n6143), .ZN(n6137) );
  OR2_X1 U7647 ( .A1(n7899), .A2(n7977), .ZN(n6136) );
  NAND2_X1 U7648 ( .A1(n6137), .A2(n6479), .ZN(n9026) );
  NAND2_X1 U7649 ( .A1(n9799), .A2(n6143), .ZN(n6434) );
  AND3_X1 U7650 ( .A1(n6136), .A2(n6165), .A3(n7262), .ZN(n6138) );
  NAND3_X1 U7651 ( .A1(n6434), .A2(n6138), .A3(n6137), .ZN(n6139) );
  INV_X1 U7652 ( .A(n9207), .ZN(n9178) );
  OR2_X1 U7653 ( .A1(n6724), .A2(n6723), .ZN(n7170) );
  OR2_X1 U7654 ( .A1(n6722), .A2(n6141), .ZN(n6142) );
  NOR2_X1 U7655 ( .A1(n7170), .A2(n6142), .ZN(n7982) );
  INV_X1 U7656 ( .A(n6143), .ZN(n6144) );
  NAND2_X1 U7657 ( .A1(n7982), .A2(n6144), .ZN(n9104) );
  AND2_X1 U7658 ( .A1(n6145), .A2(n6141), .ZN(n6147) );
  INV_X1 U7659 ( .A(n7170), .ZN(n6146) );
  AND2_X2 U7660 ( .A1(n6147), .A2(n6146), .ZN(n9101) );
  NAND2_X1 U7661 ( .A1(n6148), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6157) );
  INV_X1 U7662 ( .A(n6151), .ZN(n6149) );
  NAND2_X1 U7663 ( .A1(n6149), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n7782) );
  INV_X1 U7664 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6150) );
  NAND2_X1 U7665 ( .A1(n6151), .A2(n6150), .ZN(n6152) );
  NAND2_X1 U7666 ( .A1(n7783), .A2(n9158), .ZN(n6156) );
  NAND2_X1 U7667 ( .A1(n6153), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6155) );
  NAND2_X1 U7668 ( .A1(n7723), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6154) );
  NAND4_X1 U7669 ( .A1(n6157), .A2(n6156), .A3(n6155), .A4(n6154), .ZN(n9111)
         );
  INV_X2 U7670 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  AOI22_X1 U7671 ( .A1(n9101), .A2(n9111), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n6158) );
  OAI21_X1 U7672 ( .B1(n9178), .B2(n9104), .A(n6158), .ZN(n6159) );
  AOI21_X1 U7673 ( .B1(n9172), .B2(n9099), .A(n6159), .ZN(n6160) );
  INV_X1 U7674 ( .A(n6161), .ZN(n6162) );
  NAND2_X1 U7675 ( .A1(n6163), .A2(n6162), .ZN(P1_U3212) );
  INV_X1 U7676 ( .A(n7262), .ZN(n6164) );
  NOR2_X1 U7677 ( .A1(n6165), .A2(n6164), .ZN(n6371) );
  NAND2_X1 U7678 ( .A1(n7899), .A2(n6165), .ZN(n6166) );
  NAND2_X1 U7679 ( .A1(n6166), .A2(n7262), .ZN(n9551) );
  NAND2_X1 U7680 ( .A1(n9551), .A2(n6167), .ZN(n6168) );
  NAND2_X1 U7681 ( .A1(n6168), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U7682 ( .A(n6181), .ZN(n6169) );
  INV_X1 U7683 ( .A(n8125), .ZN(n6170) );
  AOI211_X1 U7684 ( .C1(n6172), .C2(n6171), .A(n9835), .B(n6170), .ZN(n6178)
         );
  INV_X1 U7685 ( .A(n8771), .ZN(n6173) );
  INV_X1 U7686 ( .A(n9854), .ZN(n8214) );
  NOR2_X1 U7687 ( .A1(n6173), .A2(n8214), .ZN(n6177) );
  OAI22_X1 U7688 ( .A1(n9860), .A2(n8663), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6174), .ZN(n6176) );
  INV_X1 U7689 ( .A(n8655), .ZN(n8350) );
  INV_X1 U7690 ( .A(n8657), .ZN(n8073) );
  OAI22_X1 U7691 ( .A1(n8350), .A2(n8219), .B1(n9831), .B2(n8073), .ZN(n6175)
         );
  OR4_X1 U7692 ( .A1(n6178), .A2(n6177), .A3(n6176), .A4(n6175), .ZN(P2_U3235)
         );
  NAND2_X1 U7693 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n6189) );
  XNOR2_X1 U7694 ( .A(n6212), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n6188) );
  INV_X1 U7695 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9867) );
  NOR3_X1 U7696 ( .A1(n6188), .A2(n9864), .A3(n9867), .ZN(n6204) );
  NAND2_X1 U7697 ( .A1(n9886), .A2(n6179), .ZN(n6184) );
  OR2_X1 U7698 ( .A1(n5534), .A2(n10007), .ZN(n7616) );
  OR2_X1 U7699 ( .A1(n6180), .A2(P2_U3152), .ZN(n8447) );
  OAI21_X1 U7700 ( .B1(n6181), .B2(n7616), .A(n8447), .ZN(n6182) );
  INV_X1 U7701 ( .A(n6182), .ZN(n6183) );
  NAND2_X1 U7702 ( .A1(n6184), .A2(n6183), .ZN(n6185) );
  NAND2_X1 U7703 ( .A1(n6185), .A2(n6195), .ZN(n6191) );
  NAND2_X1 U7704 ( .A1(n6191), .A2(n8466), .ZN(n6190) );
  INV_X1 U7705 ( .A(n8441), .ZN(n8082) );
  NAND2_X1 U7706 ( .A1(n6190), .A2(n8082), .ZN(n8500) );
  INV_X1 U7707 ( .A(n8500), .ZN(n6187) );
  INV_X1 U7708 ( .A(n9879), .ZN(n8490) );
  AOI211_X1 U7709 ( .C1(n6189), .C2(n6188), .A(n6204), .B(n8490), .ZN(n6203)
         );
  INV_X1 U7710 ( .A(n6212), .ZN(n6287) );
  NOR2_X1 U7711 ( .A1(n9861), .A2(n6287), .ZN(n6202) );
  NAND2_X1 U7712 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n6194) );
  XNOR2_X1 U7713 ( .A(n6212), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n6193) );
  INV_X1 U7714 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9945) );
  NOR3_X1 U7715 ( .A1(n6193), .A2(n9945), .A3(n9867), .ZN(n6211) );
  INV_X1 U7716 ( .A(n6191), .ZN(n6192) );
  AOI211_X1 U7717 ( .C1(n6194), .C2(n6193), .A(n6211), .B(n9862), .ZN(n6201)
         );
  NAND2_X1 U7718 ( .A1(n9886), .A2(n6581), .ZN(n6196) );
  NAND2_X1 U7719 ( .A1(n6196), .A2(n6195), .ZN(n6198) );
  INV_X1 U7720 ( .A(n8447), .ZN(n7258) );
  OR2_X1 U7721 ( .A1(n9886), .A2(n7258), .ZN(n6197) );
  NAND2_X1 U7722 ( .A1(n6198), .A2(n6197), .ZN(n8506) );
  INV_X1 U7723 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6199) );
  INV_X1 U7724 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6881) );
  OAI22_X1 U7725 ( .A1(n8506), .A2(n6199), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6881), .ZN(n6200) );
  OR4_X1 U7726 ( .A1(n6203), .A2(n6202), .A3(n6201), .A4(n6200), .ZN(P2_U3246)
         );
  INV_X1 U7727 ( .A(n6306), .ZN(n6216) );
  INV_X1 U7728 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6205) );
  MUX2_X1 U7729 ( .A(n6205), .B(P2_REG2_REG_2__SCAN_IN), .S(n6240), .Z(n6238)
         );
  XNOR2_X1 U7730 ( .A(n6253), .B(P2_REG2_REG_3__SCAN_IN), .ZN(n6251) );
  AOI21_X1 U7731 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(n6253), .A(n6250), .ZN(
        n6227) );
  INV_X1 U7732 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6206) );
  MUX2_X1 U7733 ( .A(n6206), .B(P2_REG2_REG_4__SCAN_IN), .S(n6228), .Z(n6226)
         );
  NOR2_X1 U7734 ( .A1(n6227), .A2(n6226), .ZN(n6225) );
  AOI21_X1 U7735 ( .B1(n6228), .B2(P2_REG2_REG_4__SCAN_IN), .A(n6225), .ZN(
        n6265) );
  XNOR2_X1 U7736 ( .A(n6266), .B(P2_REG2_REG_5__SCAN_IN), .ZN(n6264) );
  NOR2_X1 U7737 ( .A1(n6265), .A2(n6264), .ZN(n6263) );
  AOI21_X1 U7738 ( .B1(n6266), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6263), .ZN(
        n6278) );
  INV_X1 U7739 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6207) );
  MUX2_X1 U7740 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6207), .S(n6306), .Z(n6277)
         );
  NAND2_X1 U7741 ( .A1(n6631), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6208) );
  OAI21_X1 U7742 ( .B1(n6631), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6208), .ZN(
        n6209) );
  AOI211_X1 U7743 ( .C1(n6210), .C2(n6209), .A(n8490), .B(n6630), .ZN(n6224)
         );
  INV_X1 U7744 ( .A(n6631), .ZN(n6624) );
  NOR2_X1 U7745 ( .A1(n9861), .A2(n6624), .ZN(n6223) );
  AOI21_X1 U7746 ( .B1(n6212), .B2(P2_REG1_REG_1__SCAN_IN), .A(n6211), .ZN(
        n6243) );
  INV_X1 U7747 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6213) );
  MUX2_X1 U7748 ( .A(n6213), .B(P2_REG1_REG_2__SCAN_IN), .S(n6240), .Z(n6242)
         );
  NOR2_X1 U7749 ( .A1(n6243), .A2(n6242), .ZN(n6241) );
  AOI21_X1 U7750 ( .B1(n6240), .B2(P2_REG1_REG_2__SCAN_IN), .A(n6241), .ZN(
        n6256) );
  XNOR2_X1 U7751 ( .A(n6253), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n6255) );
  NOR2_X1 U7752 ( .A1(n6256), .A2(n6255), .ZN(n6254) );
  INV_X1 U7753 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6214) );
  MUX2_X1 U7754 ( .A(n6214), .B(P2_REG1_REG_4__SCAN_IN), .S(n6228), .Z(n6230)
         );
  NOR2_X1 U7755 ( .A1(n6231), .A2(n6230), .ZN(n6229) );
  AOI21_X1 U7756 ( .B1(n6228), .B2(P2_REG1_REG_4__SCAN_IN), .A(n6229), .ZN(
        n6269) );
  XNOR2_X1 U7757 ( .A(n6266), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n6268) );
  NOR2_X1 U7758 ( .A1(n6269), .A2(n6268), .ZN(n6267) );
  INV_X1 U7759 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6215) );
  MUX2_X1 U7760 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6215), .S(n6306), .Z(n6280)
         );
  NOR2_X1 U7761 ( .A1(n6281), .A2(n6280), .ZN(n6279) );
  AOI21_X1 U7762 ( .B1(n6216), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6279), .ZN(
        n6220) );
  NAND2_X1 U7763 ( .A1(n6631), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6217) );
  OAI21_X1 U7764 ( .B1(n6631), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6217), .ZN(
        n6219) );
  OR2_X1 U7765 ( .A1(n6220), .A2(n6219), .ZN(n6623) );
  INV_X1 U7766 ( .A(n6623), .ZN(n6218) );
  AOI211_X1 U7767 ( .C1(n6220), .C2(n6219), .A(n9862), .B(n6218), .ZN(n6222)
         );
  INV_X1 U7768 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n9999) );
  NAND2_X1 U7769 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6764) );
  OAI21_X1 U7770 ( .B1(n8506), .B2(n9999), .A(n6764), .ZN(n6221) );
  OR4_X1 U7771 ( .A1(n6224), .A2(n6223), .A3(n6222), .A4(n6221), .ZN(P2_U3252)
         );
  AOI211_X1 U7772 ( .C1(n6227), .C2(n6226), .A(n6225), .B(n8490), .ZN(n6236)
         );
  INV_X1 U7773 ( .A(n6228), .ZN(n6299) );
  NOR2_X1 U7774 ( .A1(n9861), .A2(n6299), .ZN(n6235) );
  AOI211_X1 U7775 ( .C1(n6231), .C2(n6230), .A(n6229), .B(n9862), .ZN(n6234)
         );
  INV_X1 U7776 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U7777 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(n10007), .ZN(n6853) );
  OAI21_X1 U7778 ( .B1(n8506), .B2(n6232), .A(n6853), .ZN(n6233) );
  OR4_X1 U7779 ( .A1(n6236), .A2(n6235), .A3(n6234), .A4(n6233), .ZN(P2_U3249)
         );
  AOI211_X1 U7780 ( .C1(n6239), .C2(n6238), .A(n6237), .B(n8490), .ZN(n6249)
         );
  INV_X1 U7781 ( .A(n6240), .ZN(n6289) );
  NOR2_X1 U7782 ( .A1(n9861), .A2(n6289), .ZN(n6248) );
  AOI211_X1 U7783 ( .C1(n6243), .C2(n6242), .A(n6241), .B(n9862), .ZN(n6247)
         );
  INV_X1 U7784 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6245) );
  INV_X1 U7785 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6244) );
  OAI22_X1 U7786 ( .A1(n8506), .A2(n6245), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6244), .ZN(n6246) );
  OR4_X1 U7787 ( .A1(n6249), .A2(n6248), .A3(n6247), .A4(n6246), .ZN(P2_U3247)
         );
  AOI211_X1 U7788 ( .C1(n6252), .C2(n6251), .A(n6250), .B(n8490), .ZN(n6262)
         );
  INV_X1 U7789 ( .A(n6253), .ZN(n6291) );
  NOR2_X1 U7790 ( .A1(n9861), .A2(n6291), .ZN(n6261) );
  AOI211_X1 U7791 ( .C1(n6256), .C2(n6255), .A(n6254), .B(n9862), .ZN(n6260)
         );
  INV_X1 U7792 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6258) );
  NAND2_X1 U7793 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3152), .ZN(n6257) );
  OAI21_X1 U7794 ( .B1(n8506), .B2(n6258), .A(n6257), .ZN(n6259) );
  OR4_X1 U7795 ( .A1(n6262), .A2(n6261), .A3(n6260), .A4(n6259), .ZN(P2_U3248)
         );
  AOI211_X1 U7796 ( .C1(n6265), .C2(n6264), .A(n6263), .B(n8490), .ZN(n6275)
         );
  INV_X1 U7797 ( .A(n6266), .ZN(n6303) );
  NOR2_X1 U7798 ( .A1(n9861), .A2(n6303), .ZN(n6274) );
  AOI211_X1 U7799 ( .C1(n6269), .C2(n6268), .A(n6267), .B(n9862), .ZN(n6273)
         );
  INV_X1 U7800 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6271) );
  NAND2_X1 U7801 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(n10007), .ZN(n6270) );
  OAI21_X1 U7802 ( .B1(n8506), .B2(n6271), .A(n6270), .ZN(n6272) );
  OR4_X1 U7803 ( .A1(n6275), .A2(n6274), .A3(n6273), .A4(n6272), .ZN(P2_U3250)
         );
  AOI211_X1 U7804 ( .C1(n6278), .C2(n6277), .A(n8490), .B(n6276), .ZN(n6286)
         );
  AOI211_X1 U7805 ( .C1(n6281), .C2(n6280), .A(n9862), .B(n6279), .ZN(n6285)
         );
  NOR2_X1 U7806 ( .A1(n9861), .A2(n6306), .ZN(n6284) );
  INV_X1 U7807 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n9985) );
  NAND2_X1 U7808 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(n10007), .ZN(n6282) );
  OAI21_X1 U7809 ( .B1(n8506), .B2(n9985), .A(n6282), .ZN(n6283) );
  OR4_X1 U7810 ( .A1(n6286), .A2(n6285), .A3(n6284), .A4(n6283), .ZN(P2_U3251)
         );
  NOR2_X1 U7811 ( .A1(n7715), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8967) );
  INV_X1 U7812 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6288) );
  NAND2_X1 U7813 ( .A1(n7715), .A2(n10007), .ZN(n8975) );
  CLKBUF_X1 U7814 ( .A(n8975), .Z(n8969) );
  OAI222_X1 U7815 ( .A1(n8971), .A2(n6288), .B1(n8969), .B2(n6292), .C1(n10007), .C2(n6287), .ZN(P2_U3357) );
  OAI222_X1 U7816 ( .A1(n8971), .A2(n6290), .B1(n8969), .B2(n6294), .C1(
        P2_U3152), .C2(n6289), .ZN(P2_U3356) );
  OAI222_X1 U7817 ( .A1(n8971), .A2(n8933), .B1(n8969), .B2(n6296), .C1(n10007), .C2(n6291), .ZN(P2_U3355) );
  NAND2_X1 U7818 ( .A1(n7715), .A2(P1_U3084), .ZN(n8045) );
  NOR2_X1 U7819 ( .A1(n7715), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9447) );
  INV_X2 U7820 ( .A(n9447), .ZN(n8048) );
  OAI222_X1 U7821 ( .A1(n8045), .A2(n6293), .B1(n8048), .B2(n6292), .C1(
        P1_U3084), .C2(n9560), .ZN(P1_U3352) );
  INV_X1 U7822 ( .A(n8045), .ZN(n7594) );
  INV_X1 U7823 ( .A(n7594), .ZN(n9444) );
  OAI222_X1 U7824 ( .A1(n9444), .A2(n6295), .B1(n8048), .B2(n6294), .C1(
        P1_U3084), .C2(n9576), .ZN(P1_U3351) );
  OAI222_X1 U7825 ( .A1(n9444), .A2(n6297), .B1(n8048), .B2(n6296), .C1(
        P1_U3084), .C2(n6412), .ZN(P1_U3350) );
  OAI222_X1 U7826 ( .A1(n9444), .A2(n6298), .B1(n8048), .B2(n6300), .C1(
        P1_U3084), .C2(n6364), .ZN(P1_U3349) );
  OAI222_X1 U7827 ( .A1(n8971), .A2(n6301), .B1(n8969), .B2(n6300), .C1(
        P2_U3152), .C2(n6299), .ZN(P2_U3354) );
  OAI222_X1 U7828 ( .A1(n9444), .A2(n6302), .B1(n8048), .B2(n6304), .C1(
        P1_U3084), .C2(n6459), .ZN(P1_U3348) );
  OAI222_X1 U7829 ( .A1(n8971), .A2(n6305), .B1(n8969), .B2(n6304), .C1(n10007), .C2(n6303), .ZN(P2_U3353) );
  OAI222_X1 U7830 ( .A1(n8971), .A2(n6307), .B1(n8969), .B2(n6308), .C1(
        P2_U3152), .C2(n6306), .ZN(P2_U3352) );
  OAI222_X1 U7831 ( .A1(n9444), .A2(n6309), .B1(n8048), .B2(n6308), .C1(
        P1_U3084), .C2(n6366), .ZN(P1_U3347) );
  INV_X1 U7832 ( .A(n6474), .ZN(n6310) );
  AOI22_X1 U7833 ( .A1(n9744), .A2(n6312), .B1(n6311), .B2(n6310), .ZN(
        P1_U3440) );
  INV_X1 U7834 ( .A(n9744), .ZN(n9743) );
  OAI22_X1 U7835 ( .A1(n9743), .A2(P1_D_REG_1__SCAN_IN), .B1(n6722), .B2(n6313), .ZN(n6314) );
  INV_X1 U7836 ( .A(n6314), .ZN(P1_U3441) );
  INV_X1 U7837 ( .A(n6315), .ZN(n6316) );
  OAI222_X1 U7838 ( .A1(n8971), .A2(n4361), .B1(n8969), .B2(n6316), .C1(n10007), .C2(n6624), .ZN(P2_U3351) );
  OAI222_X1 U7839 ( .A1(n9444), .A2(n6317), .B1(n8048), .B2(n6316), .C1(
        P1_U3084), .C2(n6394), .ZN(P1_U3346) );
  INV_X1 U7840 ( .A(n6318), .ZN(n6320) );
  INV_X1 U7841 ( .A(n6645), .ZN(n6638) );
  OAI222_X1 U7842 ( .A1(n8971), .A2(n6319), .B1(n8969), .B2(n6320), .C1(
        P2_U3152), .C2(n6638), .ZN(P2_U3350) );
  INV_X1 U7843 ( .A(n6447), .ZN(n6399) );
  OAI222_X1 U7844 ( .A1(n9444), .A2(n6321), .B1(n8048), .B2(n6320), .C1(
        P1_U3084), .C2(n6399), .ZN(P1_U3345) );
  INV_X1 U7845 ( .A(n6322), .ZN(n6324) );
  AOI22_X1 U7846 ( .A1(n6666), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n8967), .ZN(n6323) );
  OAI21_X1 U7847 ( .B1(n6324), .B2(n8969), .A(n6323), .ZN(P2_U3349) );
  INV_X1 U7848 ( .A(n9610), .ZN(n6452) );
  OAI222_X1 U7849 ( .A1(P1_U3084), .A2(n6452), .B1(n8048), .B2(n6324), .C1(
        n8890), .C2(n8045), .ZN(P1_U3344) );
  INV_X1 U7850 ( .A(n6325), .ZN(n6335) );
  AOI22_X1 U7851 ( .A1(n6694), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n8967), .ZN(n6326) );
  OAI21_X1 U7852 ( .B1(n6335), .B2(n8975), .A(n6326), .ZN(P2_U3348) );
  INV_X1 U7853 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6334) );
  NAND2_X1 U7854 ( .A1(n6327), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6332) );
  NAND2_X1 U7855 ( .A1(n6328), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6331) );
  NAND2_X1 U7856 ( .A1(n6329), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6330) );
  NAND3_X1 U7857 ( .A1(n6332), .A2(n6331), .A3(n6330), .ZN(n8508) );
  NAND2_X1 U7858 ( .A1(n8508), .A2(P2_U3966), .ZN(n6333) );
  OAI21_X1 U7859 ( .B1(n6334), .B2(P2_U3966), .A(n6333), .ZN(P2_U3583) );
  INV_X1 U7860 ( .A(n6485), .ZN(n6491) );
  OAI222_X1 U7861 ( .A1(n8045), .A2(n6336), .B1(n8048), .B2(n6335), .C1(n6491), 
        .C2(P1_U3084), .ZN(P1_U3343) );
  INV_X1 U7862 ( .A(n6337), .ZN(n6340) );
  INV_X1 U7863 ( .A(n6791), .ZN(n6700) );
  OAI222_X1 U7864 ( .A1(n8969), .A2(n6340), .B1(n6700), .B2(n10007), .C1(n6338), .C2(n8971), .ZN(P2_U3347) );
  INV_X1 U7865 ( .A(n6492), .ZN(n6517) );
  OAI222_X1 U7866 ( .A1(P1_U3084), .A2(n6517), .B1(n8048), .B2(n6340), .C1(
        n6339), .C2(n9444), .ZN(P1_U3342) );
  NOR2_X1 U7867 ( .A1(n9870), .A2(P2_U3966), .ZN(P2_U3151) );
  MUX2_X1 U7868 ( .A(n6341), .B(P1_REG2_REG_2__SCAN_IN), .S(n9576), .Z(n9586)
         );
  INV_X1 U7869 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6342) );
  MUX2_X1 U7870 ( .A(n6342), .B(P1_REG2_REG_1__SCAN_IN), .S(n9560), .Z(n9565)
         );
  AND2_X1 U7871 ( .A1(n9556), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9566) );
  NAND2_X1 U7872 ( .A1(n9565), .A2(n9566), .ZN(n9564) );
  NAND2_X1 U7873 ( .A1(n5634), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6343) );
  NAND2_X1 U7874 ( .A1(n9564), .A2(n6343), .ZN(n9587) );
  NAND2_X1 U7875 ( .A1(n9586), .A2(n9587), .ZN(n9585) );
  OR2_X1 U7876 ( .A1(n9576), .A2(n6341), .ZN(n6413) );
  NAND2_X1 U7877 ( .A1(n9585), .A2(n6413), .ZN(n6346) );
  INV_X1 U7878 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6344) );
  MUX2_X1 U7879 ( .A(n6344), .B(P1_REG2_REG_3__SCAN_IN), .S(n6412), .Z(n6345)
         );
  NAND2_X1 U7880 ( .A1(n6346), .A2(n6345), .ZN(n6416) );
  INV_X1 U7881 ( .A(n6412), .ZN(n6362) );
  NAND2_X1 U7882 ( .A1(n6362), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6347) );
  AND2_X1 U7883 ( .A1(n6416), .A2(n6347), .ZN(n9593) );
  INV_X1 U7884 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6348) );
  MUX2_X1 U7885 ( .A(n6348), .B(P1_REG2_REG_4__SCAN_IN), .S(n6364), .Z(n9592)
         );
  NAND2_X1 U7886 ( .A1(n9593), .A2(n9592), .ZN(n9591) );
  NAND2_X1 U7887 ( .A1(n6364), .A2(n6348), .ZN(n6466) );
  INV_X1 U7888 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6349) );
  NAND2_X1 U7889 ( .A1(n6459), .A2(n6349), .ZN(n6350) );
  OAI21_X1 U7890 ( .B1(n6459), .B2(n6349), .A(n6350), .ZN(n6465) );
  AOI21_X1 U7891 ( .B1(n9591), .B2(n6466), .A(n6465), .ZN(n6468) );
  INV_X1 U7892 ( .A(n6468), .ZN(n6351) );
  NAND2_X1 U7893 ( .A1(n6351), .A2(n6350), .ZN(n6376) );
  MUX2_X1 U7894 ( .A(n5736), .B(P1_REG2_REG_6__SCAN_IN), .S(n6383), .Z(n6375)
         );
  OR2_X1 U7895 ( .A1(n6376), .A2(n6375), .ZN(n6352) );
  OAI21_X1 U7896 ( .B1(n5736), .B2(n6366), .A(n6352), .ZN(n6354) );
  AOI22_X1 U7897 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6394), .B1(n6387), .B2(
        n7177), .ZN(n6353) );
  NOR2_X1 U7898 ( .A1(n6353), .A2(n6354), .ZN(n6388) );
  AOI21_X1 U7899 ( .B1(n6354), .B2(n6353), .A(n6388), .ZN(n6374) );
  NOR2_X1 U7900 ( .A1(n9546), .A2(P1_U3084), .ZN(n7593) );
  NAND2_X1 U7901 ( .A1(n9551), .A2(n7593), .ZN(n9553) );
  INV_X1 U7902 ( .A(n6141), .ZN(n6423) );
  AND2_X1 U7903 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6868) );
  OR2_X1 U7904 ( .A1(n6141), .A2(P1_U3084), .ZN(n9549) );
  INV_X1 U7905 ( .A(n9546), .ZN(n9577) );
  NOR2_X1 U7906 ( .A1(n9549), .A2(n9577), .ZN(n6355) );
  MUX2_X1 U7907 ( .A(n9820), .B(P1_REG1_REG_7__SCAN_IN), .S(n6387), .Z(n6368)
         );
  INV_X1 U7908 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9818) );
  INV_X1 U7909 ( .A(n6364), .ZN(n9594) );
  INV_X1 U7910 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6356) );
  MUX2_X1 U7911 ( .A(n6356), .B(P1_REG1_REG_1__SCAN_IN), .S(n9560), .Z(n9562)
         );
  AND2_X1 U7912 ( .A1(n9556), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9563) );
  NAND2_X1 U7913 ( .A1(n9562), .A2(n9563), .ZN(n9571) );
  OR2_X1 U7914 ( .A1(n9560), .A2(n6356), .ZN(n9570) );
  NAND2_X1 U7915 ( .A1(n9571), .A2(n9570), .ZN(n6358) );
  MUX2_X1 U7916 ( .A(n9811), .B(P1_REG1_REG_2__SCAN_IN), .S(n9576), .Z(n6357)
         );
  NAND2_X1 U7917 ( .A1(n6358), .A2(n6357), .ZN(n9574) );
  INV_X1 U7918 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9811) );
  OR2_X1 U7919 ( .A1(n9576), .A2(n9811), .ZN(n6405) );
  NAND2_X1 U7920 ( .A1(n9574), .A2(n6405), .ZN(n6361) );
  INV_X1 U7921 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6359) );
  MUX2_X1 U7922 ( .A(n6359), .B(P1_REG1_REG_3__SCAN_IN), .S(n6412), .Z(n6360)
         );
  NAND2_X1 U7923 ( .A1(n6361), .A2(n6360), .ZN(n6408) );
  NAND2_X1 U7924 ( .A1(n6362), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6363) );
  AND2_X1 U7925 ( .A1(n6408), .A2(n6363), .ZN(n9597) );
  INV_X1 U7926 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9814) );
  MUX2_X1 U7927 ( .A(n9814), .B(P1_REG1_REG_4__SCAN_IN), .S(n6364), .Z(n9598)
         );
  NAND2_X1 U7928 ( .A1(n9597), .A2(n9598), .ZN(n9596) );
  OAI21_X1 U7929 ( .B1(n9594), .B2(P1_REG1_REG_4__SCAN_IN), .A(n9596), .ZN(
        n6462) );
  INV_X1 U7930 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9816) );
  MUX2_X1 U7931 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n9816), .S(n6459), .Z(n6461)
         );
  INV_X1 U7932 ( .A(n6460), .ZN(n6365) );
  OAI21_X1 U7933 ( .B1(n9816), .B2(n6459), .A(n6365), .ZN(n6380) );
  AOI22_X1 U7934 ( .A1(n6383), .A2(n9818), .B1(P1_REG1_REG_6__SCAN_IN), .B2(
        n6366), .ZN(n6379) );
  NOR2_X1 U7935 ( .A1(n6380), .A2(n6379), .ZN(n6378) );
  NOR2_X1 U7936 ( .A1(n6367), .A2(n6368), .ZN(n6393) );
  AOI21_X1 U7937 ( .B1(n6368), .B2(n6367), .A(n6393), .ZN(n6369) );
  NOR2_X1 U7938 ( .A1(n9621), .A2(n6369), .ZN(n6370) );
  AOI211_X1 U7939 ( .C1(n9636), .C2(n6387), .A(n6868), .B(n6370), .ZN(n6373)
         );
  OR2_X1 U7940 ( .A1(P1_U3083), .A2(n6371), .ZN(n9632) );
  NAND2_X1 U7941 ( .A1(n9661), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n6372) );
  OAI211_X1 U7942 ( .C1(n6374), .C2(n9627), .A(n6373), .B(n6372), .ZN(P1_U3248) );
  XNOR2_X1 U7943 ( .A(n6376), .B(n6375), .ZN(n6386) );
  INV_X1 U7944 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6377) );
  NOR2_X1 U7945 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6377), .ZN(n6813) );
  AOI21_X1 U7946 ( .B1(n6380), .B2(n6379), .A(n6378), .ZN(n6381) );
  NOR2_X1 U7947 ( .A1(n9621), .A2(n6381), .ZN(n6382) );
  AOI211_X1 U7948 ( .C1(n9636), .C2(n6383), .A(n6813), .B(n6382), .ZN(n6385)
         );
  NAND2_X1 U7949 ( .A1(n9661), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n6384) );
  OAI211_X1 U7950 ( .C1(n6386), .C2(n9627), .A(n6385), .B(n6384), .ZN(P1_U3247) );
  NOR2_X1 U7951 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6387), .ZN(n6389) );
  NOR2_X1 U7952 ( .A1(n6389), .A2(n6388), .ZN(n6391) );
  AOI22_X1 U7953 ( .A1(n6447), .A2(n8918), .B1(P1_REG2_REG_8__SCAN_IN), .B2(
        n6399), .ZN(n6390) );
  NOR2_X1 U7954 ( .A1(n6391), .A2(n6390), .ZN(n6449) );
  AOI21_X1 U7955 ( .B1(n6391), .B2(n6390), .A(n6449), .ZN(n6402) );
  INV_X1 U7956 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6392) );
  OR2_X1 U7957 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6392), .ZN(n7036) );
  INV_X1 U7958 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9820) );
  AOI21_X1 U7959 ( .B1(n6394), .B2(n9820), .A(n6393), .ZN(n6397) );
  INV_X1 U7960 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6395) );
  MUX2_X1 U7961 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n6395), .S(n6447), .Z(n6396)
         );
  NAND2_X1 U7962 ( .A1(n6396), .A2(n6397), .ZN(n6439) );
  OAI211_X1 U7963 ( .C1(n6397), .C2(n6396), .A(n9663), .B(n6439), .ZN(n6398)
         );
  OAI211_X1 U7964 ( .C1(n9658), .C2(n6399), .A(n7036), .B(n6398), .ZN(n6400)
         );
  AOI21_X1 U7965 ( .B1(n9661), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n6400), .ZN(
        n6401) );
  OAI21_X1 U7966 ( .B1(n6402), .B2(n9627), .A(n6401), .ZN(P1_U3249) );
  INV_X1 U7967 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6404) );
  NAND2_X1 U7968 ( .A1(n9728), .A2(P1_U4006), .ZN(n6403) );
  OAI21_X1 U7969 ( .B1(P1_U4006), .B2(n6404), .A(n6403), .ZN(P1_U3555) );
  INV_X1 U7970 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6419) );
  NOR2_X1 U7971 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8917), .ZN(n6533) );
  INV_X1 U7972 ( .A(n6533), .ZN(n6410) );
  MUX2_X1 U7973 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6359), .S(n6412), .Z(n6406)
         );
  NAND3_X1 U7974 ( .A1(n6406), .A2(n9574), .A3(n6405), .ZN(n6407) );
  NAND3_X1 U7975 ( .A1(n9663), .A2(n6408), .A3(n6407), .ZN(n6409) );
  OAI211_X1 U7976 ( .C1(n9658), .C2(n6412), .A(n6410), .B(n6409), .ZN(n6411)
         );
  INV_X1 U7977 ( .A(n6411), .ZN(n6418) );
  INV_X1 U7978 ( .A(n9627), .ZN(n9667) );
  MUX2_X1 U7979 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6344), .S(n6412), .Z(n6414)
         );
  NAND3_X1 U7980 ( .A1(n6414), .A2(n9585), .A3(n6413), .ZN(n6415) );
  NAND3_X1 U7981 ( .A1(n9667), .A2(n6416), .A3(n6415), .ZN(n6417) );
  OAI211_X1 U7982 ( .C1(n6419), .C2(n9632), .A(n6418), .B(n6417), .ZN(P1_U3244) );
  INV_X1 U7983 ( .A(n6420), .ZN(n6422) );
  OAI222_X1 U7984 ( .A1(n8971), .A2(n6421), .B1(n8969), .B2(n6422), .C1(n10007), .C2(n6974), .ZN(P2_U3346) );
  INV_X1 U7985 ( .A(n6550), .ZN(n6547) );
  OAI222_X1 U7986 ( .A1(n8045), .A2(n8934), .B1(n8048), .B2(n6422), .C1(
        P1_U3084), .C2(n6547), .ZN(P1_U3341) );
  INV_X1 U7987 ( .A(n6736), .ZN(n6426) );
  INV_X1 U7988 ( .A(n9728), .ZN(n6424) );
  NAND2_X1 U7989 ( .A1(n6424), .A2(n6800), .ZN(n9725) );
  NAND2_X1 U7990 ( .A1(n9728), .A2(n4558), .ZN(n7945) );
  NAND2_X1 U7991 ( .A1(n9725), .A2(n7945), .ZN(n7906) );
  NAND3_X1 U7992 ( .A1(n7906), .A2(n6736), .A3(n7170), .ZN(n6425) );
  OAI21_X1 U7993 ( .B1(n6713), .B2(n9701), .A(n6425), .ZN(n6803) );
  AOI21_X1 U7994 ( .B1(n6800), .B2(n6426), .A(n6803), .ZN(n6484) );
  NAND2_X1 U7995 ( .A1(n7939), .A2(n9721), .ZN(n7980) );
  OR2_X1 U7996 ( .A1(n6736), .A2(n7980), .ZN(n6427) );
  NAND2_X1 U7997 ( .A1(n6427), .A2(n6719), .ZN(n6480) );
  NOR2_X1 U7998 ( .A1(n6480), .A2(n6428), .ZN(n6429) );
  INV_X1 U7999 ( .A(n9826), .ZN(n9823) );
  NAND2_X1 U8000 ( .A1(n9823), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6430) );
  OAI21_X1 U8001 ( .B1(n6484), .B2(n9823), .A(n6430), .ZN(P1_U3523) );
  OAI21_X1 U8002 ( .B1(n6433), .B2(n5630), .A(n6432), .ZN(n9579) );
  AOI22_X1 U8003 ( .A1(n9579), .A2(n9086), .B1(n6800), .B2(n9107), .ZN(n6437)
         );
  INV_X1 U8004 ( .A(n6434), .ZN(n6435) );
  OR2_X1 U8005 ( .A1(n9026), .A2(n6435), .ZN(n9025) );
  AOI22_X1 U8006 ( .A1(n9025), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n9101), .B2(
        n6715), .ZN(n6436) );
  NAND2_X1 U8007 ( .A1(n6437), .A2(n6436), .ZN(P1_U3230) );
  NAND2_X1 U8008 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n8466), .ZN(n6438) );
  OAI21_X1 U8009 ( .B1(n7602), .B2(n8466), .A(n6438), .ZN(P2_U3567) );
  NOR2_X1 U8010 ( .A1(n9610), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6442) );
  NAND2_X1 U8011 ( .A1(n6447), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6440) );
  NAND2_X1 U8012 ( .A1(n6440), .A2(n6439), .ZN(n9606) );
  INV_X1 U8013 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9824) );
  INV_X1 U8014 ( .A(n6442), .ZN(n6441) );
  OAI21_X1 U8015 ( .B1(n9824), .B2(n6452), .A(n6441), .ZN(n9605) );
  NOR2_X1 U8016 ( .A1(n9606), .A2(n9605), .ZN(n9604) );
  INV_X1 U8017 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7407) );
  AOI22_X1 U8018 ( .A1(n6485), .A2(n7407), .B1(P1_REG1_REG_10__SCAN_IN), .B2(
        n6491), .ZN(n6443) );
  NOR2_X1 U8019 ( .A1(n6444), .A2(n6443), .ZN(n6490) );
  AOI21_X1 U8020 ( .B1(n6444), .B2(n6443), .A(n6490), .ZN(n6458) );
  NOR2_X1 U8021 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6445), .ZN(n7139) );
  NOR2_X1 U8022 ( .A1(n9658), .A2(n6491), .ZN(n6446) );
  AOI211_X1 U8023 ( .C1(n9661), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n7139), .B(
        n6446), .ZN(n6457) );
  INV_X1 U8024 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6451) );
  NOR2_X1 U8025 ( .A1(n6447), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6448) );
  NOR2_X1 U8026 ( .A1(n6449), .A2(n6448), .ZN(n9613) );
  MUX2_X1 U8027 ( .A(n6451), .B(P1_REG2_REG_9__SCAN_IN), .S(n9610), .Z(n6450)
         );
  INV_X1 U8028 ( .A(n6450), .ZN(n9612) );
  NAND2_X1 U8029 ( .A1(n9613), .A2(n9612), .ZN(n9611) );
  OAI21_X1 U8030 ( .B1(n6452), .B2(n6451), .A(n9611), .ZN(n6455) );
  MUX2_X1 U8031 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n6453), .S(n6485), .Z(n6454)
         );
  NAND2_X1 U8032 ( .A1(n6454), .A2(n6455), .ZN(n6486) );
  OAI211_X1 U8033 ( .C1(n6455), .C2(n6454), .A(n9667), .B(n6486), .ZN(n6456)
         );
  OAI211_X1 U8034 ( .C1(n6458), .C2(n9621), .A(n6457), .B(n6456), .ZN(P1_U3251) );
  INV_X1 U8035 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6471) );
  INV_X1 U8036 ( .A(n6459), .ZN(n6464) );
  AND2_X1 U8037 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6705) );
  AOI211_X1 U8038 ( .C1(n6462), .C2(n6461), .A(n6460), .B(n9621), .ZN(n6463)
         );
  AOI211_X1 U8039 ( .C1(n9636), .C2(n6464), .A(n6705), .B(n6463), .ZN(n6470)
         );
  AND3_X1 U8040 ( .A1(n9591), .A2(n6466), .A3(n6465), .ZN(n6467) );
  OAI21_X1 U8041 ( .B1(n6468), .B2(n6467), .A(n9667), .ZN(n6469) );
  OAI211_X1 U8042 ( .C1(n6471), .C2(n9632), .A(n6470), .B(n6469), .ZN(P1_U3246) );
  INV_X1 U8043 ( .A(n6475), .ZN(n6473) );
  NAND2_X1 U8044 ( .A1(n6473), .A2(n6472), .ZN(n6477) );
  OAI21_X1 U8045 ( .B1(n6475), .B2(P1_D_REG_0__SCAN_IN), .A(n6474), .ZN(n6476)
         );
  AND2_X1 U8046 ( .A1(n6477), .A2(n6476), .ZN(n6478) );
  INV_X1 U8047 ( .A(n6480), .ZN(n6481) );
  INV_X1 U8048 ( .A(n9809), .ZN(n9807) );
  INV_X1 U8049 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6482) );
  OR2_X1 U8050 ( .A1(n9809), .A2(n6482), .ZN(n6483) );
  OAI21_X1 U8051 ( .B1(n6484), .B2(n9807), .A(n6483), .ZN(P1_U3454) );
  NAND2_X1 U8052 ( .A1(n6485), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6487) );
  NAND2_X1 U8053 ( .A1(n6487), .A2(n6486), .ZN(n6489) );
  MUX2_X1 U8054 ( .A(n6518), .B(P1_REG2_REG_11__SCAN_IN), .S(n6492), .Z(n6488)
         );
  NOR2_X1 U8055 ( .A1(n6489), .A2(n6488), .ZN(n6516) );
  AOI21_X1 U8056 ( .B1(n6489), .B2(n6488), .A(n6516), .ZN(n6501) );
  INV_X1 U8057 ( .A(n6490), .ZN(n6496) );
  NAND2_X1 U8058 ( .A1(n6491), .A2(n7407), .ZN(n6494) );
  INV_X1 U8059 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6493) );
  MUX2_X1 U8060 ( .A(n6493), .B(P1_REG1_REG_11__SCAN_IN), .S(n6492), .Z(n6495)
         );
  AOI21_X1 U8061 ( .B1(n6496), .B2(n6494), .A(n6495), .ZN(n6513) );
  AND3_X1 U8062 ( .A1(n6496), .A2(n6495), .A3(n6494), .ZN(n6497) );
  OAI21_X1 U8063 ( .B1(n6513), .B2(n6497), .A(n9663), .ZN(n6500) );
  AND2_X1 U8064 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7231) );
  NOR2_X1 U8065 ( .A1(n9658), .A2(n6517), .ZN(n6498) );
  AOI211_X1 U8066 ( .C1(n9661), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n7231), .B(
        n6498), .ZN(n6499) );
  OAI211_X1 U8067 ( .C1(n6501), .C2(n9627), .A(n6500), .B(n6499), .ZN(P1_U3252) );
  INV_X1 U8068 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6506) );
  NAND2_X1 U8069 ( .A1(n5675), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6504) );
  NAND2_X1 U8070 ( .A1(n6153), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6503) );
  NAND2_X1 U8071 ( .A1(n7723), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6502) );
  AND3_X1 U8072 ( .A1(n6504), .A2(n6503), .A3(n6502), .ZN(n9142) );
  INV_X1 U8073 ( .A(n9142), .ZN(n7791) );
  NAND2_X1 U8074 ( .A1(n7791), .A2(P1_U4006), .ZN(n6505) );
  OAI21_X1 U8075 ( .B1(P1_U4006), .B2(n6506), .A(n6505), .ZN(P1_U3586) );
  INV_X1 U8076 ( .A(n6507), .ZN(n6509) );
  AOI22_X1 U8077 ( .A1(n6985), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n8967), .ZN(n6508) );
  OAI21_X1 U8078 ( .B1(n6509), .B2(n8975), .A(n6508), .ZN(P2_U3345) );
  INV_X1 U8079 ( .A(n6559), .ZN(n7448) );
  OAI222_X1 U8080 ( .A1(n8045), .A2(n6510), .B1(n8048), .B2(n6509), .C1(n7448), 
        .C2(P1_U3084), .ZN(P1_U3340) );
  INV_X1 U8081 ( .A(n6511), .ZN(n6512) );
  INV_X1 U8082 ( .A(n7219), .ZN(n7416) );
  OAI222_X1 U8083 ( .A1(n8969), .A2(n6512), .B1(n7416), .B2(P2_U3152), .C1(
        n8891), .C2(n8971), .ZN(P2_U3344) );
  INV_X1 U8084 ( .A(n9624), .ZN(n7450) );
  OAI222_X1 U8085 ( .A1(n8045), .A2(n8935), .B1(n8048), .B2(n6512), .C1(n7450), 
        .C2(P1_U3084), .ZN(P1_U3339) );
  INV_X1 U8086 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9534) );
  AOI22_X1 U8087 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n6547), .B1(n6550), .B2(
        n9534), .ZN(n6514) );
  NOR2_X1 U8088 ( .A1(n6515), .A2(n6514), .ZN(n6546) );
  AOI21_X1 U8089 ( .B1(n6515), .B2(n6514), .A(n6546), .ZN(n6524) );
  INV_X1 U8090 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6518) );
  AOI21_X1 U8091 ( .B1(n6518), .B2(n6517), .A(n6516), .ZN(n6553) );
  MUX2_X1 U8092 ( .A(n5858), .B(P1_REG2_REG_12__SCAN_IN), .S(n6550), .Z(n6551)
         );
  XNOR2_X1 U8093 ( .A(n6553), .B(n6551), .ZN(n6522) );
  NAND2_X1 U8094 ( .A1(n9661), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6520) );
  NAND2_X1 U8095 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n6519) );
  OAI211_X1 U8096 ( .C1(n9658), .C2(n6547), .A(n6520), .B(n6519), .ZN(n6521)
         );
  AOI21_X1 U8097 ( .B1(n6522), .B2(n9667), .A(n6521), .ZN(n6523) );
  OAI21_X1 U8098 ( .B1(n6524), .B2(n9621), .A(n6523), .ZN(P1_U3253) );
  NAND2_X1 U8099 ( .A1(n6527), .A2(n9086), .ZN(n6530) );
  INV_X1 U8100 ( .A(n9101), .ZN(n9453) );
  OAI22_X1 U8101 ( .A1(n9453), .A2(n6928), .B1(n9104), .B2(n6713), .ZN(n6528)
         );
  AOI21_X1 U8102 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n9025), .A(n6528), .ZN(
        n6529) );
  OAI211_X1 U8103 ( .C1(n6718), .C2(n9095), .A(n6530), .B(n6529), .ZN(P1_U3235) );
  XOR2_X1 U8104 ( .A(n6532), .B(n6531), .Z(n6538) );
  AOI21_X1 U8105 ( .B1(n9101), .B2(n9675), .A(n6533), .ZN(n6535) );
  INV_X1 U8106 ( .A(n9104), .ZN(n9456) );
  NAND2_X1 U8107 ( .A1(n9456), .A2(n9727), .ZN(n6534) );
  OAI211_X1 U8108 ( .C1(n9095), .C2(n6927), .A(n6535), .B(n6534), .ZN(n6536)
         );
  AOI21_X1 U8109 ( .B1(n9099), .B2(n8917), .A(n6536), .ZN(n6537) );
  OAI21_X1 U8110 ( .B1(n6538), .B2(n9460), .A(n6537), .ZN(P1_U3216) );
  INV_X1 U8111 ( .A(n6539), .ZN(n6543) );
  AOI22_X1 U8112 ( .A1(n9635), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n7594), .ZN(n6540) );
  OAI21_X1 U8113 ( .B1(n6543), .B2(n8048), .A(n6540), .ZN(P1_U3338) );
  INV_X1 U8114 ( .A(n6541), .ZN(n6545) );
  AOI22_X1 U8115 ( .A1(n7462), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n7594), .ZN(n6542) );
  OAI21_X1 U8116 ( .B1(n6545), .B2(n8048), .A(n6542), .ZN(P1_U3337) );
  INV_X1 U8117 ( .A(n7509), .ZN(n7417) );
  OAI222_X1 U8118 ( .A1(n8971), .A2(n6544), .B1(n8969), .B2(n6543), .C1(
        P2_U3152), .C2(n7417), .ZN(P2_U3343) );
  INV_X1 U8119 ( .A(n8477), .ZN(n7505) );
  OAI222_X1 U8120 ( .A1(n8969), .A2(n6545), .B1(n7505), .B2(n10007), .C1(n8831), .C2(n8971), .ZN(P2_U3342) );
  AOI21_X1 U8121 ( .B1(n9534), .B2(n6547), .A(n6546), .ZN(n6549) );
  INV_X1 U8122 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9528) );
  AOI22_X1 U8123 ( .A1(P1_REG1_REG_13__SCAN_IN), .A2(n7448), .B1(n6559), .B2(
        n9528), .ZN(n6548) );
  NOR2_X1 U8124 ( .A1(n6549), .A2(n6548), .ZN(n7447) );
  AOI21_X1 U8125 ( .B1(n6549), .B2(n6548), .A(n7447), .ZN(n6565) );
  INV_X1 U8126 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6562) );
  NAND2_X1 U8127 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n6550), .ZN(n6555) );
  INV_X1 U8128 ( .A(n6551), .ZN(n6552) );
  NAND2_X1 U8129 ( .A1(n6553), .A2(n6552), .ZN(n6554) );
  NAND2_X1 U8130 ( .A1(n6555), .A2(n6554), .ZN(n6558) );
  OR2_X1 U8131 ( .A1(n6559), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6556) );
  NAND2_X1 U8132 ( .A1(n6559), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7465) );
  AND2_X1 U8133 ( .A1(n6556), .A2(n7465), .ZN(n6557) );
  NAND2_X1 U8134 ( .A1(n6557), .A2(n6558), .ZN(n7464) );
  OAI211_X1 U8135 ( .C1(n6558), .C2(n6557), .A(n9667), .B(n7464), .ZN(n6561)
         );
  NOR2_X1 U8136 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5877), .ZN(n7426) );
  AOI21_X1 U8137 ( .B1(n9636), .B2(n6559), .A(n7426), .ZN(n6560) );
  OAI211_X1 U8138 ( .C1(n9632), .C2(n6562), .A(n6561), .B(n6560), .ZN(n6563)
         );
  INV_X1 U8139 ( .A(n6563), .ZN(n6564) );
  OAI21_X1 U8140 ( .B1(n6565), .B2(n9621), .A(n6564), .ZN(P1_U3254) );
  INV_X1 U8141 ( .A(n6566), .ZN(n6568) );
  AOI22_X1 U8142 ( .A1(n9875), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n8967), .ZN(n6567) );
  OAI21_X1 U8143 ( .B1(n6568), .B2(n8969), .A(n6567), .ZN(P2_U3341) );
  INV_X1 U8144 ( .A(n7460), .ZN(n9657) );
  OAI222_X1 U8145 ( .A1(n8045), .A2(n6569), .B1(n8048), .B2(n6568), .C1(n9657), 
        .C2(P1_U3084), .ZN(P1_U3336) );
  NAND3_X1 U8146 ( .A1(n6570), .A2(n6877), .A3(n6878), .ZN(n6572) );
  INV_X1 U8147 ( .A(n6875), .ZN(n6573) );
  INV_X1 U8148 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6596) );
  NAND2_X1 U8149 ( .A1(n8465), .A2(n6884), .ZN(n6584) );
  OR2_X2 U8150 ( .A1(n8464), .A2(n9916), .ZN(n8274) );
  NAND2_X1 U8151 ( .A1(n7005), .A2(n8402), .ZN(n6576) );
  INV_X1 U8152 ( .A(n8464), .ZN(n6574) );
  NAND2_X1 U8153 ( .A1(n6574), .A2(n9916), .ZN(n6575) );
  NAND2_X1 U8154 ( .A1(n6576), .A2(n6575), .ZN(n6598) );
  OR2_X1 U8155 ( .A1(n8463), .A2(n6915), .ZN(n7012) );
  NAND2_X1 U8156 ( .A1(n8463), .A2(n6915), .ZN(n8250) );
  NAND2_X1 U8157 ( .A1(n7012), .A2(n8250), .ZN(n6601) );
  NAND2_X1 U8158 ( .A1(n6598), .A2(n6601), .ZN(n6597) );
  INV_X1 U8159 ( .A(n8463), .ZN(n7017) );
  NAND2_X1 U8160 ( .A1(n7017), .A2(n6915), .ZN(n6577) );
  NAND2_X1 U8161 ( .A1(n6597), .A2(n6577), .ZN(n7024) );
  NAND2_X1 U8162 ( .A1(n8462), .A2(n9920), .ZN(n6747) );
  NAND2_X1 U8163 ( .A1(n8248), .A2(n6747), .ZN(n8406) );
  NAND2_X1 U8164 ( .A1(n7024), .A2(n8406), .ZN(n7023) );
  NAND2_X1 U8165 ( .A1(n4448), .A2(n9920), .ZN(n6578) );
  NAND2_X1 U8166 ( .A1(n7023), .A2(n6578), .ZN(n6579) );
  NAND2_X1 U8167 ( .A1(n8267), .A2(n8249), .ZN(n8407) );
  OAI21_X1 U8168 ( .B1(n6579), .B2(n8407), .A(n6743), .ZN(n6997) );
  INV_X1 U8169 ( .A(n6997), .ZN(n6594) );
  OAI22_X1 U8170 ( .A1(n8442), .A2(n6581), .B1(n7088), .B2(n6580), .ZN(n6582)
         );
  NAND2_X1 U8171 ( .A1(n6582), .A2(n8399), .ZN(n7600) );
  OR3_X1 U8172 ( .A1(n5535), .A2(n8444), .A3(n8583), .ZN(n7480) );
  INV_X1 U8173 ( .A(n6995), .ZN(n7995) );
  NOR2_X1 U8174 ( .A1(n6884), .A2(n9898), .ZN(n6883) );
  NAND2_X1 U8175 ( .A1(n6883), .A2(n9916), .ZN(n9911) );
  INV_X1 U8176 ( .A(n6915), .ZN(n6655) );
  OR2_X1 U8177 ( .A1(n9911), .A2(n6655), .ZN(n6605) );
  NOR2_X1 U8178 ( .A1(n6605), .A2(n4449), .ZN(n6583) );
  INV_X1 U8179 ( .A(n6583), .ZN(n7019) );
  AOI211_X1 U8180 ( .C1(n7995), .C2(n7019), .A(n9936), .B(n7126), .ZN(n6993)
         );
  AOI21_X1 U8181 ( .B1(n9475), .B2(n7995), .A(n6993), .ZN(n6593) );
  NOR2_X1 U8182 ( .A1(n8467), .A2(n6947), .ZN(n8260) );
  OR2_X1 U8183 ( .A1(n8465), .A2(n9907), .ZN(n8273) );
  NAND2_X1 U8184 ( .A1(n7000), .A2(n8273), .ZN(n6587) );
  INV_X1 U8185 ( .A(n8402), .ZN(n6586) );
  NAND2_X1 U8186 ( .A1(n6587), .A2(n6586), .ZN(n7002) );
  NAND2_X1 U8187 ( .A1(n7002), .A2(n8274), .ZN(n6588) );
  INV_X1 U8188 ( .A(n6601), .ZN(n8405) );
  AND2_X1 U8189 ( .A1(n7012), .A2(n8248), .ZN(n8268) );
  NAND2_X1 U8190 ( .A1(n7013), .A2(n8268), .ZN(n6748) );
  NAND2_X1 U8191 ( .A1(n6748), .A2(n6747), .ZN(n6589) );
  XNOR2_X1 U8192 ( .A(n6589), .B(n8407), .ZN(n6592) );
  NAND2_X1 U8193 ( .A1(n8444), .A2(n8569), .ZN(n8434) );
  OR2_X1 U8194 ( .A1(n6751), .A2(n8564), .ZN(n6591) );
  NAND2_X1 U8195 ( .A1(n8462), .A2(n8656), .ZN(n6590) );
  NAND2_X1 U8196 ( .A1(n6591), .A2(n6590), .ZN(n7987) );
  AOI21_X1 U8197 ( .B1(n6592), .B2(n8659), .A(n7987), .ZN(n6999) );
  OAI211_X1 U8198 ( .C1(n6594), .C2(n8785), .A(n6593), .B(n6999), .ZN(n6613)
         );
  NAND2_X1 U8199 ( .A1(n6613), .A2(n9944), .ZN(n6595) );
  OAI21_X1 U8200 ( .B1(n9944), .B2(n6596), .A(n6595), .ZN(P2_U3466) );
  INV_X1 U8201 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6608) );
  OAI21_X1 U8202 ( .B1(n6598), .B2(n6601), .A(n6597), .ZN(n6604) );
  INV_X1 U8203 ( .A(n6604), .ZN(n6916) );
  INV_X1 U8204 ( .A(n7600), .ZN(n7371) );
  NAND2_X1 U8205 ( .A1(n8464), .A2(n8656), .ZN(n6600) );
  NAND2_X1 U8206 ( .A1(n8462), .A2(n8654), .ZN(n6599) );
  NAND2_X1 U8207 ( .A1(n6600), .A2(n6599), .ZN(n6652) );
  NAND3_X1 U8208 ( .A1(n7002), .A2(n8274), .A3(n6601), .ZN(n6602) );
  AOI21_X1 U8209 ( .B1(n7013), .B2(n6602), .A(n8707), .ZN(n6603) );
  AOI211_X1 U8210 ( .C1(n7371), .C2(n6604), .A(n6652), .B(n6603), .ZN(n6921)
         );
  INV_X1 U8211 ( .A(n6605), .ZN(n7020) );
  AOI21_X1 U8212 ( .B1(n6655), .B2(n9911), .A(n7020), .ZN(n6919) );
  AOI22_X1 U8213 ( .A1(n6919), .A2(n9912), .B1(n9475), .B2(n6655), .ZN(n6606)
         );
  OAI211_X1 U8214 ( .C1(n6916), .C2(n7480), .A(n6921), .B(n6606), .ZN(n6610)
         );
  NAND2_X1 U8215 ( .A1(n6610), .A2(n9944), .ZN(n6607) );
  OAI21_X1 U8216 ( .B1(n9944), .B2(n6608), .A(n6607), .ZN(P2_U3460) );
  INV_X1 U8217 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6612) );
  NAND2_X1 U8218 ( .A1(n6610), .A2(n9954), .ZN(n6611) );
  OAI21_X1 U8219 ( .B1(n9954), .B2(n6612), .A(n6611), .ZN(P2_U3523) );
  INV_X1 U8220 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6615) );
  NAND2_X1 U8221 ( .A1(n6613), .A2(n9954), .ZN(n6614) );
  OAI21_X1 U8222 ( .B1(n9954), .B2(n6615), .A(n6614), .ZN(P2_U3525) );
  INV_X1 U8223 ( .A(n6846), .ZN(n6616) );
  AOI21_X1 U8224 ( .B1(n6618), .B2(n6617), .A(n6616), .ZN(n6622) );
  AOI22_X1 U8225 ( .A1(n8194), .A2(n8467), .B1(n9828), .B2(n8464), .ZN(n6621)
         );
  NAND2_X1 U8226 ( .A1(n9478), .A2(n6619), .ZN(n6841) );
  AOI22_X1 U8227 ( .A1(n9854), .A2(n6884), .B1(n6841), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n6620) );
  OAI211_X1 U8228 ( .C1(n6622), .C2(n9835), .A(n6621), .B(n6620), .ZN(P2_U3224) );
  INV_X1 U8229 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n9983) );
  INV_X1 U8230 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6625) );
  OAI21_X1 U8231 ( .B1(n6625), .B2(n6624), .A(n6623), .ZN(n6627) );
  XOR2_X1 U8232 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6645), .Z(n6626) );
  NAND2_X1 U8233 ( .A1(n6627), .A2(n6626), .ZN(n6637) );
  OAI211_X1 U8234 ( .C1(n6627), .C2(n6626), .A(n6637), .B(n9871), .ZN(n6629)
         );
  NAND2_X1 U8235 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n6628) );
  OAI211_X1 U8236 ( .C1(n9983), .C2(n8506), .A(n6629), .B(n6628), .ZN(n6635)
         );
  XNOR2_X1 U8237 ( .A(n6645), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n6632) );
  NOR2_X1 U8238 ( .A1(n6633), .A2(n6632), .ZN(n6644) );
  AOI211_X1 U8239 ( .C1(n6633), .C2(n6632), .A(n8490), .B(n6644), .ZN(n6634)
         );
  AOI211_X1 U8240 ( .C1(n9876), .C2(n6645), .A(n6635), .B(n6634), .ZN(n6636)
         );
  INV_X1 U8241 ( .A(n6636), .ZN(P2_U3253) );
  INV_X1 U8242 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n6643) );
  INV_X1 U8243 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6639) );
  OAI21_X1 U8244 ( .B1(n6639), .B2(n6638), .A(n6637), .ZN(n6641) );
  INV_X1 U8245 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6965) );
  MUX2_X1 U8246 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n6965), .S(n6666), .Z(n6640)
         );
  NAND2_X1 U8247 ( .A1(n6641), .A2(n6640), .ZN(n6664) );
  OAI211_X1 U8248 ( .C1(n6641), .C2(n6640), .A(n6664), .B(n9871), .ZN(n6642)
         );
  NAND2_X1 U8249 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(n10007), .ZN(n8179) );
  OAI211_X1 U8250 ( .C1(n6643), .C2(n8506), .A(n6642), .B(n8179), .ZN(n6650)
         );
  AOI21_X1 U8251 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n6645), .A(n6644), .ZN(
        n6648) );
  NAND2_X1 U8252 ( .A1(P2_REG2_REG_9__SCAN_IN), .A2(n6666), .ZN(n6646) );
  OAI21_X1 U8253 ( .B1(n6666), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6646), .ZN(
        n6647) );
  NOR2_X1 U8254 ( .A1(n6648), .A2(n6647), .ZN(n6660) );
  AOI211_X1 U8255 ( .C1(n6648), .C2(n6647), .A(n8490), .B(n6660), .ZN(n6649)
         );
  AOI211_X1 U8256 ( .C1(n9876), .C2(n6666), .A(n6650), .B(n6649), .ZN(n6651)
         );
  INV_X1 U8257 ( .A(n6651), .ZN(P2_U3254) );
  INV_X1 U8258 ( .A(n8209), .ZN(n9844) );
  AOI22_X1 U8259 ( .A1(n9844), .A2(n6652), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        P2_U3152), .ZN(n6653) );
  OAI21_X1 U8260 ( .B1(n9860), .B2(P2_REG3_REG_3__SCAN_IN), .A(n6653), .ZN(
        n6654) );
  AOI21_X1 U8261 ( .B1(n9854), .B2(n6655), .A(n6654), .ZN(n6659) );
  OAI211_X1 U8262 ( .C1(n6657), .C2(n6656), .A(n6850), .B(n9845), .ZN(n6658)
         );
  NAND2_X1 U8263 ( .A1(n6659), .A2(n6658), .ZN(P2_U3220) );
  NAND2_X1 U8264 ( .A1(n6694), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6661) );
  OAI21_X1 U8265 ( .B1(n6694), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6661), .ZN(
        n6662) );
  AOI211_X1 U8266 ( .C1(n6663), .C2(n6662), .A(n6693), .B(n8490), .ZN(n6673)
         );
  INV_X1 U8267 ( .A(n6664), .ZN(n6665) );
  INV_X1 U8268 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6667) );
  MUX2_X1 U8269 ( .A(n6667), .B(P2_REG1_REG_10__SCAN_IN), .S(n6694), .Z(n6668)
         );
  NOR2_X1 U8270 ( .A1(n6669), .A2(n6668), .ZN(n6687) );
  AOI211_X1 U8271 ( .C1(n6669), .C2(n6668), .A(n6687), .B(n9862), .ZN(n6672)
         );
  INV_X1 U8272 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n8881) );
  NAND2_X1 U8273 ( .A1(n9876), .A2(n6694), .ZN(n6670) );
  NAND2_X1 U8274 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(n10007), .ZN(n9829) );
  OAI211_X1 U8275 ( .C1(n8881), .C2(n8506), .A(n6670), .B(n9829), .ZN(n6671)
         );
  OR3_X1 U8276 ( .A1(n6673), .A2(n6672), .A3(n6671), .ZN(P2_U3255) );
  INV_X1 U8277 ( .A(n6674), .ZN(n6711) );
  AOI22_X1 U8278 ( .A1(n8480), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n8967), .ZN(n6675) );
  OAI21_X1 U8279 ( .B1(n6711), .B2(n8969), .A(n6675), .ZN(P2_U3340) );
  NAND2_X1 U8280 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9602) );
  INV_X1 U8281 ( .A(n9602), .ZN(n6676) );
  AOI21_X1 U8282 ( .B1(n9101), .B2(n9124), .A(n6676), .ZN(n6678) );
  NAND2_X1 U8283 ( .A1(n9456), .A2(n9125), .ZN(n6677) );
  OAI211_X1 U8284 ( .C1(n9095), .C2(n9764), .A(n6678), .B(n6677), .ZN(n6684)
         );
  INV_X1 U8285 ( .A(n6680), .ZN(n6681) );
  AOI211_X1 U8286 ( .C1(n6682), .C2(n6679), .A(n9460), .B(n6681), .ZN(n6683)
         );
  AOI211_X1 U8287 ( .C1(n9099), .C2(n6933), .A(n6684), .B(n6683), .ZN(n6685)
         );
  INV_X1 U8288 ( .A(n6685), .ZN(P1_U3228) );
  INV_X1 U8289 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n6686) );
  NOR2_X1 U8290 ( .A1(n8506), .A2(n6686), .ZN(n6692) );
  AOI21_X1 U8291 ( .B1(n6694), .B2(P2_REG1_REG_10__SCAN_IN), .A(n6687), .ZN(
        n6690) );
  INV_X1 U8292 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6688) );
  MUX2_X1 U8293 ( .A(n6688), .B(P2_REG1_REG_11__SCAN_IN), .S(n6791), .Z(n6689)
         );
  NOR2_X1 U8294 ( .A1(n6690), .A2(n6689), .ZN(n6790) );
  AOI211_X1 U8295 ( .C1(n6690), .C2(n6689), .A(n6790), .B(n9862), .ZN(n6691)
         );
  AOI211_X1 U8296 ( .C1(P2_REG3_REG_11__SCAN_IN), .C2(n10007), .A(n6692), .B(
        n6691), .ZN(n6699) );
  INV_X1 U8297 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8850) );
  AOI22_X1 U8298 ( .A1(n6791), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n8850), .B2(
        n6700), .ZN(n6696) );
  OAI21_X1 U8299 ( .B1(n6696), .B2(n6695), .A(n6789), .ZN(n6697) );
  NAND2_X1 U8300 ( .A1(n6697), .A2(n9879), .ZN(n6698) );
  OAI211_X1 U8301 ( .C1(n9861), .C2(n6700), .A(n6699), .B(n6698), .ZN(P2_U3256) );
  INV_X1 U8302 ( .A(n9686), .ZN(n6710) );
  OAI21_X1 U8303 ( .B1(n6703), .B2(n6702), .A(n6701), .ZN(n6704) );
  NAND2_X1 U8304 ( .A1(n6704), .A2(n9086), .ZN(n6709) );
  INV_X1 U8305 ( .A(n9026), .ZN(n9464) );
  AND2_X1 U8306 ( .A1(n9422), .A2(n9687), .ZN(n9770) );
  AOI21_X1 U8307 ( .B1(n9101), .B2(n9676), .A(n6705), .ZN(n6706) );
  OAI21_X1 U8308 ( .B1(n9702), .B2(n9104), .A(n6706), .ZN(n6707) );
  AOI21_X1 U8309 ( .B1(n9464), .B2(n9770), .A(n6707), .ZN(n6708) );
  OAI211_X1 U8310 ( .C1(n9468), .C2(n6710), .A(n6709), .B(n6708), .ZN(P1_U3225) );
  INV_X1 U8311 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6712) );
  INV_X1 U8312 ( .A(n7472), .ZN(n9130) );
  OAI222_X1 U8313 ( .A1(n8045), .A2(n6712), .B1(n8048), .B2(n6711), .C1(
        P1_U3084), .C2(n9130), .ZN(P1_U3335) );
  NAND2_X1 U8314 ( .A1(n9728), .A2(n6800), .ZN(n9715) );
  NAND2_X1 U8315 ( .A1(n6726), .A2(n9715), .ZN(n6717) );
  NAND2_X1 U8316 ( .A1(n6713), .A2(n6714), .ZN(n6716) );
  NAND2_X1 U8317 ( .A1(n6717), .A2(n6716), .ZN(n6923) );
  XNOR2_X1 U8318 ( .A(n6922), .B(n6923), .ZN(n9757) );
  INV_X1 U8319 ( .A(n9757), .ZN(n6741) );
  INV_X1 U8320 ( .A(n6719), .ZN(n6720) );
  NAND2_X1 U8321 ( .A1(n6721), .A2(n6720), .ZN(n7175) );
  NOR2_X1 U8322 ( .A1(n8041), .A2(n7980), .ZN(n9736) );
  NAND2_X1 U8323 ( .A1(n9737), .A2(n9736), .ZN(n7590) );
  NAND2_X1 U8324 ( .A1(n8043), .A2(n9137), .ZN(n6725) );
  MUX2_X1 U8325 ( .A(n6725), .B(n6724), .S(n6723), .Z(n9707) );
  INV_X1 U8326 ( .A(n9707), .ZN(n9730) );
  NAND2_X1 U8327 ( .A1(n9757), .A2(n9730), .ZN(n6734) );
  NAND2_X1 U8328 ( .A1(n9722), .A2(n6727), .ZN(n6728) );
  INV_X1 U8329 ( .A(n6922), .ZN(n7908) );
  OAI21_X1 U8330 ( .B1(n6728), .B2(n7908), .A(n6938), .ZN(n6731) );
  OR2_X1 U8331 ( .A1(n8043), .A2(n9137), .ZN(n6730) );
  OR2_X1 U8332 ( .A1(n8041), .A2(n7939), .ZN(n6729) );
  NAND2_X1 U8333 ( .A1(n6731), .A2(n9704), .ZN(n6733) );
  AOI22_X1 U8334 ( .A1(n9726), .A2(n9125), .B1(n6715), .B2(n9729), .ZN(n6732)
         );
  NAND3_X1 U8335 ( .A1(n6734), .A2(n6733), .A3(n6732), .ZN(n9755) );
  MUX2_X1 U8336 ( .A(n9755), .B(P1_REG2_REG_2__SCAN_IN), .S(n9739), .Z(n6735)
         );
  INV_X1 U8337 ( .A(n6735), .ZN(n6740) );
  NOR2_X1 U8338 ( .A1(n9716), .A2(n6936), .ZN(n9694) );
  AND2_X1 U8339 ( .A1(n9716), .A2(n6936), .ZN(n6737) );
  NOR2_X1 U8340 ( .A1(n9694), .A2(n6737), .ZN(n9753) );
  OAI22_X1 U8341 ( .A1(n9710), .A2(n6718), .B1(n9709), .B2(n9590), .ZN(n6738)
         );
  AOI21_X1 U8342 ( .B1(n9696), .B2(n9753), .A(n6738), .ZN(n6739) );
  OAI211_X1 U8343 ( .C1(n6741), .C2(n7590), .A(n6740), .B(n6739), .ZN(P1_U3289) );
  INV_X1 U8344 ( .A(n8461), .ZN(n7016) );
  NAND2_X1 U8345 ( .A1(n7016), .A2(n6995), .ZN(n6742) );
  NAND2_X1 U8346 ( .A1(n6751), .A2(n7130), .ZN(n8285) );
  INV_X1 U8347 ( .A(n6751), .ZN(n8460) );
  NAND2_X1 U8348 ( .A1(n8460), .A2(n9926), .ZN(n8279) );
  NAND2_X1 U8349 ( .A1(n6751), .A2(n9926), .ZN(n6744) );
  NAND2_X1 U8350 ( .A1(n6825), .A2(n6767), .ZN(n8286) );
  INV_X1 U8351 ( .A(n6825), .ZN(n9848) );
  NAND2_X1 U8352 ( .A1(n4425), .A2(n9848), .ZN(n8287) );
  NAND2_X1 U8353 ( .A1(n8286), .A2(n8287), .ZN(n8283) );
  OAI21_X1 U8354 ( .B1(n6745), .B2(n8283), .A(n6773), .ZN(n6746) );
  INV_X1 U8355 ( .A(n6746), .ZN(n6901) );
  NAND2_X1 U8356 ( .A1(n6748), .A2(n8251), .ZN(n6749) );
  NAND2_X1 U8357 ( .A1(n6749), .A2(n8267), .ZN(n7119) );
  INV_X1 U8358 ( .A(n8408), .ZN(n7118) );
  INV_X1 U8359 ( .A(n6778), .ZN(n6774) );
  AOI211_X1 U8360 ( .C1(n6750), .C2(n8283), .A(n8707), .B(n6774), .ZN(n6754)
         );
  OR2_X1 U8361 ( .A1(n6751), .A2(n8562), .ZN(n6753) );
  OR2_X1 U8362 ( .A1(n6954), .A2(n8564), .ZN(n6752) );
  NAND2_X1 U8363 ( .A1(n6753), .A2(n6752), .ZN(n6766) );
  NOR2_X1 U8364 ( .A1(n6754), .A2(n6766), .ZN(n6896) );
  INV_X1 U8365 ( .A(n6783), .ZN(n6755) );
  AOI211_X1 U8366 ( .C1(n6767), .C2(n7125), .A(n9936), .B(n6755), .ZN(n6899)
         );
  AOI21_X1 U8367 ( .B1(n9475), .B2(n6767), .A(n6899), .ZN(n6756) );
  OAI211_X1 U8368 ( .C1(n8785), .C2(n6901), .A(n6896), .B(n6756), .ZN(n6758)
         );
  NAND2_X1 U8369 ( .A1(n6758), .A2(n9954), .ZN(n6757) );
  OAI21_X1 U8370 ( .B1(n9954), .B2(n6625), .A(n6757), .ZN(P2_U3527) );
  INV_X1 U8371 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6760) );
  NAND2_X1 U8372 ( .A1(n6758), .A2(n9944), .ZN(n6759) );
  OAI21_X1 U8373 ( .B1(n9944), .B2(n6760), .A(n6759), .ZN(P2_U3472) );
  INV_X1 U8374 ( .A(n6761), .ZN(n9847) );
  AOI211_X1 U8375 ( .C1(n6763), .C2(n6762), .A(n9835), .B(n9847), .ZN(n6772)
         );
  INV_X1 U8376 ( .A(n6894), .ZN(n6770) );
  INV_X1 U8377 ( .A(n6764), .ZN(n6765) );
  AOI21_X1 U8378 ( .B1(n9844), .B2(n6766), .A(n6765), .ZN(n6769) );
  NAND2_X1 U8379 ( .A1(n9854), .A2(n6767), .ZN(n6768) );
  OAI211_X1 U8380 ( .C1(n9860), .C2(n6770), .A(n6769), .B(n6768), .ZN(n6771)
         );
  OR2_X1 U8381 ( .A1(n6772), .A2(n6771), .ZN(P2_U3215) );
  INV_X1 U8382 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n6786) );
  OR2_X1 U8383 ( .A1(n9853), .A2(n6954), .ZN(n8290) );
  NAND2_X1 U8384 ( .A1(n9853), .A2(n6954), .ZN(n8291) );
  INV_X1 U8385 ( .A(n8410), .ZN(n6776) );
  OAI21_X1 U8386 ( .B1(n4273), .B2(n6776), .A(n6956), .ZN(n6910) );
  INV_X1 U8387 ( .A(n8287), .ZN(n6775) );
  OAI21_X1 U8388 ( .B1(n6774), .B2(n6775), .A(n6776), .ZN(n6779) );
  NOR2_X1 U8389 ( .A1(n6776), .A2(n6775), .ZN(n6777) );
  AOI21_X1 U8390 ( .B1(n6779), .B2(n6957), .A(n8707), .ZN(n6782) );
  OR2_X1 U8391 ( .A1(n6825), .A2(n8562), .ZN(n6781) );
  OR2_X1 U8392 ( .A1(n9832), .A2(n8564), .ZN(n6780) );
  NAND2_X1 U8393 ( .A1(n6781), .A2(n6780), .ZN(n9843) );
  NOR2_X1 U8394 ( .A1(n6782), .A2(n9843), .ZN(n6905) );
  AOI211_X1 U8395 ( .C1(n9853), .C2(n6783), .A(n9936), .B(n6959), .ZN(n6908)
         );
  AOI21_X1 U8396 ( .B1(n9475), .B2(n9853), .A(n6908), .ZN(n6784) );
  OAI211_X1 U8397 ( .C1(n6910), .C2(n8785), .A(n6905), .B(n6784), .ZN(n6787)
         );
  NAND2_X1 U8398 ( .A1(n6787), .A2(n9944), .ZN(n6785) );
  OAI21_X1 U8399 ( .B1(n9944), .B2(n6786), .A(n6785), .ZN(P2_U3475) );
  NAND2_X1 U8400 ( .A1(n6787), .A2(n9954), .ZN(n6788) );
  OAI21_X1 U8401 ( .B1(n9954), .B2(n6639), .A(n6788), .ZN(P2_U3528) );
  OAI21_X1 U8402 ( .B1(n6791), .B2(P2_REG2_REG_11__SCAN_IN), .A(n6789), .ZN(
        n6967) );
  XNOR2_X1 U8403 ( .A(n6968), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n6969) );
  XNOR2_X1 U8404 ( .A(n6967), .B(n6969), .ZN(n6799) );
  INV_X1 U8405 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6796) );
  INV_X1 U8406 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6973) );
  MUX2_X1 U8407 ( .A(n6973), .B(P2_REG1_REG_12__SCAN_IN), .S(n6974), .Z(n6792)
         );
  NAND2_X1 U8408 ( .A1(n6792), .A2(n6793), .ZN(n6976) );
  OAI21_X1 U8409 ( .B1(n6793), .B2(n6792), .A(n6976), .ZN(n6794) );
  NAND2_X1 U8410 ( .A1(n9871), .A2(n6794), .ZN(n6795) );
  NAND2_X1 U8411 ( .A1(P2_U3152), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7349) );
  OAI211_X1 U8412 ( .C1(n8506), .C2(n6796), .A(n6795), .B(n7349), .ZN(n6797)
         );
  AOI21_X1 U8413 ( .B1(n6968), .B2(n9876), .A(n6797), .ZN(n6798) );
  OAI21_X1 U8414 ( .B1(n6799), .B2(n8490), .A(n6798), .ZN(P2_U3257) );
  INV_X1 U8415 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6806) );
  INV_X1 U8416 ( .A(n9710), .ZN(n9498) );
  OAI21_X1 U8417 ( .B1(n9696), .B2(n9498), .A(n6800), .ZN(n6805) );
  INV_X1 U8418 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6801) );
  NOR2_X1 U8419 ( .A1(n9709), .A2(n6801), .ZN(n6802) );
  OAI21_X1 U8420 ( .B1(n6803), .B2(n6802), .A(n9737), .ZN(n6804) );
  OAI211_X1 U8421 ( .C1(n6806), .C2(n9737), .A(n6805), .B(n6804), .ZN(P1_U3291) );
  INV_X1 U8422 ( .A(n6807), .ZN(n6809) );
  OAI222_X1 U8423 ( .A1(n8971), .A2(n6808), .B1(n8969), .B2(n6809), .C1(n8583), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  OAI222_X1 U8424 ( .A1(n8045), .A2(n6810), .B1(n8048), .B2(n6809), .C1(
        P1_U3084), .C2(n9137), .ZN(P1_U3334) );
  XOR2_X1 U8425 ( .A(n6812), .B(n6811), .Z(n6819) );
  AND2_X1 U8426 ( .A1(n9422), .A2(n7053), .ZN(n9777) );
  AOI21_X1 U8427 ( .B1(n9101), .B2(n9123), .A(n6813), .ZN(n6815) );
  NAND2_X1 U8428 ( .A1(n9456), .A2(n9124), .ZN(n6814) );
  OAI211_X1 U8429 ( .C1(n9468), .C2(n6816), .A(n6815), .B(n6814), .ZN(n6817)
         );
  AOI21_X1 U8430 ( .B1(n9464), .B2(n9777), .A(n6817), .ZN(n6818) );
  OAI21_X1 U8431 ( .B1(n6819), .B2(n9460), .A(n6818), .ZN(P1_U3237) );
  INV_X1 U8432 ( .A(n8465), .ZN(n6843) );
  INV_X1 U8433 ( .A(n8467), .ZN(n6820) );
  OAI22_X1 U8434 ( .A1(n8202), .A2(n6820), .B1(n6947), .B2(n9835), .ZN(n6822)
         );
  NAND2_X1 U8435 ( .A1(n6822), .A2(n6821), .ZN(n6824) );
  AOI22_X1 U8436 ( .A1(n9854), .A2(n9898), .B1(n6841), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n6823) );
  OAI211_X1 U8437 ( .C1(n6843), .C2(n8219), .A(n6824), .B(n6823), .ZN(P2_U3234) );
  OR2_X1 U8438 ( .A1(n6825), .A2(n8564), .ZN(n6827) );
  NAND2_X1 U8439 ( .A1(n8461), .A2(n8656), .ZN(n6826) );
  AND2_X1 U8440 ( .A1(n6827), .A2(n6826), .ZN(n7121) );
  INV_X1 U8441 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6828) );
  OAI22_X1 U8442 ( .A1(n8209), .A2(n7121), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6828), .ZN(n6830) );
  NOR2_X1 U8443 ( .A1(n8214), .A2(n9926), .ZN(n6829) );
  AOI211_X1 U8444 ( .C1(n8211), .C2(n7127), .A(n6830), .B(n6829), .ZN(n6836)
         );
  INV_X1 U8445 ( .A(n6831), .ZN(n6834) );
  OAI22_X1 U8446 ( .A1(n8202), .A2(n7016), .B1(n9835), .B2(n6832), .ZN(n6833)
         );
  NAND3_X1 U8447 ( .A1(n7997), .A2(n6834), .A3(n6833), .ZN(n6835) );
  OAI211_X1 U8448 ( .C1(n6837), .C2(n9835), .A(n6836), .B(n6835), .ZN(P2_U3241) );
  NOR2_X1 U8449 ( .A1(n8214), .A2(n9916), .ZN(n6840) );
  OAI22_X1 U8450 ( .A1(n6843), .A2(n9831), .B1(n8219), .B2(n7017), .ZN(n6839)
         );
  AOI211_X1 U8451 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(n6841), .A(n6840), .B(
        n6839), .ZN(n6849) );
  OAI22_X1 U8452 ( .A1(n8202), .A2(n6843), .B1(n9835), .B2(n6842), .ZN(n6847)
         );
  INV_X1 U8453 ( .A(n6844), .ZN(n6845) );
  NAND3_X1 U8454 ( .A1(n6847), .A2(n6846), .A3(n6845), .ZN(n6848) );
  OAI211_X1 U8455 ( .C1(n9835), .C2(n6838), .A(n6849), .B(n6848), .ZN(P2_U3239) );
  INV_X1 U8456 ( .A(n6850), .ZN(n6852) );
  INV_X1 U8457 ( .A(n6858), .ZN(n6851) );
  AOI21_X1 U8458 ( .B1(n6852), .B2(n6851), .A(n4343), .ZN(n6862) );
  INV_X1 U8459 ( .A(n6853), .ZN(n6855) );
  OAI22_X1 U8460 ( .A1(n8214), .A2(n9920), .B1(n8219), .B2(n7016), .ZN(n6854)
         );
  AOI211_X1 U8461 ( .C1(n6856), .C2(n8211), .A(n6855), .B(n6854), .ZN(n6861)
         );
  NOR3_X1 U8462 ( .A1(n8202), .A2(n6858), .A3(n6857), .ZN(n6859) );
  OAI21_X1 U8463 ( .B1(n6859), .B2(n8194), .A(n8463), .ZN(n6860) );
  OAI211_X1 U8464 ( .C1(n6862), .C2(n9835), .A(n6861), .B(n6860), .ZN(P2_U3232) );
  XNOR2_X1 U8465 ( .A(n6865), .B(n6864), .ZN(n6866) );
  XNOR2_X1 U8466 ( .A(n7146), .B(n6866), .ZN(n6873) );
  INV_X1 U8467 ( .A(n7179), .ZN(n7173) );
  NOR2_X1 U8468 ( .A1(n7173), .A2(n9799), .ZN(n9784) );
  INV_X1 U8469 ( .A(n6867), .ZN(n7176) );
  AOI21_X1 U8470 ( .B1(n9101), .B2(n9122), .A(n6868), .ZN(n6870) );
  NAND2_X1 U8471 ( .A1(n9456), .A2(n9676), .ZN(n6869) );
  OAI211_X1 U8472 ( .C1(n9468), .C2(n7176), .A(n6870), .B(n6869), .ZN(n6871)
         );
  AOI21_X1 U8473 ( .B1(n9464), .B2(n9784), .A(n6871), .ZN(n6872) );
  OAI21_X1 U8474 ( .B1(n6873), .B2(n9460), .A(n6872), .ZN(P1_U3211) );
  AND2_X1 U8475 ( .A1(n6875), .A2(n6874), .ZN(n6876) );
  INV_X1 U8476 ( .A(n6878), .ZN(n6879) );
  OAI21_X1 U8477 ( .B1(n8260), .B2(n8403), .A(n7000), .ZN(n6880) );
  AOI222_X1 U8478 ( .A1(n8659), .A2(n6880), .B1(n8464), .B2(n8654), .C1(n8467), 
        .C2(n8656), .ZN(n9906) );
  OAI21_X1 U8479 ( .B1(n6881), .B2(n8679), .A(n9906), .ZN(n6892) );
  OR2_X1 U8480 ( .A1(n6882), .A2(n8569), .ZN(n6911) );
  INV_X1 U8481 ( .A(n6883), .ZN(n7007) );
  AOI21_X1 U8482 ( .B1(n9898), .B2(n6884), .A(n9936), .ZN(n6885) );
  NAND2_X1 U8483 ( .A1(n7007), .A2(n6885), .ZN(n9905) );
  INV_X1 U8484 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6886) );
  OAI22_X1 U8485 ( .A1(n6911), .A2(n9905), .B1(n8688), .B2(n6886), .ZN(n6891)
         );
  NOR2_X1 U8486 ( .A1(n8399), .A2(n7088), .ZN(n6887) );
  AND2_X1 U8487 ( .A1(n8569), .A2(n8255), .ZN(n8242) );
  NAND2_X1 U8488 ( .A1(n8242), .A2(n7088), .ZN(n6913) );
  NAND2_X1 U8489 ( .A1(n7600), .A2(n6913), .ZN(n6888) );
  XOR2_X1 U8490 ( .A(n6889), .B(n8403), .Z(n9904) );
  OAI22_X1 U8491 ( .A1(n9907), .A2(n8700), .B1(n8711), .B2(n9904), .ZN(n6890)
         );
  AOI211_X1 U8492 ( .C1(n8688), .C2(n6892), .A(n6891), .B(n6890), .ZN(n6893)
         );
  INV_X1 U8493 ( .A(n6893), .ZN(P2_U3295) );
  INV_X1 U8494 ( .A(n6911), .ZN(n8703) );
  INV_X1 U8495 ( .A(n8679), .ZN(n8697) );
  AOI22_X1 U8496 ( .A1(n7135), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n6894), .B2(
        n8697), .ZN(n6895) );
  OAI21_X1 U8497 ( .B1(n4425), .B2(n8700), .A(n6895), .ZN(n6898) );
  NOR2_X1 U8498 ( .A1(n6896), .A2(n7135), .ZN(n6897) );
  AOI211_X1 U8499 ( .C1(n6899), .C2(n8703), .A(n6898), .B(n6897), .ZN(n6900)
         );
  OAI21_X1 U8500 ( .B1(n6901), .B2(n8711), .A(n6900), .ZN(P2_U3289) );
  INV_X1 U8501 ( .A(n9853), .ZN(n6904) );
  AOI22_X1 U8502 ( .A1(n7135), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n6902), .B2(
        n8697), .ZN(n6903) );
  OAI21_X1 U8503 ( .B1(n6904), .B2(n8700), .A(n6903), .ZN(n6907) );
  NOR2_X1 U8504 ( .A1(n6905), .A2(n7135), .ZN(n6906) );
  AOI211_X1 U8505 ( .C1(n6908), .C2(n8703), .A(n6907), .B(n6906), .ZN(n6909)
         );
  OAI21_X1 U8506 ( .B1(n8711), .B2(n6910), .A(n6909), .ZN(P2_U3288) );
  NOR2_X2 U8507 ( .A1(n6911), .A2(n9936), .ZN(n8669) );
  INV_X1 U8508 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6912) );
  OAI22_X1 U8509 ( .A1(n8688), .A2(n6912), .B1(n8679), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n6918) );
  INV_X1 U8510 ( .A(n6913), .ZN(n6914) );
  NAND2_X1 U8511 ( .A1(n8688), .A2(n6914), .ZN(n7372) );
  OAI22_X1 U8512 ( .A1(n6916), .A2(n7372), .B1(n6915), .B2(n8700), .ZN(n6917)
         );
  AOI211_X1 U8513 ( .C1(n8669), .C2(n6919), .A(n6918), .B(n6917), .ZN(n6920)
         );
  OAI21_X1 U8514 ( .B1(n7135), .B2(n6921), .A(n6920), .ZN(P2_U3293) );
  INV_X1 U8515 ( .A(n7590), .ZN(n9697) );
  NAND2_X1 U8516 ( .A1(n6923), .A2(n6922), .ZN(n6925) );
  INV_X1 U8517 ( .A(n9727), .ZN(n9700) );
  NAND2_X1 U8518 ( .A1(n9700), .A2(n6718), .ZN(n6924) );
  NAND2_X1 U8519 ( .A1(n6925), .A2(n6924), .ZN(n9692) );
  NAND2_X1 U8520 ( .A1(n6928), .A2(n6926), .ZN(n7737) );
  NAND2_X1 U8521 ( .A1(n9125), .A2(n6927), .ZN(n7055) );
  NAND2_X1 U8522 ( .A1(n7737), .A2(n7055), .ZN(n9698) );
  NAND2_X1 U8523 ( .A1(n9692), .A2(n9698), .ZN(n6930) );
  NAND2_X1 U8524 ( .A1(n6928), .A2(n6927), .ZN(n6929) );
  NAND2_X1 U8525 ( .A1(n9702), .A2(n6934), .ZN(n7736) );
  NAND2_X1 U8526 ( .A1(n9675), .A2(n9764), .ZN(n7738) );
  NAND2_X1 U8527 ( .A1(n7736), .A2(n7738), .ZN(n7907) );
  INV_X1 U8528 ( .A(n7907), .ZN(n6931) );
  XNOR2_X1 U8529 ( .A(n7041), .B(n6931), .ZN(n6943) );
  INV_X1 U8530 ( .A(n6943), .ZN(n9768) );
  NAND2_X1 U8531 ( .A1(n9694), .A2(n6927), .ZN(n9693) );
  NAND2_X1 U8532 ( .A1(n9693), .A2(n6934), .ZN(n6932) );
  NAND2_X1 U8533 ( .A1(n9683), .A2(n6932), .ZN(n9765) );
  AOI22_X1 U8534 ( .A1(n9498), .A2(n6934), .B1(n6933), .B2(n9718), .ZN(n6935)
         );
  OAI21_X1 U8535 ( .B1(n9153), .B2(n9765), .A(n6935), .ZN(n6945) );
  NAND2_X1 U8536 ( .A1(n9700), .A2(n6936), .ZN(n6937) );
  NAND2_X1 U8537 ( .A1(n7056), .A2(n7055), .ZN(n6939) );
  XNOR2_X1 U8538 ( .A(n7907), .B(n6939), .ZN(n6940) );
  NAND2_X1 U8539 ( .A1(n6940), .A2(n9704), .ZN(n6942) );
  AOI22_X1 U8540 ( .A1(n9729), .A2(n9125), .B1(n9124), .B2(n9726), .ZN(n6941)
         );
  OAI211_X1 U8541 ( .C1(n6943), .C2(n9707), .A(n6942), .B(n6941), .ZN(n9766)
         );
  MUX2_X1 U8542 ( .A(n9766), .B(P1_REG2_REG_4__SCAN_IN), .S(n9739), .Z(n6944)
         );
  AOI211_X1 U8543 ( .C1(n9697), .C2(n9768), .A(n6945), .B(n6944), .ZN(n6946)
         );
  INV_X1 U8544 ( .A(n6946), .ZN(P1_U3287) );
  INV_X1 U8545 ( .A(n8260), .ZN(n6948) );
  NAND2_X1 U8546 ( .A1(n8467), .A2(n6947), .ZN(n8256) );
  NAND2_X1 U8547 ( .A1(n6948), .A2(n8256), .ZN(n9900) );
  INV_X1 U8548 ( .A(n9900), .ZN(n6953) );
  AOI22_X1 U8549 ( .A1(n9900), .A2(n8659), .B1(n8654), .B2(n8465), .ZN(n9902)
         );
  INV_X1 U8550 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6949) );
  OAI22_X1 U8551 ( .A1(n7135), .A2(n9902), .B1(n6949), .B2(n8679), .ZN(n6950)
         );
  AOI21_X1 U8552 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n7135), .A(n6950), .ZN(
        n6952) );
  OAI21_X1 U8553 ( .B1(n8669), .B2(n8666), .A(n9898), .ZN(n6951) );
  OAI211_X1 U8554 ( .C1(n6953), .C2(n8711), .A(n6952), .B(n6951), .ZN(P2_U3296) );
  INV_X1 U8555 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n6962) );
  OR2_X1 U8556 ( .A1(n8182), .A2(n9832), .ZN(n8296) );
  NAND2_X1 U8557 ( .A1(n8182), .A2(n9832), .ZN(n8294) );
  INV_X1 U8558 ( .A(n6954), .ZN(n8459) );
  NAND2_X1 U8559 ( .A1(n9853), .A2(n8459), .ZN(n6955) );
  XOR2_X1 U8560 ( .A(n7066), .B(n8411), .Z(n7117) );
  NAND2_X1 U8561 ( .A1(n6957), .A2(n8291), .ZN(n7073) );
  XNOR2_X1 U8562 ( .A(n7073), .B(n8411), .ZN(n6958) );
  INV_X1 U8563 ( .A(n8180), .ZN(n8457) );
  AOI222_X1 U8564 ( .A1(n8659), .A2(n6958), .B1(n8457), .B2(n8654), .C1(n8459), 
        .C2(n8656), .ZN(n7112) );
  INV_X1 U8565 ( .A(n8182), .ZN(n7111) );
  AOI21_X1 U8566 ( .B1(n8182), .B2(n4426), .A(n7078), .ZN(n7115) );
  AOI22_X1 U8567 ( .A1(n7115), .A2(n9912), .B1(n9475), .B2(n8182), .ZN(n6960)
         );
  OAI211_X1 U8568 ( .C1(n7117), .C2(n8785), .A(n7112), .B(n6960), .ZN(n6963)
         );
  NAND2_X1 U8569 ( .A1(n6963), .A2(n9944), .ZN(n6961) );
  OAI21_X1 U8570 ( .B1(n9944), .B2(n6962), .A(n6961), .ZN(P2_U3478) );
  NAND2_X1 U8571 ( .A1(n6963), .A2(n9954), .ZN(n6964) );
  OAI21_X1 U8572 ( .B1(n9954), .B2(n6965), .A(n6964), .ZN(P2_U3529) );
  NOR2_X1 U8573 ( .A1(n6985), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7205) );
  NAND2_X1 U8574 ( .A1(n6985), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7207) );
  INV_X1 U8575 ( .A(n7207), .ZN(n6966) );
  NOR2_X1 U8576 ( .A1(n7205), .A2(n6966), .ZN(n6971) );
  INV_X1 U8577 ( .A(n6967), .ZN(n6970) );
  XOR2_X1 U8578 ( .A(n6971), .B(n7206), .Z(n6989) );
  INV_X1 U8579 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6972) );
  NOR2_X1 U8580 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6972), .ZN(n7330) );
  NAND2_X1 U8581 ( .A1(n6974), .A2(n6973), .ZN(n6975) );
  NAND2_X1 U8582 ( .A1(n6976), .A2(n6975), .ZN(n6979) );
  INV_X1 U8583 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6977) );
  NAND2_X1 U8584 ( .A1(n6979), .A2(n6977), .ZN(n6978) );
  INV_X1 U8585 ( .A(n6978), .ZN(n6982) );
  NAND2_X1 U8586 ( .A1(n6978), .A2(n6985), .ZN(n6981) );
  INV_X1 U8587 ( .A(n6979), .ZN(n6980) );
  NAND2_X1 U8588 ( .A1(n6980), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6984) );
  NAND2_X1 U8589 ( .A1(n6981), .A2(n6984), .ZN(n7217) );
  NOR3_X1 U8590 ( .A1(n9862), .A2(n6982), .A3(n7217), .ZN(n6983) );
  AOI211_X1 U8591 ( .C1(n9870), .C2(P2_ADDR_REG_13__SCAN_IN), .A(n7330), .B(
        n6983), .ZN(n6988) );
  AOI21_X1 U8592 ( .B1(n7217), .B2(n6984), .A(n9862), .ZN(n6986) );
  OAI21_X1 U8593 ( .B1(n6986), .B2(n9876), .A(n6985), .ZN(n6987) );
  OAI211_X1 U8594 ( .C1(n6989), .C2(n8490), .A(n6988), .B(n6987), .ZN(P2_U3258) );
  INV_X1 U8595 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6991) );
  INV_X1 U8596 ( .A(n6990), .ZN(n7989) );
  OAI22_X1 U8597 ( .A1(n8688), .A2(n6991), .B1(n7989), .B2(n8679), .ZN(n6992)
         );
  AOI21_X1 U8598 ( .B1(n6993), .B2(n8703), .A(n6992), .ZN(n6994) );
  OAI21_X1 U8599 ( .B1(n6995), .B2(n8700), .A(n6994), .ZN(n6996) );
  AOI21_X1 U8600 ( .B1(n8662), .B2(n6997), .A(n6996), .ZN(n6998) );
  OAI21_X1 U8601 ( .B1(n7135), .B2(n6999), .A(n6998), .ZN(P2_U3291) );
  NAND3_X1 U8602 ( .A1(n7000), .A2(n8273), .A3(n8402), .ZN(n7001) );
  NAND2_X1 U8603 ( .A1(n7002), .A2(n7001), .ZN(n7003) );
  AOI222_X1 U8604 ( .A1(n8659), .A2(n7003), .B1(n8463), .B2(n8654), .C1(n8465), 
        .C2(n8656), .ZN(n9915) );
  OAI22_X1 U8605 ( .A1(n6205), .A2(n8688), .B1(n6244), .B2(n8679), .ZN(n7004)
         );
  INV_X1 U8606 ( .A(n7004), .ZN(n7011) );
  XNOR2_X1 U8607 ( .A(n7005), .B(n8402), .ZN(n9918) );
  INV_X1 U8608 ( .A(n9916), .ZN(n7006) );
  NAND2_X1 U8609 ( .A1(n7007), .A2(n7006), .ZN(n9913) );
  NAND3_X1 U8610 ( .A1(n8669), .A2(n9911), .A3(n9913), .ZN(n7008) );
  OAI21_X1 U8611 ( .B1(n9916), .B2(n8700), .A(n7008), .ZN(n7009) );
  AOI21_X1 U8612 ( .B1(n8662), .B2(n9918), .A(n7009), .ZN(n7010) );
  OAI211_X1 U8613 ( .C1(n7135), .C2(n9915), .A(n7011), .B(n7010), .ZN(P2_U3294) );
  NAND2_X1 U8614 ( .A1(n7013), .A2(n7012), .ZN(n7014) );
  XNOR2_X1 U8615 ( .A(n7014), .B(n8406), .ZN(n7015) );
  OAI222_X1 U8616 ( .A1(n8562), .A2(n7017), .B1(n8564), .B2(n7016), .C1(n7015), 
        .C2(n8707), .ZN(n9922) );
  INV_X1 U8617 ( .A(n9922), .ZN(n7027) );
  OAI22_X1 U8618 ( .A1(n6206), .A2(n8688), .B1(n7018), .B2(n8679), .ZN(n7022)
         );
  INV_X1 U8619 ( .A(n8669), .ZN(n8621) );
  OAI21_X1 U8620 ( .B1(n9920), .B2(n7020), .A(n7019), .ZN(n9921) );
  NOR2_X1 U8621 ( .A1(n8621), .A2(n9921), .ZN(n7021) );
  AOI211_X1 U8622 ( .C1(n8666), .C2(n4449), .A(n7022), .B(n7021), .ZN(n7026)
         );
  OAI21_X1 U8623 ( .B1(n7024), .B2(n8406), .A(n7023), .ZN(n9924) );
  NAND2_X1 U8624 ( .A1(n9924), .A2(n8662), .ZN(n7025) );
  OAI211_X1 U8625 ( .C1(n7027), .C2(n7135), .A(n7026), .B(n7025), .ZN(P2_U3292) );
  OR2_X1 U8626 ( .A1(n7146), .A2(n7028), .ZN(n7030) );
  NAND2_X1 U8627 ( .A1(n7030), .A2(n7029), .ZN(n7034) );
  XNOR2_X1 U8628 ( .A(n7032), .B(n7031), .ZN(n7033) );
  XNOR2_X1 U8629 ( .A(n7034), .B(n7033), .ZN(n7040) );
  NAND2_X1 U8630 ( .A1(n7194), .A2(n9422), .ZN(n9792) );
  NOR2_X1 U8631 ( .A1(n9792), .A2(n9026), .ZN(n7038) );
  INV_X1 U8632 ( .A(n9123), .ZN(n7093) );
  NAND2_X1 U8633 ( .A1(n9101), .A2(n9121), .ZN(n7035) );
  OAI211_X1 U8634 ( .C1(n9104), .C2(n7093), .A(n7036), .B(n7035), .ZN(n7037)
         );
  AOI211_X1 U8635 ( .C1(n9099), .C2(n7103), .A(n7038), .B(n7037), .ZN(n7039)
         );
  OAI21_X1 U8636 ( .B1(n7040), .B2(n9460), .A(n7039), .ZN(P1_U3219) );
  NAND2_X1 U8637 ( .A1(n9702), .A2(n9764), .ZN(n7042) );
  INV_X1 U8638 ( .A(n9124), .ZN(n7043) );
  NAND2_X1 U8639 ( .A1(n7043), .A2(n9687), .ZN(n7741) );
  INV_X1 U8640 ( .A(n9687), .ZN(n7044) );
  NAND2_X1 U8641 ( .A1(n9124), .A2(n7044), .ZN(n7743) );
  NAND2_X1 U8642 ( .A1(n9124), .A2(n9687), .ZN(n7045) );
  INV_X1 U8643 ( .A(n7048), .ZN(n7047) );
  INV_X1 U8644 ( .A(n9676), .ZN(n7090) );
  INV_X1 U8645 ( .A(n7909), .ZN(n7046) );
  NAND2_X1 U8646 ( .A1(n7048), .A2(n7909), .ZN(n7049) );
  AND2_X1 U8647 ( .A1(n7092), .A2(n7049), .ZN(n7062) );
  INV_X1 U8648 ( .A(n7062), .ZN(n9782) );
  INV_X1 U8649 ( .A(n7174), .ZN(n7051) );
  NAND2_X1 U8650 ( .A1(n9684), .A2(n7053), .ZN(n7050) );
  NAND2_X1 U8651 ( .A1(n7051), .A2(n7050), .ZN(n9779) );
  AOI22_X1 U8652 ( .A1(n9498), .A2(n7053), .B1(n7052), .B2(n9718), .ZN(n7054)
         );
  OAI21_X1 U8653 ( .B1(n9779), .B2(n9153), .A(n7054), .ZN(n7064) );
  NAND2_X1 U8654 ( .A1(n7056), .A2(n7744), .ZN(n7057) );
  INV_X1 U8655 ( .A(n7741), .ZN(n7058) );
  OAI21_X1 U8656 ( .B1(n7909), .B2(n7798), .A(n7794), .ZN(n7059) );
  NAND2_X1 U8657 ( .A1(n7059), .A2(n9704), .ZN(n7061) );
  AOI22_X1 U8658 ( .A1(n9729), .A2(n9124), .B1(n9123), .B2(n9726), .ZN(n7060)
         );
  OAI211_X1 U8659 ( .C1(n7062), .C2(n9707), .A(n7061), .B(n7060), .ZN(n9780)
         );
  MUX2_X1 U8660 ( .A(n9780), .B(P1_REG2_REG_6__SCAN_IN), .S(n9739), .Z(n7063)
         );
  AOI211_X1 U8661 ( .C1(n9697), .C2(n9782), .A(n7064), .B(n7063), .ZN(n7065)
         );
  INV_X1 U8662 ( .A(n7065), .ZN(P1_U3285) );
  INV_X1 U8663 ( .A(n7066), .ZN(n7068) );
  INV_X1 U8664 ( .A(n8411), .ZN(n7067) );
  INV_X1 U8665 ( .A(n9832), .ZN(n8458) );
  OR2_X1 U8666 ( .A1(n8182), .A2(n8458), .ZN(n7069) );
  OR2_X1 U8667 ( .A1(n9840), .A2(n8180), .ZN(n8298) );
  NAND2_X1 U8668 ( .A1(n9840), .A2(n8180), .ZN(n8300) );
  NAND2_X1 U8669 ( .A1(n7071), .A2(n8413), .ZN(n7072) );
  NAND2_X1 U8670 ( .A1(n7237), .A2(n7072), .ZN(n9933) );
  XNOR2_X1 U8671 ( .A(n4347), .B(n8413), .ZN(n7075) );
  OAI22_X1 U8672 ( .A1(n7345), .A2(n8564), .B1(n9832), .B2(n8562), .ZN(n7074)
         );
  AOI21_X1 U8673 ( .B1(n7075), .B2(n8659), .A(n7074), .ZN(n7076) );
  OAI21_X1 U8674 ( .B1(n9933), .B2(n7600), .A(n7076), .ZN(n9938) );
  NAND2_X1 U8675 ( .A1(n9938), .A2(n8688), .ZN(n7083) );
  INV_X1 U8676 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7077) );
  OAI22_X1 U8677 ( .A1(n8688), .A2(n7077), .B1(n9842), .B2(n8679), .ZN(n7081)
         );
  INV_X1 U8678 ( .A(n9840), .ZN(n9935) );
  NAND2_X1 U8679 ( .A1(n7078), .A2(n9935), .ZN(n7252) );
  OR2_X1 U8680 ( .A1(n7078), .A2(n9935), .ZN(n7079) );
  NAND2_X1 U8681 ( .A1(n7252), .A2(n7079), .ZN(n9937) );
  NOR2_X1 U8682 ( .A1(n9937), .A2(n8621), .ZN(n7080) );
  AOI211_X1 U8683 ( .C1(n8666), .C2(n9840), .A(n7081), .B(n7080), .ZN(n7082)
         );
  OAI211_X1 U8684 ( .C1(n9933), .C2(n7372), .A(n7083), .B(n7082), .ZN(P2_U3286) );
  INV_X1 U8685 ( .A(n7084), .ZN(n8042) );
  INV_X1 U8686 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7085) );
  OAI222_X1 U8687 ( .A1(n8969), .A2(n8042), .B1(P2_U3152), .B2(n8436), .C1(
        n7085), .C2(n8971), .ZN(P2_U3337) );
  INV_X1 U8688 ( .A(n7086), .ZN(n7702) );
  OAI222_X1 U8689 ( .A1(n8975), .A2(n7702), .B1(n10007), .B2(n7088), .C1(n7087), .C2(n8971), .ZN(P2_U3338) );
  NAND2_X1 U8690 ( .A1(n7090), .A2(n7089), .ZN(n7091) );
  NAND2_X1 U8691 ( .A1(n7093), .A2(n7179), .ZN(n7799) );
  NAND2_X1 U8692 ( .A1(n7173), .A2(n9123), .ZN(n7797) );
  NAND2_X1 U8693 ( .A1(n7799), .A2(n7797), .ZN(n7912) );
  INV_X1 U8694 ( .A(n7098), .ZN(n7097) );
  INV_X1 U8695 ( .A(n7194), .ZN(n7094) );
  NAND2_X1 U8696 ( .A1(n7094), .A2(n9122), .ZN(n7803) );
  INV_X1 U8697 ( .A(n9122), .ZN(n7095) );
  NAND2_X1 U8698 ( .A1(n7095), .A2(n7194), .ZN(n7804) );
  NAND2_X1 U8699 ( .A1(n7098), .A2(n7911), .ZN(n7099) );
  NAND2_X1 U8700 ( .A1(n7196), .A2(n7099), .ZN(n9791) );
  INV_X1 U8701 ( .A(n7912), .ZN(n7183) );
  NAND2_X1 U8702 ( .A1(n7948), .A2(n7183), .ZN(n7182) );
  NAND2_X1 U8703 ( .A1(n7182), .A2(n7799), .ZN(n7188) );
  XNOR2_X1 U8704 ( .A(n7188), .B(n7911), .ZN(n7100) );
  NAND2_X1 U8705 ( .A1(n7100), .A2(n9704), .ZN(n7102) );
  AOI22_X1 U8706 ( .A1(n9729), .A2(n9123), .B1(n9121), .B2(n9726), .ZN(n7101)
         );
  OAI211_X1 U8707 ( .C1(n9707), .C2(n9791), .A(n7102), .B(n7101), .ZN(n9794)
         );
  NAND2_X1 U8708 ( .A1(n9794), .A2(n9737), .ZN(n7109) );
  INV_X1 U8709 ( .A(n7103), .ZN(n7104) );
  OAI22_X1 U8710 ( .A1(n9737), .A2(n8918), .B1(n7104), .B2(n9709), .ZN(n7107)
         );
  NAND2_X1 U8711 ( .A1(n7172), .A2(n7194), .ZN(n7105) );
  NAND2_X1 U8712 ( .A1(n7197), .A2(n7105), .ZN(n9793) );
  NOR2_X1 U8713 ( .A1(n9793), .A2(n9153), .ZN(n7106) );
  AOI211_X1 U8714 ( .C1(n9498), .C2(n7194), .A(n7107), .B(n7106), .ZN(n7108)
         );
  OAI211_X1 U8715 ( .C1(n9791), .C2(n7590), .A(n7109), .B(n7108), .ZN(P1_U3283) );
  AOI22_X1 U8716 ( .A1(n7135), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n8177), .B2(
        n8697), .ZN(n7110) );
  OAI21_X1 U8717 ( .B1(n7111), .B2(n8700), .A(n7110), .ZN(n7114) );
  NOR2_X1 U8718 ( .A1(n7112), .A2(n7135), .ZN(n7113) );
  AOI211_X1 U8719 ( .C1(n7115), .C2(n8669), .A(n7114), .B(n7113), .ZN(n7116)
         );
  OAI21_X1 U8720 ( .B1(n8711), .B2(n7117), .A(n7116), .ZN(P2_U3287) );
  XNOR2_X1 U8721 ( .A(n7119), .B(n7118), .ZN(n7120) );
  NAND2_X1 U8722 ( .A1(n7120), .A2(n8659), .ZN(n7122) );
  NAND2_X1 U8723 ( .A1(n7122), .A2(n7121), .ZN(n9928) );
  INV_X1 U8724 ( .A(n9928), .ZN(n7134) );
  OAI21_X1 U8725 ( .B1(n7124), .B2(n8408), .A(n7123), .ZN(n9930) );
  OAI21_X1 U8726 ( .B1(n7126), .B2(n9926), .A(n7125), .ZN(n9927) );
  INV_X1 U8727 ( .A(n7127), .ZN(n7128) );
  OAI22_X1 U8728 ( .A1(n8688), .A2(n6207), .B1(n7128), .B2(n8679), .ZN(n7129)
         );
  AOI21_X1 U8729 ( .B1(n8666), .B2(n7130), .A(n7129), .ZN(n7131) );
  OAI21_X1 U8730 ( .B1(n8621), .B2(n9927), .A(n7131), .ZN(n7132) );
  AOI21_X1 U8731 ( .B1(n9930), .B2(n8662), .A(n7132), .ZN(n7133) );
  OAI21_X1 U8732 ( .B1(n7135), .B2(n7134), .A(n7133), .ZN(P2_U3290) );
  NAND2_X1 U8733 ( .A1(n4346), .A2(n7136), .ZN(n7137) );
  XNOR2_X1 U8734 ( .A(n7138), .B(n7137), .ZN(n7144) );
  INV_X1 U8735 ( .A(n9121), .ZN(n7189) );
  NAND2_X1 U8736 ( .A1(n9099), .A2(n7310), .ZN(n7141) );
  AOI21_X1 U8737 ( .B1(n9101), .B2(n9455), .A(n7139), .ZN(n7140) );
  OAI211_X1 U8738 ( .C1(n7189), .C2(n9104), .A(n7141), .B(n7140), .ZN(n7142)
         );
  AOI21_X1 U8739 ( .B1(n9107), .B2(n7402), .A(n7142), .ZN(n7143) );
  OAI21_X1 U8740 ( .B1(n7144), .B2(n9460), .A(n7143), .ZN(P1_U3215) );
  OR2_X1 U8741 ( .A1(n7146), .A2(n7145), .ZN(n7149) );
  NAND2_X1 U8742 ( .A1(n7149), .A2(n7147), .ZN(n7151) );
  AND2_X1 U8743 ( .A1(n7148), .A2(n7149), .ZN(n7150) );
  AOI21_X1 U8744 ( .B1(n7152), .B2(n7151), .A(n7150), .ZN(n7158) );
  INV_X1 U8745 ( .A(n7199), .ZN(n7155) );
  NAND2_X1 U8746 ( .A1(n9456), .A2(n9122), .ZN(n7154) );
  AND2_X1 U8747 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9609) );
  AOI21_X1 U8748 ( .B1(n9101), .B2(n9120), .A(n9609), .ZN(n7153) );
  OAI211_X1 U8749 ( .C1(n9468), .C2(n7155), .A(n7154), .B(n7153), .ZN(n7156)
         );
  AOI21_X1 U8750 ( .B1(n9107), .B2(n7315), .A(n7156), .ZN(n7157) );
  OAI21_X1 U8751 ( .B1(n7158), .B2(n9460), .A(n7157), .ZN(P1_U3229) );
  INV_X1 U8752 ( .A(n7159), .ZN(n7160) );
  AOI21_X1 U8753 ( .B1(n9833), .B2(n7160), .A(n9835), .ZN(n7163) );
  NOR3_X1 U8754 ( .A1(n7161), .A2(n8202), .A3(n8180), .ZN(n7162) );
  OAI21_X1 U8755 ( .B1(n7163), .B2(n7162), .A(n7344), .ZN(n7169) );
  INV_X1 U8756 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7164) );
  OAI22_X1 U8757 ( .A1(n9860), .A2(n7165), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7164), .ZN(n7167) );
  OAI22_X1 U8758 ( .A1(n8180), .A2(n9831), .B1(n8219), .B2(n7328), .ZN(n7166)
         );
  AOI211_X1 U8759 ( .C1(n9854), .C2(n7265), .A(n7167), .B(n7166), .ZN(n7168)
         );
  NAND2_X1 U8760 ( .A1(n7169), .A2(n7168), .ZN(P2_U3238) );
  AND2_X1 U8761 ( .A1(n7170), .A2(n8999), .ZN(n9682) );
  INV_X1 U8762 ( .A(n9329), .ZN(n9312) );
  XNOR2_X1 U8763 ( .A(n7171), .B(n7912), .ZN(n9789) );
  OAI211_X1 U8764 ( .C1(n7174), .C2(n7173), .A(n9717), .B(n7172), .ZN(n9785)
         );
  NOR2_X1 U8765 ( .A1(n7175), .A2(n9721), .ZN(n7677) );
  INV_X1 U8766 ( .A(n7677), .ZN(n7181) );
  OAI22_X1 U8767 ( .A1(n9737), .A2(n7177), .B1(n7176), .B2(n9709), .ZN(n7178)
         );
  AOI21_X1 U8768 ( .B1(n9498), .B2(n7179), .A(n7178), .ZN(n7180) );
  OAI21_X1 U8769 ( .B1(n9785), .B2(n7181), .A(n7180), .ZN(n7186) );
  OAI21_X1 U8770 ( .B1(n7183), .B2(n7948), .A(n7182), .ZN(n7184) );
  AOI222_X1 U8771 ( .A1(n9704), .A2(n7184), .B1(n9676), .B2(n9729), .C1(n9122), 
        .C2(n9726), .ZN(n9787) );
  NOR2_X1 U8772 ( .A1(n9787), .A2(n9739), .ZN(n7185) );
  AOI211_X1 U8773 ( .C1(n9312), .C2(n9789), .A(n7186), .B(n7185), .ZN(n7187)
         );
  INV_X1 U8774 ( .A(n7187), .ZN(P1_U3284) );
  INV_X1 U8775 ( .A(n7804), .ZN(n7813) );
  NAND2_X1 U8776 ( .A1(n7386), .A2(n7803), .ZN(n7190) );
  OR2_X1 U8777 ( .A1(n7189), .A2(n7315), .ZN(n7807) );
  NAND2_X1 U8778 ( .A1(n7315), .A2(n7189), .ZN(n7805) );
  NAND2_X1 U8779 ( .A1(n7807), .A2(n7805), .ZN(n7913) );
  XNOR2_X1 U8780 ( .A(n7190), .B(n7913), .ZN(n7191) );
  NAND2_X1 U8781 ( .A1(n7191), .A2(n9704), .ZN(n7193) );
  AOI22_X1 U8782 ( .A1(n9729), .A2(n9122), .B1(n9120), .B2(n9726), .ZN(n7192)
         );
  NAND2_X1 U8783 ( .A1(n7193), .A2(n7192), .ZN(n9803) );
  INV_X1 U8784 ( .A(n9803), .ZN(n7204) );
  NAND2_X1 U8785 ( .A1(n7194), .A2(n9122), .ZN(n7195) );
  XOR2_X1 U8786 ( .A(n7314), .B(n7913), .Z(n9806) );
  INV_X1 U8787 ( .A(n7315), .ZN(n9800) );
  INV_X1 U8788 ( .A(n7197), .ZN(n7198) );
  INV_X1 U8789 ( .A(n7308), .ZN(n7309) );
  OAI21_X1 U8790 ( .B1(n9800), .B2(n7198), .A(n7309), .ZN(n9802) );
  AOI22_X1 U8791 ( .A1(n9739), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7199), .B2(
        n9718), .ZN(n7201) );
  NAND2_X1 U8792 ( .A1(n9498), .A2(n7315), .ZN(n7200) );
  OAI211_X1 U8793 ( .C1(n9802), .C2(n9153), .A(n7201), .B(n7200), .ZN(n7202)
         );
  AOI21_X1 U8794 ( .B1(n9806), .B2(n9312), .A(n7202), .ZN(n7203) );
  OAI21_X1 U8795 ( .B1(n7204), .B2(n9739), .A(n7203), .ZN(P1_U3282) );
  INV_X1 U8796 ( .A(n7211), .ZN(n7213) );
  INV_X1 U8797 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7441) );
  OR2_X1 U8798 ( .A1(n7219), .A2(n7441), .ZN(n7209) );
  NAND2_X1 U8799 ( .A1(n7219), .A2(n7441), .ZN(n7208) );
  NAND2_X1 U8800 ( .A1(n7209), .A2(n7208), .ZN(n7212) );
  INV_X1 U8801 ( .A(n7212), .ZN(n7210) );
  OAI21_X1 U8802 ( .B1(n7213), .B2(n7212), .A(n7411), .ZN(n7214) );
  NAND2_X1 U8803 ( .A1(n7214), .A2(n9879), .ZN(n7225) );
  NOR2_X1 U8804 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8820), .ZN(n7223) );
  NOR2_X1 U8805 ( .A1(n7219), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7215) );
  INV_X1 U8806 ( .A(n7415), .ZN(n7221) );
  INV_X1 U8807 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7218) );
  NAND2_X1 U8808 ( .A1(n7219), .A2(n7218), .ZN(n7216) );
  OAI211_X1 U8809 ( .C1(n7219), .C2(n7218), .A(n7217), .B(n7216), .ZN(n7220)
         );
  AOI21_X1 U8810 ( .B1(n7221), .B2(n7220), .A(n9862), .ZN(n7222) );
  AOI211_X1 U8811 ( .C1(n9870), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n7223), .B(
        n7222), .ZN(n7224) );
  OAI211_X1 U8812 ( .C1(n9861), .C2(n7416), .A(n7225), .B(n7224), .ZN(P2_U3259) );
  INV_X1 U8813 ( .A(n7226), .ZN(n8044) );
  OAI222_X1 U8814 ( .A1(n8971), .A2(n7227), .B1(n8969), .B2(n8044), .C1(n8241), 
        .C2(n10007), .ZN(P2_U3336) );
  OAI211_X1 U8815 ( .C1(n7230), .C2(n7229), .A(n7228), .B(n9086), .ZN(n7235)
         );
  INV_X1 U8816 ( .A(n9120), .ZN(n9513) );
  AOI21_X1 U8817 ( .B1(n9101), .B2(n9119), .A(n7231), .ZN(n7232) );
  OAI21_X1 U8818 ( .B1(n9513), .B2(n9104), .A(n7232), .ZN(n7233) );
  AOI21_X1 U8819 ( .B1(n9518), .B2(n9099), .A(n7233), .ZN(n7234) );
  OAI211_X1 U8820 ( .C1(n9535), .C2(n9095), .A(n7235), .B(n7234), .ZN(P1_U3234) );
  OR2_X1 U8821 ( .A1(n7361), .A2(n7328), .ZN(n8416) );
  NAND2_X1 U8822 ( .A1(n7361), .A2(n7328), .ZN(n8417) );
  NAND2_X1 U8823 ( .A1(n9840), .A2(n8457), .ZN(n7236) );
  OR2_X1 U8824 ( .A1(n7265), .A2(n7345), .ZN(n8305) );
  NAND2_X1 U8825 ( .A1(n7265), .A2(n7345), .ZN(n8308) );
  NAND2_X1 U8826 ( .A1(n8305), .A2(n8308), .ZN(n8414) );
  INV_X1 U8827 ( .A(n7345), .ZN(n9827) );
  NAND2_X1 U8828 ( .A1(n7265), .A2(n9827), .ZN(n7238) );
  XOR2_X1 U8829 ( .A(n7365), .B(n7362), .Z(n7339) );
  INV_X1 U8830 ( .A(n8300), .ZN(n7239) );
  AND2_X1 U8831 ( .A1(n8305), .A2(n8298), .ZN(n8301) );
  NAND2_X1 U8832 ( .A1(n7240), .A2(n8308), .ZN(n7366) );
  XOR2_X1 U8833 ( .A(n7366), .B(n7365), .Z(n7241) );
  INV_X1 U8834 ( .A(n7434), .ZN(n8455) );
  AOI22_X1 U8835 ( .A1(n8654), .A2(n8455), .B1(n9827), .B2(n8656), .ZN(n7351)
         );
  OAI21_X1 U8836 ( .B1(n7241), .B2(n8707), .A(n7351), .ZN(n7336) );
  INV_X1 U8837 ( .A(n7373), .ZN(n7242) );
  AOI211_X1 U8838 ( .C1(n7361), .C2(n7251), .A(n9936), .B(n7242), .ZN(n7337)
         );
  NAND2_X1 U8839 ( .A1(n7337), .A2(n8703), .ZN(n7244) );
  AOI22_X1 U8840 ( .A1(n7135), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n4841), .B2(
        n8697), .ZN(n7243) );
  OAI211_X1 U8841 ( .C1(n4548), .C2(n8700), .A(n7244), .B(n7243), .ZN(n7245)
         );
  AOI21_X1 U8842 ( .B1(n7336), .B2(n8688), .A(n7245), .ZN(n7246) );
  OAI21_X1 U8843 ( .B1(n7339), .B2(n8711), .A(n7246), .ZN(P2_U3284) );
  INV_X1 U8844 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7255) );
  XNOR2_X1 U8845 ( .A(n4371), .B(n8414), .ZN(n7274) );
  NAND2_X1 U8846 ( .A1(n7248), .A2(n8298), .ZN(n7249) );
  XNOR2_X1 U8847 ( .A(n7249), .B(n8414), .ZN(n7250) );
  INV_X1 U8848 ( .A(n7328), .ZN(n8456) );
  AOI222_X1 U8849 ( .A1(n8659), .A2(n7250), .B1(n8456), .B2(n8654), .C1(n8457), 
        .C2(n8656), .ZN(n7269) );
  AOI21_X1 U8850 ( .B1(n7265), .B2(n7252), .A(n4549), .ZN(n7272) );
  AOI22_X1 U8851 ( .A1(n7272), .A2(n9912), .B1(n9475), .B2(n7265), .ZN(n7253)
         );
  OAI211_X1 U8852 ( .C1(n7274), .C2(n8785), .A(n7269), .B(n7253), .ZN(n7256)
         );
  NAND2_X1 U8853 ( .A1(n7256), .A2(n9944), .ZN(n7254) );
  OAI21_X1 U8854 ( .B1(n9944), .B2(n7255), .A(n7254), .ZN(P2_U3484) );
  NAND2_X1 U8855 ( .A1(n7256), .A2(n9954), .ZN(n7257) );
  OAI21_X1 U8856 ( .B1(n9954), .B2(n6688), .A(n7257), .ZN(P2_U3531) );
  INV_X1 U8857 ( .A(n7261), .ZN(n7260) );
  AOI21_X1 U8858 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n8967), .A(n7258), .ZN(
        n7259) );
  OAI21_X1 U8859 ( .B1(n7260), .B2(n8969), .A(n7259), .ZN(P2_U3335) );
  NAND2_X1 U8860 ( .A1(n7261), .A2(n9447), .ZN(n7263) );
  NOR2_X1 U8861 ( .A1(n7262), .A2(P1_U3084), .ZN(n7978) );
  INV_X1 U8862 ( .A(n7978), .ZN(n7984) );
  OAI211_X1 U8863 ( .C1(n7264), .C2(n9444), .A(n7263), .B(n7984), .ZN(P1_U3330) );
  INV_X1 U8864 ( .A(n7265), .ZN(n7268) );
  AOI22_X1 U8865 ( .A1(n7135), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7266), .B2(
        n8697), .ZN(n7267) );
  OAI21_X1 U8866 ( .B1(n7268), .B2(n8700), .A(n7267), .ZN(n7271) );
  NOR2_X1 U8867 ( .A1(n7269), .A2(n7135), .ZN(n7270) );
  AOI211_X1 U8868 ( .C1(n7272), .C2(n8669), .A(n7271), .B(n7270), .ZN(n7273)
         );
  OAI21_X1 U8869 ( .B1(n8711), .B2(n7274), .A(n7273), .ZN(P2_U3285) );
  INV_X1 U8870 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n9992) );
  NOR2_X1 U8871 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7275) );
  AOI21_X1 U8872 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7275), .ZN(n9961) );
  NOR2_X1 U8873 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(P2_ADDR_REG_16__SCAN_IN), 
        .ZN(n7276) );
  AOI21_X1 U8874 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n7276), .ZN(n9964) );
  NOR2_X1 U8875 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7277) );
  AOI21_X1 U8876 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7277), .ZN(n9967) );
  NOR2_X1 U8877 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7278) );
  AOI21_X1 U8878 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7278), .ZN(n9970) );
  NOR2_X1 U8879 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7279) );
  AOI21_X1 U8880 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7279), .ZN(n9973) );
  NOR2_X1 U8881 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7285) );
  XNOR2_X1 U8882 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10004) );
  NAND2_X1 U8883 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7283) );
  XOR2_X1 U8884 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10002) );
  NAND2_X1 U8885 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7281) );
  XOR2_X1 U8886 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n9998) );
  AOI21_X1 U8887 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9955) );
  NAND3_X1 U8888 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9957) );
  OAI21_X1 U8889 ( .B1(n9955), .B2(n6199), .A(n9957), .ZN(n9997) );
  NAND2_X1 U8890 ( .A1(n9998), .A2(n9997), .ZN(n7280) );
  NAND2_X1 U8891 ( .A1(n7281), .A2(n7280), .ZN(n10001) );
  NAND2_X1 U8892 ( .A1(n10002), .A2(n10001), .ZN(n7282) );
  NAND2_X1 U8893 ( .A1(n7283), .A2(n7282), .ZN(n10003) );
  NOR2_X1 U8894 ( .A1(n10004), .A2(n10003), .ZN(n7284) );
  NOR2_X1 U8895 ( .A1(n7285), .A2(n7284), .ZN(n7286) );
  NOR2_X1 U8896 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7286), .ZN(n9988) );
  AND2_X1 U8897 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7286), .ZN(n9987) );
  NOR2_X1 U8898 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n9987), .ZN(n7287) );
  NOR2_X1 U8899 ( .A1(n9988), .A2(n7287), .ZN(n7288) );
  NAND2_X1 U8900 ( .A1(n7288), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7290) );
  XOR2_X1 U8901 ( .A(n7288), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n9986) );
  NAND2_X1 U8902 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n9986), .ZN(n7289) );
  NAND2_X1 U8903 ( .A1(n7290), .A2(n7289), .ZN(n7291) );
  NAND2_X1 U8904 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7291), .ZN(n7293) );
  XOR2_X1 U8905 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7291), .Z(n10000) );
  NAND2_X1 U8906 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10000), .ZN(n7292) );
  NAND2_X1 U8907 ( .A1(n7293), .A2(n7292), .ZN(n7294) );
  NAND2_X1 U8908 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7294), .ZN(n7296) );
  XOR2_X1 U8909 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7294), .Z(n9984) );
  NAND2_X1 U8910 ( .A1(n9984), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7295) );
  NAND2_X1 U8911 ( .A1(n7296), .A2(n7295), .ZN(n7297) );
  AND2_X1 U8912 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7297), .ZN(n7298) );
  INV_X1 U8913 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9996) );
  XNOR2_X1 U8914 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7297), .ZN(n9995) );
  NAND2_X1 U8915 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7299) );
  OAI21_X1 U8916 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n7299), .ZN(n9981) );
  NAND2_X1 U8917 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7300) );
  OAI21_X1 U8918 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7300), .ZN(n9978) );
  AOI21_X1 U8919 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9977), .ZN(n9976) );
  NOR2_X1 U8920 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7301) );
  AOI21_X1 U8921 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7301), .ZN(n9975) );
  NAND2_X1 U8922 ( .A1(n9976), .A2(n9975), .ZN(n9974) );
  OAI21_X1 U8923 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9974), .ZN(n9972) );
  NAND2_X1 U8924 ( .A1(n9973), .A2(n9972), .ZN(n9971) );
  OAI21_X1 U8925 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9971), .ZN(n9969) );
  NAND2_X1 U8926 ( .A1(n9970), .A2(n9969), .ZN(n9968) );
  OAI21_X1 U8927 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9968), .ZN(n9966) );
  NAND2_X1 U8928 ( .A1(n9967), .A2(n9966), .ZN(n9965) );
  OAI21_X1 U8929 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9965), .ZN(n9963) );
  NAND2_X1 U8930 ( .A1(n9964), .A2(n9963), .ZN(n9962) );
  OAI21_X1 U8931 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9962), .ZN(n9960) );
  NAND2_X1 U8932 ( .A1(n9961), .A2(n9960), .ZN(n9959) );
  OAI21_X1 U8933 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9959), .ZN(n9991) );
  NOR2_X1 U8934 ( .A1(n9992), .A2(n9991), .ZN(n7302) );
  NAND2_X1 U8935 ( .A1(n9992), .A2(n9991), .ZN(n9990) );
  OAI21_X1 U8936 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7302), .A(n9990), .ZN(
        n7304) );
  XNOR2_X1 U8937 ( .A(n4868), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7303) );
  XNOR2_X1 U8938 ( .A(n7304), .B(n7303), .ZN(ADD_1071_U4) );
  OR2_X1 U8939 ( .A1(n7402), .A2(n9513), .ZN(n7821) );
  NAND2_X1 U8940 ( .A1(n7402), .A2(n9513), .ZN(n7808) );
  AND2_X1 U8941 ( .A1(n7807), .A2(n7803), .ZN(n7812) );
  INV_X1 U8942 ( .A(n7805), .ZN(n7305) );
  AOI21_X1 U8943 ( .B1(n7386), .B2(n7812), .A(n7305), .ZN(n7306) );
  XOR2_X1 U8944 ( .A(n7915), .B(n7306), .Z(n7307) );
  AOI222_X1 U8945 ( .A1(n9704), .A2(n7307), .B1(n9455), .B2(n9726), .C1(n9121), 
        .C2(n9729), .ZN(n7404) );
  INV_X1 U8946 ( .A(n7402), .ZN(n7312) );
  AOI211_X1 U8947 ( .C1(n7402), .C2(n7309), .A(n9801), .B(n9507), .ZN(n7401)
         );
  AOI22_X1 U8948 ( .A1(n9739), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7310), .B2(
        n9718), .ZN(n7311) );
  OAI21_X1 U8949 ( .B1(n7312), .B2(n9710), .A(n7311), .ZN(n7323) );
  OR2_X1 U8950 ( .A1(n7315), .A2(n9121), .ZN(n7313) );
  NAND2_X1 U8951 ( .A1(n7315), .A2(n9121), .ZN(n7317) );
  NAND2_X1 U8952 ( .A1(n7319), .A2(n7317), .ZN(n7321) );
  INV_X1 U8953 ( .A(n7915), .ZN(n7316) );
  AND2_X1 U8954 ( .A1(n7317), .A2(n7316), .ZN(n7318) );
  INV_X1 U8955 ( .A(n7381), .ZN(n7320) );
  AOI21_X1 U8956 ( .B1(n7915), .B2(n7321), .A(n7320), .ZN(n7405) );
  NOR2_X1 U8957 ( .A1(n7405), .A2(n9329), .ZN(n7322) );
  AOI211_X1 U8958 ( .C1(n7401), .C2(n7677), .A(n7323), .B(n7322), .ZN(n7324)
         );
  OAI21_X1 U8959 ( .B1(n9739), .B2(n7404), .A(n7324), .ZN(P1_U3281) );
  INV_X1 U8960 ( .A(n7438), .ZN(n7481) );
  AOI21_X1 U8961 ( .B1(n7326), .B2(n7325), .A(n9835), .ZN(n7327) );
  NAND2_X1 U8962 ( .A1(n7327), .A2(n9471), .ZN(n7332) );
  INV_X1 U8963 ( .A(n8454), .ZN(n8320) );
  OAI22_X1 U8964 ( .A1(n8320), .A2(n8219), .B1(n9831), .B2(n7328), .ZN(n7329)
         );
  AOI211_X1 U8965 ( .C1(n8211), .C2(n7375), .A(n7330), .B(n7329), .ZN(n7331)
         );
  OAI211_X1 U8966 ( .C1(n7481), .C2(n8214), .A(n7332), .B(n7331), .ZN(P2_U3236) );
  INV_X1 U8967 ( .A(n7333), .ZN(n7359) );
  OAI222_X1 U8968 ( .A1(n8975), .A2(n7359), .B1(n7335), .B2(P2_U3152), .C1(
        n7334), .C2(n8971), .ZN(P2_U3334) );
  INV_X1 U8969 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7341) );
  AOI211_X1 U8970 ( .C1(n9475), .C2(n7361), .A(n7337), .B(n7336), .ZN(n7338)
         );
  OAI21_X1 U8971 ( .B1(n7339), .B2(n8785), .A(n7338), .ZN(n7342) );
  NAND2_X1 U8972 ( .A1(n7342), .A2(n9944), .ZN(n7340) );
  OAI21_X1 U8973 ( .B1(n9944), .B2(n7341), .A(n7340), .ZN(P2_U3487) );
  NAND2_X1 U8974 ( .A1(n7342), .A2(n9954), .ZN(n7343) );
  OAI21_X1 U8975 ( .B1(n9954), .B2(n6973), .A(n7343), .ZN(P2_U3532) );
  INV_X1 U8976 ( .A(n7344), .ZN(n7348) );
  NOR3_X1 U8977 ( .A1(n7346), .A2(n7345), .A3(n8202), .ZN(n7347) );
  AOI21_X1 U8978 ( .B1(n7348), .B2(n9845), .A(n7347), .ZN(n7356) );
  NAND2_X1 U8979 ( .A1(n8211), .A2(n4841), .ZN(n7350) );
  OAI211_X1 U8980 ( .C1(n7351), .C2(n8209), .A(n7350), .B(n7349), .ZN(n7354)
         );
  NOR2_X1 U8981 ( .A1(n7352), .A2(n9835), .ZN(n7353) );
  AOI211_X1 U8982 ( .C1(n9854), .C2(n7361), .A(n7354), .B(n7353), .ZN(n7355)
         );
  OAI21_X1 U8983 ( .B1(n7357), .B2(n7356), .A(n7355), .ZN(P2_U3226) );
  OAI222_X1 U8984 ( .A1(n8045), .A2(n7360), .B1(n8048), .B2(n7359), .C1(n7358), 
        .C2(P1_U3084), .ZN(P1_U3329) );
  OR2_X1 U8985 ( .A1(n7438), .A2(n7434), .ZN(n8316) );
  NAND2_X1 U8986 ( .A1(n7438), .A2(n7434), .ZN(n8315) );
  NAND2_X1 U8987 ( .A1(n7363), .A2(n8419), .ZN(n7364) );
  AND2_X1 U8988 ( .A1(n7440), .A2(n7364), .ZN(n7484) );
  NAND2_X1 U8989 ( .A1(n7366), .A2(n7365), .ZN(n7367) );
  NAND2_X1 U8990 ( .A1(n7367), .A2(n8417), .ZN(n7432) );
  XNOR2_X1 U8991 ( .A(n7432), .B(n4755), .ZN(n7369) );
  AOI22_X1 U8992 ( .A1(n8456), .A2(n8656), .B1(n8654), .B2(n8454), .ZN(n7368)
         );
  OAI21_X1 U8993 ( .B1(n7369), .B2(n8707), .A(n7368), .ZN(n7370) );
  AOI21_X1 U8994 ( .B1(n7484), .B2(n7371), .A(n7370), .ZN(n7486) );
  INV_X1 U8995 ( .A(n7372), .ZN(n7613) );
  AND2_X1 U8996 ( .A1(n7373), .A2(n7438), .ZN(n7374) );
  OR2_X1 U8997 ( .A1(n7374), .A2(n7442), .ZN(n7482) );
  AOI22_X1 U8998 ( .A1(n7135), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7375), .B2(
        n8697), .ZN(n7377) );
  NAND2_X1 U8999 ( .A1(n7438), .A2(n8666), .ZN(n7376) );
  OAI211_X1 U9000 ( .C1(n7482), .C2(n8621), .A(n7377), .B(n7376), .ZN(n7378)
         );
  AOI21_X1 U9001 ( .B1(n7484), .B2(n7613), .A(n7378), .ZN(n7379) );
  OAI21_X1 U9002 ( .B1(n7486), .B2(n7135), .A(n7379), .ZN(P2_U3283) );
  OR2_X1 U9003 ( .A1(n7402), .A2(n9120), .ZN(n7380) );
  NAND2_X1 U9004 ( .A1(n7388), .A2(n9455), .ZN(n7383) );
  NOR2_X1 U9005 ( .A1(n7388), .A2(n9455), .ZN(n7382) );
  NAND2_X1 U9006 ( .A1(n7560), .A2(n9512), .ZN(n7826) );
  NAND2_X1 U9007 ( .A1(n7827), .A2(n7826), .ZN(n7917) );
  OR2_X1 U9008 ( .A1(n7384), .A2(n7917), .ZN(n7385) );
  NAND2_X1 U9009 ( .A1(n7562), .A2(n7385), .ZN(n9529) );
  AOI22_X1 U9010 ( .A1(n9726), .A2(n9118), .B1(n9455), .B2(n9729), .ZN(n7394)
         );
  AND2_X1 U9011 ( .A1(n7821), .A2(n7812), .ZN(n7757) );
  NAND2_X1 U9012 ( .A1(n7808), .A2(n7805), .ZN(n7815) );
  NAND2_X1 U9013 ( .A1(n7815), .A2(n7821), .ZN(n7746) );
  INV_X1 U9014 ( .A(n9455), .ZN(n7387) );
  OR2_X1 U9015 ( .A1(n7388), .A2(n7387), .ZN(n7563) );
  NAND2_X1 U9016 ( .A1(n7388), .A2(n7387), .ZN(n7825) );
  NAND2_X1 U9017 ( .A1(n9510), .A2(n9511), .ZN(n9509) );
  INV_X1 U9018 ( .A(n9509), .ZN(n7389) );
  INV_X1 U9019 ( .A(n7825), .ZN(n7390) );
  OAI21_X1 U9020 ( .B1(n7389), .B2(n7390), .A(n7917), .ZN(n7392) );
  NOR2_X1 U9021 ( .A1(n7917), .A2(n7390), .ZN(n7391) );
  NAND2_X1 U9022 ( .A1(n9509), .A2(n7391), .ZN(n7566) );
  NAND3_X1 U9023 ( .A1(n7392), .A2(n9704), .A3(n7566), .ZN(n7393) );
  OAI211_X1 U9024 ( .C1(n9529), .C2(n9707), .A(n7394), .B(n7393), .ZN(n9533)
         );
  NAND2_X1 U9025 ( .A1(n9533), .A2(n9737), .ZN(n7399) );
  NAND2_X1 U9026 ( .A1(n9507), .A2(n9535), .ZN(n9506) );
  OR2_X2 U9027 ( .A1(n9506), .A2(n7560), .ZN(n7569) );
  INV_X1 U9028 ( .A(n7569), .ZN(n9500) );
  AOI211_X1 U9029 ( .C1(n7560), .C2(n9506), .A(n9801), .B(n9500), .ZN(n9530)
         );
  INV_X1 U9030 ( .A(n7560), .ZN(n9457) );
  AOI22_X1 U9031 ( .A1(n9739), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7395), .B2(
        n9718), .ZN(n7396) );
  OAI21_X1 U9032 ( .B1(n9457), .B2(n9710), .A(n7396), .ZN(n7397) );
  AOI21_X1 U9033 ( .B1(n9530), .B2(n7677), .A(n7397), .ZN(n7398) );
  OAI211_X1 U9034 ( .C1(n9529), .C2(n7590), .A(n7399), .B(n7398), .ZN(P1_U3279) );
  INV_X1 U9035 ( .A(n7980), .ZN(n7400) );
  NAND2_X1 U9036 ( .A1(n8043), .A2(n7400), .ZN(n9748) );
  AOI21_X1 U9037 ( .B1(n9422), .B2(n7402), .A(n7401), .ZN(n7403) );
  OAI211_X1 U9038 ( .C1(n9425), .C2(n7405), .A(n7404), .B(n7403), .ZN(n7408)
         );
  NAND2_X1 U9039 ( .A1(n7408), .A2(n9826), .ZN(n7406) );
  OAI21_X1 U9040 ( .B1(n9826), .B2(n7407), .A(n7406), .ZN(P1_U3533) );
  INV_X1 U9041 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7410) );
  NAND2_X1 U9042 ( .A1(n7408), .A2(n9809), .ZN(n7409) );
  OAI21_X1 U9043 ( .B1(n9809), .B2(n7410), .A(n7409), .ZN(P1_U3484) );
  XOR2_X1 U9044 ( .A(n7417), .B(n7508), .Z(n7412) );
  NOR2_X1 U9045 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n7412), .ZN(n7510) );
  AOI21_X1 U9046 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n7412), .A(n7510), .ZN(
        n7421) );
  AND2_X1 U9047 ( .A1(n10007), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7414) );
  NOR2_X1 U9048 ( .A1(n9861), .A2(n7417), .ZN(n7413) );
  AOI211_X1 U9049 ( .C1(n9870), .C2(P2_ADDR_REG_15__SCAN_IN), .A(n7414), .B(
        n7413), .ZN(n7420) );
  AOI21_X1 U9050 ( .B1(n7218), .B2(n7416), .A(n7415), .ZN(n7500) );
  XNOR2_X1 U9051 ( .A(n7500), .B(n7417), .ZN(n7418) );
  NAND2_X1 U9052 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n7418), .ZN(n7501) );
  OAI211_X1 U9053 ( .C1(n7418), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9871), .B(
        n7501), .ZN(n7419) );
  OAI211_X1 U9054 ( .C1(n7421), .C2(n8490), .A(n7420), .B(n7419), .ZN(P2_U3260) );
  XNOR2_X1 U9055 ( .A(n7423), .B(n7422), .ZN(n7424) );
  XNOR2_X1 U9056 ( .A(n7425), .B(n7424), .ZN(n7431) );
  NAND2_X1 U9057 ( .A1(n9099), .A2(n9497), .ZN(n7428) );
  AOI21_X1 U9058 ( .B1(n9101), .B2(n9117), .A(n7426), .ZN(n7427) );
  OAI211_X1 U9059 ( .C1(n9512), .C2(n9104), .A(n7428), .B(n7427), .ZN(n7429)
         );
  AOI21_X1 U9060 ( .B1(n9499), .B2(n9107), .A(n7429), .ZN(n7430) );
  OAI21_X1 U9061 ( .B1(n7431), .B2(n9460), .A(n7430), .ZN(P1_U3232) );
  NAND2_X1 U9062 ( .A1(n7432), .A2(n8419), .ZN(n7433) );
  XNOR2_X1 U9063 ( .A(n9476), .B(n8454), .ZN(n7522) );
  XNOR2_X1 U9064 ( .A(n7524), .B(n7522), .ZN(n7437) );
  OR2_X1 U9065 ( .A1(n7434), .A2(n8562), .ZN(n7436) );
  OR2_X1 U9066 ( .A1(n7602), .A2(n8564), .ZN(n7435) );
  NAND2_X1 U9067 ( .A1(n7436), .A2(n7435), .ZN(n9469) );
  AOI21_X1 U9068 ( .B1(n7437), .B2(n8659), .A(n9469), .ZN(n9484) );
  NAND2_X1 U9069 ( .A1(n7438), .A2(n8455), .ZN(n7439) );
  XNOR2_X1 U9070 ( .A(n7520), .B(n7522), .ZN(n9487) );
  NAND2_X1 U9071 ( .A1(n9487), .A2(n8662), .ZN(n7446) );
  OAI22_X1 U9072 ( .A1(n8688), .A2(n7441), .B1(n9482), .B2(n8679), .ZN(n7444)
         );
  INV_X1 U9073 ( .A(n9476), .ZN(n8319) );
  OAI21_X1 U9074 ( .B1(n7442), .B2(n8319), .A(n7528), .ZN(n9485) );
  NOR2_X1 U9075 ( .A1(n9485), .A2(n8621), .ZN(n7443) );
  AOI211_X1 U9076 ( .C1(n8666), .C2(n9476), .A(n7444), .B(n7443), .ZN(n7445)
         );
  OAI211_X1 U9077 ( .C1(n7135), .C2(n9484), .A(n7446), .B(n7445), .ZN(P2_U3282) );
  AOI22_X1 U9078 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n9130), .B1(n7472), .B2(
        n9129), .ZN(n7456) );
  INV_X1 U9079 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n7454) );
  XNOR2_X1 U9080 ( .A(n9657), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9665) );
  INV_X1 U9081 ( .A(n7462), .ZN(n9645) );
  INV_X1 U9082 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7453) );
  XOR2_X1 U9083 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n7462), .Z(n9649) );
  INV_X1 U9084 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7449) );
  AOI22_X1 U9085 ( .A1(n9624), .A2(n7449), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n7450), .ZN(n9619) );
  NOR2_X1 U9086 ( .A1(n9620), .A2(n9619), .ZN(n9618) );
  NAND2_X1 U9087 ( .A1(n9635), .A2(n7451), .ZN(n7452) );
  XOR2_X1 U9088 ( .A(n9635), .B(n7451), .Z(n9638) );
  NAND2_X1 U9089 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9638), .ZN(n9637) );
  NAND2_X1 U9090 ( .A1(n7452), .A2(n9637), .ZN(n9650) );
  NAND2_X1 U9091 ( .A1(n9649), .A2(n9650), .ZN(n9648) );
  OAI21_X1 U9092 ( .B1(n9645), .B2(n7453), .A(n9648), .ZN(n9664) );
  NAND2_X1 U9093 ( .A1(n9665), .A2(n9664), .ZN(n9662) );
  OAI21_X1 U9094 ( .B1(n9657), .B2(n7454), .A(n9662), .ZN(n7455) );
  NOR2_X1 U9095 ( .A1(n7456), .A2(n7455), .ZN(n9128) );
  AOI21_X1 U9096 ( .B1(n7456), .B2(n7455), .A(n9128), .ZN(n7479) );
  INV_X1 U9097 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n7458) );
  NAND2_X1 U9098 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9089) );
  OR2_X1 U9099 ( .A1(n9658), .A2(n9130), .ZN(n7457) );
  OAI211_X1 U9100 ( .C1(n9632), .C2(n7458), .A(n9089), .B(n7457), .ZN(n7459)
         );
  INV_X1 U9101 ( .A(n7459), .ZN(n7478) );
  NAND2_X1 U9102 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n7460), .ZN(n7471) );
  INV_X1 U9103 ( .A(n7471), .ZN(n7461) );
  AOI21_X1 U9104 ( .B1(n5956), .B2(n9657), .A(n7461), .ZN(n9668) );
  NAND2_X1 U9105 ( .A1(n7462), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7470) );
  OR2_X1 U9106 ( .A1(n7462), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7463) );
  AND2_X1 U9107 ( .A1(n7463), .A2(n7470), .ZN(n9652) );
  NAND2_X1 U9108 ( .A1(n7465), .A2(n7464), .ZN(n7466) );
  NOR2_X1 U9109 ( .A1(n9624), .A2(n7466), .ZN(n7467) );
  XNOR2_X1 U9110 ( .A(n7466), .B(n9624), .ZN(n9617) );
  NOR2_X1 U9111 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(n9617), .ZN(n9616) );
  NOR2_X1 U9112 ( .A1(n7467), .A2(n9616), .ZN(n7468) );
  NAND2_X1 U9113 ( .A1(n9635), .A2(n7468), .ZN(n7469) );
  XOR2_X1 U9114 ( .A(n9635), .B(n7468), .Z(n9640) );
  NAND2_X1 U9115 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n9640), .ZN(n9639) );
  NAND2_X1 U9116 ( .A1(n7469), .A2(n9639), .ZN(n9653) );
  NAND2_X1 U9117 ( .A1(n9652), .A2(n9653), .ZN(n9651) );
  NAND2_X1 U9118 ( .A1(n7470), .A2(n9651), .ZN(n9669) );
  NAND2_X1 U9119 ( .A1(n9668), .A2(n9669), .ZN(n9666) );
  NAND2_X1 U9120 ( .A1(n7471), .A2(n9666), .ZN(n7476) );
  OR2_X1 U9121 ( .A1(n7472), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7474) );
  NAND2_X1 U9122 ( .A1(n7472), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7473) );
  AND2_X1 U9123 ( .A1(n7474), .A2(n7473), .ZN(n7475) );
  NAND2_X1 U9124 ( .A1(n7475), .A2(n7476), .ZN(n9126) );
  OAI211_X1 U9125 ( .C1(n7476), .C2(n7475), .A(n9667), .B(n9126), .ZN(n7477)
         );
  OAI211_X1 U9126 ( .C1(n7479), .C2(n9621), .A(n7478), .B(n7477), .ZN(P1_U3259) );
  INV_X1 U9127 ( .A(n7480), .ZN(n9941) );
  OAI22_X1 U9128 ( .A1(n7482), .A2(n9936), .B1(n7481), .B2(n9934), .ZN(n7483)
         );
  AOI21_X1 U9129 ( .B1(n7484), .B2(n9941), .A(n7483), .ZN(n7485) );
  AND2_X1 U9130 ( .A1(n7486), .A2(n7485), .ZN(n7488) );
  MUX2_X1 U9131 ( .A(n6977), .B(n7488), .S(n9954), .Z(n7487) );
  INV_X1 U9132 ( .A(n7487), .ZN(P2_U3533) );
  INV_X1 U9133 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7489) );
  MUX2_X1 U9134 ( .A(n7489), .B(n7488), .S(n9944), .Z(n7490) );
  INV_X1 U9135 ( .A(n7490), .ZN(P2_U3490) );
  NOR2_X1 U9136 ( .A1(n7543), .A2(n9835), .ZN(n7493) );
  NOR2_X1 U9137 ( .A1(n8202), .A2(n7602), .ZN(n7545) );
  OAI211_X1 U9138 ( .C1(n7493), .C2(n7545), .A(n7544), .B(n4512), .ZN(n7498)
         );
  INV_X1 U9139 ( .A(n7609), .ZN(n7494) );
  OAI22_X1 U9140 ( .A1(n9860), .A2(n7494), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8840), .ZN(n7496) );
  OAI22_X1 U9141 ( .A1(n7602), .A2(n9831), .B1(n8219), .B2(n8203), .ZN(n7495)
         );
  AOI211_X1 U9142 ( .C1(n8795), .C2(n9854), .A(n7496), .B(n7495), .ZN(n7497)
         );
  OAI211_X1 U9143 ( .C1(n7491), .C2(n9835), .A(n7498), .B(n7497), .ZN(P2_U3228) );
  INV_X1 U9144 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n7499) );
  AOI22_X1 U9145 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n7505), .B1(n8477), .B2(
        n7499), .ZN(n7504) );
  NAND2_X1 U9146 ( .A1(n7509), .A2(n7500), .ZN(n7502) );
  NAND2_X1 U9147 ( .A1(n7502), .A2(n7501), .ZN(n7503) );
  NOR2_X1 U9148 ( .A1(n7504), .A2(n7503), .ZN(n8479) );
  AOI21_X1 U9149 ( .B1(n7504), .B2(n7503), .A(n8479), .ZN(n7518) );
  NOR2_X1 U9150 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8840), .ZN(n7507) );
  NOR2_X1 U9151 ( .A1(n9861), .A2(n7505), .ZN(n7506) );
  AOI211_X1 U9152 ( .C1(n9870), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n7507), .B(
        n7506), .ZN(n7517) );
  NOR2_X1 U9153 ( .A1(n7509), .A2(n7508), .ZN(n7511) );
  NOR2_X1 U9154 ( .A1(n7511), .A2(n7510), .ZN(n7515) );
  INV_X1 U9155 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7512) );
  MUX2_X1 U9156 ( .A(n7512), .B(P2_REG2_REG_16__SCAN_IN), .S(n8477), .Z(n7513)
         );
  INV_X1 U9157 ( .A(n7513), .ZN(n7514) );
  NAND2_X1 U9158 ( .A1(n7514), .A2(n7515), .ZN(n8468) );
  OAI211_X1 U9159 ( .C1(n7515), .C2(n7514), .A(n9879), .B(n8468), .ZN(n7516)
         );
  OAI211_X1 U9160 ( .C1(n7518), .C2(n9862), .A(n7517), .B(n7516), .ZN(P2_U3261) );
  OR2_X1 U9161 ( .A1(n9476), .A2(n8454), .ZN(n7519) );
  OR2_X1 U9162 ( .A1(n7552), .A2(n7602), .ZN(n8333) );
  NAND2_X1 U9163 ( .A1(n7552), .A2(n7602), .ZN(n8330) );
  NAND2_X1 U9164 ( .A1(n8333), .A2(n8330), .ZN(n8422) );
  OAI21_X1 U9165 ( .B1(n7521), .B2(n8422), .A(n7599), .ZN(n7654) );
  INV_X1 U9166 ( .A(n7654), .ZN(n7534) );
  INV_X1 U9167 ( .A(n7522), .ZN(n8421) );
  OR2_X1 U9168 ( .A1(n9476), .A2(n8320), .ZN(n7523) );
  INV_X1 U9169 ( .A(n7601), .ZN(n7525) );
  AOI21_X1 U9170 ( .B1(n7526), .B2(n8422), .A(n7525), .ZN(n7527) );
  OAI222_X1 U9171 ( .A1(n8564), .A2(n8154), .B1(n8562), .B2(n8320), .C1(n8707), 
        .C2(n7527), .ZN(n7652) );
  INV_X1 U9172 ( .A(n7528), .ZN(n7529) );
  INV_X1 U9173 ( .A(n7552), .ZN(n7650) );
  OAI21_X1 U9174 ( .B1(n7529), .B2(n7650), .A(n4338), .ZN(n7651) );
  AOI22_X1 U9175 ( .A1(n7135), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n7547), .B2(
        n8697), .ZN(n7531) );
  NAND2_X1 U9176 ( .A1(n7552), .A2(n8666), .ZN(n7530) );
  OAI211_X1 U9177 ( .C1(n7651), .C2(n8621), .A(n7531), .B(n7530), .ZN(n7532)
         );
  AOI21_X1 U9178 ( .B1(n7652), .B2(n8688), .A(n7532), .ZN(n7533) );
  OAI21_X1 U9179 ( .B1(n7534), .B2(n8711), .A(n7533), .ZN(P2_U3281) );
  INV_X1 U9180 ( .A(n7535), .ZN(n7538) );
  OAI222_X1 U9181 ( .A1(n8971), .A2(n8907), .B1(n8969), .B2(n7538), .C1(n10007), .C2(n7536), .ZN(P2_U3333) );
  OAI222_X1 U9182 ( .A1(n8045), .A2(n7539), .B1(n8048), .B2(n7538), .C1(
        P1_U3084), .C2(n7537), .ZN(P1_U3328) );
  INV_X1 U9183 ( .A(n7540), .ZN(n7558) );
  OAI222_X1 U9184 ( .A1(n8975), .A2(n7558), .B1(n7542), .B2(n10007), .C1(n7541), .C2(n8971), .ZN(P2_U3332) );
  AND2_X1 U9185 ( .A1(n7544), .A2(n7543), .ZN(n7556) );
  INV_X1 U9186 ( .A(n7545), .ZN(n7555) );
  NAND3_X1 U9187 ( .A1(n7556), .A2(n9845), .A3(n7546), .ZN(n7554) );
  INV_X1 U9188 ( .A(n7547), .ZN(n7549) );
  OAI22_X1 U9189 ( .A1(n9860), .A2(n7549), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7548), .ZN(n7551) );
  OAI22_X1 U9190 ( .A1(n8320), .A2(n9831), .B1(n8219), .B2(n8154), .ZN(n7550)
         );
  AOI211_X1 U9191 ( .C1(n7552), .C2(n9854), .A(n7551), .B(n7550), .ZN(n7553)
         );
  OAI211_X1 U9192 ( .C1(n7556), .C2(n7555), .A(n7554), .B(n7553), .ZN(P2_U3243) );
  OAI222_X1 U9193 ( .A1(P1_U3084), .A2(n7559), .B1(n8048), .B2(n7558), .C1(
        n7557), .C2(n9444), .ZN(P1_U3327) );
  XNOR2_X1 U9194 ( .A(n9421), .B(n9117), .ZN(n7920) );
  NAND2_X1 U9195 ( .A1(n7560), .A2(n9119), .ZN(n7561) );
  XOR2_X1 U9196 ( .A(n7920), .B(n7575), .Z(n9424) );
  INV_X1 U9197 ( .A(n9118), .ZN(n9452) );
  INV_X1 U9198 ( .A(n7563), .ZN(n7564) );
  NAND2_X1 U9199 ( .A1(n7826), .A2(n7564), .ZN(n7565) );
  AND2_X1 U9200 ( .A1(n7565), .A2(n7827), .ZN(n7841) );
  NAND2_X1 U9201 ( .A1(n7566), .A2(n7841), .ZN(n9493) );
  OR2_X1 U9202 ( .A1(n9499), .A2(n9452), .ZN(n7840) );
  NAND2_X1 U9203 ( .A1(n9499), .A2(n9452), .ZN(n7745) );
  NAND2_X1 U9204 ( .A1(n7840), .A2(n7745), .ZN(n9494) );
  XNOR2_X1 U9205 ( .A(n7576), .B(n7920), .ZN(n7568) );
  OAI222_X1 U9206 ( .A1(n9699), .A2(n9452), .B1(n9701), .B2(n7690), .C1(n9733), 
        .C2(n7568), .ZN(n9419) );
  AOI211_X1 U9207 ( .C1(n9421), .C2(n4329), .A(n9801), .B(n7584), .ZN(n9420)
         );
  NAND2_X1 U9208 ( .A1(n9420), .A2(n7677), .ZN(n7571) );
  AOI22_X1 U9209 ( .A1(n9739), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7628), .B2(
        n9718), .ZN(n7570) );
  OAI211_X1 U9210 ( .C1(n4677), .C2(n9710), .A(n7571), .B(n7570), .ZN(n7572)
         );
  AOI21_X1 U9211 ( .B1(n9419), .B2(n9737), .A(n7572), .ZN(n7573) );
  OAI21_X1 U9212 ( .B1(n9424), .B2(n9329), .A(n7573), .ZN(P1_U3277) );
  AND2_X1 U9213 ( .A1(n9421), .A2(n9117), .ZN(n7574) );
  NAND2_X1 U9214 ( .A1(n7669), .A2(n7690), .ZN(n7834) );
  NAND2_X1 U9215 ( .A1(n7761), .A2(n7834), .ZN(n7919) );
  XNOR2_X1 U9216 ( .A(n7671), .B(n7919), .ZN(n9413) );
  INV_X1 U9217 ( .A(n9413), .ZN(n7591) );
  NAND2_X1 U9218 ( .A1(n9413), .A2(n9730), .ZN(n7582) );
  INV_X1 U9219 ( .A(n9117), .ZN(n9496) );
  NOR2_X1 U9220 ( .A1(n9421), .A2(n9496), .ZN(n7843) );
  INV_X1 U9221 ( .A(n7919), .ZN(n7832) );
  XNOR2_X1 U9222 ( .A(n7672), .B(n7832), .ZN(n7580) );
  NAND2_X1 U9223 ( .A1(n9117), .A2(n9729), .ZN(n7578) );
  NAND2_X1 U9224 ( .A1(n9115), .A2(n9726), .ZN(n7577) );
  NAND2_X1 U9225 ( .A1(n7578), .A2(n7577), .ZN(n7579) );
  AOI21_X1 U9226 ( .B1(n7580), .B2(n9704), .A(n7579), .ZN(n7581) );
  NAND2_X1 U9227 ( .A1(n7582), .A2(n7581), .ZN(n9418) );
  NAND2_X1 U9228 ( .A1(n9418), .A2(n9737), .ZN(n7589) );
  OAI22_X1 U9229 ( .A1(n9737), .A2(n7583), .B1(n7664), .B2(n9709), .ZN(n7587)
         );
  OR2_X1 U9230 ( .A1(n7584), .A2(n9414), .ZN(n7585) );
  NAND2_X1 U9231 ( .A1(n4281), .A2(n7585), .ZN(n9415) );
  NOR2_X1 U9232 ( .A1(n9415), .A2(n9153), .ZN(n7586) );
  AOI211_X1 U9233 ( .C1(n9498), .C2(n7669), .A(n7587), .B(n7586), .ZN(n7588)
         );
  OAI211_X1 U9234 ( .C1(n7591), .C2(n7590), .A(n7589), .B(n7588), .ZN(P1_U3276) );
  INV_X1 U9235 ( .A(n7592), .ZN(n7597) );
  AOI21_X1 U9236 ( .B1(n7594), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n7593), .ZN(
        n7595) );
  OAI21_X1 U9237 ( .B1(n7597), .B2(n8048), .A(n7595), .ZN(P1_U3326) );
  OAI222_X1 U9238 ( .A1(n8969), .A2(n7597), .B1(n8441), .B2(P2_U3152), .C1(
        n7596), .C2(n8971), .ZN(P2_U3331) );
  NAND2_X1 U9239 ( .A1(n7650), .A2(n7602), .ZN(n7598) );
  OR2_X1 U9240 ( .A1(n8795), .A2(n8154), .ZN(n8326) );
  NAND2_X1 U9241 ( .A1(n8795), .A2(n8154), .ZN(n8327) );
  NAND2_X1 U9242 ( .A1(n8326), .A2(n8327), .ZN(n8423) );
  OAI21_X1 U9243 ( .B1(n4340), .B2(n8423), .A(n7638), .ZN(n7607) );
  OR2_X1 U9244 ( .A1(n7607), .A2(n7600), .ZN(n7606) );
  XNOR2_X1 U9245 ( .A(n7632), .B(n4443), .ZN(n7604) );
  OAI22_X1 U9246 ( .A1(n7602), .A2(n8562), .B1(n8203), .B2(n8564), .ZN(n7603)
         );
  AOI21_X1 U9247 ( .B1(n7604), .B2(n8659), .A(n7603), .ZN(n7605) );
  INV_X1 U9248 ( .A(n7607), .ZN(n8799) );
  AND2_X1 U9249 ( .A1(n4338), .A2(n8795), .ZN(n7608) );
  OR2_X1 U9250 ( .A1(n7608), .A2(n7643), .ZN(n8797) );
  AOI22_X1 U9251 ( .A1(n7135), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n7609), .B2(
        n8697), .ZN(n7611) );
  NAND2_X1 U9252 ( .A1(n8795), .A2(n8666), .ZN(n7610) );
  OAI211_X1 U9253 ( .C1(n8797), .C2(n8621), .A(n7611), .B(n7610), .ZN(n7612)
         );
  AOI21_X1 U9254 ( .B1(n8799), .B2(n7613), .A(n7612), .ZN(n7614) );
  OAI21_X1 U9255 ( .B1(n8800), .B2(n7135), .A(n7614), .ZN(P2_U3280) );
  INV_X1 U9256 ( .A(n7772), .ZN(n7617) );
  NAND2_X1 U9257 ( .A1(n8967), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7615) );
  OAI211_X1 U9258 ( .C1(n7617), .C2(n8969), .A(n7616), .B(n7615), .ZN(P2_U3330) );
  INV_X1 U9259 ( .A(n7619), .ZN(n7624) );
  AOI21_X1 U9260 ( .B1(n7620), .B2(n7619), .A(n7618), .ZN(n7621) );
  NOR2_X1 U9261 ( .A1(n7621), .A2(n9460), .ZN(n7622) );
  OAI21_X1 U9262 ( .B1(n7624), .B2(n7623), .A(n7622), .ZN(n7630) );
  NOR2_X1 U9263 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7625), .ZN(n9623) );
  AOI21_X1 U9264 ( .B1(n9101), .B2(n9116), .A(n9623), .ZN(n7626) );
  OAI21_X1 U9265 ( .B1(n9452), .B2(n9104), .A(n7626), .ZN(n7627) );
  AOI21_X1 U9266 ( .B1(n7628), .B2(n9099), .A(n7627), .ZN(n7629) );
  OAI211_X1 U9267 ( .C1(n4677), .C2(n9095), .A(n7630), .B(n7629), .ZN(P1_U3213) );
  NAND2_X1 U9268 ( .A1(n7772), .A2(n9447), .ZN(n7631) );
  OAI211_X1 U9269 ( .C1(n9444), .C2(n7773), .A(n7631), .B(n9549), .ZN(P1_U3325) );
  NAND2_X1 U9270 ( .A1(n7632), .A2(n4443), .ZN(n7633) );
  NAND2_X1 U9271 ( .A1(n7633), .A2(n8327), .ZN(n7634) );
  NAND2_X1 U9272 ( .A1(n8787), .A2(n8203), .ZN(n8329) );
  AOI21_X1 U9273 ( .B1(n7634), .B2(n4582), .A(n8707), .ZN(n7637) );
  OAI22_X1 U9274 ( .A1(n8155), .A2(n8564), .B1(n8154), .B2(n8562), .ZN(n7636)
         );
  AOI21_X1 U9275 ( .B1(n7637), .B2(n8071), .A(n7636), .ZN(n8790) );
  INV_X1 U9276 ( .A(n8154), .ZN(n8453) );
  INV_X1 U9277 ( .A(n7641), .ZN(n7639) );
  NAND2_X1 U9278 ( .A1(n7639), .A2(n4582), .ZN(n8050) );
  NAND2_X1 U9279 ( .A1(n7641), .A2(n7640), .ZN(n7642) );
  NAND2_X1 U9280 ( .A1(n8050), .A2(n7642), .ZN(n8792) );
  NAND2_X1 U9281 ( .A1(n8792), .A2(n8662), .ZN(n7649) );
  INV_X1 U9282 ( .A(n8787), .ZN(n8160) );
  OAI21_X1 U9283 ( .B1(n7643), .B2(n8160), .A(n9912), .ZN(n7644) );
  OR2_X1 U9284 ( .A1(n7644), .A2(n8694), .ZN(n8789) );
  INV_X1 U9285 ( .A(n8789), .ZN(n7647) );
  AOI22_X1 U9286 ( .A1(n7135), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8157), .B2(
        n8697), .ZN(n7645) );
  OAI21_X1 U9287 ( .B1(n8160), .B2(n8700), .A(n7645), .ZN(n7646) );
  AOI21_X1 U9288 ( .B1(n7647), .B2(n8703), .A(n7646), .ZN(n7648) );
  OAI211_X1 U9289 ( .C1(n7135), .C2(n8790), .A(n7649), .B(n7648), .ZN(P2_U3279) );
  INV_X1 U9290 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7655) );
  OAI22_X1 U9291 ( .A1(n7651), .A2(n9936), .B1(n7650), .B2(n9934), .ZN(n7653)
         );
  AOI211_X1 U9292 ( .C1(n9931), .C2(n7654), .A(n7653), .B(n7652), .ZN(n8962)
         );
  MUX2_X1 U9293 ( .A(n7655), .B(n8962), .S(n9954), .Z(n7656) );
  INV_X1 U9294 ( .A(n7656), .ZN(P2_U3535) );
  INV_X1 U9295 ( .A(n7661), .ZN(n7658) );
  OAI21_X1 U9296 ( .B1(n7658), .B2(n7657), .A(n9086), .ZN(n7668) );
  AOI21_X1 U9297 ( .B1(n7661), .B2(n7660), .A(n7659), .ZN(n7667) );
  NAND2_X1 U9298 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9633) );
  OAI21_X1 U9299 ( .B1(n9453), .B2(n9319), .A(n9633), .ZN(n7662) );
  AOI21_X1 U9300 ( .B1(n9456), .B2(n9117), .A(n7662), .ZN(n7663) );
  OAI21_X1 U9301 ( .B1(n7664), .B2(n9468), .A(n7663), .ZN(n7665) );
  AOI21_X1 U9302 ( .B1(n7669), .B2(n9107), .A(n7665), .ZN(n7666) );
  OAI21_X1 U9303 ( .B1(n7668), .B2(n7667), .A(n7666), .ZN(P1_U3239) );
  NOR2_X1 U9304 ( .A1(n7669), .A2(n9116), .ZN(n7670) );
  OR2_X1 U9305 ( .A1(n9410), .A2(n9319), .ZN(n7836) );
  NAND2_X1 U9306 ( .A1(n9410), .A2(n9319), .ZN(n7763) );
  NAND2_X1 U9307 ( .A1(n7836), .A2(n7763), .ZN(n7998) );
  XNOR2_X1 U9308 ( .A(n7999), .B(n7998), .ZN(n9412) );
  INV_X1 U9309 ( .A(n9301), .ZN(n8000) );
  NOR2_X1 U9310 ( .A1(n7672), .A2(n7919), .ZN(n7674) );
  INV_X1 U9311 ( .A(n7761), .ZN(n7673) );
  OR2_X1 U9312 ( .A1(n7674), .A2(n7673), .ZN(n7675) );
  OR2_X1 U9313 ( .A1(n7998), .A2(n7673), .ZN(n7848) );
  NOR2_X1 U9314 ( .A1(n7674), .A2(n7848), .ZN(n8011) );
  AOI21_X1 U9315 ( .B1(n7998), .B2(n7675), .A(n8011), .ZN(n7676) );
  OAI222_X1 U9316 ( .A1(n9701), .A2(n8000), .B1(n9699), .B2(n7690), .C1(n9733), 
        .C2(n7676), .ZN(n9408) );
  INV_X1 U9317 ( .A(n9410), .ZN(n7680) );
  AOI211_X1 U9318 ( .C1(n9410), .C2(n4281), .A(n9801), .B(n4564), .ZN(n9409)
         );
  NAND2_X1 U9319 ( .A1(n9409), .A2(n7677), .ZN(n7679) );
  AOI22_X1 U9320 ( .A1(n9739), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n7687), .B2(
        n9718), .ZN(n7678) );
  OAI211_X1 U9321 ( .C1(n7680), .C2(n9710), .A(n7679), .B(n7678), .ZN(n7681)
         );
  AOI21_X1 U9322 ( .B1(n9408), .B2(n9737), .A(n7681), .ZN(n7682) );
  OAI21_X1 U9323 ( .B1(n9329), .B2(n9412), .A(n7682), .ZN(P1_U3275) );
  XOR2_X1 U9324 ( .A(n7684), .B(n7683), .Z(n7685) );
  XNOR2_X1 U9325 ( .A(n4355), .B(n7685), .ZN(n7693) );
  NAND2_X1 U9326 ( .A1(n9099), .A2(n7687), .ZN(n7689) );
  AND2_X1 U9327 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9647) );
  AOI21_X1 U9328 ( .B1(n9101), .B2(n9301), .A(n9647), .ZN(n7688) );
  OAI211_X1 U9329 ( .C1(n7690), .C2(n9104), .A(n7689), .B(n7688), .ZN(n7691)
         );
  AOI21_X1 U9330 ( .B1(n9410), .B2(n9107), .A(n7691), .ZN(n7692) );
  OAI21_X1 U9331 ( .B1(n7693), .B2(n9460), .A(n7692), .ZN(P1_U3224) );
  INV_X1 U9332 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7778) );
  INV_X1 U9333 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8972) );
  MUX2_X1 U9334 ( .A(n7778), .B(n8972), .S(n7715), .Z(n7698) );
  INV_X1 U9335 ( .A(SI_29_), .ZN(n7697) );
  NAND2_X1 U9336 ( .A1(n7698), .A2(n7697), .ZN(n7706) );
  INV_X1 U9337 ( .A(n7698), .ZN(n7699) );
  NAND2_X1 U9338 ( .A1(n7699), .A2(SI_29_), .ZN(n7700) );
  INV_X1 U9339 ( .A(n8062), .ZN(n8974) );
  OAI222_X1 U9340 ( .A1(n8045), .A2(n7778), .B1(P1_U3084), .B2(n7701), .C1(
        n8048), .C2(n8974), .ZN(P1_U3324) );
  OAI222_X1 U9341 ( .A1(n8045), .A2(n7703), .B1(n8048), .B2(n7702), .C1(n7939), 
        .C2(P1_U3084), .ZN(P1_U3333) );
  NAND2_X1 U9342 ( .A1(n7705), .A2(n7704), .ZN(n7707) );
  NAND2_X1 U9343 ( .A1(n7707), .A2(n7706), .ZN(n7709) );
  INV_X1 U9344 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8046) );
  INV_X1 U9345 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8865) );
  MUX2_X1 U9346 ( .A(n8046), .B(n8865), .S(n7715), .Z(n7710) );
  INV_X1 U9347 ( .A(n7720), .ZN(n7708) );
  NAND2_X1 U9348 ( .A1(n7708), .A2(SI_30_), .ZN(n7714) );
  INV_X1 U9349 ( .A(n7709), .ZN(n7712) );
  INV_X1 U9350 ( .A(n7710), .ZN(n7711) );
  NAND2_X1 U9351 ( .A1(n7712), .A2(n7711), .ZN(n7713) );
  NAND2_X1 U9352 ( .A1(n7714), .A2(n7713), .ZN(n7718) );
  MUX2_X1 U9353 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7715), .Z(n7716) );
  XNOR2_X1 U9354 ( .A(n7716), .B(SI_31_), .ZN(n7717) );
  NOR2_X1 U9355 ( .A1(n5663), .A2(n6334), .ZN(n7719) );
  NAND2_X1 U9356 ( .A1(n8224), .A2(n7777), .ZN(n7722) );
  OR2_X1 U9357 ( .A1(n5663), .A2(n8046), .ZN(n7721) );
  NAND2_X1 U9358 ( .A1(n7722), .A2(n7721), .ZN(n9334) );
  NAND2_X1 U9359 ( .A1(n5675), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n7726) );
  NAND2_X1 U9360 ( .A1(n6153), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7725) );
  NAND2_X1 U9361 ( .A1(n7723), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7724) );
  AND3_X1 U9362 ( .A1(n7726), .A2(n7725), .A3(n7724), .ZN(n8033) );
  OR2_X1 U9363 ( .A1(n9334), .A2(n8033), .ZN(n7929) );
  OR2_X1 U9364 ( .A1(n9145), .A2(n7929), .ZN(n7727) );
  NAND2_X1 U9365 ( .A1(n9330), .A2(n9142), .ZN(n7930) );
  NAND2_X1 U9366 ( .A1(n9360), .A2(n9105), .ZN(n8023) );
  INV_X1 U9367 ( .A(n9206), .ZN(n9236) );
  NAND2_X1 U9368 ( .A1(n9366), .A2(n9236), .ZN(n9203) );
  OR2_X1 U9369 ( .A1(n9366), .A2(n9236), .ZN(n7943) );
  NAND2_X1 U9370 ( .A1(n9370), .A2(n9251), .ZN(n7958) );
  INV_X1 U9371 ( .A(n7958), .ZN(n7728) );
  NAND2_X1 U9372 ( .A1(n7943), .A2(n7728), .ZN(n7729) );
  NAND3_X1 U9373 ( .A1(n8023), .A2(n9203), .A3(n7729), .ZN(n7875) );
  INV_X1 U9374 ( .A(n7875), .ZN(n7771) );
  NAND2_X1 U9375 ( .A1(n9377), .A2(n9258), .ZN(n8021) );
  INV_X1 U9376 ( .A(n9276), .ZN(n9250) );
  INV_X1 U9377 ( .A(n9113), .ZN(n9286) );
  NAND2_X1 U9378 ( .A1(n9385), .A2(n9286), .ZN(n8016) );
  NAND2_X1 U9379 ( .A1(n7903), .A2(n4798), .ZN(n7730) );
  NAND2_X1 U9380 ( .A1(n9382), .A2(n9250), .ZN(n8018) );
  AND2_X1 U9381 ( .A1(n7730), .A2(n8018), .ZN(n7731) );
  AND2_X1 U9382 ( .A1(n8021), .A2(n7731), .ZN(n7868) );
  NOR2_X1 U9383 ( .A1(n9385), .A2(n9286), .ZN(n8017) );
  INV_X1 U9384 ( .A(n9300), .ZN(n9090) );
  OR2_X1 U9385 ( .A1(n9391), .A2(n9090), .ZN(n7904) );
  INV_X1 U9386 ( .A(n7904), .ZN(n7732) );
  OR2_X1 U9387 ( .A1(n8017), .A2(n7732), .ZN(n7859) );
  INV_X1 U9388 ( .A(n7859), .ZN(n7734) );
  INV_X1 U9389 ( .A(n9114), .ZN(n9320) );
  OR2_X1 U9390 ( .A1(n9397), .A2(n9320), .ZN(n7905) );
  OR2_X1 U9391 ( .A1(n9405), .A2(n8000), .ZN(n9296) );
  AND2_X1 U9392 ( .A1(n7905), .A2(n9296), .ZN(n8014) );
  NAND2_X1 U9393 ( .A1(n9391), .A2(n9090), .ZN(n8015) );
  NAND2_X1 U9394 ( .A1(n9397), .A2(n9320), .ZN(n8013) );
  NAND3_X1 U9395 ( .A1(n4808), .A2(n8015), .A3(n8013), .ZN(n7733) );
  NAND3_X1 U9396 ( .A1(n7734), .A2(n7903), .A3(n7733), .ZN(n7735) );
  OR2_X1 U9397 ( .A1(n9377), .A2(n9258), .ZN(n7902) );
  INV_X1 U9398 ( .A(n7902), .ZN(n7867) );
  OR2_X1 U9399 ( .A1(n9370), .A2(n9251), .ZN(n7872) );
  INV_X1 U9400 ( .A(n7872), .ZN(n8022) );
  AOI211_X1 U9401 ( .C1(n7868), .C2(n7735), .A(n7867), .B(n8022), .ZN(n7957)
         );
  INV_X1 U9402 ( .A(n7736), .ZN(n7740) );
  INV_X1 U9403 ( .A(n7737), .ZN(n7739) );
  OAI211_X1 U9404 ( .C1(n7740), .C2(n7739), .A(n7743), .B(n7738), .ZN(n7742)
         );
  NAND3_X1 U9405 ( .A1(n7742), .A2(n7795), .A3(n7741), .ZN(n7752) );
  NAND3_X1 U9406 ( .A1(n7744), .A2(n7796), .A3(n7743), .ZN(n7952) );
  NAND2_X1 U9407 ( .A1(n9405), .A2(n8000), .ZN(n8012) );
  AND2_X1 U9408 ( .A1(n8013), .A2(n8012), .ZN(n7854) );
  INV_X1 U9409 ( .A(n7854), .ZN(n7766) );
  INV_X1 U9410 ( .A(n7763), .ZN(n8010) );
  NAND2_X1 U9411 ( .A1(n9421), .A2(n9496), .ZN(n7754) );
  AND2_X1 U9412 ( .A1(n7754), .A2(n7745), .ZN(n7829) );
  AND2_X1 U9413 ( .A1(n7746), .A2(n7825), .ZN(n7747) );
  NAND2_X1 U9414 ( .A1(n7826), .A2(n7747), .ZN(n7756) );
  NAND2_X1 U9415 ( .A1(n7804), .A2(n7799), .ZN(n7748) );
  NOR2_X1 U9416 ( .A1(n7756), .A2(n7748), .ZN(n7749) );
  NAND3_X1 U9417 ( .A1(n7834), .A2(n7829), .A3(n7749), .ZN(n7750) );
  OR3_X1 U9418 ( .A1(n7766), .A2(n8010), .A3(n7750), .ZN(n7947) );
  AOI211_X1 U9419 ( .C1(n7796), .C2(n7752), .A(n7751), .B(n7947), .ZN(n7767)
         );
  INV_X1 U9420 ( .A(n7840), .ZN(n7753) );
  OR2_X1 U9421 ( .A1(n7843), .A2(n7753), .ZN(n7755) );
  NAND2_X1 U9422 ( .A1(n7755), .A2(n7754), .ZN(n7831) );
  OAI21_X1 U9423 ( .B1(n7757), .B2(n7756), .A(n7841), .ZN(n7758) );
  NAND2_X1 U9424 ( .A1(n7829), .A2(n7758), .ZN(n7759) );
  NAND2_X1 U9425 ( .A1(n7831), .A2(n7759), .ZN(n7760) );
  NAND2_X1 U9426 ( .A1(n7760), .A2(n7834), .ZN(n7762) );
  NAND3_X1 U9427 ( .A1(n7836), .A2(n7762), .A3(n7761), .ZN(n7764) );
  NAND2_X1 U9428 ( .A1(n7764), .A2(n7763), .ZN(n7765) );
  OAI22_X1 U9429 ( .A1(n7947), .A2(n7797), .B1(n7766), .B2(n7765), .ZN(n7944)
         );
  AND2_X1 U9430 ( .A1(n7868), .A2(n8015), .ZN(n7953) );
  OAI21_X1 U9431 ( .B1(n7767), .B2(n7944), .A(n7953), .ZN(n7768) );
  NAND3_X1 U9432 ( .A1(n7957), .A2(n7768), .A3(n7943), .ZN(n7770) );
  INV_X1 U9433 ( .A(n8024), .ZN(n7769) );
  NOR2_X1 U9434 ( .A1(n9355), .A2(n9178), .ZN(n8027) );
  AOI211_X1 U9435 ( .C1(n7771), .C2(n7770), .A(n7769), .B(n8027), .ZN(n7776)
         );
  NAND2_X1 U9436 ( .A1(n7772), .A2(n7777), .ZN(n7775) );
  OR2_X1 U9437 ( .A1(n5663), .A2(n7773), .ZN(n7774) );
  NAND2_X1 U9438 ( .A1(n9345), .A2(n9179), .ZN(n8029) );
  NAND2_X1 U9439 ( .A1(n9351), .A2(n9009), .ZN(n7901) );
  NAND2_X1 U9440 ( .A1(n8029), .A2(n7901), .ZN(n7966) );
  INV_X1 U9441 ( .A(n8028), .ZN(n9160) );
  NAND2_X1 U9442 ( .A1(n9355), .A2(n9178), .ZN(n8026) );
  NOR2_X1 U9443 ( .A1(n9160), .A2(n8026), .ZN(n7965) );
  AOI211_X1 U9444 ( .C1(n7776), .C2(n8028), .A(n7966), .B(n7965), .ZN(n7790)
         );
  NAND2_X1 U9445 ( .A1(n8062), .A2(n7777), .ZN(n7781) );
  OR2_X1 U9446 ( .A1(n5663), .A2(n7778), .ZN(n7780) );
  NAND2_X1 U9447 ( .A1(n5675), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n7787) );
  INV_X1 U9448 ( .A(n7782), .ZN(n8035) );
  NAND2_X1 U9449 ( .A1(n7783), .A2(n8035), .ZN(n7786) );
  NAND2_X1 U9450 ( .A1(n7723), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7785) );
  NAND2_X1 U9451 ( .A1(n6153), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n7784) );
  NAND4_X1 U9452 ( .A1(n7787), .A2(n7786), .A3(n7785), .A4(n7784), .ZN(n9164)
         );
  INV_X1 U9453 ( .A(n9164), .ZN(n7788) );
  NAND2_X1 U9454 ( .A1(n7890), .A2(n7900), .ZN(n7972) );
  NAND2_X1 U9455 ( .A1(n9337), .A2(n7788), .ZN(n7970) );
  INV_X1 U9456 ( .A(n8033), .ZN(n9110) );
  AOI21_X1 U9457 ( .B1(n9110), .B2(n7791), .A(n9149), .ZN(n7895) );
  INV_X1 U9458 ( .A(n7895), .ZN(n7789) );
  OAI211_X1 U9459 ( .C1(n7790), .C2(n7972), .A(n7970), .B(n7789), .ZN(n7793)
         );
  AND2_X1 U9460 ( .A1(n9145), .A2(n7791), .ZN(n7974) );
  INV_X1 U9461 ( .A(n7974), .ZN(n7792) );
  NAND2_X1 U9462 ( .A1(n7792), .A2(n7931), .ZN(n7936) );
  AOI21_X1 U9463 ( .B1(n7898), .B2(n7793), .A(n7936), .ZN(n7934) );
  AND2_X1 U9464 ( .A1(n8043), .A2(n9721), .ZN(n7881) );
  INV_X1 U9465 ( .A(n7881), .ZN(n7897) );
  OAI211_X1 U9466 ( .C1(n7798), .C2(n4834), .A(n7797), .B(n7796), .ZN(n7800)
         );
  NAND2_X1 U9467 ( .A1(n7800), .A2(n7799), .ZN(n7801) );
  INV_X1 U9468 ( .A(n7803), .ZN(n7806) );
  OAI211_X1 U9469 ( .C1(n7814), .C2(n7806), .A(n7805), .B(n7804), .ZN(n7811)
         );
  AND2_X1 U9470 ( .A1(n7821), .A2(n7807), .ZN(n7810) );
  NAND2_X1 U9471 ( .A1(n7826), .A2(n7808), .ZN(n7809) );
  AOI21_X1 U9472 ( .B1(n7811), .B2(n7810), .A(n7809), .ZN(n7820) );
  OAI21_X1 U9473 ( .B1(n7814), .B2(n7813), .A(n7812), .ZN(n7818) );
  INV_X1 U9474 ( .A(n7815), .ZN(n7817) );
  INV_X1 U9475 ( .A(n7827), .ZN(n7816) );
  AOI21_X1 U9476 ( .B1(n7818), .B2(n7817), .A(n7816), .ZN(n7819) );
  MUX2_X1 U9477 ( .A(n7820), .B(n7819), .S(n7881), .Z(n7824) );
  OR2_X1 U9478 ( .A1(n7821), .A2(n7897), .ZN(n7822) );
  AND2_X1 U9479 ( .A1(n9511), .A2(n7822), .ZN(n7823) );
  NAND2_X1 U9480 ( .A1(n7826), .A2(n7825), .ZN(n7828) );
  OR2_X1 U9481 ( .A1(n7829), .A2(n7843), .ZN(n7830) );
  MUX2_X1 U9482 ( .A(n7831), .B(n7830), .S(n7897), .Z(n7833) );
  AND2_X1 U9483 ( .A1(n7833), .A2(n7832), .ZN(n7846) );
  INV_X1 U9484 ( .A(n7834), .ZN(n7835) );
  NOR2_X1 U9485 ( .A1(n7998), .A2(n7835), .ZN(n7838) );
  INV_X1 U9486 ( .A(n7836), .ZN(n7837) );
  AOI21_X1 U9487 ( .B1(n7839), .B2(n7838), .A(n7837), .ZN(n7852) );
  NAND2_X1 U9488 ( .A1(n7841), .A2(n7840), .ZN(n7842) );
  NOR2_X1 U9489 ( .A1(n7843), .A2(n7842), .ZN(n7844) );
  NAND2_X1 U9490 ( .A1(n7845), .A2(n7844), .ZN(n7847) );
  NAND2_X1 U9491 ( .A1(n7847), .A2(n7846), .ZN(n7850) );
  INV_X1 U9492 ( .A(n7848), .ZN(n7849) );
  AOI21_X1 U9493 ( .B1(n7850), .B2(n7849), .A(n8010), .ZN(n7851) );
  NAND2_X1 U9494 ( .A1(n7853), .A2(n9316), .ZN(n7856) );
  MUX2_X1 U9495 ( .A(n7854), .B(n8014), .S(n7897), .Z(n7855) );
  AND2_X1 U9496 ( .A1(n7904), .A2(n7905), .ZN(n7858) );
  NAND2_X1 U9497 ( .A1(n8016), .A2(n8015), .ZN(n7857) );
  AOI21_X1 U9498 ( .B1(n7861), .B2(n7858), .A(n7857), .ZN(n7863) );
  AND2_X1 U9499 ( .A1(n8015), .A2(n8013), .ZN(n7860) );
  AOI21_X1 U9500 ( .B1(n7861), .B2(n7860), .A(n7859), .ZN(n7862) );
  NAND2_X1 U9501 ( .A1(n4810), .A2(n7903), .ZN(n7864) );
  OAI21_X1 U9502 ( .B1(n7866), .B2(n7864), .A(n8018), .ZN(n7865) );
  AOI21_X1 U9503 ( .B1(n7865), .B2(n7902), .A(n4794), .ZN(n7871) );
  NAND2_X1 U9504 ( .A1(n7866), .A2(n7903), .ZN(n7869) );
  AOI21_X1 U9505 ( .B1(n7869), .B2(n7868), .A(n7867), .ZN(n7870) );
  NAND2_X1 U9506 ( .A1(n7872), .A2(n7958), .ZN(n9235) );
  INV_X1 U9507 ( .A(n9235), .ZN(n9227) );
  NAND3_X1 U9508 ( .A1(n9227), .A2(n7943), .A3(n9203), .ZN(n7878) );
  NAND2_X1 U9509 ( .A1(n9203), .A2(n8022), .ZN(n7873) );
  NAND3_X1 U9510 ( .A1(n8024), .A2(n7943), .A3(n7873), .ZN(n7874) );
  MUX2_X1 U9511 ( .A(n7875), .B(n7874), .S(n7897), .Z(n7876) );
  INV_X1 U9512 ( .A(n7876), .ZN(n7877) );
  OAI21_X1 U9513 ( .B1(n7879), .B2(n7878), .A(n7877), .ZN(n7885) );
  MUX2_X1 U9514 ( .A(n8024), .B(n8023), .S(n7897), .Z(n7880) );
  XNOR2_X1 U9515 ( .A(n9355), .B(n9207), .ZN(n9190) );
  AND2_X1 U9516 ( .A1(n7880), .A2(n9190), .ZN(n7884) );
  NAND2_X1 U9517 ( .A1(n7901), .A2(n8026), .ZN(n7882) );
  MUX2_X1 U9518 ( .A(n8027), .B(n7882), .S(n7881), .Z(n7883) );
  AOI21_X1 U9519 ( .B1(n7885), .B2(n7884), .A(n7883), .ZN(n7889) );
  INV_X1 U9520 ( .A(n7900), .ZN(n7886) );
  NOR2_X1 U9521 ( .A1(n7887), .A2(n4826), .ZN(n7888) );
  INV_X1 U9522 ( .A(n7890), .ZN(n7891) );
  MUX2_X1 U9523 ( .A(n7970), .B(n7892), .S(n7897), .Z(n7893) );
  OAI211_X1 U9524 ( .C1(n7894), .C2(n8030), .A(n7898), .B(n7893), .ZN(n7896)
         );
  NOR2_X1 U9525 ( .A1(n9149), .A2(n9110), .ZN(n7969) );
  NAND2_X1 U9526 ( .A1(n7900), .A2(n8029), .ZN(n9155) );
  INV_X1 U9527 ( .A(n9155), .ZN(n9162) );
  INV_X1 U9528 ( .A(n9177), .ZN(n7968) );
  XNOR2_X1 U9529 ( .A(n9366), .B(n9206), .ZN(n9219) );
  NAND2_X1 U9530 ( .A1(n7903), .A2(n8018), .ZN(n9255) );
  INV_X1 U9531 ( .A(n9255), .ZN(n8020) );
  NOR2_X1 U9532 ( .A1(n8017), .A2(n4798), .ZN(n9275) );
  NAND2_X1 U9533 ( .A1(n7904), .A2(n8015), .ZN(n9283) );
  INV_X1 U9534 ( .A(n9310), .ZN(n9298) );
  INV_X1 U9535 ( .A(n9316), .ZN(n7924) );
  INV_X1 U9536 ( .A(n7998), .ZN(n7922) );
  NOR4_X1 U9537 ( .A1(n7907), .A2(n9724), .A3(n9698), .A4(n7906), .ZN(n7910)
         );
  NAND4_X1 U9538 ( .A1(n7910), .A2(n9680), .A3(n7909), .A4(n7908), .ZN(n7914)
         );
  NOR4_X1 U9539 ( .A1(n7914), .A2(n7913), .A3(n7096), .A4(n7912), .ZN(n7916)
         );
  NAND3_X1 U9540 ( .A1(n7916), .A2(n9511), .A3(n7915), .ZN(n7918) );
  NOR4_X1 U9541 ( .A1(n7919), .A2(n9494), .A3(n7918), .A4(n7917), .ZN(n7921)
         );
  NAND3_X1 U9542 ( .A1(n7922), .A2(n7921), .A3(n7920), .ZN(n7923) );
  NOR4_X1 U9543 ( .A1(n9283), .A2(n9298), .A3(n7924), .A4(n7923), .ZN(n7925)
         );
  NAND4_X1 U9544 ( .A1(n4278), .A2(n8020), .A3(n9275), .A4(n7925), .ZN(n7926)
         );
  NOR4_X1 U9545 ( .A1(n9205), .A2(n4788), .A3(n9235), .A4(n7926), .ZN(n7927)
         );
  NAND4_X1 U9546 ( .A1(n9162), .A2(n7968), .A3(n7927), .A4(n9190), .ZN(n7928)
         );
  NOR4_X1 U9547 ( .A1(n7974), .A2(n7969), .A3(n8030), .A4(n7928), .ZN(n7932)
         );
  AND2_X1 U9548 ( .A1(n7930), .A2(n7929), .ZN(n7976) );
  AOI21_X1 U9549 ( .B1(n7932), .B2(n7976), .A(n7931), .ZN(n7935) );
  NAND2_X1 U9550 ( .A1(n7935), .A2(n9137), .ZN(n7942) );
  NOR2_X1 U9551 ( .A1(n7936), .A2(n6134), .ZN(n7937) );
  NAND2_X1 U9552 ( .A1(n7938), .A2(n7937), .ZN(n7941) );
  INV_X1 U9553 ( .A(n7943), .ZN(n7964) );
  INV_X1 U9554 ( .A(n7944), .ZN(n7956) );
  AOI21_X1 U9555 ( .B1(n9727), .B2(n6718), .A(n8041), .ZN(n7946) );
  INV_X1 U9556 ( .A(n7947), .ZN(n7950) );
  INV_X1 U9557 ( .A(n7948), .ZN(n7949) );
  OAI211_X1 U9558 ( .C1(n7952), .C2(n7951), .A(n7950), .B(n7949), .ZN(n7955)
         );
  INV_X1 U9559 ( .A(n7953), .ZN(n7954) );
  AOI21_X1 U9560 ( .B1(n7956), .B2(n7955), .A(n7954), .ZN(n7960) );
  INV_X1 U9561 ( .A(n7957), .ZN(n7959) );
  OAI211_X1 U9562 ( .C1(n7960), .C2(n7959), .A(n7958), .B(n9203), .ZN(n7962)
         );
  INV_X1 U9563 ( .A(n8023), .ZN(n7961) );
  OAI21_X1 U9564 ( .B1(n7962), .B2(n7961), .A(n8024), .ZN(n7963) );
  AOI211_X1 U9565 ( .C1(n7964), .C2(n8023), .A(n7963), .B(n8027), .ZN(n7967)
         );
  AOI211_X1 U9566 ( .C1(n7968), .C2(n7967), .A(n7966), .B(n7965), .ZN(n7973)
         );
  INV_X1 U9567 ( .A(n7969), .ZN(n7971) );
  OAI211_X1 U9568 ( .C1(n7973), .C2(n7972), .A(n7971), .B(n7970), .ZN(n7975)
         );
  AOI21_X1 U9569 ( .B1(n7976), .B2(n7975), .A(n7974), .ZN(n7981) );
  NAND2_X1 U9570 ( .A1(n7981), .A2(n7977), .ZN(n7979) );
  OAI211_X1 U9571 ( .C1(n7981), .C2(n7980), .A(n7979), .B(n7978), .ZN(n7986)
         );
  NAND2_X1 U9572 ( .A1(n7982), .A2(n9577), .ZN(n7983) );
  OAI211_X1 U9573 ( .C1(n6134), .C2(n7984), .A(n7983), .B(P1_B_REG_SCAN_IN), 
        .ZN(n7985) );
  AOI22_X1 U9574 ( .A1(n9844), .A2(n7987), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n7988) );
  OAI21_X1 U9575 ( .B1(n7989), .B2(n9860), .A(n7988), .ZN(n7994) );
  INV_X1 U9576 ( .A(n8202), .ZN(n9850) );
  AOI22_X1 U9577 ( .A1(n9850), .A2(n8462), .B1(n9845), .B2(n7990), .ZN(n7992)
         );
  NOR3_X1 U9578 ( .A1(n4343), .A2(n7992), .A3(n7991), .ZN(n7993) );
  AOI211_X1 U9579 ( .C1(n9854), .C2(n7995), .A(n7994), .B(n7993), .ZN(n7996)
         );
  OAI21_X1 U9580 ( .B1(n7997), .B2(n9835), .A(n7996), .ZN(P2_U3229) );
  INV_X1 U9581 ( .A(n9385), .ZN(n9274) );
  INV_X1 U9582 ( .A(n9405), .ZN(n8001) );
  OAI21_X1 U9583 ( .B1(n8001), .B2(n8000), .A(n9315), .ZN(n8002) );
  OAI21_X1 U9584 ( .B1(n9301), .B2(n9405), .A(n8002), .ZN(n9311) );
  NOR2_X1 U9585 ( .A1(n9391), .A2(n9300), .ZN(n8003) );
  NAND2_X1 U9586 ( .A1(n9254), .A2(n9255), .ZN(n8006) );
  NAND2_X1 U9587 ( .A1(n9382), .A2(n9276), .ZN(n8005) );
  INV_X1 U9588 ( .A(n9360), .ZN(n9202) );
  AOI22_X1 U9589 ( .A1(n9196), .A2(n9205), .B1(n9105), .B2(n9202), .ZN(n9185)
         );
  NAND2_X1 U9590 ( .A1(n4557), .A2(n9178), .ZN(n8008) );
  AOI22_X1 U9591 ( .A1(n9185), .A2(n8008), .B1(n9355), .B2(n9207), .ZN(n9169)
         );
  AOI22_X1 U9592 ( .A1(n9169), .A2(n9177), .B1(n9009), .B2(n9174), .ZN(n9156)
         );
  NAND2_X1 U9593 ( .A1(n9156), .A2(n9155), .ZN(n9154) );
  INV_X1 U9594 ( .A(P1_B_REG_SCAN_IN), .ZN(n8009) );
  OAI21_X1 U9595 ( .B1(n9546), .B2(n8009), .A(n9726), .ZN(n9143) );
  NOR2_X1 U9596 ( .A1(n8011), .A2(n8010), .ZN(n9317) );
  NAND2_X1 U9597 ( .A1(n9317), .A2(n8012), .ZN(n9297) );
  INV_X1 U9598 ( .A(n8018), .ZN(n8019) );
  AOI21_X1 U9599 ( .B1(n9256), .B2(n8020), .A(n8019), .ZN(n9248) );
  NAND3_X1 U9600 ( .A1(n9218), .A2(n8023), .A3(n9203), .ZN(n8025) );
  NAND2_X1 U9601 ( .A1(n8025), .A2(n8024), .ZN(n9189) );
  XNOR2_X1 U9602 ( .A(n8031), .B(n8030), .ZN(n8032) );
  OAI222_X1 U9603 ( .A1(n9699), .A2(n9179), .B1(n9143), .B2(n8033), .C1(n8032), 
        .C2(n9733), .ZN(n9339) );
  INV_X1 U9604 ( .A(n9337), .ZN(n8038) );
  NOR2_X1 U9605 ( .A1(n9322), .A2(n9405), .ZN(n9321) );
  INV_X1 U9606 ( .A(n9397), .ZN(n9305) );
  NAND2_X1 U9607 ( .A1(n9303), .A2(n9293), .ZN(n9287) );
  OR2_X2 U9608 ( .A1(n9287), .A2(n9385), .ZN(n9269) );
  NAND2_X1 U9609 ( .A1(n9213), .A2(n9202), .ZN(n9197) );
  INV_X1 U9610 ( .A(n9157), .ZN(n8034) );
  AOI211_X1 U9611 ( .C1(n9337), .C2(n8034), .A(n9801), .B(n4265), .ZN(n9338)
         );
  NAND2_X1 U9612 ( .A1(n9338), .A2(n9260), .ZN(n8037) );
  AOI22_X1 U9613 ( .A1(n9739), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n8035), .B2(
        n9718), .ZN(n8036) );
  OAI211_X1 U9614 ( .C1(n8038), .C2(n9710), .A(n8037), .B(n8036), .ZN(n8039)
         );
  AOI21_X1 U9615 ( .B1(n9339), .B2(n9737), .A(n8039), .ZN(n8040) );
  OAI21_X1 U9616 ( .B1(n9344), .B2(n9329), .A(n8040), .ZN(P1_U3355) );
  OAI222_X1 U9617 ( .A1(n8045), .A2(n8943), .B1(n8048), .B2(n8042), .C1(n8041), 
        .C2(P1_U3084), .ZN(P1_U3332) );
  OAI222_X1 U9618 ( .A1(n8045), .A2(n8948), .B1(n8048), .B2(n8044), .C1(
        P1_U3084), .C2(n8043), .ZN(P1_U3331) );
  INV_X1 U9619 ( .A(n8224), .ZN(n8092) );
  INV_X1 U9620 ( .A(n8144), .ZN(n8548) );
  INV_X1 U9621 ( .A(n8203), .ZN(n8452) );
  OR2_X1 U9622 ( .A1(n8787), .A2(n8452), .ZN(n8049) );
  NAND2_X1 U9623 ( .A1(n8050), .A2(n8049), .ZN(n8692) );
  NAND2_X1 U9624 ( .A1(n8783), .A2(n8155), .ZN(n8345) );
  NAND2_X1 U9625 ( .A1(n8339), .A2(n8345), .ZN(n8704) );
  INV_X1 U9626 ( .A(n8155), .ZN(n8451) );
  OR2_X1 U9627 ( .A1(n8783), .A2(n8451), .ZN(n8051) );
  NAND2_X1 U9628 ( .A1(n8778), .A2(n8657), .ZN(n8052) );
  OR2_X1 U9629 ( .A1(n8778), .A2(n8657), .ZN(n8053) );
  INV_X1 U9630 ( .A(n8647), .ZN(n8126) );
  NAND2_X1 U9631 ( .A1(n8771), .A2(n8126), .ZN(n8075) );
  OR2_X1 U9632 ( .A1(n8764), .A2(n8655), .ZN(n8055) );
  AND2_X1 U9633 ( .A1(n8764), .A2(n8655), .ZN(n8054) );
  NAND2_X1 U9634 ( .A1(n8759), .A2(n8104), .ZN(n8245) );
  NAND2_X1 U9635 ( .A1(n8076), .A2(n8245), .ZN(n8356) );
  NOR2_X1 U9636 ( .A1(n8759), .A2(n8648), .ZN(n8056) );
  AOI21_X1 U9637 ( .B1(n8624), .B2(n8356), .A(n8056), .ZN(n8603) );
  OR2_X1 U9638 ( .A1(n8618), .A2(n8057), .ZN(n8243) );
  NAND2_X1 U9639 ( .A1(n8618), .A2(n8057), .ZN(n8359) );
  NAND2_X1 U9640 ( .A1(n8243), .A2(n8359), .ZN(n8604) );
  INV_X1 U9641 ( .A(n8561), .ZN(n8450) );
  OR2_X1 U9642 ( .A1(n8737), .A2(n8144), .ZN(n8372) );
  NAND2_X1 U9643 ( .A1(n8737), .A2(n8144), .ZN(n8376) );
  NAND2_X1 U9644 ( .A1(n8372), .A2(n8376), .ZN(n8558) );
  NAND2_X1 U9645 ( .A1(n8555), .A2(n8558), .ZN(n8554) );
  OAI21_X1 U9646 ( .B1(n8548), .B2(n8737), .A(n8554), .ZN(n8537) );
  XNOR2_X1 U9647 ( .A(n8732), .B(n8563), .ZN(n8536) );
  NAND2_X1 U9648 ( .A1(n8725), .A2(n8096), .ZN(n8381) );
  INV_X1 U9649 ( .A(n8096), .ZN(n8549) );
  NAND2_X1 U9650 ( .A1(n8062), .A2(n4266), .ZN(n8064) );
  NAND2_X1 U9651 ( .A1(n5328), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8063) );
  OR2_X1 U9652 ( .A1(n8720), .A2(n8065), .ZN(n8386) );
  NAND2_X1 U9653 ( .A1(n8720), .A2(n8065), .ZN(n8387) );
  NAND2_X1 U9654 ( .A1(n8386), .A2(n8387), .ZN(n8430) );
  INV_X1 U9655 ( .A(n8783), .ZN(n8701) );
  INV_X1 U9656 ( .A(n8764), .ZN(n8644) );
  INV_X1 U9657 ( .A(n8759), .ZN(n8629) );
  INV_X1 U9658 ( .A(n8737), .ZN(n8067) );
  NAND2_X1 U9659 ( .A1(n8061), .A2(n8539), .ZN(n8522) );
  AOI21_X1 U9660 ( .B1(n8720), .B2(n8522), .A(n8513), .ZN(n8721) );
  INV_X1 U9661 ( .A(n8720), .ZN(n8070) );
  AOI22_X1 U9662 ( .A1(n8068), .A2(n8697), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n7135), .ZN(n8069) );
  OAI21_X1 U9663 ( .B1(n8070), .B2(n8700), .A(n8069), .ZN(n8089) );
  INV_X1 U9664 ( .A(n8339), .ZN(n8072) );
  OR2_X1 U9665 ( .A1(n8778), .A2(n8073), .ZN(n8348) );
  NAND2_X1 U9666 ( .A1(n8778), .A2(n8073), .ZN(n8346) );
  NAND2_X1 U9667 ( .A1(n8074), .A2(n8346), .ZN(n8653) );
  INV_X1 U9668 ( .A(n8075), .ZN(n8343) );
  XNOR2_X1 U9669 ( .A(n8764), .B(n8655), .ZN(n8646) );
  AND2_X1 U9670 ( .A1(n8764), .A2(n8350), .ZN(n8630) );
  NOR2_X1 U9671 ( .A1(n8356), .A2(n8630), .ZN(n8077) );
  INV_X1 U9672 ( .A(n8076), .ZN(n8246) );
  INV_X1 U9673 ( .A(n8604), .ZN(n8608) );
  INV_X1 U9674 ( .A(n8359), .ZN(n8589) );
  INV_X1 U9675 ( .A(n8363), .ZN(n8078) );
  OR2_X1 U9676 ( .A1(n8742), .A2(n8561), .ZN(n8371) );
  INV_X1 U9677 ( .A(n8376), .ZN(n8079) );
  INV_X1 U9678 ( .A(n8536), .ZN(n8546) );
  NAND2_X1 U9679 ( .A1(n8547), .A2(n8546), .ZN(n8545) );
  OR2_X1 U9680 ( .A1(n8732), .A2(n8563), .ZN(n8375) );
  NAND2_X1 U9681 ( .A1(n8545), .A2(n8375), .ZN(n8528) );
  INV_X1 U9682 ( .A(n8527), .ZN(n8428) );
  INV_X1 U9683 ( .A(n8380), .ZN(n8080) );
  OAI21_X1 U9684 ( .B1(n8081), .B2(n8066), .A(n8227), .ZN(n8087) );
  AOI21_X1 U9685 ( .B1(n8082), .B2(P2_B_REG_SCAN_IN), .A(n8564), .ZN(n8509) );
  INV_X1 U9686 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8942) );
  NAND2_X1 U9687 ( .A1(n4954), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8083) );
  OAI211_X1 U9688 ( .C1(n5000), .C2(n8942), .A(n8084), .B(n8083), .ZN(n8449)
         );
  AOI211_X1 U9689 ( .C1(n8721), .C2(n8669), .A(n8089), .B(n8088), .ZN(n8090)
         );
  OAI21_X1 U9690 ( .B1(n8724), .B2(n8711), .A(n8090), .ZN(P2_U3267) );
  OAI222_X1 U9691 ( .A1(n8975), .A2(n8092), .B1(n8091), .B2(n10007), .C1(n8865), .C2(n8971), .ZN(P2_U3328) );
  XNOR2_X1 U9692 ( .A(n8094), .B(n8093), .ZN(n8100) );
  OAI22_X1 U9693 ( .A1(n8542), .A2(n9860), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8095), .ZN(n8098) );
  OAI22_X1 U9694 ( .A1(n8096), .A2(n8219), .B1(n8144), .B2(n9831), .ZN(n8097)
         );
  AOI211_X1 U9695 ( .C1(n8732), .C2(n9854), .A(n8098), .B(n8097), .ZN(n8099)
         );
  OAI21_X1 U9696 ( .B1(n8100), .B2(n9835), .A(n8099), .ZN(P2_U3216) );
  INV_X1 U9697 ( .A(n8103), .ZN(n8102) );
  NOR2_X1 U9698 ( .A1(n8102), .A2(n8101), .ZN(n8162) );
  AOI22_X1 U9699 ( .A1(n8103), .A2(n9845), .B1(n9850), .B2(n8634), .ZN(n8110)
         );
  NOR2_X1 U9700 ( .A1(n8104), .A2(n8562), .ZN(n8105) );
  AOI21_X1 U9701 ( .B1(n4477), .B2(n8654), .A(n8105), .ZN(n8613) );
  OAI22_X1 U9702 ( .A1(n8613), .A2(n8209), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8106), .ZN(n8108) );
  INV_X1 U9703 ( .A(n8618), .ZN(n8753) );
  NOR2_X1 U9704 ( .A1(n8753), .A2(n8214), .ZN(n8107) );
  AOI211_X1 U9705 ( .C1(n8211), .C2(n8617), .A(n8108), .B(n8107), .ZN(n8109)
         );
  OAI21_X1 U9706 ( .B1(n8162), .B2(n8110), .A(n8109), .ZN(P2_U3218) );
  NAND3_X1 U9707 ( .A1(n8112), .A2(n9850), .A3(n8451), .ZN(n8113) );
  OAI21_X1 U9708 ( .B1(n8111), .B2(n9835), .A(n8113), .ZN(n8116) );
  INV_X1 U9709 ( .A(n8114), .ZN(n8115) );
  NAND2_X1 U9710 ( .A1(n8116), .A2(n8115), .ZN(n8121) );
  NOR2_X1 U9711 ( .A1(n9860), .A2(n8680), .ZN(n8119) );
  AOI22_X1 U9712 ( .A1(n8647), .A2(n8654), .B1(n8451), .B2(n8656), .ZN(n8686)
         );
  OAI22_X1 U9713 ( .A1(n8209), .A2(n8686), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8117), .ZN(n8118) );
  AOI211_X1 U9714 ( .C1(n8778), .C2(n9854), .A(n8119), .B(n8118), .ZN(n8120)
         );
  OAI211_X1 U9715 ( .C1(n9835), .C2(n8122), .A(n8121), .B(n8120), .ZN(P2_U3221) );
  INV_X1 U9716 ( .A(n8123), .ZN(n8124) );
  AOI21_X1 U9717 ( .B1(n8125), .B2(n8124), .A(n9835), .ZN(n8130) );
  NOR3_X1 U9718 ( .A1(n8127), .A2(n8126), .A3(n8202), .ZN(n8129) );
  OAI21_X1 U9719 ( .B1(n8130), .B2(n8129), .A(n8128), .ZN(n8134) );
  AOI22_X1 U9720 ( .A1(n8211), .A2(n8642), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        n10007), .ZN(n8133) );
  AOI22_X1 U9721 ( .A1(n8194), .A2(n8647), .B1(n9828), .B2(n8648), .ZN(n8132)
         );
  NAND2_X1 U9722 ( .A1(n8764), .A2(n9854), .ZN(n8131) );
  NAND4_X1 U9723 ( .A1(n8134), .A2(n8133), .A3(n8132), .A4(n8131), .ZN(
        P2_U3225) );
  INV_X1 U9724 ( .A(n8742), .ZN(n8150) );
  INV_X1 U9725 ( .A(n8139), .ZN(n8136) );
  NOR3_X1 U9726 ( .A1(n8136), .A2(n9835), .A3(n8135), .ZN(n8142) );
  NAND3_X1 U9727 ( .A1(n8137), .A2(n9850), .A3(n8450), .ZN(n8138) );
  OAI21_X1 U9728 ( .B1(n8139), .B2(n9835), .A(n8138), .ZN(n8141) );
  MUX2_X1 U9729 ( .A(n8142), .B(n8141), .S(n8140), .Z(n8143) );
  INV_X1 U9730 ( .A(n8143), .ZN(n8149) );
  OAI22_X1 U9731 ( .A1(n8144), .A2(n8564), .B1(n8165), .B2(n8562), .ZN(n8741)
         );
  INV_X1 U9732 ( .A(n8145), .ZN(n8578) );
  OAI22_X1 U9733 ( .A1(n8578), .A2(n9860), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8146), .ZN(n8147) );
  AOI21_X1 U9734 ( .B1(n8741), .B2(n9844), .A(n8147), .ZN(n8148) );
  OAI211_X1 U9735 ( .C1(n8150), .C2(n8214), .A(n8149), .B(n8148), .ZN(P2_U3227) );
  AOI21_X1 U9736 ( .B1(n8152), .B2(n8151), .A(n9835), .ZN(n8153) );
  NAND2_X1 U9737 ( .A1(n8153), .A2(n8201), .ZN(n8159) );
  AND2_X1 U9738 ( .A1(n10007), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9869) );
  OAI22_X1 U9739 ( .A1(n8155), .A2(n8219), .B1(n9831), .B2(n8154), .ZN(n8156)
         );
  AOI211_X1 U9740 ( .C1(n8211), .C2(n8157), .A(n9869), .B(n8156), .ZN(n8158)
         );
  OAI211_X1 U9741 ( .C1(n8160), .C2(n8214), .A(n8159), .B(n8158), .ZN(P2_U3230) );
  NOR2_X1 U9742 ( .A1(n8162), .A2(n8161), .ZN(n8164) );
  XNOR2_X1 U9743 ( .A(n8164), .B(n8163), .ZN(n8168) );
  OAI22_X1 U9744 ( .A1(n8168), .A2(n9835), .B1(n8165), .B2(n8202), .ZN(n8166)
         );
  OAI21_X1 U9745 ( .B1(n8168), .B2(n8167), .A(n8166), .ZN(n8174) );
  OR2_X1 U9746 ( .A1(n8561), .A2(n8564), .ZN(n8170) );
  NAND2_X1 U9747 ( .A1(n8634), .A2(n8656), .ZN(n8169) );
  NAND2_X1 U9748 ( .A1(n8170), .A2(n8169), .ZN(n8590) );
  OAI22_X1 U9749 ( .A1(n8598), .A2(n9860), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8171), .ZN(n8172) );
  AOI21_X1 U9750 ( .B1(n8590), .B2(n9844), .A(n8172), .ZN(n8173) );
  OAI211_X1 U9751 ( .C1(n4478), .C2(n8214), .A(n8174), .B(n8173), .ZN(P2_U3231) );
  OAI21_X1 U9752 ( .B1(n8184), .B2(n9855), .A(n8175), .ZN(n8176) );
  NAND2_X1 U9753 ( .A1(n8176), .A2(n9845), .ZN(n8188) );
  NAND2_X1 U9754 ( .A1(n8211), .A2(n8177), .ZN(n8178) );
  OAI211_X1 U9755 ( .C1(n8219), .C2(n8180), .A(n8179), .B(n8178), .ZN(n8181)
         );
  AOI21_X1 U9756 ( .B1(n9854), .B2(n8182), .A(n8181), .ZN(n8187) );
  NOR3_X1 U9757 ( .A1(n8184), .A2(n8202), .A3(n8183), .ZN(n8185) );
  OAI21_X1 U9758 ( .B1(n8185), .B2(n8194), .A(n8459), .ZN(n8186) );
  NAND3_X1 U9759 ( .A1(n8188), .A2(n8187), .A3(n8186), .ZN(P2_U3233) );
  NAND2_X1 U9760 ( .A1(n9850), .A2(n8648), .ZN(n8192) );
  NAND2_X1 U9761 ( .A1(n8189), .A2(n9845), .ZN(n8191) );
  MUX2_X1 U9762 ( .A(n8192), .B(n8191), .S(n8190), .Z(n8198) );
  INV_X1 U9763 ( .A(n8193), .ZN(n8627) );
  AOI22_X1 U9764 ( .A1(n8211), .A2(n8627), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8197) );
  AOI22_X1 U9765 ( .A1(n9828), .A2(n8634), .B1(n8194), .B2(n8655), .ZN(n8196)
         );
  NAND2_X1 U9766 ( .A1(n8759), .A2(n9854), .ZN(n8195) );
  NAND4_X1 U9767 ( .A1(n8198), .A2(n8197), .A3(n8196), .A4(n8195), .ZN(
        P2_U3237) );
  INV_X1 U9768 ( .A(n8199), .ZN(n8200) );
  AOI21_X1 U9769 ( .B1(n8201), .B2(n8200), .A(n9835), .ZN(n8206) );
  NOR3_X1 U9770 ( .A1(n8204), .A2(n8203), .A3(n8202), .ZN(n8205) );
  OAI21_X1 U9771 ( .B1(n8206), .B2(n8205), .A(n8111), .ZN(n8213) );
  INV_X1 U9772 ( .A(n8207), .ZN(n8698) );
  AOI22_X1 U9773 ( .A1(n8452), .A2(n8656), .B1(n8657), .B2(n8654), .ZN(n8706)
         );
  OAI22_X1 U9774 ( .A1(n8209), .A2(n8706), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8208), .ZN(n8210) );
  AOI21_X1 U9775 ( .B1(n8698), .B2(n8211), .A(n8210), .ZN(n8212) );
  OAI211_X1 U9776 ( .C1(n8701), .C2(n8214), .A(n8213), .B(n8212), .ZN(P2_U3240) );
  XNOR2_X1 U9777 ( .A(n8216), .B(n8215), .ZN(n8223) );
  INV_X1 U9778 ( .A(n8217), .ZN(n8568) );
  OAI22_X1 U9779 ( .A1(n8568), .A2(n9860), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8218), .ZN(n8221) );
  OAI22_X1 U9780 ( .A1(n8563), .A2(n8219), .B1(n8561), .B2(n9831), .ZN(n8220)
         );
  AOI211_X1 U9781 ( .C1(n8737), .C2(n9854), .A(n8221), .B(n8220), .ZN(n8222)
         );
  OAI21_X1 U9782 ( .B1(n8223), .B2(n9835), .A(n8222), .ZN(P2_U3242) );
  NAND2_X1 U9783 ( .A1(n8224), .A2(n8231), .ZN(n8226) );
  NAND2_X1 U9784 ( .A1(n4902), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8225) );
  INV_X1 U9785 ( .A(n8449), .ZN(n8235) );
  NOR2_X1 U9786 ( .A1(n8515), .A2(n8235), .ZN(n8384) );
  AOI21_X1 U9787 ( .B1(n8227), .B2(n8387), .A(n8384), .ZN(n8230) );
  NOR2_X1 U9788 ( .A1(n8508), .A2(n8436), .ZN(n8229) );
  NAND3_X1 U9789 ( .A1(n8227), .A2(n8719), .A3(n8387), .ZN(n8228) );
  NAND2_X1 U9790 ( .A1(n9448), .A2(n8231), .ZN(n8233) );
  NAND2_X1 U9791 ( .A1(n5328), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8232) );
  INV_X1 U9792 ( .A(n8508), .ZN(n8234) );
  OR2_X1 U9793 ( .A1(n8712), .A2(n8234), .ZN(n8392) );
  NAND2_X1 U9794 ( .A1(n8515), .A2(n8235), .ZN(n8389) );
  INV_X1 U9795 ( .A(n8712), .ZN(n8510) );
  NOR2_X1 U9796 ( .A1(n8510), .A2(n8508), .ZN(n8395) );
  XNOR2_X1 U9797 ( .A(n8237), .B(n8569), .ZN(n8238) );
  AOI21_X1 U9798 ( .B1(n8240), .B2(n8239), .A(n8238), .ZN(n8440) );
  NOR2_X1 U9799 ( .A1(n8395), .A2(n8384), .ZN(n8401) );
  NAND2_X2 U9800 ( .A1(n8242), .A2(n8241), .ZN(n8393) );
  MUX2_X1 U9801 ( .A(n8400), .B(n8401), .S(n8393), .Z(n8398) );
  INV_X1 U9802 ( .A(n8243), .ZN(n8244) );
  NOR2_X1 U9803 ( .A1(n8358), .A2(n8245), .ZN(n8247) );
  MUX2_X1 U9804 ( .A(n8247), .B(n8246), .S(n8393), .Z(n8362) );
  NAND2_X1 U9805 ( .A1(n8269), .A2(n8249), .ZN(n8254) );
  NAND2_X1 U9806 ( .A1(n8251), .A2(n8250), .ZN(n8253) );
  INV_X1 U9807 ( .A(n8279), .ZN(n8252) );
  AOI21_X1 U9808 ( .B1(n8254), .B2(n8253), .A(n8252), .ZN(n8282) );
  NAND2_X1 U9809 ( .A1(n8465), .A2(n9907), .ZN(n8263) );
  NAND2_X1 U9810 ( .A1(n8256), .A2(n8263), .ZN(n8259) );
  NAND2_X1 U9811 ( .A1(n8256), .A2(n8255), .ZN(n8257) );
  NAND2_X1 U9812 ( .A1(n8257), .A2(n8273), .ZN(n8258) );
  MUX2_X1 U9813 ( .A(n8259), .B(n8258), .S(n8393), .Z(n8262) );
  AND2_X1 U9814 ( .A1(n8260), .A2(n8436), .ZN(n8261) );
  NOR2_X1 U9815 ( .A1(n8262), .A2(n8261), .ZN(n8277) );
  NAND2_X1 U9816 ( .A1(n8275), .A2(n8263), .ZN(n8264) );
  OAI211_X1 U9817 ( .C1(n8277), .C2(n8264), .A(n8274), .B(n8393), .ZN(n8266)
         );
  NAND3_X1 U9818 ( .A1(n8266), .A2(n8265), .A3(n8405), .ZN(n8272) );
  OAI211_X1 U9819 ( .C1(n8269), .C2(n8268), .A(n8285), .B(n8267), .ZN(n8270)
         );
  NAND2_X1 U9820 ( .A1(n8270), .A2(n8393), .ZN(n8271) );
  NAND2_X1 U9821 ( .A1(n8272), .A2(n8271), .ZN(n8280) );
  NAND2_X1 U9822 ( .A1(n8274), .A2(n8273), .ZN(n8276) );
  OAI211_X1 U9823 ( .C1(n8277), .C2(n8276), .A(n8385), .B(n8275), .ZN(n8278)
         );
  NAND3_X1 U9824 ( .A1(n8280), .A2(n8279), .A3(n8278), .ZN(n8281) );
  OAI21_X1 U9825 ( .B1(n8282), .B2(n8393), .A(n8281), .ZN(n8284) );
  OAI211_X1 U9826 ( .C1(n8285), .C2(n8393), .A(n8284), .B(n4267), .ZN(n8289)
         );
  MUX2_X1 U9827 ( .A(n8287), .B(n8286), .S(n8393), .Z(n8288) );
  NAND3_X1 U9828 ( .A1(n8289), .A2(n8410), .A3(n8288), .ZN(n8293) );
  MUX2_X1 U9829 ( .A(n8291), .B(n8290), .S(n8393), .Z(n8292) );
  NAND3_X1 U9830 ( .A1(n8293), .A2(n8411), .A3(n8292), .ZN(n8299) );
  AND2_X1 U9831 ( .A1(n8300), .A2(n8294), .ZN(n8295) );
  MUX2_X1 U9832 ( .A(n8296), .B(n8295), .S(n8393), .Z(n8297) );
  NAND3_X1 U9833 ( .A1(n8299), .A2(n8298), .A3(n8297), .ZN(n8304) );
  AND2_X1 U9834 ( .A1(n8308), .A2(n8300), .ZN(n8302) );
  MUX2_X1 U9835 ( .A(n8302), .B(n8301), .S(n8393), .Z(n8303) );
  NAND2_X1 U9836 ( .A1(n8304), .A2(n8303), .ZN(n8311) );
  AND2_X1 U9837 ( .A1(n8416), .A2(n8305), .ZN(n8307) );
  INV_X1 U9838 ( .A(n8417), .ZN(n8306) );
  AOI21_X1 U9839 ( .B1(n8311), .B2(n8307), .A(n8306), .ZN(n8313) );
  AND2_X1 U9840 ( .A1(n8417), .A2(n8308), .ZN(n8310) );
  INV_X1 U9841 ( .A(n8416), .ZN(n8309) );
  AOI21_X1 U9842 ( .B1(n8311), .B2(n8310), .A(n8309), .ZN(n8312) );
  MUX2_X1 U9843 ( .A(n8313), .B(n8312), .S(n8393), .Z(n8314) );
  NAND2_X1 U9844 ( .A1(n8314), .A2(n8419), .ZN(n8318) );
  MUX2_X1 U9845 ( .A(n8316), .B(n8315), .S(n8393), .Z(n8317) );
  MUX2_X1 U9846 ( .A(n8320), .B(n8319), .S(n8385), .Z(n8325) );
  MUX2_X1 U9847 ( .A(n8454), .B(n9476), .S(n8393), .Z(n8321) );
  INV_X1 U9848 ( .A(n8333), .ZN(n8323) );
  INV_X1 U9849 ( .A(n8330), .ZN(n8322) );
  NAND2_X1 U9850 ( .A1(n8331), .A2(n8326), .ZN(n8328) );
  NAND2_X1 U9851 ( .A1(n8329), .A2(n8327), .ZN(n8332) );
  MUX2_X1 U9852 ( .A(n8328), .B(n8332), .S(n8393), .Z(n8338) );
  OAI211_X1 U9853 ( .C1(n8338), .C2(n8330), .A(n8345), .B(n8329), .ZN(n8335)
         );
  OAI211_X1 U9854 ( .C1(n8333), .C2(n8332), .A(n8339), .B(n8331), .ZN(n8334)
         );
  MUX2_X1 U9855 ( .A(n8335), .B(n8334), .S(n8393), .Z(n8336) );
  INV_X1 U9856 ( .A(n8336), .ZN(n8337) );
  NAND3_X1 U9857 ( .A1(n8347), .A2(n8339), .A3(n8348), .ZN(n8340) );
  NAND2_X1 U9858 ( .A1(n8340), .A2(n8346), .ZN(n8342) );
  OR2_X1 U9859 ( .A1(n8630), .A2(n8393), .ZN(n8341) );
  AOI21_X1 U9860 ( .B1(n8342), .B2(n8352), .A(n8341), .ZN(n8344) );
  NAND3_X1 U9861 ( .A1(n8347), .A2(n8346), .A3(n8345), .ZN(n8349) );
  NAND3_X1 U9862 ( .A1(n8349), .A2(n8348), .A3(n8393), .ZN(n8351) );
  OR2_X1 U9863 ( .A1(n8764), .A2(n8350), .ZN(n8353) );
  NAND2_X1 U9864 ( .A1(n8351), .A2(n8353), .ZN(n8355) );
  AND2_X1 U9865 ( .A1(n8353), .A2(n8352), .ZN(n8354) );
  NAND2_X1 U9866 ( .A1(n8630), .A2(n8393), .ZN(n8357) );
  AND2_X1 U9867 ( .A1(n8364), .A2(n8359), .ZN(n8360) );
  OAI22_X1 U9868 ( .A1(n8362), .A2(n8361), .B1(n8385), .B2(n8360), .ZN(n8366)
         );
  MUX2_X1 U9869 ( .A(n8364), .B(n8363), .S(n8393), .Z(n8365) );
  NAND3_X1 U9870 ( .A1(n8366), .A2(n4359), .A3(n8365), .ZN(n8369) );
  AND2_X1 U9871 ( .A1(n8742), .A2(n8561), .ZN(n8367) );
  OAI21_X1 U9872 ( .B1(n8558), .B2(n8367), .A(n8393), .ZN(n8368) );
  NAND2_X1 U9873 ( .A1(n8369), .A2(n8368), .ZN(n8370) );
  NAND2_X1 U9874 ( .A1(n8372), .A2(n8371), .ZN(n8373) );
  NAND2_X1 U9875 ( .A1(n8373), .A2(n8385), .ZN(n8374) );
  NAND3_X1 U9876 ( .A1(n8377), .A2(n8546), .A3(n8376), .ZN(n8378) );
  NAND3_X1 U9877 ( .A1(n8379), .A2(n8428), .A3(n8378), .ZN(n8383) );
  MUX2_X1 U9878 ( .A(n8381), .B(n8380), .S(n8393), .Z(n8382) );
  NAND3_X1 U9879 ( .A1(n8383), .A2(n8066), .A3(n8382), .ZN(n8391) );
  INV_X1 U9880 ( .A(n8384), .ZN(n8390) );
  MUX2_X1 U9881 ( .A(n8387), .B(n8386), .S(n8385), .Z(n8388) );
  NAND4_X1 U9882 ( .A1(n8391), .A2(n8390), .A3(n8389), .A4(n8388), .ZN(n8397)
         );
  INV_X1 U9883 ( .A(n8392), .ZN(n8394) );
  MUX2_X1 U9884 ( .A(n8395), .B(n8394), .S(n8393), .Z(n8396) );
  AOI211_X1 U9885 ( .C1(n8399), .C2(n8434), .A(n5535), .B(n8435), .ZN(n8438)
         );
  INV_X1 U9886 ( .A(n8400), .ZN(n8432) );
  INV_X1 U9887 ( .A(n8401), .ZN(n8431) );
  INV_X1 U9888 ( .A(n8674), .ZN(n8684) );
  NOR2_X1 U9889 ( .A1(n8402), .A2(n9900), .ZN(n8404) );
  NAND4_X1 U9890 ( .A1(n8405), .A2(n8404), .A3(n5535), .A4(n8403), .ZN(n8409)
         );
  NOR4_X1 U9891 ( .A1(n8409), .A2(n8408), .A3(n8407), .A4(n8406), .ZN(n8412)
         );
  NAND4_X1 U9892 ( .A1(n8412), .A2(n4267), .A3(n8411), .A4(n8410), .ZN(n8415)
         );
  NOR3_X1 U9893 ( .A1(n8415), .A2(n7070), .A3(n8414), .ZN(n8418) );
  NAND4_X1 U9894 ( .A1(n8419), .A2(n8418), .A3(n8417), .A4(n8416), .ZN(n8420)
         );
  OR4_X1 U9895 ( .A1(n8423), .A2(n8422), .A3(n8421), .A4(n8420), .ZN(n8424) );
  NOR4_X1 U9896 ( .A1(n8684), .A2(n4582), .A3(n8704), .A4(n8424), .ZN(n8425)
         );
  NAND4_X1 U9897 ( .A1(n8632), .A2(n8660), .A3(n8425), .A4(n8646), .ZN(n8426)
         );
  NOR4_X1 U9898 ( .A1(n8558), .A2(n8604), .A3(n8594), .A4(n8426), .ZN(n8427)
         );
  NAND4_X1 U9899 ( .A1(n8428), .A2(n8427), .A3(n8546), .A4(n4359), .ZN(n8429)
         );
  NOR4_X1 U9900 ( .A1(n8432), .A2(n8431), .A3(n8430), .A4(n8429), .ZN(n8433)
         );
  XNOR2_X1 U9901 ( .A(n8433), .B(n8583), .ZN(n8437) );
  NOR2_X1 U9902 ( .A1(n8440), .A2(n8439), .ZN(n8448) );
  INV_X1 U9903 ( .A(n9886), .ZN(n8443) );
  NOR4_X1 U9904 ( .A1(n8443), .A2(n8442), .A3(n8441), .A4(n8562), .ZN(n8446)
         );
  OAI21_X1 U9905 ( .B1(n8447), .B2(n8444), .A(P2_B_REG_SCAN_IN), .ZN(n8445) );
  OAI22_X1 U9906 ( .A1(n8448), .A2(n8447), .B1(n8446), .B2(n8445), .ZN(
        P2_U3244) );
  MUX2_X1 U9907 ( .A(n8449), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8466), .Z(
        P2_U3582) );
  MUX2_X1 U9908 ( .A(n8529), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8466), .Z(
        P2_U3581) );
  MUX2_X1 U9909 ( .A(n8549), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8466), .Z(
        P2_U3580) );
  MUX2_X1 U9910 ( .A(n8530), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8466), .Z(
        P2_U3579) );
  MUX2_X1 U9911 ( .A(n8548), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8466), .Z(
        P2_U3578) );
  MUX2_X1 U9912 ( .A(n8450), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8466), .Z(
        P2_U3577) );
  MUX2_X1 U9913 ( .A(n4477), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8466), .Z(
        P2_U3576) );
  MUX2_X1 U9914 ( .A(n8634), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8466), .Z(
        P2_U3575) );
  MUX2_X1 U9915 ( .A(n8648), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8466), .Z(
        P2_U3574) );
  MUX2_X1 U9916 ( .A(n8655), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8466), .Z(
        P2_U3573) );
  MUX2_X1 U9917 ( .A(n8647), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8466), .Z(
        P2_U3572) );
  MUX2_X1 U9918 ( .A(n8657), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8466), .Z(
        P2_U3571) );
  MUX2_X1 U9919 ( .A(n8451), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8466), .Z(
        P2_U3570) );
  MUX2_X1 U9920 ( .A(n8452), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8466), .Z(
        P2_U3569) );
  MUX2_X1 U9921 ( .A(n8453), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8466), .Z(
        P2_U3568) );
  MUX2_X1 U9922 ( .A(n8454), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8466), .Z(
        P2_U3566) );
  MUX2_X1 U9923 ( .A(n8455), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8466), .Z(
        P2_U3565) );
  MUX2_X1 U9924 ( .A(n8456), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8466), .Z(
        P2_U3564) );
  MUX2_X1 U9925 ( .A(n9827), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8466), .Z(
        P2_U3563) );
  MUX2_X1 U9926 ( .A(n8457), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8466), .Z(
        P2_U3562) );
  MUX2_X1 U9927 ( .A(n8458), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8466), .Z(
        P2_U3561) );
  MUX2_X1 U9928 ( .A(n8459), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8466), .Z(
        P2_U3560) );
  MUX2_X1 U9929 ( .A(n9848), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8466), .Z(
        P2_U3559) );
  MUX2_X1 U9930 ( .A(n8460), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8466), .Z(
        P2_U3558) );
  MUX2_X1 U9931 ( .A(n8461), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8466), .Z(
        P2_U3557) );
  MUX2_X1 U9932 ( .A(n8462), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8466), .Z(
        P2_U3556) );
  MUX2_X1 U9933 ( .A(n8463), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8466), .Z(
        P2_U3555) );
  MUX2_X1 U9934 ( .A(n8464), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8466), .Z(
        P2_U3554) );
  MUX2_X1 U9935 ( .A(n8465), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8466), .Z(
        P2_U3553) );
  MUX2_X1 U9936 ( .A(n8467), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8466), .Z(
        P2_U3552) );
  NAND2_X1 U9937 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8477), .ZN(n8469) );
  NAND2_X1 U9938 ( .A1(n8469), .A2(n8468), .ZN(n9877) );
  INV_X1 U9939 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8470) );
  XNOR2_X1 U9940 ( .A(n9875), .B(n8470), .ZN(n9878) );
  NAND2_X1 U9941 ( .A1(n9877), .A2(n9878), .ZN(n8472) );
  NAND2_X1 U9942 ( .A1(n9875), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8471) );
  NAND2_X1 U9943 ( .A1(n8472), .A2(n8471), .ZN(n8473) );
  AOI21_X1 U9944 ( .B1(n8474), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8493), .ZN(
        n8491) );
  NAND2_X1 U9945 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(n10007), .ZN(n8475) );
  OAI21_X1 U9946 ( .B1(n8506), .B2(n9992), .A(n8475), .ZN(n8476) );
  AOI21_X1 U9947 ( .B1(n9876), .B2(n8480), .A(n8476), .ZN(n8489) );
  NOR2_X1 U9948 ( .A1(n8477), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8478) );
  INV_X1 U9949 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8793) );
  XNOR2_X1 U9950 ( .A(n9875), .B(n8793), .ZN(n9873) );
  NAND2_X1 U9951 ( .A1(n9874), .A2(n9873), .ZN(n9872) );
  INV_X1 U9952 ( .A(n9872), .ZN(n8482) );
  AND2_X1 U9953 ( .A1(n9875), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8483) );
  OR2_X1 U9954 ( .A1(n8480), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8495) );
  NAND2_X1 U9955 ( .A1(n8480), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8481) );
  NAND2_X1 U9956 ( .A1(n8495), .A2(n8481), .ZN(n8484) );
  OAI21_X1 U9957 ( .B1(n8482), .B2(n8483), .A(n8484), .ZN(n8486) );
  NOR2_X1 U9958 ( .A1(n8484), .A2(n8483), .ZN(n8485) );
  NAND2_X1 U9959 ( .A1(n9872), .A2(n8485), .ZN(n8496) );
  NAND2_X1 U9960 ( .A1(n8486), .A2(n8496), .ZN(n8487) );
  NAND2_X1 U9961 ( .A1(n8487), .A2(n9871), .ZN(n8488) );
  OAI211_X1 U9962 ( .C1(n8491), .C2(n8490), .A(n8489), .B(n8488), .ZN(P2_U3263) );
  NOR2_X1 U9963 ( .A1(n8493), .A2(n8492), .ZN(n8494) );
  XOR2_X1 U9964 ( .A(n8494), .B(P2_REG2_REG_19__SCAN_IN), .Z(n8503) );
  NAND2_X1 U9965 ( .A1(n8496), .A2(n8495), .ZN(n8498) );
  INV_X1 U9966 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8497) );
  XNOR2_X1 U9967 ( .A(n8498), .B(n8497), .ZN(n8501) );
  AOI21_X1 U9968 ( .B1(n8501), .B2(n9871), .A(n9876), .ZN(n8499) );
  INV_X1 U9969 ( .A(n8501), .ZN(n8502) );
  AOI22_X1 U9970 ( .A1(n8503), .A2(n9879), .B1(n9871), .B2(n8502), .ZN(n8504)
         );
  NAND2_X1 U9971 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n8505) );
  NAND2_X1 U9972 ( .A1(n8719), .A2(n8513), .ZN(n8716) );
  XNOR2_X1 U9973 ( .A(n8716), .B(n8712), .ZN(n8714) );
  NAND2_X1 U9974 ( .A1(n8509), .A2(n8508), .ZN(n8717) );
  NOR2_X1 U9975 ( .A1(n7135), .A2(n8717), .ZN(n8516) );
  NOR2_X1 U9976 ( .A1(n8510), .A2(n8700), .ZN(n8511) );
  AOI211_X1 U9977 ( .C1(n7135), .C2(P2_REG2_REG_31__SCAN_IN), .A(n8516), .B(
        n8511), .ZN(n8512) );
  OAI21_X1 U9978 ( .B1(n8714), .B2(n8621), .A(n8512), .ZN(P2_U3265) );
  INV_X1 U9979 ( .A(n8513), .ZN(n8514) );
  NAND2_X1 U9980 ( .A1(n8515), .A2(n8514), .ZN(n8715) );
  NAND3_X1 U9981 ( .A1(n8716), .A2(n8669), .A3(n8715), .ZN(n8518) );
  AOI21_X1 U9982 ( .B1(n7135), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8516), .ZN(
        n8517) );
  OAI211_X1 U9983 ( .C1(n8719), .C2(n8700), .A(n8518), .B(n8517), .ZN(P2_U3266) );
  OAI21_X1 U9984 ( .B1(n8520), .B2(n8527), .A(n8519), .ZN(n8521) );
  INV_X1 U9985 ( .A(n8521), .ZN(n8729) );
  INV_X1 U9986 ( .A(n8539), .ZN(n8524) );
  INV_X1 U9987 ( .A(n8522), .ZN(n8523) );
  AOI21_X1 U9988 ( .B1(n8725), .B2(n8524), .A(n8523), .ZN(n8726) );
  AOI22_X1 U9989 ( .A1(n8525), .A2(n8697), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n7135), .ZN(n8526) );
  OAI21_X1 U9990 ( .B1(n8061), .B2(n8700), .A(n8526), .ZN(n8533) );
  XNOR2_X1 U9991 ( .A(n8528), .B(n8527), .ZN(n8531) );
  AOI222_X1 U9992 ( .A1(n8659), .A2(n8531), .B1(n8530), .B2(n8656), .C1(n8529), 
        .C2(n8654), .ZN(n8728) );
  NOR2_X1 U9993 ( .A1(n8728), .A2(n7135), .ZN(n8532) );
  AOI211_X1 U9994 ( .C1(n8726), .C2(n8669), .A(n8533), .B(n8532), .ZN(n8534)
         );
  OAI21_X1 U9995 ( .B1(n8729), .B2(n8711), .A(n8534), .ZN(P2_U3268) );
  OAI21_X1 U9996 ( .B1(n8537), .B2(n8536), .A(n8535), .ZN(n8538) );
  INV_X1 U9997 ( .A(n8538), .ZN(n8734) );
  AOI211_X1 U9998 ( .C1(n8732), .C2(n8565), .A(n9936), .B(n8539), .ZN(n8731)
         );
  INV_X1 U9999 ( .A(n8732), .ZN(n8540) );
  NOR2_X1 U10000 ( .A1(n8540), .A2(n8700), .ZN(n8544) );
  OAI22_X1 U10001 ( .A1(n8542), .A2(n8679), .B1(n8541), .B2(n8688), .ZN(n8543)
         );
  AOI211_X1 U10002 ( .C1(n8731), .C2(n8703), .A(n8544), .B(n8543), .ZN(n8553)
         );
  OAI211_X1 U10003 ( .C1(n8547), .C2(n8546), .A(n8545), .B(n8659), .ZN(n8551)
         );
  AOI22_X1 U10004 ( .A1(n8549), .A2(n8654), .B1(n8656), .B2(n8548), .ZN(n8550)
         );
  NAND2_X1 U10005 ( .A1(n8551), .A2(n8550), .ZN(n8730) );
  NAND2_X1 U10006 ( .A1(n8730), .A2(n8688), .ZN(n8552) );
  OAI211_X1 U10007 ( .C1(n8734), .C2(n8711), .A(n8553), .B(n8552), .ZN(
        P2_U3269) );
  OAI21_X1 U10008 ( .B1(n8555), .B2(n8558), .A(n8554), .ZN(n8556) );
  INV_X1 U10009 ( .A(n8556), .ZN(n8739) );
  AOI22_X1 U10010 ( .A1(n8737), .A2(n8666), .B1(n7135), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8573) );
  AOI21_X1 U10011 ( .B1(n8559), .B2(n8558), .A(n8557), .ZN(n8560) );
  OAI222_X1 U10012 ( .A1(n8564), .A2(n8563), .B1(n8562), .B2(n8561), .C1(n8707), .C2(n8560), .ZN(n8735) );
  INV_X1 U10013 ( .A(n8582), .ZN(n8567) );
  INV_X1 U10014 ( .A(n8565), .ZN(n8566) );
  AOI211_X1 U10015 ( .C1(n8737), .C2(n8567), .A(n9936), .B(n8566), .ZN(n8736)
         );
  INV_X1 U10016 ( .A(n8736), .ZN(n8570) );
  OAI22_X1 U10017 ( .A1(n8570), .A2(n8569), .B1(n8679), .B2(n8568), .ZN(n8571)
         );
  OAI21_X1 U10018 ( .B1(n8735), .B2(n8571), .A(n8688), .ZN(n8572) );
  OAI211_X1 U10019 ( .C1(n8739), .C2(n8711), .A(n8573), .B(n8572), .ZN(
        P2_U3270) );
  OAI21_X1 U10020 ( .B1(n8576), .B2(n8575), .A(n8574), .ZN(n8577) );
  INV_X1 U10021 ( .A(n8577), .ZN(n8745) );
  OAI22_X1 U10022 ( .A1(n8578), .A2(n8679), .B1(n8882), .B2(n8688), .ZN(n8586)
         );
  XNOR2_X1 U10023 ( .A(n4289), .B(n4359), .ZN(n8579) );
  NAND2_X1 U10024 ( .A1(n8579), .A2(n8659), .ZN(n8743) );
  NAND2_X1 U10025 ( .A1(n8742), .A2(n8595), .ZN(n8580) );
  NAND2_X1 U10026 ( .A1(n8580), .A2(n9912), .ZN(n8581) );
  NOR2_X1 U10027 ( .A1(n8582), .A2(n8581), .ZN(n8740) );
  AOI21_X1 U10028 ( .B1(n8740), .B2(n8583), .A(n8741), .ZN(n8584) );
  AOI21_X1 U10029 ( .B1(n8743), .B2(n8584), .A(n7135), .ZN(n8585) );
  AOI211_X1 U10030 ( .C1(n8666), .C2(n8742), .A(n8586), .B(n8585), .ZN(n8587)
         );
  OAI21_X1 U10031 ( .B1(n8745), .B2(n8711), .A(n8587), .ZN(P2_U3271) );
  NOR2_X1 U10032 ( .A1(n8588), .A2(n8707), .ZN(n8592) );
  OAI21_X1 U10033 ( .B1(n8611), .B2(n8589), .A(n8594), .ZN(n8591) );
  AOI21_X1 U10034 ( .B1(n8592), .B2(n8591), .A(n8590), .ZN(n8750) );
  OAI21_X1 U10035 ( .B1(n4294), .B2(n8594), .A(n8593), .ZN(n8746) );
  NAND2_X1 U10036 ( .A1(n8746), .A2(n8662), .ZN(n8602) );
  INV_X1 U10037 ( .A(n8595), .ZN(n8596) );
  AOI21_X1 U10038 ( .B1(n8747), .B2(n8616), .A(n8596), .ZN(n8748) );
  NOR2_X1 U10039 ( .A1(n4478), .A2(n8700), .ZN(n8600) );
  OAI22_X1 U10040 ( .A1(n8598), .A2(n8679), .B1(n8688), .B2(n8597), .ZN(n8599)
         );
  AOI211_X1 U10041 ( .C1(n8748), .C2(n8669), .A(n8600), .B(n8599), .ZN(n8601)
         );
  OAI211_X1 U10042 ( .C1(n7135), .C2(n8750), .A(n8602), .B(n8601), .ZN(
        P2_U3272) );
  NOR2_X1 U10043 ( .A1(n8605), .A2(n8604), .ZN(n8606) );
  OR2_X1 U10044 ( .A1(n8607), .A2(n8606), .ZN(n8752) );
  NOR2_X1 U10045 ( .A1(n8609), .A2(n8608), .ZN(n8610) );
  OR2_X1 U10046 ( .A1(n8611), .A2(n8610), .ZN(n8612) );
  NAND2_X1 U10047 ( .A1(n8612), .A2(n8659), .ZN(n8614) );
  NAND2_X1 U10048 ( .A1(n8614), .A2(n8613), .ZN(n8756) );
  NAND2_X1 U10049 ( .A1(n8625), .A2(n8618), .ZN(n8615) );
  NAND2_X1 U10050 ( .A1(n8616), .A2(n8615), .ZN(n8754) );
  AOI22_X1 U10051 ( .A1(n7135), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8617), .B2(
        n8697), .ZN(n8620) );
  NAND2_X1 U10052 ( .A1(n8618), .A2(n8666), .ZN(n8619) );
  OAI211_X1 U10053 ( .C1(n8754), .C2(n8621), .A(n8620), .B(n8619), .ZN(n8622)
         );
  AOI21_X1 U10054 ( .B1(n8756), .B2(n8688), .A(n8622), .ZN(n8623) );
  OAI21_X1 U10055 ( .B1(n8752), .B2(n8711), .A(n8623), .ZN(P2_U3273) );
  XNOR2_X1 U10056 ( .A(n8624), .B(n8632), .ZN(n8763) );
  INV_X1 U10057 ( .A(n8640), .ZN(n8626) );
  AOI21_X1 U10058 ( .B1(n8759), .B2(n8626), .A(n4415), .ZN(n8760) );
  AOI22_X1 U10059 ( .A1(n7135), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8627), .B2(
        n8697), .ZN(n8628) );
  OAI21_X1 U10060 ( .B1(n8629), .B2(n8700), .A(n8628), .ZN(n8637) );
  INV_X1 U10061 ( .A(n8630), .ZN(n8631) );
  NAND2_X1 U10062 ( .A1(n8645), .A2(n8631), .ZN(n8633) );
  XNOR2_X1 U10063 ( .A(n8633), .B(n8632), .ZN(n8635) );
  AOI222_X1 U10064 ( .A1(n8659), .A2(n8635), .B1(n8655), .B2(n8656), .C1(n8634), .C2(n8654), .ZN(n8762) );
  NOR2_X1 U10065 ( .A1(n8762), .A2(n7135), .ZN(n8636) );
  AOI211_X1 U10066 ( .C1(n8760), .C2(n8669), .A(n8637), .B(n8636), .ZN(n8638)
         );
  OAI21_X1 U10067 ( .B1(n8711), .B2(n8763), .A(n8638), .ZN(P2_U3274) );
  XOR2_X1 U10068 ( .A(n8646), .B(n8639), .Z(n8768) );
  INV_X1 U10069 ( .A(n8668), .ZN(n8641) );
  AOI21_X1 U10070 ( .B1(n8764), .B2(n8641), .A(n8640), .ZN(n8765) );
  AOI22_X1 U10071 ( .A1(n7135), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8642), .B2(
        n8697), .ZN(n8643) );
  OAI21_X1 U10072 ( .B1(n8644), .B2(n8700), .A(n8643), .ZN(n8651) );
  OAI21_X1 U10073 ( .B1(n4328), .B2(n8646), .A(n8645), .ZN(n8649) );
  AOI222_X1 U10074 ( .A1(n8659), .A2(n8649), .B1(n8648), .B2(n8654), .C1(n8647), .C2(n8656), .ZN(n8767) );
  NOR2_X1 U10075 ( .A1(n8767), .A2(n7135), .ZN(n8650) );
  AOI211_X1 U10076 ( .C1(n8765), .C2(n8669), .A(n8651), .B(n8650), .ZN(n8652)
         );
  OAI21_X1 U10077 ( .B1(n8768), .B2(n8711), .A(n8652), .ZN(P2_U3275) );
  XNOR2_X1 U10078 ( .A(n8653), .B(n8660), .ZN(n8658) );
  AOI222_X1 U10079 ( .A1(n8659), .A2(n8658), .B1(n8657), .B2(n8656), .C1(n8655), .C2(n8654), .ZN(n8774) );
  NAND2_X1 U10080 ( .A1(n8661), .A2(n8660), .ZN(n8769) );
  NAND3_X1 U10081 ( .A1(n8770), .A2(n8769), .A3(n8662), .ZN(n8672) );
  INV_X1 U10082 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8664) );
  OAI22_X1 U10083 ( .A1(n8688), .A2(n8664), .B1(n8663), .B2(n8679), .ZN(n8665)
         );
  AOI21_X1 U10084 ( .B1(n8771), .B2(n8666), .A(n8665), .ZN(n8671) );
  AND2_X1 U10085 ( .A1(n8676), .A2(n8771), .ZN(n8667) );
  NOR2_X1 U10086 ( .A1(n8668), .A2(n8667), .ZN(n8772) );
  NAND2_X1 U10087 ( .A1(n8772), .A2(n8669), .ZN(n8670) );
  AND3_X1 U10088 ( .A1(n8672), .A2(n8671), .A3(n8670), .ZN(n8673) );
  OAI21_X1 U10089 ( .B1(n7135), .B2(n8774), .A(n8673), .ZN(P2_U3276) );
  XNOR2_X1 U10090 ( .A(n8675), .B(n8674), .ZN(n8780) );
  INV_X1 U10091 ( .A(n8676), .ZN(n8677) );
  AOI211_X1 U10092 ( .C1(n8778), .C2(n8695), .A(n9936), .B(n8677), .ZN(n8777)
         );
  INV_X1 U10093 ( .A(n8778), .ZN(n8678) );
  NOR2_X1 U10094 ( .A1(n8678), .A2(n8700), .ZN(n8683) );
  OAI22_X1 U10095 ( .A1(n8688), .A2(n8681), .B1(n8680), .B2(n8679), .ZN(n8682)
         );
  AOI211_X1 U10096 ( .C1(n8777), .C2(n8703), .A(n8683), .B(n8682), .ZN(n8690)
         );
  XNOR2_X1 U10097 ( .A(n8685), .B(n8684), .ZN(n8687) );
  OAI21_X1 U10098 ( .B1(n8687), .B2(n8707), .A(n8686), .ZN(n8776) );
  NAND2_X1 U10099 ( .A1(n8776), .A2(n8688), .ZN(n8689) );
  OAI211_X1 U10100 ( .C1(n8780), .C2(n8711), .A(n8690), .B(n8689), .ZN(
        P2_U3277) );
  OAI21_X1 U10101 ( .B1(n8692), .B2(n8704), .A(n8691), .ZN(n8693) );
  INV_X1 U10102 ( .A(n8693), .ZN(n8786) );
  INV_X1 U10103 ( .A(n8694), .ZN(n8696) );
  AOI211_X1 U10104 ( .C1(n8783), .C2(n8696), .A(n9936), .B(n4419), .ZN(n8782)
         );
  AOI22_X1 U10105 ( .A1(n7135), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8698), .B2(
        n8697), .ZN(n8699) );
  OAI21_X1 U10106 ( .B1(n8701), .B2(n8700), .A(n8699), .ZN(n8702) );
  AOI21_X1 U10107 ( .B1(n8782), .B2(n8703), .A(n8702), .ZN(n8710) );
  XOR2_X1 U10108 ( .A(n8705), .B(n8704), .Z(n8708) );
  OAI21_X1 U10109 ( .B1(n8708), .B2(n8707), .A(n8706), .ZN(n8781) );
  NAND2_X1 U10110 ( .A1(n8781), .A2(n8688), .ZN(n8709) );
  OAI211_X1 U10111 ( .C1(n8786), .C2(n8711), .A(n8710), .B(n8709), .ZN(
        P2_U3278) );
  NAND2_X1 U10112 ( .A1(n8712), .A2(n9475), .ZN(n8713) );
  OAI211_X1 U10113 ( .C1(n8714), .C2(n9936), .A(n8713), .B(n8717), .ZN(n8802)
         );
  MUX2_X1 U10114 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8802), .S(n9954), .Z(
        P2_U3551) );
  NAND3_X1 U10115 ( .A1(n8716), .A2(n9912), .A3(n8715), .ZN(n8718) );
  OAI211_X1 U10116 ( .C1(n8719), .C2(n9934), .A(n8718), .B(n8717), .ZN(n8803)
         );
  MUX2_X1 U10117 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8803), .S(n9954), .Z(
        P2_U3550) );
  AOI22_X1 U10118 ( .A1(n8726), .A2(n9912), .B1(n9475), .B2(n8725), .ZN(n8727)
         );
  OAI211_X1 U10119 ( .C1(n8729), .C2(n8785), .A(n8728), .B(n8727), .ZN(n8804)
         );
  MUX2_X1 U10120 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8804), .S(n9954), .Z(
        P2_U3548) );
  AOI211_X1 U10121 ( .C1(n9475), .C2(n8732), .A(n8731), .B(n8730), .ZN(n8733)
         );
  OAI21_X1 U10122 ( .B1(n8734), .B2(n8785), .A(n8733), .ZN(n8805) );
  MUX2_X1 U10123 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8805), .S(n9954), .Z(
        P2_U3547) );
  AOI211_X1 U10124 ( .C1(n9475), .C2(n8737), .A(n8736), .B(n8735), .ZN(n8738)
         );
  OAI21_X1 U10125 ( .B1(n8785), .B2(n8739), .A(n8738), .ZN(n8806) );
  MUX2_X1 U10126 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8806), .S(n9954), .Z(
        P2_U3546) );
  AOI211_X1 U10127 ( .C1(n9475), .C2(n8742), .A(n8741), .B(n8740), .ZN(n8744)
         );
  OAI211_X1 U10128 ( .C1(n8745), .C2(n8785), .A(n8744), .B(n8743), .ZN(n8807)
         );
  MUX2_X1 U10129 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8807), .S(n9954), .Z(
        P2_U3545) );
  INV_X1 U10130 ( .A(n8746), .ZN(n8751) );
  AOI22_X1 U10131 ( .A1(n8748), .A2(n9912), .B1(n9475), .B2(n8747), .ZN(n8749)
         );
  OAI211_X1 U10132 ( .C1(n8751), .C2(n8785), .A(n8750), .B(n8749), .ZN(n8808)
         );
  MUX2_X1 U10133 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8808), .S(n9954), .Z(
        P2_U3544) );
  OR2_X1 U10134 ( .A1(n8752), .A2(n8785), .ZN(n8758) );
  OAI22_X1 U10135 ( .A1(n8754), .A2(n9936), .B1(n8753), .B2(n9934), .ZN(n8755)
         );
  NOR2_X1 U10136 ( .A1(n8756), .A2(n8755), .ZN(n8757) );
  NAND2_X1 U10137 ( .A1(n8758), .A2(n8757), .ZN(n8809) );
  MUX2_X1 U10138 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8809), .S(n9954), .Z(
        P2_U3543) );
  AOI22_X1 U10139 ( .A1(n8760), .A2(n9912), .B1(n9475), .B2(n8759), .ZN(n8761)
         );
  OAI211_X1 U10140 ( .C1(n8763), .C2(n8785), .A(n8762), .B(n8761), .ZN(n8810)
         );
  MUX2_X1 U10141 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8810), .S(n9954), .Z(
        P2_U3542) );
  AOI22_X1 U10142 ( .A1(n8765), .A2(n9912), .B1(n9475), .B2(n8764), .ZN(n8766)
         );
  OAI211_X1 U10143 ( .C1(n8768), .C2(n8785), .A(n8767), .B(n8766), .ZN(n8811)
         );
  MUX2_X1 U10144 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8811), .S(n9954), .Z(
        P2_U3541) );
  NAND3_X1 U10145 ( .A1(n8770), .A2(n9931), .A3(n8769), .ZN(n8775) );
  AOI22_X1 U10146 ( .A1(n8772), .A2(n9912), .B1(n9475), .B2(n8771), .ZN(n8773)
         );
  NAND3_X1 U10147 ( .A1(n8775), .A2(n8774), .A3(n8773), .ZN(n8812) );
  MUX2_X1 U10148 ( .A(n8812), .B(P2_REG1_REG_20__SCAN_IN), .S(n9952), .Z(
        P2_U3540) );
  AOI211_X1 U10149 ( .C1(n9475), .C2(n8778), .A(n8777), .B(n8776), .ZN(n8779)
         );
  OAI21_X1 U10150 ( .B1(n8780), .B2(n8785), .A(n8779), .ZN(n8813) );
  MUX2_X1 U10151 ( .A(n8813), .B(P2_REG1_REG_19__SCAN_IN), .S(n9952), .Z(
        P2_U3539) );
  AOI211_X1 U10152 ( .C1(n9475), .C2(n8783), .A(n8782), .B(n8781), .ZN(n8784)
         );
  OAI21_X1 U10153 ( .B1(n8786), .B2(n8785), .A(n8784), .ZN(n8957) );
  MUX2_X1 U10154 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8957), .S(n9954), .Z(
        P2_U3538) );
  NAND2_X1 U10155 ( .A1(n8787), .A2(n9475), .ZN(n8788) );
  NAND3_X1 U10156 ( .A1(n8790), .A2(n8789), .A3(n8788), .ZN(n8791) );
  AOI21_X1 U10157 ( .B1(n8792), .B2(n9931), .A(n8791), .ZN(n8959) );
  MUX2_X1 U10158 ( .A(n8959), .B(n8793), .S(n9952), .Z(n8794) );
  INV_X1 U10159 ( .A(n8794), .ZN(P2_U3537) );
  INV_X1 U10160 ( .A(n8795), .ZN(n8796) );
  OAI22_X1 U10161 ( .A1(n8797), .A2(n9936), .B1(n8796), .B2(n9934), .ZN(n8798)
         );
  AOI21_X1 U10162 ( .B1(n8799), .B2(n9941), .A(n8798), .ZN(n8801) );
  NAND2_X1 U10163 ( .A1(n8801), .A2(n8800), .ZN(n8961) );
  MUX2_X1 U10164 ( .A(n8961), .B(P2_REG1_REG_16__SCAN_IN), .S(n9952), .Z(
        P2_U3536) );
  MUX2_X1 U10165 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8802), .S(n9944), .Z(
        P2_U3519) );
  MUX2_X1 U10166 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8803), .S(n9944), .Z(
        P2_U3518) );
  MUX2_X1 U10167 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8804), .S(n9944), .Z(
        P2_U3516) );
  MUX2_X1 U10168 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8805), .S(n9944), .Z(
        P2_U3515) );
  MUX2_X1 U10169 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8806), .S(n9944), .Z(
        P2_U3514) );
  MUX2_X1 U10170 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8807), .S(n9944), .Z(
        P2_U3513) );
  MUX2_X1 U10171 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8808), .S(n9944), .Z(
        P2_U3512) );
  MUX2_X1 U10172 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8809), .S(n9944), .Z(
        P2_U3511) );
  MUX2_X1 U10173 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8810), .S(n9944), .Z(
        P2_U3510) );
  MUX2_X1 U10174 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8811), .S(n9944), .Z(
        P2_U3509) );
  MUX2_X1 U10175 ( .A(n8812), .B(P2_REG0_REG_20__SCAN_IN), .S(n9942), .Z(
        P2_U3508) );
  MUX2_X1 U10176 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8813), .S(n9944), .Z(n8956) );
  INV_X1 U10177 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9752) );
  AOI22_X1 U10178 ( .A1(n8815), .A2(keyinput6), .B1(keyinput5), .B2(n9752), 
        .ZN(n8814) );
  OAI221_X1 U10179 ( .B1(n8815), .B2(keyinput6), .C1(n9752), .C2(keyinput5), 
        .A(n8814), .ZN(n8824) );
  AOI22_X1 U10180 ( .A1(n8817), .A2(keyinput53), .B1(n5575), .B2(keyinput52), 
        .ZN(n8816) );
  OAI221_X1 U10181 ( .B1(n8817), .B2(keyinput53), .C1(n5575), .C2(keyinput52), 
        .A(n8816), .ZN(n8823) );
  AOI22_X1 U10182 ( .A1(n8916), .A2(keyinput40), .B1(keyinput38), .B2(n5604), 
        .ZN(n8818) );
  OAI221_X1 U10183 ( .B1(n8916), .B2(keyinput40), .C1(n5604), .C2(keyinput38), 
        .A(n8818), .ZN(n8822) );
  INV_X1 U10184 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9540) );
  AOI22_X1 U10185 ( .A1(n9540), .A2(keyinput26), .B1(keyinput49), .B2(n8820), 
        .ZN(n8819) );
  OAI221_X1 U10186 ( .B1(n9540), .B2(keyinput26), .C1(n8820), .C2(keyinput49), 
        .A(n8819), .ZN(n8821) );
  NOR4_X1 U10187 ( .A1(n8824), .A2(n8823), .A3(n8822), .A4(n8821), .ZN(n8875)
         );
  INV_X1 U10188 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8826) );
  AOI22_X1 U10189 ( .A1(n5337), .A2(keyinput39), .B1(keyinput7), .B2(n8826), 
        .ZN(n8825) );
  OAI221_X1 U10190 ( .B1(n5337), .B2(keyinput39), .C1(n8826), .C2(keyinput7), 
        .A(n8825), .ZN(n8834) );
  INV_X1 U10191 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n8828) );
  AOI22_X1 U10192 ( .A1(n8828), .A2(keyinput3), .B1(n9867), .B2(keyinput19), 
        .ZN(n8827) );
  OAI221_X1 U10193 ( .B1(n8828), .B2(keyinput3), .C1(n9867), .C2(keyinput19), 
        .A(n8827), .ZN(n8833) );
  INV_X1 U10194 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8830) );
  AOI22_X1 U10195 ( .A1(n8831), .A2(keyinput24), .B1(keyinput61), .B2(n8830), 
        .ZN(n8829) );
  OAI221_X1 U10196 ( .B1(n8831), .B2(keyinput24), .C1(n8830), .C2(keyinput61), 
        .A(n8829), .ZN(n8832) );
  NOR3_X1 U10197 ( .A1(n8834), .A2(n8833), .A3(n8832), .ZN(n8862) );
  INV_X1 U10198 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n9742) );
  AOI22_X1 U10199 ( .A1(n8918), .A2(keyinput1), .B1(n9742), .B2(keyinput10), 
        .ZN(n8835) );
  OAI221_X1 U10200 ( .B1(n8918), .B2(keyinput1), .C1(n9742), .C2(keyinput10), 
        .A(n8835), .ZN(n8838) );
  AOI22_X1 U10201 ( .A1(n9534), .A2(keyinput29), .B1(n8943), .B2(keyinput8), 
        .ZN(n8836) );
  OAI221_X1 U10202 ( .B1(n9534), .B2(keyinput29), .C1(n8943), .C2(keyinput8), 
        .A(n8836), .ZN(n8837) );
  NOR2_X1 U10203 ( .A1(n8838), .A2(n8837), .ZN(n8861) );
  AOI22_X1 U10204 ( .A1(n8840), .A2(keyinput31), .B1(keyinput20), .B2(n4462), 
        .ZN(n8839) );
  OAI221_X1 U10205 ( .B1(n8840), .B2(keyinput31), .C1(n4462), .C2(keyinput20), 
        .A(n8839), .ZN(n8844) );
  INV_X1 U10206 ( .A(SI_18_), .ZN(n8842) );
  INV_X1 U10207 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n9887) );
  AOI22_X1 U10208 ( .A1(n8842), .A2(keyinput57), .B1(keyinput41), .B2(n9887), 
        .ZN(n8841) );
  OAI221_X1 U10209 ( .B1(n8842), .B2(keyinput57), .C1(n9887), .C2(keyinput41), 
        .A(n8841), .ZN(n8843) );
  NOR2_X1 U10210 ( .A1(n8844), .A2(n8843), .ZN(n8860) );
  AOI22_X1 U10211 ( .A1(n9307), .A2(keyinput56), .B1(keyinput17), .B2(n9528), 
        .ZN(n8845) );
  OAI221_X1 U10212 ( .B1(n9307), .B2(keyinput56), .C1(n9528), .C2(keyinput17), 
        .A(n8845), .ZN(n8858) );
  XNOR2_X1 U10213 ( .A(P2_IR_REG_26__SCAN_IN), .B(keyinput63), .ZN(n8849) );
  XNOR2_X1 U10214 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(keyinput28), .ZN(n8848) );
  XNOR2_X1 U10215 ( .A(P2_REG0_REG_20__SCAN_IN), .B(keyinput22), .ZN(n8847) );
  XNOR2_X1 U10216 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput35), .ZN(n8846) );
  AND4_X1 U10217 ( .A1(n8849), .A2(n8848), .A3(n8847), .A4(n8846), .ZN(n8856)
         );
  XNOR2_X1 U10218 ( .A(keyinput23), .B(P1_REG2_REG_27__SCAN_IN), .ZN(n8855) );
  XNOR2_X1 U10219 ( .A(keyinput58), .B(n4847), .ZN(n8852) );
  XNOR2_X1 U10220 ( .A(keyinput51), .B(n8850), .ZN(n8851) );
  NOR2_X1 U10221 ( .A1(n8852), .A2(n8851), .ZN(n8854) );
  XNOR2_X1 U10222 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput47), .ZN(n8853) );
  NAND4_X1 U10223 ( .A1(n8856), .A2(n8855), .A3(n8854), .A4(n8853), .ZN(n8857)
         );
  NOR2_X1 U10224 ( .A1(n8858), .A2(n8857), .ZN(n8859) );
  AND4_X1 U10225 ( .A1(n8862), .A2(n8861), .A3(n8860), .A4(n8859), .ZN(n8874)
         );
  INV_X1 U10226 ( .A(SI_3_), .ZN(n8936) );
  AOI22_X1 U10227 ( .A1(n8936), .A2(keyinput59), .B1(n8934), .B2(keyinput14), 
        .ZN(n8863) );
  OAI221_X1 U10228 ( .B1(n8936), .B2(keyinput59), .C1(n8934), .C2(keyinput14), 
        .A(n8863), .ZN(n8872) );
  AOI22_X1 U10229 ( .A1(n8935), .A2(keyinput0), .B1(keyinput37), .B2(n8865), 
        .ZN(n8864) );
  OAI221_X1 U10230 ( .B1(n8935), .B2(keyinput0), .C1(n8865), .C2(keyinput37), 
        .A(n8864), .ZN(n8871) );
  INV_X1 U10231 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n9888) );
  INV_X1 U10232 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8867) );
  AOI22_X1 U10233 ( .A1(n9888), .A2(keyinput16), .B1(keyinput55), .B2(n8867), 
        .ZN(n8866) );
  OAI221_X1 U10234 ( .B1(n9888), .B2(keyinput16), .C1(n8867), .C2(keyinput55), 
        .A(n8866), .ZN(n8870) );
  AOI22_X1 U10235 ( .A1(n8944), .A2(keyinput15), .B1(n8933), .B2(keyinput32), 
        .ZN(n8868) );
  OAI221_X1 U10236 ( .B1(n8944), .B2(keyinput15), .C1(n8933), .C2(keyinput32), 
        .A(n8868), .ZN(n8869) );
  NOR4_X1 U10237 ( .A1(n8872), .A2(n8871), .A3(n8870), .A4(n8869), .ZN(n8873)
         );
  AND3_X1 U10238 ( .A1(n8875), .A2(n8874), .A3(n8873), .ZN(n8915) );
  INV_X1 U10239 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n9740) );
  INV_X1 U10240 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n8877) );
  AOI22_X1 U10241 ( .A1(n9740), .A2(keyinput34), .B1(keyinput12), .B2(n8877), 
        .ZN(n8876) );
  OAI221_X1 U10242 ( .B1(n9740), .B2(keyinput34), .C1(n8877), .C2(keyinput12), 
        .A(n8876), .ZN(n8886) );
  AOI22_X1 U10243 ( .A1(n8917), .A2(keyinput46), .B1(n6150), .B2(keyinput4), 
        .ZN(n8878) );
  OAI221_X1 U10244 ( .B1(n8917), .B2(keyinput46), .C1(n6150), .C2(keyinput4), 
        .A(n8878), .ZN(n8885) );
  INV_X1 U10245 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8937) );
  AOI22_X1 U10246 ( .A1(n8937), .A2(keyinput36), .B1(keyinput30), .B2(n9985), 
        .ZN(n8879) );
  OAI221_X1 U10247 ( .B1(n8937), .B2(keyinput36), .C1(n9985), .C2(keyinput30), 
        .A(n8879), .ZN(n8884) );
  INV_X1 U10248 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8882) );
  AOI22_X1 U10249 ( .A1(n8882), .A2(keyinput13), .B1(keyinput54), .B2(n8881), 
        .ZN(n8880) );
  OAI221_X1 U10250 ( .B1(n8882), .B2(keyinput13), .C1(n8881), .C2(keyinput54), 
        .A(n8880), .ZN(n8883) );
  NOR4_X1 U10251 ( .A1(n8886), .A2(n8885), .A3(n8884), .A4(n8883), .ZN(n8914)
         );
  AOI22_X1 U10252 ( .A1(n9820), .A2(keyinput45), .B1(n8888), .B2(keyinput42), 
        .ZN(n8887) );
  OAI221_X1 U10253 ( .B1(n9820), .B2(keyinput45), .C1(n8888), .C2(keyinput42), 
        .A(n8887), .ZN(n8899) );
  AOI22_X1 U10254 ( .A1(n8891), .A2(keyinput18), .B1(keyinput2), .B2(n8890), 
        .ZN(n8889) );
  OAI221_X1 U10255 ( .B1(n8891), .B2(keyinput18), .C1(n8890), .C2(keyinput2), 
        .A(n8889), .ZN(n8898) );
  INV_X1 U10256 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8893) );
  AOI22_X1 U10257 ( .A1(n8893), .A2(keyinput33), .B1(n6063), .B2(keyinput50), 
        .ZN(n8892) );
  OAI221_X1 U10258 ( .B1(n8893), .B2(keyinput33), .C1(n6063), .C2(keyinput50), 
        .A(n8892), .ZN(n8897) );
  INV_X1 U10259 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8895) );
  AOI22_X1 U10260 ( .A1(n8942), .A2(keyinput44), .B1(n8895), .B2(keyinput27), 
        .ZN(n8894) );
  OAI221_X1 U10261 ( .B1(n8942), .B2(keyinput44), .C1(n8895), .C2(keyinput27), 
        .A(n8894), .ZN(n8896) );
  NOR4_X1 U10262 ( .A1(n8899), .A2(n8898), .A3(n8897), .A4(n8896), .ZN(n8913)
         );
  INV_X1 U10263 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n9889) );
  AOI22_X1 U10264 ( .A1(n9889), .A2(keyinput9), .B1(n5877), .B2(keyinput11), 
        .ZN(n8900) );
  OAI221_X1 U10265 ( .B1(n9889), .B2(keyinput9), .C1(n5877), .C2(keyinput11), 
        .A(n8900), .ZN(n8911) );
  INV_X1 U10266 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8902) );
  INV_X1 U10267 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n9741) );
  AOI22_X1 U10268 ( .A1(n8902), .A2(keyinput43), .B1(n9741), .B2(keyinput60), 
        .ZN(n8901) );
  OAI221_X1 U10269 ( .B1(n8902), .B2(keyinput43), .C1(n9741), .C2(keyinput60), 
        .A(n8901), .ZN(n8910) );
  INV_X1 U10270 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8904) );
  AOI22_X1 U10271 ( .A1(n8948), .A2(keyinput25), .B1(keyinput21), .B2(n8904), 
        .ZN(n8903) );
  OAI221_X1 U10272 ( .B1(n8948), .B2(keyinput25), .C1(n8904), .C2(keyinput21), 
        .A(n8903), .ZN(n8909) );
  AOI22_X1 U10273 ( .A1(n8907), .A2(keyinput62), .B1(keyinput48), .B2(n8906), 
        .ZN(n8905) );
  OAI221_X1 U10274 ( .B1(n8907), .B2(keyinput62), .C1(n8906), .C2(keyinput48), 
        .A(n8905), .ZN(n8908) );
  NOR4_X1 U10275 ( .A1(n8911), .A2(n8910), .A3(n8909), .A4(n8908), .ZN(n8912)
         );
  NAND4_X1 U10276 ( .A1(n8915), .A2(n8914), .A3(n8913), .A4(n8912), .ZN(n8954)
         );
  OR4_X1 U10277 ( .A1(P1_REG0_REG_19__SCAN_IN), .A2(P1_REG2_REG_18__SCAN_IN), 
        .A3(P1_REG1_REG_13__SCAN_IN), .A4(n5337), .ZN(n8932) );
  NAND4_X1 U10278 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P2_REG2_REG_25__SCAN_IN), 
        .A3(P1_REG0_REG_30__SCAN_IN), .A4(n9740), .ZN(n8921) );
  NAND4_X1 U10279 ( .A1(n8917), .A2(n8916), .A3(P2_ADDR_REG_19__SCAN_IN), .A4(
        SI_15_), .ZN(n8920) );
  NAND4_X1 U10280 ( .A1(n8918), .A2(P2_IR_REG_26__SCAN_IN), .A3(
        P2_IR_REG_20__SCAN_IN), .A4(P1_REG0_REG_13__SCAN_IN), .ZN(n8919) );
  NOR3_X1 U10281 ( .A1(n8921), .A2(n8920), .A3(n8919), .ZN(n8930) );
  NOR3_X1 U10282 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_REG2_REG_24__SCAN_IN), 
        .A3(n9752), .ZN(n8929) );
  NOR3_X1 U10283 ( .A1(SI_18_), .A2(P1_DATAO_REG_16__SCAN_IN), .A3(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n8922) );
  AND2_X1 U10284 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(n8922), .ZN(n8923) );
  NAND4_X1 U10285 ( .A1(n8923), .A2(P2_ADDR_REG_6__SCAN_IN), .A3(n8881), .A4(
        P1_ADDR_REG_16__SCAN_IN), .ZN(n8926) );
  NAND4_X1 U10286 ( .A1(n9742), .A2(n9889), .A3(n8924), .A4(
        P2_IR_REG_0__SCAN_IN), .ZN(n8925) );
  NOR2_X1 U10287 ( .A1(n8926), .A2(n8925), .ZN(n8927) );
  NAND4_X1 U10288 ( .A1(n8930), .A2(n8929), .A3(n8928), .A4(n8927), .ZN(n8931)
         );
  NOR2_X1 U10289 ( .A1(n8932), .A2(n8931), .ZN(n8952) );
  NAND4_X1 U10290 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(n8935), .A3(n8934), .A4(
        n8933), .ZN(n8941) );
  NAND4_X1 U10291 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), 
        .A3(n8936), .A4(n4462), .ZN(n8940) );
  NAND4_X1 U10292 ( .A1(P2_REG0_REG_18__SCAN_IN), .A2(P2_REG3_REG_16__SCAN_IN), 
        .A3(P2_REG1_REG_18__SCAN_IN), .A4(n8937), .ZN(n8939) );
  NAND4_X1 U10293 ( .A1(P2_REG0_REG_20__SCAN_IN), .A2(P2_REG2_REG_11__SCAN_IN), 
        .A3(P2_REG0_REG_15__SCAN_IN), .A4(n9820), .ZN(n8938) );
  NOR4_X1 U10294 ( .A1(n8941), .A2(n8940), .A3(n8939), .A4(n8938), .ZN(n8951)
         );
  NAND3_X1 U10295 ( .A1(SI_27_), .A2(n9534), .A3(n8942), .ZN(n8947) );
  NAND4_X1 U10296 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_REG3_REG_25__SCAN_IN), 
        .A3(P1_REG3_REG_21__SCAN_IN), .A4(n8943), .ZN(n8946) );
  NAND4_X1 U10297 ( .A1(P1_REG2_REG_27__SCAN_IN), .A2(P1_DATAO_REG_30__SCAN_IN), .A3(P1_REG1_REG_30__SCAN_IN), .A4(n8944), .ZN(n8945) );
  NOR4_X1 U10298 ( .A1(P1_REG2_REG_25__SCAN_IN), .A2(n8947), .A3(n8946), .A4(
        n8945), .ZN(n8950) );
  NOR4_X1 U10299 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(SI_21_), .A3(n8948), 
        .A4(n5877), .ZN(n8949) );
  NAND4_X1 U10300 ( .A1(n8952), .A2(n8951), .A3(n8950), .A4(n8949), .ZN(n8953)
         );
  XNOR2_X1 U10301 ( .A(n8954), .B(n8953), .ZN(n8955) );
  XNOR2_X1 U10302 ( .A(n8956), .B(n8955), .ZN(P2_U3507) );
  MUX2_X1 U10303 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8957), .S(n9944), .Z(
        P2_U3505) );
  INV_X1 U10304 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8958) );
  MUX2_X1 U10305 ( .A(n8959), .B(n8958), .S(n9942), .Z(n8960) );
  INV_X1 U10306 ( .A(n8960), .ZN(P2_U3502) );
  MUX2_X1 U10307 ( .A(n8961), .B(P2_REG0_REG_16__SCAN_IN), .S(n9942), .Z(
        P2_U3499) );
  INV_X1 U10308 ( .A(n8962), .ZN(n8963) );
  MUX2_X1 U10309 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8963), .S(n9944), .Z(
        P2_U3496) );
  INV_X1 U10310 ( .A(n9448), .ZN(n8970) );
  NOR4_X1 U10311 ( .A1(n8965), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3152), .A4(
        n8964), .ZN(n8966) );
  AOI21_X1 U10312 ( .B1(n8967), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8966), .ZN(
        n8968) );
  OAI21_X1 U10313 ( .B1(n8970), .B2(n8969), .A(n8968), .ZN(P2_U3327) );
  OAI222_X1 U10314 ( .A1(n8975), .A2(n8974), .B1(n8973), .B2(P2_U3152), .C1(
        n8972), .C2(n8971), .ZN(P2_U3329) );
  MUX2_X1 U10315 ( .A(n8976), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10316 ( .A(n8978), .ZN(n8979) );
  NOR2_X1 U10317 ( .A1(n8977), .A2(n8979), .ZN(n8981) );
  XNOR2_X1 U10318 ( .A(n8981), .B(n8980), .ZN(n8986) );
  AOI22_X1 U10319 ( .A1(n9101), .A2(n9206), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8983) );
  NAND2_X1 U10320 ( .A1(n9231), .A2(n9099), .ZN(n8982) );
  OAI211_X1 U10321 ( .C1(n9258), .C2(n9104), .A(n8983), .B(n8982), .ZN(n8984)
         );
  AOI21_X1 U10322 ( .B1(n9370), .B2(n9107), .A(n8984), .ZN(n8985) );
  OAI21_X1 U10323 ( .B1(n8986), .B2(n9460), .A(n8985), .ZN(P1_U3214) );
  OAI21_X1 U10324 ( .B1(n8989), .B2(n8988), .A(n8987), .ZN(n8990) );
  NAND2_X1 U10325 ( .A1(n8990), .A2(n9086), .ZN(n8994) );
  NAND2_X1 U10326 ( .A1(n9113), .A2(n9101), .ZN(n8991) );
  NAND2_X1 U10327 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9140) );
  OAI211_X1 U10328 ( .C1(n9320), .C2(n9104), .A(n8991), .B(n9140), .ZN(n8992)
         );
  AOI21_X1 U10329 ( .B1(n9290), .B2(n9099), .A(n8992), .ZN(n8993) );
  OAI211_X1 U10330 ( .C1(n9293), .C2(n9095), .A(n8994), .B(n8993), .ZN(
        P1_U3217) );
  INV_X1 U10331 ( .A(n9013), .ZN(n9006) );
  NAND2_X1 U10332 ( .A1(n9345), .A2(n8995), .ZN(n8998) );
  NAND2_X1 U10333 ( .A1(n9111), .A2(n8996), .ZN(n8997) );
  NAND2_X1 U10334 ( .A1(n8998), .A2(n8997), .ZN(n9000) );
  XNOR2_X1 U10335 ( .A(n9000), .B(n8999), .ZN(n9004) );
  AOI22_X1 U10336 ( .A1(n9345), .A2(n9002), .B1(n9001), .B2(n9111), .ZN(n9003)
         );
  XNOR2_X1 U10337 ( .A(n9004), .B(n9003), .ZN(n9015) );
  NAND2_X1 U10338 ( .A1(n9006), .A2(n9005), .ZN(n9019) );
  NAND2_X1 U10339 ( .A1(n9099), .A2(n9158), .ZN(n9008) );
  AOI22_X1 U10340 ( .A1(n9101), .A2(n9164), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n9007) );
  OAI211_X1 U10341 ( .C1(n9009), .C2(n9104), .A(n9008), .B(n9007), .ZN(n9010)
         );
  AOI21_X1 U10342 ( .B1(n9345), .B2(n9107), .A(n9010), .ZN(n9018) );
  INV_X1 U10343 ( .A(n9014), .ZN(n9012) );
  INV_X1 U10344 ( .A(n9015), .ZN(n9011) );
  NAND4_X1 U10345 ( .A1(n9013), .A2(n9086), .A3(n9012), .A4(n9011), .ZN(n9017)
         );
  NAND3_X1 U10346 ( .A1(n9015), .A2(n9014), .A3(n9086), .ZN(n9016) );
  NAND4_X1 U10347 ( .A1(n9019), .A2(n9018), .A3(n9017), .A4(n9016), .ZN(
        P1_U3218) );
  NAND2_X1 U10348 ( .A1(n9021), .A2(n9020), .ZN(n9023) );
  XNOR2_X1 U10349 ( .A(n9023), .B(n9022), .ZN(n9024) );
  NAND2_X1 U10350 ( .A1(n9024), .A2(n9086), .ZN(n9030) );
  AOI22_X1 U10351 ( .A1(n9456), .A2(n9728), .B1(n9101), .B2(n9727), .ZN(n9029)
         );
  NAND2_X1 U10352 ( .A1(n9025), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n9028) );
  NAND2_X1 U10353 ( .A1(n9422), .A2(n9719), .ZN(n9747) );
  OR2_X1 U10354 ( .A1(n9026), .A2(n9747), .ZN(n9027) );
  NAND4_X1 U10355 ( .A1(n9030), .A2(n9029), .A3(n9028), .A4(n9027), .ZN(
        P1_U3220) );
  XOR2_X1 U10356 ( .A(n9032), .B(n9031), .Z(n9037) );
  AOI22_X1 U10357 ( .A1(n9112), .A2(n9101), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n9034) );
  NAND2_X1 U10358 ( .A1(n9456), .A2(n9113), .ZN(n9033) );
  OAI211_X1 U10359 ( .C1(n9468), .C2(n9261), .A(n9034), .B(n9033), .ZN(n9035)
         );
  AOI21_X1 U10360 ( .B1(n9382), .B2(n9107), .A(n9035), .ZN(n9036) );
  OAI21_X1 U10361 ( .B1(n9037), .B2(n9460), .A(n9036), .ZN(P1_U3221) );
  AOI22_X1 U10362 ( .A1(n9101), .A2(n9207), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9040) );
  NAND2_X1 U10363 ( .A1(n9456), .A2(n9206), .ZN(n9039) );
  OAI211_X1 U10364 ( .C1(n9468), .C2(n9041), .A(n9040), .B(n9039), .ZN(n9042)
         );
  AOI21_X1 U10365 ( .B1(n9360), .B2(n9107), .A(n9042), .ZN(n9043) );
  OAI21_X1 U10366 ( .B1(n9044), .B2(n9460), .A(n9043), .ZN(P1_U3223) );
  XOR2_X1 U10367 ( .A(n9046), .B(n9045), .Z(n9052) );
  NAND2_X1 U10368 ( .A1(n9099), .A2(n9323), .ZN(n9049) );
  NOR2_X1 U10369 ( .A1(n9047), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9660) );
  AOI21_X1 U10370 ( .B1(n9101), .B2(n9114), .A(n9660), .ZN(n9048) );
  OAI211_X1 U10371 ( .C1(n9319), .C2(n9104), .A(n9049), .B(n9048), .ZN(n9050)
         );
  AOI21_X1 U10372 ( .B1(n9405), .B2(n9107), .A(n9050), .ZN(n9051) );
  OAI21_X1 U10373 ( .B1(n9052), .B2(n9460), .A(n9051), .ZN(P1_U3226) );
  OAI21_X1 U10374 ( .B1(n9055), .B2(n9054), .A(n9053), .ZN(n9056) );
  NAND2_X1 U10375 ( .A1(n9056), .A2(n9086), .ZN(n9060) );
  AOI22_X1 U10376 ( .A1(n9101), .A2(n9221), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9057) );
  OAI21_X1 U10377 ( .B1(n9251), .B2(n9104), .A(n9057), .ZN(n9058) );
  AOI21_X1 U10378 ( .B1(n9215), .B2(n9099), .A(n9058), .ZN(n9059) );
  OAI211_X1 U10379 ( .C1(n9217), .C2(n9095), .A(n9060), .B(n9059), .ZN(
        P1_U3227) );
  INV_X1 U10380 ( .A(n9061), .ZN(n9066) );
  AOI21_X1 U10381 ( .B1(n9063), .B2(n9065), .A(n4354), .ZN(n9064) );
  AOI21_X1 U10382 ( .B1(n9066), .B2(n9065), .A(n9064), .ZN(n9071) );
  AOI22_X1 U10383 ( .A1(n9276), .A2(n9101), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9068) );
  NAND2_X1 U10384 ( .A1(n9456), .A2(n9300), .ZN(n9067) );
  OAI211_X1 U10385 ( .C1(n9468), .C2(n9271), .A(n9068), .B(n9067), .ZN(n9069)
         );
  AOI21_X1 U10386 ( .B1(n9385), .B2(n9107), .A(n9069), .ZN(n9070) );
  OAI21_X1 U10387 ( .B1(n9071), .B2(n9460), .A(n9070), .ZN(P1_U3231) );
  INV_X1 U10388 ( .A(n9072), .ZN(n9073) );
  NOR2_X1 U10389 ( .A1(n9074), .A2(n9073), .ZN(n9076) );
  XNOR2_X1 U10390 ( .A(n9076), .B(n9075), .ZN(n9081) );
  AOI22_X1 U10391 ( .A1(n9222), .A2(n9101), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n9078) );
  NAND2_X1 U10392 ( .A1(n9276), .A2(n9456), .ZN(n9077) );
  OAI211_X1 U10393 ( .C1(n9468), .C2(n9244), .A(n9078), .B(n9077), .ZN(n9079)
         );
  AOI21_X1 U10394 ( .B1(n9377), .B2(n9107), .A(n9079), .ZN(n9080) );
  OAI21_X1 U10395 ( .B1(n9081), .B2(n9460), .A(n9080), .ZN(P1_U3233) );
  INV_X1 U10396 ( .A(n9084), .ZN(n9082) );
  AOI21_X1 U10397 ( .B1(n9085), .B2(n9084), .A(n9083), .ZN(n9087) );
  OAI21_X1 U10398 ( .B1(n9088), .B2(n9087), .A(n9086), .ZN(n9094) );
  OAI21_X1 U10399 ( .B1(n9453), .B2(n9090), .A(n9089), .ZN(n9092) );
  NOR2_X1 U10400 ( .A1(n9468), .A2(n9306), .ZN(n9091) );
  AOI211_X1 U10401 ( .C1(n9456), .C2(n9301), .A(n9092), .B(n9091), .ZN(n9093)
         );
  OAI211_X1 U10402 ( .C1(n9305), .C2(n9095), .A(n9094), .B(n9093), .ZN(
        P1_U3236) );
  NOR2_X1 U10403 ( .A1(n9096), .A2(n4333), .ZN(n9097) );
  XNOR2_X1 U10404 ( .A(n9098), .B(n9097), .ZN(n9109) );
  NAND2_X1 U10405 ( .A1(n9099), .A2(n9187), .ZN(n9103) );
  AOI22_X1 U10406 ( .A1(n9101), .A2(n9191), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9102) );
  OAI211_X1 U10407 ( .C1(n9105), .C2(n9104), .A(n9103), .B(n9102), .ZN(n9106)
         );
  AOI21_X1 U10408 ( .B1(n9355), .B2(n9107), .A(n9106), .ZN(n9108) );
  OAI21_X1 U10409 ( .B1(n9109), .B2(n9460), .A(n9108), .ZN(P1_U3238) );
  MUX2_X1 U10410 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9110), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10411 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9164), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10412 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9111), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10413 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9191), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10414 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9207), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10415 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9221), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10416 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9206), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10417 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9222), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10418 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9112), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10419 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9276), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10420 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9113), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10421 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9300), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10422 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9114), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10423 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9301), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10424 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9115), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10425 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9116), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10426 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9117), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10427 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9118), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10428 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9119), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10429 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9455), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10430 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9120), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10431 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9121), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10432 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9122), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10433 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9123), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10434 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9676), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10435 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9124), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10436 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9675), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10437 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9125), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10438 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9727), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10439 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6715), .S(P1_U4006), .Z(
        P1_U3556) );
  OAI21_X1 U10440 ( .B1(n9130), .B2(n9307), .A(n9126), .ZN(n9127) );
  XOR2_X1 U10441 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9127), .Z(n9134) );
  INV_X1 U10442 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9131) );
  XOR2_X1 U10443 ( .A(n9132), .B(n9131), .Z(n9136) );
  NAND2_X1 U10444 ( .A1(n9136), .A2(n9663), .ZN(n9133) );
  OAI211_X1 U10445 ( .C1(n9134), .C2(n9553), .A(n9133), .B(n9658), .ZN(n9139)
         );
  INV_X1 U10446 ( .A(n9134), .ZN(n9135) );
  OAI22_X1 U10447 ( .A1(n9136), .A2(n9621), .B1(n9627), .B2(n9135), .ZN(n9138)
         );
  NAND2_X1 U10448 ( .A1(n9149), .A2(n4265), .ZN(n9141) );
  XNOR2_X1 U10449 ( .A(n9330), .B(n9141), .ZN(n9332) );
  NOR2_X1 U10450 ( .A1(n9143), .A2(n9142), .ZN(n9333) );
  INV_X1 U10451 ( .A(n9333), .ZN(n9144) );
  NOR2_X1 U10452 ( .A1(n9739), .A2(n9144), .ZN(n9151) );
  NOR2_X1 U10453 ( .A1(n9145), .A2(n9710), .ZN(n9146) );
  AOI211_X1 U10454 ( .C1(n9739), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9151), .B(
        n9146), .ZN(n9147) );
  OAI21_X1 U10455 ( .B1(n9332), .B2(n9153), .A(n9147), .ZN(P1_U3261) );
  XNOR2_X1 U10456 ( .A(n9149), .B(n4265), .ZN(n9336) );
  NOR2_X1 U10457 ( .A1(n9149), .A2(n9710), .ZN(n9150) );
  AOI211_X1 U10458 ( .C1(n9739), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9151), .B(
        n9150), .ZN(n9152) );
  OAI21_X1 U10459 ( .B1(n9336), .B2(n9153), .A(n9152), .ZN(P1_U3262) );
  OAI21_X1 U10460 ( .B1(n9156), .B2(n9155), .A(n9154), .ZN(n9349) );
  AOI21_X1 U10461 ( .B1(n9345), .B2(n9170), .A(n9157), .ZN(n9346) );
  AOI22_X1 U10462 ( .A1(n9739), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9158), .B2(
        n9718), .ZN(n9159) );
  OAI21_X1 U10463 ( .B1(n4553), .B2(n9710), .A(n9159), .ZN(n9167) );
  NOR2_X1 U10464 ( .A1(n9175), .A2(n9160), .ZN(n9163) );
  OAI21_X1 U10465 ( .B1(n9163), .B2(n9162), .A(n9161), .ZN(n9165) );
  AOI222_X1 U10466 ( .A1(n9704), .A2(n9165), .B1(n9191), .B2(n9729), .C1(n9164), .C2(n9726), .ZN(n9348) );
  NOR2_X1 U10467 ( .A1(n9348), .A2(n9739), .ZN(n9166) );
  AOI211_X1 U10468 ( .C1(n9696), .C2(n9346), .A(n9167), .B(n9166), .ZN(n9168)
         );
  OAI21_X1 U10469 ( .B1(n9329), .B2(n9349), .A(n9168), .ZN(P1_U3263) );
  XOR2_X1 U10470 ( .A(n9177), .B(n9169), .Z(n9354) );
  INV_X1 U10471 ( .A(n9186), .ZN(n9171) );
  AOI211_X1 U10472 ( .C1(n9351), .C2(n9171), .A(n9801), .B(n4555), .ZN(n9350)
         );
  AOI22_X1 U10473 ( .A1(n9739), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9172), .B2(
        n9718), .ZN(n9173) );
  OAI21_X1 U10474 ( .B1(n9174), .B2(n9710), .A(n9173), .ZN(n9183) );
  AOI211_X1 U10475 ( .C1(n9177), .C2(n9176), .A(n9733), .B(n9175), .ZN(n9181)
         );
  OAI22_X1 U10476 ( .A1(n9179), .A2(n9701), .B1(n9178), .B2(n9699), .ZN(n9180)
         );
  NOR2_X1 U10477 ( .A1(n9181), .A2(n9180), .ZN(n9353) );
  NOR2_X1 U10478 ( .A1(n9353), .A2(n9739), .ZN(n9182) );
  AOI211_X1 U10479 ( .C1(n9260), .C2(n9350), .A(n9183), .B(n9182), .ZN(n9184)
         );
  OAI21_X1 U10480 ( .B1(n9354), .B2(n9329), .A(n9184), .ZN(P1_U3264) );
  XOR2_X1 U10481 ( .A(n9190), .B(n9185), .Z(n9359) );
  AOI21_X1 U10482 ( .B1(n9355), .B2(n9197), .A(n9186), .ZN(n9356) );
  AOI22_X1 U10483 ( .A1(n9739), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9187), .B2(
        n9718), .ZN(n9188) );
  OAI21_X1 U10484 ( .B1(n4557), .B2(n9710), .A(n9188), .ZN(n9194) );
  XOR2_X1 U10485 ( .A(n9190), .B(n9189), .Z(n9192) );
  AOI222_X1 U10486 ( .A1(n9704), .A2(n9192), .B1(n9221), .B2(n9729), .C1(n9191), .C2(n9726), .ZN(n9358) );
  NOR2_X1 U10487 ( .A1(n9358), .A2(n9739), .ZN(n9193) );
  AOI211_X1 U10488 ( .C1(n9696), .C2(n9356), .A(n9194), .B(n9193), .ZN(n9195)
         );
  OAI21_X1 U10489 ( .B1(n9329), .B2(n9359), .A(n9195), .ZN(P1_U3265) );
  XOR2_X1 U10490 ( .A(n9205), .B(n9196), .Z(n9364) );
  INV_X1 U10491 ( .A(n9213), .ZN(n9199) );
  INV_X1 U10492 ( .A(n9197), .ZN(n9198) );
  AOI21_X1 U10493 ( .B1(n9360), .B2(n9199), .A(n9198), .ZN(n9361) );
  AOI22_X1 U10494 ( .A1(n9739), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9200), .B2(
        n9718), .ZN(n9201) );
  OAI21_X1 U10495 ( .B1(n9202), .B2(n9710), .A(n9201), .ZN(n9210) );
  NAND2_X1 U10496 ( .A1(n9218), .A2(n9203), .ZN(n9204) );
  XOR2_X1 U10497 ( .A(n9205), .B(n9204), .Z(n9208) );
  AOI222_X1 U10498 ( .A1(n9704), .A2(n9208), .B1(n9207), .B2(n9726), .C1(n9206), .C2(n9729), .ZN(n9363) );
  NOR2_X1 U10499 ( .A1(n9363), .A2(n9739), .ZN(n9209) );
  AOI211_X1 U10500 ( .C1(n9361), .C2(n9696), .A(n9210), .B(n9209), .ZN(n9211)
         );
  OAI21_X1 U10501 ( .B1(n9364), .B2(n9329), .A(n9211), .ZN(P1_U3266) );
  XNOR2_X1 U10502 ( .A(n9212), .B(n9219), .ZN(n9369) );
  INV_X1 U10503 ( .A(n9229), .ZN(n9214) );
  AOI211_X1 U10504 ( .C1(n9366), .C2(n9214), .A(n9801), .B(n9213), .ZN(n9365)
         );
  AOI22_X1 U10505 ( .A1(n9739), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9215), .B2(
        n9718), .ZN(n9216) );
  OAI21_X1 U10506 ( .B1(n9217), .B2(n9710), .A(n9216), .ZN(n9225) );
  OAI21_X1 U10507 ( .B1(n9220), .B2(n9219), .A(n9218), .ZN(n9223) );
  AOI222_X1 U10508 ( .A1(n9704), .A2(n9223), .B1(n9222), .B2(n9729), .C1(n9221), .C2(n9726), .ZN(n9368) );
  NOR2_X1 U10509 ( .A1(n9368), .A2(n9739), .ZN(n9224) );
  AOI211_X1 U10510 ( .C1(n9365), .C2(n9260), .A(n9225), .B(n9224), .ZN(n9226)
         );
  OAI21_X1 U10511 ( .B1(n9369), .B2(n9329), .A(n9226), .ZN(P1_U3267) );
  XNOR2_X1 U10512 ( .A(n9228), .B(n9227), .ZN(n9374) );
  INV_X1 U10513 ( .A(n9242), .ZN(n9230) );
  AOI21_X1 U10514 ( .B1(n9370), .B2(n9230), .A(n9229), .ZN(n9371) );
  AOI22_X1 U10515 ( .A1(n9739), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9231), .B2(
        n9718), .ZN(n9232) );
  OAI21_X1 U10516 ( .B1(n9233), .B2(n9710), .A(n9232), .ZN(n9240) );
  AOI211_X1 U10517 ( .C1(n9235), .C2(n9234), .A(n9733), .B(n4299), .ZN(n9238)
         );
  OAI22_X1 U10518 ( .A1(n9258), .A2(n9699), .B1(n9236), .B2(n9701), .ZN(n9237)
         );
  NOR2_X1 U10519 ( .A1(n9238), .A2(n9237), .ZN(n9373) );
  NOR2_X1 U10520 ( .A1(n9373), .A2(n9739), .ZN(n9239) );
  AOI211_X1 U10521 ( .C1(n9371), .C2(n9696), .A(n9240), .B(n9239), .ZN(n9241)
         );
  OAI21_X1 U10522 ( .B1(n9374), .B2(n9329), .A(n9241), .ZN(P1_U3268) );
  XNOR2_X1 U10523 ( .A(n4288), .B(n4278), .ZN(n9379) );
  AOI211_X1 U10524 ( .C1(n9377), .C2(n9259), .A(n9801), .B(n9242), .ZN(n9376)
         );
  NOR2_X1 U10525 ( .A1(n9243), .A2(n9710), .ZN(n9247) );
  OAI22_X1 U10526 ( .A1(n9737), .A2(n9245), .B1(n9244), .B2(n9709), .ZN(n9246)
         );
  AOI211_X1 U10527 ( .C1(n9376), .C2(n9260), .A(n9247), .B(n9246), .ZN(n9253)
         );
  XNOR2_X1 U10528 ( .A(n9248), .B(n4278), .ZN(n9249) );
  OAI222_X1 U10529 ( .A1(n9701), .A2(n9251), .B1(n9699), .B2(n9250), .C1(n9249), .C2(n9733), .ZN(n9375) );
  NAND2_X1 U10530 ( .A1(n9375), .A2(n9737), .ZN(n9252) );
  OAI211_X1 U10531 ( .C1(n9379), .C2(n9329), .A(n9253), .B(n9252), .ZN(
        P1_U3269) );
  XNOR2_X1 U10532 ( .A(n9254), .B(n9255), .ZN(n9384) );
  XNOR2_X1 U10533 ( .A(n9256), .B(n9255), .ZN(n9257) );
  OAI222_X1 U10534 ( .A1(n9699), .A2(n9286), .B1(n9701), .B2(n9258), .C1(n9257), .C2(n9733), .ZN(n9380) );
  INV_X1 U10535 ( .A(n9382), .ZN(n9265) );
  AOI211_X1 U10536 ( .C1(n9382), .C2(n9269), .A(n9801), .B(n4568), .ZN(n9381)
         );
  NAND2_X1 U10537 ( .A1(n9381), .A2(n9260), .ZN(n9264) );
  INV_X1 U10538 ( .A(n9261), .ZN(n9262) );
  AOI22_X1 U10539 ( .A1(n9739), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9262), .B2(
        n9718), .ZN(n9263) );
  OAI211_X1 U10540 ( .C1(n9265), .C2(n9710), .A(n9264), .B(n9263), .ZN(n9266)
         );
  AOI21_X1 U10541 ( .B1(n9380), .B2(n9737), .A(n9266), .ZN(n9267) );
  OAI21_X1 U10542 ( .B1(n9384), .B2(n9329), .A(n9267), .ZN(P1_U3270) );
  XOR2_X1 U10543 ( .A(n9275), .B(n9268), .Z(n9389) );
  INV_X1 U10544 ( .A(n9269), .ZN(n9270) );
  AOI21_X1 U10545 ( .B1(n9385), .B2(n9287), .A(n9270), .ZN(n9386) );
  INV_X1 U10546 ( .A(n9271), .ZN(n9272) );
  AOI22_X1 U10547 ( .A1(n9739), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9272), .B2(
        n9718), .ZN(n9273) );
  OAI21_X1 U10548 ( .B1(n9274), .B2(n9710), .A(n9273), .ZN(n9279) );
  XOR2_X1 U10549 ( .A(n9275), .B(n4286), .Z(n9277) );
  AOI222_X1 U10550 ( .A1(n9704), .A2(n9277), .B1(n9300), .B2(n9729), .C1(n9276), .C2(n9726), .ZN(n9388) );
  NOR2_X1 U10551 ( .A1(n9388), .A2(n9739), .ZN(n9278) );
  AOI211_X1 U10552 ( .C1(n9386), .C2(n9696), .A(n9279), .B(n9278), .ZN(n9280)
         );
  OAI21_X1 U10553 ( .B1(n9329), .B2(n9389), .A(n9280), .ZN(P1_U3271) );
  XOR2_X1 U10554 ( .A(n9283), .B(n9281), .Z(n9395) );
  AOI21_X1 U10555 ( .B1(n9284), .B2(n9283), .A(n9282), .ZN(n9285) );
  OAI222_X1 U10556 ( .A1(n9699), .A2(n9320), .B1(n9701), .B2(n9286), .C1(n9733), .C2(n9285), .ZN(n9390) );
  INV_X1 U10557 ( .A(n9303), .ZN(n9289) );
  INV_X1 U10558 ( .A(n9287), .ZN(n9288) );
  AOI21_X1 U10559 ( .B1(n9391), .B2(n9289), .A(n9288), .ZN(n9392) );
  NAND2_X1 U10560 ( .A1(n9392), .A2(n9696), .ZN(n9292) );
  AOI22_X1 U10561 ( .A1(n9739), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9290), .B2(
        n9718), .ZN(n9291) );
  OAI211_X1 U10562 ( .C1(n9293), .C2(n9710), .A(n9292), .B(n9291), .ZN(n9294)
         );
  AOI21_X1 U10563 ( .B1(n9390), .B2(n9737), .A(n9294), .ZN(n9295) );
  OAI21_X1 U10564 ( .B1(n9395), .B2(n9329), .A(n9295), .ZN(P1_U3272) );
  NAND2_X1 U10565 ( .A1(n9297), .A2(n9296), .ZN(n9299) );
  XNOR2_X1 U10566 ( .A(n9299), .B(n9298), .ZN(n9302) );
  AOI222_X1 U10567 ( .A1(n9704), .A2(n9302), .B1(n9301), .B2(n9729), .C1(n9300), .C2(n9726), .ZN(n9400) );
  INV_X1 U10568 ( .A(n9321), .ZN(n9304) );
  AOI21_X1 U10569 ( .B1(n9397), .B2(n9304), .A(n9303), .ZN(n9398) );
  NOR2_X1 U10570 ( .A1(n9305), .A2(n9710), .ZN(n9309) );
  OAI22_X1 U10571 ( .A1(n9737), .A2(n9307), .B1(n9306), .B2(n9709), .ZN(n9308)
         );
  AOI211_X1 U10572 ( .C1(n9398), .C2(n9696), .A(n9309), .B(n9308), .ZN(n9314)
         );
  NAND2_X1 U10573 ( .A1(n9311), .A2(n9310), .ZN(n9396) );
  NAND3_X1 U10574 ( .A1(n4684), .A2(n9312), .A3(n9396), .ZN(n9313) );
  OAI211_X1 U10575 ( .C1(n9400), .C2(n9739), .A(n9314), .B(n9313), .ZN(
        P1_U3273) );
  XNOR2_X1 U10576 ( .A(n9315), .B(n9316), .ZN(n9407) );
  XNOR2_X1 U10577 ( .A(n9317), .B(n9316), .ZN(n9318) );
  OAI222_X1 U10578 ( .A1(n9701), .A2(n9320), .B1(n9699), .B2(n9319), .C1(n9318), .C2(n9733), .ZN(n9403) );
  AOI211_X1 U10579 ( .C1(n9405), .C2(n9322), .A(n9801), .B(n9321), .ZN(n9404)
         );
  INV_X1 U10580 ( .A(n9404), .ZN(n9325) );
  INV_X1 U10581 ( .A(n9323), .ZN(n9324) );
  OAI22_X1 U10582 ( .A1(n9325), .A2(n9721), .B1(n9709), .B2(n9324), .ZN(n9326)
         );
  OAI21_X1 U10583 ( .B1(n9403), .B2(n9326), .A(n9737), .ZN(n9328) );
  AOI22_X1 U10584 ( .A1(n9405), .A2(n9498), .B1(n9739), .B2(
        P1_REG2_REG_17__SCAN_IN), .ZN(n9327) );
  OAI211_X1 U10585 ( .C1(n9407), .C2(n9329), .A(n9328), .B(n9327), .ZN(
        P1_U3274) );
  AOI21_X1 U10586 ( .B1(n9330), .B2(n9422), .A(n9333), .ZN(n9331) );
  OAI21_X1 U10587 ( .B1(n9332), .B2(n9801), .A(n9331), .ZN(n9426) );
  MUX2_X1 U10588 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9426), .S(n9826), .Z(
        P1_U3554) );
  AOI21_X1 U10589 ( .B1(n9334), .B2(n9422), .A(n9333), .ZN(n9335) );
  OAI21_X1 U10590 ( .B1(n9336), .B2(n9801), .A(n9335), .ZN(n9427) );
  MUX2_X1 U10591 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9427), .S(n9826), .Z(
        P1_U3553) );
  INV_X1 U10592 ( .A(n9338), .ZN(n9341) );
  INV_X1 U10593 ( .A(n9339), .ZN(n9340) );
  OAI211_X1 U10594 ( .C1(n9799), .C2(n8038), .A(n9341), .B(n9340), .ZN(n9342)
         );
  INV_X1 U10595 ( .A(n9342), .ZN(n9343) );
  AOI22_X1 U10596 ( .A1(n9346), .A2(n9717), .B1(n9422), .B2(n9345), .ZN(n9347)
         );
  OAI211_X1 U10597 ( .C1(n9349), .C2(n9425), .A(n9348), .B(n9347), .ZN(n9428)
         );
  MUX2_X1 U10598 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9428), .S(n9826), .Z(
        P1_U3551) );
  AOI21_X1 U10599 ( .B1(n9422), .B2(n9351), .A(n9350), .ZN(n9352) );
  OAI211_X1 U10600 ( .C1(n9354), .C2(n9425), .A(n9353), .B(n9352), .ZN(n9429)
         );
  MUX2_X1 U10601 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9429), .S(n9826), .Z(
        P1_U3550) );
  AOI22_X1 U10602 ( .A1(n9356), .A2(n9717), .B1(n9422), .B2(n9355), .ZN(n9357)
         );
  OAI211_X1 U10603 ( .C1(n9359), .C2(n9425), .A(n9358), .B(n9357), .ZN(n9430)
         );
  MUX2_X1 U10604 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9430), .S(n9826), .Z(
        P1_U3549) );
  AOI22_X1 U10605 ( .A1(n9361), .A2(n9717), .B1(n9422), .B2(n9360), .ZN(n9362)
         );
  OAI211_X1 U10606 ( .C1(n9364), .C2(n9425), .A(n9363), .B(n9362), .ZN(n9431)
         );
  MUX2_X1 U10607 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9431), .S(n9826), .Z(
        P1_U3548) );
  AOI21_X1 U10608 ( .B1(n9422), .B2(n9366), .A(n9365), .ZN(n9367) );
  OAI211_X1 U10609 ( .C1(n9369), .C2(n9425), .A(n9368), .B(n9367), .ZN(n9432)
         );
  MUX2_X1 U10610 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9432), .S(n9826), .Z(
        P1_U3547) );
  AOI22_X1 U10611 ( .A1(n9371), .A2(n9717), .B1(n9422), .B2(n9370), .ZN(n9372)
         );
  OAI211_X1 U10612 ( .C1(n9374), .C2(n9425), .A(n9373), .B(n9372), .ZN(n9433)
         );
  MUX2_X1 U10613 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9433), .S(n9826), .Z(
        P1_U3546) );
  AOI211_X1 U10614 ( .C1(n9422), .C2(n9377), .A(n9376), .B(n9375), .ZN(n9378)
         );
  OAI21_X1 U10615 ( .B1(n9425), .B2(n9379), .A(n9378), .ZN(n9434) );
  MUX2_X1 U10616 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9434), .S(n9826), .Z(
        P1_U3545) );
  AOI211_X1 U10617 ( .C1(n9422), .C2(n9382), .A(n9381), .B(n9380), .ZN(n9383)
         );
  OAI21_X1 U10618 ( .B1(n9425), .B2(n9384), .A(n9383), .ZN(n9435) );
  MUX2_X1 U10619 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9435), .S(n9826), .Z(
        P1_U3544) );
  AOI22_X1 U10620 ( .A1(n9386), .A2(n9717), .B1(n9422), .B2(n9385), .ZN(n9387)
         );
  OAI211_X1 U10621 ( .C1(n9389), .C2(n9425), .A(n9388), .B(n9387), .ZN(n9436)
         );
  MUX2_X1 U10622 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9436), .S(n9826), .Z(
        P1_U3543) );
  INV_X1 U10623 ( .A(n9390), .ZN(n9394) );
  AOI22_X1 U10624 ( .A1(n9392), .A2(n9717), .B1(n9422), .B2(n9391), .ZN(n9393)
         );
  OAI211_X1 U10625 ( .C1(n9395), .C2(n9425), .A(n9394), .B(n9393), .ZN(n9437)
         );
  MUX2_X1 U10626 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9437), .S(n9826), .Z(
        P1_U3542) );
  NAND2_X1 U10627 ( .A1(n9396), .A2(n9805), .ZN(n9401) );
  AOI22_X1 U10628 ( .A1(n9398), .A2(n9717), .B1(n9422), .B2(n9397), .ZN(n9399)
         );
  OAI211_X1 U10629 ( .C1(n9402), .C2(n9401), .A(n9400), .B(n9399), .ZN(n9438)
         );
  MUX2_X1 U10630 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9438), .S(n9826), .Z(
        P1_U3541) );
  AOI211_X1 U10631 ( .C1(n9422), .C2(n9405), .A(n9404), .B(n9403), .ZN(n9406)
         );
  OAI21_X1 U10632 ( .B1(n9425), .B2(n9407), .A(n9406), .ZN(n9439) );
  MUX2_X1 U10633 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9439), .S(n9826), .Z(
        P1_U3540) );
  AOI211_X1 U10634 ( .C1(n9422), .C2(n9410), .A(n9409), .B(n9408), .ZN(n9411)
         );
  OAI21_X1 U10635 ( .B1(n9425), .B2(n9412), .A(n9411), .ZN(n9440) );
  MUX2_X1 U10636 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9440), .S(n9826), .Z(
        P1_U3539) );
  INV_X1 U10637 ( .A(n9748), .ZN(n9797) );
  AND2_X1 U10638 ( .A1(n9413), .A2(n9797), .ZN(n9417) );
  OAI22_X1 U10639 ( .A1(n9415), .A2(n9801), .B1(n9414), .B2(n9799), .ZN(n9416)
         );
  MUX2_X1 U10640 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9441), .S(n9826), .Z(
        P1_U3538) );
  AOI211_X1 U10641 ( .C1(n9422), .C2(n9421), .A(n9420), .B(n9419), .ZN(n9423)
         );
  OAI21_X1 U10642 ( .B1(n9425), .B2(n9424), .A(n9423), .ZN(n9442) );
  MUX2_X1 U10643 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9442), .S(n9826), .Z(
        P1_U3537) );
  MUX2_X1 U10644 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9426), .S(n9809), .Z(
        P1_U3522) );
  MUX2_X1 U10645 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9427), .S(n9809), .Z(
        P1_U3521) );
  MUX2_X1 U10646 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9428), .S(n9809), .Z(
        P1_U3519) );
  MUX2_X1 U10647 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9429), .S(n9809), .Z(
        P1_U3518) );
  MUX2_X1 U10648 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9430), .S(n9809), .Z(
        P1_U3517) );
  MUX2_X1 U10649 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9431), .S(n9809), .Z(
        P1_U3516) );
  MUX2_X1 U10650 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9432), .S(n9809), .Z(
        P1_U3515) );
  MUX2_X1 U10651 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9433), .S(n9809), .Z(
        P1_U3514) );
  MUX2_X1 U10652 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9434), .S(n9809), .Z(
        P1_U3513) );
  MUX2_X1 U10653 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9435), .S(n9809), .Z(
        P1_U3512) );
  MUX2_X1 U10654 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9436), .S(n9809), .Z(
        P1_U3511) );
  MUX2_X1 U10655 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9437), .S(n9809), .Z(
        P1_U3510) );
  MUX2_X1 U10656 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9438), .S(n9809), .Z(
        P1_U3508) );
  MUX2_X1 U10657 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9439), .S(n9809), .Z(
        P1_U3505) );
  MUX2_X1 U10658 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9440), .S(n9809), .Z(
        P1_U3502) );
  MUX2_X1 U10659 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9441), .S(n9809), .Z(
        P1_U3499) );
  MUX2_X1 U10660 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9442), .S(n9809), .Z(
        P1_U3496) );
  NAND3_X1 U10661 ( .A1(n5594), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n9445) );
  OAI22_X1 U10662 ( .A1(n9443), .A2(n9445), .B1(n6334), .B2(n9444), .ZN(n9446)
         );
  AOI21_X1 U10663 ( .B1(n9448), .B2(n9447), .A(n9446), .ZN(n9449) );
  INV_X1 U10664 ( .A(n9449), .ZN(P1_U3322) );
  MUX2_X1 U10665 ( .A(n9450), .B(n9556), .S(P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U10666 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n9451) );
  OAI22_X1 U10667 ( .A1(n9453), .A2(n9452), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9451), .ZN(n9454) );
  AOI21_X1 U10668 ( .B1(n9456), .B2(n9455), .A(n9454), .ZN(n9466) );
  NOR2_X1 U10669 ( .A1(n9457), .A2(n9799), .ZN(n9531) );
  NAND2_X1 U10670 ( .A1(n9459), .A2(n9458), .ZN(n9461) );
  AOI21_X1 U10671 ( .B1(n9462), .B2(n9461), .A(n9460), .ZN(n9463) );
  AOI21_X1 U10672 ( .B1(n9464), .B2(n9531), .A(n9463), .ZN(n9465) );
  OAI211_X1 U10673 ( .C1(n9468), .C2(n9467), .A(n9466), .B(n9465), .ZN(
        P1_U3222) );
  AOI22_X1 U10674 ( .A1(n9844), .A2(n9469), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        n10007), .ZN(n9481) );
  AND2_X1 U10675 ( .A1(n9471), .A2(n9470), .ZN(n9474) );
  OAI21_X1 U10676 ( .B1(n9474), .B2(n9473), .A(n9472), .ZN(n9479) );
  NAND2_X1 U10677 ( .A1(n9476), .A2(n9475), .ZN(n9483) );
  INV_X1 U10678 ( .A(n9483), .ZN(n9477) );
  AOI22_X1 U10679 ( .A1(n9479), .A2(n9845), .B1(n9478), .B2(n9477), .ZN(n9480)
         );
  OAI211_X1 U10680 ( .C1(n9860), .C2(n9482), .A(n9481), .B(n9480), .ZN(
        P2_U3217) );
  OAI211_X1 U10681 ( .C1(n9936), .C2(n9485), .A(n9484), .B(n9483), .ZN(n9486)
         );
  AOI21_X1 U10682 ( .B1(n9487), .B2(n9931), .A(n9486), .ZN(n9489) );
  AOI22_X1 U10683 ( .A1(n9954), .A2(n9489), .B1(n7218), .B2(n9952), .ZN(
        P2_U3534) );
  INV_X1 U10684 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9488) );
  AOI22_X1 U10685 ( .A1(n9944), .A2(n9489), .B1(n9488), .B2(n9942), .ZN(
        P2_U3493) );
  XOR2_X1 U10686 ( .A(n9490), .B(n9494), .Z(n9527) );
  INV_X1 U10687 ( .A(n9491), .ZN(n9492) );
  AOI21_X1 U10688 ( .B1(n9494), .B2(n9493), .A(n9492), .ZN(n9495) );
  OAI222_X1 U10689 ( .A1(n9699), .A2(n9512), .B1(n9701), .B2(n9496), .C1(n9733), .C2(n9495), .ZN(n9525) );
  AOI21_X1 U10690 ( .B1(n9730), .B2(n9527), .A(n9525), .ZN(n9504) );
  AOI222_X1 U10691 ( .A1(n9499), .A2(n9498), .B1(P1_REG2_REG_13__SCAN_IN), 
        .B2(n9739), .C1(n9718), .C2(n9497), .ZN(n9503) );
  OAI21_X1 U10692 ( .B1(n4563), .B2(n9500), .A(n4329), .ZN(n9524) );
  INV_X1 U10693 ( .A(n9524), .ZN(n9501) );
  AOI22_X1 U10694 ( .A1(n9527), .A2(n9697), .B1(n9696), .B2(n9501), .ZN(n9502)
         );
  OAI211_X1 U10695 ( .C1(n9739), .C2(n9504), .A(n9503), .B(n9502), .ZN(
        P1_U3278) );
  XNOR2_X1 U10696 ( .A(n9505), .B(n9511), .ZN(n9517) );
  INV_X1 U10697 ( .A(n9517), .ZN(n9539) );
  OAI21_X1 U10698 ( .B1(n9507), .B2(n9535), .A(n9506), .ZN(n9536) );
  INV_X1 U10699 ( .A(n9536), .ZN(n9508) );
  AOI22_X1 U10700 ( .A1(n9539), .A2(n9697), .B1(n9696), .B2(n9508), .ZN(n9523)
         );
  OAI21_X1 U10701 ( .B1(n9511), .B2(n9510), .A(n9509), .ZN(n9515) );
  OAI22_X1 U10702 ( .A1(n9513), .A2(n9699), .B1(n9512), .B2(n9701), .ZN(n9514)
         );
  AOI21_X1 U10703 ( .B1(n9515), .B2(n9704), .A(n9514), .ZN(n9516) );
  OAI21_X1 U10704 ( .B1(n9517), .B2(n9707), .A(n9516), .ZN(n9537) );
  NOR2_X1 U10705 ( .A1(n9535), .A2(n9710), .ZN(n9521) );
  INV_X1 U10706 ( .A(n9518), .ZN(n9519) );
  OAI22_X1 U10707 ( .A1(n9737), .A2(n6518), .B1(n9519), .B2(n9709), .ZN(n9520)
         );
  AOI211_X1 U10708 ( .C1(n9537), .C2(n9737), .A(n9521), .B(n9520), .ZN(n9522)
         );
  NAND2_X1 U10709 ( .A1(n9523), .A2(n9522), .ZN(P1_U3280) );
  OAI22_X1 U10710 ( .A1(n9524), .A2(n9801), .B1(n4563), .B2(n9799), .ZN(n9526)
         );
  AOI211_X1 U10711 ( .C1(n9527), .C2(n9805), .A(n9526), .B(n9525), .ZN(n9541)
         );
  AOI22_X1 U10712 ( .A1(n9826), .A2(n9541), .B1(n9528), .B2(n9823), .ZN(
        P1_U3536) );
  NOR2_X1 U10713 ( .A1(n9529), .A2(n9748), .ZN(n9532) );
  NOR4_X1 U10714 ( .A1(n9533), .A2(n9532), .A3(n9531), .A4(n9530), .ZN(n9543)
         );
  AOI22_X1 U10715 ( .A1(n9826), .A2(n9543), .B1(n9534), .B2(n9823), .ZN(
        P1_U3535) );
  OAI22_X1 U10716 ( .A1(n9536), .A2(n9801), .B1(n9535), .B2(n9799), .ZN(n9538)
         );
  AOI211_X1 U10717 ( .C1(n9797), .C2(n9539), .A(n9538), .B(n9537), .ZN(n9545)
         );
  AOI22_X1 U10718 ( .A1(n9826), .A2(n9545), .B1(n6493), .B2(n9823), .ZN(
        P1_U3534) );
  AOI22_X1 U10719 ( .A1(n9809), .A2(n9541), .B1(n9540), .B2(n9807), .ZN(
        P1_U3493) );
  INV_X1 U10720 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9542) );
  AOI22_X1 U10721 ( .A1(n9809), .A2(n9543), .B1(n9542), .B2(n9807), .ZN(
        P1_U3490) );
  INV_X1 U10722 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9544) );
  AOI22_X1 U10723 ( .A1(n9809), .A2(n9545), .B1(n9544), .B2(n9807), .ZN(
        P1_U3487) );
  XNOR2_X1 U10724 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10725 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  NOR2_X1 U10726 ( .A1(n9546), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9547) );
  OR2_X1 U10727 ( .A1(n9547), .A2(n6141), .ZN(n9548) );
  XNOR2_X1 U10728 ( .A(n9548), .B(n9556), .ZN(n9581) );
  INV_X1 U10729 ( .A(n9549), .ZN(n9550) );
  NAND3_X1 U10730 ( .A1(n9551), .A2(n9550), .A3(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9552) );
  NAND2_X1 U10731 ( .A1(n9553), .A2(n9552), .ZN(n9554) );
  AOI22_X1 U10732 ( .A1(n9661), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(n9581), .B2(
        n9554), .ZN(n9558) );
  NAND3_X1 U10733 ( .A1(n9663), .A2(n9556), .A3(n9555), .ZN(n9557) );
  OAI211_X1 U10734 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n6801), .A(n9558), .B(
        n9557), .ZN(P1_U3241) );
  INV_X1 U10735 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9559) );
  OAI22_X1 U10736 ( .A1(n9658), .A2(n9560), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9559), .ZN(n9561) );
  AOI21_X1 U10737 ( .B1(n9661), .B2(P1_ADDR_REG_1__SCAN_IN), .A(n9561), .ZN(
        n9569) );
  OAI211_X1 U10738 ( .C1(n9563), .C2(n9562), .A(n9663), .B(n9571), .ZN(n9568)
         );
  OAI211_X1 U10739 ( .C1(n9566), .C2(n9565), .A(n9667), .B(n9564), .ZN(n9567)
         );
  NAND3_X1 U10740 ( .A1(n9569), .A2(n9568), .A3(n9567), .ZN(P1_U3242) );
  INV_X1 U10741 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9590) );
  MUX2_X1 U10742 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9811), .S(n9576), .Z(n9572)
         );
  NAND3_X1 U10743 ( .A1(n9572), .A2(n9571), .A3(n9570), .ZN(n9573) );
  NAND3_X1 U10744 ( .A1(n9663), .A2(n9574), .A3(n9573), .ZN(n9575) );
  OAI21_X1 U10745 ( .B1(n9658), .B2(n9576), .A(n9575), .ZN(n9584) );
  OR2_X1 U10746 ( .A1(n9577), .A2(n6141), .ZN(n9578) );
  INV_X1 U10747 ( .A(n9578), .ZN(n9582) );
  OR2_X1 U10748 ( .A1(n9579), .A2(n9578), .ZN(n9580) );
  OAI211_X1 U10749 ( .C1(n9582), .C2(n9581), .A(n9580), .B(P1_U4006), .ZN(
        n9601) );
  INV_X1 U10750 ( .A(n9601), .ZN(n9583) );
  AOI211_X1 U10751 ( .C1(n9661), .C2(P1_ADDR_REG_2__SCAN_IN), .A(n9584), .B(
        n9583), .ZN(n9589) );
  OAI211_X1 U10752 ( .C1(n9587), .C2(n9586), .A(n9667), .B(n9585), .ZN(n9588)
         );
  OAI211_X1 U10753 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n9590), .A(n9589), .B(
        n9588), .ZN(P1_U3243) );
  OAI21_X1 U10754 ( .B1(n9593), .B2(n9592), .A(n9591), .ZN(n9595) );
  AOI222_X1 U10755 ( .A1(n9595), .A2(n9667), .B1(n9661), .B2(
        P1_ADDR_REG_4__SCAN_IN), .C1(n9594), .C2(n9636), .ZN(n9603) );
  OAI21_X1 U10756 ( .B1(n9598), .B2(n9597), .A(n9596), .ZN(n9599) );
  NAND2_X1 U10757 ( .A1(n9663), .A2(n9599), .ZN(n9600) );
  NAND4_X1 U10758 ( .A1(n9603), .A2(n9602), .A3(n9601), .A4(n9600), .ZN(
        P1_U3245) );
  AOI21_X1 U10759 ( .B1(n9606), .B2(n9605), .A(n9604), .ZN(n9607) );
  NOR2_X1 U10760 ( .A1(n9607), .A2(n9621), .ZN(n9608) );
  AOI211_X1 U10761 ( .C1(n9636), .C2(n9610), .A(n9609), .B(n9608), .ZN(n9615)
         );
  OAI211_X1 U10762 ( .C1(n9613), .C2(n9612), .A(n9611), .B(n9667), .ZN(n9614)
         );
  OAI211_X1 U10763 ( .C1(n9996), .C2(n9632), .A(n9615), .B(n9614), .ZN(
        P1_U3250) );
  INV_X1 U10764 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9631) );
  AOI21_X1 U10765 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9617), .A(n9616), .ZN(
        n9628) );
  AOI21_X1 U10766 ( .B1(n9620), .B2(n9619), .A(n9618), .ZN(n9622) );
  OR2_X1 U10767 ( .A1(n9622), .A2(n9621), .ZN(n9626) );
  AOI21_X1 U10768 ( .B1(n9636), .B2(n9624), .A(n9623), .ZN(n9625) );
  OAI211_X1 U10769 ( .C1(n9628), .C2(n9627), .A(n9626), .B(n9625), .ZN(n9629)
         );
  INV_X1 U10770 ( .A(n9629), .ZN(n9630) );
  OAI21_X1 U10771 ( .B1(n9632), .B2(n9631), .A(n9630), .ZN(P1_U3255) );
  INV_X1 U10772 ( .A(n9633), .ZN(n9634) );
  AOI21_X1 U10773 ( .B1(n9636), .B2(n9635), .A(n9634), .ZN(n9644) );
  OAI211_X1 U10774 ( .C1(n9638), .C2(P1_REG1_REG_15__SCAN_IN), .A(n9663), .B(
        n9637), .ZN(n9643) );
  NAND2_X1 U10775 ( .A1(n9661), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n9642) );
  OAI211_X1 U10776 ( .C1(n9640), .C2(P1_REG2_REG_15__SCAN_IN), .A(n9667), .B(
        n9639), .ZN(n9641) );
  NAND4_X1 U10777 ( .A1(n9644), .A2(n9643), .A3(n9642), .A4(n9641), .ZN(
        P1_U3256) );
  NOR2_X1 U10778 ( .A1(n9658), .A2(n9645), .ZN(n9646) );
  AOI211_X1 U10779 ( .C1(P1_ADDR_REG_16__SCAN_IN), .C2(n9661), .A(n9647), .B(
        n9646), .ZN(n9656) );
  OAI211_X1 U10780 ( .C1(n9650), .C2(n9649), .A(n9663), .B(n9648), .ZN(n9655)
         );
  OAI211_X1 U10781 ( .C1(n9653), .C2(n9652), .A(n9667), .B(n9651), .ZN(n9654)
         );
  NAND3_X1 U10782 ( .A1(n9656), .A2(n9655), .A3(n9654), .ZN(P1_U3257) );
  NOR2_X1 U10783 ( .A1(n9658), .A2(n9657), .ZN(n9659) );
  AOI211_X1 U10784 ( .C1(n9661), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n9660), .B(
        n9659), .ZN(n9672) );
  OAI211_X1 U10785 ( .C1(n9665), .C2(n9664), .A(n9663), .B(n9662), .ZN(n9671)
         );
  OAI211_X1 U10786 ( .C1(n9669), .C2(n9668), .A(n9667), .B(n9666), .ZN(n9670)
         );
  NAND3_X1 U10787 ( .A1(n9672), .A2(n9671), .A3(n9670), .ZN(P1_U3258) );
  XNOR2_X1 U10788 ( .A(n9673), .B(n9680), .ZN(n9674) );
  NAND2_X1 U10789 ( .A1(n9674), .A2(n9704), .ZN(n9678) );
  AOI22_X1 U10790 ( .A1(n9726), .A2(n9676), .B1(n9675), .B2(n9729), .ZN(n9677)
         );
  NAND2_X1 U10791 ( .A1(n9678), .A2(n9677), .ZN(n9775) );
  INV_X1 U10792 ( .A(n9680), .ZN(n9681) );
  XNOR2_X1 U10793 ( .A(n9679), .B(n9681), .ZN(n9769) );
  AND2_X1 U10794 ( .A1(n9769), .A2(n9682), .ZN(n9690) );
  AOI21_X1 U10795 ( .B1(n9683), .B2(n9687), .A(n9801), .ZN(n9685) );
  NAND2_X1 U10796 ( .A1(n9685), .A2(n9684), .ZN(n9772) );
  AOI22_X1 U10797 ( .A1(n4342), .A2(n9687), .B1(n9718), .B2(n9686), .ZN(n9688)
         );
  OAI21_X1 U10798 ( .B1(n9772), .B2(n9721), .A(n9688), .ZN(n9689) );
  NOR3_X1 U10799 ( .A1(n9775), .A2(n9690), .A3(n9689), .ZN(n9691) );
  AOI22_X1 U10800 ( .A1(n9739), .A2(n6349), .B1(n9691), .B2(n9737), .ZN(
        P1_U3286) );
  XOR2_X1 U10801 ( .A(n9692), .B(n9698), .Z(n9708) );
  INV_X1 U10802 ( .A(n9708), .ZN(n9762) );
  OAI21_X1 U10803 ( .B1(n9694), .B2(n6927), .A(n9693), .ZN(n9759) );
  INV_X1 U10804 ( .A(n9759), .ZN(n9695) );
  AOI22_X1 U10805 ( .A1(n9762), .A2(n9697), .B1(n9696), .B2(n9695), .ZN(n9714)
         );
  OAI22_X1 U10806 ( .A1(n9702), .A2(n9701), .B1(n9700), .B2(n9699), .ZN(n9703)
         );
  AOI21_X1 U10807 ( .B1(n9705), .B2(n9704), .A(n9703), .ZN(n9706) );
  OAI21_X1 U10808 ( .B1(n9708), .B2(n9707), .A(n9706), .ZN(n9760) );
  MUX2_X1 U10809 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n9760), .S(n9737), .Z(n9712)
         );
  OAI22_X1 U10810 ( .A1(n9710), .A2(n6927), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9709), .ZN(n9711) );
  NOR2_X1 U10811 ( .A1(n9712), .A2(n9711), .ZN(n9713) );
  NAND2_X1 U10812 ( .A1(n9714), .A2(n9713), .ZN(P1_U3288) );
  XNOR2_X1 U10813 ( .A(n9724), .B(n9715), .ZN(n9745) );
  OAI211_X1 U10814 ( .C1(n6714), .C2(n4558), .A(n9717), .B(n9716), .ZN(n9746)
         );
  AOI22_X1 U10815 ( .A1(n4342), .A2(n9719), .B1(n9718), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n9720) );
  OAI21_X1 U10816 ( .B1(n9746), .B2(n9721), .A(n9720), .ZN(n9735) );
  INV_X1 U10817 ( .A(n9722), .ZN(n9723) );
  AOI21_X1 U10818 ( .B1(n9725), .B2(n9724), .A(n9723), .ZN(n9734) );
  AOI22_X1 U10819 ( .A1(n9729), .A2(n9728), .B1(n9727), .B2(n9726), .ZN(n9732)
         );
  NAND2_X1 U10820 ( .A1(n9745), .A2(n9730), .ZN(n9731) );
  OAI211_X1 U10821 ( .C1(n9734), .C2(n9733), .A(n9732), .B(n9731), .ZN(n9751)
         );
  AOI211_X1 U10822 ( .C1(n9736), .C2(n9745), .A(n9735), .B(n9751), .ZN(n9738)
         );
  AOI22_X1 U10823 ( .A1(n9739), .A2(n6342), .B1(n9738), .B2(n9737), .ZN(
        P1_U3290) );
  AND2_X1 U10824 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9744), .ZN(P1_U3292) );
  AND2_X1 U10825 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9744), .ZN(P1_U3293) );
  AND2_X1 U10826 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9744), .ZN(P1_U3294) );
  AND2_X1 U10827 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9744), .ZN(P1_U3295) );
  AND2_X1 U10828 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9744), .ZN(P1_U3296) );
  NOR2_X1 U10829 ( .A1(n9743), .A2(n9740), .ZN(P1_U3297) );
  AND2_X1 U10830 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9744), .ZN(P1_U3298) );
  AND2_X1 U10831 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9744), .ZN(P1_U3299) );
  AND2_X1 U10832 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9744), .ZN(P1_U3300) );
  AND2_X1 U10833 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9744), .ZN(P1_U3301) );
  AND2_X1 U10834 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9744), .ZN(P1_U3302) );
  AND2_X1 U10835 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9744), .ZN(P1_U3303) );
  AND2_X1 U10836 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9744), .ZN(P1_U3304) );
  AND2_X1 U10837 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9744), .ZN(P1_U3305) );
  AND2_X1 U10838 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9744), .ZN(P1_U3306) );
  AND2_X1 U10839 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9744), .ZN(P1_U3307) );
  AND2_X1 U10840 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9744), .ZN(P1_U3308) );
  AND2_X1 U10841 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9744), .ZN(P1_U3309) );
  AND2_X1 U10842 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9744), .ZN(P1_U3310) );
  NOR2_X1 U10843 ( .A1(n9743), .A2(n9741), .ZN(P1_U3311) );
  AND2_X1 U10844 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9744), .ZN(P1_U3312) );
  AND2_X1 U10845 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9744), .ZN(P1_U3313) );
  AND2_X1 U10846 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9744), .ZN(P1_U3314) );
  NOR2_X1 U10847 ( .A1(n9743), .A2(n9742), .ZN(P1_U3315) );
  AND2_X1 U10848 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9744), .ZN(P1_U3316) );
  AND2_X1 U10849 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9744), .ZN(P1_U3317) );
  AND2_X1 U10850 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9744), .ZN(P1_U3318) );
  AND2_X1 U10851 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9744), .ZN(P1_U3319) );
  AND2_X1 U10852 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9744), .ZN(P1_U3320) );
  AND2_X1 U10853 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9744), .ZN(P1_U3321) );
  INV_X1 U10854 ( .A(n9745), .ZN(n9749) );
  OAI211_X1 U10855 ( .C1(n9749), .C2(n9748), .A(n9747), .B(n9746), .ZN(n9750)
         );
  NOR2_X1 U10856 ( .A1(n9751), .A2(n9750), .ZN(n9810) );
  AOI22_X1 U10857 ( .A1(n9809), .A2(n9810), .B1(n9752), .B2(n9807), .ZN(
        P1_U3457) );
  INV_X1 U10858 ( .A(n9753), .ZN(n9754) );
  OAI22_X1 U10859 ( .A1(n9754), .A2(n9801), .B1(n6718), .B2(n9799), .ZN(n9756)
         );
  AOI211_X1 U10860 ( .C1(n9797), .C2(n9757), .A(n9756), .B(n9755), .ZN(n9812)
         );
  INV_X1 U10861 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9758) );
  AOI22_X1 U10862 ( .A1(n9809), .A2(n9812), .B1(n9758), .B2(n9807), .ZN(
        P1_U3460) );
  OAI22_X1 U10863 ( .A1(n9759), .A2(n9801), .B1(n6927), .B2(n9799), .ZN(n9761)
         );
  AOI211_X1 U10864 ( .C1(n9797), .C2(n9762), .A(n9761), .B(n9760), .ZN(n9813)
         );
  INV_X1 U10865 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9763) );
  AOI22_X1 U10866 ( .A1(n9809), .A2(n9813), .B1(n9763), .B2(n9807), .ZN(
        P1_U3463) );
  OAI22_X1 U10867 ( .A1(n9765), .A2(n9801), .B1(n9764), .B2(n9799), .ZN(n9767)
         );
  AOI211_X1 U10868 ( .C1(n9797), .C2(n9768), .A(n9767), .B(n9766), .ZN(n9815)
         );
  AOI22_X1 U10869 ( .A1(n9809), .A2(n9815), .B1(n5695), .B2(n9807), .ZN(
        P1_U3466) );
  AND2_X1 U10870 ( .A1(n9769), .A2(n9805), .ZN(n9774) );
  INV_X1 U10871 ( .A(n9770), .ZN(n9771) );
  NAND2_X1 U10872 ( .A1(n9772), .A2(n9771), .ZN(n9773) );
  NOR3_X1 U10873 ( .A1(n9775), .A2(n9774), .A3(n9773), .ZN(n9817) );
  INV_X1 U10874 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9776) );
  AOI22_X1 U10875 ( .A1(n9809), .A2(n9817), .B1(n9776), .B2(n9807), .ZN(
        P1_U3469) );
  INV_X1 U10876 ( .A(n9777), .ZN(n9778) );
  OAI21_X1 U10877 ( .B1(n9779), .B2(n9801), .A(n9778), .ZN(n9781) );
  AOI211_X1 U10878 ( .C1(n9797), .C2(n9782), .A(n9781), .B(n9780), .ZN(n9819)
         );
  INV_X1 U10879 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9783) );
  AOI22_X1 U10880 ( .A1(n9809), .A2(n9819), .B1(n9783), .B2(n9807), .ZN(
        P1_U3472) );
  INV_X1 U10881 ( .A(n9784), .ZN(n9786) );
  NAND3_X1 U10882 ( .A1(n9787), .A2(n9786), .A3(n9785), .ZN(n9788) );
  AOI21_X1 U10883 ( .B1(n9805), .B2(n9789), .A(n9788), .ZN(n9821) );
  INV_X1 U10884 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9790) );
  AOI22_X1 U10885 ( .A1(n9809), .A2(n9821), .B1(n9790), .B2(n9807), .ZN(
        P1_U3475) );
  INV_X1 U10886 ( .A(n9791), .ZN(n9796) );
  OAI21_X1 U10887 ( .B1(n9793), .B2(n9801), .A(n9792), .ZN(n9795) );
  AOI211_X1 U10888 ( .C1(n9797), .C2(n9796), .A(n9795), .B(n9794), .ZN(n9822)
         );
  INV_X1 U10889 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9798) );
  AOI22_X1 U10890 ( .A1(n9809), .A2(n9822), .B1(n9798), .B2(n9807), .ZN(
        P1_U3478) );
  OAI22_X1 U10891 ( .A1(n9802), .A2(n9801), .B1(n9800), .B2(n9799), .ZN(n9804)
         );
  AOI211_X1 U10892 ( .C1(n9806), .C2(n9805), .A(n9804), .B(n9803), .ZN(n9825)
         );
  INV_X1 U10893 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9808) );
  AOI22_X1 U10894 ( .A1(n9809), .A2(n9825), .B1(n9808), .B2(n9807), .ZN(
        P1_U3481) );
  AOI22_X1 U10895 ( .A1(n9826), .A2(n9810), .B1(n6356), .B2(n9823), .ZN(
        P1_U3524) );
  AOI22_X1 U10896 ( .A1(n9826), .A2(n9812), .B1(n9811), .B2(n9823), .ZN(
        P1_U3525) );
  AOI22_X1 U10897 ( .A1(n9826), .A2(n9813), .B1(n6359), .B2(n9823), .ZN(
        P1_U3526) );
  AOI22_X1 U10898 ( .A1(n9826), .A2(n9815), .B1(n9814), .B2(n9823), .ZN(
        P1_U3527) );
  AOI22_X1 U10899 ( .A1(n9826), .A2(n9817), .B1(n9816), .B2(n9823), .ZN(
        P1_U3528) );
  AOI22_X1 U10900 ( .A1(n9826), .A2(n9819), .B1(n9818), .B2(n9823), .ZN(
        P1_U3529) );
  AOI22_X1 U10901 ( .A1(n9826), .A2(n9821), .B1(n9820), .B2(n9823), .ZN(
        P1_U3530) );
  AOI22_X1 U10902 ( .A1(n9826), .A2(n9822), .B1(n6395), .B2(n9823), .ZN(
        P1_U3531) );
  AOI22_X1 U10903 ( .A1(n9826), .A2(n9825), .B1(n9824), .B2(n9823), .ZN(
        P1_U3532) );
  NAND2_X1 U10904 ( .A1(n9828), .A2(n9827), .ZN(n9830) );
  OAI211_X1 U10905 ( .C1(n9832), .C2(n9831), .A(n9830), .B(n9829), .ZN(n9839)
         );
  INV_X1 U10906 ( .A(n9833), .ZN(n9834) );
  AOI211_X1 U10907 ( .C1(n9837), .C2(n9836), .A(n9835), .B(n9834), .ZN(n9838)
         );
  AOI211_X1 U10908 ( .C1(n9854), .C2(n9840), .A(n9839), .B(n9838), .ZN(n9841)
         );
  OAI21_X1 U10909 ( .B1(n9860), .B2(n9842), .A(n9841), .ZN(P2_U3219) );
  AOI22_X1 U10910 ( .A1(n9844), .A2(n9843), .B1(P2_REG3_REG_8__SCAN_IN), .B2(
        P2_U3152), .ZN(n9858) );
  OAI21_X1 U10911 ( .B1(n9847), .B2(n9846), .A(n9845), .ZN(n9852) );
  NAND3_X1 U10912 ( .A1(n9850), .A2(n9849), .A3(n9848), .ZN(n9851) );
  NAND2_X1 U10913 ( .A1(n9852), .A2(n9851), .ZN(n9856) );
  AOI22_X1 U10914 ( .A1(n9856), .A2(n9855), .B1(n9854), .B2(n9853), .ZN(n9857)
         );
  OAI211_X1 U10915 ( .C1(n9860), .C2(n9859), .A(n9858), .B(n9857), .ZN(
        P2_U3223) );
  AOI22_X1 U10916 ( .A1(n9879), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9871), .ZN(n9868) );
  INV_X1 U10917 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9864) );
  OAI21_X1 U10918 ( .B1(n9862), .B2(P2_REG1_REG_0__SCAN_IN), .A(n9861), .ZN(
        n9863) );
  AOI21_X1 U10919 ( .B1(n9879), .B2(n9864), .A(n9863), .ZN(n9866) );
  AOI22_X1 U10920 ( .A1(n9870), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9865) );
  OAI221_X1 U10921 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9868), .C1(n9867), .C2(
        n9866), .A(n9865), .ZN(P2_U3245) );
  AOI21_X1 U10922 ( .B1(n9870), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n9869), .ZN(
        n9884) );
  OAI211_X1 U10923 ( .C1(n9874), .C2(n9873), .A(n9872), .B(n9871), .ZN(n9883)
         );
  NAND2_X1 U10924 ( .A1(n9876), .A2(n9875), .ZN(n9882) );
  XOR2_X1 U10925 ( .A(n9878), .B(n9877), .Z(n9880) );
  NAND2_X1 U10926 ( .A1(n9880), .A2(n9879), .ZN(n9881) );
  NAND4_X1 U10927 ( .A1(n9884), .A2(n9883), .A3(n9882), .A4(n9881), .ZN(
        P2_U3262) );
  AND2_X1 U10928 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9890), .ZN(P2_U3297) );
  AND2_X1 U10929 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9890), .ZN(P2_U3298) );
  AND2_X1 U10930 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9890), .ZN(P2_U3299) );
  AND2_X1 U10931 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9890), .ZN(P2_U3300) );
  AND2_X1 U10932 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9890), .ZN(P2_U3301) );
  AND2_X1 U10933 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9890), .ZN(P2_U3302) );
  INV_X1 U10934 ( .A(n9890), .ZN(n9894) );
  NOR2_X1 U10935 ( .A1(n9894), .A2(n9887), .ZN(P2_U3303) );
  AND2_X1 U10936 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9890), .ZN(P2_U3304) );
  AND2_X1 U10937 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9890), .ZN(P2_U3305) );
  AND2_X1 U10938 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9890), .ZN(P2_U3306) );
  AND2_X1 U10939 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9890), .ZN(P2_U3307) );
  AND2_X1 U10940 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9890), .ZN(P2_U3308) );
  AND2_X1 U10941 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9890), .ZN(P2_U3309) );
  NOR2_X1 U10942 ( .A1(n9894), .A2(n9888), .ZN(P2_U3310) );
  AND2_X1 U10943 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9890), .ZN(P2_U3311) );
  AND2_X1 U10944 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9890), .ZN(P2_U3312) );
  NOR2_X1 U10945 ( .A1(n9894), .A2(n9889), .ZN(P2_U3313) );
  AND2_X1 U10946 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9890), .ZN(P2_U3314) );
  AND2_X1 U10947 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9890), .ZN(P2_U3315) );
  AND2_X1 U10948 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9890), .ZN(P2_U3316) );
  AND2_X1 U10949 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9890), .ZN(P2_U3317) );
  AND2_X1 U10950 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9890), .ZN(P2_U3318) );
  AND2_X1 U10951 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9890), .ZN(P2_U3319) );
  AND2_X1 U10952 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9890), .ZN(P2_U3320) );
  AND2_X1 U10953 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9890), .ZN(P2_U3321) );
  AND2_X1 U10954 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9890), .ZN(P2_U3322) );
  AND2_X1 U10955 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9890), .ZN(P2_U3323) );
  AND2_X1 U10956 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9890), .ZN(P2_U3324) );
  AND2_X1 U10957 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9890), .ZN(P2_U3325) );
  AND2_X1 U10958 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9890), .ZN(P2_U3326) );
  INV_X1 U10959 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9891) );
  AOI22_X1 U10960 ( .A1(n9893), .A2(n9892), .B1(n9891), .B2(n9890), .ZN(
        P2_U3437) );
  INV_X1 U10961 ( .A(n9893), .ZN(n9896) );
  OAI22_X1 U10962 ( .A1(n9896), .A2(n9895), .B1(P2_D_REG_1__SCAN_IN), .B2(
        n9894), .ZN(n9897) );
  INV_X1 U10963 ( .A(n9897), .ZN(P2_U3438) );
  AOI22_X1 U10964 ( .A1(n9900), .A2(n9931), .B1(n9899), .B2(n9898), .ZN(n9901)
         );
  AND2_X1 U10965 ( .A1(n9902), .A2(n9901), .ZN(n9946) );
  INV_X1 U10966 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9903) );
  AOI22_X1 U10967 ( .A1(n9944), .A2(n9946), .B1(n9903), .B2(n9942), .ZN(
        P2_U3451) );
  INV_X1 U10968 ( .A(n9904), .ZN(n9909) );
  OAI211_X1 U10969 ( .C1(n9907), .C2(n9934), .A(n9906), .B(n9905), .ZN(n9908)
         );
  AOI21_X1 U10970 ( .B1(n9909), .B2(n9931), .A(n9908), .ZN(n9948) );
  INV_X1 U10971 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9910) );
  AOI22_X1 U10972 ( .A1(n9944), .A2(n9948), .B1(n9910), .B2(n9942), .ZN(
        P2_U3454) );
  NAND3_X1 U10973 ( .A1(n9913), .A2(n9912), .A3(n9911), .ZN(n9914) );
  OAI211_X1 U10974 ( .C1(n9916), .C2(n9934), .A(n9915), .B(n9914), .ZN(n9917)
         );
  AOI21_X1 U10975 ( .B1(n9918), .B2(n9931), .A(n9917), .ZN(n9949) );
  INV_X1 U10976 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9919) );
  AOI22_X1 U10977 ( .A1(n9944), .A2(n9949), .B1(n9919), .B2(n9942), .ZN(
        P2_U3457) );
  OAI22_X1 U10978 ( .A1(n9921), .A2(n9936), .B1(n9920), .B2(n9934), .ZN(n9923)
         );
  AOI211_X1 U10979 ( .C1(n9931), .C2(n9924), .A(n9923), .B(n9922), .ZN(n9950)
         );
  INV_X1 U10980 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9925) );
  AOI22_X1 U10981 ( .A1(n9944), .A2(n9950), .B1(n9925), .B2(n9942), .ZN(
        P2_U3463) );
  OAI22_X1 U10982 ( .A1(n9927), .A2(n9936), .B1(n9926), .B2(n9934), .ZN(n9929)
         );
  AOI211_X1 U10983 ( .C1(n9931), .C2(n9930), .A(n9929), .B(n9928), .ZN(n9951)
         );
  INV_X1 U10984 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9932) );
  AOI22_X1 U10985 ( .A1(n9944), .A2(n9951), .B1(n9932), .B2(n9942), .ZN(
        P2_U3469) );
  INV_X1 U10986 ( .A(n9933), .ZN(n9940) );
  OAI22_X1 U10987 ( .A1(n9937), .A2(n9936), .B1(n9935), .B2(n9934), .ZN(n9939)
         );
  AOI211_X1 U10988 ( .C1(n9941), .C2(n9940), .A(n9939), .B(n9938), .ZN(n9953)
         );
  INV_X1 U10989 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9943) );
  AOI22_X1 U10990 ( .A1(n9944), .A2(n9953), .B1(n9943), .B2(n9942), .ZN(
        P2_U3481) );
  AOI22_X1 U10991 ( .A1(n9954), .A2(n9946), .B1(n9945), .B2(n9952), .ZN(
        P2_U3520) );
  INV_X1 U10992 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9947) );
  AOI22_X1 U10993 ( .A1(n9954), .A2(n9948), .B1(n9947), .B2(n9952), .ZN(
        P2_U3521) );
  AOI22_X1 U10994 ( .A1(n9954), .A2(n9949), .B1(n6213), .B2(n9952), .ZN(
        P2_U3522) );
  AOI22_X1 U10995 ( .A1(n9954), .A2(n9950), .B1(n6214), .B2(n9952), .ZN(
        P2_U3524) );
  AOI22_X1 U10996 ( .A1(n9954), .A2(n9951), .B1(n6215), .B2(n9952), .ZN(
        P2_U3526) );
  AOI22_X1 U10997 ( .A1(n9954), .A2(n9953), .B1(n6667), .B2(n9952), .ZN(
        P2_U3530) );
  INV_X1 U10998 ( .A(n9955), .ZN(n9956) );
  NAND2_X1 U10999 ( .A1(n9957), .A2(n9956), .ZN(n9958) );
  XNOR2_X1 U11000 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9958), .ZN(ADD_1071_U5) );
  XOR2_X1 U11001 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11002 ( .B1(n9961), .B2(n9960), .A(n9959), .ZN(ADD_1071_U56) );
  OAI21_X1 U11003 ( .B1(n9964), .B2(n9963), .A(n9962), .ZN(ADD_1071_U57) );
  OAI21_X1 U11004 ( .B1(n9967), .B2(n9966), .A(n9965), .ZN(ADD_1071_U58) );
  OAI21_X1 U11005 ( .B1(n9970), .B2(n9969), .A(n9968), .ZN(ADD_1071_U59) );
  OAI21_X1 U11006 ( .B1(n9973), .B2(n9972), .A(n9971), .ZN(ADD_1071_U60) );
  OAI21_X1 U11007 ( .B1(n9976), .B2(n9975), .A(n9974), .ZN(ADD_1071_U61) );
  AOI21_X1 U11008 ( .B1(n9979), .B2(n9978), .A(n9977), .ZN(ADD_1071_U62) );
  AOI21_X1 U11009 ( .B1(n9982), .B2(n9981), .A(n9980), .ZN(ADD_1071_U63) );
  XNOR2_X1 U11010 ( .A(n9984), .B(n9983), .ZN(ADD_1071_U48) );
  XNOR2_X1 U11011 ( .A(n9986), .B(n9985), .ZN(ADD_1071_U50) );
  NOR2_X1 U11012 ( .A1(n9988), .A2(n9987), .ZN(n9989) );
  XOR2_X1 U11013 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n9989), .Z(ADD_1071_U51) );
  OAI21_X1 U11014 ( .B1(n9992), .B2(n9991), .A(n9990), .ZN(n9993) );
  XNOR2_X1 U11015 ( .A(n9993), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11016 ( .B1(n9996), .B2(n9995), .A(n9994), .ZN(ADD_1071_U47) );
  XOR2_X1 U11017 ( .A(n9998), .B(n9997), .Z(ADD_1071_U54) );
  XNOR2_X1 U11018 ( .A(n10000), .B(n9999), .ZN(ADD_1071_U49) );
  XOR2_X1 U11019 ( .A(n10002), .B(n10001), .Z(ADD_1071_U53) );
  XNOR2_X1 U11020 ( .A(n10004), .B(n10003), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4772 ( .A(n5663), .Z(n7779) );
  CLKBUF_X1 U4773 ( .A(n5443), .Z(n5532) );
  INV_X2 U4779 ( .A(n6153), .ZN(n6098) );
  CLKBUF_X1 U4804 ( .A(n7686), .Z(n4355) );
  CLKBUF_X1 U4820 ( .A(n9148), .Z(n4265) );
endmodule

