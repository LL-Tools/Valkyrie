

module b17_C_gen_AntiSAT_k_128_1 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput_f0, keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, 
        keyinput_f5, keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, 
        keyinput_f10, keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, 
        keyinput_f15, keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, 
        keyinput_f20, keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, 
        keyinput_f25, keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, 
        keyinput_f30, keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, 
        keyinput_f35, keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, 
        keyinput_f40, keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, 
        keyinput_f45, keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, 
        keyinput_f50, keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, 
        keyinput_f55, keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, 
        keyinput_f60, keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, 
        keyinput_g1, keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, 
        keyinput_g6, keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, 
        keyinput_g11, keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, 
        keyinput_g16, keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, 
        keyinput_g21, keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, 
        keyinput_g26, keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, 
        keyinput_g31, keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, 
        keyinput_g36, keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, 
        keyinput_g41, keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, 
        keyinput_g46, keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, 
        keyinput_g51, keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, 
        keyinput_g56, keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, 
        keyinput_g61, keyinput_g62, keyinput_g63, U355, U356, U357, U358, U359, 
        U360, U361, U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, 
        U373, U374, U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, 
        U376, U247, U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, 
        U236, U235, U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, 
        U224, U223, U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, 
        U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, 
        U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, 
        U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274, 
        P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, 
        P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, 
        P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, 
        P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, 
        P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, 
        P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, 
        P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, 
        P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, 
        P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, 
        P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, 
        P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, 
        P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, 
        P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, 
        P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, 
        P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, 
        P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, 
        P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, 
        P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, 
        P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, 
        P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, 
        P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, 
        P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, 
        P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, 
        P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, 
        P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, 
        P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, 
        P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, 
        P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, 
        P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, 
        P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, 
        P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, 
        P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, 
        P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, 
        P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, 
        P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, 
        P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, 
        P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, 
        P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, 
        P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, 
        P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, 
        P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, 
        P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, 
        P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, 
        P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, 
        P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, 
        P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, 
        P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, 
        P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, 
        P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, 
        P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, 
        P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, 
        P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, 
        P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, 
        P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, 
        P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, 
        P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, 
        P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, 
        P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, 
        P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, 
        P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, 
        P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, 
        P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, 
        P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, 
        P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, 
        P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, 
        P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, 
        P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, 
        P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, 
        P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, 
        P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, 
        P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, 
        P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, 
        P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, 
        P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, 
        P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, 
        P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, 
        P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, 
        P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, 
        P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, 
        P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, 
        P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, 
        P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, 
        P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, 
        P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, 
        P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, 
        P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, 
        P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, 
        P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, 
        P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, 
        P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, 
        P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, 
        P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, 
        P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, 
        P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, 
        P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, 
        P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, 
        P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, 
        P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, 
        P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, 
        P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, 
        P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, 
        P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, 
        P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, 
        P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, 
        P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, 
        P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, 
        P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, 
        P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, 
        P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, 
        P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, 
        P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, 
        P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, 
        P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, 
        P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, 
        P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, 
        P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, 
        P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, 
        P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, 
        P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, 
        P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, 
        P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, 
        P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, 
        P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, 
        P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, 
        P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, 
        P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, 
        P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, 
        P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, 
        P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, 
        P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, 
        P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, 
        P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, 
        P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, 
        P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, 
        P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, 
        P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, 
        P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, 
        P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, 
        P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, 
        P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, 
        P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, 
        P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, 
        P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, 
        P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, 
        P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, 
        P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, 
        P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, 
        P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, 
        P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, 
        P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, 
        P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, 
        P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, 
        P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, 
        P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, 
        P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, 
        P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, 
        P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, 
        P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, 
        P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, 
        P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, 
        P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, 
        P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, 
        P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, 
        P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, 
        P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, 
        P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, 
        P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, 
        P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, 
        P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, 
        P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, 
        P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, 
        P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, 
        P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, 
        P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, 
        P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, 
        P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, 
        P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, 
        P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, 
        P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, 
        P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, 
        P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9636, n9638, n9639, n9640, n9641, n9642, n9643, n9645, n9647, n9648,
         n9649, n9651, n9652, n9653, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
         n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
         n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
         n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,
         n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778,
         n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
         n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,
         n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802,
         n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810,
         n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818,
         n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
         n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834,
         n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842,
         n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850,
         n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
         n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
         n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874,
         n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882,
         n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890,
         n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
         n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906,
         n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914,
         n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922,
         n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,
         n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938,
         n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
         n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,
         n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962,
         n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,
         n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978,
         n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986,
         n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,
         n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
         n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,
         n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
         n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
         n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034,
         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
         n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
         n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058,
         n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
         n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
         n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
         n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
         n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106,
         n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,
         n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
         n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,
         n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
         n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
         n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154,
         n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
         n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,
         n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178,
         n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186,
         n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194,
         n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202,
         n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
         n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218,
         n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226,
         n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
         n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
         n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,
         n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258,
         n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266,
         n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,
         n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
         n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
         n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,
         n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
         n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,
         n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322,
         n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,
         n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
         n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,
         n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
         n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
         n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,
         n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
         n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394,
         n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
         n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
         n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
         n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
         n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
         n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
         n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
         n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458,
         n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,
         n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
         n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
         n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
         n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,
         n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
         n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
         n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,
         n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
         n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
         n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
         n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
         n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602,
         n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610,
         n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
         n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
         n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,
         n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
         n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
         n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,
         n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
         n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674,
         n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682,
         n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,
         n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
         n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706,
         n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,
         n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,
         n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730,
         n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
         n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746,
         n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754,
         n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762,
         n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770,
         n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778,
         n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,
         n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
         n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
         n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
         n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818,
         n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826,
         n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,
         n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,
         n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850,
         n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
         n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866,
         n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874,
         n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
         n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,
         n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,
         n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906,
         n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914,
         n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922,
         n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
         n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,
         n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,
         n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
         n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,
         n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970,
         n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978,
         n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
         n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
         n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
         n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
         n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,
         n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
         n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
         n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,
         n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,
         n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058,
         n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
         n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,
         n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
         n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
         n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
         n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106,
         n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114,
         n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,
         n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
         n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,
         n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
         n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
         n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,
         n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
         n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
         n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
         n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250,
         n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258,
         n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,
         n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
         n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
         n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290,
         n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
         n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306,
         n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314,
         n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322,
         n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330,
         n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338,
         n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
         n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
         n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362,
         n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
         n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378,
         n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,
         n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394,
         n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402,
         n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410,
         n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
         n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,
         n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434,
         n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
         n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450,
         n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458,
         n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466,
         n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474,
         n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482,
         n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490,
         n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498,
         n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506,
         n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,
         n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522,
         n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
         n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538,
         n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,
         n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,
         n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
         n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,
         n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578,
         n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,
         n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594,
         n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602,
         n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610,
         n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618,
         n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626,
         n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634,
         n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642,
         n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650,
         n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658,
         n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666,
         n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674,
         n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682,
         n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690,
         n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698,
         n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,
         n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714,
         n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722,
         n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,
         n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738,
         n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746,
         n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754,
         n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762,
         n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,
         n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778,
         n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786,
         n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794,
         n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
         n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810,
         n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818,
         n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826,
         n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834,
         n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842,
         n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850,
         n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858,
         n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866,
         n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874,
         n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882,
         n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890,
         n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898,
         n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906,
         n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914,
         n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922,
         n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930,
         n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938,
         n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946,
         n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954,
         n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962,
         n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970,
         n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978,
         n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986,
         n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994,
         n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002,
         n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010,
         n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018,
         n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026,
         n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034,
         n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042,
         n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050,
         n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058,
         n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066,
         n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074,
         n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082,
         n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090,
         n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098,
         n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106,
         n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114,
         n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122,
         n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130,
         n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138,
         n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146,
         n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154,
         n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162,
         n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170,
         n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178,
         n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186,
         n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194,
         n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202,
         n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210,
         n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218,
         n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226,
         n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234,
         n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242,
         n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250,
         n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258,
         n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266,
         n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274,
         n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282,
         n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290,
         n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298,
         n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306,
         n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314,
         n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322,
         n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330,
         n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338,
         n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346,
         n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354,
         n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362,
         n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370,
         n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378,
         n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386,
         n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394,
         n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402,
         n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410,
         n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418,
         n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426,
         n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434,
         n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442,
         n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450,
         n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458,
         n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466,
         n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474,
         n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482,
         n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490,
         n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498,
         n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506,
         n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514,
         n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522,
         n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530,
         n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538,
         n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546,
         n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554,
         n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562,
         n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570,
         n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578,
         n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586,
         n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594,
         n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602,
         n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610,
         n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618,
         n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626,
         n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634,
         n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642,
         n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650,
         n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658,
         n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666,
         n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674,
         n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682,
         n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690,
         n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698,
         n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706,
         n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714,
         n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722,
         n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730,
         n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738,
         n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746,
         n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754,
         n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762,
         n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770,
         n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778,
         n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786,
         n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794,
         n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802,
         n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810,
         n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818,
         n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826,
         n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834,
         n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842,
         n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850,
         n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858,
         n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866,
         n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874,
         n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
         n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890,
         n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898,
         n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906,
         n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914,
         n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922,
         n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930,
         n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938,
         n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946,
         n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954,
         n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962,
         n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970,
         n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978,
         n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986,
         n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994,
         n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002,
         n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010,
         n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018,
         n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026,
         n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034,
         n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042,
         n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050,
         n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058,
         n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066,
         n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
         n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082,
         n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090,
         n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098,
         n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106,
         n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114,
         n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122,
         n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130,
         n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
         n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
         n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154,
         n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162,
         n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170,
         n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178,
         n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186,
         n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194,
         n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202,
         n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210,
         n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218,
         n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226,
         n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234,
         n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242,
         n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250,
         n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258,
         n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266,
         n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274,
         n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282,
         n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290,
         n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298,
         n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306,
         n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314,
         n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322,
         n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330,
         n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338,
         n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346,
         n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354,
         n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362,
         n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370,
         n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378,
         n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386,
         n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394,
         n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402,
         n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410,
         n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418,
         n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426,
         n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
         n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442,
         n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450,
         n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458,
         n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466,
         n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474,
         n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482,
         n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490,
         n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498,
         n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506,
         n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514,
         n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522,
         n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530,
         n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538,
         n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546,
         n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554,
         n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562,
         n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570,
         n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578,
         n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586,
         n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594,
         n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
         n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610,
         n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618,
         n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626,
         n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634,
         n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642,
         n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650,
         n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658,
         n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666,
         n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674,
         n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682,
         n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690,
         n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698,
         n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706,
         n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714,
         n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
         n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730,
         n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738,
         n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746,
         n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754,
         n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762,
         n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770,
         n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778,
         n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786,
         n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
         n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802,
         n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810,
         n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818,
         n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826,
         n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834,
         n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842,
         n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850,
         n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858,
         n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
         n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874,
         n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882,
         n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890,
         n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898,
         n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906,
         n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914,
         n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922,
         n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
         n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
         n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946,
         n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954,
         n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962,
         n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970,
         n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978,
         n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986,
         n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994,
         n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002,
         n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010,
         n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018,
         n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026,
         n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034,
         n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042,
         n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050,
         n21051, n21052, n21053, n21054;

  OAI21_X2 U11080 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19130), .A(n16787), 
        .ZN(n18144) );
  OR2_X1 U11081 ( .A1(n10019), .A2(n12436), .ZN(n19528) );
  NAND2_X1 U11082 ( .A1(n12452), .A2(n12423), .ZN(n19830) );
  NAND2_X1 U11083 ( .A1(n11270), .A2(n11269), .ZN(n11962) );
  CLKBUF_X2 U11084 ( .A(n15894), .Z(n15864) );
  BUF_X1 U11085 ( .A(n17211), .Z(n9657) );
  CLKBUF_X2 U11086 ( .A(n10654), .Z(n10774) );
  BUF_X2 U11087 ( .A(n10631), .Z(n12727) );
  CLKBUF_X2 U11088 ( .A(n10659), .Z(n10775) );
  CLKBUF_X2 U11089 ( .A(n13964), .Z(n17433) );
  CLKBUF_X2 U11090 ( .A(n13948), .Z(n17432) );
  CLKBUF_X2 U11091 ( .A(n15940), .Z(n17380) );
  CLKBUF_X2 U11092 ( .A(n11117), .Z(n11754) );
  CLKBUF_X1 U11093 ( .A(n11805), .Z(n9645) );
  AND2_X1 U11094 ( .A1(n10371), .A2(n10489), .ZN(n12150) );
  AND2_X1 U11095 ( .A1(n10371), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12088) );
  AND2_X1 U11096 ( .A1(n9641), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12087) );
  CLKBUF_X1 U11097 ( .A(n15894), .Z(n17450) );
  AND2_X1 U11098 ( .A1(n12337), .A2(n10648), .ZN(n12767) );
  INV_X1 U11099 ( .A(n13129), .ZN(n14166) );
  CLKBUF_X2 U11100 ( .A(n11055), .Z(n11775) );
  CLKBUF_X1 U11101 ( .A(n10615), .Z(n19486) );
  BUF_X2 U11105 ( .A(n11227), .Z(n9647) );
  AND2_X1 U11107 ( .A1(n11014), .A2(n11015), .ZN(n11117) );
  AND2_X2 U11108 ( .A1(n13333), .A2(n11009), .ZN(n11050) );
  NOR2_X2 U11109 ( .A1(n18512), .A2(n17653), .ZN(n17603) );
  OAI21_X1 U11110 ( .B1(n16124), .B2(n16123), .A(n19131), .ZN(n17653) );
  INV_X1 U11111 ( .A(n19981), .ZN(n9636) );
  INV_X1 U11113 ( .A(n9636), .ZN(n9638) );
  CLKBUF_X2 U11114 ( .A(n11198), .Z(n9648) );
  CLKBUF_X2 U11115 ( .A(n11586), .Z(n11776) );
  OR2_X1 U11116 ( .A1(n10774), .A2(n12785), .ZN(n10687) );
  AND2_X1 U11117 ( .A1(n9642), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10516) );
  AND2_X1 U11118 ( .A1(n10687), .A2(n10686), .ZN(n10691) );
  AND4_X1 U11119 ( .A1(n10233), .A2(n10234), .A3(n12555), .A4(n9791), .ZN(
        n10031) );
  OR2_X1 U11120 ( .A1(n10019), .A2(n12444), .ZN(n19494) );
  AND2_X1 U11121 ( .A1(n9890), .A2(n9738), .ZN(n16016) );
  INV_X1 U11122 ( .A(n10659), .ZN(n10680) );
  OR2_X1 U11123 ( .A1(n15014), .A2(n10243), .ZN(n9834) );
  AND2_X1 U11124 ( .A1(n12287), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10811) );
  INV_X1 U11125 ( .A(n12495), .ZN(n12843) );
  CLKBUF_X3 U11127 ( .A(n10617), .Z(n12755) );
  CLKBUF_X2 U11129 ( .A(n15911), .Z(n9655) );
  INV_X1 U11131 ( .A(n13660), .ZN(n9900) );
  AOI21_X1 U11132 ( .B1(n14979), .B2(n14973), .A(n12293), .ZN(n14967) );
  CLKBUF_X3 U11133 ( .A(n10601), .Z(n12012) );
  INV_X1 U11134 ( .A(n19136), .ZN(n16806) );
  NAND2_X1 U11135 ( .A1(n13308), .A2(n9713), .ZN(n13446) );
  XNOR2_X1 U11136 ( .A(n12559), .B(n15660), .ZN(n15416) );
  INV_X1 U11137 ( .A(n17661), .ZN(n18482) );
  INV_X1 U11138 ( .A(n18144), .ZN(n18101) );
  INV_X1 U11139 ( .A(n15709), .ZN(n15707) );
  INV_X1 U11140 ( .A(n20197), .ZN(n20189) );
  XNOR2_X1 U11141 ( .A(n11990), .B(n11827), .ZN(n14186) );
  NAND2_X2 U11142 ( .A1(n13536), .A2(n13522), .ZN(n12307) );
  AND2_X2 U11143 ( .A1(n11014), .A2(n13344), .ZN(n11055) );
  NAND2_X2 U11144 ( .A1(n12685), .A2(n12684), .ZN(n15319) );
  NAND2_X2 U11145 ( .A1(n10122), .A2(n11867), .ZN(n13722) );
  NOR2_X2 U11146 ( .A1(n17799), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17798) );
  INV_X2 U11147 ( .A(n12771), .ZN(n10640) );
  NAND2_X2 U11148 ( .A1(n12952), .A2(n13482), .ZN(n12377) );
  AND2_X4 U11149 ( .A1(n11009), .A2(n11015), .ZN(n9672) );
  INV_X1 U11150 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9639) );
  NOR2_X1 U11151 ( .A1(n11828), .A2(n11141), .ZN(n13329) );
  AOI211_X2 U11152 ( .C1(n16204), .C2(n14555), .A(n14554), .B(n14553), .ZN(
        n14556) );
  NAND2_X2 U11153 ( .A1(n19115), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13939) );
  AND2_X2 U11154 ( .A1(n12001), .A2(n10262), .ZN(n11990) );
  NAND2_X2 U11155 ( .A1(n10630), .A2(n10235), .ZN(n12340) );
  AND2_X2 U11156 ( .A1(n10640), .A2(n10639), .ZN(n10630) );
  INV_X4 U11157 ( .A(n13959), .ZN(n17447) );
  INV_X2 U11158 ( .A(n11352), .ZN(n9951) );
  NAND2_X2 U11159 ( .A1(n10144), .A2(n10143), .ZN(n11352) );
  AND2_X4 U11160 ( .A1(n12741), .A2(n10352), .ZN(n10372) );
  AND4_X2 U11161 ( .A1(n11027), .A2(n11026), .A3(n11025), .A4(n11024), .ZN(
        n11028) );
  AND4_X2 U11162 ( .A1(n11066), .A2(n11065), .A3(n11064), .A4(n11063), .ZN(
        n9737) );
  INV_X2 U11163 ( .A(n12307), .ZN(n9640) );
  INV_X2 U11164 ( .A(n12307), .ZN(n9641) );
  NOR4_X4 U11165 ( .A1(n17653), .A2(n17595), .A3(n17596), .A4(n17506), .ZN(
        n17594) );
  BUF_X4 U11166 ( .A(n10824), .Z(n10994) );
  AOI21_X2 U11167 ( .B1(n20106), .B2(n10642), .A(n12755), .ZN(n12410) );
  OR2_X4 U11168 ( .A1(n13888), .A2(n11903), .ZN(n14626) );
  INV_X1 U11169 ( .A(n12266), .ZN(n9642) );
  INV_X1 U11170 ( .A(n12266), .ZN(n9643) );
  AND2_X4 U11171 ( .A1(n11005), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13333) );
  AOI221_X2 U11172 ( .B1(n18217), .B2(n18931), .C1(n18246), .C2(n18931), .A(
        n18207), .ZN(n18225) );
  INV_X2 U11173 ( .A(n20115), .ZN(n12733) );
  NAND2_X4 U11174 ( .A1(n10454), .A2(n10453), .ZN(n20115) );
  OAI21_X1 U11176 ( .B1(n14525), .B2(n11916), .A(n16174), .ZN(n14517) );
  INV_X1 U11177 ( .A(n12373), .ZN(n11144) );
  NOR3_X2 U11178 ( .A1(n14231), .A2(n20887), .A3(n21005), .ZN(n14210) );
  BUF_X4 U11179 ( .A(n11198), .Z(n9682) );
  NAND2_X2 U11181 ( .A1(n11029), .A2(n11028), .ZN(n11133) );
  AND2_X2 U11182 ( .A1(n13346), .A2(n13344), .ZN(n11227) );
  AND2_X1 U11183 ( .A1(n13346), .A2(n13330), .ZN(n11670) );
  NOR3_X1 U11184 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n18944), .ZN(n9649) );
  NOR3_X1 U11185 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n18944), .ZN(n13948) );
  NOR2_X2 U11187 ( .A1(n18044), .A2(n9856), .ZN(n17906) );
  OR2_X1 U11188 ( .A1(n10111), .A2(n15255), .ZN(n15270) );
  AND3_X1 U11189 ( .A1(n10110), .A2(n10109), .A3(n15256), .ZN(n15463) );
  AND4_X1 U11190 ( .A1(n12703), .A2(n15279), .A3(n12702), .A4(n10231), .ZN(
        n15255) );
  CLKBUF_X1 U11191 ( .A(n14979), .Z(n14980) );
  INV_X1 U11192 ( .A(n15345), .ZN(n9653) );
  AND2_X1 U11193 ( .A1(n9916), .A2(n9914), .ZN(n9752) );
  NOR3_X1 U11194 ( .A1(n14604), .A2(n10088), .A3(n11909), .ZN(n9947) );
  NAND2_X1 U11195 ( .A1(n12558), .A2(n14909), .ZN(n12559) );
  OR2_X1 U11196 ( .A1(n15156), .A2(n15155), .ZN(n15158) );
  AND2_X1 U11197 ( .A1(n10014), .A2(n10013), .ZN(n17789) );
  AND2_X1 U11198 ( .A1(n12803), .A2(n12849), .ZN(n15545) );
  OR2_X1 U11199 ( .A1(n14628), .A2(n16273), .ZN(n11906) );
  NAND2_X1 U11200 ( .A1(n13367), .A2(n13369), .ZN(n13368) );
  AOI22_X1 U11201 ( .A1(n18132), .A2(n18329), .B1(n18012), .B2(n18331), .ZN(
        n18044) );
  NAND2_X1 U11202 ( .A1(n10028), .A2(n12424), .ZN(n15728) );
  CLKBUF_X2 U11203 ( .A(n13359), .Z(n9673) );
  NAND2_X1 U11204 ( .A1(n10028), .A2(n12423), .ZN(n19732) );
  OR2_X2 U11205 ( .A1(n12445), .A2(n12444), .ZN(n12531) );
  OR2_X1 U11206 ( .A1(n20848), .A2(n13647), .ZN(n13734) );
  NAND2_X1 U11207 ( .A1(n13034), .A2(n13033), .ZN(n13035) );
  NOR2_X1 U11208 ( .A1(n18921), .A2(n18459), .ZN(n18463) );
  NOR2_X1 U11209 ( .A1(n18096), .A2(n18097), .ZN(n18095) );
  NOR2_X1 U11210 ( .A1(n18110), .A2(n16002), .ZN(n16005) );
  AND3_X1 U11211 ( .A1(n10611), .A2(n12346), .A3(n10610), .ZN(n12409) );
  NOR2_X1 U11212 ( .A1(n18123), .A2(n18124), .ZN(n15999) );
  XNOR2_X1 U11214 ( .A(n15994), .B(n18436), .ZN(n18124) );
  CLKBUF_X2 U11215 ( .A(n10605), .Z(n10508) );
  INV_X2 U11216 ( .A(n10601), .ZN(n10606) );
  BUF_X2 U11217 ( .A(n11215), .Z(n11800) );
  BUF_X1 U11218 ( .A(n15912), .Z(n17448) );
  CLKBUF_X2 U11219 ( .A(n9672), .Z(n11638) );
  CLKBUF_X2 U11220 ( .A(n11072), .Z(n11782) );
  CLKBUF_X3 U11221 ( .A(n15756), .Z(n9656) );
  BUF_X2 U11222 ( .A(n11073), .Z(n11091) );
  INV_X4 U11224 ( .A(n10487), .ZN(n12308) );
  CLKBUF_X1 U11225 ( .A(n11227), .Z(n9674) );
  BUF_X2 U11226 ( .A(n11197), .Z(n11783) );
  CLKBUF_X3 U11227 ( .A(n15913), .Z(n9658) );
  NOR2_X1 U11229 ( .A1(n17178), .A2(n13940), .ZN(n13964) );
  NOR2_X1 U11230 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13938), .ZN(
        n17211) );
  CLKBUF_X2 U11231 ( .A(n10487), .Z(n12282) );
  INV_X2 U11232 ( .A(n18447), .ZN(n9652) );
  AND2_X2 U11233 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12741) );
  NAND2_X1 U11234 ( .A1(n15270), .A2(n15453), .ZN(n15450) );
  AOI21_X1 U11235 ( .B1(n12877), .B2(n16205), .A(n9785), .ZN(n10130) );
  NAND2_X1 U11236 ( .A1(n14517), .A2(n11998), .ZN(n11999) );
  AOI211_X1 U11237 ( .C1(n14546), .C2(n16205), .A(n14545), .B(n14544), .ZN(
        n14547) );
  AOI21_X1 U11238 ( .B1(n14200), .B2(n11991), .A(n11990), .ZN(n14387) );
  OR2_X1 U11239 ( .A1(n15282), .A2(n15281), .ZN(n15473) );
  NAND2_X1 U11240 ( .A1(n12723), .A2(n9956), .ZN(n15247) );
  AND2_X1 U11241 ( .A1(n14101), .A2(n14100), .ZN(n14102) );
  AND2_X1 U11242 ( .A1(n14112), .A2(n14111), .ZN(n14113) );
  NAND2_X1 U11243 ( .A1(n11914), .A2(n16174), .ZN(n14557) );
  NAND2_X1 U11244 ( .A1(n9945), .A2(n9944), .ZN(n11914) );
  OAI21_X1 U11245 ( .B1(n15443), .B2(n15442), .A(n15441), .ZN(n15444) );
  AND2_X1 U11246 ( .A1(n9846), .A2(n9845), .ZN(n15443) );
  AND2_X2 U11247 ( .A1(n10226), .A2(n10224), .ZN(n10072) );
  NAND2_X1 U11248 ( .A1(n16102), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16613) );
  OR2_X1 U11249 ( .A1(n16045), .A2(n16651), .ZN(n10167) );
  NAND2_X1 U11250 ( .A1(n12599), .A2(n9697), .ZN(n10226) );
  NAND2_X1 U11251 ( .A1(n16043), .A2(n16042), .ZN(n16044) );
  NOR2_X1 U11252 ( .A1(n17780), .A2(n17779), .ZN(n17778) );
  OR2_X1 U11253 ( .A1(n14759), .A2(n14756), .ZN(n11910) );
  AOI21_X1 U11254 ( .B1(n17791), .B2(n17952), .A(n17789), .ZN(n17779) );
  NAND2_X1 U11255 ( .A1(n9864), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17791) );
  AND2_X1 U11256 ( .A1(n13747), .A2(n9788), .ZN(n9903) );
  OR2_X1 U11257 ( .A1(n11892), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16197) );
  NOR2_X1 U11258 ( .A1(n17818), .A2(n18158), .ZN(n18155) );
  OR2_X1 U11259 ( .A1(n10031), .A2(n12838), .ZN(n10030) );
  NOR2_X1 U11260 ( .A1(n10222), .A2(n9963), .ZN(n9962) );
  INV_X1 U11261 ( .A(n12493), .ZN(n10234) );
  AND2_X1 U11262 ( .A1(n14858), .A2(n10192), .ZN(n15224) );
  NAND2_X1 U11263 ( .A1(n11343), .A2(n11342), .ZN(n13147) );
  NOR2_X1 U11264 ( .A1(n14372), .A2(n13764), .ZN(n20190) );
  NAND2_X1 U11265 ( .A1(n17888), .A2(n17874), .ZN(n17915) );
  NOR2_X1 U11266 ( .A1(n17725), .A2(n17531), .ZN(n17527) );
  NOR2_X1 U11267 ( .A1(n13661), .A2(n13662), .ZN(n13763) );
  CLKBUF_X1 U11268 ( .A(n12402), .Z(n14491) );
  NAND2_X1 U11269 ( .A1(n11265), .A2(n11264), .ZN(n11331) );
  NAND2_X1 U11270 ( .A1(n12633), .A2(n12686), .ZN(n12694) );
  OR2_X1 U11271 ( .A1(n13136), .A2(n13137), .ZN(n13138) );
  AOI21_X1 U11272 ( .B1(n16034), .B2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n9857), .ZN(n17927) );
  AND2_X1 U11273 ( .A1(n11282), .A2(n11281), .ZN(n13390) );
  OR2_X1 U11274 ( .A1(n17719), .A2(n17540), .ZN(n17541) );
  OR2_X1 U11275 ( .A1(n12047), .A2(n12046), .ZN(n10272) );
  OR2_X1 U11276 ( .A1(n13181), .A2(n10199), .ZN(n16527) );
  INV_X1 U11277 ( .A(n12439), .ZN(n10028) );
  AND2_X1 U11278 ( .A1(n13044), .A2(n12044), .ZN(n13159) );
  XNOR2_X1 U11279 ( .A(n11207), .B(n11206), .ZN(n11332) );
  AND2_X1 U11280 ( .A1(n13049), .A2(n13048), .ZN(n13051) );
  NAND2_X1 U11281 ( .A1(n12028), .A2(n12027), .ZN(n12045) );
  NOR2_X1 U11282 ( .A1(n12853), .A2(n13563), .ZN(n15567) );
  OR2_X1 U11283 ( .A1(n12853), .A2(n12783), .ZN(n15569) );
  AND2_X1 U11284 ( .A1(n9895), .A2(n9891), .ZN(n11207) );
  OR2_X1 U11285 ( .A1(n12645), .A2(n10590), .ZN(n12659) );
  OR2_X1 U11286 ( .A1(n13059), .A2(n16591), .ZN(n12450) );
  NAND2_X1 U11287 ( .A1(n12764), .A2(n13010), .ZN(n12853) );
  NAND2_X1 U11288 ( .A1(n13109), .A2(n12991), .ZN(n20848) );
  AND2_X1 U11289 ( .A1(n9893), .A2(n9892), .ZN(n9891) );
  XNOR2_X1 U11290 ( .A(n11263), .B(n11261), .ZN(n11339) );
  NOR2_X1 U11291 ( .A1(n15709), .A2(n15708), .ZN(n19479) );
  XNOR2_X1 U11292 ( .A(n11344), .B(n10085), .ZN(n13419) );
  NAND2_X1 U11293 ( .A1(n10083), .A2(n11235), .ZN(n11344) );
  OAI21_X1 U11294 ( .B1(n19322), .B2(n12859), .A(n12041), .ZN(n15684) );
  NAND2_X1 U11295 ( .A1(n11240), .A2(n11893), .ZN(n11263) );
  NAND2_X1 U11296 ( .A1(n11257), .A2(n11256), .ZN(n20325) );
  AND2_X1 U11297 ( .A1(n9695), .A2(n18380), .ZN(n10012) );
  OR2_X1 U11298 ( .A1(n18067), .A2(n18373), .ZN(n10154) );
  INV_X1 U11299 ( .A(n12422), .ZN(n12418) );
  NOR2_X2 U11300 ( .A1(n16806), .A2(n16787), .ZN(n18132) );
  NOR2_X1 U11301 ( .A1(n12601), .A2(n10118), .ZN(n12617) );
  NAND2_X1 U11302 ( .A1(n11268), .A2(n11267), .ZN(n13470) );
  NAND2_X1 U11303 ( .A1(n11189), .A2(n11188), .ZN(n11190) );
  NOR2_X1 U11304 ( .A1(n18072), .A2(n15979), .ZN(n15981) );
  OR2_X1 U11305 ( .A1(n12601), .A2(n12727), .ZN(n12706) );
  NOR2_X1 U11306 ( .A1(n18074), .A2(n18073), .ZN(n18072) );
  AOI21_X1 U11307 ( .B1(n10780), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n10682), .ZN(n12022) );
  NAND2_X1 U11308 ( .A1(n9851), .A2(n9747), .ZN(n15682) );
  NAND2_X1 U11309 ( .A1(n12605), .A2(n12603), .ZN(n12601) );
  CLKBUF_X1 U11310 ( .A(n11165), .Z(n11166) );
  INV_X2 U11311 ( .A(n10614), .ZN(n10780) );
  NOR2_X1 U11312 ( .A1(n12593), .A2(n12592), .ZN(n12605) );
  INV_X1 U11313 ( .A(n18914), .ZN(n18943) );
  NAND2_X1 U11314 ( .A1(n11146), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11165) );
  NOR2_X2 U11315 ( .A1(n18265), .A2(n18951), .ZN(n18267) );
  NAND2_X1 U11316 ( .A1(n18953), .A2(n18949), .ZN(n18265) );
  NOR2_X1 U11317 ( .A1(n18113), .A2(n15972), .ZN(n18100) );
  NAND2_X1 U11318 ( .A1(n10653), .A2(n10649), .ZN(n10676) );
  NOR2_X1 U11319 ( .A1(n12511), .A2(n12512), .ZN(n12557) );
  XNOR2_X1 U11320 ( .A(n16005), .B(n16006), .ZN(n18096) );
  AND2_X1 U11321 ( .A1(n10645), .A2(n10644), .ZN(n10653) );
  OAI21_X1 U11322 ( .B1(n9841), .B2(n12331), .A(n12738), .ZN(n9840) );
  NOR2_X2 U11323 ( .A1(n18929), .A2(n15987), .ZN(n18953) );
  OAI21_X1 U11324 ( .B1(n12963), .B2(n10822), .A(n10821), .ZN(n13496) );
  NAND2_X1 U11325 ( .A1(n14034), .A2(n18915), .ZN(n15987) );
  AND2_X1 U11326 ( .A1(n11151), .A2(n11150), .ZN(n13076) );
  AOI21_X1 U11327 ( .B1(n12767), .B2(n12771), .A(n10616), .ZN(n10661) );
  NOR2_X1 U11328 ( .A1(n14046), .A2(n14054), .ZN(n18915) );
  NAND2_X2 U11329 ( .A1(n19136), .A2(n17701), .ZN(n17767) );
  AOI21_X1 U11330 ( .B1(n11235), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n10085), 
        .ZN(n10084) );
  INV_X1 U11331 ( .A(n11378), .ZN(n11379) );
  AOI21_X1 U11332 ( .B1(n13070), .B2(n14788), .A(n11156), .ZN(n11174) );
  NOR2_X1 U11333 ( .A1(n19136), .A2(n17700), .ZN(n14054) );
  MUX2_X1 U11334 ( .A(n12745), .B(n14944), .S(n12727), .Z(n12508) );
  OR2_X1 U11335 ( .A1(n12816), .A2(n20122), .ZN(n12963) );
  NOR4_X1 U11336 ( .A1(n18482), .A2(n14047), .A3(n14032), .A4(n17511), .ZN(
        n18976) );
  CLKBUF_X1 U11337 ( .A(n11176), .Z(n13649) );
  NAND2_X1 U11338 ( .A1(n13482), .A2(n13660), .ZN(n13656) );
  AND4_X2 U11339 ( .A1(n12727), .A2(n13571), .A3(n19486), .A4(n20089), .ZN(
        n10998) );
  INV_X1 U11340 ( .A(n10608), .ZN(n20103) );
  CLKBUF_X1 U11341 ( .A(n13129), .Z(n14188) );
  AND2_X1 U11342 ( .A1(n20115), .A2(n13571), .ZN(n12329) );
  AND3_X1 U11343 ( .A1(n12413), .A2(n10631), .A3(n9741), .ZN(n12775) );
  NOR2_X1 U11344 ( .A1(n10643), .A2(n15751), .ZN(n10665) );
  AND4_X1 U11345 ( .A1(n10601), .A2(n10615), .A3(n10647), .A4(n10605), .ZN(
        n10639) );
  INV_X2 U11346 ( .A(n20116), .ZN(n15751) );
  INV_X1 U11347 ( .A(n20116), .ZN(n13571) );
  INV_X1 U11348 ( .A(n10615), .ZN(n12413) );
  AND2_X2 U11349 ( .A1(n10479), .A2(n10478), .ZN(n20116) );
  CLKBUF_X2 U11350 ( .A(n10455), .Z(n19459) );
  INV_X2 U11351 ( .A(n13658), .ZN(n9666) );
  INV_X1 U11352 ( .A(n13658), .ZN(n9665) );
  AND2_X2 U11353 ( .A1(n10430), .A2(n10429), .ZN(n12771) );
  INV_X1 U11354 ( .A(n10455), .ZN(n12777) );
  NAND4_X2 U11355 ( .A1(n9997), .A2(n15965), .A3(n9723), .A4(n15963), .ZN(
        n18142) );
  CLKBUF_X1 U11356 ( .A(n11170), .Z(n13689) );
  CLKBUF_X1 U11357 ( .A(n11143), .Z(n13212) );
  OR2_X1 U11358 ( .A1(n10507), .A2(n10506), .ZN(n12815) );
  OR2_X1 U11359 ( .A1(n10522), .A2(n10521), .ZN(n12490) );
  NAND2_X1 U11360 ( .A1(n10273), .A2(n15925), .ZN(n17654) );
  INV_X2 U11361 ( .A(U212), .ZN(n16735) );
  OR2_X1 U11362 ( .A1(n10535), .A2(n10534), .ZN(n12827) );
  AND2_X1 U11363 ( .A1(n10003), .A2(n9998), .ZN(n9997) );
  NAND2_X1 U11364 ( .A1(n10440), .A2(n10441), .ZN(n10615) );
  NAND2_X1 U11365 ( .A1(n10370), .A2(n10369), .ZN(n10601) );
  NAND3_X1 U11366 ( .A1(n10283), .A2(n10452), .A3(n10451), .ZN(n10453) );
  NAND2_X2 U11367 ( .A1(n9737), .A2(n11071), .ZN(n11141) );
  OR2_X1 U11368 ( .A1(n11062), .A2(n11061), .ZN(n11306) );
  AND4_X1 U11369 ( .A1(n11095), .A2(n11094), .A3(n11093), .A4(n11092), .ZN(
        n11106) );
  NAND2_X1 U11370 ( .A1(n10447), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10454) );
  AND4_X1 U11371 ( .A1(n11129), .A2(n11128), .A3(n11127), .A4(n11126), .ZN(
        n13658) );
  INV_X1 U11372 ( .A(n10306), .ZN(n10301) );
  NAND2_X1 U11373 ( .A1(n9939), .A2(n9691), .ZN(n11134) );
  OR2_X2 U11374 ( .A1(n16736), .A2(n16680), .ZN(n16738) );
  AND4_X1 U11375 ( .A1(n10446), .A2(n10445), .A3(n10444), .A4(n10443), .ZN(
        n10447) );
  AND4_X1 U11376 ( .A1(n11099), .A2(n11098), .A3(n11097), .A4(n11096), .ZN(
        n11105) );
  AND4_X1 U11377 ( .A1(n11125), .A2(n11124), .A3(n11123), .A4(n11122), .ZN(
        n11126) );
  AND4_X1 U11378 ( .A1(n11121), .A2(n11120), .A3(n11119), .A4(n11118), .ZN(
        n11127) );
  AND4_X1 U11379 ( .A1(n11116), .A2(n11115), .A3(n11114), .A4(n11113), .ZN(
        n11128) );
  AND4_X1 U11380 ( .A1(n11090), .A2(n11089), .A3(n11088), .A4(n11087), .ZN(
        n11107) );
  AND4_X1 U11381 ( .A1(n11111), .A2(n11110), .A3(n11109), .A4(n11108), .ZN(
        n11129) );
  AND3_X1 U11382 ( .A1(n9740), .A2(n10286), .A3(n11037), .ZN(n11049) );
  AND4_X1 U11383 ( .A1(n11023), .A2(n11022), .A3(n11021), .A4(n11020), .ZN(
        n11029) );
  NAND2_X2 U11384 ( .A1(n20034), .A2(n19997), .ZN(n20043) );
  CLKBUF_X2 U11385 ( .A(n11050), .Z(n9681) );
  AND4_X1 U11386 ( .A1(n11103), .A2(n11102), .A3(n11101), .A4(n11100), .ZN(
        n11104) );
  CLKBUF_X1 U11387 ( .A(n10450), .Z(n12309) );
  AND2_X2 U11388 ( .A1(n10488), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10515) );
  AND2_X2 U11389 ( .A1(n10488), .A2(n10489), .ZN(n10514) );
  AND2_X2 U11390 ( .A1(n9671), .A2(n10489), .ZN(n10544) );
  INV_X4 U11391 ( .A(n15839), .ZN(n17212) );
  CLKBUF_X3 U11392 ( .A(n17455), .Z(n15860) );
  BUF_X2 U11393 ( .A(n13971), .Z(n17407) );
  INV_X1 U11394 ( .A(n20054), .ZN(n19981) );
  BUF_X4 U11395 ( .A(n11226), .Z(n11784) );
  BUF_X2 U11396 ( .A(n15912), .Z(n17334) );
  CLKBUF_X1 U11397 ( .A(n11226), .Z(n11806) );
  INV_X2 U11398 ( .A(n16772), .ZN(U215) );
  OR2_X1 U11399 ( .A1(n10465), .A2(n10464), .ZN(n10466) );
  OAI22_X1 U11400 ( .A1(n12132), .A2(n12464), .B1(n12275), .B2(n12471), .ZN(
        n10422) );
  OR2_X1 U11401 ( .A1(n10417), .A2(n10416), .ZN(n10418) );
  INV_X1 U11402 ( .A(n12266), .ZN(n9671) );
  INV_X2 U11403 ( .A(n16776), .ZN(n16778) );
  CLKBUF_X1 U11404 ( .A(n12266), .Z(n12275) );
  INV_X2 U11405 ( .A(n13974), .ZN(n9667) );
  INV_X4 U11406 ( .A(n12133), .ZN(n10488) );
  INV_X4 U11407 ( .A(n17150), .ZN(n17449) );
  INV_X2 U11408 ( .A(n20098), .ZN(n20034) );
  OR2_X1 U11409 ( .A1(n18944), .A2(n13940), .ZN(n15839) );
  AND2_X2 U11410 ( .A1(n13333), .A2(n13346), .ZN(n11078) );
  NOR2_X1 U11411 ( .A1(n19095), .A2(n17977), .ZN(n19133) );
  AND2_X2 U11412 ( .A1(n13333), .A2(n13083), .ZN(n11226) );
  AND2_X2 U11413 ( .A1(n13330), .A2(n11009), .ZN(n11586) );
  AND2_X1 U11414 ( .A1(n13083), .A2(n13330), .ZN(n11073) );
  AND2_X2 U11415 ( .A1(n11006), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11009) );
  NAND2_X1 U11416 ( .A1(n19115), .A2(n19108), .ZN(n17178) );
  AND2_X4 U11417 ( .A1(n11015), .A2(n13346), .ZN(n11197) );
  NAND3_X2 U11418 ( .A1(n19111), .A2(n18986), .A3(n18978), .ZN(n18447) );
  AND2_X2 U11419 ( .A1(n11007), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13330) );
  OR2_X1 U11420 ( .A1(n18944), .A2(n14035), .ZN(n17150) );
  NOR2_X2 U11421 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10351) );
  NOR2_X1 U11422 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10350) );
  INV_X1 U11423 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11007) );
  AND2_X1 U11424 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13521) );
  CLKBUF_X1 U11425 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n15690) );
  NAND2_X1 U11426 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18944) );
  AND2_X2 U11427 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13344) );
  INV_X1 U11428 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15754) );
  INV_X1 U11429 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12440) );
  INV_X1 U11430 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12437) );
  INV_X1 U11431 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12482) );
  INV_X1 U11432 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12441) );
  INV_X1 U11433 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12462) );
  NAND2_X1 U11434 ( .A1(n11874), .A2(n9662), .ZN(n9659) );
  AND2_X2 U11435 ( .A1(n9659), .A2(n9660), .ZN(n16195) );
  OR2_X1 U11436 ( .A1(n9661), .A2(n13835), .ZN(n9660) );
  INV_X1 U11437 ( .A(n11882), .ZN(n9661) );
  AND2_X1 U11438 ( .A1(n11873), .A2(n11882), .ZN(n9662) );
  NAND2_X1 U11439 ( .A1(n13425), .A2(n11255), .ZN(n9663) );
  NAND2_X1 U11440 ( .A1(n11282), .A2(n11281), .ZN(n9664) );
  NAND2_X1 U11441 ( .A1(n13425), .A2(n11255), .ZN(n11258) );
  NOR2_X1 U11442 ( .A1(n11999), .A2(n11918), .ZN(n14508) );
  CLKBUF_X1 U11443 ( .A(n11142), .Z(n14432) );
  NAND2_X1 U11445 ( .A1(n11142), .A2(n11134), .ZN(n12387) );
  INV_X1 U11446 ( .A(n11133), .ZN(n11142) );
  AOI21_X2 U11447 ( .B1(n11260), .B2(n20846), .A(n9784), .ZN(n11832) );
  INV_X1 U11448 ( .A(n12972), .ZN(n11085) );
  OR4_X1 U11449 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(n19115), .A4(n19092), .ZN(
        n13974) );
  AND2_X1 U11450 ( .A1(n13330), .A2(n11009), .ZN(n9668) );
  AND2_X1 U11451 ( .A1(n13083), .A2(n13330), .ZN(n9669) );
  INV_X1 U11452 ( .A(n11091), .ZN(n9670) );
  NOR2_X2 U11453 ( .A1(n15033), .A2(n15035), .ZN(n15029) );
  NAND2_X2 U11454 ( .A1(n11165), .A2(n11161), .ZN(n11184) );
  AND2_X2 U11455 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13083) );
  NAND2_X1 U11456 ( .A1(n14507), .A2(n11920), .ZN(n11995) );
  NAND2_X1 U11457 ( .A1(n11258), .A2(n11191), .ZN(n9899) );
  NOR2_X1 U11458 ( .A1(n13390), .A2(n9949), .ZN(n9948) );
  OR2_X1 U11459 ( .A1(n11263), .A2(n11262), .ZN(n11264) );
  XNOR2_X1 U11460 ( .A(n11852), .B(n13293), .ZN(n13284) );
  NAND2_X1 U11461 ( .A1(n11841), .A2(n11840), .ZN(n11852) );
  AND2_X4 U11462 ( .A1(n13536), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10371) );
  NAND2_X1 U11463 ( .A1(n9951), .A2(n9948), .ZN(n11377) );
  NAND2_X2 U11464 ( .A1(n9951), .A2(n9664), .ZN(n11364) );
  NAND2_X2 U11465 ( .A1(n10675), .A2(n10674), .ZN(n10020) );
  INV_X2 U11466 ( .A(n19244), .ZN(n19310) );
  NAND2_X1 U11467 ( .A1(n14557), .A2(n11917), .ZN(n14549) );
  AOI21_X1 U11468 ( .B1(n11858), .B2(n11495), .A(n11373), .ZN(n13606) );
  AND2_X2 U11469 ( .A1(n12387), .A2(n11306), .ZN(n11152) );
  NOR2_X2 U11470 ( .A1(n15019), .A2(n15021), .ZN(n12166) );
  INV_X1 U11471 ( .A(n13660), .ZN(n9676) );
  INV_X2 U11472 ( .A(n11141), .ZN(n13616) );
  NAND2_X2 U11473 ( .A1(n11364), .A2(n11353), .ZN(n13387) );
  XNOR2_X1 U11474 ( .A(n11856), .B(n13405), .ZN(n13402) );
  XNOR2_X1 U11475 ( .A(n11832), .B(n11339), .ZN(n13359) );
  AND2_X4 U11476 ( .A1(n13333), .A2(n11014), .ZN(n11072) );
  AND2_X1 U11477 ( .A1(n13344), .A2(n13083), .ZN(n9677) );
  AND2_X1 U11478 ( .A1(n13344), .A2(n13083), .ZN(n9678) );
  AND2_X1 U11479 ( .A1(n11014), .A2(n11015), .ZN(n9679) );
  AND2_X1 U11480 ( .A1(n11014), .A2(n11015), .ZN(n9680) );
  AND2_X2 U11481 ( .A1(n13346), .A2(n13330), .ZN(n9684) );
  OAI21_X1 U11482 ( .B1(n11347), .B2(n11234), .A(n10084), .ZN(n11240) );
  AND2_X4 U11483 ( .A1(n11015), .A2(n13083), .ZN(n11198) );
  AND2_X1 U11484 ( .A1(n13346), .A2(n13330), .ZN(n9683) );
  INV_X2 U11485 ( .A(n14551), .ZN(n16205) );
  AND2_X1 U11486 ( .A1(n9735), .A2(n12846), .ZN(n9917) );
  OAI22_X1 U11487 ( .A1(n10607), .A2(n12771), .B1(n10640), .B2(n10819), .ZN(
        n10611) );
  OR2_X1 U11488 ( .A1(n17791), .A2(n18050), .ZN(n16043) );
  OR2_X1 U11489 ( .A1(n16371), .A2(n12495), .ZN(n15257) );
  AND2_X1 U11490 ( .A1(n16394), .A2(n12721), .ZN(n15291) );
  AND4_X1 U11491 ( .A1(n10572), .A2(n10571), .A3(n10570), .A4(n10569), .ZN(
        n10583) );
  AND4_X1 U11492 ( .A1(n10580), .A2(n10579), .A3(n10578), .A4(n10577), .ZN(
        n10581) );
  AND4_X1 U11493 ( .A1(n10576), .A2(n10575), .A3(n10574), .A4(n10573), .ZN(
        n10582) );
  OR2_X1 U11494 ( .A1(n11292), .A2(n11291), .ZN(n11869) );
  AOI21_X1 U11495 ( .B1(n10819), .B2(n12771), .A(n12413), .ZN(n10633) );
  NAND2_X1 U11496 ( .A1(n9687), .A2(n9907), .ZN(n9906) );
  INV_X1 U11497 ( .A(n9908), .ZN(n9907) );
  NAND2_X1 U11498 ( .A1(n16174), .A2(n9827), .ZN(n10089) );
  INV_X1 U11499 ( .A(n14788), .ZN(n13218) );
  OR2_X1 U11500 ( .A1(n12282), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10867) );
  NAND2_X1 U11501 ( .A1(n12233), .A2(n12235), .ZN(n12236) );
  NAND2_X1 U11502 ( .A1(n15092), .A2(n9836), .ZN(n15033) );
  AND2_X1 U11503 ( .A1(n10248), .A2(n12054), .ZN(n9836) );
  AND2_X1 U11504 ( .A1(n9771), .A2(n15043), .ZN(n10248) );
  NAND2_X1 U11505 ( .A1(n15604), .A2(n10197), .ZN(n10196) );
  INV_X1 U11506 ( .A(n15242), .ZN(n10197) );
  NOR2_X1 U11507 ( .A1(n10131), .A2(n9918), .ZN(n9915) );
  INV_X1 U11508 ( .A(n12846), .ZN(n9918) );
  AND2_X1 U11509 ( .A1(n15044), .A2(n15036), .ZN(n10185) );
  NAND2_X1 U11510 ( .A1(n10051), .A2(n15572), .ZN(n10050) );
  INV_X1 U11511 ( .A(n10054), .ZN(n10051) );
  AOI21_X1 U11512 ( .B1(n10057), .B2(n10056), .A(n10055), .ZN(n10054) );
  INV_X1 U11513 ( .A(n15571), .ZN(n10055) );
  AND2_X2 U11514 ( .A1(n12842), .A2(n10030), .ZN(n12834) );
  NAND2_X1 U11515 ( .A1(n15668), .A2(n9731), .ZN(n12836) );
  AND4_X1 U11516 ( .A1(n10568), .A2(n10567), .A3(n10566), .A4(n10565), .ZN(
        n10584) );
  AND2_X1 U11517 ( .A1(n10508), .A2(n20089), .ZN(n10818) );
  AND2_X1 U11518 ( .A1(n10818), .A2(n13571), .ZN(n10959) );
  NAND2_X1 U11519 ( .A1(n10023), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10370) );
  NOR2_X1 U11520 ( .A1(n16786), .A2(n19148), .ZN(n14046) );
  NOR2_X1 U11521 ( .A1(n17178), .A2(n14035), .ZN(n15912) );
  NAND2_X1 U11522 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n9639), .ZN(
        n13940) );
  NOR2_X1 U11523 ( .A1(n14028), .A2(n15886), .ZN(n14048) );
  INV_X1 U11524 ( .A(n11819), .ZN(n11791) );
  AND2_X1 U11525 ( .A1(n13219), .A2(n13231), .ZN(n13132) );
  INV_X2 U11526 ( .A(n11544), .ZN(n11825) );
  NOR2_X1 U11527 ( .A1(n10257), .A2(n9807), .ZN(n10256) );
  INV_X1 U11528 ( .A(n14140), .ZN(n14163) );
  AND2_X1 U11529 ( .A1(n14549), .A2(n10129), .ZN(n12870) );
  NAND2_X1 U11530 ( .A1(n16173), .A2(n14647), .ZN(n10129) );
  AND2_X1 U11531 ( .A1(n20279), .A2(n13235), .ZN(n14648) );
  INV_X1 U11532 ( .A(n14648), .ZN(n14652) );
  OR2_X1 U11533 ( .A1(n12756), .A2(n12345), .ZN(n13563) );
  INV_X1 U11534 ( .A(n15682), .ZN(n13568) );
  AND2_X1 U11535 ( .A1(n12754), .A2(n12753), .ZN(n12856) );
  INV_X1 U11536 ( .A(n10593), .ZN(n12710) );
  XNOR2_X1 U11537 ( .A(n10290), .B(n10289), .ZN(n14096) );
  AND2_X1 U11538 ( .A1(n15617), .A2(n10071), .ZN(n10068) );
  AND2_X1 U11539 ( .A1(n9739), .A2(n16483), .ZN(n10224) );
  NOR2_X1 U11540 ( .A1(n15430), .A2(n15434), .ZN(n10240) );
  AOI21_X1 U11541 ( .B1(n15278), .B2(n9734), .A(n9957), .ZN(n9956) );
  INV_X1 U11542 ( .A(n15459), .ZN(n9845) );
  NAND2_X1 U11543 ( .A1(n15454), .A2(n15430), .ZN(n9846) );
  AND2_X1 U11544 ( .A1(n10755), .A2(n10754), .ZN(n15022) );
  AND2_X1 U11545 ( .A1(n10185), .A2(n10184), .ZN(n10183) );
  INV_X1 U11546 ( .A(n14837), .ZN(n10184) );
  NOR2_X1 U11547 ( .A1(n10132), .A2(n15382), .ZN(n10131) );
  INV_X1 U11548 ( .A(n9726), .ZN(n10132) );
  INV_X1 U11549 ( .A(n15567), .ZN(n13027) );
  NAND2_X1 U11550 ( .A1(n9980), .A2(n9808), .ZN(n16843) );
  NAND2_X1 U11551 ( .A1(n9989), .A2(n9987), .ZN(n16864) );
  NOR2_X1 U11552 ( .A1(n9985), .A2(n9988), .ZN(n9987) );
  INV_X1 U11553 ( .A(n9990), .ZN(n9988) );
  CLKBUF_X1 U11554 ( .A(n17146), .Z(n9985) );
  NAND2_X1 U11555 ( .A1(n16820), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16809) );
  NOR2_X1 U11556 ( .A1(n16821), .A2(n17773), .ZN(n16820) );
  NAND2_X1 U11557 ( .A1(n16044), .A2(n9859), .ZN(n16609) );
  NAND2_X1 U11558 ( .A1(n9865), .A2(n9743), .ZN(n10014) );
  INV_X1 U11559 ( .A(n17798), .ZN(n9865) );
  NAND2_X1 U11560 ( .A1(n16037), .A2(n10278), .ZN(n16038) );
  NAND2_X1 U11561 ( .A1(n16666), .A2(n15960), .ZN(n18050) );
  NOR3_X1 U11562 ( .A1(n18497), .A2(n14048), .A3(n14047), .ZN(n15983) );
  NOR2_X1 U11563 ( .A1(n15463), .A2(n15260), .ZN(n15263) );
  OAI21_X1 U11564 ( .B1(n17778), .B2(n9751), .A(n9699), .ZN(n10018) );
  NAND2_X1 U11565 ( .A1(n11017), .A2(n11018), .ZN(n9940) );
  NAND2_X1 U11566 ( .A1(n9936), .A2(n11970), .ZN(n9935) );
  OAI22_X1 U11567 ( .A1(n11969), .A2(n11968), .B1(n11967), .B2(n11966), .ZN(
        n9936) );
  NAND2_X1 U11568 ( .A1(n11971), .A2(n12379), .ZN(n9934) );
  NAND2_X1 U11569 ( .A1(n20846), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n9932) );
  NAND2_X1 U11570 ( .A1(n10484), .A2(n10483), .ZN(n10485) );
  NAND2_X1 U11571 ( .A1(n12329), .A2(n12737), .ZN(n9844) );
  NAND2_X1 U11572 ( .A1(n11131), .A2(n11143), .ZN(n11136) );
  OR2_X1 U11573 ( .A1(n11951), .A2(n11950), .ZN(n11953) );
  NAND2_X1 U11574 ( .A1(n11170), .A2(n11133), .ZN(n11130) );
  OR2_X1 U11575 ( .A1(n11362), .A2(n9787), .ZN(n9949) );
  NAND2_X1 U11576 ( .A1(n13622), .A2(n11897), .ZN(n11236) );
  INV_X1 U11577 ( .A(n11940), .ZN(n11974) );
  NOR2_X1 U11578 ( .A1(n11940), .A2(n11927), .ZN(n11971) );
  NAND2_X1 U11579 ( .A1(n10330), .A2(n10339), .ZN(n10337) );
  NAND2_X1 U11580 ( .A1(n12811), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10654) );
  NAND2_X1 U11581 ( .A1(n9954), .A2(n12461), .ZN(n12493) );
  INV_X1 U11582 ( .A(n10647), .ZN(n12732) );
  NOR2_X1 U11583 ( .A1(n17642), .A2(n15969), .ZN(n15973) );
  NOR2_X1 U11584 ( .A1(n11171), .A2(n10271), .ZN(n11172) );
  INV_X1 U11585 ( .A(n13232), .ZN(n11171) );
  NAND2_X1 U11586 ( .A1(n14320), .A2(n9909), .ZN(n9908) );
  INV_X1 U11587 ( .A(n14335), .ZN(n9909) );
  NAND2_X1 U11588 ( .A1(n13218), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11819) );
  INV_X1 U11589 ( .A(n10277), .ZN(n10254) );
  NOR2_X1 U11590 ( .A1(n11134), .A2(n20753), .ZN(n11495) );
  NOR2_X1 U11591 ( .A1(n10103), .A2(n9810), .ZN(n10102) );
  INV_X1 U11592 ( .A(n9803), .ZN(n10103) );
  INV_X1 U11593 ( .A(n14237), .ZN(n10106) );
  NAND2_X1 U11594 ( .A1(n14626), .A2(n10091), .ZN(n10090) );
  OAI21_X1 U11595 ( .B1(n9689), .B2(n10152), .A(n16173), .ZN(n10150) );
  NOR2_X1 U11596 ( .A1(n10098), .A2(n14311), .ZN(n10097) );
  INV_X1 U11597 ( .A(n10099), .ZN(n10098) );
  INV_X1 U11598 ( .A(n14415), .ZN(n10108) );
  INV_X1 U11599 ( .A(n11900), .ZN(n10080) );
  NAND2_X1 U11600 ( .A1(n9693), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9894) );
  INV_X1 U11601 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20602) );
  INV_X1 U11602 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20528) );
  NAND2_X1 U11603 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20096), .ZN(
        n12322) );
  NAND2_X1 U11604 ( .A1(n12712), .A2(n12706), .ZN(n10593) );
  NAND2_X1 U11605 ( .A1(n12688), .A2(n12706), .ZN(n12633) );
  INV_X1 U11606 ( .A(n12648), .ZN(n10117) );
  INV_X1 U11607 ( .A(n12600), .ZN(n10586) );
  INV_X1 U11608 ( .A(n12601), .ZN(n10120) );
  NAND2_X1 U11609 ( .A1(n12755), .A2(n10665), .ZN(n10659) );
  NAND2_X1 U11610 ( .A1(n15139), .A2(n10211), .ZN(n10210) );
  INV_X1 U11611 ( .A(n15145), .ZN(n10211) );
  AOI211_X1 U11612 ( .C1(n12257), .C2(n12260), .A(n12256), .B(n14971), .ZN(
        n12258) );
  NAND2_X1 U11613 ( .A1(n9833), .A2(n12212), .ZN(n12216) );
  INV_X1 U11614 ( .A(n15172), .ZN(n10205) );
  INV_X1 U11615 ( .A(n15050), .ZN(n10249) );
  NOR2_X1 U11616 ( .A1(n12997), .A2(n15751), .ZN(n12229) );
  NOR2_X1 U11617 ( .A1(n16500), .A2(n10170), .ZN(n10169) );
  AND2_X1 U11618 ( .A1(n9717), .A2(n10180), .ZN(n10179) );
  AOI21_X1 U11619 ( .B1(n15311), .B2(n10221), .A(n9728), .ZN(n10220) );
  INV_X1 U11620 ( .A(n15317), .ZN(n10221) );
  INV_X1 U11621 ( .A(n15318), .ZN(n9963) );
  INV_X1 U11622 ( .A(n15311), .ZN(n10222) );
  INV_X1 U11623 ( .A(n10220), .ZN(n9959) );
  NAND2_X1 U11624 ( .A1(n10070), .A2(n9694), .ZN(n15328) );
  INV_X1 U11625 ( .A(n15232), .ZN(n10194) );
  AND2_X1 U11626 ( .A1(n15074), .A2(n10176), .ZN(n10175) );
  NOR2_X1 U11627 ( .A1(n15095), .A2(n15096), .ZN(n14855) );
  INV_X1 U11628 ( .A(n16468), .ZN(n10071) );
  OR2_X1 U11629 ( .A1(n12842), .A2(n12844), .ZN(n12846) );
  AND2_X1 U11630 ( .A1(n10188), .A2(n10187), .ZN(n10186) );
  INV_X1 U11631 ( .A(n13586), .ZN(n10187) );
  INV_X1 U11632 ( .A(n10784), .ZN(n10777) );
  NOR2_X1 U11633 ( .A1(n10564), .A2(n10563), .ZN(n12589) );
  NAND2_X1 U11634 ( .A1(n13702), .A2(n9967), .ZN(n9966) );
  AOI21_X1 U11635 ( .B1(n9970), .B2(n9967), .A(n9965), .ZN(n9964) );
  INV_X1 U11636 ( .A(n15672), .ZN(n9965) );
  AOI21_X1 U11637 ( .B1(n14936), .B2(n10861), .A(n12785), .ZN(n9974) );
  AND2_X1 U11638 ( .A1(n13703), .A2(n9972), .ZN(n9971) );
  NAND2_X1 U11639 ( .A1(n14936), .A2(n9973), .ZN(n9972) );
  AND2_X1 U11640 ( .A1(n12843), .A2(n12785), .ZN(n9973) );
  NAND2_X1 U11641 ( .A1(n10234), .A2(n10233), .ZN(n12829) );
  NAND2_X1 U11642 ( .A1(n9919), .A2(n12493), .ZN(n12494) );
  INV_X1 U11643 ( .A(n10233), .ZN(n9919) );
  INV_X1 U11644 ( .A(n13492), .ZN(n10190) );
  INV_X1 U11645 ( .A(n10998), .ZN(n10989) );
  NOR2_X1 U11646 ( .A1(n10422), .A2(n10421), .ZN(n10428) );
  AND2_X1 U11647 ( .A1(n12229), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12018) );
  INV_X1 U11648 ( .A(n12444), .ZN(n12423) );
  NAND2_X1 U11649 ( .A1(n10348), .A2(n10347), .ZN(n12334) );
  NAND2_X1 U11650 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19092), .ZN(
        n13941) );
  NAND2_X1 U11651 ( .A1(n19092), .A2(n19102), .ZN(n9994) );
  AND2_X1 U11652 ( .A1(n15929), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n9873) );
  NAND2_X1 U11653 ( .A1(n9658), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n9863) );
  NOR4_X1 U11654 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A4(n19115), .ZN(n15913) );
  NOR2_X1 U11655 ( .A1(n13940), .A2(n13939), .ZN(n15940) );
  NAND2_X1 U11656 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10001) );
  AOI22_X1 U11657 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10002) );
  NOR2_X1 U11658 ( .A1(n13941), .A2(n13939), .ZN(n15911) );
  NAND2_X1 U11659 ( .A1(n10154), .A2(n9695), .ZN(n15982) );
  NAND2_X1 U11660 ( .A1(n10008), .A2(n18099), .ZN(n10006) );
  NOR2_X1 U11661 ( .A1(n18085), .A2(n10010), .ZN(n10009) );
  INV_X1 U11662 ( .A(n10009), .ZN(n10007) );
  INV_X1 U11663 ( .A(n15975), .ZN(n10008) );
  XNOR2_X1 U11664 ( .A(n15995), .B(n17647), .ZN(n15967) );
  INV_X1 U11665 ( .A(n14236), .ZN(n10255) );
  INV_X1 U11666 ( .A(n13656), .ZN(n20842) );
  AND3_X1 U11667 ( .A1(n14181), .A2(n14286), .A3(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n14254) );
  AND2_X1 U11668 ( .A1(n10264), .A2(n10263), .ZN(n10262) );
  INV_X1 U11669 ( .A(n11991), .ZN(n10263) );
  INV_X1 U11670 ( .A(n14349), .ZN(n11547) );
  NAND2_X1 U11671 ( .A1(n9901), .A2(n11452), .ZN(n13895) );
  NAND2_X1 U11672 ( .A1(n9902), .A2(n9905), .ZN(n9901) );
  NAND2_X1 U11673 ( .A1(n13633), .A2(n9903), .ZN(n9902) );
  NAND2_X1 U11674 ( .A1(n11842), .A2(n11338), .ZN(n10251) );
  AOI21_X1 U11675 ( .B1(n11338), .B2(n11529), .A(n10253), .ZN(n10252) );
  INV_X1 U11676 ( .A(n11351), .ZN(n10253) );
  NAND2_X1 U11677 ( .A1(n13147), .A2(n13146), .ZN(n13399) );
  NAND2_X1 U11678 ( .A1(n9943), .A2(n9942), .ZN(n11998) );
  NAND2_X1 U11679 ( .A1(n14549), .A2(n14647), .ZN(n9943) );
  AND2_X1 U11680 ( .A1(n14526), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9942) );
  NOR2_X1 U11681 ( .A1(n10087), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10086) );
  INV_X1 U11682 ( .A(n11917), .ZN(n10087) );
  INV_X1 U11683 ( .A(n14549), .ZN(n14536) );
  OR2_X1 U11684 ( .A1(n14300), .A2(n14283), .ZN(n14285) );
  OAI21_X1 U11685 ( .B1(n9947), .B2(n10091), .A(n14626), .ZN(n9946) );
  NOR2_X1 U11686 ( .A1(n14411), .A2(n14352), .ZN(n14351) );
  AND2_X1 U11687 ( .A1(n10094), .A2(n10093), .ZN(n13373) );
  INV_X1 U11688 ( .A(n13299), .ZN(n10093) );
  INV_X1 U11689 ( .A(n13300), .ZN(n10094) );
  AND2_X1 U11690 ( .A1(n13218), .A2(n12973), .ZN(n13231) );
  AND2_X1 U11691 ( .A1(n20287), .A2(n14643), .ZN(n16284) );
  AND2_X1 U11692 ( .A1(n13660), .A2(n9666), .ZN(n14140) );
  INV_X1 U11693 ( .A(n9673), .ZN(n13389) );
  AND2_X1 U11694 ( .A1(n12952), .A2(n9666), .ZN(n14793) );
  NOR2_X1 U11695 ( .A1(n20601), .A2(n20298), .ZN(n20536) );
  INV_X1 U11696 ( .A(n20569), .ZN(n20560) );
  NAND2_X1 U11697 ( .A1(n20846), .A2(n13421), .ZN(n20298) );
  AOI21_X1 U11698 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20643), .A(n20298), 
        .ZN(n20650) );
  NOR2_X1 U11699 ( .A1(n13219), .A2(n16112), .ZN(n16087) );
  INV_X1 U11700 ( .A(n19985), .ZN(n20123) );
  NAND2_X1 U11701 ( .A1(n10120), .A2(n10586), .ZN(n12610) );
  AND2_X1 U11702 ( .A1(n13589), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10247) );
  INV_X1 U11703 ( .A(n13446), .ZN(n10246) );
  OR2_X1 U11704 ( .A1(n15014), .A2(n15016), .ZN(n10245) );
  NOR2_X1 U11705 ( .A1(n15199), .A2(n15201), .ZN(n15200) );
  INV_X1 U11706 ( .A(n10643), .ZN(n13014) );
  AND2_X1 U11707 ( .A1(n15053), .A2(n9792), .ZN(n15025) );
  INV_X1 U11708 ( .A(n15022), .ZN(n10182) );
  NAND2_X1 U11709 ( .A1(n9848), .A2(n9780), .ZN(n15523) );
  INV_X1 U11710 ( .A(n15553), .ZN(n9848) );
  AOI21_X1 U11711 ( .B1(n10045), .B2(n10052), .A(n9786), .ZN(n10044) );
  OR2_X1 U11712 ( .A1(n15068), .A2(n15059), .ZN(n15061) );
  NOR2_X2 U11713 ( .A1(n15061), .A2(n15051), .ZN(n15053) );
  AND2_X1 U11714 ( .A1(n15373), .A2(n16435), .ZN(n10059) );
  AND2_X1 U11715 ( .A1(n14855), .A2(n10175), .ZN(n15076) );
  AOI21_X1 U11716 ( .B1(n10066), .B2(n10065), .A(n10064), .ZN(n10063) );
  AND3_X1 U11717 ( .A1(n10803), .A2(n10802), .A3(n10801), .ZN(n16528) );
  INV_X1 U11718 ( .A(n12609), .ZN(n10225) );
  INV_X1 U11719 ( .A(n15396), .ZN(n10239) );
  NAND2_X1 U11720 ( .A1(n12836), .A2(n10275), .ZN(n9921) );
  NOR2_X1 U11722 ( .A1(n12835), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15418) );
  INV_X1 U11723 ( .A(n12836), .ZN(n15423) );
  NAND2_X1 U11724 ( .A1(n12034), .A2(n12033), .ZN(n12038) );
  NAND2_X1 U11725 ( .A1(n12013), .A2(n20089), .ZN(n12040) );
  XNOR2_X1 U11726 ( .A(n12045), .B(n12046), .ZN(n13160) );
  NAND2_X1 U11727 ( .A1(n19727), .A2(n15723), .ZN(n19636) );
  NAND2_X1 U11728 ( .A1(n20075), .A2(n15724), .ZN(n19728) );
  INV_X1 U11729 ( .A(n20064), .ZN(n19553) );
  NAND2_X2 U11730 ( .A1(n10399), .A2(n10398), .ZN(n10647) );
  NAND2_X1 U11731 ( .A1(n10279), .A2(n10384), .ZN(n10399) );
  NAND2_X1 U11732 ( .A1(n10397), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10398) );
  NOR2_X1 U11733 ( .A1(n10383), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10384) );
  NAND2_X1 U11734 ( .A1(n19440), .A2(n20082), .ZN(n19864) );
  NAND2_X1 U11735 ( .A1(n15702), .A2(n15701), .ZN(n19919) );
  OR2_X1 U11736 ( .A1(n16602), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15702) );
  AND2_X1 U11737 ( .A1(n13519), .A2(n13518), .ZN(n15685) );
  AND2_X1 U11738 ( .A1(n17803), .A2(n17816), .ZN(n9991) );
  INV_X1 U11739 ( .A(n17858), .ZN(n9986) );
  OR2_X1 U11740 ( .A1(n16938), .A2(n17146), .ZN(n16927) );
  INV_X1 U11741 ( .A(n18501), .ZN(n17511) );
  NAND2_X1 U11742 ( .A1(n19092), .A2(n19102), .ZN(n10155) );
  NAND2_X1 U11743 ( .A1(n15921), .A2(n15920), .ZN(n15922) );
  NAND2_X1 U11744 ( .A1(n13964), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n15920) );
  NAND2_X1 U11745 ( .A1(n17769), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16821) );
  NAND2_X1 U11746 ( .A1(n9861), .A2(n16610), .ZN(n16102) );
  NAND2_X1 U11747 ( .A1(n16044), .A2(n9809), .ZN(n9861) );
  INV_X1 U11748 ( .A(n10014), .ZN(n9864) );
  INV_X1 U11749 ( .A(n9867), .ZN(n17830) );
  NAND2_X1 U11750 ( .A1(n9853), .A2(n9852), .ZN(n9857) );
  AOI21_X1 U11751 ( .B1(n18050), .B2(n16032), .A(n9768), .ZN(n9852) );
  NAND2_X1 U11752 ( .A1(n16033), .A2(n18050), .ZN(n9853) );
  OAI21_X1 U11753 ( .B1(n16033), .B2(n16032), .A(n18050), .ZN(n16035) );
  NOR2_X1 U11754 ( .A1(n16021), .A2(n18048), .ZN(n18309) );
  NAND2_X1 U11755 ( .A1(n9889), .A2(n16009), .ZN(n9887) );
  NOR2_X1 U11756 ( .A1(n18100), .A2(n18099), .ZN(n18098) );
  OAI21_X1 U11757 ( .B1(n14064), .B2(n17660), .A(n14063), .ZN(n18950) );
  AOI21_X1 U11758 ( .B1(n11772), .B2(n11771), .A(n11770), .ZN(n12868) );
  NAND2_X1 U11759 ( .A1(n9692), .A2(n11144), .ZN(n13109) );
  NAND2_X1 U11760 ( .A1(n14331), .A2(n9825), .ZN(n14250) );
  AND2_X1 U11761 ( .A1(n14331), .A2(n9822), .ZN(n14277) );
  AND2_X1 U11762 ( .A1(n14331), .A2(n14180), .ZN(n14305) );
  NAND3_X1 U11763 ( .A1(n16147), .A2(P1_REIP_REG_14__SCAN_IN), .A3(
        P1_REIP_REG_13__SCAN_IN), .ZN(n16146) );
  INV_X1 U11764 ( .A(n20178), .ZN(n20151) );
  INV_X2 U11765 ( .A(n13163), .ZN(n20274) );
  XNOR2_X1 U11766 ( .A(n11985), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13669) );
  OR2_X1 U11767 ( .A1(n11984), .A2(n11993), .ZN(n11985) );
  NAND2_X1 U11768 ( .A1(n9910), .A2(n12003), .ZN(n14447) );
  OR2_X1 U11769 ( .A1(n9686), .A2(n12002), .ZN(n12003) );
  INV_X1 U11770 ( .A(n16202), .ZN(n16204) );
  NAND2_X1 U11771 ( .A1(n13643), .A2(n13476), .ZN(n14551) );
  NAND2_X1 U11772 ( .A1(n20135), .A2(n11981), .ZN(n16209) );
  XNOR2_X1 U11773 ( .A(n11924), .B(n11923), .ZN(n14668) );
  XNOR2_X1 U11774 ( .A(n10082), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14677) );
  NAND2_X1 U11775 ( .A1(n11995), .A2(n11996), .ZN(n10082) );
  XNOR2_X1 U11776 ( .A(n12873), .B(n14160), .ZN(n14696) );
  AND2_X1 U11777 ( .A1(n14661), .A2(n14657), .ZN(n14735) );
  NAND2_X1 U11778 ( .A1(n13238), .A2(n14793), .ZN(n20287) );
  INV_X1 U11779 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20643) );
  INV_X1 U11780 ( .A(n13419), .ZN(n13781) );
  CLKBUF_X1 U11781 ( .A(n13651), .Z(n13652) );
  INV_X1 U11782 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20532) );
  INV_X1 U11783 ( .A(n20681), .ZN(n20729) );
  INV_X1 U11784 ( .A(n20068), .ZN(n19868) );
  AND2_X1 U11785 ( .A1(n14917), .A2(n10596), .ZN(n19153) );
  AND2_X1 U11786 ( .A1(n14917), .A2(n12796), .ZN(n20111) );
  AND2_X1 U11787 ( .A1(n12707), .A2(n12706), .ZN(n16394) );
  INV_X1 U11788 ( .A(n19301), .ZN(n19325) );
  NOR2_X1 U11789 ( .A1(n15121), .A2(n12366), .ZN(n11000) );
  AND2_X1 U11790 ( .A1(n19357), .A2(n12353), .ZN(n16417) );
  AND2_X1 U11791 ( .A1(n12351), .A2(n13010), .ZN(n19357) );
  OR2_X1 U11792 ( .A1(n13514), .A2(n12350), .ZN(n12351) );
  OAI21_X1 U11793 ( .B1(n11002), .B2(n16433), .A(n14098), .ZN(n14099) );
  OAI21_X1 U11794 ( .B1(n9685), .B2(n10180), .A(n9725), .ZN(n16348) );
  NAND2_X1 U11795 ( .A1(n15276), .A2(n19435), .ZN(n10138) );
  INV_X1 U11796 ( .A(n15275), .ZN(n10137) );
  INV_X1 U11797 ( .A(n15452), .ZN(n10140) );
  NOR2_X1 U11798 ( .A1(n15451), .A2(n19429), .ZN(n10139) );
  NAND2_X1 U11799 ( .A1(n12913), .A2(n12857), .ZN(n19438) );
  NAND2_X1 U11800 ( .A1(n12864), .A2(n20122), .ZN(n19431) );
  INV_X1 U11801 ( .A(n19431), .ZN(n16495) );
  NOR2_X1 U11802 ( .A1(n14093), .A2(n14092), .ZN(n14094) );
  NAND2_X1 U11803 ( .A1(n10212), .A2(n14086), .ZN(n14091) );
  XNOR2_X1 U11804 ( .A(n9725), .B(n12414), .ZN(n14807) );
  XNOR2_X1 U11805 ( .A(n14093), .B(n14092), .ZN(n12865) );
  NAND2_X1 U11806 ( .A1(n14093), .A2(n10022), .ZN(n9925) );
  NAND2_X1 U11807 ( .A1(n9724), .A2(n15434), .ZN(n10022) );
  AND2_X1 U11808 ( .A1(n15258), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10110) );
  NOR2_X1 U11809 ( .A1(n15274), .A2(n15453), .ZN(n15451) );
  NOR2_X1 U11810 ( .A1(n15285), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15452) );
  AND2_X1 U11811 ( .A1(n15486), .A2(n12792), .ZN(n15481) );
  OR2_X1 U11812 ( .A1(n16525), .A2(n12847), .ZN(n12788) );
  INV_X1 U11813 ( .A(n16563), .ZN(n16582) );
  INV_X1 U11814 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20096) );
  INV_X1 U11815 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20089) );
  NOR2_X2 U11816 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20068) );
  NAND2_X1 U11817 ( .A1(n16865), .A2(n17786), .ZN(n9979) );
  NAND2_X1 U11818 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n17189), .ZN(n17180) );
  INV_X1 U11819 ( .A(n18512), .ZN(n17489) );
  INV_X1 U11820 ( .A(n16648), .ZN(n10166) );
  NAND2_X1 U11821 ( .A1(n16609), .A2(n10167), .ZN(n16645) );
  AND2_X1 U11822 ( .A1(n16044), .A2(n17780), .ZN(n16045) );
  INV_X1 U11823 ( .A(n10016), .ZN(n10015) );
  AOI21_X1 U11824 ( .B1(n18214), .B2(n17783), .A(n17774), .ZN(n10016) );
  NOR2_X1 U11825 ( .A1(n18211), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9879) );
  NAND2_X1 U11826 ( .A1(n18218), .A2(n9881), .ZN(n9880) );
  AND2_X1 U11827 ( .A1(n9882), .A2(n18209), .ZN(n9881) );
  AOI21_X1 U11828 ( .B1(n18265), .B2(n18205), .A(n18210), .ZN(n9882) );
  AND2_X1 U11829 ( .A1(n18225), .A2(n9884), .ZN(n18218) );
  AOI21_X1 U11830 ( .B1(n18333), .B2(n18208), .A(n9885), .ZN(n9884) );
  NOR2_X1 U11831 ( .A1(n18953), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9885) );
  AOI211_X1 U11832 ( .C1(n15882), .C2(n16607), .A(n15881), .B(n15880), .ZN(
        n15889) );
  OAI21_X1 U11833 ( .B1(n9929), .B2(n9928), .A(n9926), .ZN(n11956) );
  INV_X1 U11834 ( .A(n12380), .ZN(n9928) );
  NAND2_X1 U11835 ( .A1(n11962), .A2(n9927), .ZN(n9926) );
  AND2_X1 U11836 ( .A1(n9666), .A2(n12380), .ZN(n9927) );
  NOR2_X1 U11837 ( .A1(n13649), .A2(n11944), .ZN(n11967) );
  NAND2_X1 U11838 ( .A1(n11962), .A2(n9666), .ZN(n9930) );
  AND2_X1 U11839 ( .A1(n9666), .A2(n11949), .ZN(n9929) );
  OAI22_X1 U11840 ( .A1(n10659), .A2(n10624), .B1(n10677), .B2(n14954), .ZN(
        n10625) );
  NAND2_X1 U11841 ( .A1(n10679), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10627) );
  INV_X1 U11842 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12468) );
  CLKBUF_X1 U11843 ( .A(n12275), .Z(n12283) );
  CLKBUF_X1 U11844 ( .A(n12132), .Z(n12284) );
  CLKBUF_X1 U11845 ( .A(n12133), .Z(n12281) );
  INV_X1 U11846 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12471) );
  INV_X1 U11847 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12465) );
  INV_X1 U11848 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12481) );
  AOI22_X1 U11849 ( .A1(n10450), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9642), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10357) );
  NAND2_X1 U11850 ( .A1(n11932), .A2(n11931), .ZN(n11939) );
  INV_X1 U11851 ( .A(n14223), .ZN(n10105) );
  NOR2_X1 U11852 ( .A1(n11236), .A2(n20846), .ZN(n11239) );
  OR2_X1 U11853 ( .A1(n11322), .A2(n11321), .ZN(n11885) );
  OR2_X1 U11854 ( .A1(n11302), .A2(n11301), .ZN(n11876) );
  OR2_X1 U11855 ( .A1(n11251), .A2(n11250), .ZN(n11843) );
  NOR2_X1 U11856 ( .A1(n11190), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9897) );
  NAND2_X1 U11857 ( .A1(n11138), .A2(n11306), .ZN(n11131) );
  NOR2_X1 U11858 ( .A1(n9941), .A2(n9940), .ZN(n9939) );
  OR2_X1 U11859 ( .A1(n11280), .A2(n11279), .ZN(n11859) );
  AOI21_X1 U11860 ( .B1(n9933), .B2(n9778), .A(n9931), .ZN(n11976) );
  NAND2_X1 U11861 ( .A1(n11975), .A2(n9932), .ZN(n9931) );
  NAND2_X1 U11862 ( .A1(n9935), .A2(n9934), .ZN(n9933) );
  AND2_X1 U11863 ( .A1(n10333), .A2(n10332), .ZN(n10344) );
  OR2_X1 U11864 ( .A1(n10337), .A2(n10335), .ZN(n10333) );
  AND2_X1 U11865 ( .A1(n10592), .A2(n10116), .ZN(n10115) );
  INV_X1 U11866 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10114) );
  INV_X1 U11867 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12464) );
  INV_X1 U11868 ( .A(n10058), .ZN(n10056) );
  AND2_X1 U11869 ( .A1(n12591), .A2(n12590), .ZN(n12838) );
  NOR2_X1 U11870 ( .A1(n10486), .A2(n10485), .ZN(n10494) );
  INV_X2 U11871 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13522) );
  INV_X1 U11872 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12432) );
  INV_X1 U11873 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12430) );
  INV_X1 U11874 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12453) );
  AOI22_X1 U11875 ( .A1(n10372), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12287), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10024) );
  AOI22_X1 U11876 ( .A1(n10371), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9640), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10361) );
  AOI22_X1 U11877 ( .A1(n10372), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12287), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n9955) );
  AND2_X1 U11878 ( .A1(n9842), .A2(n12327), .ZN(n9841) );
  INV_X1 U11879 ( .A(n9843), .ZN(n9842) );
  OAI21_X1 U11880 ( .B1(n12765), .B2(n12328), .A(n9844), .ZN(n9843) );
  NAND2_X1 U11881 ( .A1(n12771), .A2(n10615), .ZN(n12335) );
  NOR2_X1 U11882 ( .A1(n17635), .A2(n15976), .ZN(n15977) );
  AND2_X1 U11883 ( .A1(n11937), .A2(n11936), .ZN(n12378) );
  OR2_X1 U11884 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20294), .ZN(
        n11936) );
  OR2_X1 U11885 ( .A1(n11972), .A2(n11935), .ZN(n11937) );
  AND2_X1 U11886 ( .A1(n14254), .A2(n14173), .ZN(n14227) );
  AOI22_X1 U11887 ( .A1(n11050), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9672), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11053) );
  AOI21_X1 U11888 ( .B1(n11055), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n11056), .ZN(n11060) );
  AND2_X1 U11889 ( .A1(n11112), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11056) );
  AOI22_X1 U11890 ( .A1(n11072), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9669), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11059) );
  AND2_X1 U11891 ( .A1(n11766), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11767) );
  OR2_X1 U11892 ( .A1(n10260), .A2(n10258), .ZN(n10257) );
  NAND2_X1 U11893 ( .A1(n10261), .A2(n13930), .ZN(n10260) );
  INV_X1 U11894 ( .A(n14360), .ZN(n10261) );
  INV_X1 U11895 ( .A(n13928), .ZN(n10259) );
  NOR2_X1 U11896 ( .A1(n11368), .A2(n16210), .ZN(n11323) );
  NAND2_X1 U11897 ( .A1(n9911), .A2(n9787), .ZN(n11305) );
  NAND2_X1 U11898 ( .A1(n9951), .A2(n9950), .ZN(n9911) );
  NOR2_X1 U11899 ( .A1(n13390), .A2(n11362), .ZN(n9950) );
  INV_X1 U11900 ( .A(n13606), .ZN(n11374) );
  CLKBUF_X1 U11901 ( .A(n11925), .Z(n11926) );
  INV_X1 U11902 ( .A(n14262), .ZN(n10104) );
  NOR2_X1 U11903 ( .A1(n14323), .A2(n10100), .ZN(n10099) );
  INV_X1 U11904 ( .A(n14336), .ZN(n10100) );
  INV_X1 U11905 ( .A(n11904), .ZN(n10088) );
  AND2_X1 U11906 ( .A1(n16174), .A2(n11904), .ZN(n10091) );
  AND2_X1 U11907 ( .A1(n16170), .A2(n11907), .ZN(n14757) );
  AND2_X1 U11908 ( .A1(n14166), .A2(n13292), .ZN(n14164) );
  INV_X1 U11909 ( .A(n11239), .ZN(n11893) );
  OR2_X1 U11910 ( .A1(n11221), .A2(n11220), .ZN(n11897) );
  NOR2_X1 U11911 ( .A1(n13757), .A2(n10096), .ZN(n10095) );
  INV_X1 U11912 ( .A(n13723), .ZN(n10096) );
  NOR2_X1 U11913 ( .A1(n14188), .A2(n14163), .ZN(n14154) );
  NAND2_X1 U11914 ( .A1(n11133), .A2(n9666), .ZN(n11927) );
  NAND2_X1 U11915 ( .A1(n11586), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11037) );
  AND2_X1 U11916 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11042) );
  OR2_X1 U11917 ( .A1(n11233), .A2(n11232), .ZN(n11844) );
  NAND2_X1 U11918 ( .A1(n13622), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11270) );
  NAND3_X1 U11919 ( .A1(n11138), .A2(n13660), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11940) );
  NOR2_X1 U11920 ( .A1(n11204), .A2(n11203), .ZN(n11846) );
  NAND2_X1 U11921 ( .A1(n11154), .A2(n11132), .ZN(n11155) );
  INV_X1 U11922 ( .A(n11131), .ZN(n11132) );
  CLKBUF_X1 U11923 ( .A(n13078), .Z(n13079) );
  INV_X1 U11924 ( .A(n11134), .ZN(n11170) );
  AND4_X1 U11925 ( .A1(n11070), .A2(n11069), .A3(n11068), .A4(n11067), .ZN(
        n11071) );
  INV_X1 U11926 ( .A(n13357), .ZN(n13421) );
  AOI21_X1 U11927 ( .B1(n20845), .B2(n16341), .A(n16095), .ZN(n13357) );
  AND2_X1 U11928 ( .A1(n16062), .A2(n16345), .ZN(n13349) );
  AOI21_X1 U11929 ( .B1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n20088), .A(
        n10329), .ZN(n10341) );
  NOR2_X1 U11930 ( .A1(n12716), .A2(n12717), .ZN(n12725) );
  INV_X1 U11931 ( .A(n12694), .ZN(n10113) );
  NAND2_X1 U11932 ( .A1(n10593), .A2(n12711), .ZN(n12716) );
  AND2_X1 U11933 ( .A1(n12656), .A2(n12639), .ZN(n12664) );
  INV_X1 U11934 ( .A(n10538), .ZN(n12512) );
  AND2_X1 U11935 ( .A1(n10727), .A2(n10177), .ZN(n10176) );
  INV_X1 U11936 ( .A(n15080), .ZN(n10177) );
  AND2_X1 U11937 ( .A1(n12166), .A2(n12187), .ZN(n12167) );
  INV_X1 U11938 ( .A(n15192), .ZN(n10206) );
  NAND2_X1 U11939 ( .A1(n15029), .A2(n15030), .ZN(n15019) );
  AND2_X1 U11940 ( .A1(n12076), .A2(n12055), .ZN(n10250) );
  INV_X1 U11941 ( .A(n14858), .ZN(n10195) );
  NOR2_X1 U11942 ( .A1(n10159), .A2(n10157), .ZN(n10156) );
  AND2_X1 U11943 ( .A1(n10295), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10292) );
  NOR2_X1 U11944 ( .A1(n14840), .A2(n10300), .ZN(n10295) );
  NOR2_X1 U11945 ( .A1(n16428), .A2(n10162), .ZN(n10161) );
  INV_X1 U11946 ( .A(n14856), .ZN(n10727) );
  INV_X1 U11947 ( .A(n15258), .ZN(n9957) );
  INV_X1 U11948 ( .A(n14976), .ZN(n10181) );
  AND2_X1 U11949 ( .A1(n10983), .A2(n10982), .ZN(n15145) );
  NAND2_X1 U11950 ( .A1(n9710), .A2(n14827), .ZN(n10204) );
  NAND2_X1 U11951 ( .A1(n9653), .A2(n9824), .ZN(n10142) );
  NOR2_X1 U11952 ( .A1(n15536), .A2(n12634), .ZN(n10236) );
  INV_X1 U11953 ( .A(n15333), .ZN(n10046) );
  AND2_X1 U11954 ( .A1(n12848), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10238) );
  INV_X1 U11955 ( .A(n10068), .ZN(n10065) );
  INV_X1 U11956 ( .A(n16452), .ZN(n10064) );
  OR2_X1 U11957 ( .A1(n10202), .A2(n13273), .ZN(n10201) );
  AND2_X1 U11958 ( .A1(n10716), .A2(n10715), .ZN(n14870) );
  NAND2_X1 U11959 ( .A1(n10203), .A2(n16560), .ZN(n10202) );
  INV_X1 U11960 ( .A(n13180), .ZN(n10203) );
  AND2_X1 U11961 ( .A1(n13443), .A2(n13457), .ZN(n10188) );
  INV_X1 U11962 ( .A(n15418), .ZN(n10237) );
  OR2_X1 U11963 ( .A1(n10550), .A2(n10549), .ZN(n12552) );
  NAND2_X1 U11964 ( .A1(n10025), .A2(n12826), .ZN(n12830) );
  INV_X1 U11965 ( .A(n13701), .ZN(n10026) );
  NAND2_X1 U11966 ( .A1(n10689), .A2(n10688), .ZN(n10690) );
  NAND2_X1 U11967 ( .A1(n10020), .A2(n12020), .ZN(n10683) );
  XNOR2_X1 U11968 ( .A(n12022), .B(n12021), .ZN(n12023) );
  INV_X1 U11969 ( .A(n13517), .ZN(n12736) );
  INV_X1 U11970 ( .A(n19459), .ZN(n10632) );
  NAND2_X1 U11971 ( .A1(n10382), .A2(n10381), .ZN(n10383) );
  NAND3_X1 U11972 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n20068), .A3(n19919), 
        .ZN(n15708) );
  AOI21_X1 U11974 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n18968), .A(
        n14044), .ZN(n14052) );
  NAND3_X1 U11975 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(n19108), .ZN(n13938) );
  NOR4_X1 U11976 ( .A1(n18054), .A2(n17081), .A3(n18022), .A4(n18009), .ZN(
        n17018) );
  NOR2_X1 U11977 ( .A1(n9860), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9859) );
  INV_X1 U11978 ( .A(n17780), .ZN(n9860) );
  OAI211_X1 U11979 ( .C1(n16033), .C2(n9856), .A(n9855), .B(n9854), .ZN(n9858)
         );
  OR2_X1 U11980 ( .A1(n17952), .A2(n9856), .ZN(n9854) );
  NAND2_X1 U11981 ( .A1(n15982), .A2(n9806), .ZN(n9855) );
  AND2_X1 U11982 ( .A1(n15977), .A2(n16010), .ZN(n15960) );
  INV_X1 U11983 ( .A(n16013), .ZN(n9889) );
  AND2_X1 U11984 ( .A1(n12952), .A2(n12953), .ZN(n12959) );
  AND2_X1 U11985 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n14172), .ZN(n14286) );
  NOR2_X1 U11986 ( .A1(n20753), .A2(n13768), .ZN(n13663) );
  INV_X1 U11987 ( .A(n13734), .ZN(n13768) );
  AND2_X1 U11988 ( .A1(n13076), .A2(n10282), .ZN(n11180) );
  INV_X1 U11989 ( .A(n13763), .ZN(n13736) );
  NAND2_X1 U11990 ( .A1(n12386), .A2(n12385), .ZN(n13101) );
  AND2_X1 U11991 ( .A1(n20753), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11824) );
  NAND2_X1 U11992 ( .A1(n11767), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11821) );
  AND2_X1 U11993 ( .A1(n14226), .A2(n13644), .ZN(n11745) );
  OR2_X1 U11994 ( .A1(n14519), .A2(n9799), .ZN(n11728) );
  NOR2_X1 U11995 ( .A1(n11681), .A2(n14550), .ZN(n11682) );
  NAND2_X1 U11996 ( .A1(n11682), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11723) );
  AND2_X1 U11997 ( .A1(n14555), .A2(n13644), .ZN(n11661) );
  INV_X1 U11998 ( .A(n11631), .ZN(n11632) );
  NAND2_X1 U11999 ( .A1(n11633), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11681) );
  CLKBUF_X1 U12000 ( .A(n14280), .Z(n14281) );
  NAND2_X1 U12001 ( .A1(n11598), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11631) );
  AND2_X1 U12002 ( .A1(n11581), .A2(n11580), .ZN(n14320) );
  AND2_X1 U12003 ( .A1(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n11563), .ZN(
        n11564) );
  NAND2_X1 U12004 ( .A1(n11564), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11597) );
  INV_X1 U12005 ( .A(n11542), .ZN(n11563) );
  NOR2_X1 U12006 ( .A1(n11515), .A2(n16141), .ZN(n11499) );
  NAND2_X1 U12007 ( .A1(n11499), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11542) );
  NOR2_X1 U12008 ( .A1(n11483), .A2(n14621), .ZN(n11498) );
  NAND2_X1 U12009 ( .A1(n11468), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11483) );
  INV_X1 U12010 ( .A(n11467), .ZN(n11468) );
  INV_X1 U12011 ( .A(n13895), .ZN(n11451) );
  NOR2_X1 U12012 ( .A1(n11430), .A2(n20155), .ZN(n11434) );
  OR2_X1 U12013 ( .A1(n11404), .A2(n11400), .ZN(n11430) );
  AND2_X1 U12014 ( .A1(n13747), .A2(n9769), .ZN(n9904) );
  NAND2_X1 U12015 ( .A1(n11384), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11404) );
  NAND2_X1 U12016 ( .A1(n11369), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11368) );
  NOR2_X1 U12017 ( .A1(n11354), .A2(n11307), .ZN(n11369) );
  INV_X1 U12018 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11307) );
  AND2_X1 U12019 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n20596), .ZN(n13476) );
  INV_X1 U12020 ( .A(n14164), .ZN(n14153) );
  AND2_X1 U12021 ( .A1(n14272), .A2(n9812), .ZN(n14212) );
  INV_X1 U12022 ( .A(n14213), .ZN(n10101) );
  NAND2_X1 U12023 ( .A1(n14272), .A2(n10102), .ZN(n14222) );
  NAND2_X1 U12024 ( .A1(n14272), .A2(n14262), .ZN(n14261) );
  NOR2_X1 U12025 ( .A1(n14285), .A2(n14271), .ZN(n14272) );
  NAND2_X1 U12026 ( .A1(n10149), .A2(n10148), .ZN(n14558) );
  AOI21_X1 U12027 ( .B1(n11913), .B2(n10151), .A(n10150), .ZN(n10148) );
  NOR3_X1 U12028 ( .A1(n14566), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n9944) );
  INV_X1 U12029 ( .A(n14595), .ZN(n9945) );
  NAND2_X1 U12030 ( .A1(n14351), .A2(n9712), .ZN(n14300) );
  NAND2_X1 U12031 ( .A1(n14351), .A2(n10099), .ZN(n14325) );
  NAND2_X1 U12032 ( .A1(n14351), .A2(n14336), .ZN(n14337) );
  NAND2_X1 U12033 ( .A1(n14595), .A2(n14594), .ZN(n14593) );
  NAND2_X1 U12034 ( .A1(n14363), .A2(n9782), .ZN(n14411) );
  INV_X1 U12035 ( .A(n14413), .ZN(n10107) );
  NAND2_X1 U12036 ( .A1(n14363), .A2(n9760), .ZN(n14426) );
  NAND2_X1 U12037 ( .A1(n14363), .A2(n9764), .ZN(n14417) );
  AND2_X1 U12038 ( .A1(n14363), .A2(n14362), .ZN(n14424) );
  NOR2_X1 U12039 ( .A1(n13918), .A2(n13917), .ZN(n14363) );
  AOI21_X1 U12040 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n16174), .ZN(n14617) );
  OR2_X1 U12041 ( .A1(n13900), .A2(n13901), .ZN(n13918) );
  AND2_X1 U12042 ( .A1(n13724), .A2(n9711), .ZN(n16295) );
  AND2_X1 U12043 ( .A1(n10075), .A2(n11902), .ZN(n10074) );
  NAND2_X1 U12044 ( .A1(n16195), .A2(n10077), .ZN(n10076) );
  INV_X1 U12045 ( .A(n16287), .ZN(n16312) );
  NAND2_X1 U12046 ( .A1(n13724), .A2(n13723), .ZN(n13758) );
  NAND2_X1 U12047 ( .A1(n10073), .A2(n13461), .ZN(n10122) );
  NAND2_X1 U12048 ( .A1(n13373), .A2(n9819), .ZN(n13464) );
  INV_X1 U12049 ( .A(n16284), .ZN(n14764) );
  CLKBUF_X1 U12050 ( .A(n13083), .Z(n14795) );
  OR2_X1 U12051 ( .A1(n9673), .A2(n13420), .ZN(n20411) );
  NAND2_X1 U12052 ( .A1(n13387), .A2(n11842), .ZN(n20386) );
  AND2_X1 U12053 ( .A1(n9673), .A2(n13420), .ZN(n20559) );
  CLKBUF_X1 U12054 ( .A(n13419), .Z(n13420) );
  OR2_X1 U12055 ( .A1(n9673), .A2(n13781), .ZN(n20642) );
  INV_X1 U12056 ( .A(n20559), .ZN(n20385) );
  OR2_X1 U12057 ( .A1(n11842), .A2(n13390), .ZN(n20648) );
  CLKBUF_X1 U12058 ( .A(n10604), .Z(n10456) );
  AOI22_X1 U12059 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n20088), .B2(n13539), .ZN(
        n12747) );
  AND2_X1 U12060 ( .A1(n10536), .A2(n10523), .ZN(n12738) );
  NOR2_X1 U12061 ( .A1(n10326), .A2(n15273), .ZN(n10327) );
  NAND2_X1 U12062 ( .A1(n10327), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10328) );
  NAND2_X1 U12063 ( .A1(n12656), .A2(n9762), .ZN(n12631) );
  NAND2_X1 U12064 ( .A1(n10315), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10318) );
  AND2_X1 U12065 ( .A1(n12637), .A2(n12658), .ZN(n19232) );
  AND2_X1 U12066 ( .A1(n12621), .A2(n9714), .ZN(n12643) );
  NAND2_X1 U12067 ( .A1(n12621), .A2(n9706), .ZN(n12651) );
  NAND2_X1 U12068 ( .A1(n12621), .A2(n10587), .ZN(n12649) );
  NAND2_X1 U12069 ( .A1(n9709), .A2(n15115), .ZN(n10118) );
  AND2_X1 U12070 ( .A1(n13562), .A2(n13010), .ZN(n14917) );
  AND2_X1 U12071 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10303) );
  INV_X1 U12072 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14954) );
  AND2_X1 U12073 ( .A1(n10179), .A2(n12414), .ZN(n10178) );
  NOR2_X1 U12074 ( .A1(n10210), .A2(n10209), .ZN(n10208) );
  INV_X1 U12075 ( .A(n15129), .ZN(n10209) );
  NOR2_X1 U12076 ( .A1(n15158), .A2(n10210), .ZN(n15128) );
  NOR2_X1 U12077 ( .A1(n15158), .A2(n15145), .ZN(n15147) );
  NAND2_X1 U12078 ( .A1(n14988), .A2(n9744), .ZN(n10241) );
  INV_X1 U12079 ( .A(n12258), .ZN(n9832) );
  NAND2_X1 U12080 ( .A1(n14988), .A2(n12236), .ZN(n12259) );
  OR2_X1 U12081 ( .A1(n15005), .A2(n15016), .ZN(n10243) );
  NAND2_X1 U12082 ( .A1(n12167), .A2(n10244), .ZN(n9835) );
  INV_X1 U12083 ( .A(n15005), .ZN(n10244) );
  INV_X1 U12084 ( .A(n12167), .ZN(n10242) );
  AND2_X1 U12085 ( .A1(n10975), .A2(n10974), .ZN(n15172) );
  NAND2_X1 U12086 ( .A1(n10206), .A2(n10973), .ZN(n15173) );
  CLKBUF_X1 U12087 ( .A(n15019), .Z(n15020) );
  AND2_X1 U12088 ( .A1(n10970), .A2(n10969), .ZN(n15201) );
  CLKBUF_X1 U12089 ( .A(n15033), .Z(n15034) );
  AND3_X1 U12090 ( .A1(n10962), .A2(n10961), .A3(n10960), .ZN(n15242) );
  NOR2_X1 U12091 ( .A1(n10195), .A2(n10196), .ZN(n15241) );
  AND2_X1 U12092 ( .A1(n12229), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13310) );
  AND2_X1 U12093 ( .A1(n10602), .A2(n12329), .ZN(n12347) );
  NAND2_X1 U12094 ( .A1(n19357), .A2(n12369), .ZN(n13052) );
  AND2_X1 U12095 ( .A1(n13013), .A2(n20123), .ZN(n19391) );
  INV_X1 U12096 ( .A(n12363), .ZN(n15709) );
  OAI21_X1 U12097 ( .B1(n12362), .B2(n12361), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12363) );
  NAND2_X1 U12098 ( .A1(n10292), .A2(n9716), .ZN(n10325) );
  AND2_X1 U12099 ( .A1(n10292), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10324) );
  NAND2_X1 U12100 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n10320), .ZN(
        n10300) );
  AND2_X1 U12101 ( .A1(n10315), .A2(n10160), .ZN(n10320) );
  AND2_X1 U12102 ( .A1(n9707), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10160) );
  NAND2_X1 U12103 ( .A1(n10315), .A2(n9707), .ZN(n10321) );
  NOR2_X1 U12104 ( .A1(n9915), .A2(n9719), .ZN(n9914) );
  NOR2_X1 U12105 ( .A1(n10316), .A2(n19249), .ZN(n10315) );
  NAND2_X1 U12106 ( .A1(n10313), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10316) );
  NOR2_X1 U12107 ( .A1(n16458), .A2(n10314), .ZN(n10313) );
  NAND2_X1 U12108 ( .A1(n14855), .A2(n10727), .ZN(n15081) );
  AND2_X1 U12109 ( .A1(n10301), .A2(n9793), .ZN(n10310) );
  NOR2_X1 U12110 ( .A1(n14871), .A2(n14870), .ZN(n15103) );
  NAND2_X1 U12111 ( .A1(n10301), .A2(n9696), .ZN(n10311) );
  NAND2_X1 U12112 ( .A1(n10301), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10309) );
  AND2_X1 U12113 ( .A1(n10301), .A2(n10169), .ZN(n10308) );
  INV_X1 U12114 ( .A(n9915), .ZN(n9913) );
  NOR2_X1 U12115 ( .A1(n15411), .A2(n10304), .ZN(n10307) );
  AND2_X1 U12116 ( .A1(n13319), .A2(n13320), .ZN(n13444) );
  NAND2_X1 U12117 ( .A1(n10303), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10302) );
  NOR2_X1 U12118 ( .A1(n10302), .A2(n19439), .ZN(n10305) );
  NAND4_X1 U12119 ( .A1(n10653), .A2(n10664), .A3(n10663), .A4(n10662), .ZN(
        n12034) );
  NOR2_X1 U12120 ( .A1(n14087), .A2(n10214), .ZN(n10213) );
  NOR2_X1 U12121 ( .A1(n15257), .A2(n15292), .ZN(n10231) );
  NAND2_X1 U12122 ( .A1(n9753), .A2(n10027), .ZN(n15274) );
  NOR2_X1 U12123 ( .A1(n10141), .A2(n15507), .ZN(n10027) );
  NAND2_X1 U12124 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n12850), .ZN(
        n10141) );
  OR2_X1 U12125 ( .A1(n15011), .A2(n14998), .ZN(n15000) );
  NOR2_X1 U12126 ( .A1(n15000), .A2(n14990), .ZN(n14991) );
  AND2_X1 U12127 ( .A1(n15025), .A2(n14824), .ZN(n15009) );
  NAND2_X1 U12128 ( .A1(n15009), .A2(n15008), .ZN(n15011) );
  AOI21_X1 U12129 ( .B1(n9962), .B2(n9960), .A(n9959), .ZN(n9958) );
  INV_X1 U12130 ( .A(n9962), .ZN(n9961) );
  INV_X1 U12131 ( .A(n12684), .ZN(n9960) );
  AND2_X1 U12132 ( .A1(n10751), .A2(n10750), .ZN(n14837) );
  NAND2_X1 U12133 ( .A1(n15053), .A2(n10185), .ZN(n15038) );
  AND2_X1 U12134 ( .A1(n15053), .A2(n15044), .ZN(n15046) );
  NOR2_X1 U12135 ( .A1(n9705), .A2(n10193), .ZN(n10192) );
  INV_X1 U12136 ( .A(n15222), .ZN(n10193) );
  NAND2_X1 U12137 ( .A1(n10047), .A2(n10050), .ZN(n15365) );
  NAND2_X1 U12138 ( .A1(n10049), .A2(n10048), .ZN(n10047) );
  NAND2_X1 U12139 ( .A1(n10072), .A2(n10071), .ZN(n10070) );
  OR2_X1 U12140 ( .A1(n10201), .A2(n10200), .ZN(n10199) );
  INV_X1 U12141 ( .A(n13324), .ZN(n10200) );
  OR2_X1 U12142 ( .A1(n13181), .A2(n10202), .ZN(n16559) );
  AND2_X1 U12143 ( .A1(n10713), .A2(n10712), .ZN(n13586) );
  AND2_X1 U12144 ( .A1(n13444), .A2(n10186), .ZN(n13599) );
  AND2_X1 U12145 ( .A1(n13444), .A2(n13443), .ZN(n13458) );
  NAND2_X1 U12146 ( .A1(n13444), .A2(n10188), .ZN(n13585) );
  NAND2_X1 U12147 ( .A1(n13505), .A2(n10857), .ZN(n13049) );
  NAND2_X1 U12148 ( .A1(n12517), .A2(n12516), .ZN(n15417) );
  NAND2_X1 U12149 ( .A1(n9966), .A2(n9964), .ZN(n12517) );
  AOI21_X1 U12150 ( .B1(n9971), .B2(n9781), .A(n9968), .ZN(n9967) );
  AND2_X1 U12151 ( .A1(n9974), .A2(n9969), .ZN(n9968) );
  NOR2_X1 U12152 ( .A1(n9971), .A2(n9974), .ZN(n9970) );
  AND2_X1 U12153 ( .A1(n10842), .A2(n9755), .ZN(n10189) );
  AND2_X1 U12154 ( .A1(n10698), .A2(n10697), .ZN(n13311) );
  NOR2_X1 U12155 ( .A1(n13312), .A2(n13311), .ZN(n13319) );
  AND2_X2 U12157 ( .A1(n9839), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13536) );
  INV_X1 U12158 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9839) );
  AOI21_X1 U12159 ( .B1(n13059), .B2(n12039), .A(n12032), .ZN(n13046) );
  NAND2_X1 U12160 ( .A1(n13158), .A2(n10272), .ZN(n13267) );
  NAND2_X1 U12161 ( .A1(n12017), .A2(n9775), .ZN(n12019) );
  INV_X1 U12162 ( .A(n12018), .ZN(n9838) );
  NAND2_X1 U12163 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19919), .ZN(n19468) );
  OR2_X1 U12164 ( .A1(n19727), .A2(n15723), .ZN(n19836) );
  OR2_X1 U12165 ( .A1(n19727), .A2(n20093), .ZN(n19865) );
  INV_X1 U12166 ( .A(n19479), .ZN(n19481) );
  INV_X1 U12167 ( .A(n19468), .ZN(n19485) );
  NOR2_X1 U12168 ( .A1(n15707), .A2(n15708), .ZN(n19480) );
  INV_X1 U12169 ( .A(n12734), .ZN(n9851) );
  NAND2_X1 U12170 ( .A1(n9985), .A2(n17803), .ZN(n9990) );
  AND2_X1 U12171 ( .A1(n16885), .A2(n17816), .ZN(n16886) );
  NAND2_X1 U12172 ( .A1(n17882), .A2(n9765), .ZN(n16816) );
  NOR2_X1 U12173 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16930), .ZN(n16919) );
  NOR2_X1 U12174 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16952), .ZN(n16939) );
  NAND2_X1 U12175 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14035) );
  AOI21_X1 U12176 ( .B1(n18915), .B2(n18914), .A(n17699), .ZN(n17130) );
  INV_X1 U12177 ( .A(n17168), .ZN(n17190) );
  AOI21_X1 U12178 ( .B1(n17334), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A(
        n9874), .ZN(n17299) );
  AOI21_X1 U12179 ( .B1(n15756), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A(n9876), .ZN(n17321) );
  AND2_X1 U12180 ( .A1(n9872), .A2(n9871), .ZN(n17351) );
  NAND2_X1 U12181 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n9871) );
  AOI21_X1 U12182 ( .B1(n9656), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A(n9877), 
        .ZN(n17382) );
  NAND2_X1 U12183 ( .A1(n15929), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n9870) );
  NAND2_X1 U12184 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n9869) );
  NAND2_X1 U12185 ( .A1(n15936), .A2(n9863), .ZN(n9862) );
  AOI22_X1 U12186 ( .A1(n18922), .A2(n15983), .B1(n15831), .B2(n15830), .ZN(
        n16122) );
  AOI21_X1 U12187 ( .B1(n9658), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(n9875), 
        .ZN(n9996) );
  NAND2_X1 U12188 ( .A1(n9656), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n9995) );
  NAND2_X1 U12189 ( .A1(n17447), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10003) );
  NOR2_X1 U12190 ( .A1(n10000), .A2(n9999), .ZN(n9998) );
  NOR2_X1 U12191 ( .A1(n13974), .A2(n15962), .ZN(n9999) );
  AOI211_X1 U12192 ( .C1(n15864), .C2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n13980), .B(n13979), .ZN(n13981) );
  NOR2_X1 U12193 ( .A1(n17699), .A2(n17660), .ZN(n17679) );
  NOR2_X1 U12194 ( .A1(n17700), .A2(n17699), .ZN(n17701) );
  NOR2_X1 U12195 ( .A1(n16809), .A2(n16845), .ZN(n16639) );
  AND2_X1 U12196 ( .A1(n17882), .A2(n9794), .ZN(n17769) );
  INV_X1 U12197 ( .A(n17814), .ZN(n9992) );
  OAI21_X1 U12198 ( .B1(n18139), .B2(n17881), .A(n18819), .ZN(n17837) );
  INV_X1 U12199 ( .A(n16946), .ZN(n17850) );
  NAND2_X1 U12200 ( .A1(n17882), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17852) );
  NOR2_X1 U12201 ( .A1(n17893), .A2(n17894), .ZN(n17882) );
  NOR2_X1 U12202 ( .A1(n17934), .A2(n17935), .ZN(n17919) );
  NAND2_X1 U12203 ( .A1(n17964), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17934) );
  AND2_X1 U12204 ( .A1(n9976), .A2(n17018), .ZN(n17964) );
  NOR2_X1 U12205 ( .A1(n18075), .A2(n9977), .ZN(n9976) );
  NAND2_X1 U12206 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n9978), .ZN(
        n9977) );
  INV_X1 U12207 ( .A(n17987), .ZN(n9978) );
  NAND2_X1 U12208 ( .A1(n18046), .A2(n17018), .ZN(n17985) );
  INV_X1 U12209 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18022) );
  NAND2_X1 U12210 ( .A1(n15982), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18011) );
  NOR2_X1 U12211 ( .A1(n18075), .A2(n18082), .ZN(n18046) );
  NAND2_X1 U12212 ( .A1(n17789), .A2(n17776), .ZN(n16042) );
  INV_X1 U12213 ( .A(n16043), .ZN(n16669) );
  NOR2_X1 U12214 ( .A1(n18158), .A2(n17819), .ZN(n18154) );
  NAND2_X1 U12215 ( .A1(n17915), .A2(n16039), .ZN(n17841) );
  NOR2_X1 U12217 ( .A1(n17962), .A2(n17957), .ZN(n17956) );
  INV_X1 U12218 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17957) );
  NOR2_X1 U12219 ( .A1(n9767), .A2(n18017), .ZN(n17948) );
  NOR2_X1 U12220 ( .A1(n18300), .A2(n17970), .ZN(n17969) );
  NOR2_X1 U12221 ( .A1(n18309), .A2(n18292), .ZN(n17963) );
  NAND2_X1 U12222 ( .A1(n17963), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17962) );
  INV_X1 U12223 ( .A(n18011), .ZN(n18331) );
  NAND2_X1 U12224 ( .A1(n15872), .A2(n15871), .ZN(n16666) );
  NAND2_X1 U12225 ( .A1(n18011), .A2(n16033), .ZN(n18382) );
  INV_X1 U12226 ( .A(n18917), .ZN(n16780) );
  INV_X1 U12227 ( .A(n18078), .ZN(n9888) );
  NAND2_X1 U12228 ( .A1(n9868), .A2(n10004), .ZN(n18074) );
  INV_X1 U12229 ( .A(n10005), .ZN(n10004) );
  OAI22_X1 U12230 ( .A1(n10009), .A2(n10006), .B1(n10011), .B2(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10005) );
  NOR2_X1 U12231 ( .A1(n18095), .A2(n16007), .ZN(n18089) );
  INV_X1 U12232 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18436) );
  XNOR2_X1 U12233 ( .A(n15967), .B(n18436), .ZN(n18121) );
  INV_X1 U12234 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18978) );
  NOR2_X1 U12235 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18479), .ZN(n18766) );
  INV_X1 U12236 ( .A(n15883), .ZN(n18489) );
  NOR2_X1 U12237 ( .A1(n13958), .A2(n13957), .ZN(n18493) );
  NOR2_X1 U12238 ( .A1(n13947), .A2(n13946), .ZN(n18497) );
  NOR2_X1 U12239 ( .A1(n14003), .A2(n14002), .ZN(n18501) );
  NOR2_X1 U12240 ( .A1(n13993), .A2(n13992), .ZN(n18506) );
  INV_X1 U12241 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19095) );
  OR2_X1 U12242 ( .A1(n14250), .A2(n14183), .ZN(n14231) );
  INV_X1 U12243 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14328) );
  NOR2_X1 U12244 ( .A1(n16146), .A2(n14179), .ZN(n14331) );
  NOR2_X1 U12245 ( .A1(n16159), .A2(n14177), .ZN(n16147) );
  NOR2_X1 U12246 ( .A1(n20173), .A2(n13869), .ZN(n20158) );
  AND2_X1 U12247 ( .A1(n13669), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13648) );
  INV_X1 U12248 ( .A(n20196), .ZN(n20177) );
  NAND2_X1 U12249 ( .A1(n13763), .A2(n9826), .ZN(n14372) );
  AND2_X1 U12250 ( .A1(n13734), .A2(n13670), .ZN(n20197) );
  AND2_X1 U12251 ( .A1(n13734), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20196) );
  INV_X1 U12252 ( .A(n20183), .ZN(n20193) );
  NAND2_X1 U12253 ( .A1(n13734), .A2(n13736), .ZN(n20185) );
  NOR2_X1 U12254 ( .A1(n13373), .A2(n9820), .ZN(n13739) );
  AND2_X1 U12255 ( .A1(n20216), .A2(n13433), .ZN(n14430) );
  NAND2_X1 U12256 ( .A1(n13135), .A2(n13134), .ZN(n20216) );
  NAND2_X1 U12257 ( .A1(n13132), .A2(n9937), .ZN(n13135) );
  INV_X1 U12258 ( .A(n14430), .ZN(n20209) );
  INV_X1 U12259 ( .A(n11306), .ZN(n13433) );
  OAI21_X1 U12260 ( .B1(n9783), .B2(n14201), .A(n14200), .ZN(n14202) );
  INV_X1 U12261 ( .A(n14481), .ZN(n14490) );
  INV_X1 U12262 ( .A(n14437), .ZN(n14488) );
  INV_X1 U12263 ( .A(n14500), .ZN(n14503) );
  NAND2_X1 U12264 ( .A1(n12391), .A2(n12390), .ZN(n14498) );
  OR2_X1 U12265 ( .A1(n13133), .A2(n12954), .ZN(n12390) );
  NAND2_X1 U12266 ( .A1(n13101), .A2(n9937), .ZN(n12391) );
  OR2_X1 U12267 ( .A1(n14502), .A2(n13157), .ZN(n14500) );
  OAI21_X1 U12268 ( .B1(n13109), .B2(n13108), .A(n13107), .ZN(n20220) );
  AND2_X1 U12269 ( .A1(n13656), .A2(n20840), .ZN(n13020) );
  INV_X1 U12270 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14550) );
  CLKBUF_X1 U12271 ( .A(n14347), .Z(n14348) );
  INV_X1 U12272 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16210) );
  INV_X1 U12273 ( .A(n16209), .ZN(n16194) );
  NAND2_X1 U12274 ( .A1(n10251), .A2(n10252), .ZN(n13400) );
  OR3_X1 U12275 ( .A1(n14654), .A2(n14653), .A3(n14652), .ZN(n16230) );
  NAND2_X1 U12276 ( .A1(n10081), .A2(n16196), .ZN(n13860) );
  INV_X1 U12277 ( .A(n20282), .ZN(n16259) );
  NAND2_X1 U12278 ( .A1(n13238), .A2(n13231), .ZN(n14715) );
  INV_X1 U12279 ( .A(n16260), .ZN(n20285) );
  AND2_X2 U12280 ( .A1(n13238), .A2(n13230), .ZN(n20282) );
  INV_X1 U12281 ( .A(n20324), .ZN(n20347) );
  OR2_X1 U12282 ( .A1(n20386), .A2(n20525), .ZN(n20380) );
  INV_X1 U12283 ( .A(n20373), .ZN(n20375) );
  INV_X1 U12284 ( .A(n13691), .ZN(n13625) );
  OAI21_X1 U12285 ( .B1(n13479), .B2(n13478), .A(n20650), .ZN(n13699) );
  OAI211_X1 U12286 ( .C1(n20488), .C2(n20609), .A(n20473), .B(n20536), .ZN(
        n20491) );
  OAI211_X1 U12287 ( .C1(n20538), .C2(n20537), .A(n20536), .B(n20535), .ZN(
        n20555) );
  OAI21_X1 U12288 ( .B1(n20574), .B2(n20573), .A(n20572), .ZN(n20592) );
  OAI211_X1 U12289 ( .C1(n20724), .C2(n20687), .A(n20686), .B(n20685), .ZN(
        n20730) );
  INV_X1 U12290 ( .A(n20295), .ZN(n20745) );
  OR2_X1 U12291 ( .A1(n20648), .A2(n20385), .ZN(n20295) );
  INV_X1 U12292 ( .A(n20749), .ZN(n20682) );
  AND2_X1 U12293 ( .A1(n16085), .A2(n16084), .ZN(n16101) );
  NOR2_X1 U12294 ( .A1(n13219), .A2(n20609), .ZN(n16095) );
  INV_X1 U12295 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n16345) );
  INV_X1 U12296 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20609) );
  NOR2_X1 U12297 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20755), .ZN(n20817) );
  CLKBUF_X1 U12298 ( .A(n12346), .Z(n12883) );
  INV_X1 U12299 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19986) );
  NAND2_X1 U12300 ( .A1(n10639), .A2(n10641), .ZN(n20106) );
  NAND2_X1 U12301 ( .A1(n14809), .A2(n14808), .ZN(n10153) );
  NAND2_X1 U12302 ( .A1(n16365), .A2(n16366), .ZN(n16364) );
  NAND2_X1 U12303 ( .A1(n16377), .A2(n16378), .ZN(n16376) );
  NAND2_X1 U12304 ( .A1(n12704), .A2(n10592), .ZN(n12708) );
  NAND2_X1 U12305 ( .A1(n16399), .A2(n16400), .ZN(n16398) );
  NAND2_X1 U12306 ( .A1(n16410), .A2(n16411), .ZN(n16409) );
  NAND2_X1 U12307 ( .A1(n10173), .A2(n10171), .ZN(n19179) );
  NOR2_X1 U12308 ( .A1(n10174), .A2(n9700), .ZN(n10171) );
  AND2_X1 U12309 ( .A1(n20111), .A2(n10481), .ZN(n19324) );
  AND2_X1 U12310 ( .A1(n10121), .A2(n12612), .ZN(n14883) );
  AND2_X1 U12311 ( .A1(n12949), .A2(n13509), .ZN(n19327) );
  OR2_X1 U12312 ( .A1(n20111), .A2(n10459), .ZN(n19301) );
  INV_X1 U12313 ( .A(n19327), .ZN(n19320) );
  NAND2_X1 U12314 ( .A1(n14813), .A2(n14812), .ZN(n19326) );
  NAND2_X1 U12315 ( .A1(n20111), .A2(n10788), .ZN(n19321) );
  INV_X1 U12316 ( .A(n19308), .ZN(n19334) );
  OR2_X1 U12317 ( .A1(n10944), .A2(n10943), .ZN(n15084) );
  OR2_X1 U12318 ( .A1(n10800), .A2(n10799), .ZN(n15101) );
  OR2_X1 U12319 ( .A1(n10875), .A2(n10874), .ZN(n13589) );
  INV_X2 U12320 ( .A(n15116), .ZN(n15089) );
  INV_X1 U12321 ( .A(n15106), .ZN(n15109) );
  INV_X1 U12322 ( .A(n20082), .ZN(n15724) );
  INV_X1 U12323 ( .A(n20093), .ZN(n15723) );
  AND2_X2 U12324 ( .A1(n12412), .A2(n13010), .ZN(n15116) );
  OR2_X1 U12325 ( .A1(n15089), .A2(n12413), .ZN(n15106) );
  INV_X1 U12326 ( .A(n19358), .ZN(n19383) );
  INV_X1 U12327 ( .A(n19357), .ZN(n19382) );
  INV_X1 U12328 ( .A(n15230), .ZN(n19385) );
  AND2_X2 U12329 ( .A1(n19153), .A2(n13571), .ZN(n12949) );
  OAI21_X1 U12330 ( .B1(n10042), .B2(n10038), .A(n10037), .ZN(n10036) );
  NOR2_X1 U12331 ( .A1(n15342), .A2(n10039), .ZN(n10038) );
  NAND2_X1 U12332 ( .A1(n10042), .A2(n15341), .ZN(n10037) );
  NAND2_X1 U12333 ( .A1(n10062), .A2(n10066), .ZN(n16454) );
  NAND2_X1 U12334 ( .A1(n10072), .A2(n10068), .ZN(n10062) );
  INV_X1 U12335 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n15411) );
  INV_X1 U12336 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19439) );
  AND2_X1 U12337 ( .A1(n19438), .A2(n12965), .ZN(n19426) );
  CLKBUF_X1 U12338 ( .A(n13269), .Z(n13270) );
  INV_X1 U12339 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14943) );
  INV_X1 U12340 ( .A(n19426), .ZN(n16491) );
  OAI211_X1 U12341 ( .C1(n15443), .C2(n15434), .A(n9746), .B(n10021), .ZN(
        n9924) );
  NOR2_X1 U12342 ( .A1(n15435), .A2(n9736), .ZN(n10021) );
  NAND2_X1 U12343 ( .A1(n15481), .A2(n12793), .ZN(n15459) );
  INV_X1 U12344 ( .A(n15259), .ZN(n15281) );
  NAND2_X1 U12345 ( .A1(n12703), .A2(n12702), .ZN(n15294) );
  AND2_X1 U12346 ( .A1(n15513), .A2(n12791), .ZN(n15486) );
  NAND2_X1 U12347 ( .A1(n12692), .A2(n15317), .ZN(n15310) );
  NAND2_X1 U12348 ( .A1(n15523), .A2(n16526), .ZN(n15513) );
  NAND2_X1 U12349 ( .A1(n15053), .A2(n10183), .ZN(n15023) );
  OR2_X1 U12350 ( .A1(n9722), .A2(n10040), .ZN(n10034) );
  NAND2_X1 U12351 ( .A1(n15334), .A2(n15341), .ZN(n10040) );
  AND2_X1 U12352 ( .A1(n10042), .A2(n15342), .ZN(n10035) );
  AND2_X1 U12353 ( .A1(n10036), .A2(n16584), .ZN(n10033) );
  NAND2_X1 U12354 ( .A1(n9849), .A2(n12789), .ZN(n15553) );
  INV_X1 U12355 ( .A(n15559), .ZN(n9849) );
  NAND2_X1 U12356 ( .A1(n10053), .A2(n10057), .ZN(n15573) );
  NAND2_X1 U12357 ( .A1(n16437), .A2(n10058), .ZN(n10053) );
  AND2_X1 U12358 ( .A1(n15069), .A2(n15068), .ZN(n19238) );
  AND2_X1 U12359 ( .A1(n10223), .A2(n9739), .ZN(n16481) );
  NAND2_X1 U12360 ( .A1(n16562), .A2(n9745), .ZN(n16525) );
  NAND2_X1 U12361 ( .A1(n10133), .A2(n9726), .ZN(n15381) );
  CLKBUF_X1 U12362 ( .A(n15409), .Z(n15410) );
  NAND2_X1 U12363 ( .A1(n15668), .A2(n12833), .ZN(n15421) );
  OAI21_X1 U12364 ( .B1(n13702), .B2(n10861), .A(n14936), .ZN(n13705) );
  AND2_X1 U12365 ( .A1(n13023), .A2(n13024), .ZN(n9850) );
  OR2_X1 U12366 ( .A1(n12853), .A2(n12797), .ZN(n16563) );
  INV_X1 U12367 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15692) );
  INV_X1 U12368 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20088) );
  INV_X1 U12369 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20079) );
  NAND2_X1 U12370 ( .A1(n13035), .A2(n10842), .ZN(n13491) );
  OAI21_X1 U12371 ( .B1(n13046), .B2(n13045), .A(n13044), .ZN(n20082) );
  AND2_X1 U12372 ( .A1(n13158), .A2(n13161), .ZN(n19440) );
  INV_X1 U12373 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15859) );
  INV_X1 U12374 ( .A(n19970), .ZN(n19488) );
  AND2_X1 U12375 ( .A1(n19594), .A2(n19590), .ZN(n19599) );
  NOR2_X1 U12376 ( .A1(n19553), .A2(n19667), .ZN(n19595) );
  OAI21_X1 U12377 ( .B1(n19643), .B2(n19868), .A(n19642), .ZN(n19661) );
  AOI22_X1 U12378 ( .A1(n19705), .A2(n19704), .B1(n19703), .B2(n19702), .ZN(
        n19721) );
  INV_X1 U12379 ( .A(n19757), .ZN(n19743) );
  OAI21_X1 U12380 ( .B1(n19736), .B2(n19735), .A(n19734), .ZN(n19753) );
  NOR2_X1 U12381 ( .A1(n19836), .A2(n19728), .ZN(n19769) );
  NOR2_X1 U12382 ( .A1(n19865), .A2(n19553), .ZN(n19801) );
  NOR2_X1 U12383 ( .A1(n19836), .A2(n19553), .ZN(n19816) );
  INV_X1 U12384 ( .A(n19823), .ZN(n19862) );
  INV_X1 U12385 ( .A(n19930), .ZN(n19883) );
  INV_X1 U12386 ( .A(n19948), .ZN(n19892) );
  INV_X1 U12387 ( .A(n19954), .ZN(n19895) );
  INV_X1 U12388 ( .A(n19960), .ZN(n19898) );
  OAI21_X1 U12389 ( .B1(n19879), .B2(n19878), .A(n19877), .ZN(n19904) );
  INV_X1 U12390 ( .A(n19971), .ZN(n19903) );
  NOR2_X2 U12391 ( .A1(n19836), .A2(n19835), .ZN(n19902) );
  OAI22_X1 U12392 ( .A1(n16689), .A2(n19483), .B1(n18485), .B2(n19481), .ZN(
        n19927) );
  AND2_X1 U12393 ( .A1(n19459), .A2(n19485), .ZN(n19931) );
  OAI22_X1 U12394 ( .A1(n19464), .A2(n19483), .B1(n19463), .B2(n19481), .ZN(
        n19939) );
  OAI22_X1 U12395 ( .A1(n19473), .A2(n19483), .B1(n19472), .B2(n19481), .ZN(
        n19951) );
  AND2_X1 U12396 ( .A1(n10508), .A2(n19485), .ZN(n19949) );
  AND2_X1 U12397 ( .A1(n12012), .A2(n19485), .ZN(n19955) );
  OAI22_X1 U12398 ( .A1(n16682), .A2(n19483), .B1(n17512), .B2(n19481), .ZN(
        n19957) );
  NOR2_X2 U12399 ( .A1(n19865), .A2(n19864), .ZN(n19966) );
  OAI22_X1 U12400 ( .A1(n19484), .A2(n19483), .B1(n19482), .B2(n19481), .ZN(
        n19965) );
  AND2_X1 U12401 ( .A1(n19486), .A2(n19485), .ZN(n19962) );
  OR2_X1 U12402 ( .A1(n19980), .A2(n19591), .ZN(n16605) );
  NAND2_X1 U12403 ( .A1(n15682), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16602) );
  AND3_X1 U12404 ( .A1(n13582), .A2(n20110), .A3(n13581), .ZN(n19976) );
  NAND2_X1 U12405 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19986), .ZN(n20098) );
  XOR2_X1 U12406 ( .A(n19136), .B(n17661), .Z(n19148) );
  INV_X1 U12407 ( .A(n17130), .ZN(n19147) );
  NAND2_X1 U12408 ( .A1(n19131), .A2(n16780), .ZN(n17699) );
  INV_X1 U12409 ( .A(n9982), .ZN(n16857) );
  AND2_X1 U12410 ( .A1(n16864), .A2(n16822), .ZN(n16865) );
  NAND2_X1 U12411 ( .A1(n9989), .A2(n9990), .ZN(n16875) );
  AND2_X1 U12412 ( .A1(n16908), .A2(n16817), .ZN(n16909) );
  NAND2_X1 U12413 ( .A1(n9984), .A2(n9983), .ZN(n16920) );
  NAND2_X1 U12414 ( .A1(n9985), .A2(n9986), .ZN(n9983) );
  AND2_X1 U12415 ( .A1(n16927), .A2(n16815), .ZN(n16928) );
  NOR2_X1 U12416 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17099), .ZN(n17086) );
  INV_X1 U12417 ( .A(n17180), .ZN(n17145) );
  AND2_X1 U12418 ( .A1(n17261), .A2(n17201), .ZN(n17241) );
  NOR4_X2 U12419 ( .A1(n19136), .A2(n18482), .A3(n16122), .A4(n18983), .ZN(
        n17496) );
  INV_X1 U12420 ( .A(n17522), .ZN(n17519) );
  NOR2_X1 U12421 ( .A1(n17705), .A2(n17576), .ZN(n17577) );
  NOR2_X2 U12422 ( .A1(n17511), .A2(n17646), .ZN(n17584) );
  AND2_X1 U12423 ( .A1(n9870), .A2(n9869), .ZN(n17453) );
  NOR2_X1 U12424 ( .A1(n15910), .A2(n15909), .ZN(n17642) );
  INV_X1 U12425 ( .A(n17655), .ZN(n17648) );
  NOR3_X1 U12426 ( .A1(n15924), .A2(n15923), .A3(n15922), .ZN(n15925) );
  INV_X1 U12427 ( .A(n15919), .ZN(n15923) );
  NOR2_X2 U12428 ( .A1(n13970), .A2(n13969), .ZN(n18512) );
  NOR2_X1 U12429 ( .A1(n19133), .A2(n17679), .ZN(n17676) );
  CLKBUF_X1 U12430 ( .A(n17676), .Z(n17695) );
  OAI21_X1 U12431 ( .B1(n19136), .B2(n19137), .A(n17701), .ZN(n17758) );
  NOR2_X1 U12432 ( .A1(n19136), .A2(n17764), .ZN(n17761) );
  BUF_X1 U12433 ( .A(n17758), .Z(n17764) );
  INV_X1 U12435 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17773) );
  INV_X1 U12436 ( .A(n17980), .ZN(n17996) );
  NAND2_X1 U12437 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17969), .ZN(
        n18277) );
  NOR2_X1 U12438 ( .A1(n19095), .A2(n18071), .ZN(n17980) );
  INV_X1 U12439 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n18009) );
  INV_X1 U12440 ( .A(n18819), .ZN(n18858) );
  NOR2_X1 U12441 ( .A1(n18102), .A2(n18104), .ZN(n18083) );
  NOR2_X1 U12442 ( .A1(n17920), .A2(n17980), .ZN(n18126) );
  INV_X1 U12443 ( .A(n18126), .ZN(n18135) );
  NAND2_X1 U12444 ( .A1(n17888), .A2(n16038), .ZN(n17831) );
  AOI22_X1 U12445 ( .A1(n18286), .A2(n18317), .B1(n18278), .B2(n18277), .ZN(
        n18266) );
  INV_X1 U12446 ( .A(n17956), .ZN(n18286) );
  OAI21_X2 U12447 ( .B1(n18934), .B2(n15987), .A(n18933), .ZN(n18951) );
  INV_X1 U12448 ( .A(n10154), .ZN(n18066) );
  NAND2_X1 U12449 ( .A1(n9805), .A2(n18085), .ZN(n18084) );
  INV_X1 U12450 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18430) );
  NAND2_X1 U12451 ( .A1(n15983), .A2(n19148), .ZN(n18949) );
  INV_X1 U12452 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18957) );
  INV_X1 U12453 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18964) );
  INV_X1 U12454 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18968) );
  INV_X1 U12455 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n19092) );
  AOI211_X2 U12456 ( .C1(n19131), .C2(n18950), .A(n18481), .B(n14065), .ZN(
        n19116) );
  INV_X1 U12457 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19086) );
  INV_X1 U12458 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n19007) );
  NOR2_X1 U12460 ( .A1(n10266), .A2(n10265), .ZN(n10264) );
  INV_X1 U12461 ( .A(n9783), .ZN(n10266) );
  INV_X1 U12462 ( .A(n12868), .ZN(n10265) );
  OAI21_X1 U12463 ( .B1(n14668), .B2(n20135), .A(n10145), .ZN(P1_U2968) );
  INV_X1 U12464 ( .A(n10146), .ZN(n10145) );
  OAI21_X1 U12465 ( .B1(n14186), .B2(n14551), .A(n11989), .ZN(n10146) );
  OAI21_X1 U12466 ( .B1(n14677), .B2(n20135), .A(n11997), .ZN(P1_U2969) );
  OAI21_X1 U12467 ( .B1(n14696), .B2(n20135), .A(n10130), .ZN(P1_U2971) );
  OAI21_X1 U12468 ( .B1(n14704), .B2(n20135), .A(n12010), .ZN(P1_U2972) );
  NOR2_X1 U12469 ( .A1(n12009), .A2(n12008), .ZN(n12010) );
  AND2_X1 U12470 ( .A1(n12371), .A2(n12370), .ZN(n12372) );
  INV_X1 U12471 ( .A(n14099), .ZN(n14100) );
  AOI21_X1 U12472 ( .B1(n14807), .B2(n19435), .A(n12863), .ZN(n12866) );
  INV_X1 U12473 ( .A(n9925), .ZN(n15436) );
  AOI21_X1 U12474 ( .B1(n15268), .B2(n16496), .A(n15267), .ZN(n15269) );
  AOI21_X1 U12475 ( .B1(n16363), .B2(n19435), .A(n15265), .ZN(n15266) );
  OAI21_X1 U12476 ( .B1(n15277), .B2(n15463), .A(n10135), .ZN(P2_U2987) );
  AOI21_X1 U12477 ( .B1(n10140), .B2(n10139), .A(n10136), .ZN(n10135) );
  NAND2_X1 U12478 ( .A1(n10138), .A2(n10137), .ZN(n10136) );
  AND2_X1 U12479 ( .A1(n14110), .A2(n14109), .ZN(n14111) );
  NOR2_X1 U12480 ( .A1(n12813), .A2(n10276), .ZN(n12854) );
  OAI21_X1 U12481 ( .B1(n15437), .B2(n16570), .A(n10191), .ZN(P2_U3017) );
  INV_X1 U12482 ( .A(n9922), .ZN(n10191) );
  OAI21_X1 U12483 ( .B1(n9925), .B2(n16587), .A(n9923), .ZN(n9922) );
  INV_X1 U12484 ( .A(n9924), .ZN(n9923) );
  OR2_X1 U12485 ( .A1(n16849), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n9975) );
  AOI21_X1 U12486 ( .B1(n16645), .B2(n18041), .A(n10164), .ZN(n16650) );
  OAI211_X1 U12487 ( .C1(n16647), .C2(n16646), .A(n10166), .B(n10165), .ZN(
        n10164) );
  NAND2_X1 U12488 ( .A1(n16649), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10165) );
  AOI21_X1 U12489 ( .B1(n10018), .B2(n10017), .A(n10015), .ZN(n16676) );
  NAND2_X1 U12490 ( .A1(n9880), .A2(n9878), .ZN(n18212) );
  NOR2_X1 U12491 ( .A1(n9879), .A2(n18459), .ZN(n9878) );
  NAND2_X1 U12492 ( .A1(n12001), .A2(n10264), .ZN(n14200) );
  AND2_X1 U12493 ( .A1(n14991), .A2(n9717), .ZN(n9685) );
  NAND2_X1 U12494 ( .A1(n12733), .A2(n20116), .ZN(n10608) );
  AND2_X1 U12495 ( .A1(n14258), .A2(n9763), .ZN(n9686) );
  NOR2_X1 U12496 ( .A1(n14297), .A2(n14309), .ZN(n9687) );
  AND3_X1 U12497 ( .A1(n9993), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n9688) );
  NOR2_X2 U12498 ( .A1(n13941), .A2(n17178), .ZN(n15756) );
  NOR2_X1 U12499 ( .A1(n10259), .A2(n10257), .ZN(n14407) );
  AND2_X1 U12500 ( .A1(n14605), .A2(n14603), .ZN(n9689) );
  AND2_X1 U12501 ( .A1(n14272), .A2(n9803), .ZN(n9690) );
  NAND2_X1 U12502 ( .A1(n15283), .A2(n9823), .ZN(n14093) );
  NAND2_X1 U12503 ( .A1(n14258), .A2(n9761), .ZN(n14235) );
  NAND2_X1 U12504 ( .A1(n9653), .A2(n10236), .ZN(n15321) );
  NOR2_X1 U12505 ( .A1(n10259), .A2(n10260), .ZN(n14359) );
  NOR2_X1 U12506 ( .A1(n14334), .A2(n14335), .ZN(n14319) );
  AND3_X1 U12507 ( .A1(n11010), .A2(n11011), .A3(n11013), .ZN(n9691) );
  AND2_X1 U12508 ( .A1(n9938), .A2(n9937), .ZN(n9692) );
  OR2_X1 U12509 ( .A1(n11270), .A2(n11846), .ZN(n9693) );
  INV_X1 U12510 ( .A(n16174), .ZN(n16173) );
  NAND3_X1 U12511 ( .A1(n9835), .A2(n9811), .A3(n9834), .ZN(n9833) );
  AND2_X1 U12512 ( .A1(n12626), .A2(n10069), .ZN(n9694) );
  OR2_X1 U12513 ( .A1(n15981), .A2(n15980), .ZN(n9695) );
  AND2_X1 U12514 ( .A1(n10169), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n9696) );
  XNOR2_X1 U12515 ( .A(n9833), .B(n12215), .ZN(n14995) );
  XNOR2_X1 U12516 ( .A(n12233), .B(n12234), .ZN(n14987) );
  AND2_X1 U12517 ( .A1(n10242), .A2(n10245), .ZN(n15003) );
  INV_X1 U12518 ( .A(n10142), .ZN(n15301) );
  AND2_X1 U12519 ( .A1(n12598), .A2(n9779), .ZN(n9697) );
  AND2_X1 U12520 ( .A1(n9689), .A2(n10089), .ZN(n9698) );
  NOR2_X1 U12521 ( .A1(n16674), .A2(n16673), .ZN(n9699) );
  NOR2_X1 U12522 ( .A1(n19180), .A2(n19186), .ZN(n9700) );
  AND2_X1 U12523 ( .A1(n10060), .A2(n16435), .ZN(n9701) );
  AND2_X1 U12524 ( .A1(n13071), .A2(n9676), .ZN(n9702) );
  OR2_X1 U12525 ( .A1(n9694), .A2(n10067), .ZN(n10066) );
  AND2_X1 U12526 ( .A1(n15092), .A2(n12054), .ZN(n9703) );
  AND2_X1 U12527 ( .A1(n9813), .A2(n13035), .ZN(n13493) );
  AND2_X1 U12528 ( .A1(n9703), .A2(n9771), .ZN(n15042) );
  AND2_X1 U12529 ( .A1(n13633), .A2(n13747), .ZN(n9704) );
  OR2_X1 U12530 ( .A1(n10196), .A2(n10194), .ZN(n9705) );
  AND2_X1 U12531 ( .A1(n10587), .A2(n10117), .ZN(n9706) );
  NOR2_X1 U12532 ( .A1(n10195), .A2(n9705), .ZN(n15221) );
  AND2_X1 U12533 ( .A1(n10161), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9707) );
  INV_X1 U12534 ( .A(n10198), .ZN(n13274) );
  AND2_X1 U12535 ( .A1(n13310), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n9708) );
  AND2_X1 U12536 ( .A1(n10586), .A2(n10119), .ZN(n9709) );
  AND2_X1 U12537 ( .A1(n10973), .A2(n10205), .ZN(n9710) );
  AND2_X1 U12538 ( .A1(n10095), .A2(n9777), .ZN(n9711) );
  AND2_X1 U12539 ( .A1(n10097), .A2(n14298), .ZN(n9712) );
  INV_X1 U12540 ( .A(n10052), .ZN(n10048) );
  NAND2_X1 U12541 ( .A1(n10057), .A2(n15572), .ZN(n10052) );
  AND2_X1 U12542 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n9713)
         );
  AND2_X1 U12543 ( .A1(n9706), .A2(n9804), .ZN(n9714) );
  AND2_X1 U12544 ( .A1(n12052), .A2(n10247), .ZN(n9715) );
  NAND2_X1 U12545 ( .A1(n10246), .A2(n10247), .ZN(n13588) );
  NAND2_X1 U12546 ( .A1(n13308), .A2(n13310), .ZN(n13309) );
  OR2_X1 U12547 ( .A1(n12853), .A2(n12812), .ZN(n16574) );
  INV_X1 U12548 ( .A(n16574), .ZN(n16592) );
  AND2_X1 U12549 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n9716) );
  AND2_X1 U12550 ( .A1(n14982), .A2(n10181), .ZN(n9717) );
  AND2_X1 U12551 ( .A1(n9716), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9718) );
  NAND2_X1 U12552 ( .A1(n10238), .A2(n12849), .ZN(n9719) );
  AND2_X1 U12553 ( .A1(n10236), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9720) );
  INV_X2 U12554 ( .A(n10679), .ZN(n10784) );
  OR2_X1 U12555 ( .A1(n19486), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n9721) );
  NAND2_X1 U12556 ( .A1(n15622), .A2(n10238), .ZN(n15377) );
  AND2_X2 U12557 ( .A1(n12309), .A2(n10489), .ZN(n10501) );
  AND2_X1 U12558 ( .A1(n10043), .A2(n10044), .ZN(n9722) );
  NOR2_X1 U12559 ( .A1(n10142), .A2(n10218), .ZN(n15283) );
  AND3_X1 U12560 ( .A1(n15964), .A2(n9996), .A3(n9995), .ZN(n9723) );
  NAND2_X1 U12561 ( .A1(n15622), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15592) );
  OR2_X1 U12562 ( .A1(n15274), .A2(n15430), .ZN(n9724) );
  OR2_X1 U12563 ( .A1(n14307), .A2(n14309), .ZN(n14295) );
  NAND2_X1 U12564 ( .A1(n14258), .A2(n14260), .ZN(n14244) );
  OR2_X1 U12565 ( .A1(n14334), .A2(n9908), .ZN(n14307) );
  NAND2_X1 U12566 ( .A1(n14991), .A2(n10179), .ZN(n9725) );
  NOR2_X1 U12567 ( .A1(n15345), .A2(n15536), .ZN(n15337) );
  NOR2_X1 U12568 ( .A1(n14280), .A2(n14282), .ZN(n14268) );
  INV_X1 U12569 ( .A(n9938), .ZN(n13219) );
  NAND2_X1 U12570 ( .A1(n11978), .A2(n11979), .ZN(n9938) );
  OR2_X1 U12571 ( .A1(n10239), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9726) );
  INV_X1 U12572 ( .A(n10152), .ZN(n10151) );
  NAND2_X1 U12573 ( .A1(n14594), .A2(n9818), .ZN(n10152) );
  INV_X1 U12574 ( .A(n11345), .ZN(n10085) );
  AND2_X1 U12575 ( .A1(n10206), .A2(n9710), .ZN(n9727) );
  NAND2_X1 U12576 ( .A1(n12980), .A2(n13269), .ZN(n12449) );
  INV_X1 U12577 ( .A(n9910), .ZN(n12001) );
  NAND2_X1 U12578 ( .A1(n14258), .A2(n9776), .ZN(n9910) );
  AND3_X1 U12579 ( .A1(n14834), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n12843), .ZN(n9728) );
  OR2_X1 U12580 ( .A1(n12865), .A2(n19429), .ZN(n9729) );
  OR2_X1 U12581 ( .A1(n12865), .A2(n16587), .ZN(n9730) );
  INV_X1 U12582 ( .A(n12436), .ZN(n12424) );
  NAND2_X1 U12583 ( .A1(n10223), .A2(n12609), .ZN(n15630) );
  AND2_X1 U12584 ( .A1(n12833), .A2(n10237), .ZN(n9731) );
  NAND2_X1 U12585 ( .A1(n10070), .A2(n12626), .ZN(n15616) );
  NAND2_X1 U12586 ( .A1(n12733), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10643) );
  AND3_X1 U12587 ( .A1(n14818), .A2(n10861), .A3(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n9732) );
  INV_X2 U12588 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10489) );
  AND2_X1 U12589 ( .A1(n12555), .A2(n12554), .ZN(n9733) );
  AND2_X1 U12590 ( .A1(n15279), .A2(n12806), .ZN(n9734) );
  INV_X1 U12591 ( .A(n17654), .ZN(n15995) );
  INV_X1 U12592 ( .A(n19668), .ZN(n12518) );
  OR2_X1 U12593 ( .A1(n15396), .A2(n16558), .ZN(n9735) );
  AOI21_X1 U12594 ( .B1(n10676), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10678), .ZN(n12020) );
  OR3_X1 U12595 ( .A1(n9862), .A2(n15934), .A3(n15935), .ZN(n15988) );
  INV_X1 U12596 ( .A(n15988), .ZN(n17647) );
  AND2_X1 U12597 ( .A1(n16349), .A2(n16582), .ZN(n9736) );
  OR2_X1 U12598 ( .A1(n16012), .A2(n16013), .ZN(n9738) );
  NAND2_X1 U12599 ( .A1(n14987), .A2(n14989), .ZN(n14988) );
  NOR2_X1 U12600 ( .A1(n10225), .A2(n15632), .ZN(n9739) );
  XNOR2_X1 U12601 ( .A(n11895), .B(n11383), .ZN(n11883) );
  AND4_X1 U12602 ( .A1(n11033), .A2(n11032), .A3(n11031), .A4(n11030), .ZN(
        n9740) );
  OR2_X1 U12603 ( .A1(n17178), .A2(n9994), .ZN(n13959) );
  AND2_X1 U12604 ( .A1(n10601), .A2(n10647), .ZN(n9741) );
  INV_X1 U12605 ( .A(n10072), .ZN(n16465) );
  INV_X1 U12606 ( .A(n15292), .ZN(n10232) );
  AND2_X1 U12607 ( .A1(n11191), .A2(n9693), .ZN(n9742) );
  NOR2_X1 U12608 ( .A1(n16041), .A2(n16040), .ZN(n9743) );
  AND2_X1 U12609 ( .A1(n12236), .A2(n9832), .ZN(n9744) );
  AND2_X1 U12610 ( .A1(n12786), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9745) );
  INV_X1 U12611 ( .A(n9912), .ZN(n15622) );
  NAND2_X1 U12612 ( .A1(n9916), .A2(n9913), .ZN(n9912) );
  NOR2_X1 U12613 ( .A1(n15432), .A2(n15433), .ZN(n9746) );
  INV_X1 U12614 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n19102) );
  NAND2_X1 U12615 ( .A1(n12334), .A2(n13014), .ZN(n9747) );
  OAI21_X1 U12616 ( .B1(n12685), .B2(n9961), .A(n9958), .ZN(n15303) );
  AND2_X1 U12617 ( .A1(n10133), .A2(n10131), .ZN(n9748) );
  AND2_X1 U12618 ( .A1(n9930), .A2(n9929), .ZN(n9749) );
  NOR2_X1 U12619 ( .A1(n15192), .A2(n10204), .ZN(n14826) );
  AND2_X1 U12620 ( .A1(n9930), .A2(n11949), .ZN(n9750) );
  OR2_X1 U12621 ( .A1(n16669), .A2(n10287), .ZN(n9751) );
  AND2_X1 U12622 ( .A1(n9653), .A2(n9720), .ZN(n9753) );
  NAND2_X1 U12623 ( .A1(n14996), .A2(n12216), .ZN(n12233) );
  INV_X1 U12624 ( .A(n9665), .ZN(n13482) );
  NAND2_X1 U12625 ( .A1(n10154), .A2(n10012), .ZN(n16033) );
  OR2_X1 U12626 ( .A1(n9889), .A2(n16009), .ZN(n9754) );
  AND2_X1 U12627 ( .A1(n12019), .A2(n12049), .ZN(n13266) );
  INV_X1 U12628 ( .A(n9847), .ZN(n16562) );
  OR2_X1 U12629 ( .A1(n15652), .A2(n15647), .ZN(n9847) );
  AND2_X1 U12630 ( .A1(n10190), .A2(n13499), .ZN(n9755) );
  AND2_X1 U12631 ( .A1(n10186), .A2(n13598), .ZN(n9756) );
  NOR2_X1 U12632 ( .A1(n14604), .A2(n11909), .ZN(n9757) );
  AND2_X1 U12633 ( .A1(n10241), .A2(n14973), .ZN(n9758) );
  AND2_X1 U12634 ( .A1(n13633), .A2(n9904), .ZN(n13854) );
  NAND2_X1 U12635 ( .A1(n9703), .A2(n10250), .ZN(n15049) );
  NAND2_X1 U12636 ( .A1(n15224), .A2(n15213), .ZN(n15199) );
  AOI21_X1 U12637 ( .B1(n11312), .B2(n11495), .A(n11311), .ZN(n13631) );
  AND2_X1 U12638 ( .A1(n10315), .A2(n10161), .ZN(n9759) );
  AND2_X1 U12639 ( .A1(n14362), .A2(n14423), .ZN(n9760) );
  AND2_X1 U12640 ( .A1(n11707), .A2(n14260), .ZN(n9761) );
  AND2_X1 U12641 ( .A1(n12639), .A2(n19181), .ZN(n9762) );
  AND2_X1 U12642 ( .A1(n9761), .A2(n10255), .ZN(n9763) );
  AND2_X1 U12643 ( .A1(n9760), .A2(n10108), .ZN(n9764) );
  AND2_X1 U12644 ( .A1(n9688), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9765) );
  NAND2_X1 U12645 ( .A1(n17925), .A2(n18050), .ZN(n17888) );
  NOR2_X1 U12646 ( .A1(n14859), .A2(n14860), .ZN(n14858) );
  AND2_X1 U12647 ( .A1(n9703), .A2(n12055), .ZN(n15056) );
  AND2_X1 U12648 ( .A1(n14855), .A2(n10176), .ZN(n9766) );
  INV_X1 U12649 ( .A(n15341), .ZN(n10039) );
  INV_X1 U12650 ( .A(n14936), .ZN(n9969) );
  AND3_X1 U12651 ( .A1(n18011), .A2(n17952), .A3(n16033), .ZN(n9767) );
  OAI21_X1 U12652 ( .B1(n13702), .B2(n9970), .A(n9967), .ZN(n15671) );
  AND2_X1 U12653 ( .A1(n17952), .A2(n18272), .ZN(n9768) );
  NAND2_X1 U12654 ( .A1(n12841), .A2(n15406), .ZN(n15395) );
  NOR2_X1 U12655 ( .A1(n13853), .A2(n10254), .ZN(n9769) );
  AND2_X1 U12656 ( .A1(n14351), .A2(n10097), .ZN(n9770) );
  NAND2_X1 U12657 ( .A1(n15669), .A2(n15676), .ZN(n15668) );
  AND2_X1 U12658 ( .A1(n10250), .A2(n10249), .ZN(n9771) );
  AND2_X1 U12659 ( .A1(n9979), .A2(n9981), .ZN(n9772) );
  NAND2_X1 U12660 ( .A1(n9834), .A2(n9835), .ZN(n15004) );
  NOR2_X1 U12661 ( .A1(n16886), .A2(n9985), .ZN(n9773) );
  NOR2_X1 U12662 ( .A1(n13181), .A2(n13180), .ZN(n9774) );
  AND2_X1 U12663 ( .A1(n9838), .A2(n12016), .ZN(n9775) );
  AND2_X1 U12664 ( .A1(n9763), .A2(n12002), .ZN(n9776) );
  AND2_X1 U12665 ( .A1(n16293), .A2(n16294), .ZN(n9777) );
  OR2_X1 U12666 ( .A1(n11974), .A2(n11973), .ZN(n9778) );
  OR2_X1 U12667 ( .A1(n13181), .A2(n10201), .ZN(n10198) );
  AND2_X1 U12668 ( .A1(n15386), .A2(n15399), .ZN(n9779) );
  NAND2_X1 U12669 ( .A1(n10120), .A2(n9709), .ZN(n10121) );
  AND2_X1 U12670 ( .A1(n12790), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9780) );
  OR2_X1 U12671 ( .A1(n9969), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9781) );
  AND2_X1 U12672 ( .A1(n9764), .A2(n10107), .ZN(n9782) );
  AND2_X1 U12673 ( .A1(n11797), .A2(n11796), .ZN(n9783) );
  NOR2_X1 U12674 ( .A1(n11270), .A2(n11259), .ZN(n9784) );
  OR2_X1 U12675 ( .A1(n12876), .A2(n12875), .ZN(n9785) );
  NAND2_X1 U12676 ( .A1(n15354), .A2(n15363), .ZN(n9786) );
  INV_X1 U12677 ( .A(n15334), .ZN(n10042) );
  INV_X1 U12678 ( .A(n15617), .ZN(n10067) );
  OR2_X1 U12679 ( .A1(n10059), .A2(n15332), .ZN(n10057) );
  AND2_X1 U12680 ( .A1(n11304), .A2(n11303), .ZN(n9787) );
  AND2_X1 U12681 ( .A1(n9769), .A2(n13867), .ZN(n9788) );
  AND2_X1 U12682 ( .A1(n14788), .A2(n9900), .ZN(n9789) );
  AND2_X1 U12683 ( .A1(n9982), .A2(n17786), .ZN(n9790) );
  AND2_X1 U12684 ( .A1(n12554), .A2(n12827), .ZN(n9791) );
  AND2_X1 U12685 ( .A1(n10183), .A2(n10182), .ZN(n9792) );
  AND2_X1 U12686 ( .A1(n9696), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9793) );
  AND2_X1 U12687 ( .A1(n9765), .A2(n9992), .ZN(n9794) );
  AND2_X1 U12688 ( .A1(n9714), .A2(n12642), .ZN(n9795) );
  AND2_X1 U12689 ( .A1(n10175), .A2(n15067), .ZN(n9796) );
  AND2_X1 U12690 ( .A1(n9986), .A2(n16815), .ZN(n9797) );
  AND2_X1 U12691 ( .A1(n9762), .A2(n14844), .ZN(n9798) );
  AND2_X1 U12692 ( .A1(n10050), .A2(n10046), .ZN(n10045) );
  INV_X1 U12693 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20846) );
  INV_X2 U12694 ( .A(n19144), .ZN(n19127) );
  OR2_X1 U12695 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n9799) );
  INV_X1 U12696 ( .A(n16570), .ZN(n16584) );
  AND2_X1 U12697 ( .A1(n13724), .A2(n10095), .ZN(n9800) );
  AOI21_X2 U12698 ( .B1(n15889), .B2(n15888), .A(n18983), .ZN(n18391) );
  INV_X1 U12699 ( .A(n18391), .ZN(n18459) );
  AND2_X1 U12700 ( .A1(n10327), .A2(n10156), .ZN(n9801) );
  NOR2_X1 U12701 ( .A1(n17146), .A2(n16812), .ZN(n16937) );
  NAND2_X1 U12702 ( .A1(n13308), .A2(n9708), .ZN(n13317) );
  INV_X1 U12703 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10170) );
  AND2_X1 U12704 ( .A1(n10292), .A2(n9718), .ZN(n9802) );
  NOR2_X1 U12705 ( .A1(n14247), .A2(n10104), .ZN(n9803) );
  AND2_X1 U12706 ( .A1(n17882), .A2(n9688), .ZN(n16619) );
  OR2_X1 U12707 ( .A1(n10508), .A2(n10729), .ZN(n9804) );
  NAND2_X1 U12708 ( .A1(n10124), .A2(n10126), .ZN(n13209) );
  NOR2_X1 U12709 ( .A1(n18098), .A2(n15975), .ZN(n9805) );
  AND2_X1 U12710 ( .A1(n18243), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9806) );
  NAND2_X1 U12711 ( .A1(n13265), .A2(n12050), .ZN(n13308) );
  OR2_X1 U12712 ( .A1(n14410), .A2(n14418), .ZN(n9807) );
  OR2_X1 U12713 ( .A1(n9981), .A2(n16844), .ZN(n9808) );
  OR2_X1 U12714 ( .A1(n20751), .A2(n20846), .ZN(n16100) );
  INV_X1 U12715 ( .A(n16100), .ZN(n9937) );
  NOR2_X1 U12716 ( .A1(n13446), .A2(n12051), .ZN(n13587) );
  AND2_X1 U12717 ( .A1(n9859), .A2(n18050), .ZN(n9809) );
  INV_X1 U12718 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11006) );
  INV_X1 U12719 ( .A(n17146), .ZN(n17133) );
  OR2_X1 U12720 ( .A1(n10105), .A2(n10106), .ZN(n9810) );
  OR2_X1 U12721 ( .A1(n10270), .A2(n12188), .ZN(n9811) );
  INV_X1 U12722 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11005) );
  AND2_X1 U12723 ( .A1(n10102), .A2(n10101), .ZN(n9812) );
  AND2_X1 U12724 ( .A1(n10842), .A2(n10190), .ZN(n9813) );
  NOR2_X1 U12725 ( .A1(n16928), .A2(n9985), .ZN(n9814) );
  AND2_X1 U12726 ( .A1(n16823), .A2(n17786), .ZN(n9815) );
  AND2_X1 U12727 ( .A1(n9718), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9816) );
  INV_X1 U12728 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n19197) );
  INV_X1 U12729 ( .A(n14438), .ZN(n13418) );
  AND2_X2 U12730 ( .A1(n12401), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14438)
         );
  NOR2_X1 U12731 ( .A1(n17957), .A2(n18274), .ZN(n18243) );
  INV_X1 U12732 ( .A(n18243), .ZN(n9856) );
  INV_X1 U12733 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10162) );
  NOR2_X1 U12734 ( .A1(n13080), .A2(n13212), .ZN(n13225) );
  INV_X1 U12735 ( .A(n14965), .ZN(n10180) );
  AND2_X1 U12736 ( .A1(n10115), .A2(n10114), .ZN(n9817) );
  INV_X1 U12737 ( .A(n14421), .ZN(n10258) );
  AND2_X1 U12738 ( .A1(n14656), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9818) );
  AND2_X1 U12739 ( .A1(n13372), .A2(n13371), .ZN(n9819) );
  AND2_X1 U12740 ( .A1(n13300), .A2(n13299), .ZN(n9820) );
  INV_X1 U12741 ( .A(n10174), .ZN(n10172) );
  AND2_X1 U12742 ( .A1(n10291), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10174) );
  AND2_X1 U12743 ( .A1(n10156), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9821) );
  AND2_X1 U12744 ( .A1(n14181), .A2(n14180), .ZN(n9822) );
  AND2_X1 U12745 ( .A1(n10240), .A2(n12850), .ZN(n9823) );
  AND2_X1 U12746 ( .A1(n9720), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9824) );
  AND2_X1 U12747 ( .A1(n9822), .A2(n14182), .ZN(n9825) );
  AND2_X1 U12748 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .ZN(n9826) );
  OR2_X1 U12749 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n9827) );
  INV_X1 U12750 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n10116) );
  INV_X1 U12751 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10013) );
  INV_X1 U12752 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10218) );
  INV_X1 U12753 ( .A(n17853), .ZN(n9993) );
  INV_X1 U12754 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10157) );
  INV_X1 U12755 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10159) );
  INV_X1 U12756 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10163) );
  INV_X1 U12757 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10010) );
  INV_X1 U12758 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10168) );
  INV_X1 U12759 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10119) );
  INV_X1 U12760 ( .A(n13687), .ZN(n13694) );
  OAI221_X1 U12761 ( .B1(n20433), .B2(n20609), .C1(n20433), .C2(n20418), .A(
        n20686), .ZN(n20436) );
  NOR2_X1 U12762 ( .A1(n9652), .A2(n17776), .ZN(n10017) );
  INV_X1 U12763 ( .A(n20705), .ZN(n9828) );
  INV_X1 U12764 ( .A(n9828), .ZN(n9829) );
  INV_X1 U12765 ( .A(n20717), .ZN(n9830) );
  INV_X1 U12766 ( .A(n9830), .ZN(n9831) );
  AOI22_X2 U12767 ( .A1(DATAI_23_), .A2(n13686), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n13687), .ZN(n20733) );
  NOR2_X1 U12768 ( .A1(n14551), .A2(n13418), .ZN(n13687) );
  NOR3_X2 U12769 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18852), .A3(
        n18604), .ZN(n18620) );
  NOR3_X2 U12770 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18852), .A3(
        n18740), .ZN(n18711) );
  NOR3_X2 U12771 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18852), .A3(
        n18556), .ZN(n18531) );
  AOI22_X2 U12772 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n13687), .B1(DATAI_16_), 
        .B2(n13686), .ZN(n20691) );
  NOR2_X1 U12773 ( .A1(n14438), .A2(n14551), .ZN(n13686) );
  INV_X1 U12774 ( .A(n12693), .ZN(n10112) );
  OR2_X1 U12775 ( .A1(n12694), .A2(n12693), .ZN(n12697) );
  NOR2_X2 U12776 ( .A1(n13690), .A2(n9900), .ZN(n20680) );
  NAND3_X1 U12777 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20846), .A3(n13421), 
        .ZN(n13690) );
  NAND2_X1 U12778 ( .A1(n10029), .A2(n12022), .ZN(n10134) );
  NAND2_X1 U12779 ( .A1(n15319), .A2(n15318), .ZN(n12692) );
  NAND2_X1 U12780 ( .A1(n10219), .A2(n10217), .ZN(n12700) );
  NAND2_X1 U12781 ( .A1(n9837), .A2(n12018), .ZN(n12049) );
  NAND2_X1 U12782 ( .A1(n12017), .A2(n12016), .ZN(n9837) );
  AOI21_X1 U12783 ( .B1(n9840), .B2(n12332), .A(n12334), .ZN(n12333) );
  NAND2_X1 U12784 ( .A1(n15567), .A2(n9850), .ZN(n13037) );
  NAND2_X1 U12785 ( .A1(n15682), .A2(n20122), .ZN(n13517) );
  NAND2_X1 U12786 ( .A1(n16033), .A2(n9858), .ZN(n16034) );
  NAND2_X1 U12787 ( .A1(n9867), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9866) );
  NAND3_X1 U12788 ( .A1(n17888), .A2(n16038), .A3(n17836), .ZN(n9867) );
  NOR2_X1 U12789 ( .A1(n17841), .A2(n9866), .ZN(n17810) );
  NOR2_X4 U12790 ( .A1(n13939), .A2(n14035), .ZN(n15929) );
  INV_X2 U12791 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n19115) );
  NAND3_X1 U12792 ( .A1(n18100), .A2(n10008), .A3(n10007), .ZN(n9868) );
  NAND2_X1 U12793 ( .A1(n15929), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n9872) );
  AOI22_X1 U12794 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n15929), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15944) );
  AOI22_X1 U12795 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n15929), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17220) );
  AOI22_X1 U12796 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n15929), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17273) );
  AOI22_X1 U12797 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n15929), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17363) );
  AOI22_X1 U12798 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n15929), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17313) );
  AOI21_X1 U12799 ( .B1(n17448), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A(
        n9873), .ZN(n15930) );
  AND2_X1 U12800 ( .A1(n15929), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n9874) );
  AND2_X1 U12801 ( .A1(n15929), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n9875) );
  AND2_X1 U12802 ( .A1(n15929), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n9876) );
  AND2_X1 U12803 ( .A1(n15929), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n9877) );
  OAI211_X1 U12804 ( .C1(n18087), .C2(n9754), .A(n9887), .B(n9886), .ZN(n18078) );
  NAND2_X1 U12805 ( .A1(n18087), .A2(n9889), .ZN(n9886) );
  NAND2_X1 U12806 ( .A1(n9888), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9890) );
  NOR2_X1 U12807 ( .A1(n18087), .A2(n16009), .ZN(n16012) );
  INV_X1 U12808 ( .A(n9890), .ZN(n18077) );
  XNOR2_X2 U12809 ( .A(n15993), .B(n15988), .ZN(n15994) );
  NAND3_X1 U12810 ( .A1(n9663), .A2(n11192), .A3(n11191), .ZN(n9898) );
  NAND3_X1 U12811 ( .A1(n11258), .A2(n11192), .A3(n9742), .ZN(n9892) );
  OR2_X1 U12812 ( .A1(n9897), .A2(n9894), .ZN(n9893) );
  NAND3_X1 U12813 ( .A1(n9896), .A2(n9899), .A3(n9693), .ZN(n9895) );
  INV_X1 U12814 ( .A(n9897), .ZN(n9896) );
  NAND2_X1 U12815 ( .A1(n13347), .A2(n9898), .ZN(n13068) );
  NAND2_X1 U12816 ( .A1(n9899), .A2(n11190), .ZN(n13347) );
  OR2_X1 U12817 ( .A1(n13660), .A2(n20846), .ZN(n11269) );
  NAND2_X1 U12818 ( .A1(n9900), .A2(n11828), .ZN(n11847) );
  NAND2_X1 U12819 ( .A1(n9900), .A2(n9666), .ZN(n13654) );
  AOI21_X1 U12820 ( .B1(n11844), .B2(n9900), .A(n20846), .ZN(n11237) );
  AOI21_X1 U12821 ( .B1(n11154), .B2(n9666), .A(n9900), .ZN(n13069) );
  OAI21_X1 U12822 ( .B1(n11149), .B2(n11148), .A(n9900), .ZN(n11151) );
  AOI21_X1 U12823 ( .B1(n13079), .B2(n20850), .A(n9900), .ZN(n13214) );
  NAND3_X1 U12824 ( .A1(n9903), .A2(n13633), .A3(n11438), .ZN(n11452) );
  INV_X1 U12825 ( .A(n11438), .ZN(n9905) );
  OR2_X2 U12826 ( .A1(n14334), .A2(n9906), .ZN(n14280) );
  NAND2_X1 U12827 ( .A1(n12001), .A2(n12868), .ZN(n14199) );
  NAND3_X1 U12828 ( .A1(n15406), .A2(n12841), .A3(n9735), .ZN(n10133) );
  NAND3_X1 U12829 ( .A1(n15406), .A2(n12841), .A3(n9917), .ZN(n9916) );
  AND2_X2 U12830 ( .A1(n9953), .A2(n12492), .ZN(n10233) );
  NAND3_X1 U12831 ( .A1(n9921), .A2(n12840), .A3(n9920), .ZN(n15407) );
  NAND3_X1 U12832 ( .A1(n9731), .A2(n15668), .A3(n12837), .ZN(n9920) );
  AND2_X4 U12833 ( .A1(n13344), .A2(n13083), .ZN(n11690) );
  NAND3_X1 U12834 ( .A1(n11019), .A2(n11016), .A3(n11012), .ZN(n9941) );
  NAND2_X2 U12835 ( .A1(n9946), .A2(n9698), .ZN(n14595) );
  INV_X4 U12836 ( .A(n14628), .ZN(n16174) );
  NAND2_X2 U12837 ( .A1(n11895), .A2(n11894), .ZN(n14628) );
  NAND2_X2 U12838 ( .A1(n11380), .A2(n11379), .ZN(n11895) );
  NAND2_X1 U12839 ( .A1(n14628), .A2(n14640), .ZN(n13906) );
  XNOR2_X2 U12840 ( .A(n9952), .B(n12011), .ZN(n13269) );
  NAND2_X2 U12841 ( .A1(n10134), .A2(n10683), .ZN(n9952) );
  NAND2_X1 U12842 ( .A1(n12011), .A2(n9952), .ZN(n10694) );
  NAND4_X1 U12843 ( .A1(n12489), .A2(n12487), .A3(n12486), .A4(n12488), .ZN(
        n9953) );
  NAND4_X1 U12844 ( .A1(n12457), .A2(n12458), .A3(n12459), .A4(n12456), .ZN(
        n9954) );
  NAND4_X1 U12845 ( .A1(n10438), .A2(n10437), .A3(n10436), .A4(n9955), .ZN(
        n10439) );
  INV_X4 U12846 ( .A(n13524), .ZN(n12287) );
  NAND2_X1 U12847 ( .A1(n15278), .A2(n15279), .ZN(n15259) );
  INV_X1 U12848 ( .A(n15303), .ZN(n12701) );
  NAND3_X1 U12849 ( .A1(n16842), .A2(n16841), .A3(n9975), .ZN(P3_U2641) );
  NAND2_X1 U12850 ( .A1(n16865), .A2(n9815), .ZN(n9980) );
  AOI21_X1 U12851 ( .B1(n17146), .B2(n17786), .A(n9985), .ZN(n9981) );
  OR2_X1 U12852 ( .A1(n16865), .A2(n17146), .ZN(n9982) );
  NAND2_X1 U12853 ( .A1(n16927), .A2(n9797), .ZN(n9984) );
  NAND2_X1 U12854 ( .A1(n16885), .A2(n9991), .ZN(n9989) );
  INV_X2 U12855 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19108) );
  NAND3_X1 U12856 ( .A1(n15961), .A2(n10002), .A3(n10001), .ZN(n10000) );
  INV_X1 U12857 ( .A(n18085), .ZN(n10011) );
  OR2_X2 U12858 ( .A1(n10019), .A2(n12448), .ZN(n12532) );
  OR2_X2 U12859 ( .A1(n12450), .A2(n10019), .ZN(n19448) );
  OR2_X2 U12860 ( .A1(n13269), .A2(n12980), .ZN(n10019) );
  NAND4_X1 U12861 ( .A1(n10024), .A2(n10361), .A3(n10362), .A4(n10363), .ZN(
        n10023) );
  NAND2_X1 U12862 ( .A1(n12829), .A2(n12494), .ZN(n13702) );
  NAND3_X1 U12863 ( .A1(n12829), .A2(n10026), .A3(n12494), .ZN(n10025) );
  NAND3_X1 U12864 ( .A1(n10675), .A2(n10674), .A3(n12021), .ZN(n10029) );
  NAND3_X1 U12865 ( .A1(n10233), .A2(n10234), .A3(n12827), .ZN(n12562) );
  NAND2_X1 U12866 ( .A1(n10031), .A2(n12838), .ZN(n12842) );
  NAND3_X1 U12867 ( .A1(n10034), .A2(n10033), .A3(n10032), .ZN(n10041) );
  NAND2_X1 U12868 ( .A1(n9722), .A2(n10035), .ZN(n10032) );
  NAND2_X1 U12869 ( .A1(n9722), .A2(n15342), .ZN(n15344) );
  NAND3_X1 U12870 ( .A1(n10034), .A2(n10036), .A3(n10032), .ZN(n15535) );
  NAND2_X1 U12871 ( .A1(n10041), .A2(n15534), .ZN(P2_U3025) );
  INV_X1 U12872 ( .A(n16437), .ZN(n10049) );
  NAND2_X1 U12873 ( .A1(n16437), .A2(n10045), .ZN(n10043) );
  NAND2_X1 U12874 ( .A1(n16437), .A2(n16434), .ZN(n10060) );
  AND2_X1 U12875 ( .A1(n15331), .A2(n16434), .ZN(n10058) );
  NAND2_X1 U12876 ( .A1(n16465), .A2(n10066), .ZN(n10061) );
  NAND2_X1 U12877 ( .A1(n10061), .A2(n10063), .ZN(n15329) );
  INV_X1 U12878 ( .A(n15618), .ZN(n10069) );
  XNOR2_X1 U12879 ( .A(n10073), .B(n13461), .ZN(n13611) );
  NAND2_X1 U12880 ( .A1(n10123), .A2(n11857), .ZN(n10073) );
  INV_X1 U12881 ( .A(n16197), .ZN(n10078) );
  NAND2_X1 U12882 ( .A1(n16195), .A2(n16197), .ZN(n10081) );
  NAND2_X1 U12883 ( .A1(n10076), .A2(n10074), .ZN(n13888) );
  NAND2_X1 U12884 ( .A1(n11900), .A2(n10079), .ZN(n10075) );
  NOR2_X1 U12885 ( .A1(n10080), .A2(n10078), .ZN(n10077) );
  INV_X1 U12886 ( .A(n16196), .ZN(n10079) );
  NAND2_X1 U12887 ( .A1(n11347), .A2(n20846), .ZN(n10083) );
  XNOR2_X2 U12888 ( .A(n11210), .B(n11209), .ZN(n11347) );
  NAND2_X1 U12889 ( .A1(n10086), .A2(n14557), .ZN(n14525) );
  NAND2_X2 U12890 ( .A1(n14626), .A2(n11904), .ZN(n16186) );
  NAND2_X1 U12891 ( .A1(n10090), .A2(n10089), .ZN(n11913) );
  NAND3_X1 U12892 ( .A1(n14185), .A2(n14184), .A3(n10092), .ZN(P1_U2809) );
  OR2_X1 U12893 ( .A1(n14186), .A2(n20178), .ZN(n10092) );
  NAND3_X1 U12894 ( .A1(n13724), .A2(n9711), .A3(n13877), .ZN(n13900) );
  INV_X1 U12895 ( .A(n15255), .ZN(n10109) );
  NAND2_X1 U12896 ( .A1(n15256), .A2(n15258), .ZN(n10111) );
  NOR3_X1 U12897 ( .A1(n12694), .A2(P2_EBX_REG_24__SCAN_IN), .A3(n12693), .ZN(
        n12704) );
  NAND3_X1 U12898 ( .A1(n10113), .A2(n9817), .A3(n10112), .ZN(n12712) );
  NAND2_X1 U12899 ( .A1(n12621), .A2(n9795), .ZN(n12645) );
  NAND2_X1 U12900 ( .A1(n12656), .A2(n9798), .ZN(n12688) );
  INV_X1 U12901 ( .A(n10121), .ZN(n12613) );
  NAND2_X1 U12902 ( .A1(n13403), .A2(n13402), .ZN(n10123) );
  NAND2_X1 U12903 ( .A1(n11831), .A2(n11830), .ZN(n13182) );
  NAND2_X1 U12904 ( .A1(n13209), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11841) );
  NAND2_X1 U12905 ( .A1(n10125), .A2(n11838), .ZN(n10124) );
  NAND2_X1 U12906 ( .A1(n13182), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10125) );
  NAND2_X1 U12907 ( .A1(n10127), .A2(n13182), .ZN(n10126) );
  NOR2_X1 U12908 ( .A1(n11838), .A2(n10128), .ZN(n10127) );
  NAND2_X1 U12909 ( .A1(n13182), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11837) );
  INV_X1 U12910 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n10128) );
  INV_X1 U12911 ( .A(n11331), .ZN(n10143) );
  INV_X1 U12912 ( .A(n11332), .ZN(n10144) );
  NAND2_X1 U12913 ( .A1(n9757), .A2(n10147), .ZN(n10149) );
  NOR2_X2 U12914 ( .A1(n16186), .A2(n10152), .ZN(n10147) );
  OAI211_X1 U12915 ( .C1(n14809), .C2(n14808), .A(n10153), .B(n19315), .ZN(
        n14820) );
  OAI21_X1 U12916 ( .B1(n10153), .B2(n19339), .A(n10280), .ZN(n11004) );
  XNOR2_X1 U12917 ( .A(n15981), .B(n15980), .ZN(n18067) );
  NOR2_X2 U12918 ( .A1(n13939), .A2(n10155), .ZN(n13971) );
  NAND2_X1 U12919 ( .A1(n10327), .A2(n9821), .ZN(n10290) );
  INV_X1 U12920 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10158) );
  NAND2_X1 U12921 ( .A1(n10292), .A2(n9816), .ZN(n10326) );
  NAND2_X1 U12922 ( .A1(n14096), .A2(n19974), .ZN(n10173) );
  NAND2_X1 U12923 ( .A1(n10173), .A2(n10172), .ZN(n19244) );
  NAND2_X1 U12924 ( .A1(n14855), .A2(n9796), .ZN(n15068) );
  NAND2_X1 U12925 ( .A1(n14991), .A2(n10178), .ZN(n10786) );
  NAND2_X1 U12926 ( .A1(n14991), .A2(n14982), .ZN(n14984) );
  NAND2_X1 U12927 ( .A1(n13444), .A2(n9756), .ZN(n14871) );
  NAND2_X1 U12928 ( .A1(n13035), .A2(n10189), .ZN(n13503) );
  NAND2_X1 U12929 ( .A1(n14858), .A2(n15604), .ZN(n15240) );
  INV_X1 U12930 ( .A(n15158), .ZN(n10207) );
  NAND2_X1 U12931 ( .A1(n10207), .A2(n10208), .ZN(n15131) );
  INV_X1 U12932 ( .A(n15131), .ZN(n10993) );
  NAND2_X1 U12933 ( .A1(n15247), .A2(n15246), .ZN(n10215) );
  NAND2_X1 U12934 ( .A1(n15247), .A2(n10213), .ZN(n10212) );
  INV_X1 U12935 ( .A(n15246), .ZN(n10214) );
  NAND2_X1 U12936 ( .A1(n10215), .A2(n15245), .ZN(n12731) );
  INV_X1 U12937 ( .A(n10216), .ZN(n10217) );
  OAI21_X1 U12938 ( .B1(n15311), .B2(n9728), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10216) );
  NAND2_X1 U12939 ( .A1(n12692), .A2(n10220), .ZN(n10219) );
  CLKBUF_X1 U12940 ( .A(n10226), .Z(n10223) );
  NAND2_X1 U12941 ( .A1(n12599), .A2(n12598), .ZN(n15383) );
  INV_X2 U12942 ( .A(n10605), .ZN(n10631) );
  NAND2_X2 U12943 ( .A1(n10229), .A2(n10227), .ZN(n10605) );
  NAND2_X1 U12944 ( .A1(n10228), .A2(n10489), .ZN(n10227) );
  NAND4_X1 U12945 ( .A1(n10360), .A2(n10357), .A3(n10359), .A4(n10358), .ZN(
        n10228) );
  NAND2_X1 U12946 ( .A1(n10230), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10229) );
  NAND4_X1 U12947 ( .A1(n10355), .A2(n10354), .A3(n10353), .A4(n10356), .ZN(
        n10230) );
  AND3_X2 U12948 ( .A1(n12703), .A2(n12702), .A3(n10232), .ZN(n15278) );
  AND2_X2 U12949 ( .A1(n12340), .A2(n10595), .ZN(n10604) );
  NAND2_X1 U12950 ( .A1(n10617), .A2(n12733), .ZN(n10595) );
  NOR2_X2 U12951 ( .A1(n10442), .A2(n12335), .ZN(n10617) );
  AND2_X1 U12952 ( .A1(n19459), .A2(n20115), .ZN(n10235) );
  NAND3_X1 U12953 ( .A1(n10241), .A2(n14973), .A3(n14981), .ZN(n14979) );
  INV_X1 U12954 ( .A(n10245), .ZN(n15015) );
  NAND2_X1 U12955 ( .A1(n10246), .A2(n9715), .ZN(n15108) );
  NAND4_X1 U12956 ( .A1(n10251), .A2(n13146), .A3(n10252), .A4(n13147), .ZN(
        n13397) );
  NAND3_X1 U12957 ( .A1(n13633), .A2(n13747), .A3(n10277), .ZN(n13762) );
  NAND2_X1 U12958 ( .A1(n13928), .A2(n10256), .ZN(n14347) );
  NAND2_X1 U12959 ( .A1(n13928), .A2(n13930), .ZN(n13929) );
  INV_X1 U12960 ( .A(n12834), .ZN(n12837) );
  OR2_X1 U12961 ( .A1(n13266), .A2(n13267), .ZN(n13268) );
  AOI22_X1 U12962 ( .A1(n10450), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9671), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10452) );
  NAND2_X1 U12963 ( .A1(n10636), .A2(n10635), .ZN(n12780) );
  OR2_X1 U12964 ( .A1(n14103), .A2(n16587), .ZN(n14112) );
  NAND2_X1 U12965 ( .A1(n15259), .A2(n15257), .ZN(n15256) );
  NAND2_X1 U12966 ( .A1(n12701), .A2(n10218), .ZN(n12702) );
  NAND2_X2 U12967 ( .A1(n10351), .A2(n13522), .ZN(n12132) );
  OR2_X1 U12968 ( .A1(n13160), .A2(n13159), .ZN(n13161) );
  NAND2_X1 U12969 ( .A1(n10652), .A2(n10651), .ZN(n10671) );
  INV_X1 U12970 ( .A(n11377), .ZN(n11380) );
  NAND2_X1 U12971 ( .A1(n11305), .A2(n11377), .ZN(n11871) );
  NAND2_X1 U12972 ( .A1(n13893), .A2(n11452), .ZN(n13928) );
  AND2_X1 U12973 ( .A1(n20216), .A2(n11306), .ZN(n20212) );
  INV_X1 U12974 ( .A(n20135), .ZN(n11980) );
  NOR2_X1 U12975 ( .A1(n13101), .A2(n13100), .ZN(n16067) );
  NAND2_X2 U12976 ( .A1(n14498), .A2(n13157), .ZN(n14505) );
  AND2_X1 U12977 ( .A1(n12416), .A2(n12415), .ZN(n10267) );
  OR2_X1 U12978 ( .A1(n12853), .A2(n12852), .ZN(n16587) );
  NOR2_X1 U12979 ( .A1(n20162), .A2(n20161), .ZN(n10268) );
  NOR2_X1 U12980 ( .A1(n14075), .A2(n20161), .ZN(n10269) );
  OR2_X1 U12981 ( .A1(n15007), .A2(n12186), .ZN(n10270) );
  OR2_X1 U12982 ( .A1(n14804), .A2(n20846), .ZN(n10271) );
  INV_X1 U12983 ( .A(n20678), .ZN(n20596) );
  NAND2_X1 U12984 ( .A1(n20753), .A2(n20609), .ZN(n20678) );
  AND4_X1 U12985 ( .A1(n15917), .A2(n15916), .A3(n15915), .A4(n15914), .ZN(
        n10273) );
  AND2_X1 U12986 ( .A1(n10371), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n10274) );
  INV_X1 U12987 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11923) );
  NAND2_X1 U12988 ( .A1(n12864), .A2(n15751), .ZN(n19429) );
  INV_X1 U12989 ( .A(n19429), .ZN(n16496) );
  AND2_X1 U12990 ( .A1(n12834), .A2(n15422), .ZN(n10275) );
  AND2_X1 U12991 ( .A1(n14807), .A2(n16592), .ZN(n10276) );
  NAND3_X1 U12992 ( .A1(n11403), .A2(n11402), .A3(n11401), .ZN(n10277) );
  OR3_X1 U12993 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n17859), .ZN(n10278) );
  AND4_X1 U12994 ( .A1(n10376), .A2(n10375), .A3(n10374), .A4(n10373), .ZN(
        n10279) );
  INV_X1 U12995 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20155) );
  NOR2_X1 U12996 ( .A1(n10600), .A2(n10599), .ZN(n10280) );
  AND2_X1 U12997 ( .A1(n19438), .A2(n20080), .ZN(n19435) );
  INV_X1 U12998 ( .A(n19435), .ZN(n16433) );
  AND4_X1 U12999 ( .A1(n10493), .A2(n10492), .A3(n10491), .A4(n10490), .ZN(
        n10281) );
  INV_X2 U13000 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20753) );
  AND2_X1 U13001 ( .A1(n13654), .A2(n11172), .ZN(n10282) );
  AND3_X1 U13002 ( .A1(n10449), .A2(n10448), .A3(n10489), .ZN(n10283) );
  INV_X1 U13003 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16476) );
  INV_X1 U13004 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16428) );
  INV_X1 U13005 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11919) );
  OAI21_X1 U13006 ( .B1(n15451), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n9724), .ZN(n15438) );
  OR3_X1 U13007 ( .A1(n17022), .A2(n17014), .A3(n19034), .ZN(n10284) );
  NAND2_X1 U13008 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18991), .ZN(n17137) );
  NOR2_X1 U13009 ( .A1(n17977), .A2(n18101), .ZN(n17920) );
  INV_X1 U13010 ( .A(n17920), .ZN(n17881) );
  OR2_X1 U13011 ( .A1(n13344), .A2(n13349), .ZN(n10285) );
  AND3_X1 U13012 ( .A1(n11036), .A2(n11035), .A3(n11034), .ZN(n10286) );
  OR2_X1 U13013 ( .A1(n16668), .A2(n17628), .ZN(n10287) );
  OR2_X1 U13014 ( .A1(n16103), .A2(n16651), .ZN(n10288) );
  AND2_X1 U13015 ( .A1(n17496), .A2(n17489), .ZN(n17500) );
  INV_X2 U13016 ( .A(n17500), .ZN(n17494) );
  NAND2_X1 U13017 ( .A1(n12429), .A2(n13269), .ZN(n12439) );
  OR2_X1 U13018 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20532), .ZN(
        n11930) );
  NOR2_X1 U13019 ( .A1(n11963), .A2(n12381), .ZN(n11965) );
  INV_X1 U13020 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10331) );
  AOI22_X1 U13021 ( .A1(n12308), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10488), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10360) );
  XNOR2_X1 U13022 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11938) );
  INV_X1 U13023 ( .A(n11843), .ZN(n11259) );
  INV_X1 U13024 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12470) );
  INV_X1 U13025 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12438) );
  NOR2_X1 U13026 ( .A1(n12747), .A2(n12322), .ZN(n10329) );
  NOR3_X1 U13027 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20294), .A3(
        n11972), .ZN(n12382) );
  NAND2_X1 U13028 ( .A1(n11934), .A2(n11933), .ZN(n11972) );
  AOI22_X1 U13029 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11112), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11011) );
  AND3_X1 U13030 ( .A1(n11254), .A2(n11253), .A3(n11252), .ZN(n11261) );
  INV_X1 U13031 ( .A(n10344), .ZN(n10346) );
  INV_X1 U13032 ( .A(n12187), .ZN(n12188) );
  INV_X1 U13033 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10352) );
  OAI22_X1 U13034 ( .A1(n12426), .A2(n19830), .B1(n19875), .B2(n12425), .ZN(
        n12427) );
  INV_X1 U13035 ( .A(n14246), .ZN(n11707) );
  OAI21_X1 U13036 ( .B1(n11544), .B2(n11386), .A(n11385), .ZN(n11387) );
  AND2_X1 U13037 ( .A1(n11210), .A2(n11208), .ZN(n11255) );
  AND4_X1 U13038 ( .A1(n11046), .A2(n11045), .A3(n11044), .A4(n11043), .ZN(
        n11047) );
  INV_X1 U13039 ( .A(n11234), .ZN(n11235) );
  NAND2_X1 U13040 ( .A1(n10346), .A2(n10345), .ZN(n10348) );
  INV_X1 U13041 ( .A(n13597), .ZN(n12052) );
  INV_X1 U13042 ( .A(n12234), .ZN(n12235) );
  AOI22_X1 U13043 ( .A1(n9643), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10488), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10444) );
  OAI21_X1 U13044 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n19108), .A(
        n14036), .ZN(n14041) );
  NAND2_X1 U13045 ( .A1(n11306), .A2(n11134), .ZN(n11143) );
  INV_X1 U13046 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13332) );
  AND2_X1 U13047 ( .A1(n11724), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11725) );
  NAND2_X1 U13048 ( .A1(n13433), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11544) );
  INV_X1 U13049 ( .A(n14154), .ZN(n14151) );
  AND2_X1 U13050 ( .A1(n10981), .A2(n10980), .ZN(n15155) );
  AND2_X1 U13051 ( .A1(n15101), .A2(n15093), .ZN(n12054) );
  OR2_X1 U13052 ( .A1(n12230), .A2(n12232), .ZN(n12257) );
  INV_X1 U13053 ( .A(n12310), .ZN(n12302) );
  INV_X1 U13054 ( .A(n12215), .ZN(n12212) );
  AND2_X1 U13055 ( .A1(n10765), .A2(n10764), .ZN(n14998) );
  INV_X1 U13056 ( .A(n12847), .ZN(n12848) );
  NOR2_X1 U13057 ( .A1(n18944), .A2(n13941), .ZN(n15894) );
  AND2_X1 U13058 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15978), .ZN(
        n15979) );
  NOR2_X1 U13059 ( .A1(n18512), .A2(n18493), .ZN(n15984) );
  NOR2_X1 U13060 ( .A1(n9665), .A2(n13660), .ZN(n11176) );
  OR2_X1 U13061 ( .A1(n11821), .A2(n14511), .ZN(n11984) );
  NAND2_X1 U13062 ( .A1(n11725), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11765) );
  AND2_X1 U13063 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n11632), .ZN(
        n11633) );
  NOR2_X1 U13064 ( .A1(n11597), .A2(n14328), .ZN(n11598) );
  INV_X1 U13065 ( .A(n9799), .ZN(n13644) );
  NOR2_X1 U13066 ( .A1(n20643), .A2(n13780), .ZN(n13691) );
  OR2_X2 U13067 ( .A1(n11084), .A2(n11083), .ZN(n11828) );
  NAND2_X1 U13068 ( .A1(n20467), .A2(n20846), .ZN(n11282) );
  NAND2_X1 U13069 ( .A1(n10435), .A2(n10489), .ZN(n10441) );
  AND2_X1 U13070 ( .A1(n12210), .A2(n12209), .ZN(n12213) );
  AND2_X1 U13071 ( .A1(n10972), .A2(n10971), .ZN(n14838) );
  AND2_X1 U13072 ( .A1(n10372), .A2(n10489), .ZN(n12152) );
  OAI21_X1 U13073 ( .B1(n15423), .B2(n15419), .A(n12834), .ZN(n12841) );
  NAND2_X1 U13075 ( .A1(n10606), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12997) );
  AND2_X1 U13076 ( .A1(n19974), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12039) );
  NOR2_X1 U13077 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13510) );
  INV_X1 U13078 ( .A(n17787), .ZN(n16822) );
  INV_X1 U13079 ( .A(n15987), .ZN(n18927) );
  INV_X1 U13080 ( .A(n18497), .ZN(n15877) );
  NOR2_X1 U13081 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17952), .ZN(
        n17914) );
  NOR2_X1 U13082 ( .A1(n18120), .A2(n15968), .ZN(n15971) );
  INV_X1 U13083 ( .A(n18949), .ZN(n18931) );
  INV_X1 U13084 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16141) );
  INV_X1 U13085 ( .A(n20175), .ZN(n20192) );
  INV_X1 U13086 ( .A(n11495), .ZN(n11529) );
  NAND2_X1 U13087 ( .A1(n11498), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11515) );
  OR2_X1 U13088 ( .A1(n11986), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14779) );
  INV_X1 U13089 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14792) );
  OR2_X1 U13090 ( .A1(n11842), .A2(n9664), .ZN(n20442) );
  AND2_X1 U13091 ( .A1(n13473), .A2(n13472), .ZN(n13624) );
  OR2_X1 U13092 ( .A1(n20442), .A2(n13389), .ZN(n13477) );
  OR2_X1 U13093 ( .A1(n13387), .A2(n13388), .ZN(n20569) );
  NOR2_X1 U13094 ( .A1(n20530), .A2(n20298), .ZN(n20686) );
  INV_X1 U13095 ( .A(n13686), .ZN(n13693) );
  INV_X1 U13096 ( .A(n19326), .ZN(n19303) );
  AND2_X1 U13097 ( .A1(n10349), .A2(n12751), .ZN(n13562) );
  OR2_X1 U13098 ( .A1(n10917), .A2(n10916), .ZN(n15093) );
  AND3_X1 U13099 ( .A1(n10890), .A2(n10889), .A3(n10888), .ZN(n13273) );
  NAND2_X1 U13100 ( .A1(n19357), .A2(n12413), .ZN(n19358) );
  INV_X1 U13101 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15273) );
  AND2_X1 U13102 ( .A1(n10932), .A2(n10931), .ZN(n14860) );
  OR2_X1 U13103 ( .A1(n12799), .A2(n12798), .ZN(n16556) );
  XNOR2_X1 U13104 ( .A(n15684), .B(n12042), .ZN(n13045) );
  AND2_X1 U13105 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19779) );
  INV_X1 U13106 ( .A(n12543), .ZN(n19641) );
  NOR2_X1 U13107 ( .A1(n19440), .A2(n15724), .ZN(n20064) );
  NAND2_X1 U13108 ( .A1(n19440), .A2(n15724), .ZN(n19835) );
  INV_X1 U13109 ( .A(n19480), .ZN(n19483) );
  INV_X1 U13110 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19974) );
  OAI21_X1 U13111 ( .B1(n14045), .B2(n14051), .A(n14052), .ZN(n18917) );
  INV_X1 U13112 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16845) );
  NOR2_X1 U13113 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17026), .ZN(n17006) );
  INV_X1 U13114 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17102) );
  NOR2_X1 U13115 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17124), .ZN(n17106) );
  NAND2_X1 U13116 ( .A1(n18929), .A2(n18927), .ZN(n18914) );
  NOR2_X1 U13117 ( .A1(n14030), .A2(n18934), .ZN(n15831) );
  NOR2_X1 U13118 ( .A1(n17717), .A2(n17548), .ZN(n17547) );
  NOR2_X1 U13119 ( .A1(n17703), .A2(n17590), .ZN(n17585) );
  INV_X1 U13120 ( .A(n17837), .ZN(n17986) );
  AOI21_X1 U13121 ( .B1(n18143), .B2(n18468), .A(n19109), .ZN(n18479) );
  OR2_X1 U13122 ( .A1(n18172), .A2(n18277), .ZN(n17819) );
  NOR2_X1 U13123 ( .A1(n18173), .A2(n18242), .ZN(n18204) );
  INV_X1 U13124 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17993) );
  INV_X1 U13125 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18959) );
  INV_X1 U13126 ( .A(n20185), .ZN(n20161) );
  AND2_X1 U13127 ( .A1(n14140), .A2(n13665), .ZN(n20183) );
  INV_X1 U13128 ( .A(n20216), .ZN(n14429) );
  OR2_X1 U13129 ( .A1(n13133), .A2(n14163), .ZN(n13134) );
  INV_X1 U13130 ( .A(n14498), .ZN(n14502) );
  INV_X1 U13131 ( .A(n13164), .ZN(n20260) );
  NAND2_X1 U13132 ( .A1(n12007), .A2(n12006), .ZN(n12008) );
  NAND2_X1 U13133 ( .A1(n11435), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11467) );
  AND2_X1 U13134 ( .A1(n11434), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11435) );
  AND2_X1 U13135 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n11323), .ZN(
        n11384) );
  INV_X1 U13136 ( .A(n14715), .ZN(n14765) );
  NAND2_X1 U13137 ( .A1(n16284), .A2(n14715), .ZN(n16287) );
  AND2_X1 U13138 ( .A1(n13223), .A2(n9937), .ZN(n13238) );
  NOR2_X1 U13139 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n16336) );
  OAI22_X1 U13140 ( .A1(n20304), .A2(n20303), .B1(n20469), .B2(n20414), .ZN(
        n20320) );
  OAI22_X1 U13141 ( .A1(n20358), .A2(n20357), .B1(n20356), .B2(n20469), .ZN(
        n20376) );
  INV_X1 U13142 ( .A(n20380), .ZN(n20406) );
  NOR2_X2 U13143 ( .A1(n20386), .A2(n20385), .ZN(n20435) );
  NOR2_X2 U13144 ( .A1(n20442), .A2(n20642), .ZN(n20461) );
  NOR2_X1 U13145 ( .A1(n13477), .A2(n13420), .ZN(n13790) );
  NOR2_X1 U13146 ( .A1(n13477), .A2(n13781), .ZN(n20490) );
  INV_X1 U13147 ( .A(n20411), .ZN(n20466) );
  NOR2_X2 U13148 ( .A1(n20569), .A2(n20642), .ZN(n20554) );
  NOR2_X2 U13149 ( .A1(n20569), .A2(n20525), .ZN(n20591) );
  INV_X1 U13150 ( .A(n20610), .ZN(n20636) );
  NOR2_X2 U13151 ( .A1(n20595), .A2(n13420), .ZN(n20669) );
  NOR2_X1 U13152 ( .A1(n20643), .A2(n20673), .ZN(n20742) );
  NAND2_X1 U13153 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20850) );
  INV_X1 U13154 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20129) );
  INV_X1 U13155 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20755) );
  NAND2_X1 U13156 ( .A1(n16352), .A2(n16353), .ZN(n16351) );
  NAND2_X1 U13157 ( .A1(n16388), .A2(n16389), .ZN(n16387) );
  INV_X1 U13158 ( .A(n19321), .ZN(n19314) );
  INV_X1 U13159 ( .A(n15056), .ZN(n15083) );
  OR2_X1 U13160 ( .A1(n10930), .A2(n10929), .ZN(n15088) );
  INV_X1 U13161 ( .A(n12317), .ZN(n12318) );
  INV_X1 U13162 ( .A(n16605), .ZN(n13010) );
  INV_X1 U13163 ( .A(n12951), .ZN(n12941) );
  AND2_X1 U13164 ( .A1(n15098), .A2(n15097), .ZN(n19274) );
  AND2_X1 U13165 ( .A1(n13314), .A2(n13313), .ZN(n19434) );
  INV_X1 U13166 ( .A(n19438), .ZN(n16477) );
  OR2_X1 U13167 ( .A1(n15570), .A2(n9847), .ZN(n16526) );
  INV_X1 U13168 ( .A(n16587), .ZN(n16566) );
  NOR2_X1 U13169 ( .A1(n15684), .A2(n12999), .ZN(n20093) );
  OAI21_X1 U13170 ( .B1(n19452), .B2(n19451), .A(n19450), .ZN(n19490) );
  NOR2_X1 U13171 ( .A1(n19553), .A2(n19636), .ZN(n19578) );
  INV_X1 U13172 ( .A(n19599), .ZN(n19614) );
  NOR2_X2 U13173 ( .A1(n19636), .A2(n19835), .ZN(n19630) );
  NOR2_X2 U13174 ( .A1(n19667), .A2(n19835), .ZN(n19662) );
  NAND2_X1 U13175 ( .A1(n19727), .A2(n20093), .ZN(n19667) );
  INV_X1 U13176 ( .A(n19919), .ZN(n19639) );
  INV_X1 U13177 ( .A(n19758), .ZN(n19774) );
  AND2_X1 U13178 ( .A1(n19785), .A2(n19783), .ZN(n19805) );
  NOR2_X1 U13179 ( .A1(n19865), .A2(n19835), .ZN(n19823) );
  INV_X1 U13180 ( .A(n19942), .ZN(n19889) );
  NOR2_X1 U13181 ( .A1(n19591), .A2(n10677), .ZN(n13583) );
  INV_X1 U13182 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19997) );
  NAND2_X1 U13183 ( .A1(n19136), .A2(n18267), .ZN(n18921) );
  NOR2_X1 U13184 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16890), .ZN(n16874) );
  NOR2_X1 U13185 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16913), .ZN(n16898) );
  NOR2_X1 U13186 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16981), .ZN(n16959) );
  NOR2_X1 U13187 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16994), .ZN(n16984) );
  NOR2_X1 U13188 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17051), .ZN(n17032) );
  NOR2_X1 U13189 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17077), .ZN(n17061) );
  NAND4_X1 U13190 ( .A1(n18447), .A2(n19147), .A3(n17137), .A4(n18979), .ZN(
        n17189) );
  NOR2_X2 U13191 ( .A1(n16804), .A2(n16808), .ZN(n17168) );
  NOR2_X1 U13192 ( .A1(n17199), .A2(n17279), .ZN(n17261) );
  INV_X1 U13193 ( .A(n17478), .ZN(n17468) );
  NOR2_X1 U13194 ( .A1(n17499), .A2(n17473), .ZN(n17478) );
  INV_X1 U13195 ( .A(n17496), .ZN(n17499) );
  NOR2_X1 U13196 ( .A1(n17721), .A2(n17541), .ZN(n17536) );
  NOR2_X1 U13197 ( .A1(n17552), .A2(n17572), .ZN(n17562) );
  INV_X1 U13198 ( .A(n17553), .ZN(n17583) );
  INV_X1 U13199 ( .A(n17603), .ZN(n17646) );
  AND2_X1 U13200 ( .A1(n18952), .A2(n16127), .ZN(n17655) );
  NAND3_X1 U13201 ( .A1(n13983), .A2(n13982), .A3(n13981), .ZN(n17661) );
  INV_X1 U13202 ( .A(n18052), .ZN(n18041) );
  NAND2_X1 U13203 ( .A1(n18144), .A2(n18045), .ZN(n18071) );
  INV_X1 U13204 ( .A(n18050), .ZN(n17952) );
  NOR2_X1 U13205 ( .A1(n18204), .A2(n18459), .ZN(n18214) );
  INV_X1 U13206 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17926) );
  INV_X1 U13207 ( .A(n18388), .ZN(n18362) );
  INV_X1 U13208 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18380) );
  INV_X1 U13209 ( .A(n18460), .ZN(n18454) );
  NOR2_X1 U13210 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19086), .ZN(
        n19109) );
  INV_X1 U13211 ( .A(n18617), .ZN(n18621) );
  INV_X1 U13212 ( .A(n18646), .ZN(n18635) );
  INV_X1 U13213 ( .A(n18665), .ZN(n18667) );
  INV_X1 U13214 ( .A(n18734), .ZN(n18736) );
  INV_X1 U13215 ( .A(n18755), .ZN(n18759) );
  INV_X1 U13216 ( .A(n18803), .ZN(n18815) );
  INV_X1 U13217 ( .A(n18825), .ZN(n18847) );
  INV_X1 U13218 ( .A(n18790), .ZN(n18906) );
  NOR2_X1 U13219 ( .A1(n16802), .A2(n18978), .ZN(n19131) );
  INV_X1 U13220 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20841) );
  NAND2_X1 U13221 ( .A1(n13734), .A2(n13648), .ZN(n20178) );
  INV_X1 U13222 ( .A(n14613), .ZN(n14487) );
  AND2_X1 U13223 ( .A1(n13169), .A2(n13168), .ZN(n13623) );
  OR2_X1 U13224 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16341), .ZN(n20218) );
  INV_X1 U13225 ( .A(n20220), .ZN(n20246) );
  NOR2_X1 U13226 ( .A1(n13109), .A2(n13020), .ZN(n13163) );
  NAND2_X1 U13227 ( .A1(n16209), .A2(n13185), .ZN(n16202) );
  NAND2_X2 U13228 ( .A1(n12971), .A2(n9692), .ZN(n20135) );
  NAND2_X1 U13229 ( .A1(n13238), .A2(n13228), .ZN(n16260) );
  INV_X1 U13230 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20294) );
  OR2_X1 U13231 ( .A1(n16334), .A2(n13104), .ZN(n16340) );
  OR2_X1 U13232 ( .A1(n20386), .A2(n20411), .ZN(n20324) );
  OR2_X1 U13233 ( .A1(n20386), .A2(n20642), .ZN(n20373) );
  AOI22_X1 U13234 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20384), .B1(n20389), 
        .B2(n20383), .ZN(n20410) );
  NAND2_X1 U13235 ( .A1(n20412), .A2(n20466), .ZN(n20465) );
  INV_X1 U13236 ( .A(n13785), .ZN(n13826) );
  INV_X1 U13237 ( .A(n20490), .ZN(n13697) );
  NAND2_X1 U13238 ( .A1(n20560), .A2(n20466), .ZN(n20522) );
  AOI22_X1 U13239 ( .A1(n20533), .A2(n20537), .B1(n20531), .B2(n20530), .ZN(
        n20558) );
  NAND2_X1 U13240 ( .A1(n20560), .A2(n20559), .ZN(n20610) );
  AOI22_X1 U13241 ( .A1(n20607), .A2(n20604), .B1(n20601), .B2(n20600), .ZN(
        n20641) );
  OR2_X1 U13242 ( .A1(n20648), .A2(n20642), .ZN(n20681) );
  OR2_X1 U13243 ( .A1(n20648), .A2(n20525), .ZN(n20749) );
  INV_X1 U13244 ( .A(n20746), .ZN(n13715) );
  NAND2_X1 U13245 ( .A1(n16345), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20751) );
  INV_X1 U13246 ( .A(n20831), .ZN(n20827) );
  INV_X1 U13247 ( .A(n20791), .ZN(n20816) );
  INV_X1 U13248 ( .A(n20817), .ZN(n20854) );
  NAND2_X1 U13249 ( .A1(n12856), .A2(n12855), .ZN(n12913) );
  INV_X1 U13250 ( .A(n19324), .ZN(n19304) );
  NAND2_X1 U13251 ( .A1(n13265), .A2(n13268), .ZN(n19727) );
  INV_X1 U13252 ( .A(n19440), .ZN(n20075) );
  NAND2_X1 U13253 ( .A1(n19357), .A2(n12352), .ZN(n15230) );
  NOR2_X1 U13254 ( .A1(n19385), .A2(n19383), .ZN(n19355) );
  AND2_X1 U13255 ( .A1(n15134), .A2(n13052), .ZN(n19389) );
  NAND2_X1 U13256 ( .A1(n19391), .A2(n13014), .ZN(n13207) );
  INV_X1 U13257 ( .A(n19391), .ZN(n19423) );
  INV_X1 U13258 ( .A(n12949), .ZN(n13011) );
  INV_X1 U13259 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n19249) );
  INV_X1 U13260 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16458) );
  INV_X1 U13261 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16500) );
  AOI21_X1 U13262 ( .B1(n15268), .B2(n16566), .A(n15447), .ZN(n15448) );
  OR2_X1 U13263 ( .A1(n12853), .A2(n12766), .ZN(n16570) );
  INV_X1 U13264 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16121) );
  OR2_X1 U13265 ( .A1(n19728), .A2(n19636), .ZN(n19522) );
  INV_X1 U13266 ( .A(n19578), .ZN(n19576) );
  INV_X1 U13267 ( .A(n19595), .ZN(n19617) );
  AOI21_X1 U13268 ( .B1(n15705), .B2(n19583), .A(n15704), .ZN(n19635) );
  AOI211_X2 U13269 ( .C1(n19640), .C2(n19643), .A(n19639), .B(n19638), .ZN(
        n19666) );
  OR2_X1 U13270 ( .A1(n19864), .A2(n19667), .ZN(n19725) );
  NAND2_X1 U13271 ( .A1(n19695), .A2(n19694), .ZN(n19757) );
  INV_X1 U13272 ( .A(n19769), .ZN(n19777) );
  INV_X1 U13273 ( .A(n19801), .ZN(n19809) );
  INV_X1 U13274 ( .A(n19816), .ZN(n19827) );
  INV_X1 U13275 ( .A(n19927), .ZN(n19842) );
  INV_X1 U13276 ( .A(n19957), .ZN(n19857) );
  AOI21_X1 U13277 ( .B1(n19874), .B2(n19878), .A(n19872), .ZN(n19908) );
  NAND2_X1 U13278 ( .A1(n19441), .A2(n19914), .ZN(n19970) );
  OR4_X1 U13279 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), 
        .A3(P2_STATEBS16_REG_SCAN_IN), .A4(n10677), .ZN(n19977) );
  NAND2_X1 U13280 ( .A1(n19131), .A2(n18974), .ZN(n16787) );
  INV_X1 U13281 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17839) );
  INV_X1 U13282 ( .A(n17196), .ZN(n17182) );
  INV_X1 U13283 ( .A(n17195), .ZN(n17188) );
  NOR2_X1 U13284 ( .A1(n16953), .A2(n17306), .ZN(n17319) );
  AND2_X1 U13285 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17349), .ZN(n17361) );
  NOR2_X1 U13286 ( .A1(n17751), .A2(n17619), .ZN(n17622) );
  NOR2_X1 U13287 ( .A1(n15900), .A2(n15899), .ZN(n17635) );
  INV_X1 U13288 ( .A(n17656), .ZN(n17651) );
  INV_X1 U13289 ( .A(n17679), .ZN(n17698) );
  INV_X1 U13290 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17733) );
  INV_X1 U13291 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18190) );
  NAND2_X1 U13292 ( .A1(n18136), .A2(n16666), .ZN(n18052) );
  INV_X1 U13293 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18082) );
  NAND2_X1 U13294 ( .A1(n18766), .A2(n18535), .ZN(n18819) );
  INV_X1 U13295 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18238) );
  INV_X1 U13296 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18272) );
  NAND3_X1 U13297 ( .A1(n18919), .A2(n18391), .A3(n16666), .ZN(n18388) );
  NAND2_X1 U13298 ( .A1(n18447), .A2(n18459), .ZN(n18460) );
  AND2_X1 U13299 ( .A1(n19146), .A2(n16782), .ZN(n19130) );
  INV_X1 U13300 ( .A(n18793), .ZN(n18862) );
  INV_X1 U13301 ( .A(n18840), .ZN(n18902) );
  INV_X1 U13302 ( .A(n19131), .ZN(n18983) );
  INV_X1 U13303 ( .A(n19083), .ZN(n18992) );
  CLKBUF_X1 U13304 ( .A(n18992), .Z(n19080) );
  INV_X1 U13305 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n19009) );
  NAND2_X1 U13306 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n19007), .ZN(n19144) );
  NOR2_X1 U13307 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12882), .ZN(n16768)
         );
  INV_X1 U13308 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20001) );
  OR2_X1 U13309 ( .A1(n11004), .A2(n11003), .ZN(P2_U2824) );
  INV_X1 U13310 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10291) );
  INV_X1 U13311 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15295) );
  INV_X1 U13312 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14840) );
  NAND2_X1 U13313 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n10305), .ZN(
        n10304) );
  NAND2_X1 U13314 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n10307), .ZN(
        n10306) );
  NAND2_X1 U13315 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n10310), .ZN(
        n10314) );
  INV_X1 U13316 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n10289) );
  INV_X1 U13317 ( .A(n10324), .ZN(n10294) );
  INV_X1 U13318 ( .A(n10292), .ZN(n10297) );
  INV_X1 U13319 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14829) );
  NAND2_X1 U13320 ( .A1(n10297), .A2(n14829), .ZN(n10293) );
  NAND2_X1 U13321 ( .A1(n10294), .A2(n10293), .ZN(n15313) );
  INV_X1 U13322 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10752) );
  INV_X1 U13323 ( .A(n10295), .ZN(n10298) );
  NAND2_X1 U13324 ( .A1(n10752), .A2(n10298), .ZN(n10296) );
  NAND2_X1 U13325 ( .A1(n10297), .A2(n10296), .ZN(n16057) );
  NAND2_X1 U13326 ( .A1(n14840), .A2(n10300), .ZN(n10299) );
  AND2_X1 U13327 ( .A1(n10299), .A2(n10298), .ZN(n14846) );
  INV_X1 U13328 ( .A(n14846), .ZN(n15336) );
  OAI21_X1 U13329 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n10320), .A(
        n10300), .ZN(n15348) );
  INV_X1 U13330 ( .A(n15348), .ZN(n19186) );
  OAI21_X1 U13331 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n9759), .A(
        n10321), .ZN(n15367) );
  INV_X1 U13332 ( .A(n15367), .ZN(n19214) );
  OAI21_X1 U13333 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n10315), .A(
        n10318), .ZN(n15374) );
  INV_X1 U13334 ( .A(n15374), .ZN(n19237) );
  OAI21_X1 U13335 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n10313), .A(
        n10316), .ZN(n16446) );
  INV_X1 U13336 ( .A(n16446), .ZN(n19261) );
  OAI21_X1 U13337 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n10310), .A(
        n10314), .ZN(n19267) );
  INV_X1 U13338 ( .A(n19267), .ZN(n10312) );
  OAI21_X1 U13339 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n10308), .A(
        n10311), .ZN(n16490) );
  INV_X1 U13340 ( .A(n16490), .ZN(n14869) );
  OAI21_X1 U13341 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n10301), .A(
        n10309), .ZN(n15389) );
  INV_X1 U13342 ( .A(n15389), .ZN(n19295) );
  AOI21_X1 U13343 ( .B1(n15411), .B2(n10304), .A(n10307), .ZN(n19312) );
  AOI21_X1 U13344 ( .B1(n19439), .B2(n10302), .A(n10305), .ZN(n19425) );
  AOI21_X1 U13345 ( .B1(n14954), .B2(n14943), .A(n10303), .ZN(n14941) );
  AOI22_X1 U13346 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n19974), .ZN(n19340) );
  AOI22_X1 U13347 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n14954), .B2(n19974), .ZN(
        n14960) );
  NAND2_X1 U13348 ( .A1(n19340), .A2(n14960), .ZN(n14959) );
  NOR2_X1 U13349 ( .A1(n14941), .A2(n14959), .ZN(n14929) );
  OAI21_X1 U13350 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n10303), .A(
        n10302), .ZN(n14930) );
  NAND2_X1 U13351 ( .A1(n14929), .A2(n14930), .ZN(n14918) );
  NOR2_X1 U13352 ( .A1(n19425), .A2(n14918), .ZN(n14906) );
  OAI21_X1 U13353 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n10305), .A(
        n10304), .ZN(n15424) );
  NAND2_X1 U13354 ( .A1(n14906), .A2(n15424), .ZN(n19309) );
  NOR2_X1 U13355 ( .A1(n19312), .A2(n19309), .ZN(n14895) );
  OAI21_X1 U13356 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n10307), .A(
        n10306), .ZN(n15401) );
  NAND2_X1 U13357 ( .A1(n14895), .A2(n15401), .ZN(n19293) );
  NOR2_X1 U13358 ( .A1(n19295), .A2(n19293), .ZN(n14884) );
  AOI21_X1 U13359 ( .B1(n16500), .B2(n10309), .A(n10308), .ZN(n16492) );
  INV_X1 U13360 ( .A(n16492), .ZN(n14885) );
  NAND2_X1 U13361 ( .A1(n14884), .A2(n14885), .ZN(n14867) );
  NOR2_X1 U13362 ( .A1(n14869), .A2(n14867), .ZN(n19286) );
  AOI21_X1 U13363 ( .B1(n16476), .B2(n10311), .A(n10310), .ZN(n16464) );
  INV_X1 U13364 ( .A(n16464), .ZN(n19289) );
  NAND2_X1 U13365 ( .A1(n19286), .A2(n19289), .ZN(n19266) );
  NOR2_X1 U13366 ( .A1(n10312), .A2(n19266), .ZN(n14851) );
  AOI21_X1 U13367 ( .B1(n16458), .B2(n10314), .A(n10313), .ZN(n16447) );
  INV_X1 U13368 ( .A(n16447), .ZN(n14852) );
  NAND2_X1 U13369 ( .A1(n14851), .A2(n14852), .ZN(n19259) );
  NOR2_X1 U13370 ( .A1(n19261), .A2(n19259), .ZN(n19243) );
  AOI21_X1 U13371 ( .B1(n19249), .B2(n10316), .A(n10315), .ZN(n19246) );
  INV_X1 U13372 ( .A(n19246), .ZN(n10317) );
  NAND2_X1 U13373 ( .A1(n19243), .A2(n10317), .ZN(n19235) );
  NOR2_X1 U13374 ( .A1(n19237), .A2(n19235), .ZN(n19220) );
  AOI21_X1 U13375 ( .B1(n16428), .B2(n10318), .A(n9759), .ZN(n19222) );
  INV_X1 U13376 ( .A(n19222), .ZN(n10319) );
  NAND2_X1 U13377 ( .A1(n19220), .A2(n10319), .ZN(n19212) );
  NOR2_X1 U13378 ( .A1(n19214), .A2(n19212), .ZN(n19194) );
  AOI21_X1 U13379 ( .B1(n10321), .B2(n19197), .A(n10320), .ZN(n19196) );
  INV_X1 U13380 ( .A(n19196), .ZN(n10322) );
  NAND2_X1 U13381 ( .A1(n19194), .A2(n10322), .ZN(n19180) );
  NAND2_X1 U13382 ( .A1(n15336), .A2(n19179), .ZN(n10323) );
  NAND2_X1 U13383 ( .A1(n10323), .A2(n19310), .ZN(n16056) );
  NAND2_X1 U13384 ( .A1(n16057), .A2(n16056), .ZN(n16055) );
  NAND2_X1 U13385 ( .A1(n19310), .A2(n16055), .ZN(n14823) );
  NAND2_X1 U13386 ( .A1(n15313), .A2(n14823), .ZN(n14822) );
  NAND2_X1 U13387 ( .A1(n19310), .A2(n14822), .ZN(n16410) );
  OAI21_X1 U13388 ( .B1(n10324), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n10325), .ZN(n16411) );
  NAND2_X1 U13389 ( .A1(n19310), .A2(n16409), .ZN(n16399) );
  AOI21_X1 U13390 ( .B1(n10325), .B2(n15295), .A(n9802), .ZN(n15297) );
  INV_X1 U13391 ( .A(n15297), .ZN(n16400) );
  NAND2_X1 U13392 ( .A1(n19310), .A2(n16398), .ZN(n16388) );
  OAI21_X1 U13393 ( .B1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n9802), .A(
        n10326), .ZN(n16389) );
  NAND2_X1 U13394 ( .A1(n19310), .A2(n16387), .ZN(n16377) );
  AOI21_X1 U13395 ( .B1(n15273), .B2(n10326), .A(n10327), .ZN(n15271) );
  INV_X1 U13396 ( .A(n15271), .ZN(n16378) );
  NAND2_X1 U13397 ( .A1(n19310), .A2(n16376), .ZN(n16365) );
  OAI21_X1 U13398 ( .B1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n10327), .A(
        n10328), .ZN(n16366) );
  NAND2_X1 U13399 ( .A1(n19310), .A2(n16364), .ZN(n16352) );
  AOI21_X1 U13400 ( .B1(n10328), .B2(n10159), .A(n9801), .ZN(n15250) );
  INV_X1 U13401 ( .A(n15250), .ZN(n16353) );
  NAND2_X1 U13402 ( .A1(n19310), .A2(n16351), .ZN(n14809) );
  XNOR2_X1 U13403 ( .A(n9801), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14808) );
  INV_X2 U13404 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n10677) );
  INV_X2 U13405 ( .A(n19977), .ZN(n19315) );
  NAND2_X1 U13406 ( .A1(n19315), .A2(n19310), .ZN(n19339) );
  NAND2_X1 U13407 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20079), .ZN(
        n10338) );
  NAND2_X1 U13408 ( .A1(n10341), .A2(n10338), .ZN(n10330) );
  NAND2_X1 U13409 ( .A1(n13522), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10339) );
  MUX2_X1 U13410 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n10331), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10335) );
  NAND2_X1 U13411 ( .A1(n10331), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10332) );
  NOR2_X1 U13412 ( .A1(n16121), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10334) );
  NAND2_X1 U13413 ( .A1(n10344), .A2(n10334), .ZN(n10536) );
  INV_X1 U13414 ( .A(n10335), .ZN(n10336) );
  XNOR2_X1 U13415 ( .A(n10337), .B(n10336), .ZN(n10523) );
  AND2_X1 U13416 ( .A1(n10339), .A2(n10338), .ZN(n10340) );
  XNOR2_X1 U13417 ( .A(n10341), .B(n10340), .ZN(n12737) );
  INV_X1 U13418 ( .A(n12737), .ZN(n10342) );
  XNOR2_X1 U13419 ( .A(n12747), .B(n12322), .ZN(n12324) );
  NOR2_X1 U13420 ( .A1(n10342), .A2(n12324), .ZN(n10343) );
  NAND2_X1 U13421 ( .A1(n12738), .A2(n10343), .ZN(n10349) );
  NAND2_X1 U13422 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n15859), .ZN(
        n10345) );
  NAND2_X1 U13423 ( .A1(n16121), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10347) );
  INV_X1 U13424 ( .A(n12334), .ZN(n12751) );
  NAND2_X1 U13425 ( .A1(n10677), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19980) );
  NAND2_X2 U13426 ( .A1(n10351), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10487) );
  NAND2_X2 U13427 ( .A1(n10350), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12133) );
  AOI22_X1 U13428 ( .A1(n12308), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10488), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10356) );
  INV_X2 U13429 ( .A(n12307), .ZN(n12299) );
  AOI22_X1 U13430 ( .A1(n10371), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9640), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10355) );
  INV_X2 U13431 ( .A(n12132), .ZN(n10450) );
  NAND2_X4 U13432 ( .A1(n13521), .A2(n13522), .ZN(n12266) );
  AOI22_X1 U13433 ( .A1(n10450), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9643), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10354) );
  AOI22_X1 U13434 ( .A1(n10372), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12287), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10353) );
  AOI22_X1 U13435 ( .A1(n10372), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12287), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10359) );
  AOI22_X1 U13436 ( .A1(n12299), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__5__SCAN_IN), .B2(n10371), .ZN(n10358) );
  AOI22_X1 U13437 ( .A1(n12308), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10488), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10363) );
  AOI22_X1 U13438 ( .A1(n10450), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9642), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10362) );
  AOI22_X1 U13439 ( .A1(n10450), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9671), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10367) );
  AOI22_X1 U13440 ( .A1(n12308), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10488), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10366) );
  AOI22_X1 U13441 ( .A1(n10371), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9641), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10365) );
  AOI22_X1 U13442 ( .A1(n10372), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12287), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10364) );
  NAND4_X1 U13443 ( .A1(n10367), .A2(n10366), .A3(n10365), .A4(n10364), .ZN(
        n10368) );
  NAND2_X1 U13444 ( .A1(n10368), .A2(n10489), .ZN(n10369) );
  NAND2_X1 U13445 ( .A1(n10371), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10376) );
  NAND2_X1 U13446 ( .A1(n12299), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10375) );
  CLKBUF_X2 U13447 ( .A(n10372), .Z(n12171) );
  NAND2_X1 U13448 ( .A1(n10372), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10374) );
  NAND2_X1 U13449 ( .A1(n12287), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10373) );
  INV_X1 U13450 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12237) );
  INV_X1 U13451 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10377) );
  OAI22_X1 U13452 ( .A1(n10487), .A2(n12237), .B1(n12133), .B2(n10377), .ZN(
        n10378) );
  INV_X1 U13453 ( .A(n10378), .ZN(n10382) );
  INV_X1 U13454 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10379) );
  OAI22_X1 U13455 ( .A1(n12132), .A2(n12238), .B1(n12266), .B2(n10379), .ZN(
        n10380) );
  INV_X1 U13456 ( .A(n10380), .ZN(n10381) );
  NAND2_X1 U13457 ( .A1(n10371), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10388) );
  NAND2_X1 U13458 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10387) );
  NAND2_X1 U13459 ( .A1(n10372), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10386) );
  NAND2_X1 U13460 ( .A1(n12287), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10385) );
  NAND4_X1 U13461 ( .A1(n10388), .A2(n10387), .A3(n10386), .A4(n10385), .ZN(
        n10396) );
  INV_X1 U13462 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12248) );
  INV_X1 U13463 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10389) );
  OAI22_X1 U13464 ( .A1(n10487), .A2(n12248), .B1(n12133), .B2(n10389), .ZN(
        n10390) );
  INV_X1 U13465 ( .A(n10390), .ZN(n10394) );
  INV_X1 U13466 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12246) );
  INV_X1 U13467 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10391) );
  OAI22_X1 U13468 ( .A1(n12132), .A2(n12246), .B1(n12266), .B2(n10391), .ZN(
        n10392) );
  INV_X1 U13469 ( .A(n10392), .ZN(n10393) );
  NAND2_X1 U13470 ( .A1(n10394), .A2(n10393), .ZN(n10395) );
  NOR2_X1 U13471 ( .A1(n10396), .A2(n10395), .ZN(n10397) );
  AOI22_X1 U13472 ( .A1(n12308), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10488), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10403) );
  AOI22_X1 U13473 ( .A1(n10450), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9671), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10402) );
  AOI22_X1 U13474 ( .A1(n10371), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9641), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10401) );
  AOI22_X1 U13475 ( .A1(n10372), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12287), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10400) );
  NAND4_X1 U13476 ( .A1(n10403), .A2(n10402), .A3(n10401), .A4(n10400), .ZN(
        n10404) );
  NAND2_X1 U13477 ( .A1(n10404), .A2(n10489), .ZN(n10411) );
  AOI22_X1 U13478 ( .A1(n12308), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10488), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10408) );
  AOI22_X1 U13479 ( .A1(n10450), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9643), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10407) );
  AOI22_X1 U13480 ( .A1(n10372), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12287), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10406) );
  AOI22_X1 U13481 ( .A1(n10371), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9640), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10405) );
  NAND4_X1 U13482 ( .A1(n10408), .A2(n10407), .A3(n10406), .A4(n10405), .ZN(
        n10409) );
  NAND2_X1 U13483 ( .A1(n10409), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10410) );
  NAND2_X1 U13484 ( .A1(n10411), .A2(n10410), .ZN(n10455) );
  NAND4_X1 U13485 ( .A1(n10631), .A2(n10606), .A3(n10647), .A4(n12777), .ZN(
        n10442) );
  NAND2_X1 U13486 ( .A1(n10371), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n10415) );
  NAND2_X1 U13487 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n10414) );
  NAND2_X1 U13488 ( .A1(n10372), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10413) );
  NAND2_X1 U13489 ( .A1(n12287), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10412) );
  NAND4_X1 U13490 ( .A1(n10415), .A2(n10414), .A3(n10413), .A4(n10412), .ZN(
        n10419) );
  OAI22_X1 U13491 ( .A1(n10487), .A2(n12482), .B1(n12133), .B2(n12470), .ZN(
        n10417) );
  OAI22_X1 U13492 ( .A1(n12132), .A2(n12462), .B1(n12266), .B2(n12468), .ZN(
        n10416) );
  NOR2_X1 U13493 ( .A1(n10419), .A2(n10418), .ZN(n10420) );
  NAND2_X1 U13494 ( .A1(n10420), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10430) );
  OAI22_X1 U13495 ( .A1(n10487), .A2(n12481), .B1(n12133), .B2(n12465), .ZN(
        n10421) );
  NAND2_X1 U13496 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n10425) );
  NAND2_X1 U13497 ( .A1(n12287), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n10424) );
  NAND2_X1 U13498 ( .A1(n10372), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n10423) );
  NAND3_X1 U13499 ( .A1(n10425), .A2(n10424), .A3(n10423), .ZN(n10426) );
  NOR2_X1 U13500 ( .A1(n10426), .A2(n10274), .ZN(n10427) );
  NAND3_X1 U13501 ( .A1(n10428), .A2(n10427), .A3(n10489), .ZN(n10429) );
  AOI22_X1 U13502 ( .A1(n10450), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9642), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10434) );
  AOI22_X1 U13503 ( .A1(n12308), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10488), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10433) );
  AOI22_X1 U13504 ( .A1(n10371), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12299), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10432) );
  AOI22_X1 U13505 ( .A1(n10372), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12287), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10431) );
  NAND4_X1 U13506 ( .A1(n10434), .A2(n10433), .A3(n10432), .A4(n10431), .ZN(
        n10435) );
  AOI22_X1 U13507 ( .A1(n10371), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12299), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10436) );
  AOI22_X1 U13508 ( .A1(n12308), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10488), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10438) );
  AOI22_X1 U13509 ( .A1(n10450), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9671), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10437) );
  NAND2_X1 U13510 ( .A1(n10439), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10440) );
  AOI22_X1 U13511 ( .A1(n10450), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12308), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10446) );
  AOI22_X1 U13512 ( .A1(n10371), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12299), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10445) );
  AOI22_X1 U13513 ( .A1(n10372), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12287), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10443) );
  AOI22_X1 U13514 ( .A1(n10372), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12287), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10449) );
  AOI22_X1 U13515 ( .A1(n10371), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12299), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10448) );
  AOI22_X1 U13516 ( .A1(n12308), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10488), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10451) );
  INV_X1 U13517 ( .A(n10456), .ZN(n12796) );
  NOR2_X1 U13518 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20059) );
  INV_X1 U13519 ( .A(n20059), .ZN(n20065) );
  NOR2_X1 U13520 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20065), .ZN(n10457) );
  AND2_X2 U13521 ( .A1(n10457), .A2(n19974), .ZN(n19427) );
  INV_X2 U13522 ( .A(n19427), .ZN(n19300) );
  NAND2_X1 U13523 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19591), .ZN(n19972) );
  NOR2_X1 U13524 ( .A1(n19980), .A2(n19972), .ZN(n16599) );
  NOR2_X1 U13525 ( .A1(n19315), .A2(n16599), .ZN(n10458) );
  NAND2_X1 U13526 ( .A1(n19300), .A2(n10458), .ZN(n10459) );
  INV_X1 U13527 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n20042) );
  NAND2_X1 U13528 ( .A1(n10371), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10463) );
  NAND2_X1 U13529 ( .A1(n12299), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10462) );
  NAND2_X1 U13530 ( .A1(n10372), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10461) );
  NAND2_X1 U13531 ( .A1(n12287), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10460) );
  NAND4_X1 U13532 ( .A1(n10463), .A2(n10462), .A3(n10461), .A4(n10460), .ZN(
        n10467) );
  OAI22_X1 U13533 ( .A1(n12132), .A2(n12440), .B1(n12133), .B2(n12430), .ZN(
        n10465) );
  OAI22_X1 U13534 ( .A1(n10487), .A2(n15754), .B1(n12266), .B2(n12432), .ZN(
        n10464) );
  NOR2_X1 U13535 ( .A1(n10467), .A2(n10466), .ZN(n10468) );
  NAND2_X1 U13536 ( .A1(n10468), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10479) );
  NAND2_X1 U13537 ( .A1(n10371), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10472) );
  NAND2_X1 U13538 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10471) );
  NAND2_X1 U13539 ( .A1(n10372), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10470) );
  NAND2_X1 U13540 ( .A1(n12287), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10469) );
  NAND4_X1 U13541 ( .A1(n10472), .A2(n10471), .A3(n10470), .A4(n10469), .ZN(
        n10476) );
  OAI22_X1 U13542 ( .A1(n12132), .A2(n12441), .B1(n12266), .B2(n12453), .ZN(
        n10474) );
  OAI22_X1 U13543 ( .A1(n10487), .A2(n12437), .B1(n12133), .B2(n12438), .ZN(
        n10473) );
  OR2_X1 U13544 ( .A1(n10474), .A2(n10473), .ZN(n10475) );
  NOR2_X1 U13545 ( .A1(n10476), .A2(n10475), .ZN(n10477) );
  NAND2_X1 U13546 ( .A1(n10477), .A2(n10489), .ZN(n10478) );
  NAND2_X1 U13547 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20114) );
  INV_X1 U13548 ( .A(n20114), .ZN(n20118) );
  NOR2_X1 U13549 ( .A1(n20118), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n14810) );
  INV_X1 U13550 ( .A(n14810), .ZN(n10787) );
  NAND2_X1 U13551 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n10787), .ZN(n10480) );
  NOR2_X1 U13552 ( .A1(n12765), .A2(n10480), .ZN(n10481) );
  AOI22_X1 U13553 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n12150), .B1(
        n12087), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10495) );
  AND2_X2 U13554 ( .A1(n9641), .A2(n10489), .ZN(n12151) );
  AOI22_X1 U13555 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n12151), .B1(
        n12088), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10482) );
  INV_X1 U13556 ( .A(n10482), .ZN(n10486) );
  AND2_X2 U13557 ( .A1(n12287), .A2(n10489), .ZN(n10806) );
  AOI22_X1 U13558 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12152), .B1(
        n10806), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10484) );
  AND2_X2 U13559 ( .A1(n12171), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10552) );
  AOI22_X1 U13560 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10811), .B1(
        n10552), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10483) );
  INV_X2 U13561 ( .A(n10867), .ZN(n12157) );
  AND2_X2 U13562 ( .A1(n12309), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10558) );
  AOI22_X1 U13563 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12157), .B1(
        n10558), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10493) );
  AOI22_X1 U13564 ( .A1(n10501), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10492) );
  OR2_X1 U13565 ( .A1(n12282), .A2(n10489), .ZN(n10868) );
  INV_X2 U13566 ( .A(n10868), .ZN(n12158) );
  AOI22_X1 U13567 ( .A1(n12158), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10491) );
  AOI22_X1 U13568 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10544), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10490) );
  NAND3_X1 U13569 ( .A1(n10495), .A2(n10494), .A3(n10281), .ZN(n12460) );
  MUX2_X1 U13570 ( .A(n12460), .B(n12737), .S(n12765), .Z(n12745) );
  INV_X1 U13571 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n14944) );
  INV_X1 U13572 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n14953) );
  NOR2_X1 U13573 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), 
        .ZN(n10509) );
  AOI22_X1 U13574 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12150), .B1(
        n12088), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10499) );
  AOI22_X1 U13575 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12151), .B1(
        n12087), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10498) );
  AOI22_X1 U13576 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10811), .B1(
        n10552), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10497) );
  AOI22_X1 U13577 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12152), .B1(
        n10806), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10496) );
  NAND4_X1 U13578 ( .A1(n10499), .A2(n10498), .A3(n10497), .A4(n10496), .ZN(
        n10507) );
  INV_X1 U13579 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12447) );
  INV_X1 U13580 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12426) );
  OAI22_X1 U13581 ( .A1(n12447), .A2(n10867), .B1(n10868), .B2(n12426), .ZN(
        n10500) );
  INV_X1 U13582 ( .A(n10500), .ZN(n10505) );
  AOI22_X1 U13583 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10544), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10504) );
  AOI22_X1 U13584 ( .A1(n10501), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10503) );
  AOI22_X1 U13585 ( .A1(n10558), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10502) );
  NAND4_X1 U13586 ( .A1(n10505), .A2(n10504), .A3(n10503), .A4(n10502), .ZN(
        n10506) );
  MUX2_X1 U13587 ( .A(n10509), .B(n12815), .S(n10508), .Z(n12507) );
  NAND2_X1 U13588 ( .A1(n12508), .A2(n12507), .ZN(n12506) );
  INV_X1 U13589 ( .A(n12506), .ZN(n10525) );
  AOI22_X1 U13590 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12088), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10513) );
  AOI22_X1 U13591 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12087), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10512) );
  AOI22_X1 U13592 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10811), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10511) );
  AOI22_X1 U13593 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12152), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10510) );
  NAND4_X1 U13594 ( .A1(n10513), .A2(n10512), .A3(n10511), .A4(n10510), .ZN(
        n10522) );
  AOI22_X1 U13595 ( .A1(n12158), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12157), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10520) );
  AOI22_X1 U13596 ( .A1(n10501), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10519) );
  AOI22_X1 U13597 ( .A1(n10558), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10518) );
  AOI22_X1 U13598 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10517) );
  NAND4_X1 U13599 ( .A1(n10520), .A2(n10519), .A3(n10518), .A4(n10517), .ZN(
        n10521) );
  MUX2_X1 U13600 ( .A(n12490), .B(n10523), .S(n12765), .Z(n12320) );
  INV_X1 U13601 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n10524) );
  MUX2_X1 U13602 ( .A(n12320), .B(n10524), .S(n12727), .Z(n12496) );
  NAND2_X1 U13603 ( .A1(n10525), .A2(n12496), .ZN(n12511) );
  AOI22_X1 U13604 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12088), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10529) );
  AOI22_X1 U13605 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12087), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10528) );
  INV_X1 U13606 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12238) );
  AOI22_X1 U13607 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10811), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10527) );
  AOI22_X1 U13608 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12152), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10526) );
  NAND4_X1 U13609 ( .A1(n10529), .A2(n10528), .A3(n10527), .A4(n10526), .ZN(
        n10535) );
  AOI22_X1 U13610 ( .A1(n12158), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12157), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10533) );
  AOI22_X1 U13611 ( .A1(n10501), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10532) );
  AOI22_X1 U13612 ( .A1(n10558), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10531) );
  AOI22_X1 U13613 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10530) );
  NAND4_X1 U13614 ( .A1(n10533), .A2(n10532), .A3(n10531), .A4(n10530), .ZN(
        n10534) );
  MUX2_X1 U13615 ( .A(n10536), .B(n12827), .S(n20103), .Z(n12321) );
  INV_X1 U13616 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n10537) );
  MUX2_X1 U13617 ( .A(n12321), .B(n10537), .S(n12727), .Z(n10538) );
  INV_X1 U13618 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n10551) );
  AOI22_X1 U13619 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12088), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10542) );
  AOI22_X1 U13620 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12087), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10541) );
  AOI22_X1 U13621 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10811), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10540) );
  AOI22_X1 U13622 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12152), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10539) );
  NAND4_X1 U13623 ( .A1(n10542), .A2(n10541), .A3(n10540), .A4(n10539), .ZN(
        n10550) );
  INV_X1 U13624 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12528) );
  INV_X1 U13625 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12534) );
  OAI22_X1 U13626 ( .A1(n10868), .A2(n12528), .B1(n10867), .B2(n12534), .ZN(
        n10543) );
  INV_X1 U13627 ( .A(n10543), .ZN(n10548) );
  AOI22_X1 U13628 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10547) );
  AOI22_X1 U13629 ( .A1(n10501), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10546) );
  AOI22_X1 U13630 ( .A1(n10558), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10545) );
  NAND4_X1 U13631 ( .A1(n10548), .A2(n10547), .A3(n10546), .A4(n10545), .ZN(
        n10549) );
  MUX2_X1 U13632 ( .A(n10551), .B(n12552), .S(n10508), .Z(n12556) );
  NAND2_X1 U13633 ( .A1(n12557), .A2(n12556), .ZN(n12593) );
  AOI22_X1 U13634 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12150), .B1(
        n12088), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10556) );
  AOI22_X1 U13635 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n12151), .B1(
        n12087), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10555) );
  AOI22_X1 U13636 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10811), .B1(
        n10552), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10554) );
  AOI22_X1 U13637 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n10806), .B1(
        n12152), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10553) );
  NAND4_X1 U13638 ( .A1(n10556), .A2(n10555), .A3(n10554), .A4(n10553), .ZN(
        n10564) );
  INV_X1 U13639 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n15720) );
  INV_X1 U13640 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12572) );
  OAI22_X1 U13641 ( .A1(n15720), .A2(n10867), .B1(n10868), .B2(n12572), .ZN(
        n10557) );
  INV_X1 U13642 ( .A(n10557), .ZN(n10562) );
  AOI22_X1 U13643 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10544), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10561) );
  AOI22_X1 U13644 ( .A1(n10501), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10560) );
  AOI22_X1 U13645 ( .A1(n10558), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10559) );
  NAND4_X1 U13646 ( .A1(n10562), .A2(n10561), .A3(n10560), .A4(n10559), .ZN(
        n10563) );
  MUX2_X1 U13647 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n12589), .S(n10508), .Z(
        n12592) );
  INV_X1 U13648 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n10585) );
  NAND2_X1 U13649 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10568) );
  NAND2_X1 U13650 ( .A1(n12088), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10567) );
  NAND2_X1 U13651 ( .A1(n12087), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10566) );
  NAND2_X1 U13652 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10565) );
  NAND2_X1 U13653 ( .A1(n12157), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10572) );
  NAND2_X1 U13654 ( .A1(n12158), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10571) );
  NAND2_X1 U13655 ( .A1(n10501), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10570) );
  NAND2_X1 U13656 ( .A1(n10514), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10569) );
  NAND2_X1 U13657 ( .A1(n10558), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10576) );
  NAND2_X1 U13658 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10575) );
  NAND2_X1 U13659 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10574) );
  NAND2_X1 U13660 ( .A1(n10516), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10573) );
  NAND2_X1 U13661 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10580) );
  NAND2_X1 U13662 ( .A1(n10811), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10579) );
  NAND2_X1 U13663 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10578) );
  NAND2_X1 U13664 ( .A1(n12152), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10577) );
  NAND4_X1 U13665 ( .A1(n10584), .A2(n10583), .A3(n10582), .A4(n10581), .ZN(
        n10861) );
  MUX2_X1 U13666 ( .A(n10585), .B(n10861), .S(n10508), .Z(n12603) );
  INV_X1 U13667 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n19291) );
  NOR2_X1 U13668 ( .A1(n10508), .A2(n19291), .ZN(n12600) );
  INV_X1 U13669 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n15115) );
  INV_X1 U13670 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n15104) );
  NAND2_X1 U13671 ( .A1(n12617), .A2(n15104), .ZN(n12627) );
  NAND2_X1 U13672 ( .A1(n12706), .A2(n12627), .ZN(n12621) );
  NAND2_X1 U13673 ( .A1(n12727), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10587) );
  INV_X1 U13674 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n10725) );
  NOR2_X1 U13675 ( .A1(n10508), .A2(n10725), .ZN(n12648) );
  INV_X1 U13676 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n10729) );
  NAND2_X1 U13677 ( .A1(n12727), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n12642) );
  INV_X1 U13678 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n15072) );
  INV_X1 U13679 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n10588) );
  AND2_X1 U13680 ( .A1(n15072), .A2(n10588), .ZN(n10589) );
  NOR2_X1 U13681 ( .A1(n10508), .A2(n10589), .ZN(n10590) );
  INV_X1 U13682 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n19208) );
  NOR2_X1 U13683 ( .A1(n10508), .A2(n19208), .ZN(n12654) );
  NOR2_X2 U13684 ( .A1(n12659), .A2(n12654), .ZN(n12656) );
  NAND2_X1 U13685 ( .A1(n12727), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n12639) );
  INV_X1 U13686 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n19181) );
  NAND2_X1 U13687 ( .A1(n12727), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12686) );
  INV_X1 U13688 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n10591) );
  NOR2_X1 U13689 ( .A1(n10508), .A2(n10591), .ZN(n12693) );
  INV_X1 U13690 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n10592) );
  NAND2_X1 U13691 ( .A1(n12727), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12711) );
  INV_X1 U13692 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n10772) );
  NOR2_X1 U13693 ( .A1(n10508), .A2(n10772), .ZN(n12717) );
  NAND2_X1 U13694 ( .A1(n12727), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12724) );
  NAND2_X1 U13695 ( .A1(n12725), .A2(n12724), .ZN(n12729) );
  NOR2_X1 U13696 ( .A1(n12729), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10594) );
  MUX2_X1 U13697 ( .A(n12710), .B(n10594), .S(n12727), .Z(n14088) );
  INV_X1 U13698 ( .A(n14088), .ZN(n10598) );
  INV_X1 U13699 ( .A(n10595), .ZN(n10596) );
  NAND2_X2 U13700 ( .A1(n20034), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n20038) );
  INV_X1 U13701 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19156) );
  NAND2_X1 U13702 ( .A1(n19156), .A2(n19997), .ZN(n19991) );
  NAND3_X1 U13703 ( .A1(n19986), .A2(n20038), .A3(n19991), .ZN(n19985) );
  NAND2_X1 U13704 ( .A1(n20123), .A2(n20114), .ZN(n12735) );
  NOR2_X1 U13705 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n12735), .ZN(n13509) );
  INV_X1 U13706 ( .A(n13509), .ZN(n10597) );
  NAND2_X1 U13707 ( .A1(n12949), .A2(n10597), .ZN(n14813) );
  INV_X1 U13708 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n10783) );
  OAI222_X1 U13709 ( .A1(n19301), .A2(n20042), .B1(n19304), .B2(n10598), .C1(
        n14813), .C2(n10783), .ZN(n10600) );
  NOR2_X2 U13710 ( .A1(n19325), .A2(n20089), .ZN(n19308) );
  AND2_X1 U13711 ( .A1(n19308), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10599) );
  NAND2_X1 U13712 ( .A1(n12012), .A2(n10631), .ZN(n10646) );
  NOR2_X1 U13713 ( .A1(n10646), .A2(n19459), .ZN(n10602) );
  NAND3_X1 U13714 ( .A1(n12347), .A2(n10640), .A3(n19486), .ZN(n10603) );
  NAND2_X2 U13715 ( .A1(n10604), .A2(n10603), .ZN(n10650) );
  NAND2_X1 U13716 ( .A1(n10650), .A2(n15751), .ZN(n10613) );
  NAND3_X1 U13717 ( .A1(n10631), .A2(n20115), .A3(n10606), .ZN(n10607) );
  NAND2_X2 U13718 ( .A1(n10606), .A2(n10605), .ZN(n10819) );
  INV_X1 U13719 ( .A(n12329), .ZN(n10609) );
  NAND2_X1 U13720 ( .A1(n10609), .A2(n10608), .ZN(n12346) );
  AND2_X1 U13721 ( .A1(n12732), .A2(n19486), .ZN(n10610) );
  NOR2_X1 U13722 ( .A1(n12771), .A2(n19459), .ZN(n10612) );
  NAND2_X1 U13723 ( .A1(n12409), .A2(n10612), .ZN(n10668) );
  NAND2_X1 U13724 ( .A1(n10613), .A2(n10668), .ZN(n12811) );
  BUF_X1 U13725 ( .A(n10654), .Z(n10614) );
  NAND2_X1 U13726 ( .A1(n12775), .A2(n10640), .ZN(n12348) );
  INV_X1 U13727 ( .A(n12348), .ZN(n10616) );
  NAND3_X1 U13728 ( .A1(n10616), .A2(n12777), .A3(n20103), .ZN(n12782) );
  NOR2_X2 U13729 ( .A1(n12782), .A2(n19974), .ZN(n10679) );
  INV_X1 U13730 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n10619) );
  AOI22_X1 U13731 ( .A1(n10680), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n10618) );
  OAI21_X1 U13732 ( .B1(n10784), .B2(n10619), .A(n10618), .ZN(n10620) );
  AOI21_X1 U13733 ( .B1(n10780), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n10620), .ZN(n14965) );
  INV_X1 U13734 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15624) );
  OR2_X1 U13735 ( .A1(n10774), .A2(n15624), .ZN(n10623) );
  INV_X1 U13736 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n15625) );
  OAI22_X1 U13737 ( .A1(n10775), .A2(n15625), .B1(n10677), .B2(n16500), .ZN(
        n10621) );
  AOI21_X1 U13738 ( .B1(n10777), .B2(P2_EBX_REG_9__SCAN_IN), .A(n10621), .ZN(
        n10622) );
  NAND2_X1 U13739 ( .A1(n10623), .A2(n10622), .ZN(n13598) );
  NOR2_X1 U13740 ( .A1(n10654), .A2(n15692), .ZN(n10629) );
  INV_X1 U13741 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n10624) );
  INV_X1 U13742 ( .A(n10625), .ZN(n10626) );
  NAND2_X1 U13743 ( .A1(n10627), .A2(n10626), .ZN(n10628) );
  NOR2_X1 U13744 ( .A1(n10629), .A2(n10628), .ZN(n10672) );
  AOI21_X1 U13745 ( .B1(n10630), .B2(n19459), .A(n12733), .ZN(n10636) );
  MUX2_X1 U13746 ( .A(n12732), .B(n10631), .S(n12012), .Z(n10634) );
  NAND3_X1 U13747 ( .A1(n10634), .A2(n10633), .A3(n10632), .ZN(n10635) );
  NAND2_X1 U13748 ( .A1(n10819), .A2(n15751), .ZN(n12773) );
  NAND2_X1 U13749 ( .A1(n12773), .A2(n20115), .ZN(n10637) );
  NAND2_X1 U13750 ( .A1(n12780), .A2(n10637), .ZN(n10638) );
  NAND2_X1 U13751 ( .A1(n10638), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10645) );
  NOR2_X1 U13752 ( .A1(n19459), .A2(n10640), .ZN(n10641) );
  NOR2_X1 U13753 ( .A1(n19459), .A2(n15751), .ZN(n10642) );
  NAND2_X1 U13754 ( .A1(n12410), .A2(n13014), .ZN(n10644) );
  NAND2_X1 U13755 ( .A1(n10646), .A2(n10819), .ZN(n12336) );
  NAND2_X1 U13756 ( .A1(n12336), .A2(n10647), .ZN(n12337) );
  NAND2_X1 U13757 ( .A1(n10819), .A2(n12732), .ZN(n12341) );
  AND2_X1 U13758 ( .A1(n12341), .A2(n19486), .ZN(n10648) );
  NAND2_X1 U13759 ( .A1(n10661), .A2(n10665), .ZN(n10649) );
  NAND2_X1 U13760 ( .A1(n10676), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10652) );
  AOI22_X1 U13761 ( .A1(n13549), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n13510), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10651) );
  XNOR2_X1 U13762 ( .A(n10672), .B(n10671), .ZN(n12029) );
  INV_X1 U13763 ( .A(n10654), .ZN(n10655) );
  NAND2_X1 U13764 ( .A1(n10655), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10664) );
  INV_X1 U13765 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n10658) );
  INV_X1 U13766 ( .A(n13510), .ZN(n10657) );
  NAND2_X1 U13767 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10656) );
  OAI211_X1 U13768 ( .C1(n10659), .C2(n10658), .A(n10657), .B(n10656), .ZN(
        n10660) );
  AOI21_X1 U13769 ( .B1(n10679), .B2(P2_EBX_REG_0__SCAN_IN), .A(n10660), .ZN(
        n10663) );
  NAND3_X1 U13770 ( .A1(n10661), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n12773), 
        .ZN(n10662) );
  INV_X1 U13771 ( .A(n10665), .ZN(n10666) );
  NOR2_X1 U13772 ( .A1(n10666), .A2(n12771), .ZN(n10667) );
  OAI22_X1 U13773 ( .A1(n10676), .A2(n10667), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n10679), .ZN(n10670) );
  INV_X1 U13774 ( .A(n10668), .ZN(n13526) );
  AOI22_X1 U13775 ( .A1(n13526), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n13510), .ZN(n10669) );
  NAND2_X1 U13776 ( .A1(n10670), .A2(n10669), .ZN(n12033) );
  NAND2_X1 U13777 ( .A1(n12029), .A2(n12038), .ZN(n10675) );
  INV_X1 U13778 ( .A(n10671), .ZN(n10673) );
  NAND2_X1 U13779 ( .A1(n10673), .A2(n10672), .ZN(n10674) );
  OAI21_X1 U13780 ( .B1(n20079), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10677), 
        .ZN(n10678) );
  AOI22_X1 U13781 ( .A1(n10680), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10681) );
  OAI21_X1 U13782 ( .B1(n10784), .B2(n14944), .A(n10681), .ZN(n10682) );
  INV_X1 U13783 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12785) );
  INV_X1 U13784 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n10684) );
  INV_X1 U13785 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13706) );
  OAI22_X1 U13786 ( .A1(n10775), .A2(n10684), .B1(n10677), .B2(n13706), .ZN(
        n10685) );
  AOI21_X1 U13787 ( .B1(n10679), .B2(P2_EBX_REG_3__SCAN_IN), .A(n10685), .ZN(
        n10686) );
  NAND2_X1 U13788 ( .A1(n10676), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10689) );
  NAND2_X1 U13789 ( .A1(n13510), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10688) );
  XNOR2_X2 U13790 ( .A(n10691), .B(n10690), .ZN(n12011) );
  INV_X1 U13791 ( .A(n10690), .ZN(n10692) );
  NAND2_X1 U13792 ( .A1(n10692), .A2(n10691), .ZN(n10693) );
  NAND2_X1 U13793 ( .A1(n10694), .A2(n10693), .ZN(n13312) );
  INV_X1 U13794 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15676) );
  OR2_X1 U13795 ( .A1(n10774), .A2(n15676), .ZN(n10698) );
  INV_X1 U13796 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n10695) );
  OAI22_X1 U13797 ( .A1(n10775), .A2(n10695), .B1(n10677), .B2(n19439), .ZN(
        n10696) );
  AOI21_X1 U13798 ( .B1(n10777), .B2(P2_EBX_REG_4__SCAN_IN), .A(n10696), .ZN(
        n10697) );
  INV_X1 U13799 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15660) );
  OR2_X1 U13800 ( .A1(n10774), .A2(n15660), .ZN(n10702) );
  INV_X1 U13801 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n15426) );
  INV_X1 U13802 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10699) );
  OAI22_X1 U13803 ( .A1(n10775), .A2(n15426), .B1(n10677), .B2(n10699), .ZN(
        n10700) );
  AOI21_X1 U13804 ( .B1(n10777), .B2(P2_EBX_REG_5__SCAN_IN), .A(n10700), .ZN(
        n10701) );
  NAND2_X1 U13805 ( .A1(n10702), .A2(n10701), .ZN(n13320) );
  INV_X1 U13806 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12799) );
  OR2_X1 U13807 ( .A1(n10774), .A2(n12799), .ZN(n10705) );
  INV_X1 U13808 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n10860) );
  OAI22_X1 U13809 ( .A1(n10775), .A2(n10860), .B1(n10677), .B2(n15411), .ZN(
        n10703) );
  AOI21_X1 U13810 ( .B1(n10777), .B2(P2_EBX_REG_6__SCAN_IN), .A(n10703), .ZN(
        n10704) );
  NAND2_X1 U13811 ( .A1(n10705), .A2(n10704), .ZN(n13443) );
  INV_X1 U13812 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16558) );
  OR2_X1 U13813 ( .A1(n10774), .A2(n16558), .ZN(n10709) );
  INV_X1 U13814 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n15402) );
  INV_X1 U13815 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10706) );
  OAI22_X1 U13816 ( .A1(n10775), .A2(n15402), .B1(n10677), .B2(n10706), .ZN(
        n10707) );
  AOI21_X1 U13817 ( .B1(n10777), .B2(P2_EBX_REG_7__SCAN_IN), .A(n10707), .ZN(
        n10708) );
  NAND2_X1 U13818 ( .A1(n10709), .A2(n10708), .ZN(n13457) );
  INV_X1 U13819 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16561) );
  OR2_X1 U13820 ( .A1(n10774), .A2(n16561), .ZN(n10713) );
  INV_X1 U13821 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n10710) );
  OAI22_X1 U13822 ( .A1(n10775), .A2(n10710), .B1(n10677), .B2(n10170), .ZN(
        n10711) );
  AOI21_X1 U13823 ( .B1(n10777), .B2(P2_EBX_REG_8__SCAN_IN), .A(n10711), .ZN(
        n10712) );
  INV_X1 U13824 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16545) );
  OR2_X1 U13825 ( .A1(n10774), .A2(n16545), .ZN(n10716) );
  INV_X1 U13826 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n10905) );
  INV_X1 U13827 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n14873) );
  OAI22_X1 U13828 ( .A1(n10775), .A2(n10905), .B1(n10677), .B2(n14873), .ZN(
        n10714) );
  AOI21_X1 U13829 ( .B1(n10777), .B2(P2_EBX_REG_10__SCAN_IN), .A(n10714), .ZN(
        n10715) );
  OR2_X1 U13830 ( .A1(n10774), .A2(n16542), .ZN(n10720) );
  INV_X1 U13831 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n10717) );
  OAI22_X1 U13832 ( .A1(n10775), .A2(n10717), .B1(n10677), .B2(n16476), .ZN(
        n10718) );
  AOI21_X1 U13833 ( .B1(n10777), .B2(P2_EBX_REG_11__SCAN_IN), .A(n10718), .ZN(
        n10719) );
  NAND2_X1 U13834 ( .A1(n10720), .A2(n10719), .ZN(n15102) );
  NAND2_X1 U13835 ( .A1(n15103), .A2(n15102), .ZN(n15095) );
  INV_X1 U13836 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n10722) );
  AOI22_X1 U13837 ( .A1(n10680), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n10721) );
  OAI21_X1 U13838 ( .B1(n10784), .B2(n10722), .A(n10721), .ZN(n10723) );
  AOI21_X1 U13839 ( .B1(n10780), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n10723), .ZN(n15096) );
  AOI22_X1 U13840 ( .A1(n10680), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n10724) );
  OAI21_X1 U13841 ( .B1(n10784), .B2(n10725), .A(n10724), .ZN(n10726) );
  AOI21_X1 U13842 ( .B1(n10780), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n10726), .ZN(n14856) );
  AOI22_X1 U13843 ( .A1(n10680), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n10728) );
  OAI21_X1 U13844 ( .B1(n10784), .B2(n10729), .A(n10728), .ZN(n10730) );
  AOI21_X1 U13845 ( .B1(n10780), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n10730), .ZN(n15080) );
  INV_X1 U13846 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16505) );
  OR2_X1 U13847 ( .A1(n10774), .A2(n16505), .ZN(n10734) );
  INV_X1 U13848 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n10731) );
  OAI22_X1 U13849 ( .A1(n10775), .A2(n10731), .B1(n10677), .B2(n19249), .ZN(
        n10732) );
  AOI21_X1 U13850 ( .B1(n10777), .B2(P2_EBX_REG_15__SCAN_IN), .A(n10732), .ZN(
        n10733) );
  NAND2_X1 U13851 ( .A1(n10734), .A2(n10733), .ZN(n15074) );
  INV_X1 U13852 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15577) );
  OR2_X1 U13853 ( .A1(n10774), .A2(n15577), .ZN(n10737) );
  INV_X1 U13854 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n15584) );
  OAI22_X1 U13855 ( .A1(n10775), .A2(n15584), .B1(n10677), .B2(n10162), .ZN(
        n10735) );
  AOI21_X1 U13856 ( .B1(n10777), .B2(P2_EBX_REG_16__SCAN_IN), .A(n10735), .ZN(
        n10736) );
  NAND2_X1 U13857 ( .A1(n10737), .A2(n10736), .ZN(n15067) );
  AOI22_X1 U13858 ( .A1(n10680), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n10738) );
  OAI21_X1 U13859 ( .B1(n10784), .B2(n10588), .A(n10738), .ZN(n10739) );
  AOI21_X1 U13860 ( .B1(n10780), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n10739), .ZN(n15059) );
  AOI22_X1 U13861 ( .A1(n10680), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n10740) );
  OAI21_X1 U13862 ( .B1(n10784), .B2(n19208), .A(n10740), .ZN(n10741) );
  AOI21_X1 U13863 ( .B1(n10780), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n10741), .ZN(n15051) );
  INV_X1 U13864 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12641) );
  OR2_X1 U13865 ( .A1(n10774), .A2(n12641), .ZN(n10744) );
  INV_X1 U13866 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n15357) );
  OAI22_X1 U13867 ( .A1(n10775), .A2(n15357), .B1(n10677), .B2(n19197), .ZN(
        n10742) );
  AOI21_X1 U13868 ( .B1(n10777), .B2(P2_EBX_REG_19__SCAN_IN), .A(n10742), .ZN(
        n10743) );
  NAND2_X1 U13869 ( .A1(n10744), .A2(n10743), .ZN(n15044) );
  INV_X1 U13870 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15346) );
  OR2_X1 U13871 ( .A1(n10774), .A2(n15346), .ZN(n10748) );
  INV_X1 U13872 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n20020) );
  INV_X1 U13873 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10745) );
  OAI22_X1 U13874 ( .A1(n10775), .A2(n20020), .B1(n10677), .B2(n10745), .ZN(
        n10746) );
  AOI21_X1 U13875 ( .B1(n10777), .B2(P2_EBX_REG_20__SCAN_IN), .A(n10746), .ZN(
        n10747) );
  NAND2_X1 U13876 ( .A1(n10748), .A2(n10747), .ZN(n15036) );
  INV_X1 U13877 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12634) );
  OR2_X1 U13878 ( .A1(n10774), .A2(n12634), .ZN(n10751) );
  INV_X1 U13879 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20022) );
  OAI22_X1 U13880 ( .A1(n10775), .A2(n20022), .B1(n10677), .B2(n14840), .ZN(
        n10749) );
  AOI21_X1 U13881 ( .B1(n10777), .B2(P2_EBX_REG_21__SCAN_IN), .A(n10749), .ZN(
        n10750) );
  INV_X1 U13882 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15515) );
  OR2_X1 U13883 ( .A1(n10774), .A2(n15515), .ZN(n10755) );
  INV_X1 U13884 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n20024) );
  OAI22_X1 U13885 ( .A1(n10775), .A2(n20024), .B1(n10677), .B2(n10752), .ZN(
        n10753) );
  AOI21_X1 U13886 ( .B1(n10777), .B2(P2_EBX_REG_22__SCAN_IN), .A(n10753), .ZN(
        n10754) );
  INV_X1 U13887 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15507) );
  OR2_X1 U13888 ( .A1(n10774), .A2(n15507), .ZN(n10758) );
  INV_X1 U13889 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20026) );
  OAI22_X1 U13890 ( .A1(n10775), .A2(n20026), .B1(n10677), .B2(n14829), .ZN(
        n10756) );
  AOI21_X1 U13891 ( .B1(n10777), .B2(P2_EBX_REG_23__SCAN_IN), .A(n10756), .ZN(
        n10757) );
  NAND2_X1 U13892 ( .A1(n10758), .A2(n10757), .ZN(n14824) );
  OR2_X1 U13893 ( .A1(n10774), .A2(n10218), .ZN(n10762) );
  INV_X1 U13894 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20028) );
  INV_X1 U13895 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10759) );
  OAI22_X1 U13896 ( .A1(n10775), .A2(n20028), .B1(n10677), .B2(n10759), .ZN(
        n10760) );
  AOI21_X1 U13897 ( .B1(n10777), .B2(P2_EBX_REG_24__SCAN_IN), .A(n10760), .ZN(
        n10761) );
  NAND2_X1 U13898 ( .A1(n10762), .A2(n10761), .ZN(n15008) );
  INV_X1 U13899 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15480) );
  OR2_X1 U13900 ( .A1(n10774), .A2(n15480), .ZN(n10765) );
  INV_X1 U13901 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20030) );
  OAI22_X1 U13902 ( .A1(n10775), .A2(n20030), .B1(n10677), .B2(n15295), .ZN(
        n10763) );
  AOI21_X1 U13903 ( .B1(n10777), .B2(P2_EBX_REG_25__SCAN_IN), .A(n10763), .ZN(
        n10764) );
  AOI22_X1 U13904 ( .A1(n10680), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n10766) );
  OAI21_X1 U13905 ( .B1(n10784), .B2(n10116), .A(n10766), .ZN(n10767) );
  AOI21_X1 U13906 ( .B1(n10780), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n10767), .ZN(n14990) );
  INV_X1 U13907 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15453) );
  OR2_X1 U13908 ( .A1(n10774), .A2(n15453), .ZN(n10770) );
  INV_X1 U13909 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n10986) );
  OAI22_X1 U13910 ( .A1(n10775), .A2(n10986), .B1(n10677), .B2(n15273), .ZN(
        n10768) );
  AOI21_X1 U13911 ( .B1(n10777), .B2(P2_EBX_REG_27__SCAN_IN), .A(n10768), .ZN(
        n10769) );
  NAND2_X1 U13912 ( .A1(n10770), .A2(n10769), .ZN(n14982) );
  AOI22_X1 U13913 ( .A1(n10680), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n10771) );
  OAI21_X1 U13914 ( .B1(n10784), .B2(n10772), .A(n10771), .ZN(n10773) );
  AOI21_X1 U13915 ( .B1(n10780), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n10773), .ZN(n14976) );
  INV_X1 U13916 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14092) );
  OR2_X1 U13917 ( .A1(n10774), .A2(n14092), .ZN(n10779) );
  INV_X1 U13918 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n20040) );
  OAI22_X1 U13919 ( .A1(n10775), .A2(n20040), .B1(n10677), .B2(n10158), .ZN(
        n10776) );
  AOI21_X1 U13920 ( .B1(n10777), .B2(P2_EBX_REG_30__SCAN_IN), .A(n10776), .ZN(
        n10778) );
  NAND2_X1 U13921 ( .A1(n10779), .A2(n10778), .ZN(n12414) );
  NAND2_X1 U13922 ( .A1(n10780), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10782) );
  AOI22_X1 U13923 ( .A1(n10680), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n10781) );
  OAI211_X1 U13924 ( .C1(n10784), .C2(n10783), .A(n10782), .B(n10781), .ZN(
        n10785) );
  XNOR2_X1 U13925 ( .A(n10786), .B(n10785), .ZN(n14964) );
  INV_X1 U13926 ( .A(n14964), .ZN(n11002) );
  NOR2_X1 U13927 ( .A1(n12765), .A2(n10787), .ZN(n10788) );
  NAND2_X1 U13928 ( .A1(n10995), .A2(P2_EAX_REG_20__SCAN_IN), .ZN(n10790) );
  NOR2_X2 U13929 ( .A1(n15751), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10824) );
  NAND2_X1 U13930 ( .A1(n10824), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10789) );
  OAI211_X1 U13931 ( .C1(n10989), .C2(n20020), .A(n10790), .B(n10789), .ZN(
        n15190) );
  INV_X2 U13932 ( .A(n9721), .ZN(n10995) );
  AOI22_X1 U13933 ( .A1(n10995), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n10824), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10803) );
  NAND2_X1 U13934 ( .A1(n10998), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n10802) );
  AOI22_X1 U13935 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12088), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10794) );
  AOI22_X1 U13936 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12087), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10793) );
  AOI22_X1 U13937 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10811), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10792) );
  AOI22_X1 U13938 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12152), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10791) );
  NAND4_X1 U13939 ( .A1(n10794), .A2(n10793), .A3(n10792), .A4(n10791), .ZN(
        n10800) );
  AOI22_X1 U13940 ( .A1(n12158), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12157), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10798) );
  AOI22_X1 U13941 ( .A1(n10501), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10797) );
  AOI22_X1 U13942 ( .A1(n10558), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10796) );
  AOI22_X1 U13943 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10795) );
  NAND4_X1 U13944 ( .A1(n10798), .A2(n10797), .A3(n10796), .A4(n10795), .ZN(
        n10799) );
  NAND2_X1 U13945 ( .A1(n10959), .A2(n15101), .ZN(n10801) );
  INV_X1 U13946 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n16585) );
  NAND2_X1 U13947 ( .A1(n12413), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n10804) );
  OAI211_X1 U13948 ( .C1(n15751), .C2(n16585), .A(n10804), .B(n20089), .ZN(
        n10805) );
  AOI21_X1 U13949 ( .B1(n10998), .B2(P2_REIP_REG_0__SCAN_IN), .A(n10805), .ZN(
        n13497) );
  INV_X1 U13950 ( .A(n13497), .ZN(n10823) );
  AOI22_X1 U13951 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10810) );
  AOI22_X1 U13952 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12152), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10809) );
  AOI22_X1 U13953 ( .A1(n12157), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10806), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10808) );
  AOI22_X1 U13954 ( .A1(n12158), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10558), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10807) );
  NAND4_X1 U13955 ( .A1(n10810), .A2(n10809), .A3(n10808), .A4(n10807), .ZN(
        n10817) );
  AOI22_X1 U13956 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10815) );
  AOI22_X1 U13957 ( .A1(n10501), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10544), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10814) );
  AOI22_X1 U13958 ( .A1(n12088), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12087), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10813) );
  AOI22_X1 U13959 ( .A1(n10811), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10812) );
  NAND4_X1 U13960 ( .A1(n10815), .A2(n10814), .A3(n10813), .A4(n10812), .ZN(
        n10816) );
  NOR2_X1 U13961 ( .A1(n10817), .A2(n10816), .ZN(n12816) );
  INV_X1 U13963 ( .A(n10818), .ZN(n10822) );
  INV_X1 U13964 ( .A(n10819), .ZN(n12352) );
  NAND2_X1 U13965 ( .A1(n10824), .A2(n12352), .ZN(n10835) );
  OAI211_X1 U13966 ( .C1(n20089), .C2(n20096), .A(n10835), .B(n9721), .ZN(
        n10820) );
  INV_X1 U13967 ( .A(n10820), .ZN(n10821) );
  NAND2_X1 U13968 ( .A1(n10823), .A2(n13496), .ZN(n10832) );
  AOI22_X1 U13969 ( .A1(n10995), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n10994), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10826) );
  NAND2_X1 U13970 ( .A1(n10998), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10825) );
  AND2_X1 U13971 ( .A1(n10826), .A2(n10825), .ZN(n10833) );
  INV_X1 U13972 ( .A(n10833), .ZN(n10827) );
  XNOR2_X1 U13973 ( .A(n10832), .B(n10827), .ZN(n13054) );
  NAND2_X1 U13974 ( .A1(n10819), .A2(n19486), .ZN(n10828) );
  MUX2_X1 U13975 ( .A(n10828), .B(n20088), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n10830) );
  NAND2_X1 U13976 ( .A1(n10959), .A2(n12815), .ZN(n10829) );
  NAND2_X1 U13977 ( .A1(n10830), .A2(n10829), .ZN(n13055) );
  INV_X1 U13978 ( .A(n13055), .ZN(n10831) );
  NAND2_X1 U13979 ( .A1(n13054), .A2(n10831), .ZN(n13053) );
  NAND2_X1 U13980 ( .A1(n10833), .A2(n10832), .ZN(n10834) );
  NAND2_X1 U13981 ( .A1(n13053), .A2(n10834), .ZN(n10840) );
  NAND2_X1 U13982 ( .A1(n10959), .A2(n12460), .ZN(n10836) );
  OAI211_X1 U13983 ( .C1(n20089), .C2(n20079), .A(n10836), .B(n10835), .ZN(
        n10839) );
  XNOR2_X1 U13984 ( .A(n10840), .B(n10839), .ZN(n13034) );
  AOI22_X1 U13985 ( .A1(n10995), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n10994), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10838) );
  NAND2_X1 U13986 ( .A1(n10998), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10837) );
  AND2_X1 U13987 ( .A1(n10838), .A2(n10837), .ZN(n13033) );
  INV_X1 U13988 ( .A(n10839), .ZN(n10841) );
  NAND2_X1 U13989 ( .A1(n10841), .A2(n10840), .ZN(n10842) );
  NAND2_X1 U13990 ( .A1(n10959), .A2(n12490), .ZN(n10845) );
  NOR2_X1 U13991 ( .A1(n10331), .A2(n20089), .ZN(n10843) );
  AOI21_X1 U13992 ( .B1(n10994), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n10843), .ZN(n10844) );
  NAND2_X1 U13993 ( .A1(n10845), .A2(n10844), .ZN(n10848) );
  NAND2_X1 U13994 ( .A1(n10995), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n10846) );
  OAI21_X1 U13995 ( .B1(n10989), .B2(n10684), .A(n10846), .ZN(n10847) );
  NOR2_X1 U13996 ( .A1(n10848), .A2(n10847), .ZN(n13492) );
  AOI22_X1 U13997 ( .A1(n10998), .A2(P2_REIP_REG_4__SCAN_IN), .B1(n10995), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n10850) );
  AOI22_X1 U13998 ( .A1(n10959), .A2(n12827), .B1(n10994), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10849) );
  NAND2_X1 U13999 ( .A1(n10850), .A2(n10849), .ZN(n13499) );
  INV_X1 U14000 ( .A(n13503), .ZN(n10855) );
  NAND2_X1 U14001 ( .A1(n10995), .A2(P2_EAX_REG_5__SCAN_IN), .ZN(n10852) );
  NAND2_X1 U14002 ( .A1(n10994), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10851) );
  AND2_X1 U14003 ( .A1(n10852), .A2(n10851), .ZN(n10854) );
  NAND2_X1 U14004 ( .A1(n10959), .A2(n12552), .ZN(n10853) );
  OAI211_X1 U14005 ( .C1(n15426), .C2(n10989), .A(n10854), .B(n10853), .ZN(
        n13501) );
  NAND2_X1 U14006 ( .A1(n10855), .A2(n13501), .ZN(n13505) );
  INV_X1 U14007 ( .A(n12589), .ZN(n10856) );
  NAND2_X1 U14008 ( .A1(n10959), .A2(n10856), .ZN(n10857) );
  NAND2_X1 U14009 ( .A1(n10824), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10859) );
  NAND2_X1 U14010 ( .A1(n10995), .A2(P2_EAX_REG_6__SCAN_IN), .ZN(n10858) );
  OAI211_X1 U14011 ( .C1(n10989), .C2(n10860), .A(n10859), .B(n10858), .ZN(
        n13048) );
  INV_X1 U14012 ( .A(n10861), .ZN(n12495) );
  AND2_X1 U14013 ( .A1(n10959), .A2(n12843), .ZN(n10862) );
  NOR2_X1 U14014 ( .A1(n13051), .A2(n10862), .ZN(n13181) );
  AOI222_X1 U14015 ( .A1(n10998), .A2(P2_REIP_REG_7__SCAN_IN), .B1(n10995), 
        .B2(P2_EAX_REG_7__SCAN_IN), .C1(n10994), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n13180) );
  AOI22_X1 U14016 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12088), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10866) );
  AOI22_X1 U14017 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12087), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10865) );
  AOI22_X1 U14018 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12152), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10864) );
  AOI22_X1 U14019 ( .A1(n10811), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10806), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10863) );
  NAND4_X1 U14020 ( .A1(n10866), .A2(n10865), .A3(n10864), .A4(n10863), .ZN(
        n10875) );
  INV_X1 U14021 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n19882) );
  INV_X1 U14022 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n19646) );
  OAI22_X1 U14023 ( .A1(n10868), .A2(n19882), .B1(n10867), .B2(n19646), .ZN(
        n10869) );
  INV_X1 U14024 ( .A(n10869), .ZN(n10873) );
  AOI22_X1 U14025 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10872) );
  AOI22_X1 U14026 ( .A1(n10501), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10871) );
  AOI22_X1 U14027 ( .A1(n10558), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10870) );
  NAND4_X1 U14028 ( .A1(n10873), .A2(n10872), .A3(n10871), .A4(n10870), .ZN(
        n10874) );
  AOI22_X1 U14029 ( .A1(n10998), .A2(P2_REIP_REG_8__SCAN_IN), .B1(n10959), 
        .B2(n13589), .ZN(n10877) );
  AOI22_X1 U14030 ( .A1(n10995), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n10994), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10876) );
  NAND2_X1 U14031 ( .A1(n10877), .A2(n10876), .ZN(n16560) );
  AOI22_X1 U14032 ( .A1(n10995), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n10994), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10890) );
  NAND2_X1 U14033 ( .A1(n10998), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n10889) );
  AOI22_X1 U14034 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12150), .B1(
        n12088), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10881) );
  AOI22_X1 U14035 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12151), .B1(
        n12087), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10880) );
  AOI22_X1 U14036 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10811), .B1(
        n10552), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10879) );
  AOI22_X1 U14037 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n10806), .B1(
        n12152), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10878) );
  NAND4_X1 U14038 ( .A1(n10881), .A2(n10880), .A3(n10879), .A4(n10878), .ZN(
        n10887) );
  AOI22_X1 U14039 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12157), .B1(
        n12158), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10885) );
  AOI22_X1 U14040 ( .A1(n10501), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10884) );
  AOI22_X1 U14041 ( .A1(n10558), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10883) );
  AOI22_X1 U14042 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10544), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10882) );
  NAND4_X1 U14043 ( .A1(n10885), .A2(n10884), .A3(n10883), .A4(n10882), .ZN(
        n10886) );
  NOR2_X1 U14044 ( .A1(n10887), .A2(n10886), .ZN(n13597) );
  NAND2_X1 U14045 ( .A1(n10959), .A2(n12052), .ZN(n10888) );
  NAND2_X1 U14046 ( .A1(n10995), .A2(P2_EAX_REG_10__SCAN_IN), .ZN(n10892) );
  NAND2_X1 U14047 ( .A1(n10824), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10891) );
  AND2_X1 U14048 ( .A1(n10892), .A2(n10891), .ZN(n10904) );
  AOI22_X1 U14049 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12150), .B1(
        n12088), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10896) );
  AOI22_X1 U14050 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n12151), .B1(
        n12087), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10895) );
  AOI22_X1 U14051 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10552), .B1(
        n10806), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10894) );
  AOI22_X1 U14052 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10811), .B1(
        n12152), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10893) );
  NAND4_X1 U14053 ( .A1(n10896), .A2(n10895), .A3(n10894), .A4(n10893), .ZN(
        n10902) );
  AOI22_X1 U14054 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n10558), .B1(
        n12158), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10900) );
  AOI22_X1 U14055 ( .A1(n10501), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10899) );
  AOI22_X1 U14056 ( .A1(n12157), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10898) );
  AOI22_X1 U14057 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10544), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10897) );
  NAND4_X1 U14058 ( .A1(n10900), .A2(n10899), .A3(n10898), .A4(n10897), .ZN(
        n10901) );
  NOR2_X1 U14059 ( .A1(n10902), .A2(n10901), .ZN(n12053) );
  INV_X1 U14060 ( .A(n12053), .ZN(n15111) );
  NAND2_X1 U14061 ( .A1(n10959), .A2(n15111), .ZN(n10903) );
  OAI211_X1 U14062 ( .C1(n10989), .C2(n10905), .A(n10904), .B(n10903), .ZN(
        n13324) );
  NOR2_X2 U14063 ( .A1(n16528), .A2(n16527), .ZN(n16529) );
  INV_X1 U14064 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n10920) );
  NAND2_X1 U14065 ( .A1(n10995), .A2(P2_EAX_REG_12__SCAN_IN), .ZN(n10907) );
  NAND2_X1 U14066 ( .A1(n10824), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10906) );
  AND2_X1 U14067 ( .A1(n10907), .A2(n10906), .ZN(n10919) );
  AOI22_X1 U14068 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12088), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10911) );
  AOI22_X1 U14069 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12087), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10910) );
  AOI22_X1 U14070 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12152), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10909) );
  AOI22_X1 U14071 ( .A1(n10811), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10806), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10908) );
  NAND4_X1 U14072 ( .A1(n10911), .A2(n10910), .A3(n10909), .A4(n10908), .ZN(
        n10917) );
  AOI22_X1 U14073 ( .A1(n12157), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10558), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10915) );
  AOI22_X1 U14074 ( .A1(n10501), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10914) );
  AOI22_X1 U14075 ( .A1(n12158), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10913) );
  AOI22_X1 U14076 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10912) );
  NAND4_X1 U14077 ( .A1(n10915), .A2(n10914), .A3(n10913), .A4(n10912), .ZN(
        n10916) );
  NAND2_X1 U14078 ( .A1(n10959), .A2(n15093), .ZN(n10918) );
  OAI211_X1 U14079 ( .C1(n10989), .C2(n10920), .A(n10919), .B(n10918), .ZN(
        n13451) );
  NAND2_X1 U14080 ( .A1(n16529), .A2(n13451), .ZN(n14859) );
  AOI22_X1 U14081 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12088), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10924) );
  AOI22_X1 U14082 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12087), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10923) );
  INV_X1 U14083 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12111) );
  AOI22_X1 U14084 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10811), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10922) );
  AOI22_X1 U14085 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12152), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10921) );
  NAND4_X1 U14086 ( .A1(n10924), .A2(n10923), .A3(n10922), .A4(n10921), .ZN(
        n10930) );
  AOI22_X1 U14087 ( .A1(n12158), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12157), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10928) );
  AOI22_X1 U14088 ( .A1(n10501), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10927) );
  AOI22_X1 U14089 ( .A1(n10558), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10926) );
  AOI22_X1 U14090 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10925) );
  NAND4_X1 U14091 ( .A1(n10928), .A2(n10927), .A3(n10926), .A4(n10925), .ZN(
        n10929) );
  AOI22_X1 U14092 ( .A1(n10998), .A2(P2_REIP_REG_13__SCAN_IN), .B1(n10959), 
        .B2(n15088), .ZN(n10932) );
  AOI22_X1 U14093 ( .A1(n10995), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n10994), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10931) );
  INV_X1 U14094 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n10947) );
  NAND2_X1 U14095 ( .A1(n10995), .A2(P2_EAX_REG_14__SCAN_IN), .ZN(n10934) );
  NAND2_X1 U14096 ( .A1(n10824), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10933) );
  AND2_X1 U14097 ( .A1(n10934), .A2(n10933), .ZN(n10946) );
  AOI22_X1 U14098 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n12087), .B1(
        n12088), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10938) );
  AOI22_X1 U14099 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n12151), .B1(
        n12150), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10937) );
  AOI22_X1 U14100 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10552), .B1(
        n12152), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10936) );
  AOI22_X1 U14101 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10811), .B1(
        n10806), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10935) );
  NAND4_X1 U14102 ( .A1(n10938), .A2(n10937), .A3(n10936), .A4(n10935), .ZN(
        n10944) );
  AOI22_X1 U14103 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12157), .B1(
        n10558), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10942) );
  AOI22_X1 U14104 ( .A1(n10501), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10941) );
  AOI22_X1 U14105 ( .A1(n12158), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10940) );
  AOI22_X1 U14106 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10544), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10939) );
  NAND4_X1 U14107 ( .A1(n10942), .A2(n10941), .A3(n10940), .A4(n10939), .ZN(
        n10943) );
  NAND2_X1 U14108 ( .A1(n10959), .A2(n15084), .ZN(n10945) );
  OAI211_X1 U14109 ( .C1(n10989), .C2(n10947), .A(n10946), .B(n10945), .ZN(
        n15604) );
  AOI22_X1 U14110 ( .A1(n10995), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n10994), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10962) );
  NAND2_X1 U14111 ( .A1(n10998), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n10961) );
  AOI22_X1 U14112 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n12150), .B1(
        n12088), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10951) );
  AOI22_X1 U14113 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12151), .B1(
        n12087), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10950) );
  AOI22_X1 U14114 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10811), .B1(
        n10552), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10949) );
  AOI22_X1 U14115 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n10806), .B1(
        n12152), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10948) );
  NAND4_X1 U14116 ( .A1(n10951), .A2(n10950), .A3(n10949), .A4(n10948), .ZN(
        n10957) );
  AOI22_X1 U14117 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n12157), .B1(
        n12158), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10955) );
  AOI22_X1 U14118 ( .A1(n10501), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10954) );
  AOI22_X1 U14119 ( .A1(n10558), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10953) );
  AOI22_X1 U14120 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10544), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10952) );
  NAND4_X1 U14121 ( .A1(n10955), .A2(n10954), .A3(n10953), .A4(n10952), .ZN(
        n10956) );
  NOR2_X1 U14122 ( .A1(n10957), .A2(n10956), .ZN(n15073) );
  INV_X1 U14123 ( .A(n15073), .ZN(n10958) );
  NAND2_X1 U14124 ( .A1(n10959), .A2(n10958), .ZN(n10960) );
  NAND2_X1 U14125 ( .A1(n10995), .A2(P2_EAX_REG_16__SCAN_IN), .ZN(n10964) );
  NAND2_X1 U14126 ( .A1(n10824), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10963) );
  OAI211_X1 U14127 ( .C1(n10989), .C2(n15584), .A(n10964), .B(n10963), .ZN(
        n15232) );
  INV_X1 U14128 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n15575) );
  NAND2_X1 U14129 ( .A1(n10995), .A2(P2_EAX_REG_17__SCAN_IN), .ZN(n10966) );
  NAND2_X1 U14130 ( .A1(n10994), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10965) );
  OAI211_X1 U14131 ( .C1(n10989), .C2(n15575), .A(n10966), .B(n10965), .ZN(
        n15222) );
  INV_X1 U14132 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n20017) );
  NAND2_X1 U14133 ( .A1(n10995), .A2(P2_EAX_REG_18__SCAN_IN), .ZN(n10968) );
  NAND2_X1 U14134 ( .A1(n10994), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10967) );
  OAI211_X1 U14135 ( .C1(n10989), .C2(n20017), .A(n10968), .B(n10967), .ZN(
        n15213) );
  AOI22_X1 U14136 ( .A1(n10995), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n10994), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10970) );
  NAND2_X1 U14137 ( .A1(n10998), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n10969) );
  NAND2_X1 U14138 ( .A1(n15190), .A2(n15200), .ZN(n15192) );
  AOI22_X1 U14139 ( .A1(n10995), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n10994), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10972) );
  NAND2_X1 U14140 ( .A1(n10998), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n10971) );
  INV_X1 U14141 ( .A(n14838), .ZN(n10973) );
  AOI22_X1 U14142 ( .A1(n10995), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n10994), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10975) );
  NAND2_X1 U14143 ( .A1(n10998), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n10974) );
  NAND2_X1 U14144 ( .A1(n10995), .A2(P2_EAX_REG_23__SCAN_IN), .ZN(n10977) );
  NAND2_X1 U14145 ( .A1(n10824), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10976) );
  OAI211_X1 U14146 ( .C1(n10989), .C2(n20026), .A(n10977), .B(n10976), .ZN(
        n14827) );
  NAND2_X1 U14147 ( .A1(n10995), .A2(P2_EAX_REG_24__SCAN_IN), .ZN(n10979) );
  NAND2_X1 U14148 ( .A1(n10824), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10978) );
  OAI211_X1 U14149 ( .C1(n10989), .C2(n20028), .A(n10979), .B(n10978), .ZN(
        n15165) );
  NAND2_X1 U14150 ( .A1(n14826), .A2(n15165), .ZN(n15156) );
  AOI22_X1 U14151 ( .A1(n10995), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n10994), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n10981) );
  NAND2_X1 U14152 ( .A1(n10998), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n10980) );
  AOI22_X1 U14153 ( .A1(n10995), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n10994), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10983) );
  NAND2_X1 U14154 ( .A1(n10998), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n10982) );
  NAND2_X1 U14155 ( .A1(n10995), .A2(P2_EAX_REG_27__SCAN_IN), .ZN(n10985) );
  NAND2_X1 U14156 ( .A1(n10824), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10984) );
  OAI211_X1 U14157 ( .C1(n10989), .C2(n10986), .A(n10985), .B(n10984), .ZN(
        n15139) );
  INV_X1 U14158 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n20036) );
  NAND2_X1 U14159 ( .A1(n10995), .A2(P2_EAX_REG_28__SCAN_IN), .ZN(n10988) );
  NAND2_X1 U14160 ( .A1(n10824), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10987) );
  OAI211_X1 U14161 ( .C1(n10989), .C2(n20036), .A(n10988), .B(n10987), .ZN(
        n15129) );
  AOI22_X1 U14162 ( .A1(n10995), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n10994), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n10991) );
  NAND2_X1 U14163 ( .A1(n10998), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n10990) );
  AND2_X1 U14164 ( .A1(n10991), .A2(n10990), .ZN(n15123) );
  INV_X1 U14165 ( .A(n15123), .ZN(n10992) );
  NAND2_X1 U14166 ( .A1(n10993), .A2(n10992), .ZN(n15121) );
  AOI22_X1 U14167 ( .A1(n10995), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n10994), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10997) );
  NAND2_X1 U14168 ( .A1(n10998), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n10996) );
  AND2_X1 U14169 ( .A1(n10997), .A2(n10996), .ZN(n12366) );
  AOI222_X1 U14170 ( .A1(n10998), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n10995), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n10824), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10999) );
  XNOR2_X1 U14171 ( .A(n11000), .B(n10999), .ZN(n15117) );
  INV_X1 U14172 ( .A(n15117), .ZN(n11001) );
  OAI22_X1 U14173 ( .A1(n11002), .A2(n19321), .B1(n11001), .B2(n19320), .ZN(
        n11003) );
  AOI22_X1 U14174 ( .A1(n11050), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11073), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11013) );
  INV_X1 U14175 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11008) );
  AOI22_X1 U14177 ( .A1(n11072), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11055), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11012) );
  NOR2_X4 U14178 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11015) );
  AOI22_X1 U14179 ( .A1(n11586), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11010) );
  AND2_X2 U14180 ( .A1(n11014), .A2(n13330), .ZN(n11215) );
  NOR2_X4 U14181 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13346) );
  AOI22_X1 U14182 ( .A1(n11215), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9683), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11019) );
  AOI22_X1 U14183 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9679), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11018) );
  AOI22_X1 U14184 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11198), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11017) );
  AOI22_X1 U14185 ( .A1(n11078), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11197), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11016) );
  AOI22_X1 U14186 ( .A1(n11198), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9677), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11023) );
  AOI22_X1 U14187 ( .A1(n9668), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11073), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11022) );
  AOI22_X1 U14188 ( .A1(n11078), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11226), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11021) );
  AOI22_X1 U14189 ( .A1(n11072), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9672), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11020) );
  AOI22_X1 U14190 ( .A1(n11112), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11055), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11027) );
  AOI22_X1 U14191 ( .A1(n11215), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11026) );
  AOI22_X1 U14192 ( .A1(n11050), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11025) );
  AOI22_X1 U14193 ( .A1(n9680), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11197), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11024) );
  NAND2_X1 U14194 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11033) );
  NAND2_X1 U14195 ( .A1(n11050), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11032) );
  NAND2_X1 U14196 ( .A1(n11072), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11031) );
  NAND2_X1 U14197 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11030) );
  NAND2_X1 U14198 ( .A1(n11055), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11036) );
  NAND2_X1 U14199 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11035) );
  NAND2_X1 U14200 ( .A1(n11112), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11034) );
  NAND2_X1 U14201 ( .A1(n11197), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11040) );
  NAND2_X1 U14202 ( .A1(n11117), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11039) );
  NAND2_X1 U14203 ( .A1(n11078), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11038) );
  NAND3_X1 U14204 ( .A1(n11040), .A2(n11039), .A3(n11038), .ZN(n11041) );
  NOR2_X1 U14205 ( .A1(n11042), .A2(n11041), .ZN(n11048) );
  NAND2_X1 U14206 ( .A1(n11215), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11046) );
  NAND2_X1 U14207 ( .A1(n11670), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11045) );
  NAND2_X1 U14208 ( .A1(n9648), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11044) );
  NAND2_X1 U14209 ( .A1(n11690), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11043) );
  NAND3_X2 U14210 ( .A1(n11049), .A2(n11048), .A3(n11047), .ZN(n11138) );
  AOI22_X1 U14211 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11117), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11054) );
  AOI22_X1 U14212 ( .A1(n11078), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11197), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11052) );
  AOI22_X1 U14213 ( .A1(n11670), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11198), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11051) );
  NAND4_X1 U14214 ( .A1(n11054), .A2(n11053), .A3(n11052), .A4(n11051), .ZN(
        n11062) );
  AOI22_X1 U14215 ( .A1(n11586), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11058) );
  AOI22_X1 U14216 ( .A1(n11215), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11057) );
  NAND4_X1 U14217 ( .A1(n11060), .A2(n11059), .A3(n11058), .A4(n11057), .ZN(
        n11061) );
  OAI21_X1 U14218 ( .B1(n11130), .B2(n11138), .A(n11152), .ZN(n13073) );
  INV_X1 U14219 ( .A(n13073), .ZN(n11086) );
  AOI22_X1 U14220 ( .A1(n11050), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11072), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11066) );
  BUF_X4 U14221 ( .A(n11078), .Z(n11777) );
  AOI22_X1 U14222 ( .A1(n11777), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11226), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11065) );
  AOI22_X1 U14223 ( .A1(n11586), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9669), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11064) );
  AOI22_X1 U14224 ( .A1(n11215), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9678), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11063) );
  AOI22_X1 U14225 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11112), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11070) );
  AOI22_X1 U14226 ( .A1(n11055), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11069) );
  AOI22_X1 U14227 ( .A1(n11117), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11197), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11068) );
  AOI22_X1 U14228 ( .A1(n11670), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11198), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11067) );
  AOI22_X1 U14229 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11805), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11077) );
  AOI22_X1 U14230 ( .A1(n11072), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11055), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11076) );
  AOI22_X1 U14231 ( .A1(n11050), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9669), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11075) );
  AOI22_X1 U14232 ( .A1(n11586), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11074) );
  NAND4_X1 U14233 ( .A1(n11077), .A2(n11076), .A3(n11075), .A4(n11074), .ZN(
        n11084) );
  AOI22_X1 U14234 ( .A1(n11215), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9683), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11082) );
  AOI22_X1 U14235 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11117), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11081) );
  BUF_X4 U14236 ( .A(n11078), .Z(n11807) );
  AOI22_X1 U14237 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11197), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11080) );
  AOI22_X1 U14238 ( .A1(n9647), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11198), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11079) );
  NAND4_X1 U14239 ( .A1(n11082), .A2(n11081), .A3(n11080), .A4(n11079), .ZN(
        n11083) );
  NAND2_X1 U14240 ( .A1(n13616), .A2(n11828), .ZN(n12972) );
  NAND2_X1 U14241 ( .A1(n11086), .A2(n11085), .ZN(n11925) );
  NOR2_X1 U14242 ( .A1(n11925), .A2(n11136), .ZN(n13078) );
  NAND2_X1 U14243 ( .A1(n11805), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11090) );
  NAND2_X1 U14244 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11089) );
  NAND2_X1 U14245 ( .A1(n11072), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11088) );
  NAND2_X1 U14246 ( .A1(n11055), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11087) );
  NAND2_X1 U14247 ( .A1(n11050), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11095) );
  NAND2_X1 U14248 ( .A1(n11586), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11094) );
  NAND2_X1 U14249 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11093) );
  NAND2_X1 U14250 ( .A1(n11690), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11092) );
  NAND2_X1 U14251 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11099) );
  NAND2_X1 U14252 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11098) );
  NAND2_X1 U14253 ( .A1(n11117), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11097) );
  NAND2_X1 U14254 ( .A1(n11197), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11096) );
  NAND2_X1 U14255 ( .A1(n11215), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11103) );
  NAND2_X1 U14256 ( .A1(n11670), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11102) );
  NAND2_X1 U14257 ( .A1(n9682), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11101) );
  NAND2_X1 U14258 ( .A1(n9647), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11100) );
  NAND4_X4 U14259 ( .A1(n11107), .A2(n11106), .A3(n11105), .A4(n11104), .ZN(
        n13660) );
  NAND2_X1 U14260 ( .A1(n13078), .A2(n13660), .ZN(n12373) );
  NAND2_X1 U14261 ( .A1(n11050), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11111) );
  NAND2_X1 U14262 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11110) );
  NAND2_X1 U14263 ( .A1(n11055), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11109) );
  NAND2_X1 U14264 ( .A1(n9647), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11108) );
  NAND2_X1 U14265 ( .A1(n11072), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11116) );
  NAND2_X1 U14266 ( .A1(n11805), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11115) );
  NAND2_X1 U14267 ( .A1(n11586), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11114) );
  NAND2_X1 U14268 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11113) );
  NAND2_X1 U14269 ( .A1(n11215), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11121) );
  NAND2_X1 U14270 ( .A1(n11777), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11120) );
  NAND2_X1 U14271 ( .A1(n11117), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11119) );
  NAND2_X1 U14272 ( .A1(n11197), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11118) );
  NAND2_X1 U14273 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11125) );
  NAND2_X1 U14274 ( .A1(n11670), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11124) );
  NAND2_X1 U14275 ( .A1(n9682), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11123) );
  NAND2_X1 U14276 ( .A1(n11690), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11122) );
  INV_X1 U14277 ( .A(n11130), .ZN(n11154) );
  NAND3_X1 U14278 ( .A1(n13616), .A2(n11133), .A3(n11134), .ZN(n11135) );
  NAND2_X1 U14279 ( .A1(n11136), .A2(n11135), .ZN(n11137) );
  AOI21_X2 U14280 ( .B1(n11155), .B2(n11828), .A(n11137), .ZN(n11147) );
  INV_X1 U14281 ( .A(n11138), .ZN(n11153) );
  AND2_X2 U14282 ( .A1(n11147), .A2(n9702), .ZN(n12952) );
  INV_X1 U14283 ( .A(n12377), .ZN(n11139) );
  AOI21_X1 U14284 ( .B1(n11144), .B2(n9666), .A(n11139), .ZN(n13224) );
  INV_X1 U14285 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n11140) );
  XNOR2_X1 U14286 ( .A(n11140), .B(P1_STATE_REG_1__SCAN_IN), .ZN(n12968) );
  NAND3_X1 U14287 ( .A1(n13329), .A2(n11176), .A3(n14432), .ZN(n13080) );
  AOI21_X1 U14288 ( .B1(n11144), .B2(n12968), .A(n13225), .ZN(n11145) );
  NAND2_X1 U14289 ( .A1(n13224), .A2(n11145), .ZN(n11146) );
  INV_X1 U14290 ( .A(n11147), .ZN(n11149) );
  NOR2_X1 U14291 ( .A1(n13071), .A2(n13616), .ZN(n11148) );
  NAND2_X1 U14292 ( .A1(n11141), .A2(n13660), .ZN(n11150) );
  NAND2_X1 U14293 ( .A1(n11152), .A2(n13622), .ZN(n11173) );
  OR2_X1 U14294 ( .A1(n11173), .A2(n11154), .ZN(n13070) );
  AND2_X2 U14295 ( .A1(n11828), .A2(n9665), .ZN(n13129) );
  AND2_X1 U14296 ( .A1(n13071), .A2(n13129), .ZN(n11156) );
  INV_X1 U14297 ( .A(n13329), .ZN(n11157) );
  OAI211_X1 U14298 ( .C1(n13656), .C2(n13622), .A(n13654), .B(n11157), .ZN(
        n11158) );
  INV_X1 U14299 ( .A(n11158), .ZN(n11159) );
  NAND3_X1 U14300 ( .A1(n13076), .A2(n11174), .A3(n11159), .ZN(n11160) );
  NAND2_X1 U14301 ( .A1(n11160), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11161) );
  NAND2_X1 U14302 ( .A1(n11184), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11164) );
  NAND2_X1 U14303 ( .A1(n16336), .A2(n20846), .ZN(n11986) );
  NAND2_X1 U14304 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11186) );
  OAI21_X1 U14305 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n11186), .ZN(n20529) );
  NAND2_X1 U14306 ( .A1(n20751), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11181) );
  OAI21_X1 U14307 ( .B1(n11986), .B2(n20529), .A(n11181), .ZN(n11162) );
  INV_X1 U14308 ( .A(n11162), .ZN(n11163) );
  NAND2_X1 U14309 ( .A1(n11164), .A2(n11163), .ZN(n11167) );
  XNOR2_X2 U14310 ( .A(n11167), .B(n11166), .ZN(n13425) );
  NAND2_X1 U14311 ( .A1(n11184), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11169) );
  INV_X1 U14312 ( .A(n20751), .ZN(n16089) );
  MUX2_X1 U14313 ( .A(n16089), .B(n11986), .S(n20643), .Z(n11168) );
  NAND2_X1 U14314 ( .A1(n11169), .A2(n11168), .ZN(n11210) );
  NAND2_X1 U14315 ( .A1(n13329), .A2(n13689), .ZN(n13232) );
  INV_X1 U14316 ( .A(n16336), .ZN(n14804) );
  NAND2_X1 U14317 ( .A1(n11173), .A2(n20842), .ZN(n11179) );
  INV_X1 U14318 ( .A(n11174), .ZN(n11175) );
  NAND2_X1 U14319 ( .A1(n11175), .A2(n9666), .ZN(n11178) );
  INV_X1 U14320 ( .A(n11828), .ZN(n13422) );
  INV_X1 U14321 ( .A(n13649), .ZN(n12954) );
  AND2_X1 U14322 ( .A1(n12954), .A2(n14166), .ZN(n12995) );
  OAI21_X1 U14323 ( .B1(n11154), .B2(n13422), .A(n12995), .ZN(n11177) );
  NAND4_X1 U14324 ( .A1(n11180), .A2(n11179), .A3(n11178), .A4(n11177), .ZN(
        n11208) );
  INV_X1 U14325 ( .A(n11166), .ZN(n11183) );
  NAND2_X1 U14326 ( .A1(n11181), .A2(n14792), .ZN(n11182) );
  NAND2_X1 U14327 ( .A1(n11183), .A2(n11182), .ZN(n11191) );
  NAND2_X1 U14328 ( .A1(n11184), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11189) );
  INV_X1 U14329 ( .A(n11986), .ZN(n11266) );
  INV_X1 U14330 ( .A(n11186), .ZN(n11185) );
  NAND2_X1 U14331 ( .A1(n11185), .A2(n20532), .ZN(n20562) );
  NAND2_X1 U14332 ( .A1(n11186), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11187) );
  NAND2_X1 U14333 ( .A1(n20562), .A2(n11187), .ZN(n13786) );
  AOI22_X1 U14334 ( .A1(n11266), .A2(n13786), .B1(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n20751), .ZN(n11188) );
  INV_X1 U14335 ( .A(n11190), .ZN(n11192) );
  AOI22_X1 U14336 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(n9645), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11196) );
  AOI22_X1 U14337 ( .A1(n11782), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11195) );
  AOI22_X1 U14338 ( .A1(n11050), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11194) );
  AOI22_X1 U14339 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11193) );
  NAND4_X1 U14340 ( .A1(n11196), .A2(n11195), .A3(n11194), .A4(n11193), .ZN(
        n11204) );
  AOI22_X1 U14341 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9684), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11202) );
  AOI22_X1 U14342 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11201) );
  AOI22_X1 U14343 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11197), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11200) );
  AOI22_X1 U14344 ( .A1(n9647), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9682), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11199) );
  NAND4_X1 U14345 ( .A1(n11202), .A2(n11201), .A3(n11200), .A4(n11199), .ZN(
        n11203) );
  INV_X1 U14346 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11205) );
  OAI22_X1 U14347 ( .A1(n11269), .A2(n11846), .B1(n11940), .B2(n11205), .ZN(
        n11206) );
  INV_X1 U14348 ( .A(n11208), .ZN(n11209) );
  AOI22_X1 U14349 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11805), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11214) );
  AOI22_X1 U14350 ( .A1(n11072), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11213) );
  AOI22_X1 U14351 ( .A1(n11050), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11212) );
  AOI22_X1 U14352 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11211) );
  NAND4_X1 U14353 ( .A1(n11214), .A2(n11213), .A3(n11212), .A4(n11211), .ZN(
        n11221) );
  AOI22_X1 U14354 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9684), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11219) );
  AOI22_X1 U14355 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11117), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11218) );
  AOI22_X1 U14356 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11197), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11217) );
  AOI22_X1 U14357 ( .A1(n9647), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9682), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11216) );
  NAND4_X1 U14358 ( .A1(n11219), .A2(n11218), .A3(n11217), .A4(n11216), .ZN(
        n11220) );
  NOR2_X1 U14359 ( .A1(n11270), .A2(n11897), .ZN(n11241) );
  AOI22_X1 U14360 ( .A1(n11782), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9672), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11225) );
  AOI22_X1 U14361 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11224) );
  AOI22_X1 U14362 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11117), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11223) );
  AOI22_X1 U14363 ( .A1(n9682), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11222) );
  NAND4_X1 U14364 ( .A1(n11225), .A2(n11224), .A3(n11223), .A4(n11222), .ZN(
        n11233) );
  AOI22_X1 U14365 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11806), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11231) );
  AOI22_X1 U14366 ( .A1(n11805), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11230) );
  AOI22_X1 U14367 ( .A1(n9684), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11197), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11229) );
  AOI22_X1 U14368 ( .A1(n11050), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9647), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11228) );
  NAND4_X1 U14369 ( .A1(n11231), .A2(n11230), .A3(n11229), .A4(n11228), .ZN(
        n11232) );
  MUX2_X1 U14370 ( .A(n11239), .B(n11241), .S(n11844), .Z(n11234) );
  INV_X1 U14371 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11238) );
  OAI211_X1 U14372 ( .C1(n11940), .C2(n11238), .A(n11237), .B(n11236), .ZN(
        n11345) );
  NAND2_X1 U14373 ( .A1(n11974), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11254) );
  INV_X1 U14374 ( .A(n11241), .ZN(n11253) );
  AOI22_X1 U14375 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(n9645), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11245) );
  AOI22_X1 U14376 ( .A1(n11782), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11244) );
  AOI22_X1 U14377 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11243) );
  AOI22_X1 U14378 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9647), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11242) );
  NAND4_X1 U14379 ( .A1(n11245), .A2(n11244), .A3(n11243), .A4(n11242), .ZN(
        n11251) );
  AOI22_X1 U14380 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11249) );
  AOI22_X1 U14381 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11197), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11248) );
  AOI22_X1 U14382 ( .A1(n9684), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(n9682), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11247) );
  AOI22_X1 U14383 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11246) );
  NAND4_X1 U14384 ( .A1(n11249), .A2(n11248), .A3(n11247), .A4(n11246), .ZN(
        n11250) );
  OR2_X1 U14385 ( .A1(n11269), .A2(n11259), .ZN(n11252) );
  INV_X1 U14386 ( .A(n13425), .ZN(n11257) );
  INV_X1 U14387 ( .A(n11255), .ZN(n11256) );
  NAND2_X1 U14388 ( .A1(n20325), .A2(n9663), .ZN(n13651) );
  INV_X1 U14389 ( .A(n13651), .ZN(n11260) );
  NAND2_X1 U14390 ( .A1(n11339), .A2(n11832), .ZN(n11265) );
  INV_X1 U14391 ( .A(n11261), .ZN(n11262) );
  NAND2_X1 U14392 ( .A1(n11184), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11268) );
  NOR3_X1 U14393 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20532), .A3(
        n20602), .ZN(n13478) );
  INV_X1 U14394 ( .A(n13478), .ZN(n13780) );
  NAND3_X1 U14395 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20673) );
  AOI21_X1 U14396 ( .B1(n20528), .B2(n13625), .A(n20742), .ZN(n20468) );
  AOI22_X1 U14397 ( .A1(n11266), .A2(n20468), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20751), .ZN(n11267) );
  XNOR2_X2 U14398 ( .A(n13347), .B(n13470), .ZN(n20467) );
  AOI22_X1 U14399 ( .A1(n9645), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11274) );
  AOI22_X1 U14400 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11782), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11273) );
  AOI22_X1 U14401 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11272) );
  AOI22_X1 U14402 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9682), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11271) );
  NAND4_X1 U14403 ( .A1(n11274), .A2(n11273), .A3(n11272), .A4(n11271), .ZN(
        n11280) );
  AOI22_X1 U14404 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11278) );
  AOI22_X1 U14405 ( .A1(n9684), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11783), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11277) );
  AOI22_X1 U14406 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9647), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11276) );
  AOI22_X1 U14407 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11275) );
  NAND4_X1 U14408 ( .A1(n11278), .A2(n11277), .A3(n11276), .A4(n11275), .ZN(
        n11279) );
  AOI22_X1 U14409 ( .A1(n11962), .A2(n11859), .B1(n11974), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11281) );
  AOI22_X1 U14410 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9645), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11286) );
  AOI22_X1 U14411 ( .A1(n11782), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11285) );
  AOI22_X1 U14412 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11284) );
  AOI22_X1 U14413 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11283) );
  NAND4_X1 U14414 ( .A1(n11286), .A2(n11285), .A3(n11284), .A4(n11283), .ZN(
        n11292) );
  AOI22_X1 U14415 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11800), .B1(
        n9684), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11290) );
  AOI22_X1 U14416 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11806), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11289) );
  AOI22_X1 U14417 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11777), .B1(
        n11783), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11288) );
  AOI22_X1 U14418 ( .A1(n9647), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9682), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11287) );
  NAND4_X1 U14419 ( .A1(n11290), .A2(n11289), .A3(n11288), .A4(n11287), .ZN(
        n11291) );
  AOI22_X1 U14420 ( .A1(n11962), .A2(n11869), .B1(n11974), .B2(
        P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11362) );
  AOI22_X1 U14421 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11782), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11296) );
  AOI22_X1 U14422 ( .A1(n11777), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11784), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11295) );
  AOI22_X1 U14423 ( .A1(n11805), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11294) );
  AOI22_X1 U14424 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9684), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11293) );
  NAND4_X1 U14425 ( .A1(n11296), .A2(n11295), .A3(n11294), .A4(n11293), .ZN(
        n11302) );
  AOI22_X1 U14426 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11300) );
  AOI22_X1 U14427 ( .A1(n11754), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11783), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11299) );
  AOI22_X1 U14428 ( .A1(n9647), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9682), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11298) );
  AOI22_X1 U14429 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11297) );
  NAND4_X1 U14430 ( .A1(n11300), .A2(n11299), .A3(n11298), .A4(n11297), .ZN(
        n11301) );
  NAND2_X1 U14431 ( .A1(n11962), .A2(n11876), .ZN(n11304) );
  NAND2_X1 U14432 ( .A1(n11974), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11303) );
  INV_X1 U14433 ( .A(n11871), .ZN(n11312) );
  INV_X1 U14434 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n11310) );
  NAND2_X1 U14435 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11354) );
  INV_X1 U14436 ( .A(n11368), .ZN(n11308) );
  INV_X1 U14437 ( .A(n11323), .ZN(n11324) );
  OAI21_X1 U14438 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n11308), .A(
        n11324), .ZN(n16203) );
  AOI22_X1 U14439 ( .A1(n13644), .A2(n16203), .B1(n11824), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11309) );
  OAI21_X1 U14440 ( .B1(n11544), .B2(n11310), .A(n11309), .ZN(n11311) );
  AOI22_X1 U14441 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9645), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11316) );
  AOI22_X1 U14442 ( .A1(n11782), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11315) );
  AOI22_X1 U14443 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11314) );
  AOI22_X1 U14444 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9678), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11313) );
  NAND4_X1 U14445 ( .A1(n11316), .A2(n11315), .A3(n11314), .A4(n11313), .ZN(
        n11322) );
  AOI22_X1 U14446 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9684), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11320) );
  AOI22_X1 U14447 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11319) );
  AOI22_X1 U14448 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11783), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11318) );
  AOI22_X1 U14449 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9682), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11317) );
  NAND4_X1 U14450 ( .A1(n11320), .A2(n11319), .A3(n11318), .A4(n11317), .ZN(
        n11321) );
  AOI22_X1 U14451 ( .A1(n11962), .A2(n11885), .B1(n11974), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11378) );
  NAND2_X1 U14452 ( .A1(n11377), .A2(n11378), .ZN(n11875) );
  INV_X1 U14453 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11329) );
  INV_X1 U14454 ( .A(n11384), .ZN(n11327) );
  INV_X1 U14455 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11325) );
  NAND2_X1 U14456 ( .A1(n11325), .A2(n11324), .ZN(n11326) );
  NAND2_X1 U14457 ( .A1(n11327), .A2(n11326), .ZN(n20188) );
  AOI22_X1 U14458 ( .A1(n20188), .A2(n13644), .B1(n11824), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11328) );
  OAI21_X1 U14459 ( .B1(n11544), .B2(n11329), .A(n11328), .ZN(n11330) );
  AOI21_X1 U14460 ( .B1(n11875), .B2(n11495), .A(n11330), .ZN(n13632) );
  NOR2_X1 U14461 ( .A1(n13631), .A2(n13632), .ZN(n11376) );
  NAND2_X1 U14462 ( .A1(n11332), .A2(n11331), .ZN(n11333) );
  NAND2_X1 U14463 ( .A1(n11352), .A2(n11333), .ZN(n11842) );
  INV_X1 U14464 ( .A(n13212), .ZN(n11334) );
  NAND2_X1 U14465 ( .A1(n11334), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11359) );
  XNOR2_X1 U14466 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13742) );
  AOI21_X1 U14467 ( .B1(n13644), .B2(n13742), .A(n11824), .ZN(n11336) );
  NAND2_X1 U14468 ( .A1(n11825), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11335) );
  OAI211_X1 U14469 ( .C1(n11359), .C2(n11005), .A(n11336), .B(n11335), .ZN(
        n11337) );
  INV_X1 U14470 ( .A(n11337), .ZN(n11338) );
  NAND2_X1 U14471 ( .A1(n11824), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11351) );
  NAND2_X1 U14472 ( .A1(n9673), .A2(n11495), .ZN(n11343) );
  INV_X1 U14473 ( .A(n11359), .ZN(n11365) );
  NAND2_X1 U14474 ( .A1(n11365), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11341) );
  AOI22_X1 U14475 ( .A1(n11825), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20753), .ZN(n11340) );
  AND2_X1 U14476 ( .A1(n11341), .A2(n11340), .ZN(n11342) );
  NAND2_X1 U14477 ( .A1(n13781), .A2(n13689), .ZN(n11346) );
  NAND2_X1 U14478 ( .A1(n11346), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13136) );
  AOI22_X1 U14479 ( .A1(n11825), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20753), .ZN(n11348) );
  OAI21_X1 U14480 ( .B1(n11006), .B2(n11359), .A(n11348), .ZN(n11349) );
  AOI21_X1 U14481 ( .B1(n11347), .B2(n11495), .A(n11349), .ZN(n13137) );
  NAND2_X1 U14482 ( .A1(n13137), .A2(n13644), .ZN(n11350) );
  NAND2_X1 U14483 ( .A1(n13138), .A2(n11350), .ZN(n13146) );
  NAND2_X1 U14484 ( .A1(n13397), .A2(n11351), .ZN(n13367) );
  NAND2_X1 U14485 ( .A1(n11352), .A2(n13390), .ZN(n11353) );
  INV_X1 U14486 ( .A(n11354), .ZN(n11356) );
  INV_X1 U14487 ( .A(n11369), .ZN(n11355) );
  OAI21_X1 U14488 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11356), .A(
        n11355), .ZN(n14373) );
  AOI22_X1 U14489 ( .A1(n13644), .A2(n14373), .B1(n11824), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11358) );
  NAND2_X1 U14490 ( .A1(n11825), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11357) );
  OAI211_X1 U14491 ( .C1(n11359), .C2(n13332), .A(n11358), .B(n11357), .ZN(
        n11360) );
  INV_X1 U14492 ( .A(n11360), .ZN(n11361) );
  OAI21_X1 U14493 ( .B1(n13387), .B2(n11529), .A(n11361), .ZN(n13369) );
  INV_X1 U14494 ( .A(n13368), .ZN(n11375) );
  INV_X1 U14495 ( .A(n11362), .ZN(n11363) );
  XNOR2_X1 U14496 ( .A(n11364), .B(n11363), .ZN(n11858) );
  NAND2_X1 U14497 ( .A1(n11365), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11372) );
  INV_X1 U14498 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11366) );
  AOI21_X1 U14499 ( .B1(n11366), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11367) );
  AOI21_X1 U14500 ( .B1(n11825), .B2(P1_EAX_REG_4__SCAN_IN), .A(n11367), .ZN(
        n11371) );
  OAI21_X1 U14501 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n11369), .A(
        n11368), .ZN(n13842) );
  NOR2_X1 U14502 ( .A1(n13842), .A2(n9799), .ZN(n11370) );
  AOI21_X1 U14503 ( .B1(n11372), .B2(n11371), .A(n11370), .ZN(n11373) );
  NAND2_X1 U14504 ( .A1(n11375), .A2(n11374), .ZN(n13630) );
  INV_X1 U14505 ( .A(n13630), .ZN(n13605) );
  AND2_X2 U14506 ( .A1(n11376), .A2(n13605), .ZN(n13633) );
  NAND2_X1 U14507 ( .A1(n11962), .A2(n11897), .ZN(n11382) );
  NAND2_X1 U14508 ( .A1(n11974), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11381) );
  NAND2_X1 U14509 ( .A1(n11382), .A2(n11381), .ZN(n11383) );
  NAND2_X1 U14510 ( .A1(n11883), .A2(n11495), .ZN(n11389) );
  INV_X1 U14511 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n11386) );
  OAI21_X1 U14512 ( .B1(n11384), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n11404), .ZN(n20163) );
  AOI22_X1 U14513 ( .A1(n20163), .A2(n13644), .B1(n11824), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11385) );
  INV_X1 U14514 ( .A(n11387), .ZN(n11388) );
  NAND2_X1 U14515 ( .A1(n11389), .A2(n11388), .ZN(n13747) );
  AOI22_X1 U14516 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11782), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11393) );
  AOI22_X1 U14517 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11392) );
  AOI22_X1 U14518 ( .A1(n9684), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11783), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11391) );
  AOI22_X1 U14519 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9647), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11390) );
  NAND4_X1 U14520 ( .A1(n11393), .A2(n11392), .A3(n11391), .A4(n11390), .ZN(
        n11399) );
  AOI22_X1 U14521 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9645), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11397) );
  AOI22_X1 U14522 ( .A1(n11775), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11396) );
  AOI22_X1 U14523 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11395) );
  AOI22_X1 U14524 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9682), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11394) );
  NAND4_X1 U14525 ( .A1(n11397), .A2(n11396), .A3(n11395), .A4(n11394), .ZN(
        n11398) );
  OAI21_X1 U14526 ( .B1(n11399), .B2(n11398), .A(n11495), .ZN(n11403) );
  INV_X1 U14527 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11400) );
  XNOR2_X1 U14528 ( .A(n11404), .B(n11400), .ZN(n13862) );
  AOI22_X1 U14529 ( .A1(n13862), .A2(n13644), .B1(n11824), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11402) );
  NAND2_X1 U14530 ( .A1(n11825), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11401) );
  XNOR2_X1 U14531 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n11430), .ZN(
        n20150) );
  INV_X1 U14532 ( .A(n20150), .ZN(n11419) );
  AOI22_X1 U14533 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11805), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11408) );
  AOI22_X1 U14534 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11782), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11407) );
  AOI22_X1 U14535 ( .A1(n11754), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9684), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11406) );
  AOI22_X1 U14536 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9647), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11405) );
  NAND4_X1 U14537 ( .A1(n11408), .A2(n11407), .A3(n11406), .A4(n11405), .ZN(
        n11414) );
  AOI22_X1 U14538 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11806), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11412) );
  AOI22_X1 U14539 ( .A1(n11775), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11411) );
  AOI22_X1 U14540 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11410) );
  AOI22_X1 U14541 ( .A1(n11783), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9682), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11409) );
  NAND4_X1 U14542 ( .A1(n11412), .A2(n11411), .A3(n11410), .A4(n11409), .ZN(
        n11413) );
  NOR2_X1 U14543 ( .A1(n11414), .A2(n11413), .ZN(n11417) );
  NAND2_X1 U14544 ( .A1(n11825), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11416) );
  NAND2_X1 U14545 ( .A1(n11824), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11415) );
  OAI211_X1 U14546 ( .C1(n11529), .C2(n11417), .A(n11416), .B(n11415), .ZN(
        n11418) );
  AOI21_X1 U14547 ( .B1(n11419), .B2(n13644), .A(n11418), .ZN(n13853) );
  AOI22_X1 U14548 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11638), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11423) );
  AOI22_X1 U14549 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11422) );
  AOI22_X1 U14550 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11421) );
  AOI22_X1 U14551 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9678), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11420) );
  NAND4_X1 U14552 ( .A1(n11423), .A2(n11422), .A3(n11421), .A4(n11420), .ZN(
        n11429) );
  AOI22_X1 U14553 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11806), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11427) );
  AOI22_X1 U14554 ( .A1(n11805), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11426) );
  AOI22_X1 U14555 ( .A1(n9684), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11783), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11425) );
  AOI22_X1 U14556 ( .A1(n11072), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9682), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11424) );
  NAND4_X1 U14557 ( .A1(n11427), .A2(n11426), .A3(n11425), .A4(n11424), .ZN(
        n11428) );
  NOR2_X1 U14558 ( .A1(n11429), .A2(n11428), .ZN(n11433) );
  XNOR2_X1 U14559 ( .A(n11434), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14634) );
  NAND2_X1 U14560 ( .A1(n14634), .A2(n13644), .ZN(n11432) );
  AOI22_X1 U14561 ( .A1(n11825), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n11824), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11431) );
  OAI211_X1 U14562 ( .C1(n11433), .C2(n11529), .A(n11432), .B(n11431), .ZN(
        n13867) );
  NAND2_X1 U14563 ( .A1(n11825), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n11437) );
  OAI21_X1 U14564 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11435), .A(
        n11467), .ZN(n16193) );
  AOI22_X1 U14565 ( .A1(n13644), .A2(n16193), .B1(n11824), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11436) );
  NAND2_X1 U14566 ( .A1(n11437), .A2(n11436), .ZN(n11438) );
  AOI22_X1 U14567 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11442) );
  AOI22_X1 U14568 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11800), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11441) );
  AOI22_X1 U14569 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11440) );
  AOI22_X1 U14570 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9678), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11439) );
  NAND4_X1 U14571 ( .A1(n11442), .A2(n11441), .A3(n11440), .A4(n11439), .ZN(
        n11448) );
  AOI22_X1 U14572 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11782), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11446) );
  AOI22_X1 U14573 ( .A1(n11805), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11445) );
  AOI22_X1 U14574 ( .A1(n9684), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11783), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11444) );
  AOI22_X1 U14575 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9648), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11443) );
  NAND4_X1 U14576 ( .A1(n11446), .A2(n11445), .A3(n11444), .A4(n11443), .ZN(
        n11447) );
  OR2_X1 U14577 ( .A1(n11448), .A2(n11447), .ZN(n11449) );
  NAND2_X1 U14578 ( .A1(n11495), .A2(n11449), .ZN(n13896) );
  INV_X1 U14579 ( .A(n13896), .ZN(n11450) );
  NAND2_X1 U14580 ( .A1(n11451), .A2(n11450), .ZN(n13893) );
  AOI22_X1 U14581 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11805), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11456) );
  AOI22_X1 U14582 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n11777), .B1(
        n11806), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11455) );
  AOI22_X1 U14583 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11800), .B1(
        n9684), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11454) );
  AOI22_X1 U14584 ( .A1(n11775), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9674), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11453) );
  NAND4_X1 U14585 ( .A1(n11456), .A2(n11455), .A3(n11454), .A4(n11453), .ZN(
        n11462) );
  AOI22_X1 U14586 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n9681), .B1(
        n11782), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11460) );
  AOI22_X1 U14587 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11776), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11459) );
  AOI22_X1 U14588 ( .A1(n11754), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11783), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11458) );
  AOI22_X1 U14589 ( .A1(n9648), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(n9678), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11457) );
  NAND4_X1 U14590 ( .A1(n11460), .A2(n11459), .A3(n11458), .A4(n11457), .ZN(
        n11461) );
  NOR2_X1 U14591 ( .A1(n11462), .A2(n11461), .ZN(n11466) );
  XNOR2_X1 U14592 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n11467), .ZN(
        n16181) );
  INV_X1 U14593 ( .A(n16181), .ZN(n11463) );
  AOI22_X1 U14594 ( .A1(n11824), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n13644), .B2(n11463), .ZN(n11465) );
  NAND2_X1 U14595 ( .A1(n11825), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n11464) );
  OAI211_X1 U14596 ( .C1(n11529), .C2(n11466), .A(n11465), .B(n11464), .ZN(
        n13930) );
  INV_X1 U14597 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14621) );
  XNOR2_X1 U14598 ( .A(n11483), .B(n14621), .ZN(n14620) );
  AOI22_X1 U14599 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9645), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11472) );
  AOI22_X1 U14600 ( .A1(n11072), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11471) );
  AOI22_X1 U14601 ( .A1(n11754), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9684), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11470) );
  AOI22_X1 U14602 ( .A1(n9647), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9682), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11469) );
  NAND4_X1 U14603 ( .A1(n11472), .A2(n11471), .A3(n11470), .A4(n11469), .ZN(
        n11478) );
  AOI22_X1 U14604 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11806), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11476) );
  AOI22_X1 U14605 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11475) );
  AOI22_X1 U14606 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11783), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11474) );
  AOI22_X1 U14607 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11473) );
  NAND4_X1 U14608 ( .A1(n11476), .A2(n11475), .A3(n11474), .A4(n11473), .ZN(
        n11477) );
  NOR2_X1 U14609 ( .A1(n11478), .A2(n11477), .ZN(n11481) );
  NAND2_X1 U14610 ( .A1(n11825), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11480) );
  NAND2_X1 U14611 ( .A1(n11824), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11479) );
  OAI211_X1 U14612 ( .C1(n11529), .C2(n11481), .A(n11480), .B(n11479), .ZN(
        n11482) );
  AOI21_X1 U14613 ( .B1(n14620), .B2(n13644), .A(n11482), .ZN(n14360) );
  XOR2_X1 U14614 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n11498), .Z(
        n16177) );
  AOI22_X1 U14615 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11782), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11487) );
  AOI22_X1 U14616 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11486) );
  AOI22_X1 U14617 ( .A1(n11754), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9684), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11485) );
  AOI22_X1 U14618 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11484) );
  NAND4_X1 U14619 ( .A1(n11487), .A2(n11486), .A3(n11485), .A4(n11484), .ZN(
        n11493) );
  AOI22_X1 U14620 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9645), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11491) );
  AOI22_X1 U14621 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11806), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11490) );
  AOI22_X1 U14622 ( .A1(n11775), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9674), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11489) );
  AOI22_X1 U14623 ( .A1(n11783), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9682), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11488) );
  NAND4_X1 U14624 ( .A1(n11491), .A2(n11490), .A3(n11489), .A4(n11488), .ZN(
        n11492) );
  OR2_X1 U14625 ( .A1(n11493), .A2(n11492), .ZN(n11494) );
  AOI22_X1 U14626 ( .A1(n11495), .A2(n11494), .B1(n11824), .B2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11497) );
  NAND2_X1 U14627 ( .A1(n11825), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11496) );
  OAI211_X1 U14628 ( .C1(n16177), .C2(n9799), .A(n11497), .B(n11496), .ZN(
        n14421) );
  OR2_X1 U14629 ( .A1(n11499), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11500) );
  NAND2_X1 U14630 ( .A1(n11500), .A2(n11542), .ZN(n16164) );
  AOI22_X1 U14631 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11805), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11504) );
  AOI22_X1 U14632 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9684), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11503) );
  AOI22_X1 U14633 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11502) );
  AOI22_X1 U14634 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9682), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11501) );
  NAND4_X1 U14635 ( .A1(n11504), .A2(n11503), .A3(n11502), .A4(n11501), .ZN(
        n11510) );
  AOI22_X1 U14636 ( .A1(n11072), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11508) );
  AOI22_X1 U14637 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11507) );
  AOI22_X1 U14638 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11783), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11506) );
  AOI22_X1 U14639 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9678), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11505) );
  NAND4_X1 U14640 ( .A1(n11508), .A2(n11507), .A3(n11506), .A4(n11505), .ZN(
        n11509) );
  NOR2_X1 U14641 ( .A1(n11510), .A2(n11509), .ZN(n11513) );
  OAI21_X1 U14642 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20841), .A(
        n20753), .ZN(n11512) );
  NAND2_X1 U14643 ( .A1(n11825), .A2(P1_EAX_REG_16__SCAN_IN), .ZN(n11511) );
  OAI211_X1 U14644 ( .C1(n11819), .C2(n11513), .A(n11512), .B(n11511), .ZN(
        n11514) );
  OAI21_X1 U14645 ( .B1(n16164), .B2(n9799), .A(n11514), .ZN(n14410) );
  XNOR2_X1 U14646 ( .A(n11515), .B(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16165) );
  INV_X1 U14647 ( .A(n16165), .ZN(n11531) );
  AOI22_X1 U14648 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11519) );
  AOI22_X1 U14649 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9684), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11518) );
  AOI22_X1 U14650 ( .A1(n11777), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11517) );
  AOI22_X1 U14651 ( .A1(n11782), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9674), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11516) );
  NAND4_X1 U14652 ( .A1(n11519), .A2(n11518), .A3(n11517), .A4(n11516), .ZN(
        n11525) );
  AOI22_X1 U14653 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11805), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11523) );
  AOI22_X1 U14654 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11522) );
  AOI22_X1 U14655 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11783), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11521) );
  AOI22_X1 U14656 ( .A1(n9648), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11520) );
  NAND4_X1 U14657 ( .A1(n11523), .A2(n11522), .A3(n11521), .A4(n11520), .ZN(
        n11524) );
  NOR2_X1 U14658 ( .A1(n11525), .A2(n11524), .ZN(n11528) );
  NAND2_X1 U14659 ( .A1(n11825), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11527) );
  NAND2_X1 U14660 ( .A1(n11824), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11526) );
  OAI211_X1 U14661 ( .C1(n11529), .C2(n11528), .A(n11527), .B(n11526), .ZN(
        n11530) );
  AOI21_X1 U14662 ( .B1(n11531), .B2(n13644), .A(n11530), .ZN(n14418) );
  INV_X1 U14663 ( .A(n14347), .ZN(n11548) );
  AOI22_X1 U14664 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9645), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11535) );
  AOI22_X1 U14665 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11534) );
  AOI22_X1 U14666 ( .A1(n11777), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9684), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11533) );
  AOI22_X1 U14667 ( .A1(n9682), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(n9678), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11532) );
  NAND4_X1 U14668 ( .A1(n11535), .A2(n11534), .A3(n11533), .A4(n11532), .ZN(
        n11541) );
  AOI22_X1 U14669 ( .A1(n11072), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11539) );
  AOI22_X1 U14670 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11538) );
  AOI22_X1 U14671 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11783), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11537) );
  AOI22_X1 U14672 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9674), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11536) );
  NAND4_X1 U14673 ( .A1(n11539), .A2(n11538), .A3(n11537), .A4(n11536), .ZN(
        n11540) );
  OR2_X1 U14674 ( .A1(n11541), .A2(n11540), .ZN(n11546) );
  INV_X1 U14675 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14479) );
  XNOR2_X1 U14676 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n11563), .ZN(
        n14611) );
  AOI22_X1 U14677 ( .A1(n13644), .A2(n14611), .B1(n11824), .B2(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11543) );
  OAI21_X1 U14678 ( .B1(n11544), .B2(n14479), .A(n11543), .ZN(n11545) );
  AOI21_X1 U14679 ( .B1(n11791), .B2(n11546), .A(n11545), .ZN(n14349) );
  NAND2_X1 U14680 ( .A1(n11548), .A2(n11547), .ZN(n14334) );
  AOI22_X1 U14681 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9645), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11552) );
  AOI22_X1 U14682 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11551) );
  AOI22_X1 U14683 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11550) );
  AOI22_X1 U14684 ( .A1(n11783), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11549) );
  NAND4_X1 U14685 ( .A1(n11552), .A2(n11551), .A3(n11550), .A4(n11549), .ZN(
        n11558) );
  AOI22_X1 U14686 ( .A1(n11072), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11556) );
  AOI22_X1 U14687 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9684), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11555) );
  AOI22_X1 U14688 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9674), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11554) );
  AOI22_X1 U14689 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9682), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11553) );
  NAND4_X1 U14690 ( .A1(n11556), .A2(n11555), .A3(n11554), .A4(n11553), .ZN(
        n11557) );
  NOR2_X1 U14691 ( .A1(n11558), .A2(n11557), .ZN(n11562) );
  NAND2_X1 U14692 ( .A1(n20753), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11559) );
  NAND2_X1 U14693 ( .A1(n9799), .A2(n11559), .ZN(n11560) );
  AOI21_X1 U14694 ( .B1(n11825), .B2(P1_EAX_REG_18__SCAN_IN), .A(n11560), .ZN(
        n11561) );
  OAI21_X1 U14695 ( .B1(n11819), .B2(n11562), .A(n11561), .ZN(n11566) );
  OAI21_X1 U14696 ( .B1(n11564), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n11597), .ZN(n14596) );
  OR2_X1 U14697 ( .A1(n14596), .A2(n9799), .ZN(n11565) );
  NAND2_X1 U14698 ( .A1(n11566), .A2(n11565), .ZN(n14335) );
  AOI22_X1 U14699 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9645), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11570) );
  AOI22_X1 U14700 ( .A1(n11072), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11569) );
  AOI22_X1 U14701 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11568) );
  AOI22_X1 U14702 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11783), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11567) );
  NAND4_X1 U14703 ( .A1(n11570), .A2(n11569), .A3(n11568), .A4(n11567), .ZN(
        n11576) );
  AOI22_X1 U14704 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11574) );
  AOI22_X1 U14705 ( .A1(n11777), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9684), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11573) );
  AOI22_X1 U14706 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9678), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11572) );
  AOI22_X1 U14707 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9682), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11571) );
  NAND4_X1 U14708 ( .A1(n11574), .A2(n11573), .A3(n11572), .A4(n11571), .ZN(
        n11575) );
  NOR2_X1 U14709 ( .A1(n11576), .A2(n11575), .ZN(n11579) );
  AOI21_X1 U14710 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14328), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11577) );
  AOI21_X1 U14711 ( .B1(n11825), .B2(P1_EAX_REG_19__SCAN_IN), .A(n11577), .ZN(
        n11578) );
  OAI21_X1 U14712 ( .B1(n11819), .B2(n11579), .A(n11578), .ZN(n11581) );
  XNOR2_X1 U14713 ( .A(n11597), .B(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14587) );
  NAND2_X1 U14714 ( .A1(n14587), .A2(n13644), .ZN(n11580) );
  AOI22_X1 U14715 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11805), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11585) );
  AOI22_X1 U14716 ( .A1(n11777), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11806), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11584) );
  AOI22_X1 U14717 ( .A1(n11782), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9682), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11583) );
  AOI22_X1 U14718 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11800), .B1(
        n11783), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11582) );
  NAND4_X1 U14719 ( .A1(n11585), .A2(n11584), .A3(n11583), .A4(n11582), .ZN(
        n11592) );
  AOI22_X1 U14720 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11590) );
  AOI22_X1 U14721 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11776), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11589) );
  AOI22_X1 U14722 ( .A1(n11754), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9684), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11588) );
  AOI22_X1 U14723 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11587) );
  NAND4_X1 U14724 ( .A1(n11590), .A2(n11589), .A3(n11588), .A4(n11587), .ZN(
        n11591) );
  NOR2_X1 U14725 ( .A1(n11592), .A2(n11591), .ZN(n11596) );
  NAND2_X1 U14726 ( .A1(n20753), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11593) );
  NAND2_X1 U14727 ( .A1(n9799), .A2(n11593), .ZN(n11594) );
  AOI21_X1 U14728 ( .B1(n11825), .B2(P1_EAX_REG_20__SCAN_IN), .A(n11594), .ZN(
        n11595) );
  OAI21_X1 U14729 ( .B1(n11819), .B2(n11596), .A(n11595), .ZN(n11601) );
  OR2_X1 U14730 ( .A1(n11598), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11599) );
  AND2_X1 U14731 ( .A1(n11599), .A2(n11631), .ZN(n14581) );
  NAND2_X1 U14732 ( .A1(n14581), .A2(n13644), .ZN(n11600) );
  NAND2_X1 U14733 ( .A1(n11601), .A2(n11600), .ZN(n14309) );
  AOI22_X1 U14734 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11605) );
  AOI22_X1 U14735 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11782), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U14736 ( .A1(n11777), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11603) );
  AOI22_X1 U14737 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9674), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11602) );
  NAND4_X1 U14738 ( .A1(n11605), .A2(n11604), .A3(n11603), .A4(n11602), .ZN(
        n11611) );
  AOI22_X1 U14739 ( .A1(n9645), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11609) );
  AOI22_X1 U14740 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11783), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11608) );
  AOI22_X1 U14741 ( .A1(n9684), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(n9648), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11607) );
  AOI22_X1 U14742 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9678), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11606) );
  NAND4_X1 U14743 ( .A1(n11609), .A2(n11608), .A3(n11607), .A4(n11606), .ZN(
        n11610) );
  NOR2_X1 U14744 ( .A1(n11611), .A2(n11610), .ZN(n11614) );
  INV_X1 U14745 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14571) );
  AOI21_X1 U14746 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14571), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11612) );
  AOI21_X1 U14747 ( .B1(n11825), .B2(P1_EAX_REG_21__SCAN_IN), .A(n11612), .ZN(
        n11613) );
  OAI21_X1 U14748 ( .B1(n11819), .B2(n11614), .A(n11613), .ZN(n11616) );
  XNOR2_X1 U14749 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n11631), .ZN(
        n14569) );
  NAND2_X1 U14750 ( .A1(n13644), .A2(n14569), .ZN(n11615) );
  NAND2_X1 U14751 ( .A1(n11616), .A2(n11615), .ZN(n14297) );
  AOI22_X1 U14752 ( .A1(n9645), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11620) );
  AOI22_X1 U14753 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11782), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11619) );
  AOI22_X1 U14754 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9684), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11618) );
  AOI22_X1 U14755 ( .A1(n11777), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11617) );
  NAND4_X1 U14756 ( .A1(n11620), .A2(n11619), .A3(n11618), .A4(n11617), .ZN(
        n11626) );
  AOI22_X1 U14757 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11624) );
  AOI22_X1 U14758 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11783), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11623) );
  AOI22_X1 U14759 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9648), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11622) );
  AOI22_X1 U14760 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9678), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11621) );
  NAND4_X1 U14761 ( .A1(n11624), .A2(n11623), .A3(n11622), .A4(n11621), .ZN(
        n11625) );
  NOR2_X1 U14762 ( .A1(n11626), .A2(n11625), .ZN(n11630) );
  NAND2_X1 U14763 ( .A1(n20753), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11627) );
  NAND2_X1 U14764 ( .A1(n9799), .A2(n11627), .ZN(n11628) );
  AOI21_X1 U14765 ( .B1(n11825), .B2(P1_EAX_REG_22__SCAN_IN), .A(n11628), .ZN(
        n11629) );
  OAI21_X1 U14766 ( .B1(n11819), .B2(n11630), .A(n11629), .ZN(n11637) );
  INV_X1 U14767 ( .A(n11633), .ZN(n11634) );
  INV_X1 U14768 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14561) );
  NAND2_X1 U14769 ( .A1(n11634), .A2(n14561), .ZN(n11635) );
  AND2_X1 U14770 ( .A1(n11681), .A2(n11635), .ZN(n14563) );
  NAND2_X1 U14771 ( .A1(n14563), .A2(n13644), .ZN(n11636) );
  NAND2_X1 U14772 ( .A1(n11637), .A2(n11636), .ZN(n14282) );
  AOI22_X1 U14773 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9645), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11642) );
  AOI22_X1 U14774 ( .A1(n11782), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11641) );
  AOI22_X1 U14775 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11640) );
  AOI22_X1 U14776 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11639) );
  NAND4_X1 U14777 ( .A1(n11642), .A2(n11641), .A3(n11640), .A4(n11639), .ZN(
        n11648) );
  AOI22_X1 U14778 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9684), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11646) );
  AOI22_X1 U14779 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11645) );
  AOI22_X1 U14780 ( .A1(n11777), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11783), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11644) );
  AOI22_X1 U14781 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9682), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11643) );
  NAND4_X1 U14782 ( .A1(n11646), .A2(n11645), .A3(n11644), .A4(n11643), .ZN(
        n11647) );
  NOR2_X1 U14783 ( .A1(n11648), .A2(n11647), .ZN(n11665) );
  AOI22_X1 U14784 ( .A1(n11775), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11652) );
  AOI22_X1 U14785 ( .A1(n11754), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11783), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11651) );
  AOI22_X1 U14786 ( .A1(n9684), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(n9647), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11650) );
  AOI22_X1 U14787 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9678), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11649) );
  NAND4_X1 U14788 ( .A1(n11652), .A2(n11651), .A3(n11650), .A4(n11649), .ZN(
        n11658) );
  AOI22_X1 U14789 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9645), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11656) );
  AOI22_X1 U14790 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11782), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11655) );
  AOI22_X1 U14791 ( .A1(n11777), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11806), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11654) );
  AOI22_X1 U14792 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9682), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11653) );
  NAND4_X1 U14793 ( .A1(n11656), .A2(n11655), .A3(n11654), .A4(n11653), .ZN(
        n11657) );
  NOR2_X1 U14794 ( .A1(n11658), .A2(n11657), .ZN(n11664) );
  XOR2_X1 U14795 ( .A(n11665), .B(n11664), .Z(n11659) );
  NAND2_X1 U14796 ( .A1(n11659), .A2(n11791), .ZN(n11663) );
  AOI21_X1 U14797 ( .B1(n14550), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11660) );
  AOI21_X1 U14798 ( .B1(n11825), .B2(P1_EAX_REG_23__SCAN_IN), .A(n11660), .ZN(
        n11662) );
  XNOR2_X1 U14799 ( .A(n11681), .B(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14555) );
  AOI21_X1 U14800 ( .B1(n11663), .B2(n11662), .A(n11661), .ZN(n14270) );
  AND2_X2 U14801 ( .A1(n14268), .A2(n14270), .ZN(n14258) );
  NOR2_X1 U14802 ( .A1(n11665), .A2(n11664), .ZN(n11689) );
  AOI22_X1 U14803 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9645), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11669) );
  AOI22_X1 U14804 ( .A1(n11782), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11668) );
  AOI22_X1 U14805 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11667) );
  AOI22_X1 U14806 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11666) );
  NAND4_X1 U14807 ( .A1(n11669), .A2(n11668), .A3(n11667), .A4(n11666), .ZN(
        n11676) );
  AOI22_X1 U14808 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9684), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11674) );
  AOI22_X1 U14809 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11673) );
  AOI22_X1 U14810 ( .A1(n11777), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11783), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11672) );
  AOI22_X1 U14811 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(n9682), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11671) );
  NAND4_X1 U14812 ( .A1(n11674), .A2(n11673), .A3(n11672), .A4(n11671), .ZN(
        n11675) );
  OR2_X1 U14813 ( .A1(n11676), .A2(n11675), .ZN(n11688) );
  INV_X1 U14814 ( .A(n11688), .ZN(n11677) );
  XNOR2_X1 U14815 ( .A(n11689), .B(n11677), .ZN(n11678) );
  NAND2_X1 U14816 ( .A1(n11678), .A2(n11791), .ZN(n11687) );
  NAND2_X1 U14817 ( .A1(n20753), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11679) );
  NAND2_X1 U14818 ( .A1(n9799), .A2(n11679), .ZN(n11680) );
  AOI21_X1 U14819 ( .B1(n11825), .B2(P1_EAX_REG_24__SCAN_IN), .A(n11680), .ZN(
        n11686) );
  INV_X1 U14820 ( .A(n11682), .ZN(n11683) );
  INV_X1 U14821 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14543) );
  NAND2_X1 U14822 ( .A1(n11683), .A2(n14543), .ZN(n11684) );
  NAND2_X1 U14823 ( .A1(n11723), .A2(n11684), .ZN(n14542) );
  NOR2_X1 U14824 ( .A1(n14542), .A2(n9799), .ZN(n11685) );
  AOI21_X1 U14825 ( .B1(n11687), .B2(n11686), .A(n11685), .ZN(n14260) );
  NAND2_X1 U14826 ( .A1(n11689), .A2(n11688), .ZN(n11708) );
  AOI22_X1 U14827 ( .A1(n11775), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U14828 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11693) );
  AOI22_X1 U14829 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11783), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11692) );
  AOI22_X1 U14830 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11691) );
  NAND4_X1 U14831 ( .A1(n11694), .A2(n11693), .A3(n11692), .A4(n11691), .ZN(
        n11700) );
  AOI22_X1 U14832 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9645), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11698) );
  AOI22_X1 U14833 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11782), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11697) );
  AOI22_X1 U14834 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9684), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11696) );
  AOI22_X1 U14835 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(n9682), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11695) );
  NAND4_X1 U14836 ( .A1(n11698), .A2(n11697), .A3(n11696), .A4(n11695), .ZN(
        n11699) );
  NOR2_X1 U14837 ( .A1(n11700), .A2(n11699), .ZN(n11709) );
  XOR2_X1 U14838 ( .A(n11708), .B(n11709), .Z(n11701) );
  NAND2_X1 U14839 ( .A1(n11701), .A2(n11791), .ZN(n11704) );
  INV_X1 U14840 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14531) );
  AOI21_X1 U14841 ( .B1(n14531), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11702) );
  AOI21_X1 U14842 ( .B1(n11825), .B2(P1_EAX_REG_25__SCAN_IN), .A(n11702), .ZN(
        n11703) );
  NAND2_X1 U14843 ( .A1(n11704), .A2(n11703), .ZN(n11706) );
  XNOR2_X1 U14844 ( .A(n11723), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14533) );
  NAND2_X1 U14845 ( .A1(n14533), .A2(n13644), .ZN(n11705) );
  NAND2_X1 U14846 ( .A1(n11706), .A2(n11705), .ZN(n14246) );
  NOR2_X1 U14847 ( .A1(n11709), .A2(n11708), .ZN(n11731) );
  AOI22_X1 U14848 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9645), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11713) );
  AOI22_X1 U14849 ( .A1(n11782), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11712) );
  AOI22_X1 U14850 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11711) );
  AOI22_X1 U14851 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9677), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11710) );
  NAND4_X1 U14852 ( .A1(n11713), .A2(n11712), .A3(n11711), .A4(n11710), .ZN(
        n11719) );
  AOI22_X1 U14853 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9684), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11717) );
  AOI22_X1 U14854 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11716) );
  AOI22_X1 U14855 ( .A1(n11777), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11783), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11715) );
  AOI22_X1 U14856 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(n9648), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11714) );
  NAND4_X1 U14857 ( .A1(n11717), .A2(n11716), .A3(n11715), .A4(n11714), .ZN(
        n11718) );
  OR2_X1 U14858 ( .A1(n11719), .A2(n11718), .ZN(n11730) );
  XNOR2_X1 U14859 ( .A(n11731), .B(n11730), .ZN(n11722) );
  INV_X1 U14860 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14520) );
  AOI21_X1 U14861 ( .B1(n14520), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11720) );
  AOI21_X1 U14862 ( .B1(n11825), .B2(P1_EAX_REG_26__SCAN_IN), .A(n11720), .ZN(
        n11721) );
  OAI21_X1 U14863 ( .B1(n11722), .B2(n11819), .A(n11721), .ZN(n11729) );
  INV_X1 U14864 ( .A(n11723), .ZN(n11724) );
  INV_X1 U14865 ( .A(n11725), .ZN(n11726) );
  NAND2_X1 U14866 ( .A1(n11726), .A2(n14520), .ZN(n11727) );
  NAND2_X1 U14867 ( .A1(n11765), .A2(n11727), .ZN(n14519) );
  NAND2_X1 U14868 ( .A1(n11729), .A2(n11728), .ZN(n14236) );
  NAND2_X1 U14869 ( .A1(n11731), .A2(n11730), .ZN(n11748) );
  AOI22_X1 U14870 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11782), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11735) );
  AOI22_X1 U14871 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11777), .B1(
        n11806), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11734) );
  AOI22_X1 U14872 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n11776), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11733) );
  AOI22_X1 U14873 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(n9678), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11732) );
  NAND4_X1 U14874 ( .A1(n11735), .A2(n11734), .A3(n11733), .A4(n11732), .ZN(
        n11741) );
  AOI22_X1 U14875 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9645), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11739) );
  AOI22_X1 U14876 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11800), .B1(
        n9684), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11738) );
  AOI22_X1 U14877 ( .A1(n11754), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11783), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11737) );
  AOI22_X1 U14878 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11775), .B1(
        n9648), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11736) );
  NAND4_X1 U14879 ( .A1(n11739), .A2(n11738), .A3(n11737), .A4(n11736), .ZN(
        n11740) );
  NOR2_X1 U14880 ( .A1(n11741), .A2(n11740), .ZN(n11749) );
  XOR2_X1 U14881 ( .A(n11748), .B(n11749), .Z(n11742) );
  NAND2_X1 U14882 ( .A1(n11742), .A2(n11791), .ZN(n11747) );
  NAND2_X1 U14883 ( .A1(n20753), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11743) );
  NAND2_X1 U14884 ( .A1(n9799), .A2(n11743), .ZN(n11744) );
  AOI21_X1 U14885 ( .B1(n11825), .B2(P1_EAX_REG_27__SCAN_IN), .A(n11744), .ZN(
        n11746) );
  XNOR2_X1 U14886 ( .A(n11765), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14226) );
  AOI21_X1 U14887 ( .B1(n11747), .B2(n11746), .A(n11745), .ZN(n12002) );
  NOR2_X1 U14888 ( .A1(n11749), .A2(n11748), .ZN(n11774) );
  AOI22_X1 U14889 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9645), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11753) );
  AOI22_X1 U14890 ( .A1(n11782), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11752) );
  AOI22_X1 U14891 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11751) );
  AOI22_X1 U14892 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9677), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11750) );
  NAND4_X1 U14893 ( .A1(n11753), .A2(n11752), .A3(n11751), .A4(n11750), .ZN(
        n11760) );
  AOI22_X1 U14894 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9684), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11758) );
  AOI22_X1 U14895 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11757) );
  AOI22_X1 U14896 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11783), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11756) );
  AOI22_X1 U14897 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(n9648), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11755) );
  NAND4_X1 U14898 ( .A1(n11758), .A2(n11757), .A3(n11756), .A4(n11755), .ZN(
        n11759) );
  OR2_X1 U14899 ( .A1(n11760), .A2(n11759), .ZN(n11773) );
  INV_X1 U14900 ( .A(n11773), .ZN(n11761) );
  XNOR2_X1 U14901 ( .A(n11774), .B(n11761), .ZN(n11762) );
  NAND2_X1 U14902 ( .A1(n11762), .A2(n11791), .ZN(n11772) );
  NAND2_X1 U14903 ( .A1(n20753), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11763) );
  NAND2_X1 U14904 ( .A1(n9799), .A2(n11763), .ZN(n11764) );
  AOI21_X1 U14905 ( .B1(n11825), .B2(P1_EAX_REG_28__SCAN_IN), .A(n11764), .ZN(
        n11771) );
  INV_X1 U14906 ( .A(n11765), .ZN(n11766) );
  INV_X1 U14907 ( .A(n11767), .ZN(n11768) );
  INV_X1 U14908 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12874) );
  NAND2_X1 U14909 ( .A1(n11768), .A2(n12874), .ZN(n11769) );
  NAND2_X1 U14910 ( .A1(n11821), .A2(n11769), .ZN(n14214) );
  NOR2_X1 U14911 ( .A1(n14214), .A2(n9799), .ZN(n11770) );
  NAND2_X1 U14912 ( .A1(n11774), .A2(n11773), .ZN(n11798) );
  AOI22_X1 U14913 ( .A1(n9645), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11781) );
  AOI22_X1 U14914 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11780) );
  AOI22_X1 U14915 ( .A1(n11777), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11779) );
  AOI22_X1 U14916 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11778) );
  NAND4_X1 U14917 ( .A1(n11781), .A2(n11780), .A3(n11779), .A4(n11778), .ZN(
        n11790) );
  AOI22_X1 U14918 ( .A1(n11782), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11638), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11788) );
  AOI22_X1 U14919 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9684), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11787) );
  AOI22_X1 U14920 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11783), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11786) );
  AOI22_X1 U14921 ( .A1(n9681), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9648), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11785) );
  NAND4_X1 U14922 ( .A1(n11788), .A2(n11787), .A3(n11786), .A4(n11785), .ZN(
        n11789) );
  NOR2_X1 U14923 ( .A1(n11790), .A2(n11789), .ZN(n11799) );
  XOR2_X1 U14924 ( .A(n11798), .B(n11799), .Z(n11792) );
  NAND2_X1 U14925 ( .A1(n11792), .A2(n11791), .ZN(n11795) );
  INV_X1 U14926 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14511) );
  AOI21_X1 U14927 ( .B1(n14511), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11793) );
  AOI21_X1 U14928 ( .B1(n11825), .B2(P1_EAX_REG_29__SCAN_IN), .A(n11793), .ZN(
        n11794) );
  NAND2_X1 U14929 ( .A1(n11795), .A2(n11794), .ZN(n11797) );
  XNOR2_X1 U14930 ( .A(n11821), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14513) );
  NAND2_X1 U14931 ( .A1(n14513), .A2(n13644), .ZN(n11796) );
  NOR2_X1 U14932 ( .A1(n11799), .A2(n11798), .ZN(n11815) );
  AOI22_X1 U14933 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11091), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11804) );
  AOI22_X1 U14934 ( .A1(n9684), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11783), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11803) );
  AOI22_X1 U14935 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9674), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11802) );
  AOI22_X1 U14936 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11801) );
  NAND4_X1 U14937 ( .A1(n11804), .A2(n11803), .A3(n11802), .A4(n11801), .ZN(
        n11813) );
  AOI22_X1 U14938 ( .A1(n9645), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11811) );
  AOI22_X1 U14939 ( .A1(n11050), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11782), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11810) );
  AOI22_X1 U14940 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11809) );
  AOI22_X1 U14941 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9648), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11808) );
  NAND4_X1 U14942 ( .A1(n11811), .A2(n11810), .A3(n11809), .A4(n11808), .ZN(
        n11812) );
  NOR2_X1 U14943 ( .A1(n11813), .A2(n11812), .ZN(n11814) );
  XOR2_X1 U14944 ( .A(n11815), .B(n11814), .Z(n11820) );
  NAND2_X1 U14945 ( .A1(n20753), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11816) );
  NAND2_X1 U14946 ( .A1(n9799), .A2(n11816), .ZN(n11817) );
  AOI21_X1 U14947 ( .B1(n11825), .B2(P1_EAX_REG_30__SCAN_IN), .A(n11817), .ZN(
        n11818) );
  OAI21_X1 U14948 ( .B1(n11820), .B2(n11819), .A(n11818), .ZN(n11823) );
  XNOR2_X1 U14949 ( .A(n11984), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14191) );
  NAND2_X1 U14950 ( .A1(n14191), .A2(n13644), .ZN(n11822) );
  NAND2_X1 U14951 ( .A1(n11823), .A2(n11822), .ZN(n11991) );
  AOI22_X1 U14952 ( .A1(n11825), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n11824), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11826) );
  INV_X1 U14953 ( .A(n11826), .ZN(n11827) );
  NOR2_X1 U14954 ( .A1(n16345), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13643) );
  INV_X1 U14955 ( .A(n11927), .ZN(n11884) );
  NAND2_X1 U14956 ( .A1(n13419), .A2(n11884), .ZN(n11831) );
  OAI21_X1 U14957 ( .B1(n13656), .B2(n11844), .A(n11847), .ZN(n11829) );
  INV_X1 U14958 ( .A(n11829), .ZN(n11830) );
  NAND2_X1 U14959 ( .A1(n11832), .A2(n9666), .ZN(n11836) );
  XNOR2_X1 U14960 ( .A(n11844), .B(n11843), .ZN(n11833) );
  OAI211_X1 U14961 ( .C1(n11833), .C2(n13656), .A(n11085), .B(n11133), .ZN(
        n11834) );
  INV_X1 U14962 ( .A(n11834), .ZN(n11835) );
  NAND2_X1 U14963 ( .A1(n11836), .A2(n11835), .ZN(n11838) );
  INV_X1 U14964 ( .A(n11838), .ZN(n11839) );
  OR2_X1 U14965 ( .A1(n11837), .A2(n11839), .ZN(n11840) );
  INV_X1 U14966 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13293) );
  OR2_X1 U14967 ( .A1(n11842), .A2(n11927), .ZN(n11851) );
  NAND2_X1 U14968 ( .A1(n11844), .A2(n11843), .ZN(n11845) );
  NAND2_X1 U14969 ( .A1(n11845), .A2(n11846), .ZN(n11860) );
  OAI21_X1 U14970 ( .B1(n11846), .B2(n11845), .A(n11860), .ZN(n11849) );
  INV_X1 U14971 ( .A(n11847), .ZN(n11848) );
  AOI21_X1 U14972 ( .B1(n11849), .B2(n20842), .A(n11848), .ZN(n11850) );
  NAND2_X1 U14973 ( .A1(n11851), .A2(n11850), .ZN(n13283) );
  NAND2_X1 U14974 ( .A1(n13284), .A2(n13283), .ZN(n11854) );
  NAND2_X1 U14975 ( .A1(n11852), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11853) );
  NAND2_X1 U14976 ( .A1(n11854), .A2(n11853), .ZN(n13403) );
  XNOR2_X1 U14977 ( .A(n11860), .B(n11859), .ZN(n11855) );
  OAI22_X2 U14978 ( .A1(n13387), .A2(n11927), .B1(n13656), .B2(n11855), .ZN(
        n11856) );
  INV_X1 U14979 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13405) );
  NAND2_X1 U14980 ( .A1(n11856), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11857) );
  NAND2_X1 U14981 ( .A1(n11858), .A2(n11884), .ZN(n11864) );
  AND2_X1 U14982 ( .A1(n11860), .A2(n11859), .ZN(n11868) );
  INV_X1 U14983 ( .A(n11869), .ZN(n11861) );
  XNOR2_X1 U14984 ( .A(n11868), .B(n11861), .ZN(n11862) );
  NAND2_X1 U14985 ( .A1(n11862), .A2(n20842), .ZN(n11863) );
  NAND2_X1 U14986 ( .A1(n11864), .A2(n11863), .ZN(n11866) );
  INV_X1 U14987 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11865) );
  XNOR2_X1 U14988 ( .A(n11866), .B(n11865), .ZN(n13461) );
  NAND2_X1 U14989 ( .A1(n11866), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11867) );
  AND2_X1 U14990 ( .A1(n11869), .A2(n11868), .ZN(n11877) );
  XNOR2_X1 U14991 ( .A(n11876), .B(n11877), .ZN(n11870) );
  OAI22_X1 U14992 ( .A1(n11871), .A2(n11927), .B1(n11870), .B2(n13656), .ZN(
        n11872) );
  INV_X1 U14993 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13636) );
  XNOR2_X1 U14994 ( .A(n11872), .B(n13636), .ZN(n13721) );
  NAND2_X1 U14995 ( .A1(n13722), .A2(n13721), .ZN(n11874) );
  NAND2_X1 U14996 ( .A1(n11872), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11873) );
  NAND2_X1 U14997 ( .A1(n11874), .A2(n11873), .ZN(n13834) );
  NAND3_X1 U14998 ( .A1(n11895), .A2(n11875), .A3(n11884), .ZN(n11880) );
  NAND2_X1 U14999 ( .A1(n11877), .A2(n11876), .ZN(n11886) );
  XNOR2_X1 U15000 ( .A(n11885), .B(n11886), .ZN(n11878) );
  NAND2_X1 U15001 ( .A1(n20842), .A2(n11878), .ZN(n11879) );
  NAND2_X1 U15002 ( .A1(n11880), .A2(n11879), .ZN(n11881) );
  INV_X1 U15003 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16332) );
  XNOR2_X1 U15004 ( .A(n11881), .B(n16332), .ZN(n13835) );
  NAND2_X1 U15005 ( .A1(n11881), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11882) );
  NAND2_X1 U15006 ( .A1(n11883), .A2(n11884), .ZN(n11891) );
  INV_X1 U15007 ( .A(n11885), .ZN(n11887) );
  NOR2_X1 U15008 ( .A1(n11887), .A2(n11886), .ZN(n11896) );
  INV_X1 U15009 ( .A(n11896), .ZN(n11888) );
  XNOR2_X1 U15010 ( .A(n11897), .B(n11888), .ZN(n11889) );
  NAND2_X1 U15011 ( .A1(n20842), .A2(n11889), .ZN(n11890) );
  NAND2_X1 U15012 ( .A1(n11891), .A2(n11890), .ZN(n11892) );
  NAND2_X1 U15013 ( .A1(n11892), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16196) );
  NOR2_X1 U15014 ( .A1(n11893), .A2(n11927), .ZN(n11894) );
  NAND2_X1 U15015 ( .A1(n11897), .A2(n11896), .ZN(n11898) );
  NOR2_X1 U15016 ( .A1(n13656), .A2(n11898), .ZN(n11899) );
  NOR2_X2 U15017 ( .A1(n16174), .A2(n11899), .ZN(n13858) );
  NAND2_X1 U15018 ( .A1(n13858), .A2(n16314), .ZN(n11900) );
  INV_X1 U15019 ( .A(n13858), .ZN(n11901) );
  NAND2_X1 U15020 ( .A1(n11901), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11902) );
  AND2_X1 U15021 ( .A1(n16174), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11903) );
  OR2_X1 U15022 ( .A1(n16174), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11904) );
  AND2_X1 U15023 ( .A1(n16174), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14759) );
  NAND2_X1 U15024 ( .A1(n16174), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11905) );
  NAND2_X1 U15025 ( .A1(n11906), .A2(n11905), .ZN(n14756) );
  INV_X1 U15026 ( .A(n13906), .ZN(n14616) );
  OAI21_X1 U15027 ( .B1(n16174), .B2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n11906), .ZN(n14619) );
  NOR3_X1 U15028 ( .A1(n14617), .A2(n14616), .A3(n14619), .ZN(n16170) );
  OR2_X1 U15029 ( .A1(n16174), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11907) );
  INV_X1 U15030 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14124) );
  XNOR2_X1 U15031 ( .A(n16174), .B(n14124), .ZN(n14761) );
  NOR2_X1 U15032 ( .A1(n16174), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14760) );
  INV_X1 U15033 ( .A(n14760), .ZN(n11908) );
  OAI211_X2 U15034 ( .C1(n11910), .C2(n14757), .A(n14761), .B(n11908), .ZN(
        n14604) );
  INV_X1 U15035 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11909) );
  INV_X1 U15036 ( .A(n11910), .ZN(n14605) );
  NAND2_X1 U15037 ( .A1(n16174), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13907) );
  INV_X1 U15038 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14627) );
  INV_X1 U15039 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11911) );
  NAND2_X1 U15040 ( .A1(n14627), .A2(n11911), .ZN(n11912) );
  NAND2_X1 U15041 ( .A1(n16174), .A2(n11912), .ZN(n13908) );
  AND2_X1 U15042 ( .A1(n13907), .A2(n13908), .ZN(n14603) );
  INV_X1 U15043 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16248) );
  XNOR2_X1 U15044 ( .A(n16174), .B(n16248), .ZN(n14594) );
  NAND2_X1 U15045 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14646) );
  INV_X1 U15046 ( .A(n14646), .ZN(n14656) );
  NAND2_X1 U15047 ( .A1(n14558), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11917) );
  INV_X1 U15048 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14746) );
  NAND2_X1 U15049 ( .A1(n14746), .A2(n16248), .ZN(n14566) );
  INV_X1 U15050 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11915) );
  INV_X1 U15051 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14539) );
  INV_X1 U15052 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14709) );
  NAND2_X1 U15053 ( .A1(n14539), .A2(n14709), .ZN(n11916) );
  AND2_X1 U15054 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14705) );
  NAND2_X1 U15055 ( .A1(n14705), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14647) );
  NAND2_X1 U15056 ( .A1(n11917), .A2(n16173), .ZN(n14526) );
  NOR2_X1 U15057 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14690) );
  NAND2_X1 U15058 ( .A1(n16174), .A2(n14690), .ZN(n11918) );
  INV_X1 U15059 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14682) );
  NAND2_X1 U15060 ( .A1(n14508), .A2(n14682), .ZN(n11996) );
  NAND2_X1 U15061 ( .A1(n11996), .A2(n11919), .ZN(n11922) );
  AND2_X1 U15062 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14689) );
  AND2_X2 U15063 ( .A1(n11999), .A2(n14689), .ZN(n14507) );
  NOR2_X1 U15064 ( .A1(n16174), .A2(n14682), .ZN(n11920) );
  NAND2_X1 U15065 ( .A1(n11995), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11921) );
  NAND2_X1 U15066 ( .A1(n11922), .A2(n11921), .ZN(n11924) );
  NOR2_X1 U15067 ( .A1(n11926), .A2(n9789), .ZN(n13095) );
  AND2_X1 U15068 ( .A1(n13095), .A2(n13071), .ZN(n12971) );
  NAND2_X1 U15069 ( .A1(n20602), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11929) );
  NAND2_X1 U15070 ( .A1(n14792), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11928) );
  NAND2_X1 U15071 ( .A1(n11929), .A2(n11928), .ZN(n11951) );
  NAND2_X1 U15072 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20643), .ZN(
        n11950) );
  NAND2_X1 U15073 ( .A1(n11953), .A2(n11929), .ZN(n11961) );
  NAND2_X1 U15074 ( .A1(n11961), .A2(n11930), .ZN(n11932) );
  NAND2_X1 U15075 ( .A1(n20532), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11931) );
  NAND2_X1 U15076 ( .A1(n11939), .A2(n11938), .ZN(n11934) );
  NAND2_X1 U15077 ( .A1(n20528), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11933) );
  INV_X1 U15078 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16339) );
  NOR2_X1 U15079 ( .A1(n16339), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11935) );
  NAND2_X1 U15080 ( .A1(n11971), .A2(n12378), .ZN(n11979) );
  NAND2_X1 U15081 ( .A1(n12378), .A2(n11962), .ZN(n11977) );
  XNOR2_X1 U15082 ( .A(n11939), .B(n11938), .ZN(n12379) );
  NAND2_X1 U15083 ( .A1(n11940), .A2(n12379), .ZN(n11970) );
  INV_X1 U15084 ( .A(n11971), .ZN(n11943) );
  OAI21_X1 U15085 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20643), .A(
        n11950), .ZN(n11945) );
  INV_X1 U15086 ( .A(n11945), .ZN(n11941) );
  NAND2_X1 U15087 ( .A1(n11962), .A2(n11941), .ZN(n11942) );
  NAND2_X1 U15088 ( .A1(n11943), .A2(n11942), .ZN(n11948) );
  AND2_X1 U15089 ( .A1(n13482), .A2(n11133), .ZN(n11944) );
  AOI21_X1 U15090 ( .B1(n13071), .B2(n13660), .A(n11945), .ZN(n11946) );
  NAND2_X1 U15091 ( .A1(n11967), .A2(n11946), .ZN(n11947) );
  NAND2_X1 U15092 ( .A1(n11948), .A2(n11947), .ZN(n11955) );
  INV_X1 U15093 ( .A(n11955), .ZN(n11959) );
  NAND2_X1 U15094 ( .A1(n14432), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11949) );
  NAND2_X1 U15095 ( .A1(n11951), .A2(n11950), .ZN(n11952) );
  NAND2_X1 U15096 ( .A1(n11953), .A2(n11952), .ZN(n12380) );
  INV_X1 U15097 ( .A(n11956), .ZN(n11958) );
  NAND2_X1 U15098 ( .A1(n11974), .A2(n12380), .ZN(n11954) );
  AOI22_X1 U15099 ( .A1(n11956), .A2(n11955), .B1(n9750), .B2(n11954), .ZN(
        n11957) );
  AOI21_X1 U15100 ( .B1(n11959), .B2(n11958), .A(n11957), .ZN(n11969) );
  XNOR2_X1 U15101 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11960) );
  XNOR2_X1 U15102 ( .A(n11961), .B(n11960), .ZN(n12381) );
  INV_X1 U15103 ( .A(n11962), .ZN(n11963) );
  INV_X1 U15104 ( .A(n11967), .ZN(n11964) );
  AOI211_X1 U15105 ( .C1(n11974), .C2(n12381), .A(n11965), .B(n11964), .ZN(
        n11968) );
  INV_X1 U15106 ( .A(n11965), .ZN(n11966) );
  INV_X1 U15107 ( .A(n12382), .ZN(n11973) );
  NAND3_X1 U15108 ( .A1(n11974), .A2(n9749), .A3(n12382), .ZN(n11975) );
  NAND2_X1 U15109 ( .A1(n11977), .A2(n11976), .ZN(n11978) );
  NAND2_X1 U15110 ( .A1(n11986), .A2(n20678), .ZN(n20849) );
  NAND2_X1 U15111 ( .A1(n20849), .A2(n20846), .ZN(n11981) );
  NAND2_X1 U15112 ( .A1(n20846), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11983) );
  NAND2_X1 U15113 ( .A1(n20841), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n11982) );
  NAND2_X1 U15114 ( .A1(n11983), .A2(n11982), .ZN(n13185) );
  INV_X1 U15115 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n11993) );
  INV_X1 U15116 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11987) );
  INV_X1 U15117 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21036) );
  OR2_X1 U15118 ( .A1(n14779), .A2(n21036), .ZN(n14662) );
  OAI21_X1 U15119 ( .B1(n16209), .B2(n11987), .A(n14662), .ZN(n11988) );
  AOI21_X1 U15120 ( .B1(n16204), .B2(n13669), .A(n11988), .ZN(n11989) );
  NAND2_X1 U15121 ( .A1(n16204), .A2(n14191), .ZN(n11992) );
  INV_X2 U15122 ( .A(n14779), .ZN(n16319) );
  NAND2_X1 U15123 ( .A1(n16319), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14669) );
  OAI211_X1 U15124 ( .C1(n11993), .C2(n16209), .A(n11992), .B(n14669), .ZN(
        n11994) );
  AOI21_X1 U15125 ( .B1(n14387), .B2(n16205), .A(n11994), .ZN(n11997) );
  MUX2_X1 U15126 ( .A(n11999), .B(n11998), .S(n16173), .Z(n12000) );
  INV_X1 U15127 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14156) );
  XNOR2_X1 U15128 ( .A(n12000), .B(n14156), .ZN(n14704) );
  NOR2_X1 U15129 ( .A1(n14447), .A2(n14551), .ZN(n12009) );
  NAND2_X1 U15130 ( .A1(n16204), .A2(n14226), .ZN(n12007) );
  INV_X1 U15131 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12004) );
  INV_X1 U15132 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20887) );
  OR2_X1 U15133 ( .A1(n14779), .A2(n20887), .ZN(n14698) );
  OAI21_X1 U15134 ( .B1(n16209), .B2(n12004), .A(n14698), .ZN(n12005) );
  INV_X1 U15135 ( .A(n12005), .ZN(n12006) );
  NAND2_X1 U15136 ( .A1(n13269), .A2(n12039), .ZN(n12017) );
  NAND2_X1 U15137 ( .A1(n12012), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12013) );
  NAND2_X1 U15138 ( .A1(n19779), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19444) );
  NAND2_X1 U15139 ( .A1(n19444), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12014) );
  NAND3_X1 U15140 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n10331), .ZN(n19670) );
  INV_X1 U15141 ( .A(n19670), .ZN(n19673) );
  NAND2_X1 U15142 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19673), .ZN(
        n19702) );
  NAND2_X1 U15143 ( .A1(n12014), .A2(n19702), .ZN(n12015) );
  AND2_X1 U15144 ( .A1(n12015), .A2(n20068), .ZN(n15743) );
  AOI21_X1 U15145 ( .B1(n12040), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n15743), .ZN(n12016) );
  INV_X1 U15146 ( .A(n12020), .ZN(n12021) );
  NAND2_X1 U15147 ( .A1(n12421), .A2(n12039), .ZN(n12028) );
  INV_X1 U15148 ( .A(n19779), .ZN(n12024) );
  NAND2_X1 U15149 ( .A1(n12024), .A2(n20079), .ZN(n12025) );
  NAND2_X1 U15150 ( .A1(n19444), .A2(n12025), .ZN(n15738) );
  NOR2_X1 U15151 ( .A1(n19868), .A2(n15738), .ZN(n12026) );
  AOI21_X1 U15152 ( .B1(n12040), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12026), .ZN(n12027) );
  NAND2_X1 U15153 ( .A1(n12229), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12046) );
  INV_X1 U15154 ( .A(n12038), .ZN(n12030) );
  XNOR2_X2 U15155 ( .A(n12418), .B(n12030), .ZN(n13059) );
  NAND2_X1 U15156 ( .A1(n12040), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12031) );
  NAND2_X1 U15157 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20088), .ZN(
        n19495) );
  NAND2_X1 U15158 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20096), .ZN(
        n19523) );
  NAND2_X1 U15159 ( .A1(n19495), .A2(n19523), .ZN(n15737) );
  NAND2_X1 U15160 ( .A1(n20068), .A2(n15737), .ZN(n19526) );
  NAND2_X1 U15161 ( .A1(n12031), .A2(n19526), .ZN(n12032) );
  INV_X1 U15162 ( .A(n12033), .ZN(n12036) );
  INV_X1 U15163 ( .A(n12034), .ZN(n12035) );
  NAND2_X1 U15164 ( .A1(n12036), .A2(n12035), .ZN(n12037) );
  NAND2_X2 U15165 ( .A1(n12038), .A2(n12037), .ZN(n19322) );
  INV_X1 U15166 ( .A(n12039), .ZN(n12859) );
  AOI22_X1 U15167 ( .A1(n12040), .A2(n15690), .B1(n20068), .B2(n20096), .ZN(
        n12041) );
  NAND2_X1 U15168 ( .A1(n12229), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12042) );
  NAND2_X1 U15169 ( .A1(n13046), .A2(n13045), .ZN(n13044) );
  INV_X1 U15170 ( .A(n15684), .ZN(n12043) );
  NAND2_X1 U15171 ( .A1(n12043), .A2(n12042), .ZN(n12044) );
  NAND2_X1 U15172 ( .A1(n13160), .A2(n13159), .ZN(n13158) );
  INV_X1 U15173 ( .A(n12045), .ZN(n12047) );
  NAND2_X1 U15174 ( .A1(n13266), .A2(n13267), .ZN(n13265) );
  NAND2_X1 U15175 ( .A1(n12012), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12048) );
  AND2_X1 U15176 ( .A1(n12049), .A2(n12048), .ZN(n12050) );
  INV_X1 U15177 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12575) );
  INV_X1 U15178 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12051) );
  NOR2_X2 U15179 ( .A1(n15108), .A2(n12053), .ZN(n15092) );
  AND2_X1 U15180 ( .A1(n15088), .A2(n15084), .ZN(n12055) );
  AOI22_X1 U15181 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12088), .B1(
        n12150), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12059) );
  AOI22_X1 U15182 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12151), .B1(
        n12087), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12058) );
  AOI22_X1 U15183 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10552), .B1(
        n10811), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12057) );
  AOI22_X1 U15184 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n12152), .B1(
        n10806), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12056) );
  NAND4_X1 U15185 ( .A1(n12059), .A2(n12058), .A3(n12057), .A4(n12056), .ZN(
        n12065) );
  AOI22_X1 U15186 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12157), .B1(
        n12158), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12063) );
  AOI22_X1 U15187 ( .A1(n10501), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12062) );
  AOI22_X1 U15188 ( .A1(n10558), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12061) );
  AOI22_X1 U15189 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10544), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12060) );
  NAND4_X1 U15190 ( .A1(n12063), .A2(n12062), .A3(n12061), .A4(n12060), .ZN(
        n12064) );
  OR2_X1 U15191 ( .A1(n12065), .A2(n12064), .ZN(n15058) );
  AOI22_X1 U15192 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12088), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12069) );
  AOI22_X1 U15193 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12087), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12068) );
  AOI22_X1 U15194 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10811), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12067) );
  AOI22_X1 U15195 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12152), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12066) );
  NAND4_X1 U15196 ( .A1(n12069), .A2(n12068), .A3(n12067), .A4(n12066), .ZN(
        n12075) );
  AOI22_X1 U15197 ( .A1(n12158), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12157), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12073) );
  AOI22_X1 U15198 ( .A1(n10501), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12072) );
  AOI22_X1 U15199 ( .A1(n10558), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12071) );
  AOI22_X1 U15200 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12070) );
  NAND4_X1 U15201 ( .A1(n12073), .A2(n12072), .A3(n12071), .A4(n12070), .ZN(
        n12074) );
  NOR2_X1 U15202 ( .A1(n12075), .A2(n12074), .ZN(n15066) );
  NOR2_X1 U15203 ( .A1(n15066), .A2(n15073), .ZN(n15057) );
  AND2_X1 U15204 ( .A1(n15058), .A2(n15057), .ZN(n12076) );
  AOI22_X1 U15205 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n12088), .B1(
        n12150), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12080) );
  AOI22_X1 U15206 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12151), .B1(
        n12087), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12079) );
  AOI22_X1 U15207 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10552), .B1(
        n10811), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12078) );
  AOI22_X1 U15208 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n12152), .B1(
        n10806), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12077) );
  NAND4_X1 U15209 ( .A1(n12080), .A2(n12079), .A3(n12078), .A4(n12077), .ZN(
        n12086) );
  AOI22_X1 U15210 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12157), .B1(
        n12158), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12084) );
  AOI22_X1 U15211 ( .A1(n10501), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12083) );
  AOI22_X1 U15212 ( .A1(n10558), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12082) );
  AOI22_X1 U15213 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10544), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12081) );
  NAND4_X1 U15214 ( .A1(n12084), .A2(n12083), .A3(n12082), .A4(n12081), .ZN(
        n12085) );
  NOR2_X1 U15215 ( .A1(n12086), .A2(n12085), .ZN(n15050) );
  INV_X1 U15216 ( .A(n12087), .ZN(n12109) );
  NOR2_X1 U15217 ( .A1(n12109), .A2(n12482), .ZN(n12090) );
  INV_X1 U15218 ( .A(n12088), .ZN(n12742) );
  INV_X1 U15219 ( .A(n12150), .ZN(n12110) );
  OAI22_X1 U15220 ( .A1(n12464), .A2(n12742), .B1(n12110), .B2(n12462), .ZN(
        n12089) );
  AOI211_X1 U15221 ( .C1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .C2(n12151), .A(
        n12090), .B(n12089), .ZN(n12098) );
  AOI22_X1 U15222 ( .A1(n12158), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12157), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12094) );
  AOI22_X1 U15223 ( .A1(n10501), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12093) );
  AOI22_X1 U15224 ( .A1(n10558), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12092) );
  AOI22_X1 U15225 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12091) );
  AND4_X1 U15226 ( .A1(n12094), .A2(n12093), .A3(n12092), .A4(n12091), .ZN(
        n12097) );
  AOI22_X1 U15227 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10811), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12096) );
  AOI22_X1 U15228 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12152), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12095) );
  NAND4_X1 U15229 ( .A1(n12098), .A2(n12097), .A3(n12096), .A4(n12095), .ZN(
        n15043) );
  AOI22_X1 U15230 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12088), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12102) );
  AOI22_X1 U15231 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12087), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12101) );
  AOI22_X1 U15232 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10811), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12100) );
  AOI22_X1 U15233 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12152), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12099) );
  NAND4_X1 U15234 ( .A1(n12102), .A2(n12101), .A3(n12100), .A4(n12099), .ZN(
        n12108) );
  AOI22_X1 U15235 ( .A1(n12158), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12157), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12106) );
  AOI22_X1 U15236 ( .A1(n10501), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12105) );
  AOI22_X1 U15237 ( .A1(n10558), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12104) );
  AOI22_X1 U15238 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12103) );
  NAND4_X1 U15239 ( .A1(n12106), .A2(n12105), .A3(n12104), .A4(n12103), .ZN(
        n12107) );
  NOR2_X1 U15240 ( .A1(n12108), .A2(n12107), .ZN(n15035) );
  INV_X1 U15241 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12536) );
  NOR2_X1 U15242 ( .A1(n12109), .A2(n12536), .ZN(n12113) );
  INV_X1 U15243 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12537) );
  OAI22_X1 U15244 ( .A1(n12111), .A2(n12742), .B1(n12110), .B2(n12537), .ZN(
        n12112) );
  AOI211_X1 U15245 ( .C1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .C2(n12151), .A(
        n12113), .B(n12112), .ZN(n12121) );
  AOI22_X1 U15246 ( .A1(n12158), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12157), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12117) );
  AOI22_X1 U15247 ( .A1(n10501), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12116) );
  AOI22_X1 U15248 ( .A1(n10558), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12115) );
  AOI22_X1 U15249 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12114) );
  AND4_X1 U15250 ( .A1(n12117), .A2(n12116), .A3(n12115), .A4(n12114), .ZN(
        n12120) );
  AOI22_X1 U15251 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10811), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12119) );
  AOI22_X1 U15252 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12152), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12118) );
  NAND4_X1 U15253 ( .A1(n12121), .A2(n12120), .A3(n12119), .A4(n12118), .ZN(
        n15030) );
  AOI22_X1 U15254 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n12088), .B1(
        n12150), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12125) );
  AOI22_X1 U15255 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12151), .B1(
        n12087), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12124) );
  AOI22_X1 U15256 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10552), .B1(
        n10811), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12123) );
  AOI22_X1 U15257 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n12152), .B1(
        n10806), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12122) );
  NAND4_X1 U15258 ( .A1(n12125), .A2(n12124), .A3(n12123), .A4(n12122), .ZN(
        n12131) );
  AOI22_X1 U15259 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n12158), .B1(
        n12157), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12129) );
  AOI22_X1 U15260 ( .A1(n10501), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12128) );
  AOI22_X1 U15261 ( .A1(n10558), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12127) );
  AOI22_X1 U15262 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10544), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12126) );
  NAND4_X1 U15263 ( .A1(n12129), .A2(n12128), .A3(n12127), .A4(n12126), .ZN(
        n12130) );
  NOR2_X1 U15264 ( .A1(n12131), .A2(n12130), .ZN(n15021) );
  INV_X1 U15265 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n19598) );
  INV_X1 U15266 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12996) );
  OAI22_X1 U15267 ( .A1(n12284), .A2(n19598), .B1(n12282), .B2(n12996), .ZN(
        n12136) );
  INV_X1 U15268 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12134) );
  OAI22_X1 U15269 ( .A1(n12283), .A2(n12134), .B1(n12281), .B2(n19646), .ZN(
        n12135) );
  NOR2_X1 U15270 ( .A1(n12136), .A2(n12135), .ZN(n12140) );
  CLKBUF_X1 U15271 ( .A(n10371), .Z(n12137) );
  AOI22_X1 U15272 ( .A1(n12137), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9640), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12139) );
  AOI22_X1 U15273 ( .A1(n12171), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12287), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12138) );
  XNOR2_X1 U15274 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12310) );
  NAND4_X1 U15275 ( .A1(n12140), .A2(n12139), .A3(n12138), .A4(n12310), .ZN(
        n12149) );
  INV_X1 U15276 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15750) );
  INV_X1 U15277 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12141) );
  OAI22_X1 U15278 ( .A1(n12284), .A2(n15750), .B1(n12282), .B2(n12141), .ZN(
        n12144) );
  INV_X1 U15279 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12142) );
  OAI22_X1 U15280 ( .A1(n12283), .A2(n12142), .B1(n12281), .B2(n19882), .ZN(
        n12143) );
  NOR2_X1 U15281 ( .A1(n12144), .A2(n12143), .ZN(n12147) );
  AOI22_X1 U15282 ( .A1(n12137), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12299), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12146) );
  AOI22_X1 U15283 ( .A1(n12171), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12287), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12145) );
  NAND4_X1 U15284 ( .A1(n12147), .A2(n12302), .A3(n12146), .A4(n12145), .ZN(
        n12148) );
  AND2_X1 U15285 ( .A1(n12149), .A2(n12148), .ZN(n12185) );
  NAND2_X1 U15286 ( .A1(n20122), .A2(n12185), .ZN(n12165) );
  AOI22_X1 U15287 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12151), .B1(
        n12150), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12156) );
  AOI22_X1 U15288 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n12088), .B1(
        n12087), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12155) );
  AOI22_X1 U15289 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10552), .B1(
        n10811), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12154) );
  AOI22_X1 U15290 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n12152), .B1(
        n10806), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12153) );
  NAND4_X1 U15291 ( .A1(n12156), .A2(n12155), .A3(n12154), .A4(n12153), .ZN(
        n12164) );
  AOI22_X1 U15292 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n12157), .B1(
        n10558), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12162) );
  AOI22_X1 U15293 ( .A1(n10501), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12161) );
  AOI22_X1 U15294 ( .A1(n12158), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12160) );
  AOI22_X1 U15295 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10544), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12159) );
  NAND4_X1 U15296 ( .A1(n12162), .A2(n12161), .A3(n12160), .A4(n12159), .ZN(
        n12163) );
  OR2_X1 U15297 ( .A1(n12164), .A2(n12163), .ZN(n12182) );
  XNOR2_X1 U15298 ( .A(n12165), .B(n12182), .ZN(n12187) );
  XNOR2_X1 U15299 ( .A(n12166), .B(n12187), .ZN(n15014) );
  NAND2_X1 U15300 ( .A1(n15751), .A2(n12185), .ZN(n15016) );
  INV_X1 U15301 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12420) );
  OAI22_X1 U15302 ( .A1(n12282), .A2(n12441), .B1(n12281), .B2(n12420), .ZN(
        n12170) );
  INV_X1 U15303 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12168) );
  OAI22_X1 U15304 ( .A1(n12284), .A2(n12437), .B1(n12283), .B2(n12168), .ZN(
        n12169) );
  NOR2_X1 U15305 ( .A1(n12170), .A2(n12169), .ZN(n12174) );
  AOI22_X1 U15306 ( .A1(n12137), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9640), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12173) );
  AOI22_X1 U15307 ( .A1(n12171), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12287), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12172) );
  NAND4_X1 U15308 ( .A1(n12174), .A2(n12173), .A3(n12172), .A4(n12310), .ZN(
        n12181) );
  INV_X1 U15309 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12425) );
  OAI22_X1 U15310 ( .A1(n12282), .A2(n12440), .B1(n12281), .B2(n12425), .ZN(
        n12176) );
  INV_X1 U15311 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12446) );
  OAI22_X1 U15312 ( .A1(n12284), .A2(n15754), .B1(n12283), .B2(n12446), .ZN(
        n12175) );
  NOR2_X1 U15313 ( .A1(n12176), .A2(n12175), .ZN(n12179) );
  AOI22_X1 U15314 ( .A1(n12137), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9640), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12178) );
  AOI22_X1 U15315 ( .A1(n12171), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12287), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12177) );
  NAND4_X1 U15316 ( .A1(n12179), .A2(n12178), .A3(n12302), .A4(n12177), .ZN(
        n12180) );
  NAND2_X1 U15317 ( .A1(n12181), .A2(n12180), .ZN(n12189) );
  NAND2_X1 U15318 ( .A1(n12182), .A2(n12185), .ZN(n12190) );
  XOR2_X1 U15319 ( .A(n12189), .B(n12190), .Z(n12183) );
  NAND2_X1 U15320 ( .A1(n12183), .A2(n12229), .ZN(n15005) );
  INV_X1 U15321 ( .A(n12189), .ZN(n12184) );
  NAND2_X1 U15322 ( .A1(n15751), .A2(n12184), .ZN(n15007) );
  INV_X1 U15323 ( .A(n12185), .ZN(n12186) );
  NOR2_X1 U15324 ( .A1(n12190), .A2(n12189), .ZN(n12211) );
  INV_X1 U15325 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12192) );
  INV_X1 U15326 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12191) );
  OAI22_X1 U15327 ( .A1(n12282), .A2(n12192), .B1(n12281), .B2(n12191), .ZN(
        n12196) );
  INV_X1 U15328 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12194) );
  INV_X1 U15329 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12193) );
  OAI22_X1 U15330 ( .A1(n12284), .A2(n12194), .B1(n12283), .B2(n12193), .ZN(
        n12195) );
  NOR2_X1 U15331 ( .A1(n12196), .A2(n12195), .ZN(n12199) );
  AOI22_X1 U15332 ( .A1(n12137), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9641), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12198) );
  AOI22_X1 U15333 ( .A1(n12171), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12287), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12197) );
  NAND4_X1 U15334 ( .A1(n12199), .A2(n12198), .A3(n12197), .A4(n12310), .ZN(
        n12210) );
  INV_X1 U15335 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12201) );
  INV_X1 U15336 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12200) );
  OAI22_X1 U15337 ( .A1(n12282), .A2(n12201), .B1(n12281), .B2(n12200), .ZN(
        n12205) );
  INV_X1 U15338 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12203) );
  INV_X1 U15339 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12202) );
  OAI22_X1 U15340 ( .A1(n12284), .A2(n12203), .B1(n12283), .B2(n12202), .ZN(
        n12204) );
  NOR2_X1 U15341 ( .A1(n12205), .A2(n12204), .ZN(n12208) );
  AOI22_X1 U15342 ( .A1(n12137), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12299), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12207) );
  AOI22_X1 U15343 ( .A1(n12171), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12287), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12206) );
  NAND4_X1 U15344 ( .A1(n12208), .A2(n12207), .A3(n12302), .A4(n12206), .ZN(
        n12209) );
  NAND2_X1 U15345 ( .A1(n12211), .A2(n12213), .ZN(n12230) );
  OAI211_X1 U15346 ( .C1(n12211), .C2(n12213), .A(n12229), .B(n12230), .ZN(
        n12215) );
  INV_X1 U15347 ( .A(n12213), .ZN(n12214) );
  NOR2_X1 U15348 ( .A1(n20122), .A2(n12214), .ZN(n14997) );
  NAND2_X1 U15349 ( .A1(n14995), .A2(n14997), .ZN(n14996) );
  INV_X1 U15350 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12477) );
  OAI22_X1 U15351 ( .A1(n12282), .A2(n12464), .B1(n12281), .B2(n12477), .ZN(
        n12218) );
  INV_X1 U15352 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12463) );
  OAI22_X1 U15353 ( .A1(n12284), .A2(n12481), .B1(n12283), .B2(n12463), .ZN(
        n12217) );
  NOR2_X1 U15354 ( .A1(n12218), .A2(n12217), .ZN(n12221) );
  AOI22_X1 U15355 ( .A1(n12137), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12299), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12220) );
  AOI22_X1 U15356 ( .A1(n12171), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12287), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12219) );
  NAND4_X1 U15357 ( .A1(n12221), .A2(n12220), .A3(n12219), .A4(n12310), .ZN(
        n12228) );
  INV_X1 U15358 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12474) );
  OAI22_X1 U15359 ( .A1(n12282), .A2(n12462), .B1(n12281), .B2(n12474), .ZN(
        n12223) );
  INV_X1 U15360 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12480) );
  OAI22_X1 U15361 ( .A1(n12284), .A2(n12482), .B1(n12283), .B2(n12480), .ZN(
        n12222) );
  NOR2_X1 U15362 ( .A1(n12223), .A2(n12222), .ZN(n12226) );
  AOI22_X1 U15363 ( .A1(n12137), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9640), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12225) );
  AOI22_X1 U15364 ( .A1(n12171), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12287), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12224) );
  NAND4_X1 U15365 ( .A1(n12226), .A2(n12225), .A3(n12302), .A4(n12224), .ZN(
        n12227) );
  NAND2_X1 U15366 ( .A1(n12228), .A2(n12227), .ZN(n12232) );
  INV_X1 U15367 ( .A(n12229), .ZN(n12256) );
  AOI21_X1 U15368 ( .B1(n12230), .B2(n12232), .A(n12256), .ZN(n12231) );
  NAND2_X1 U15369 ( .A1(n12231), .A2(n12257), .ZN(n12234) );
  NOR2_X1 U15370 ( .A1(n20122), .A2(n12232), .ZN(n14989) );
  OAI22_X1 U15371 ( .A1(n12238), .A2(n12282), .B1(n12284), .B2(n12237), .ZN(
        n12241) );
  INV_X1 U15372 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12239) );
  INV_X1 U15373 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n19655) );
  OAI22_X1 U15374 ( .A1(n12283), .A2(n12239), .B1(n12281), .B2(n19655), .ZN(
        n12240) );
  NOR2_X1 U15375 ( .A1(n12241), .A2(n12240), .ZN(n12244) );
  AOI22_X1 U15376 ( .A1(n12137), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9641), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12243) );
  AOI22_X1 U15377 ( .A1(n12171), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12287), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12242) );
  NAND4_X1 U15378 ( .A1(n12244), .A2(n12243), .A3(n12242), .A4(n12310), .ZN(
        n12255) );
  INV_X1 U15379 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12245) );
  OAI22_X1 U15380 ( .A1(n12282), .A2(n12246), .B1(n12281), .B2(n12245), .ZN(
        n12250) );
  INV_X1 U15381 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12247) );
  OAI22_X1 U15382 ( .A1(n12284), .A2(n12248), .B1(n12283), .B2(n12247), .ZN(
        n12249) );
  NOR2_X1 U15383 ( .A1(n12250), .A2(n12249), .ZN(n12253) );
  AOI22_X1 U15384 ( .A1(n12137), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9641), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12252) );
  AOI22_X1 U15385 ( .A1(n12171), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12287), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12251) );
  NAND4_X1 U15386 ( .A1(n12253), .A2(n12252), .A3(n12302), .A4(n12251), .ZN(
        n12254) );
  NAND2_X1 U15387 ( .A1(n12255), .A2(n12254), .ZN(n12260) );
  NOR2_X1 U15388 ( .A1(n12257), .A2(n12260), .ZN(n14971) );
  NAND2_X2 U15389 ( .A1(n12259), .A2(n12258), .ZN(n14973) );
  NOR2_X1 U15390 ( .A1(n20122), .A2(n12260), .ZN(n14981) );
  INV_X1 U15391 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12545) );
  OAI22_X1 U15392 ( .A1(n12282), .A2(n12111), .B1(n12281), .B2(n12545), .ZN(
        n12262) );
  INV_X1 U15393 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12526) );
  INV_X1 U15394 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12519) );
  OAI22_X1 U15395 ( .A1(n12284), .A2(n12526), .B1(n12283), .B2(n12519), .ZN(
        n12261) );
  NOR2_X1 U15396 ( .A1(n12262), .A2(n12261), .ZN(n12265) );
  AOI22_X1 U15397 ( .A1(n12137), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12299), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12264) );
  AOI22_X1 U15398 ( .A1(n12171), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12287), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12263) );
  NAND4_X1 U15399 ( .A1(n12265), .A2(n12264), .A3(n12263), .A4(n12310), .ZN(
        n12273) );
  INV_X1 U15400 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12527) );
  OAI22_X1 U15401 ( .A1(n12282), .A2(n12537), .B1(n12281), .B2(n12527), .ZN(
        n12268) );
  INV_X1 U15402 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12522) );
  OAI22_X1 U15403 ( .A1(n12284), .A2(n12536), .B1(n12283), .B2(n12522), .ZN(
        n12267) );
  NOR2_X1 U15404 ( .A1(n12268), .A2(n12267), .ZN(n12271) );
  AOI22_X1 U15405 ( .A1(n12137), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9640), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12270) );
  AOI22_X1 U15406 ( .A1(n12171), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12287), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12269) );
  NAND4_X1 U15407 ( .A1(n12271), .A2(n12270), .A3(n12302), .A4(n12269), .ZN(
        n12272) );
  NAND2_X1 U15408 ( .A1(n12273), .A2(n12272), .ZN(n12293) );
  INV_X1 U15409 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12566) );
  INV_X1 U15410 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12582) );
  OAI22_X1 U15411 ( .A1(n12284), .A2(n12566), .B1(n12281), .B2(n12582), .ZN(
        n12277) );
  INV_X1 U15412 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12274) );
  OAI22_X1 U15413 ( .A1(n12282), .A2(n12575), .B1(n12283), .B2(n12274), .ZN(
        n12276) );
  NOR2_X1 U15414 ( .A1(n12277), .A2(n12276), .ZN(n12280) );
  AOI22_X1 U15415 ( .A1(n12137), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12299), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12279) );
  AOI22_X1 U15416 ( .A1(n12171), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12287), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12278) );
  NAND4_X1 U15417 ( .A1(n12280), .A2(n12279), .A3(n12278), .A4(n12310), .ZN(
        n12292) );
  INV_X1 U15418 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12563) );
  INV_X1 U15419 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12571) );
  OAI22_X1 U15420 ( .A1(n12282), .A2(n12563), .B1(n12281), .B2(n12571), .ZN(
        n12286) );
  INV_X1 U15421 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12576) );
  INV_X1 U15422 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12577) );
  OAI22_X1 U15423 ( .A1(n12284), .A2(n12576), .B1(n12283), .B2(n12577), .ZN(
        n12285) );
  NOR2_X1 U15424 ( .A1(n12286), .A2(n12285), .ZN(n12290) );
  AOI22_X1 U15425 ( .A1(n12137), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9640), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12289) );
  AOI22_X1 U15426 ( .A1(n12171), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12287), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12288) );
  NAND4_X1 U15427 ( .A1(n12290), .A2(n12289), .A3(n12302), .A4(n12288), .ZN(
        n12291) );
  NAND2_X1 U15428 ( .A1(n12292), .A2(n12291), .ZN(n12296) );
  INV_X1 U15429 ( .A(n12293), .ZN(n14974) );
  AND2_X1 U15430 ( .A1(n20122), .A2(n14974), .ZN(n12294) );
  NAND2_X1 U15431 ( .A1(n14971), .A2(n12294), .ZN(n12295) );
  NOR2_X1 U15432 ( .A1(n12295), .A2(n12296), .ZN(n12297) );
  AOI21_X1 U15433 ( .B1(n12296), .B2(n12295), .A(n12297), .ZN(n14966) );
  NAND2_X1 U15434 ( .A1(n14967), .A2(n14966), .ZN(n14968) );
  INV_X1 U15435 ( .A(n12297), .ZN(n12298) );
  NAND2_X1 U15436 ( .A1(n14968), .A2(n12298), .ZN(n12319) );
  AOI22_X1 U15437 ( .A1(n12137), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9641), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12301) );
  AOI22_X1 U15438 ( .A1(n12171), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12287), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12300) );
  NAND2_X1 U15439 ( .A1(n12301), .A2(n12300), .ZN(n12316) );
  AOI22_X1 U15440 ( .A1(n12309), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9643), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12304) );
  AOI22_X1 U15441 ( .A1(n12308), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10488), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12303) );
  NAND3_X1 U15442 ( .A1(n12304), .A2(n12303), .A3(n12302), .ZN(n12315) );
  INV_X1 U15443 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n19634) );
  AOI22_X1 U15444 ( .A1(n12171), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12287), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12306) );
  NAND2_X1 U15445 ( .A1(n12137), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12305) );
  OAI211_X1 U15446 ( .C1(n12307), .C2(n19634), .A(n12306), .B(n12305), .ZN(
        n12314) );
  AOI22_X1 U15447 ( .A1(n12308), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9643), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12312) );
  AOI22_X1 U15448 ( .A1(n12309), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10488), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12311) );
  NAND3_X1 U15449 ( .A1(n12312), .A2(n12311), .A3(n12310), .ZN(n12313) );
  OAI22_X1 U15450 ( .A1(n12316), .A2(n12315), .B1(n12314), .B2(n12313), .ZN(
        n12317) );
  XNOR2_X1 U15451 ( .A(n12319), .B(n12318), .ZN(n12417) );
  NAND2_X1 U15452 ( .A1(n12321), .A2(n12320), .ZN(n12744) );
  NAND2_X1 U15453 ( .A1(n12744), .A2(n12765), .ZN(n12332) );
  OAI21_X1 U15454 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20096), .A(
        n12322), .ZN(n12740) );
  INV_X1 U15455 ( .A(n12740), .ZN(n12326) );
  INV_X1 U15456 ( .A(n12747), .ZN(n12323) );
  AND2_X1 U15457 ( .A1(n12326), .A2(n12323), .ZN(n12328) );
  INV_X1 U15458 ( .A(n12324), .ZN(n12325) );
  OAI211_X1 U15459 ( .C1(n20122), .C2(n12326), .A(n20115), .B(n12325), .ZN(
        n12327) );
  AND2_X1 U15460 ( .A1(n10643), .A2(n20122), .ZN(n12330) );
  MUX2_X1 U15461 ( .A(n12330), .B(n20103), .S(n12737), .Z(n12331) );
  MUX2_X1 U15462 ( .A(n15859), .B(n12333), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n12734) );
  NAND2_X1 U15463 ( .A1(n12732), .A2(n15751), .ZN(n12345) );
  AOI21_X1 U15464 ( .B1(n12345), .B2(n20115), .A(n12335), .ZN(n12338) );
  NOR2_X1 U15465 ( .A1(n20122), .A2(n20115), .ZN(n20100) );
  OAI21_X1 U15466 ( .B1(n12336), .B2(n12413), .A(n20100), .ZN(n12769) );
  OAI211_X1 U15467 ( .C1(n12338), .C2(n19459), .A(n12769), .B(n12337), .ZN(
        n12339) );
  INV_X1 U15468 ( .A(n12339), .ZN(n12344) );
  NAND2_X1 U15469 ( .A1(n12341), .A2(n12777), .ZN(n12342) );
  NAND2_X1 U15470 ( .A1(n12340), .A2(n12342), .ZN(n12343) );
  NAND2_X1 U15471 ( .A1(n12344), .A2(n12343), .ZN(n12756) );
  NAND2_X1 U15472 ( .A1(n13562), .A2(n12796), .ZN(n12912) );
  NAND2_X1 U15473 ( .A1(n12883), .A2(n20114), .ZN(n12910) );
  OAI22_X1 U15474 ( .A1(n13568), .A2(n13563), .B1(n12912), .B2(n12910), .ZN(
        n13514) );
  INV_X1 U15475 ( .A(n12347), .ZN(n12349) );
  NOR2_X1 U15476 ( .A1(n12349), .A2(n12348), .ZN(n12350) );
  AND2_X1 U15477 ( .A1(n12727), .A2(n19486), .ZN(n12353) );
  NOR4_X1 U15478 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12357) );
  NOR4_X1 U15479 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12356) );
  NOR4_X1 U15480 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12355) );
  NOR4_X1 U15481 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12354) );
  NAND4_X1 U15482 ( .A1(n12357), .A2(n12356), .A3(n12355), .A4(n12354), .ZN(
        n12362) );
  NOR4_X1 U15483 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n12360) );
  NOR4_X1 U15484 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12359) );
  NOR4_X1 U15485 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12358) );
  NAND4_X1 U15486 ( .A1(n12360), .A2(n12359), .A3(n12358), .A4(n20001), .ZN(
        n12361) );
  INV_X1 U15487 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n16708) );
  OR2_X1 U15488 ( .A1(n15707), .A2(n16708), .ZN(n12365) );
  NAND2_X1 U15489 ( .A1(n15707), .A2(BUF2_REG_14__SCAN_IN), .ZN(n12364) );
  NAND2_X1 U15490 ( .A1(n12365), .A2(n12364), .ZN(n19341) );
  XNOR2_X1 U15491 ( .A(n15121), .B(n12366), .ZN(n14815) );
  INV_X1 U15492 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n12367) );
  OAI22_X1 U15493 ( .A1(n14815), .A2(n19358), .B1(n19357), .B2(n12367), .ZN(
        n12368) );
  AOI21_X1 U15494 ( .B1(n16417), .B2(n19341), .A(n12368), .ZN(n12371) );
  AND2_X1 U15495 ( .A1(n12012), .A2(n19486), .ZN(n12369) );
  NOR2_X2 U15496 ( .A1(n13052), .A2(n15709), .ZN(n16418) );
  NOR2_X2 U15497 ( .A1(n13052), .A2(n15707), .ZN(n16419) );
  AOI22_X1 U15498 ( .A1(n16418), .A2(BUF2_REG_30__SCAN_IN), .B1(n16419), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n12370) );
  OAI21_X1 U15499 ( .B1(n12417), .B2(n15230), .A(n12372), .ZN(P2_U2889) );
  NAND2_X1 U15500 ( .A1(n9666), .A2(n20850), .ZN(n12375) );
  AND2_X1 U15501 ( .A1(n11085), .A2(n13649), .ZN(n12374) );
  NAND2_X1 U15502 ( .A1(n13218), .A2(n12374), .ZN(n13227) );
  OAI21_X1 U15503 ( .B1(n12373), .B2(n12375), .A(n13227), .ZN(n12376) );
  NAND2_X1 U15504 ( .A1(n12376), .A2(n9938), .ZN(n12386) );
  INV_X1 U15505 ( .A(n12377), .ZN(n16335) );
  INV_X1 U15506 ( .A(n20850), .ZN(n20840) );
  INV_X1 U15507 ( .A(n12378), .ZN(n12384) );
  OR4_X1 U15508 ( .A1(n12382), .A2(n12381), .A3(n12380), .A4(n12379), .ZN(
        n12383) );
  NAND2_X1 U15509 ( .A1(n12384), .A2(n12383), .ZN(n12974) );
  NOR2_X1 U15510 ( .A1(n20840), .A2(n12974), .ZN(n13210) );
  NAND2_X1 U15511 ( .A1(n16335), .A2(n13210), .ZN(n12385) );
  INV_X1 U15512 ( .A(n12387), .ZN(n12389) );
  NOR2_X1 U15513 ( .A1(n11138), .A2(n16100), .ZN(n12388) );
  NAND4_X1 U15514 ( .A1(n12389), .A2(n13433), .A3(n13329), .A4(n12388), .ZN(
        n13133) );
  NAND2_X1 U15515 ( .A1(n14498), .A2(n13433), .ZN(n12408) );
  NOR4_X1 U15516 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12395) );
  NOR4_X1 U15517 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12394) );
  NOR4_X1 U15518 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12393) );
  NOR4_X1 U15519 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12392) );
  AND4_X1 U15520 ( .A1(n12395), .A2(n12394), .A3(n12393), .A4(n12392), .ZN(
        n12400) );
  NOR4_X1 U15521 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n12398) );
  NOR4_X1 U15522 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12397) );
  NOR4_X1 U15523 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12396) );
  INV_X1 U15524 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20770) );
  AND4_X1 U15525 ( .A1(n12398), .A2(n12397), .A3(n12396), .A4(n20770), .ZN(
        n12399) );
  NAND2_X1 U15526 ( .A1(n12400), .A2(n12399), .ZN(n12401) );
  NOR3_X1 U15527 ( .A1(n14502), .A2(n14438), .A3(n13212), .ZN(n12402) );
  AOI22_X1 U15528 ( .A1(n14491), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14502), .ZN(n12403) );
  INV_X1 U15529 ( .A(n12403), .ZN(n12406) );
  NOR2_X1 U15530 ( .A1(n13212), .A2(n13418), .ZN(n12404) );
  NAND2_X1 U15531 ( .A1(n14498), .A2(n12404), .ZN(n14437) );
  INV_X1 U15532 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n19484) );
  NOR2_X1 U15533 ( .A1(n14437), .A2(n19484), .ZN(n12405) );
  NOR2_X1 U15534 ( .A1(n12406), .A2(n12405), .ZN(n12407) );
  OAI21_X1 U15535 ( .B1(n14186), .B2(n12408), .A(n12407), .ZN(P1_U2873) );
  INV_X1 U15536 ( .A(n12410), .ZN(n12411) );
  AND2_X1 U15537 ( .A1(n12409), .A2(n12411), .ZN(n13520) );
  NAND2_X1 U15538 ( .A1(n13568), .A2(n13520), .ZN(n13512) );
  NAND2_X1 U15539 ( .A1(n13512), .A2(n12782), .ZN(n12412) );
  NAND2_X1 U15540 ( .A1(n14807), .A2(n15116), .ZN(n12416) );
  NAND2_X1 U15541 ( .A1(n15089), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12415) );
  OAI21_X1 U15542 ( .B1(n12417), .B2(n15106), .A(n10267), .ZN(P2_U2857) );
  INV_X1 U15543 ( .A(n12421), .ZN(n12429) );
  OR2_X2 U15544 ( .A1(n13269), .A2(n12429), .ZN(n12445) );
  NAND2_X1 U15545 ( .A1(n13059), .A2(n19322), .ZN(n12436) );
  OR2_X2 U15546 ( .A1(n12445), .A2(n12436), .ZN(n12543) );
  OR2_X1 U15547 ( .A1(n12418), .A2(n19322), .ZN(n12448) );
  NOR2_X2 U15548 ( .A1(n12445), .A2(n12448), .ZN(n19668) );
  NAND2_X1 U15549 ( .A1(n19668), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12419) );
  OAI211_X1 U15550 ( .C1(n12420), .C2(n12543), .A(n12419), .B(n20122), .ZN(
        n12428) );
  OR2_X1 U15551 ( .A1(n12422), .A2(n19322), .ZN(n12444) );
  NOR2_X1 U15553 ( .A1(n12428), .A2(n12427), .ZN(n12459) );
  INV_X1 U15554 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12431) );
  OAI22_X1 U15555 ( .A1(n12431), .A2(n19494), .B1(n15728), .B2(n12430), .ZN(
        n12435) );
  INV_X1 U15556 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12433) );
  OAI22_X1 U15558 ( .A1(n12433), .A2(n19732), .B1(n12540), .B2(n12432), .ZN(
        n12434) );
  NOR2_X1 U15559 ( .A1(n12435), .A2(n12434), .ZN(n12458) );
  INV_X1 U15560 ( .A(n19322), .ZN(n16591) );
  OR2_X2 U15561 ( .A1(n12445), .A2(n12450), .ZN(n19585) );
  OAI22_X1 U15562 ( .A1(n12438), .A2(n19528), .B1(n19585), .B2(n12437), .ZN(
        n12443) );
  OAI22_X1 U15564 ( .A1(n12441), .A2(n19448), .B1(n19697), .B2(n12440), .ZN(
        n12442) );
  NOR2_X1 U15565 ( .A1(n12443), .A2(n12442), .ZN(n12457) );
  OAI22_X1 U15567 ( .A1(n12447), .A2(n12531), .B1(n12521), .B2(n12446), .ZN(
        n12455) );
  INV_X1 U15568 ( .A(n12450), .ZN(n12451) );
  OAI22_X1 U15570 ( .A1(n12453), .A2(n12532), .B1(n12535), .B2(n15754), .ZN(
        n12454) );
  NOR2_X1 U15571 ( .A1(n12455), .A2(n12454), .ZN(n12456) );
  INV_X1 U15572 ( .A(n12963), .ZN(n12814) );
  NAND2_X1 U15573 ( .A1(n12814), .A2(n12815), .ZN(n12821) );
  INV_X1 U15574 ( .A(n12460), .ZN(n12820) );
  NAND2_X1 U15575 ( .A1(n12821), .A2(n12820), .ZN(n12461) );
  OAI22_X1 U15576 ( .A1(n12463), .A2(n12518), .B1(n19697), .B2(n12462), .ZN(
        n12467) );
  OAI22_X1 U15577 ( .A1(n12465), .A2(n19528), .B1(n19448), .B2(n12464), .ZN(
        n12466) );
  NOR2_X1 U15578 ( .A1(n12467), .A2(n12466), .ZN(n12489) );
  INV_X1 U15579 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12469) );
  OAI22_X1 U15580 ( .A1(n12469), .A2(n19494), .B1(n12540), .B2(n12468), .ZN(
        n12473) );
  OAI22_X1 U15581 ( .A1(n12471), .A2(n12532), .B1(n15728), .B2(n12470), .ZN(
        n12472) );
  NOR2_X1 U15582 ( .A1(n12473), .A2(n12472), .ZN(n12488) );
  INV_X1 U15583 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12475) );
  OAI22_X1 U15584 ( .A1(n12475), .A2(n19732), .B1(n19875), .B2(n12474), .ZN(
        n12479) );
  INV_X1 U15585 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12476) );
  OAI22_X1 U15586 ( .A1(n12477), .A2(n12543), .B1(n19830), .B2(n12476), .ZN(
        n12478) );
  NOR2_X1 U15587 ( .A1(n12479), .A2(n12478), .ZN(n12487) );
  OAI22_X1 U15588 ( .A1(n12481), .A2(n19585), .B1(n12521), .B2(n12480), .ZN(
        n12485) );
  INV_X1 U15589 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12483) );
  OAI22_X1 U15590 ( .A1(n12483), .A2(n12531), .B1(n12535), .B2(n12482), .ZN(
        n12484) );
  NOR2_X1 U15591 ( .A1(n12485), .A2(n12484), .ZN(n12486) );
  INV_X1 U15592 ( .A(n12490), .ZN(n12491) );
  NAND2_X1 U15593 ( .A1(n12491), .A2(n15751), .ZN(n12492) );
  INV_X1 U15594 ( .A(n12496), .ZN(n12497) );
  NAND2_X1 U15595 ( .A1(n12497), .A2(n12506), .ZN(n12498) );
  NAND2_X1 U15596 ( .A1(n12511), .A2(n12498), .ZN(n14936) );
  MUX2_X1 U15597 ( .A(n12740), .B(n12816), .S(n20103), .Z(n12748) );
  INV_X1 U15598 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13000) );
  MUX2_X1 U15599 ( .A(n12748), .B(n13000), .S(n12727), .Z(n12961) );
  NOR2_X1 U15600 ( .A1(n12961), .A2(n16585), .ZN(n13006) );
  INV_X1 U15601 ( .A(n13006), .ZN(n12505) );
  INV_X1 U15602 ( .A(n12507), .ZN(n12501) );
  AND2_X1 U15603 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n12499) );
  NAND2_X1 U15604 ( .A1(n12727), .A2(n12499), .ZN(n12500) );
  NAND2_X1 U15605 ( .A1(n12501), .A2(n12500), .ZN(n14952) );
  INV_X1 U15606 ( .A(n14952), .ZN(n12502) );
  NAND2_X1 U15607 ( .A1(n12502), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12504) );
  AND2_X1 U15608 ( .A1(n14952), .A2(n15692), .ZN(n12503) );
  AOI21_X1 U15609 ( .B1(n12505), .B2(n12504), .A(n12503), .ZN(n12982) );
  OAI21_X1 U15610 ( .B1(n12508), .B2(n12507), .A(n12506), .ZN(n14942) );
  XNOR2_X1 U15611 ( .A(n14942), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12981) );
  NAND2_X1 U15612 ( .A1(n12982), .A2(n12981), .ZN(n12983) );
  INV_X1 U15613 ( .A(n14942), .ZN(n12509) );
  NAND2_X1 U15614 ( .A1(n12509), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12510) );
  NAND2_X1 U15615 ( .A1(n12983), .A2(n12510), .ZN(n13703) );
  INV_X1 U15616 ( .A(n12557), .ZN(n12514) );
  NAND2_X1 U15617 ( .A1(n12512), .A2(n12511), .ZN(n12513) );
  NAND2_X1 U15618 ( .A1(n12514), .A2(n12513), .ZN(n14925) );
  XNOR2_X1 U15619 ( .A(n14925), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n15672) );
  INV_X1 U15620 ( .A(n14925), .ZN(n12515) );
  NAND2_X1 U15621 ( .A1(n12515), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12516) );
  INV_X1 U15622 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12520) );
  OAI22_X1 U15623 ( .A1(n12520), .A2(n19528), .B1(n12518), .B2(n12519), .ZN(
        n12524) );
  OAI22_X1 U15624 ( .A1(n12111), .A2(n19448), .B1(n12521), .B2(n12522), .ZN(
        n12523) );
  NOR2_X1 U15625 ( .A1(n12524), .A2(n12523), .ZN(n12551) );
  INV_X1 U15626 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12525) );
  OAI22_X1 U15627 ( .A1(n12526), .A2(n19585), .B1(n15728), .B2(n12525), .ZN(
        n12530) );
  OAI22_X1 U15628 ( .A1(n12528), .A2(n19830), .B1(n19875), .B2(n12527), .ZN(
        n12529) );
  NOR2_X1 U15629 ( .A1(n12530), .A2(n12529), .ZN(n12550) );
  INV_X1 U15630 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12533) );
  OAI22_X1 U15631 ( .A1(n12534), .A2(n12531), .B1(n12532), .B2(n12533), .ZN(
        n12539) );
  OAI22_X1 U15632 ( .A1(n12537), .A2(n19697), .B1(n12535), .B2(n12536), .ZN(
        n12538) );
  NOR2_X1 U15633 ( .A1(n12539), .A2(n12538), .ZN(n12549) );
  INV_X1 U15634 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12542) );
  INV_X1 U15635 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12541) );
  OAI22_X1 U15636 ( .A1(n12542), .A2(n19494), .B1(n12540), .B2(n12541), .ZN(
        n12547) );
  INV_X1 U15637 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12544) );
  OAI22_X1 U15638 ( .A1(n12545), .A2(n12543), .B1(n19732), .B2(n12544), .ZN(
        n12546) );
  NOR2_X1 U15639 ( .A1(n12547), .A2(n12546), .ZN(n12548) );
  NAND4_X1 U15640 ( .A1(n12551), .A2(n12550), .A3(n12549), .A4(n12548), .ZN(
        n12555) );
  INV_X1 U15641 ( .A(n12552), .ZN(n12553) );
  NAND2_X1 U15642 ( .A1(n12553), .A2(n15751), .ZN(n12554) );
  XNOR2_X2 U15643 ( .A(n12562), .B(n9733), .ZN(n12835) );
  NAND2_X1 U15644 ( .A1(n12835), .A2(n12495), .ZN(n12558) );
  XNOR2_X1 U15645 ( .A(n12557), .B(n12556), .ZN(n14909) );
  NAND2_X1 U15646 ( .A1(n15417), .A2(n15416), .ZN(n12561) );
  NAND2_X1 U15647 ( .A1(n12559), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12560) );
  NAND2_X1 U15648 ( .A1(n12561), .A2(n12560), .ZN(n15409) );
  INV_X1 U15649 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12564) );
  OAI22_X1 U15650 ( .A1(n12564), .A2(n19528), .B1(n19697), .B2(n12563), .ZN(
        n12568) );
  INV_X1 U15651 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12565) );
  OAI22_X1 U15652 ( .A1(n12566), .A2(n19585), .B1(n15728), .B2(n12565), .ZN(
        n12567) );
  NOR2_X1 U15653 ( .A1(n12568), .A2(n12567), .ZN(n12588) );
  INV_X1 U15654 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12570) );
  INV_X1 U15655 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12569) );
  OAI22_X1 U15656 ( .A1(n12570), .A2(n19494), .B1(n12540), .B2(n12569), .ZN(
        n12574) );
  OAI22_X1 U15657 ( .A1(n12572), .A2(n19830), .B1(n19875), .B2(n12571), .ZN(
        n12573) );
  NOR2_X1 U15658 ( .A1(n12574), .A2(n12573), .ZN(n12587) );
  OAI22_X1 U15659 ( .A1(n12575), .A2(n19448), .B1(n12518), .B2(n12274), .ZN(
        n12579) );
  OAI22_X1 U15660 ( .A1(n12577), .A2(n12521), .B1(n12535), .B2(n12576), .ZN(
        n12578) );
  NOR2_X1 U15661 ( .A1(n12579), .A2(n12578), .ZN(n12586) );
  INV_X1 U15662 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12580) );
  OAI22_X1 U15663 ( .A1(n15720), .A2(n12531), .B1(n12532), .B2(n12580), .ZN(
        n12584) );
  INV_X1 U15664 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12581) );
  OAI22_X1 U15665 ( .A1(n12582), .A2(n12543), .B1(n19732), .B2(n12581), .ZN(
        n12583) );
  NOR2_X1 U15666 ( .A1(n12584), .A2(n12583), .ZN(n12585) );
  NAND4_X1 U15667 ( .A1(n12588), .A2(n12587), .A3(n12586), .A4(n12585), .ZN(
        n12591) );
  NAND2_X1 U15668 ( .A1(n12589), .A2(n15751), .ZN(n12590) );
  NAND2_X1 U15669 ( .A1(n12834), .A2(n12495), .ZN(n12596) );
  INV_X1 U15670 ( .A(n12605), .ZN(n12595) );
  NAND2_X1 U15671 ( .A1(n12593), .A2(n12592), .ZN(n12594) );
  NAND2_X1 U15672 ( .A1(n12595), .A2(n12594), .ZN(n19305) );
  NAND2_X1 U15673 ( .A1(n12596), .A2(n19305), .ZN(n12597) );
  XNOR2_X1 U15674 ( .A(n12597), .B(n12799), .ZN(n15408) );
  NAND2_X1 U15675 ( .A1(n15409), .A2(n15408), .ZN(n12599) );
  NAND2_X1 U15676 ( .A1(n12597), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12598) );
  NAND2_X1 U15677 ( .A1(n12601), .A2(n12600), .ZN(n12602) );
  NAND2_X1 U15678 ( .A1(n12610), .A2(n12602), .ZN(n19290) );
  NOR2_X1 U15679 ( .A1(n19290), .A2(n12495), .ZN(n12606) );
  NAND2_X1 U15680 ( .A1(n12606), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15386) );
  INV_X1 U15681 ( .A(n12603), .ZN(n12604) );
  XNOR2_X1 U15682 ( .A(n12605), .B(n12604), .ZN(n14898) );
  NAND2_X1 U15683 ( .A1(n14898), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15399) );
  INV_X1 U15684 ( .A(n12606), .ZN(n12607) );
  NAND2_X1 U15685 ( .A1(n12607), .A2(n16561), .ZN(n15385) );
  INV_X1 U15686 ( .A(n14898), .ZN(n12608) );
  NAND2_X1 U15687 ( .A1(n12608), .A2(n16558), .ZN(n15398) );
  AND2_X1 U15688 ( .A1(n15385), .A2(n15398), .ZN(n12609) );
  NAND2_X1 U15689 ( .A1(n12727), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12611) );
  MUX2_X1 U15690 ( .A(n12727), .B(n12611), .S(n12610), .Z(n12612) );
  AOI21_X1 U15691 ( .B1(n14883), .B2(n10861), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15632) );
  NAND2_X1 U15692 ( .A1(n12727), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12614) );
  MUX2_X1 U15693 ( .A(n12614), .B(P2_EBX_REG_10__SCAN_IN), .S(n12613), .Z(
        n12615) );
  NAND2_X1 U15694 ( .A1(n12615), .A2(n12706), .ZN(n14874) );
  OR2_X1 U15695 ( .A1(n14874), .A2(n12495), .ZN(n12616) );
  NAND2_X1 U15696 ( .A1(n12616), .A2(n16545), .ZN(n16483) );
  INV_X1 U15697 ( .A(n12617), .ZN(n12618) );
  NAND2_X1 U15698 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n12618), .ZN(n12619) );
  NOR2_X1 U15699 ( .A1(n10508), .A2(n12619), .ZN(n12620) );
  NOR2_X1 U15700 ( .A1(n12621), .A2(n12620), .ZN(n19283) );
  AOI21_X1 U15701 ( .B1(n19283), .B2(n10861), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16468) );
  NAND2_X1 U15702 ( .A1(n12843), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12622) );
  OR2_X1 U15703 ( .A1(n14874), .A2(n12622), .ZN(n16482) );
  AND2_X1 U15704 ( .A1(n12843), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12623) );
  NAND2_X1 U15705 ( .A1(n14883), .A2(n12623), .ZN(n15631) );
  NAND2_X1 U15706 ( .A1(n16482), .A2(n15631), .ZN(n16466) );
  INV_X1 U15707 ( .A(n19283), .ZN(n12625) );
  NAND2_X1 U15708 ( .A1(n12843), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12624) );
  NOR2_X1 U15709 ( .A1(n12625), .A2(n12624), .ZN(n16467) );
  NOR2_X1 U15710 ( .A1(n16466), .A2(n16467), .ZN(n12626) );
  NAND3_X1 U15711 ( .A1(n12727), .A2(n12627), .A3(P2_EBX_REG_12__SCAN_IN), 
        .ZN(n12628) );
  NAND2_X1 U15712 ( .A1(n12649), .A2(n12628), .ZN(n19268) );
  NAND2_X1 U15713 ( .A1(n12843), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12629) );
  NOR2_X1 U15714 ( .A1(n19268), .A2(n12629), .ZN(n15618) );
  INV_X1 U15715 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n14844) );
  NOR2_X1 U15716 ( .A1(n10508), .A2(n14844), .ZN(n12630) );
  AND2_X1 U15717 ( .A1(n12631), .A2(n12630), .ZN(n12632) );
  OR2_X1 U15718 ( .A1(n12633), .A2(n12632), .ZN(n12668) );
  OAI21_X1 U15719 ( .B1(n12668), .B2(n12495), .A(n12634), .ZN(n15327) );
  NOR2_X1 U15720 ( .A1(n10508), .A2(n15072), .ZN(n12636) );
  INV_X1 U15721 ( .A(n12706), .ZN(n12635) );
  AOI21_X1 U15722 ( .B1(n12645), .B2(n12636), .A(n12635), .ZN(n12637) );
  OR2_X1 U15723 ( .A1(n12645), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12658) );
  NAND2_X1 U15724 ( .A1(n19232), .A2(n10861), .ZN(n12638) );
  XNOR2_X1 U15725 ( .A(n12638), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15373) );
  NOR2_X1 U15726 ( .A1(n12656), .A2(n12639), .ZN(n12640) );
  OR2_X1 U15727 ( .A1(n12664), .A2(n12640), .ZN(n19199) );
  OAI21_X1 U15728 ( .B1(n19199), .B2(n12495), .A(n12641), .ZN(n15354) );
  OR2_X1 U15729 ( .A1(n12643), .A2(n12642), .ZN(n12644) );
  AND2_X1 U15730 ( .A1(n12645), .A2(n12644), .ZN(n19247) );
  NAND2_X1 U15731 ( .A1(n19247), .A2(n12843), .ZN(n12646) );
  NAND2_X1 U15732 ( .A1(n12646), .A2(n16505), .ZN(n16435) );
  XNOR2_X1 U15733 ( .A(n12651), .B(n9804), .ZN(n19256) );
  NAND2_X1 U15734 ( .A1(n19256), .A2(n12843), .ZN(n12647) );
  INV_X1 U15735 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15601) );
  NAND2_X1 U15736 ( .A1(n12647), .A2(n15601), .ZN(n15595) );
  NAND2_X1 U15737 ( .A1(n12649), .A2(n12648), .ZN(n12650) );
  NAND2_X1 U15738 ( .A1(n12651), .A2(n12650), .ZN(n14866) );
  INV_X1 U15739 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12652) );
  OAI21_X1 U15740 ( .B1(n14866), .B2(n12495), .A(n12652), .ZN(n16452) );
  OR2_X1 U15741 ( .A1(n19268), .A2(n12495), .ZN(n12653) );
  INV_X1 U15742 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16515) );
  NAND2_X1 U15743 ( .A1(n12653), .A2(n16515), .ZN(n15617) );
  AND4_X1 U15744 ( .A1(n16435), .A2(n15595), .A3(n16452), .A4(n15617), .ZN(
        n12662) );
  AND2_X1 U15745 ( .A1(n12659), .A2(n12654), .ZN(n12655) );
  NOR2_X1 U15746 ( .A1(n12656), .A2(n12655), .ZN(n19207) );
  NAND2_X1 U15747 ( .A1(n19207), .A2(n12843), .ZN(n12672) );
  INV_X1 U15748 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12802) );
  NAND2_X1 U15749 ( .A1(n12672), .A2(n12802), .ZN(n15363) );
  NOR2_X1 U15750 ( .A1(n10508), .A2(n10588), .ZN(n12657) );
  NAND2_X1 U15751 ( .A1(n12658), .A2(n12657), .ZN(n12660) );
  AND2_X1 U15752 ( .A1(n12660), .A2(n12659), .ZN(n19223) );
  NAND2_X1 U15753 ( .A1(n19223), .A2(n12843), .ZN(n12661) );
  INV_X1 U15754 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16426) );
  NAND2_X1 U15755 ( .A1(n12661), .A2(n16426), .ZN(n15572) );
  AND4_X1 U15756 ( .A1(n15354), .A2(n12662), .A3(n15363), .A4(n15572), .ZN(
        n12666) );
  NOR2_X1 U15757 ( .A1(n10508), .A2(n19181), .ZN(n12663) );
  XNOR2_X1 U15758 ( .A(n12664), .B(n12663), .ZN(n19184) );
  NAND2_X1 U15759 ( .A1(n19184), .A2(n10861), .ZN(n12665) );
  NAND2_X1 U15760 ( .A1(n12665), .A2(n15346), .ZN(n15342) );
  AND4_X1 U15761 ( .A1(n15327), .A2(n15373), .A3(n12666), .A4(n15342), .ZN(
        n12667) );
  NAND2_X1 U15762 ( .A1(n15328), .A2(n12667), .ZN(n12685) );
  INV_X1 U15763 ( .A(n12668), .ZN(n14849) );
  AND2_X1 U15764 ( .A1(n12843), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12669) );
  NAND2_X1 U15765 ( .A1(n14849), .A2(n12669), .ZN(n15326) );
  INV_X1 U15766 ( .A(n19199), .ZN(n12671) );
  AND2_X1 U15767 ( .A1(n12843), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12670) );
  NAND2_X1 U15768 ( .A1(n12671), .A2(n12670), .ZN(n15353) );
  INV_X1 U15769 ( .A(n12672), .ZN(n12673) );
  NAND2_X1 U15770 ( .A1(n12673), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15364) );
  NAND2_X1 U15771 ( .A1(n15353), .A2(n15364), .ZN(n15333) );
  AND2_X1 U15772 ( .A1(n12843), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12674) );
  NAND2_X1 U15773 ( .A1(n19223), .A2(n12674), .ZN(n15571) );
  AND2_X1 U15774 ( .A1(n12843), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12675) );
  NAND2_X1 U15775 ( .A1(n19247), .A2(n12675), .ZN(n16434) );
  INV_X1 U15776 ( .A(n14866), .ZN(n12677) );
  AND2_X1 U15777 ( .A1(n12843), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12676) );
  NAND2_X1 U15778 ( .A1(n12677), .A2(n12676), .ZN(n16451) );
  AND2_X1 U15779 ( .A1(n16434), .A2(n16451), .ZN(n12680) );
  AND2_X1 U15780 ( .A1(n12843), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12678) );
  NAND2_X1 U15781 ( .A1(n19256), .A2(n12678), .ZN(n15594) );
  AND2_X1 U15782 ( .A1(n12843), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12679) );
  NAND2_X1 U15783 ( .A1(n19232), .A2(n12679), .ZN(n15331) );
  NAND4_X1 U15784 ( .A1(n15571), .A2(n12680), .A3(n15594), .A4(n15331), .ZN(
        n12681) );
  NOR2_X1 U15785 ( .A1(n15333), .A2(n12681), .ZN(n12683) );
  AND2_X1 U15786 ( .A1(n12843), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12682) );
  NAND2_X1 U15787 ( .A1(n19184), .A2(n12682), .ZN(n15341) );
  AND3_X1 U15788 ( .A1(n15326), .A2(n12683), .A3(n15341), .ZN(n12684) );
  INV_X1 U15789 ( .A(n12686), .ZN(n12687) );
  NAND2_X1 U15790 ( .A1(n12688), .A2(n12687), .ZN(n12689) );
  NAND2_X1 U15791 ( .A1(n12694), .A2(n12689), .ZN(n16053) );
  OR2_X1 U15792 ( .A1(n16053), .A2(n12495), .ZN(n12690) );
  NAND2_X1 U15793 ( .A1(n12690), .A2(n15515), .ZN(n15318) );
  NAND2_X1 U15794 ( .A1(n12843), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12691) );
  OR2_X1 U15795 ( .A1(n16053), .A2(n12691), .ZN(n15317) );
  NAND2_X1 U15796 ( .A1(n12694), .A2(n12693), .ZN(n12695) );
  AND2_X1 U15797 ( .A1(n12697), .A2(n12695), .ZN(n14834) );
  NAND2_X1 U15798 ( .A1(n14834), .A2(n12843), .ZN(n12696) );
  XNOR2_X1 U15799 ( .A(n12696), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15311) );
  NAND3_X1 U15800 ( .A1(n12697), .A2(P2_EBX_REG_24__SCAN_IN), .A3(n12727), 
        .ZN(n12698) );
  NAND2_X1 U15801 ( .A1(n12698), .A2(n12706), .ZN(n12699) );
  NOR2_X1 U15802 ( .A1(n12704), .A2(n12699), .ZN(n16405) );
  NAND2_X1 U15803 ( .A1(n16405), .A2(n10861), .ZN(n15304) );
  NAND2_X1 U15804 ( .A1(n12700), .A2(n15304), .ZN(n12703) );
  NAND2_X1 U15805 ( .A1(n12727), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12705) );
  MUX2_X1 U15806 ( .A(n12705), .B(P2_EBX_REG_25__SCAN_IN), .S(n12704), .Z(
        n12707) );
  AOI21_X1 U15807 ( .B1(n16394), .B2(n10861), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15292) );
  NAND3_X1 U15808 ( .A1(n12727), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n12708), 
        .ZN(n12709) );
  AND2_X1 U15809 ( .A1(n12710), .A2(n12709), .ZN(n16383) );
  NAND2_X1 U15810 ( .A1(n16383), .A2(n10861), .ZN(n12720) );
  XNOR2_X1 U15811 ( .A(n12720), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15279) );
  INV_X1 U15812 ( .A(n12711), .ZN(n12713) );
  NAND2_X1 U15813 ( .A1(n12713), .A2(n12712), .ZN(n12714) );
  NAND2_X1 U15814 ( .A1(n12716), .A2(n12714), .ZN(n16371) );
  INV_X1 U15815 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12715) );
  NAND2_X1 U15816 ( .A1(n15453), .A2(n12715), .ZN(n12719) );
  AOI21_X1 U15817 ( .B1(n12717), .B2(n12716), .A(n12725), .ZN(n16360) );
  NAND2_X1 U15818 ( .A1(n16360), .A2(n10861), .ZN(n15261) );
  INV_X1 U15819 ( .A(n15261), .ZN(n12718) );
  OAI21_X1 U15820 ( .B1(n15255), .B2(n12719), .A(n12718), .ZN(n12723) );
  NAND2_X1 U15821 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15430) );
  INV_X1 U15822 ( .A(n15430), .ZN(n12806) );
  INV_X1 U15823 ( .A(n12720), .ZN(n12722) );
  AND2_X1 U15824 ( .A1(n12843), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12721) );
  AOI21_X1 U15825 ( .B1(n12722), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15291), .ZN(n15258) );
  XNOR2_X1 U15826 ( .A(n12725), .B(n12724), .ZN(n12726) );
  INV_X1 U15827 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15434) );
  OAI21_X1 U15828 ( .B1(n12726), .B2(n12495), .A(n15434), .ZN(n15246) );
  INV_X1 U15829 ( .A(n12726), .ZN(n16347) );
  NAND3_X1 U15830 ( .A1(n16347), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n12843), .ZN(n15245) );
  NAND2_X1 U15831 ( .A1(n12727), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12728) );
  XNOR2_X1 U15832 ( .A(n12729), .B(n12728), .ZN(n14818) );
  AOI21_X1 U15833 ( .B1(n14818), .B2(n10861), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14087) );
  NOR2_X1 U15834 ( .A1(n14087), .A2(n9732), .ZN(n12730) );
  XNOR2_X1 U15835 ( .A(n12731), .B(n12730), .ZN(n12867) );
  OAI211_X1 U15836 ( .C1(n12734), .C2(n12733), .A(n13517), .B(n12732), .ZN(
        n12763) );
  INV_X1 U15837 ( .A(n12735), .ZN(n13515) );
  NAND3_X1 U15838 ( .A1(n12736), .A2(n13515), .A3(n19459), .ZN(n12762) );
  NAND2_X1 U15839 ( .A1(n12738), .A2(n12737), .ZN(n12739) );
  OAI21_X1 U15840 ( .B1(n12740), .B2(n12739), .A(n13562), .ZN(n12743) );
  AOI21_X1 U15841 ( .B1(n12741), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15856) );
  AOI21_X1 U15842 ( .B1(n12742), .B2(n15856), .A(P2_FLUSH_REG_SCAN_IN), .ZN(
        n16597) );
  MUX2_X1 U15843 ( .A(n12743), .B(n16597), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n20102) );
  INV_X1 U15844 ( .A(n12744), .ZN(n12750) );
  INV_X1 U15845 ( .A(n12745), .ZN(n12746) );
  OAI21_X1 U15846 ( .B1(n12748), .B2(n12747), .A(n12746), .ZN(n12749) );
  NAND2_X1 U15847 ( .A1(n12750), .A2(n12749), .ZN(n12752) );
  NAND2_X1 U15848 ( .A1(n12752), .A2(n12751), .ZN(n20101) );
  INV_X1 U15849 ( .A(n20100), .ZN(n12851) );
  OAI22_X1 U15850 ( .A1(n15751), .A2(n20102), .B1(n20101), .B2(n12851), .ZN(
        n12754) );
  INV_X1 U15851 ( .A(n20106), .ZN(n12753) );
  AND2_X1 U15852 ( .A1(n12755), .A2(n13515), .ZN(n12757) );
  AOI21_X1 U15853 ( .B1(n13562), .B2(n12757), .A(n12756), .ZN(n13511) );
  MUX2_X1 U15854 ( .A(n12755), .B(n19459), .S(n15751), .Z(n12758) );
  NAND3_X1 U15855 ( .A1(n13562), .A2(n20114), .A3(n12758), .ZN(n12759) );
  NAND2_X1 U15856 ( .A1(n13511), .A2(n12759), .ZN(n12760) );
  NOR2_X1 U15857 ( .A1(n12856), .A2(n12760), .ZN(n12761) );
  NAND3_X1 U15858 ( .A1(n12763), .A2(n12762), .A3(n12761), .ZN(n12764) );
  OR2_X1 U15859 ( .A1(n20106), .A2(n12765), .ZN(n12766) );
  INV_X1 U15860 ( .A(n12767), .ZN(n12768) );
  NAND2_X1 U15861 ( .A1(n12768), .A2(n20122), .ZN(n13535) );
  NAND2_X1 U15862 ( .A1(n13535), .A2(n12769), .ZN(n12772) );
  NOR2_X1 U15863 ( .A1(n12883), .A2(n10647), .ZN(n12770) );
  AOI21_X1 U15864 ( .B1(n12772), .B2(n12771), .A(n12770), .ZN(n12781) );
  INV_X1 U15865 ( .A(n12773), .ZN(n12774) );
  OAI21_X1 U15866 ( .B1(n12775), .B2(n12774), .A(n12883), .ZN(n12776) );
  NAND2_X1 U15867 ( .A1(n12776), .A2(n10640), .ZN(n12778) );
  MUX2_X1 U15868 ( .A(n20115), .B(n12778), .S(n12777), .Z(n12779) );
  NAND3_X1 U15869 ( .A1(n12781), .A2(n12780), .A3(n12779), .ZN(n13559) );
  INV_X1 U15870 ( .A(n12782), .ZN(n13525) );
  NOR2_X1 U15871 ( .A1(n13559), .A2(n13525), .ZN(n12783) );
  NAND2_X2 U15872 ( .A1(n13027), .A2(n15569), .ZN(n15570) );
  NAND2_X1 U15873 ( .A1(n15570), .A2(n12802), .ZN(n12789) );
  AND3_X1 U15874 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12849) );
  INV_X1 U15875 ( .A(n15570), .ZN(n16595) );
  NOR2_X1 U15876 ( .A1(n16558), .A2(n16561), .ZN(n16557) );
  INV_X1 U15877 ( .A(n16557), .ZN(n12800) );
  NAND2_X1 U15878 ( .A1(n15570), .A2(n12800), .ZN(n12786) );
  INV_X1 U15879 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13024) );
  NAND2_X1 U15880 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13023) );
  NOR2_X1 U15881 ( .A1(n13024), .A2(n13023), .ZN(n13025) );
  NAND2_X1 U15882 ( .A1(n13024), .A2(n13023), .ZN(n12784) );
  OAI211_X1 U15883 ( .C1(n15567), .C2(n13025), .A(n12784), .B(n15570), .ZN(
        n16575) );
  NOR2_X1 U15884 ( .A1(n12785), .A2(n16575), .ZN(n15677) );
  NOR2_X1 U15885 ( .A1(n15676), .A2(n15660), .ZN(n15656) );
  NAND2_X1 U15886 ( .A1(n15677), .A2(n15656), .ZN(n12798) );
  NOR2_X1 U15887 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12798), .ZN(
        n15652) );
  NAND2_X1 U15888 ( .A1(n12853), .A2(n19300), .ZN(n16586) );
  OAI211_X1 U15889 ( .C1(n15569), .C2(n13025), .A(n13037), .B(n16586), .ZN(
        n16572) );
  AOI21_X1 U15890 ( .B1(n12785), .B2(n15570), .A(n16572), .ZN(n15673) );
  OAI21_X1 U15891 ( .B1(n16595), .B2(n15656), .A(n15673), .ZN(n15647) );
  NOR2_X1 U15892 ( .A1(n16515), .A2(n12652), .ZN(n15599) );
  INV_X1 U15893 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16542) );
  NOR2_X1 U15894 ( .A1(n16545), .A2(n16542), .ZN(n16532) );
  NAND2_X1 U15895 ( .A1(n15599), .A2(n16532), .ZN(n12801) );
  INV_X1 U15896 ( .A(n12801), .ZN(n12787) );
  NAND2_X1 U15897 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n12787), .ZN(
        n12847) );
  NAND2_X1 U15898 ( .A1(n12788), .A2(n16526), .ZN(n16506) );
  OAI21_X1 U15899 ( .B1(n12849), .B2(n16595), .A(n16506), .ZN(n15559) );
  AND2_X1 U15900 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15524) );
  INV_X1 U15901 ( .A(n15524), .ZN(n15536) );
  NAND2_X1 U15902 ( .A1(n15570), .A2(n15536), .ZN(n12790) );
  NAND2_X1 U15903 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15500) );
  NAND2_X1 U15904 ( .A1(n15570), .A2(n15500), .ZN(n12791) );
  NAND2_X1 U15905 ( .A1(n15570), .A2(n10218), .ZN(n12792) );
  AND2_X1 U15906 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12850) );
  INV_X1 U15907 ( .A(n12850), .ZN(n12805) );
  NAND2_X1 U15908 ( .A1(n12805), .A2(n16526), .ZN(n12793) );
  AND2_X1 U15909 ( .A1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12794) );
  NAND2_X1 U15910 ( .A1(n12806), .A2(n12794), .ZN(n14104) );
  AND2_X1 U15911 ( .A1(n15570), .A2(n14104), .ZN(n12795) );
  NOR2_X1 U15912 ( .A1(n15459), .A2(n12795), .ZN(n14107) );
  INV_X1 U15913 ( .A(n14815), .ZN(n12809) );
  AOI21_X1 U15914 ( .B1(n20122), .B2(n12796), .A(n13520), .ZN(n12797) );
  NOR2_X1 U15915 ( .A1(n12800), .A2(n16556), .ZN(n15634) );
  NAND2_X1 U15916 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15634), .ZN(
        n16546) );
  NOR2_X1 U15917 ( .A1(n12801), .A2(n16546), .ZN(n15602) );
  NAND2_X1 U15918 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15602), .ZN(
        n16502) );
  NOR2_X1 U15919 ( .A1(n16502), .A2(n12802), .ZN(n12803) );
  AND2_X1 U15920 ( .A1(n15524), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12804) );
  NAND2_X1 U15921 ( .A1(n15545), .A2(n12804), .ZN(n15499) );
  NOR2_X1 U15922 ( .A1(n15499), .A2(n15500), .ZN(n15489) );
  NAND2_X1 U15923 ( .A1(n15489), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15475) );
  OR2_X2 U15924 ( .A1(n15475), .A2(n12805), .ZN(n15431) );
  NAND3_X1 U15925 ( .A1(n12806), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14092), .ZN(n12807) );
  NAND2_X1 U15926 ( .A1(n19427), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12861) );
  OAI21_X1 U15927 ( .B1(n15431), .B2(n12807), .A(n12861), .ZN(n12808) );
  AOI21_X1 U15928 ( .B1(n12809), .B2(n16582), .A(n12808), .ZN(n12810) );
  OAI21_X1 U15929 ( .B1(n14107), .B2(n14092), .A(n12810), .ZN(n12813) );
  INV_X1 U15930 ( .A(n12811), .ZN(n12812) );
  NOR2_X1 U15931 ( .A1(n12814), .A2(n16585), .ZN(n12818) );
  XNOR2_X1 U15932 ( .A(n12816), .B(n12815), .ZN(n12817) );
  NAND2_X1 U15933 ( .A1(n12818), .A2(n12817), .ZN(n12819) );
  XOR2_X1 U15934 ( .A(n12818), .B(n12817), .Z(n13003) );
  NAND2_X1 U15935 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13003), .ZN(
        n13002) );
  NAND2_X1 U15936 ( .A1(n12819), .A2(n13002), .ZN(n12822) );
  XNOR2_X1 U15937 ( .A(n13024), .B(n12822), .ZN(n12985) );
  XNOR2_X1 U15938 ( .A(n12821), .B(n12820), .ZN(n12984) );
  NAND2_X1 U15939 ( .A1(n12985), .A2(n12984), .ZN(n12824) );
  NAND2_X1 U15940 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12822), .ZN(
        n12823) );
  NAND2_X1 U15941 ( .A1(n12824), .A2(n12823), .ZN(n12825) );
  XNOR2_X1 U15942 ( .A(n12825), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13701) );
  NAND2_X1 U15943 ( .A1(n12825), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12826) );
  INV_X1 U15944 ( .A(n12827), .ZN(n12828) );
  XNOR2_X1 U15945 ( .A(n12829), .B(n12828), .ZN(n12831) );
  XNOR2_X1 U15946 ( .A(n12830), .B(n12831), .ZN(n15669) );
  INV_X1 U15947 ( .A(n12830), .ZN(n12832) );
  NAND2_X1 U15948 ( .A1(n12832), .A2(n12831), .ZN(n12833) );
  NAND2_X1 U15949 ( .A1(n12835), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15422) );
  INV_X1 U15950 ( .A(n15422), .ZN(n15419) );
  INV_X1 U15951 ( .A(n12838), .ZN(n12839) );
  NAND2_X1 U15952 ( .A1(n15419), .A2(n12839), .ZN(n12840) );
  NAND2_X1 U15953 ( .A1(n15407), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15406) );
  XNOR2_X1 U15954 ( .A(n12842), .B(n12495), .ZN(n15396) );
  OAI21_X1 U15955 ( .B1(n12842), .B2(n12495), .A(n16561), .ZN(n12845) );
  NAND2_X1 U15956 ( .A1(n12843), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12844) );
  NAND2_X1 U15957 ( .A1(n12845), .A2(n12846), .ZN(n15382) );
  INV_X1 U15958 ( .A(n12849), .ZN(n15556) );
  NAND2_X1 U15959 ( .A1(n9752), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15345) );
  OR2_X1 U15960 ( .A1(n20106), .A2(n12851), .ZN(n12852) );
  OAI211_X1 U15961 ( .C1(n12867), .C2(n16570), .A(n12854), .B(n9730), .ZN(
        P2_U3016) );
  NOR2_X1 U15962 ( .A1(n20115), .A2(n16605), .ZN(n12855) );
  INV_X1 U15963 ( .A(n12913), .ZN(n12864) );
  OR2_X1 U15964 ( .A1(n20068), .A2(n20059), .ZN(n20092) );
  NAND2_X1 U15965 ( .A1(n20092), .A2(n19974), .ZN(n12857) );
  AND2_X1 U15966 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20080) );
  NAND2_X1 U15967 ( .A1(n19726), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12858) );
  NAND2_X1 U15968 ( .A1(n12859), .A2(n12858), .ZN(n12965) );
  INV_X1 U15969 ( .A(n14808), .ZN(n12860) );
  NAND2_X1 U15970 ( .A1(n19426), .A2(n12860), .ZN(n12862) );
  OAI211_X1 U15971 ( .C1(n19438), .C2(n10158), .A(n12862), .B(n12861), .ZN(
        n12863) );
  OAI211_X1 U15972 ( .C1(n12867), .C2(n19431), .A(n12866), .B(n9729), .ZN(
        P2_U2984) );
  OAI21_X1 U15973 ( .B1(n12001), .B2(n12868), .A(n14199), .ZN(n14444) );
  INV_X1 U15974 ( .A(n14444), .ZN(n12877) );
  NOR3_X1 U15975 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12869) );
  NAND4_X1 U15976 ( .A1(n16174), .A2(n12869), .A3(n14539), .A4(n11915), .ZN(
        n12872) );
  NAND3_X1 U15977 ( .A1(n16173), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12871) );
  MUX2_X1 U15978 ( .A(n12872), .B(n12871), .S(n12870), .Z(n12873) );
  INV_X1 U15979 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14160) );
  NOR2_X1 U15980 ( .A1(n16202), .A2(n14214), .ZN(n12876) );
  INV_X1 U15981 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n21005) );
  OR2_X1 U15982 ( .A1(n14779), .A2(n21005), .ZN(n14688) );
  OAI21_X1 U15983 ( .B1(n16209), .B2(n12874), .A(n14688), .ZN(n12875) );
  NOR2_X1 U15984 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12879) );
  NOR4_X1 U15985 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12878) );
  NAND4_X1 U15986 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12879), .A4(n12878), .ZN(n12882) );
  INV_X1 U15987 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n20992) );
  NOR3_X1 U15988 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_D_C_N_REG_SCAN_IN), .A3(
        n20992), .ZN(n12881) );
  NOR4_X1 U15989 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(P1_BE_N_REG_2__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n12880)
         );
  NAND4_X1 U15990 ( .A1(n14438), .A2(P1_W_R_N_REG_SCAN_IN), .A3(n12881), .A4(
        n12880), .ZN(U214) );
  NOR2_X1 U15991 ( .A1(n15707), .A2(n12882), .ZN(n16680) );
  NAND2_X1 U15992 ( .A1(n16680), .A2(U214), .ZN(U212) );
  AOI21_X1 U15993 ( .B1(n20068), .B2(n10677), .A(P2_READREQUEST_REG_SCAN_IN), 
        .ZN(n12885) );
  NAND2_X1 U15994 ( .A1(n20111), .A2(n12883), .ZN(n12884) );
  OAI21_X1 U15995 ( .B1(n20111), .B2(n12885), .A(n12884), .ZN(P2_U3612) );
  OAI21_X1 U15996 ( .B1(n15751), .B2(n20114), .A(n19153), .ZN(n12914) );
  CLKBUF_X1 U15997 ( .A(n12914), .Z(n12908) );
  AOI22_X1 U15998 ( .A1(P2_EAX_REG_19__SCAN_IN), .A2(n12949), .B1(n12908), 
        .B2(P2_UWORD_REG_3__SCAN_IN), .ZN(n12886) );
  NAND3_X1 U15999 ( .A1(n19153), .A2(n20114), .A3(n20122), .ZN(n12951) );
  AOI22_X1 U16000 ( .A1(n15709), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n15707), .ZN(n19465) );
  INV_X1 U16001 ( .A(n19465), .ZN(n15202) );
  NAND2_X1 U16002 ( .A1(n12941), .A2(n15202), .ZN(n12947) );
  NAND2_X1 U16003 ( .A1(n12886), .A2(n12947), .ZN(P2_U2955) );
  AOI22_X1 U16004 ( .A1(P2_EAX_REG_23__SCAN_IN), .A2(n12949), .B1(n12908), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n12887) );
  OAI22_X1 U16005 ( .A1(n15707), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n15709), .ZN(n19489) );
  INV_X1 U16006 ( .A(n19489), .ZN(n16416) );
  NAND2_X1 U16007 ( .A1(n12941), .A2(n16416), .ZN(n12931) );
  NAND2_X1 U16008 ( .A1(n12887), .A2(n12931), .ZN(P2_U2959) );
  AOI22_X1 U16009 ( .A1(P2_EAX_REG_21__SCAN_IN), .A2(n12949), .B1(n12908), 
        .B2(P2_UWORD_REG_5__SCAN_IN), .ZN(n12888) );
  AOI22_X1 U16010 ( .A1(n15709), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n15707), .ZN(n19474) );
  INV_X1 U16011 ( .A(n19474), .ZN(n15181) );
  NAND2_X1 U16012 ( .A1(n12941), .A2(n15181), .ZN(n12937) );
  NAND2_X1 U16013 ( .A1(n12888), .A2(n12937), .ZN(P2_U2957) );
  AOI22_X1 U16014 ( .A1(P2_EAX_REG_17__SCAN_IN), .A2(n12949), .B1(n12908), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n12889) );
  AOI22_X1 U16015 ( .A1(n15709), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n15707), .ZN(n19381) );
  INV_X1 U16016 ( .A(n19381), .ZN(n15225) );
  NAND2_X1 U16017 ( .A1(n12941), .A2(n15225), .ZN(n12939) );
  NAND2_X1 U16018 ( .A1(n12889), .A2(n12939), .ZN(P2_U2953) );
  NAND2_X1 U16019 ( .A1(n12941), .A2(n19341), .ZN(n12898) );
  NAND2_X1 U16020 ( .A1(n12908), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n12890) );
  OAI211_X1 U16021 ( .C1(n13011), .C2(n12367), .A(n12898), .B(n12890), .ZN(
        P2_U2966) );
  INV_X1 U16022 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19407) );
  INV_X1 U16023 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16720) );
  OR2_X1 U16024 ( .A1(n15707), .A2(n16720), .ZN(n12892) );
  NAND2_X1 U16025 ( .A1(n15707), .A2(BUF2_REG_8__SCAN_IN), .ZN(n12891) );
  NAND2_X1 U16026 ( .A1(n12892), .A2(n12891), .ZN(n19351) );
  NAND2_X1 U16027 ( .A1(n12941), .A2(n19351), .ZN(n12920) );
  NAND2_X1 U16028 ( .A1(n12914), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n12893) );
  OAI211_X1 U16029 ( .C1(n13011), .C2(n19407), .A(n12920), .B(n12893), .ZN(
        P2_U2975) );
  INV_X1 U16030 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19401) );
  INV_X1 U16031 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16714) );
  OR2_X1 U16032 ( .A1(n15707), .A2(n16714), .ZN(n12895) );
  NAND2_X1 U16033 ( .A1(n15707), .A2(BUF2_REG_11__SCAN_IN), .ZN(n12894) );
  NAND2_X1 U16034 ( .A1(n12895), .A2(n12894), .ZN(n19348) );
  NAND2_X1 U16035 ( .A1(n12941), .A2(n19348), .ZN(n12903) );
  NAND2_X1 U16036 ( .A1(n12914), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n12896) );
  OAI211_X1 U16037 ( .C1(n13011), .C2(n19401), .A(n12903), .B(n12896), .ZN(
        P2_U2978) );
  INV_X1 U16038 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19395) );
  NAND2_X1 U16039 ( .A1(n12914), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n12897) );
  OAI211_X1 U16040 ( .C1(n13011), .C2(n19395), .A(n12898), .B(n12897), .ZN(
        P2_U2981) );
  INV_X1 U16041 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19397) );
  INV_X1 U16042 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16710) );
  OR2_X1 U16043 ( .A1(n15707), .A2(n16710), .ZN(n12900) );
  NAND2_X1 U16044 ( .A1(n15707), .A2(BUF2_REG_13__SCAN_IN), .ZN(n12899) );
  NAND2_X1 U16045 ( .A1(n12900), .A2(n12899), .ZN(n19345) );
  NAND2_X1 U16046 ( .A1(n12941), .A2(n19345), .ZN(n12905) );
  NAND2_X1 U16047 ( .A1(n12914), .A2(P2_LWORD_REG_13__SCAN_IN), .ZN(n12901) );
  OAI211_X1 U16048 ( .C1(n13011), .C2(n19397), .A(n12905), .B(n12901), .ZN(
        P2_U2980) );
  INV_X1 U16049 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n13018) );
  NAND2_X1 U16050 ( .A1(n12914), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n12902) );
  OAI211_X1 U16051 ( .C1(n13011), .C2(n13018), .A(n12903), .B(n12902), .ZN(
        P2_U2963) );
  INV_X1 U16052 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n13203) );
  NAND2_X1 U16053 ( .A1(n12914), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n12904) );
  OAI211_X1 U16054 ( .C1(n13011), .C2(n13203), .A(n12905), .B(n12904), .ZN(
        P2_U2965) );
  AOI22_X1 U16055 ( .A1(n12949), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12908), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n12906) );
  AOI22_X1 U16056 ( .A1(n15709), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n15707), .ZN(n15717) );
  INV_X1 U16057 ( .A(n15717), .ZN(n15175) );
  NAND2_X1 U16058 ( .A1(n12941), .A2(n15175), .ZN(n12929) );
  NAND2_X1 U16059 ( .A1(n12906), .A2(n12929), .ZN(P2_U2958) );
  AOI22_X1 U16060 ( .A1(n12949), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n12908), 
        .B2(P2_UWORD_REG_4__SCAN_IN), .ZN(n12907) );
  AOI22_X1 U16061 ( .A1(n15709), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n15707), .ZN(n19469) );
  INV_X1 U16062 ( .A(n19469), .ZN(n15193) );
  NAND2_X1 U16063 ( .A1(n12941), .A2(n15193), .ZN(n12924) );
  NAND2_X1 U16064 ( .A1(n12907), .A2(n12924), .ZN(P2_U2956) );
  AOI22_X1 U16065 ( .A1(n12949), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n12908), 
        .B2(P2_UWORD_REG_2__SCAN_IN), .ZN(n12909) );
  AOI22_X1 U16066 ( .A1(n15709), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n15707), .ZN(n19460) );
  INV_X1 U16067 ( .A(n19460), .ZN(n15215) );
  NAND2_X1 U16068 ( .A1(n12941), .A2(n15215), .ZN(n12945) );
  NAND2_X1 U16069 ( .A1(n12909), .A2(n12945), .ZN(P2_U2954) );
  INV_X1 U16070 ( .A(n12910), .ZN(n12911) );
  NOR3_X1 U16071 ( .A1(n12912), .A2(n12911), .A3(n13515), .ZN(n13569) );
  NOR2_X1 U16072 ( .A1(n13569), .A2(n16605), .ZN(n20108) );
  INV_X1 U16073 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n16120) );
  OAI21_X1 U16074 ( .B1(n20108), .B2(n16120), .A(n12913), .ZN(P2_U2819) );
  AOI22_X1 U16075 ( .A1(P2_EAX_REG_26__SCAN_IN), .A2(n12949), .B1(n12908), 
        .B2(P2_UWORD_REG_10__SCAN_IN), .ZN(n12917) );
  INV_X1 U16076 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16716) );
  OR2_X1 U16077 ( .A1(n15707), .A2(n16716), .ZN(n12916) );
  NAND2_X1 U16078 ( .A1(n15707), .A2(BUF2_REG_10__SCAN_IN), .ZN(n12915) );
  NAND2_X1 U16079 ( .A1(n12916), .A2(n12915), .ZN(n15151) );
  NAND2_X1 U16080 ( .A1(n12941), .A2(n15151), .ZN(n12933) );
  NAND2_X1 U16081 ( .A1(n12917), .A2(n12933), .ZN(P2_U2962) );
  AOI22_X1 U16082 ( .A1(P2_EAX_REG_28__SCAN_IN), .A2(n12949), .B1(n12908), 
        .B2(P2_UWORD_REG_12__SCAN_IN), .ZN(n12919) );
  AOI22_X1 U16083 ( .A1(n15709), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n15707), .ZN(n15133) );
  INV_X1 U16084 ( .A(n15133), .ZN(n12918) );
  NAND2_X1 U16085 ( .A1(n12941), .A2(n12918), .ZN(n12922) );
  NAND2_X1 U16086 ( .A1(n12919), .A2(n12922), .ZN(P2_U2964) );
  AOI22_X1 U16087 ( .A1(P2_EAX_REG_24__SCAN_IN), .A2(n12949), .B1(n12908), 
        .B2(P2_UWORD_REG_8__SCAN_IN), .ZN(n12921) );
  NAND2_X1 U16088 ( .A1(n12921), .A2(n12920), .ZN(P2_U2960) );
  AOI22_X1 U16089 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n12949), .B1(n12908), 
        .B2(P2_LWORD_REG_12__SCAN_IN), .ZN(n12923) );
  NAND2_X1 U16090 ( .A1(n12923), .A2(n12922), .ZN(P2_U2979) );
  AOI22_X1 U16091 ( .A1(n12949), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n12914), .B2(
        P2_LWORD_REG_4__SCAN_IN), .ZN(n12925) );
  NAND2_X1 U16092 ( .A1(n12925), .A2(n12924), .ZN(P2_U2971) );
  AOI22_X1 U16093 ( .A1(P2_EAX_REG_25__SCAN_IN), .A2(n12949), .B1(n12908), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n12928) );
  INV_X1 U16094 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16718) );
  OR2_X1 U16095 ( .A1(n15707), .A2(n16718), .ZN(n12927) );
  NAND2_X1 U16096 ( .A1(n15707), .A2(BUF2_REG_9__SCAN_IN), .ZN(n12926) );
  NAND2_X1 U16097 ( .A1(n12927), .A2(n12926), .ZN(n15161) );
  NAND2_X1 U16098 ( .A1(n12941), .A2(n15161), .ZN(n12935) );
  NAND2_X1 U16099 ( .A1(n12928), .A2(n12935), .ZN(P2_U2961) );
  AOI22_X1 U16100 ( .A1(n12949), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n12914), .B2(
        P2_LWORD_REG_6__SCAN_IN), .ZN(n12930) );
  NAND2_X1 U16101 ( .A1(n12930), .A2(n12929), .ZN(P2_U2973) );
  AOI22_X1 U16102 ( .A1(n12949), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n12914), .B2(
        P2_LWORD_REG_7__SCAN_IN), .ZN(n12932) );
  NAND2_X1 U16103 ( .A1(n12932), .A2(n12931), .ZN(P2_U2974) );
  AOI22_X1 U16104 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n12949), .B1(n12908), 
        .B2(P2_LWORD_REG_10__SCAN_IN), .ZN(n12934) );
  NAND2_X1 U16105 ( .A1(n12934), .A2(n12933), .ZN(P2_U2977) );
  AOI22_X1 U16106 ( .A1(P2_EAX_REG_9__SCAN_IN), .A2(n12949), .B1(n12908), .B2(
        P2_LWORD_REG_9__SCAN_IN), .ZN(n12936) );
  NAND2_X1 U16107 ( .A1(n12936), .A2(n12935), .ZN(P2_U2976) );
  AOI22_X1 U16108 ( .A1(n12949), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n12908), .B2(
        P2_LWORD_REG_5__SCAN_IN), .ZN(n12938) );
  NAND2_X1 U16109 ( .A1(n12938), .A2(n12937), .ZN(P2_U2972) );
  AOI22_X1 U16110 ( .A1(n12949), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12908), .B2(
        P2_LWORD_REG_1__SCAN_IN), .ZN(n12940) );
  NAND2_X1 U16111 ( .A1(n12940), .A2(n12939), .ZN(P2_U2968) );
  AOI22_X1 U16112 ( .A1(n12949), .A2(P2_EAX_REG_0__SCAN_IN), .B1(n12908), .B2(
        P2_LWORD_REG_0__SCAN_IN), .ZN(n12942) );
  AOI22_X1 U16113 ( .A1(n15709), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n15707), .ZN(n19390) );
  INV_X1 U16114 ( .A(n19390), .ZN(n15234) );
  NAND2_X1 U16115 ( .A1(n12941), .A2(n15234), .ZN(n12943) );
  NAND2_X1 U16116 ( .A1(n12942), .A2(n12943), .ZN(P2_U2967) );
  AOI22_X1 U16117 ( .A1(n12949), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n12908), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n12944) );
  NAND2_X1 U16118 ( .A1(n12944), .A2(n12943), .ZN(P2_U2952) );
  AOI22_X1 U16119 ( .A1(n12949), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n12908), .B2(
        P2_LWORD_REG_2__SCAN_IN), .ZN(n12946) );
  NAND2_X1 U16120 ( .A1(n12946), .A2(n12945), .ZN(P2_U2969) );
  AOI22_X1 U16121 ( .A1(n12949), .A2(P2_EAX_REG_3__SCAN_IN), .B1(n12908), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n12948) );
  NAND2_X1 U16122 ( .A1(n12948), .A2(n12947), .ZN(P2_U2970) );
  AOI22_X1 U16123 ( .A1(n15709), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n15707), .ZN(n15243) );
  AOI22_X1 U16124 ( .A1(n12949), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n12914), 
        .B2(P2_LWORD_REG_15__SCAN_IN), .ZN(n12950) );
  OAI21_X1 U16125 ( .B1(n15243), .B2(n12951), .A(n12950), .ZN(P2_U2982) );
  INV_X1 U16126 ( .A(n12974), .ZN(n12953) );
  INV_X1 U16127 ( .A(n12959), .ZN(n12956) );
  AND2_X1 U16128 ( .A1(n13219), .A2(n12954), .ZN(n12955) );
  AOI21_X1 U16129 ( .B1(n12956), .B2(n12373), .A(n12955), .ZN(n12970) );
  AND2_X1 U16130 ( .A1(n12970), .A2(n9937), .ZN(n12958) );
  INV_X1 U16131 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n21031) );
  NOR2_X1 U16132 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20678), .ZN(n12992) );
  NAND2_X1 U16133 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n12992), .ZN(n12957) );
  OAI21_X1 U16134 ( .B1(n12958), .B2(n21031), .A(n12957), .ZN(P1_U2803) );
  NAND2_X1 U16135 ( .A1(n12959), .A2(n9937), .ZN(n12991) );
  INV_X1 U16136 ( .A(n12991), .ZN(n12960) );
  INV_X1 U16137 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n21033) );
  INV_X1 U16138 ( .A(n12992), .ZN(n13769) );
  OAI211_X1 U16139 ( .C1(n12960), .C2(n21033), .A(n13769), .B(n13109), .ZN(
        P1_U2801) );
  INV_X1 U16140 ( .A(n12961), .ZN(n19323) );
  NOR2_X1 U16141 ( .A1(n19323), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12962) );
  NOR2_X1 U16142 ( .A1(n12962), .A2(n13006), .ZN(n16583) );
  AND2_X1 U16143 ( .A1(n19427), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n16590) );
  XNOR2_X1 U16144 ( .A(n12963), .B(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16588) );
  NOR2_X1 U16145 ( .A1(n19429), .A2(n16588), .ZN(n12964) );
  AOI211_X1 U16146 ( .C1(n16495), .C2(n16583), .A(n16590), .B(n12964), .ZN(
        n12967) );
  OAI21_X1 U16147 ( .B1(n16477), .B2(n12965), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12966) );
  OAI211_X1 U16148 ( .C1(n16433), .C2(n19322), .A(n12967), .B(n12966), .ZN(
        P2_U3014) );
  NAND2_X1 U16149 ( .A1(n12968), .A2(n20129), .ZN(n16112) );
  INV_X1 U16150 ( .A(n16112), .ZN(n13657) );
  OR3_X1 U16151 ( .A1(n14140), .A2(n13649), .A3(n13657), .ZN(n20843) );
  NAND2_X1 U16152 ( .A1(n20843), .A2(n20850), .ZN(n12969) );
  NAND2_X1 U16153 ( .A1(n12970), .A2(n12969), .ZN(n16079) );
  AND2_X1 U16154 ( .A1(n16079), .A2(n9937), .ZN(n20136) );
  INV_X1 U16155 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n21039) );
  INV_X1 U16156 ( .A(n12971), .ZN(n16076) );
  NAND3_X1 U16157 ( .A1(n16076), .A2(n12373), .A3(n13227), .ZN(n12977) );
  NOR2_X1 U16158 ( .A1(n14163), .A2(n12972), .ZN(n12973) );
  INV_X1 U16159 ( .A(n13231), .ZN(n13084) );
  NAND2_X1 U16160 ( .A1(n12952), .A2(n12974), .ZN(n12975) );
  OAI21_X1 U16161 ( .B1(n13219), .B2(n13084), .A(n12975), .ZN(n12976) );
  AOI21_X1 U16162 ( .B1(n12977), .B2(n13219), .A(n12976), .ZN(n16077) );
  INV_X1 U16163 ( .A(n16077), .ZN(n12978) );
  NAND2_X1 U16164 ( .A1(n20136), .A2(n12978), .ZN(n12979) );
  OAI21_X1 U16165 ( .B1(n20136), .B2(n21039), .A(n12979), .ZN(P1_U3484) );
  INV_X1 U16166 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20000) );
  OAI22_X1 U16167 ( .A1(n14943), .A2(n19438), .B1(n20000), .B2(n19300), .ZN(
        n12989) );
  NOR2_X1 U16168 ( .A1(n12982), .A2(n12981), .ZN(n13038) );
  INV_X1 U16169 ( .A(n12983), .ZN(n13039) );
  NOR3_X1 U16170 ( .A1(n19431), .A2(n13038), .A3(n13039), .ZN(n12988) );
  INV_X1 U16171 ( .A(n14941), .ZN(n12986) );
  XNOR2_X1 U16172 ( .A(n12985), .B(n12984), .ZN(n13028) );
  OAI22_X1 U16173 ( .A1(n16491), .A2(n12986), .B1(n19429), .B2(n13028), .ZN(
        n12987) );
  NOR3_X1 U16174 ( .A1(n12989), .A2(n12988), .A3(n12987), .ZN(n12990) );
  OAI21_X1 U16175 ( .B1(n12429), .B2(n16433), .A(n12990), .ZN(P2_U3012) );
  INV_X1 U16176 ( .A(n20848), .ZN(n12994) );
  OAI21_X1 U16177 ( .B1(n12992), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n12994), 
        .ZN(n12993) );
  OAI21_X1 U16178 ( .B1(n12995), .B2(n12994), .A(n12993), .ZN(P1_U3487) );
  OAI21_X1 U16179 ( .B1(n15751), .B2(n12996), .A(n20089), .ZN(n12998) );
  NOR2_X1 U16180 ( .A1(n12998), .A2(n12997), .ZN(n12999) );
  MUX2_X1 U16181 ( .A(n13000), .B(n19322), .S(n15116), .Z(n13001) );
  OAI21_X1 U16182 ( .B1(n15723), .B2(n15106), .A(n13001), .ZN(P2_U2887) );
  INV_X1 U16183 ( .A(n13059), .ZN(n14958) );
  OAI21_X1 U16184 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13003), .A(
        n13002), .ZN(n13061) );
  AND2_X1 U16185 ( .A1(n19427), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n13065) );
  INV_X1 U16186 ( .A(n13065), .ZN(n13004) );
  OAI21_X1 U16187 ( .B1(n19429), .B2(n13061), .A(n13004), .ZN(n13008) );
  XNOR2_X1 U16188 ( .A(n14952), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13005) );
  XNOR2_X1 U16189 ( .A(n13006), .B(n13005), .ZN(n13062) );
  OAI22_X1 U16190 ( .A1(n16491), .A2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n13062), .B2(n19431), .ZN(n13007) );
  AOI211_X1 U16191 ( .C1(n16477), .C2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13008), .B(n13007), .ZN(n13009) );
  OAI21_X1 U16192 ( .B1(n14958), .B2(n16433), .A(n13009), .ZN(P2_U3013) );
  INV_X1 U16193 ( .A(n12340), .ZN(n14916) );
  NAND2_X1 U16194 ( .A1(n14916), .A2(n13010), .ZN(n13012) );
  OAI21_X1 U16195 ( .B1(n13517), .B2(n13012), .A(n13011), .ZN(n13013) );
  INV_X1 U16196 ( .A(n13583), .ZN(n16596) );
  NOR2_X1 U16197 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16596), .ZN(n13200) );
  CLKBUF_X2 U16198 ( .A(n13200), .Z(n20113) );
  NOR2_X4 U16199 ( .A1(n19391), .A2(n20113), .ZN(n19410) );
  AOI22_X1 U16200 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n19410), .B1(n20113), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13015) );
  OAI21_X1 U16201 ( .B1(n12367), .B2(n13207), .A(n13015), .ZN(P2_U2921) );
  INV_X1 U16202 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n15159) );
  AOI22_X1 U16203 ( .A1(n13200), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13016) );
  OAI21_X1 U16204 ( .B1(n15159), .B2(n13207), .A(n13016), .ZN(P2_U2926) );
  AOI22_X1 U16205 ( .A1(n13200), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13017) );
  OAI21_X1 U16206 ( .B1(n13018), .B2(n13207), .A(n13017), .ZN(P2_U2924) );
  INV_X1 U16207 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n15132) );
  AOI22_X1 U16208 ( .A1(n20113), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13019) );
  OAI21_X1 U16209 ( .B1(n15132), .B2(n13207), .A(n13019), .ZN(P2_U2923) );
  NAND2_X1 U16210 ( .A1(n13163), .A2(n13482), .ZN(n13241) );
  INV_X1 U16211 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14495) );
  NAND2_X1 U16212 ( .A1(n13163), .A2(n9666), .ZN(n13164) );
  INV_X1 U16213 ( .A(DATAI_15_), .ZN(n13022) );
  INV_X1 U16214 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13021) );
  MUX2_X1 U16215 ( .A(n13022), .B(n13021), .S(n14438), .Z(n14496) );
  INV_X1 U16216 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20219) );
  OAI222_X1 U16217 ( .A1(n13241), .A2(n14495), .B1(n13164), .B2(n14496), .C1(
        n13163), .C2(n20219), .ZN(P1_U2967) );
  INV_X1 U16218 ( .A(n15569), .ZN(n13032) );
  INV_X1 U16219 ( .A(n13023), .ZN(n13060) );
  OAI22_X1 U16220 ( .A1(n13024), .A2(n13060), .B1(n13025), .B2(n13023), .ZN(
        n13031) );
  NOR2_X1 U16221 ( .A1(n16586), .A2(n13024), .ZN(n13030) );
  INV_X1 U16222 ( .A(n13025), .ZN(n13026) );
  OAI22_X1 U16223 ( .A1(n16587), .A2(n13028), .B1(n13027), .B2(n13026), .ZN(
        n13029) );
  AOI211_X1 U16224 ( .C1(n13032), .C2(n13031), .A(n13030), .B(n13029), .ZN(
        n13043) );
  OR2_X1 U16225 ( .A1(n13034), .A2(n13033), .ZN(n13036) );
  NAND2_X1 U16226 ( .A1(n13036), .A2(n13035), .ZN(n20077) );
  OAI21_X1 U16227 ( .B1(n19300), .B2(n20000), .A(n13037), .ZN(n13041) );
  NOR3_X1 U16228 ( .A1(n16570), .A2(n13039), .A3(n13038), .ZN(n13040) );
  AOI211_X1 U16229 ( .C1(n16582), .C2(n20077), .A(n13041), .B(n13040), .ZN(
        n13042) );
  OAI211_X1 U16230 ( .C1(n12429), .C2(n16574), .A(n13043), .B(n13042), .ZN(
        P2_U3044) );
  MUX2_X1 U16231 ( .A(n14953), .B(n14958), .S(n15116), .Z(n13047) );
  OAI21_X1 U16232 ( .B1(n15724), .B2(n15106), .A(n13047), .ZN(P2_U2886) );
  NOR2_X1 U16233 ( .A1(n13049), .A2(n13048), .ZN(n13050) );
  OR2_X1 U16234 ( .A1(n13051), .A2(n13050), .ZN(n19319) );
  INV_X1 U16235 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19412) );
  INV_X1 U16236 ( .A(n16417), .ZN(n15134) );
  OAI222_X1 U16237 ( .A1(n19319), .A2(n19355), .B1(n19357), .B2(n19412), .C1(
        n19389), .C2(n15717), .ZN(P2_U2913) );
  INV_X1 U16238 ( .A(n13054), .ZN(n13056) );
  NAND2_X1 U16239 ( .A1(n13056), .A2(n13055), .ZN(n13057) );
  NAND2_X1 U16240 ( .A1(n13053), .A2(n13057), .ZN(n20086) );
  INV_X1 U16241 ( .A(n20086), .ZN(n13498) );
  INV_X1 U16242 ( .A(n16586), .ZN(n13058) );
  AOI22_X1 U16243 ( .A1(n13059), .A2(n16592), .B1(n13058), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13067) );
  AOI211_X1 U16244 ( .C1(n15692), .C2(n16585), .A(n13060), .B(n16595), .ZN(
        n13064) );
  OAI22_X1 U16245 ( .A1(n16570), .A2(n13062), .B1(n16587), .B2(n13061), .ZN(
        n13063) );
  NOR3_X1 U16246 ( .A1(n13065), .A2(n13064), .A3(n13063), .ZN(n13066) );
  OAI211_X1 U16247 ( .C1(n13498), .C2(n16563), .A(n13067), .B(n13066), .ZN(
        P2_U3045) );
  NAND2_X1 U16248 ( .A1(n13070), .A2(n13069), .ZN(n13094) );
  NAND2_X1 U16249 ( .A1(n13422), .A2(n13660), .ZN(n13292) );
  OAI22_X1 U16250 ( .A1(n14164), .A2(n11085), .B1(n13071), .B2(n13654), .ZN(
        n13072) );
  INV_X1 U16251 ( .A(n13072), .ZN(n13075) );
  NAND2_X1 U16252 ( .A1(n13073), .A2(n9666), .ZN(n13074) );
  AND3_X1 U16253 ( .A1(n13094), .A2(n13075), .A3(n13074), .ZN(n13077) );
  AND2_X1 U16254 ( .A1(n13077), .A2(n13076), .ZN(n13233) );
  INV_X1 U16255 ( .A(n13080), .ZN(n13081) );
  NOR2_X1 U16256 ( .A1(n13079), .A2(n13081), .ZN(n13082) );
  NAND3_X1 U16257 ( .A1(n13233), .A2(n13082), .A3(n12377), .ZN(n13326) );
  INV_X1 U16258 ( .A(n13326), .ZN(n14789) );
  OR2_X1 U16259 ( .A1(n13068), .A2(n14789), .ZN(n13091) );
  XNOR2_X1 U16260 ( .A(n14795), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13085) );
  INV_X1 U16261 ( .A(n13085), .ZN(n13092) );
  NAND2_X1 U16262 ( .A1(n13329), .A2(n13092), .ZN(n13088) );
  XNOR2_X1 U16263 ( .A(n14792), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13086) );
  NAND2_X1 U16264 ( .A1(n13084), .A2(n13227), .ZN(n13334) );
  AOI22_X1 U16265 ( .A1(n14793), .A2(n13086), .B1(n13334), .B2(n13085), .ZN(
        n13087) );
  OAI21_X1 U16266 ( .B1(n13326), .B2(n13088), .A(n13087), .ZN(n13089) );
  INV_X1 U16267 ( .A(n13089), .ZN(n13090) );
  NAND2_X1 U16268 ( .A1(n13091), .A2(n13090), .ZN(n16063) );
  NOR2_X1 U16269 ( .A1(n16345), .A2(n10128), .ZN(n14797) );
  INV_X1 U16270 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13286) );
  AOI22_X1 U16271 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n13286), .B2(n11923), .ZN(
        n14794) );
  AOI222_X1 U16272 ( .A1(n16063), .A2(n16336), .B1(n14797), .B2(n14794), .C1(
        n13092), .C2(n16095), .ZN(n13106) );
  OAI211_X1 U16273 ( .C1(n14793), .C2(n13079), .A(n20850), .B(n16087), .ZN(
        n13099) );
  NOR2_X1 U16274 ( .A1(n13654), .A2(n11141), .ZN(n13093) );
  NOR2_X1 U16275 ( .A1(n13132), .A2(n13093), .ZN(n13098) );
  NAND2_X1 U16276 ( .A1(n13095), .A2(n13094), .ZN(n13097) );
  INV_X1 U16277 ( .A(n12952), .ZN(n13096) );
  NAND2_X1 U16278 ( .A1(n13097), .A2(n13096), .ZN(n13221) );
  NAND3_X1 U16279 ( .A1(n13099), .A2(n13098), .A3(n13221), .ZN(n13100) );
  OR2_X1 U16280 ( .A1(n16067), .A2(n16100), .ZN(n13103) );
  NAND2_X1 U16281 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16341) );
  OR2_X1 U16282 ( .A1(n20846), .A2(n16341), .ZN(n16346) );
  INV_X1 U16283 ( .A(n16346), .ZN(n13356) );
  NAND2_X1 U16284 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n13356), .ZN(n13102) );
  NAND2_X1 U16285 ( .A1(n13103), .A2(n13102), .ZN(n16334) );
  AND2_X1 U16286 ( .A1(n20846), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n13104) );
  INV_X1 U16287 ( .A(n16340), .ZN(n13144) );
  NAND2_X1 U16288 ( .A1(n13144), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13105) );
  OAI21_X1 U16289 ( .B1(n13106), .B2(n13144), .A(n13105), .ZN(P1_U3472) );
  INV_X1 U16290 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13111) );
  NAND2_X1 U16291 ( .A1(n13482), .A2(n13657), .ZN(n13108) );
  NAND3_X1 U16292 ( .A1(n14793), .A2(n9937), .A3(n16087), .ZN(n13107) );
  NAND2_X1 U16293 ( .A1(n20220), .A2(n13660), .ZN(n13385) );
  INV_X2 U16294 ( .A(n20218), .ZN(n20851) );
  NOR2_X4 U16295 ( .A1(n20220), .A2(n20851), .ZN(n16114) );
  AOI22_X1 U16296 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13110) );
  OAI21_X1 U16297 ( .B1(n13111), .B2(n13385), .A(n13110), .ZN(P1_U2912) );
  AOI22_X1 U16298 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13112) );
  OAI21_X1 U16299 ( .B1(n14479), .B2(n13385), .A(n13112), .ZN(P1_U2919) );
  INV_X1 U16300 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13114) );
  AOI22_X1 U16301 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13113) );
  OAI21_X1 U16302 ( .B1(n13114), .B2(n13385), .A(n13113), .ZN(P1_U2909) );
  INV_X1 U16303 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13116) );
  AOI22_X1 U16304 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13115) );
  OAI21_X1 U16305 ( .B1(n13116), .B2(n13385), .A(n13115), .ZN(P1_U2915) );
  INV_X1 U16306 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13118) );
  AOI22_X1 U16307 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13117) );
  OAI21_X1 U16308 ( .B1(n13118), .B2(n13385), .A(n13117), .ZN(P1_U2916) );
  INV_X1 U16309 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13120) );
  AOI22_X1 U16310 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13119) );
  OAI21_X1 U16311 ( .B1(n13120), .B2(n13385), .A(n13119), .ZN(P1_U2914) );
  INV_X1 U16312 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13122) );
  AOI22_X1 U16313 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13121) );
  OAI21_X1 U16314 ( .B1(n13122), .B2(n13385), .A(n13121), .ZN(P1_U2911) );
  INV_X1 U16315 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13124) );
  AOI22_X1 U16316 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13123) );
  OAI21_X1 U16317 ( .B1(n13124), .B2(n13385), .A(n13123), .ZN(P1_U2920) );
  INV_X1 U16318 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13126) );
  AOI22_X1 U16319 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13125) );
  OAI21_X1 U16320 ( .B1(n13126), .B2(n13385), .A(n13125), .ZN(P1_U2918) );
  INV_X1 U16321 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13128) );
  AOI22_X1 U16322 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13127) );
  OAI21_X1 U16323 ( .B1(n13128), .B2(n13385), .A(n13127), .ZN(P1_U2917) );
  INV_X1 U16324 ( .A(n13292), .ZN(n13130) );
  NAND2_X1 U16325 ( .A1(n13292), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13131) );
  OAI21_X1 U16326 ( .B1(n13129), .B2(P1_EBX_REG_0__SCAN_IN), .A(n13131), .ZN(
        n13153) );
  OAI21_X1 U16327 ( .B1(n14153), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13153), .ZN(n20278) );
  INV_X1 U16328 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13827) );
  INV_X1 U16329 ( .A(n13136), .ZN(n13140) );
  INV_X1 U16330 ( .A(n13137), .ZN(n13139) );
  OAI21_X1 U16331 ( .B1(n13140), .B2(n13139), .A(n13138), .ZN(n13833) );
  INV_X2 U16332 ( .A(n20212), .ZN(n14420) );
  OAI222_X1 U16333 ( .A1(n20278), .A2(n20209), .B1(n20216), .B2(n13827), .C1(
        n13833), .C2(n14420), .ZN(P1_U2872) );
  INV_X1 U16334 ( .A(n11347), .ZN(n13364) );
  OAI22_X1 U16335 ( .A1(n13364), .A2(n14789), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14788), .ZN(n16065) );
  INV_X1 U16336 ( .A(n16095), .ZN(n14802) );
  OAI22_X1 U16337 ( .A1(n16345), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14802), .ZN(n13141) );
  AOI21_X1 U16338 ( .B1(n16065), .B2(n16336), .A(n13141), .ZN(n13145) );
  AND2_X1 U16339 ( .A1(n14793), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n16064) );
  NAND2_X1 U16340 ( .A1(n16064), .A2(n16336), .ZN(n13143) );
  NAND2_X1 U16341 ( .A1(n13144), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13142) );
  OAI211_X1 U16342 ( .C1(n13145), .C2(n13144), .A(n13143), .B(n13142), .ZN(
        P1_U3474) );
  OAI21_X1 U16343 ( .B1(n13147), .B2(n13146), .A(n13399), .ZN(n13674) );
  NAND2_X1 U16344 ( .A1(n13292), .A2(n13286), .ZN(n13149) );
  INV_X1 U16345 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13150) );
  NAND2_X1 U16346 ( .A1(n14140), .A2(n13150), .ZN(n13148) );
  NAND3_X1 U16347 ( .A1(n13149), .A2(n14166), .A3(n13148), .ZN(n13152) );
  NAND2_X1 U16348 ( .A1(n13129), .A2(n13150), .ZN(n13151) );
  NAND2_X1 U16349 ( .A1(n13152), .A2(n13151), .ZN(n13290) );
  XNOR2_X1 U16350 ( .A(n13290), .B(n13153), .ZN(n13154) );
  NAND2_X1 U16351 ( .A1(n13154), .A2(n14140), .ZN(n13291) );
  OAI21_X1 U16352 ( .B1(n13154), .B2(n14140), .A(n13291), .ZN(n13666) );
  AOI22_X1 U16353 ( .A1(n14430), .A2(n13666), .B1(n14429), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13155) );
  OAI21_X1 U16354 ( .B1(n13674), .B2(n14420), .A(n13155), .ZN(P1_U2871) );
  INV_X1 U16355 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16739) );
  NAND2_X1 U16356 ( .A1(n14438), .A2(n16739), .ZN(n13156) );
  OAI21_X1 U16357 ( .B1(n14438), .B2(DATAI_0_), .A(n13156), .ZN(n13438) );
  OR2_X1 U16358 ( .A1(n11154), .A2(n13433), .ZN(n13157) );
  INV_X1 U16359 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20247) );
  OAI222_X1 U16360 ( .A1(n13438), .A2(n14500), .B1(n14498), .B2(n20247), .C1(
        n14505), .C2(n13833), .ZN(P1_U2904) );
  MUX2_X1 U16361 ( .A(n14944), .B(n12429), .S(n15116), .Z(n13162) );
  OAI21_X1 U16362 ( .B1(n20075), .B2(n15106), .A(n13162), .ZN(P2_U2885) );
  AOI22_X1 U16363 ( .A1(n20275), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n20274), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n13167) );
  INV_X1 U16364 ( .A(DATAI_7_), .ZN(n13166) );
  NAND2_X1 U16365 ( .A1(n14438), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13165) );
  OAI21_X1 U16366 ( .B1(n14438), .B2(n13166), .A(n13165), .ZN(n14457) );
  NAND2_X1 U16367 ( .A1(n20260), .A2(n14457), .ZN(n13250) );
  NAND2_X1 U16368 ( .A1(n13167), .A2(n13250), .ZN(P1_U2959) );
  AOI22_X1 U16369 ( .A1(n20275), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20274), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n13170) );
  NAND2_X1 U16370 ( .A1(n13418), .A2(DATAI_4_), .ZN(n13169) );
  NAND2_X1 U16371 ( .A1(n14438), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13168) );
  INV_X1 U16372 ( .A(n13623), .ZN(n14468) );
  NAND2_X1 U16373 ( .A1(n20260), .A2(n14468), .ZN(n13259) );
  NAND2_X1 U16374 ( .A1(n13170), .A2(n13259), .ZN(P1_U2956) );
  AOI22_X1 U16375 ( .A1(n20275), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n20274), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n13172) );
  INV_X1 U16376 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16726) );
  NAND2_X1 U16377 ( .A1(n14438), .A2(n16726), .ZN(n13171) );
  OAI21_X1 U16378 ( .B1(n14438), .B2(DATAI_5_), .A(n13171), .ZN(n13720) );
  INV_X1 U16379 ( .A(n13720), .ZN(n14464) );
  NAND2_X1 U16380 ( .A1(n20260), .A2(n14464), .ZN(n13245) );
  NAND2_X1 U16381 ( .A1(n13172), .A2(n13245), .ZN(P1_U2957) );
  AOI22_X1 U16382 ( .A1(n20275), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n20274), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n13174) );
  INV_X1 U16383 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16732) );
  NAND2_X1 U16384 ( .A1(n14438), .A2(n16732), .ZN(n13173) );
  OAI21_X1 U16385 ( .B1(n14438), .B2(DATAI_2_), .A(n13173), .ZN(n13617) );
  INV_X1 U16386 ( .A(n13617), .ZN(n14475) );
  NAND2_X1 U16387 ( .A1(n20260), .A2(n14475), .ZN(n13261) );
  NAND2_X1 U16388 ( .A1(n13174), .A2(n13261), .ZN(P1_U2954) );
  AOI22_X1 U16389 ( .A1(n20275), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n20274), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n13177) );
  NAND2_X1 U16390 ( .A1(n13418), .A2(DATAI_3_), .ZN(n13176) );
  NAND2_X1 U16391 ( .A1(n14438), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13175) );
  AND2_X1 U16392 ( .A1(n13176), .A2(n13175), .ZN(n13423) );
  INV_X1 U16393 ( .A(n13423), .ZN(n14472) );
  NAND2_X1 U16394 ( .A1(n20260), .A2(n14472), .ZN(n13263) );
  NAND2_X1 U16395 ( .A1(n13177), .A2(n13263), .ZN(P1_U2955) );
  AOI22_X1 U16396 ( .A1(n20275), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n20274), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n13179) );
  INV_X1 U16397 ( .A(DATAI_6_), .ZN(n20960) );
  NAND2_X1 U16398 ( .A1(n14438), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13178) );
  OAI21_X1 U16399 ( .B1(n14438), .B2(n20960), .A(n13178), .ZN(n14460) );
  NAND2_X1 U16400 ( .A1(n20260), .A2(n14460), .ZN(n13252) );
  NAND2_X1 U16401 ( .A1(n13179), .A2(n13252), .ZN(P1_U2958) );
  AOI21_X1 U16402 ( .B1(n13181), .B2(n13180), .A(n9774), .ZN(n14903) );
  INV_X1 U16403 ( .A(n14903), .ZN(n15641) );
  INV_X1 U16404 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19409) );
  OAI222_X1 U16405 ( .A1(n15641), .A2(n19355), .B1(n19357), .B2(n19409), .C1(
        n19489), .C2(n19389), .ZN(P2_U2912) );
  INV_X1 U16406 ( .A(n13182), .ZN(n13184) );
  INV_X1 U16407 ( .A(n11837), .ZN(n13183) );
  AOI21_X1 U16408 ( .B1(n13184), .B2(n10128), .A(n13183), .ZN(n20286) );
  AND2_X1 U16409 ( .A1(n16319), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n20284) );
  INV_X1 U16410 ( .A(n13185), .ZN(n13186) );
  INV_X1 U16411 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13828) );
  AOI21_X1 U16412 ( .B1(n16209), .B2(n13186), .A(n13828), .ZN(n13187) );
  AOI211_X1 U16413 ( .C1(n20286), .C2(n11980), .A(n20284), .B(n13187), .ZN(
        n13188) );
  OAI21_X1 U16414 ( .B1(n14551), .B2(n13833), .A(n13188), .ZN(P1_U2999) );
  INV_X1 U16415 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n15167) );
  AOI22_X1 U16416 ( .A1(n13200), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13189) );
  OAI21_X1 U16417 ( .B1(n15167), .B2(n13207), .A(n13189), .ZN(P2_U2927) );
  INV_X1 U16418 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13191) );
  AOI22_X1 U16419 ( .A1(n13200), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13190) );
  OAI21_X1 U16420 ( .B1(n13191), .B2(n13207), .A(n13190), .ZN(P2_U2931) );
  INV_X1 U16421 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13193) );
  AOI22_X1 U16422 ( .A1(n13200), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13192) );
  OAI21_X1 U16423 ( .B1(n13193), .B2(n13207), .A(n13192), .ZN(P2_U2929) );
  INV_X1 U16424 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n13195) );
  AOI22_X1 U16425 ( .A1(n13200), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13194) );
  OAI21_X1 U16426 ( .B1(n13195), .B2(n13207), .A(n13194), .ZN(P2_U2928) );
  INV_X1 U16427 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n15183) );
  AOI22_X1 U16428 ( .A1(n13200), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13196) );
  OAI21_X1 U16429 ( .B1(n15183), .B2(n13207), .A(n13196), .ZN(P2_U2930) );
  INV_X1 U16430 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n15204) );
  AOI22_X1 U16431 ( .A1(n13200), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13197) );
  OAI21_X1 U16432 ( .B1(n15204), .B2(n13207), .A(n13197), .ZN(P2_U2932) );
  INV_X1 U16433 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13199) );
  AOI22_X1 U16434 ( .A1(n13200), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13198) );
  OAI21_X1 U16435 ( .B1(n13199), .B2(n13207), .A(n13198), .ZN(P2_U2933) );
  INV_X1 U16436 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n15148) );
  AOI22_X1 U16437 ( .A1(n13200), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13201) );
  OAI21_X1 U16438 ( .B1(n15148), .B2(n13207), .A(n13201), .ZN(P2_U2925) );
  AOI22_X1 U16439 ( .A1(n20113), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13202) );
  OAI21_X1 U16440 ( .B1(n13203), .B2(n13207), .A(n13202), .ZN(P2_U2922) );
  INV_X1 U16441 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13205) );
  AOI22_X1 U16442 ( .A1(n20113), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13204) );
  OAI21_X1 U16443 ( .B1(n13205), .B2(n13207), .A(n13204), .ZN(P2_U2934) );
  INV_X1 U16444 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13208) );
  AOI22_X1 U16445 ( .A1(n20113), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13206) );
  OAI21_X1 U16446 ( .B1(n13208), .B2(n13207), .A(n13206), .ZN(P2_U2935) );
  XNOR2_X1 U16447 ( .A(n13209), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13282) );
  NAND2_X1 U16448 ( .A1(n9666), .A2(n16112), .ZN(n13211) );
  NAND2_X1 U16449 ( .A1(n13211), .A2(n13210), .ZN(n13217) );
  NOR2_X1 U16450 ( .A1(n13656), .A2(n13657), .ZN(n13213) );
  OAI21_X1 U16451 ( .B1(n13214), .B2(n13213), .A(n13212), .ZN(n13215) );
  NAND2_X1 U16452 ( .A1(n13215), .A2(n9938), .ZN(n13216) );
  MUX2_X1 U16453 ( .A(n13217), .B(n13216), .S(n13616), .Z(n13222) );
  NAND3_X1 U16454 ( .A1(n13219), .A2(n13218), .A3(n9666), .ZN(n13220) );
  NAND3_X1 U16455 ( .A1(n13222), .A2(n13221), .A3(n13220), .ZN(n13223) );
  NAND2_X1 U16456 ( .A1(n13225), .A2(n11138), .ZN(n13226) );
  NAND4_X1 U16457 ( .A1(n13224), .A2(n13227), .A3(n16076), .A4(n13226), .ZN(
        n13228) );
  OR2_X1 U16458 ( .A1(n12373), .A2(n9666), .ZN(n16091) );
  NAND2_X1 U16459 ( .A1(n13225), .A2(n13622), .ZN(n13229) );
  NAND2_X1 U16460 ( .A1(n16091), .A2(n13229), .ZN(n13230) );
  INV_X1 U16461 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20832) );
  OR2_X1 U16462 ( .A1(n14779), .A2(n20832), .ZN(n13277) );
  NOR2_X1 U16463 ( .A1(n14715), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n20283) );
  NAND2_X1 U16464 ( .A1(n13233), .A2(n13232), .ZN(n13234) );
  NAND2_X1 U16465 ( .A1(n13238), .A2(n13234), .ZN(n14643) );
  OR2_X1 U16466 ( .A1(n14643), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n20279) );
  NOR2_X1 U16467 ( .A1(n16319), .A2(n13238), .ZN(n20289) );
  INV_X1 U16468 ( .A(n20289), .ZN(n13235) );
  OAI21_X1 U16469 ( .B1(n20283), .B2(n14652), .A(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13236) );
  NAND2_X1 U16470 ( .A1(n13277), .A2(n13236), .ZN(n13237) );
  AOI21_X1 U16471 ( .B1(n20282), .B2(n13666), .A(n13237), .ZN(n13240) );
  NAND2_X1 U16472 ( .A1(n20287), .A2(n10128), .ZN(n13285) );
  NAND3_X1 U16473 ( .A1(n16287), .A2(n13286), .A3(n13285), .ZN(n13239) );
  OAI211_X1 U16474 ( .C1(n13282), .C2(n16260), .A(n13240), .B(n13239), .ZN(
        P1_U3030) );
  INV_X2 U16475 ( .A(n13241), .ZN(n20275) );
  AOI22_X1 U16476 ( .A1(n20275), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n20274), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n13244) );
  INV_X1 U16477 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16734) );
  NAND2_X1 U16478 ( .A1(n14438), .A2(n16734), .ZN(n13242) );
  OAI21_X1 U16479 ( .B1(n14438), .B2(DATAI_1_), .A(n13242), .ZN(n14480) );
  INV_X1 U16480 ( .A(n14480), .ZN(n13243) );
  NAND2_X1 U16481 ( .A1(n20260), .A2(n13243), .ZN(n13248) );
  NAND2_X1 U16482 ( .A1(n13244), .A2(n13248), .ZN(P1_U2953) );
  AOI22_X1 U16483 ( .A1(n20275), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n20274), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n13246) );
  NAND2_X1 U16484 ( .A1(n13246), .A2(n13245), .ZN(P1_U2942) );
  AOI22_X1 U16485 ( .A1(n20275), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n20274), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13247) );
  INV_X1 U16486 ( .A(n13438), .ZN(n14489) );
  NAND2_X1 U16487 ( .A1(n20260), .A2(n14489), .ZN(n13257) );
  NAND2_X1 U16488 ( .A1(n13247), .A2(n13257), .ZN(P1_U2937) );
  AOI22_X1 U16489 ( .A1(n20275), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n20274), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13249) );
  NAND2_X1 U16490 ( .A1(n13249), .A2(n13248), .ZN(P1_U2938) );
  AOI22_X1 U16491 ( .A1(n20275), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n20274), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13251) );
  NAND2_X1 U16492 ( .A1(n13251), .A2(n13250), .ZN(P1_U2944) );
  AOI22_X1 U16493 ( .A1(n20275), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n20274), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n13253) );
  NAND2_X1 U16494 ( .A1(n13253), .A2(n13252), .ZN(P1_U2943) );
  AOI22_X1 U16495 ( .A1(n20275), .A2(P1_EAX_REG_26__SCAN_IN), .B1(n20274), 
        .B2(P1_UWORD_REG_10__SCAN_IN), .ZN(n13256) );
  INV_X1 U16496 ( .A(DATAI_10_), .ZN(n13255) );
  NAND2_X1 U16497 ( .A1(n14438), .A2(BUF1_REG_10__SCAN_IN), .ZN(n13254) );
  OAI21_X1 U16498 ( .B1(n14438), .B2(n13255), .A(n13254), .ZN(n14448) );
  NAND2_X1 U16499 ( .A1(n20260), .A2(n14448), .ZN(n20266) );
  NAND2_X1 U16500 ( .A1(n13256), .A2(n20266), .ZN(P1_U2947) );
  AOI22_X1 U16501 ( .A1(n20275), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n20274), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n13258) );
  NAND2_X1 U16502 ( .A1(n13258), .A2(n13257), .ZN(P1_U2952) );
  AOI22_X1 U16503 ( .A1(n20275), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n20274), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13260) );
  NAND2_X1 U16504 ( .A1(n13260), .A2(n13259), .ZN(P1_U2941) );
  AOI22_X1 U16505 ( .A1(n20275), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n20274), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n13262) );
  NAND2_X1 U16506 ( .A1(n13262), .A2(n13261), .ZN(P1_U2939) );
  AOI22_X1 U16507 ( .A1(n20275), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n20274), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13264) );
  NAND2_X1 U16508 ( .A1(n13264), .A2(n13263), .ZN(P1_U2940) );
  INV_X1 U16509 ( .A(n19727), .ZN(n20070) );
  MUX2_X1 U16510 ( .A(P2_EBX_REG_3__SCAN_IN), .B(n13270), .S(n15116), .Z(
        n13271) );
  AOI21_X1 U16511 ( .B1(n20070), .B2(n15109), .A(n13271), .ZN(n13272) );
  INV_X1 U16512 ( .A(n13272), .ZN(P2_U2884) );
  NAND2_X1 U16513 ( .A1(n13273), .A2(n16559), .ZN(n13275) );
  NAND2_X1 U16514 ( .A1(n13275), .A2(n10198), .ZN(n15627) );
  INV_X1 U16515 ( .A(n15161), .ZN(n13276) );
  INV_X1 U16516 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19405) );
  OAI222_X1 U16517 ( .A1(n15627), .A2(n19355), .B1(n13276), .B2(n19389), .C1(
        n19405), .C2(n19357), .ZN(P2_U2910) );
  INV_X1 U16518 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13280) );
  OAI21_X1 U16519 ( .B1(n16209), .B2(n13280), .A(n13277), .ZN(n13279) );
  NOR2_X1 U16520 ( .A1(n13674), .A2(n14551), .ZN(n13278) );
  AOI211_X1 U16521 ( .C1(n16204), .C2(n13280), .A(n13279), .B(n13278), .ZN(
        n13281) );
  OAI21_X1 U16522 ( .B1(n13282), .B2(n20135), .A(n13281), .ZN(P1_U2998) );
  XNOR2_X1 U16523 ( .A(n13284), .B(n13283), .ZN(n13414) );
  NAND2_X1 U16524 ( .A1(n14764), .A2(n13285), .ZN(n16308) );
  NOR2_X1 U16525 ( .A1(n13286), .A2(n16308), .ZN(n13306) );
  OAI21_X1 U16526 ( .B1(n10128), .B2(n13286), .A(n13293), .ZN(n13726) );
  INV_X1 U16527 ( .A(n13726), .ZN(n13404) );
  NOR2_X1 U16528 ( .A1(n10128), .A2(n13286), .ZN(n13287) );
  AND2_X1 U16529 ( .A1(n13287), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13288) );
  NOR2_X1 U16530 ( .A1(n13404), .A2(n13288), .ZN(n13289) );
  NOR2_X1 U16531 ( .A1(n14715), .A2(n13289), .ZN(n13305) );
  NAND2_X1 U16532 ( .A1(n13291), .A2(n13290), .ZN(n13300) );
  NAND2_X1 U16533 ( .A1(n13292), .A2(n13293), .ZN(n13295) );
  INV_X1 U16534 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13296) );
  NAND2_X1 U16535 ( .A1(n14140), .A2(n13296), .ZN(n13294) );
  NAND3_X1 U16536 ( .A1(n13295), .A2(n14166), .A3(n13294), .ZN(n13298) );
  NAND2_X1 U16537 ( .A1(n13129), .A2(n13296), .ZN(n13297) );
  AND2_X1 U16538 ( .A1(n13298), .A2(n13297), .ZN(n13299) );
  NAND2_X1 U16539 ( .A1(n20282), .A2(n13739), .ZN(n13303) );
  NAND2_X1 U16540 ( .A1(n16319), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n13409) );
  OAI21_X1 U16541 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n16284), .A(
        n14648), .ZN(n13301) );
  NAND2_X1 U16542 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13301), .ZN(
        n13302) );
  NAND3_X1 U16543 ( .A1(n13303), .A2(n13409), .A3(n13302), .ZN(n13304) );
  AOI211_X1 U16544 ( .C1(n13306), .C2(n13293), .A(n13305), .B(n13304), .ZN(
        n13307) );
  OAI21_X1 U16545 ( .B1(n16260), .B2(n13414), .A(n13307), .ZN(P1_U3029) );
  OAI21_X1 U16546 ( .B1(n13308), .B2(n13310), .A(n13309), .ZN(n19361) );
  NAND2_X1 U16547 ( .A1(n13312), .A2(n13311), .ZN(n13314) );
  INV_X1 U16548 ( .A(n13319), .ZN(n13313) );
  MUX2_X1 U16549 ( .A(P2_EBX_REG_4__SCAN_IN), .B(n19434), .S(n15116), .Z(
        n13315) );
  INV_X1 U16550 ( .A(n13315), .ZN(n13316) );
  OAI21_X1 U16551 ( .B1(n19361), .B2(n15106), .A(n13316), .ZN(P2_U2883) );
  INV_X1 U16552 ( .A(n13309), .ZN(n13318) );
  OAI211_X1 U16553 ( .C1(n13318), .C2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        n15109), .B(n13317), .ZN(n13323) );
  NOR2_X1 U16554 ( .A1(n13320), .A2(n13319), .ZN(n13321) );
  NOR2_X1 U16555 ( .A1(n13444), .A2(n13321), .ZN(n15425) );
  NAND2_X1 U16556 ( .A1(n15116), .A2(n15425), .ZN(n13322) );
  OAI211_X1 U16557 ( .C1(n15116), .C2(n10551), .A(n13323), .B(n13322), .ZN(
        P2_U2882) );
  INV_X1 U16558 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19403) );
  INV_X1 U16559 ( .A(n15151), .ZN(n13325) );
  XNOR2_X1 U16560 ( .A(n13274), .B(n13324), .ZN(n16548) );
  OAI222_X1 U16561 ( .A1(n19357), .A2(n19403), .B1(n13325), .B2(n19389), .C1(
        n16548), .C2(n19355), .ZN(P2_U2909) );
  INV_X1 U16562 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20244) );
  OAI222_X1 U16563 ( .A1(n14480), .A2(n14500), .B1(n14498), .B2(n20244), .C1(
        n14505), .C2(n13674), .ZN(P1_U2903) );
  NAND2_X1 U16564 ( .A1(n20467), .A2(n13326), .ZN(n13341) );
  NAND2_X1 U16565 ( .A1(n14795), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13327) );
  NAND2_X1 U16566 ( .A1(n13327), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13328) );
  NAND2_X1 U16567 ( .A1(n9670), .A2(n13328), .ZN(n14801) );
  AND2_X1 U16568 ( .A1(n13329), .A2(n14801), .ZN(n13339) );
  MUX2_X1 U16569 ( .A(n13330), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n14792), .Z(n13331) );
  OAI21_X1 U16570 ( .B1(n13333), .B2(n13331), .A(n14793), .ZN(n13337) );
  MUX2_X1 U16571 ( .A(n13333), .B(n13332), .S(n14795), .Z(n13335) );
  OAI21_X1 U16572 ( .B1(n13330), .B2(n13335), .A(n13334), .ZN(n13336) );
  NAND2_X1 U16573 ( .A1(n13337), .A2(n13336), .ZN(n13338) );
  AOI21_X1 U16574 ( .B1(n14789), .B2(n13339), .A(n13338), .ZN(n13340) );
  NAND2_X1 U16575 ( .A1(n13341), .A2(n13340), .ZN(n16061) );
  AOI21_X1 U16576 ( .B1(n16061), .B2(n16063), .A(n16067), .ZN(n13343) );
  INV_X1 U16577 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n21037) );
  NAND2_X1 U16578 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21037), .ZN(n13342) );
  OAI21_X1 U16579 ( .B1(n13343), .B2(P1_STATE2_REG_1__SCAN_IN), .A(n13342), 
        .ZN(n13345) );
  INV_X1 U16580 ( .A(n16067), .ZN(n16062) );
  NAND2_X1 U16581 ( .A1(n13345), .A2(n10285), .ZN(n16083) );
  OR2_X1 U16582 ( .A1(n16083), .A2(n13346), .ZN(n13355) );
  INV_X1 U16583 ( .A(n13470), .ZN(n13424) );
  OR2_X1 U16584 ( .A1(n13347), .A2(n13424), .ZN(n13348) );
  XNOR2_X1 U16585 ( .A(n13348), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n16337) );
  NAND3_X1 U16586 ( .A1(n16337), .A2(n16335), .A3(n13349), .ZN(n13353) );
  INV_X1 U16587 ( .A(n13349), .ZN(n13351) );
  NOR2_X1 U16588 ( .A1(n16339), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n13350) );
  NAND2_X1 U16589 ( .A1(n13351), .A2(n13350), .ZN(n13352) );
  NAND2_X1 U16590 ( .A1(n13353), .A2(n13352), .ZN(n16081) );
  INV_X1 U16591 ( .A(n16081), .ZN(n13354) );
  NAND2_X1 U16592 ( .A1(n13355), .A2(n13354), .ZN(n13363) );
  OAI21_X1 U16593 ( .B1(n13363), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13356), .ZN(
        n13358) );
  NAND2_X1 U16594 ( .A1(n20753), .A2(n16345), .ZN(n20845) );
  NAND2_X1 U16595 ( .A1(n13358), .A2(n20298), .ZN(n20293) );
  NAND2_X1 U16596 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20609), .ZN(n13391) );
  INV_X1 U16597 ( .A(n13391), .ZN(n14786) );
  NOR2_X1 U16598 ( .A1(n13068), .A2(n14786), .ZN(n13361) );
  AOI21_X1 U16599 ( .B1(n9673), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20678), 
        .ZN(n20568) );
  NOR3_X1 U16600 ( .A1(n13389), .A2(n20841), .A3(n20678), .ZN(n13415) );
  MUX2_X1 U16601 ( .A(n20568), .B(n13415), .S(n11842), .Z(n13360) );
  OAI21_X1 U16602 ( .B1(n13361), .B2(n13360), .A(n20293), .ZN(n13362) );
  OAI21_X1 U16603 ( .B1(n20293), .B2(n20532), .A(n13362), .ZN(P1_U3476) );
  NOR2_X1 U16604 ( .A1(n13363), .A2(n16341), .ZN(n16098) );
  OAI22_X1 U16605 ( .A1(n13781), .A2(n20678), .B1(n13364), .B2(n14786), .ZN(
        n13365) );
  OAI21_X1 U16606 ( .B1(n16098), .B2(n13365), .A(n20293), .ZN(n13366) );
  OAI21_X1 U16607 ( .B1(n20293), .B2(n20643), .A(n13366), .ZN(P1_U3478) );
  OAI21_X1 U16608 ( .B1(n13367), .B2(n13369), .A(n13368), .ZN(n14383) );
  INV_X1 U16609 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n14371) );
  NAND2_X1 U16610 ( .A1(n14154), .A2(n14371), .ZN(n13372) );
  NAND2_X1 U16611 ( .A1(n14140), .A2(n14371), .ZN(n13370) );
  OAI211_X1 U16612 ( .C1(n13129), .C2(n13405), .A(n13370), .B(n13292), .ZN(
        n13371) );
  OAI21_X1 U16613 ( .B1(n13373), .B2(n9819), .A(n13464), .ZN(n14377) );
  INV_X1 U16614 ( .A(n14377), .ZN(n13374) );
  AOI22_X1 U16615 ( .A1(n13374), .A2(n14430), .B1(n14429), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n13375) );
  OAI21_X1 U16616 ( .B1(n14383), .B2(n14420), .A(n13375), .ZN(P1_U2869) );
  INV_X1 U16617 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13377) );
  AOI22_X1 U16618 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20851), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n16114), .ZN(n13376) );
  OAI21_X1 U16619 ( .B1(n13377), .B2(n13385), .A(n13376), .ZN(P1_U2906) );
  INV_X1 U16620 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13379) );
  AOI22_X1 U16621 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13378) );
  OAI21_X1 U16622 ( .B1(n13379), .B2(n13385), .A(n13378), .ZN(P1_U2907) );
  INV_X1 U16623 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13381) );
  AOI22_X1 U16624 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13380) );
  OAI21_X1 U16625 ( .B1(n13381), .B2(n13385), .A(n13380), .ZN(P1_U2913) );
  INV_X1 U16626 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13383) );
  AOI22_X1 U16627 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13382) );
  OAI21_X1 U16628 ( .B1(n13383), .B2(n13385), .A(n13382), .ZN(P1_U2908) );
  INV_X1 U16629 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13386) );
  AOI22_X1 U16630 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13384) );
  OAI21_X1 U16631 ( .B1(n13386), .B2(n13385), .A(n13384), .ZN(P1_U2910) );
  INV_X1 U16632 ( .A(n20293), .ZN(n13396) );
  INV_X1 U16633 ( .A(n11842), .ZN(n13388) );
  OR2_X1 U16634 ( .A1(n20648), .A2(n9673), .ZN(n20595) );
  NAND4_X1 U16635 ( .A1(n20569), .A2(n13477), .A3(n20595), .A4(
        P1_STATEBS16_REG_SCAN_IN), .ZN(n13393) );
  AOI21_X1 U16636 ( .B1(n13387), .B2(n20841), .A(n20678), .ZN(n13392) );
  AOI22_X1 U16637 ( .A1(n13393), .A2(n13392), .B1(n13391), .B2(n20467), .ZN(
        n13395) );
  NAND2_X1 U16638 ( .A1(n13396), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13394) );
  OAI21_X1 U16639 ( .B1(n13396), .B2(n13395), .A(n13394), .ZN(P1_U3475) );
  INV_X1 U16640 ( .A(n13397), .ZN(n13398) );
  AOI21_X1 U16641 ( .B1(n13400), .B2(n13399), .A(n13398), .ZN(n13738) );
  INV_X1 U16642 ( .A(n13738), .ZN(n13450) );
  AOI22_X1 U16643 ( .A1(n13739), .A2(n14430), .B1(n14429), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n13401) );
  OAI21_X1 U16644 ( .B1(n13450), .B2(n14420), .A(n13401), .ZN(P1_U2870) );
  XNOR2_X1 U16645 ( .A(n13403), .B(n13402), .ZN(n13456) );
  NAND2_X1 U16646 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13922) );
  OAI22_X1 U16647 ( .A1(n13404), .A2(n14715), .B1(n13922), .B2(n16308), .ZN(
        n13911) );
  NAND2_X1 U16648 ( .A1(n13911), .A2(n13405), .ZN(n13408) );
  NAND2_X1 U16649 ( .A1(n14764), .A2(n13922), .ZN(n13727) );
  OAI211_X1 U16650 ( .C1(n14715), .C2(n13726), .A(n14648), .B(n13727), .ZN(
        n13467) );
  INV_X1 U16651 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20771) );
  OAI22_X1 U16652 ( .A1(n16259), .A2(n14377), .B1(n20771), .B2(n14779), .ZN(
        n13406) );
  AOI21_X1 U16653 ( .B1(n13467), .B2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n13406), .ZN(n13407) );
  OAI211_X1 U16654 ( .C1(n13456), .C2(n16260), .A(n13408), .B(n13407), .ZN(
        P1_U3028) );
  NOR2_X1 U16655 ( .A1(n16202), .A2(n13742), .ZN(n13412) );
  INV_X1 U16656 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13410) );
  OAI21_X1 U16657 ( .B1(n16209), .B2(n13410), .A(n13409), .ZN(n13411) );
  AOI211_X1 U16658 ( .C1(n13738), .C2(n16205), .A(n13412), .B(n13411), .ZN(
        n13413) );
  OAI21_X1 U16659 ( .B1(n20135), .B2(n13414), .A(n13413), .ZN(P1_U2997) );
  INV_X1 U16660 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20240) );
  OAI222_X1 U16661 ( .A1(n14383), .A2(n14505), .B1(n14500), .B2(n13423), .C1(
        n14498), .C2(n20240), .ZN(P1_U2901) );
  INV_X1 U16662 ( .A(n13415), .ZN(n13416) );
  OAI21_X1 U16663 ( .B1(n13416), .B2(n20648), .A(n20673), .ZN(n13417) );
  NAND2_X1 U16664 ( .A1(n13417), .A2(n20650), .ZN(n20746) );
  INV_X1 U16665 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13432) );
  INV_X1 U16666 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n19464) );
  INV_X1 U16667 ( .A(DATAI_27_), .ZN(n20885) );
  OAI22_X2 U16668 ( .A1(n19464), .A2(n13694), .B1(n20885), .B2(n13693), .ZN(
        n20702) );
  NAND2_X1 U16669 ( .A1(n9673), .A2(n13781), .ZN(n20525) );
  AOI22_X1 U16670 ( .A1(DATAI_19_), .A2(n13686), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n13687), .ZN(n20705) );
  NOR2_X2 U16671 ( .A1(n13690), .A2(n13422), .ZN(n20701) );
  NOR2_X2 U16672 ( .A1(n13423), .A2(n20298), .ZN(n20700) );
  OR2_X1 U16673 ( .A1(n13068), .A2(n13424), .ZN(n20644) );
  NAND3_X1 U16674 ( .A1(n11347), .A2(n13425), .A3(n20596), .ZN(n13471) );
  OR2_X1 U16675 ( .A1(n20644), .A2(n13471), .ZN(n13428) );
  INV_X1 U16676 ( .A(n20673), .ZN(n13426) );
  AOI22_X1 U16677 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n13426), .B1(n20742), 
        .B2(n20596), .ZN(n13427) );
  NAND2_X1 U16678 ( .A1(n13428), .A2(n13427), .ZN(n20740) );
  AOI22_X1 U16679 ( .A1(n20701), .A2(n20742), .B1(n20700), .B2(n20740), .ZN(
        n13429) );
  OAI21_X1 U16680 ( .B1(n9829), .B2(n20295), .A(n13429), .ZN(n13430) );
  AOI21_X1 U16681 ( .B1(n20702), .B2(n20682), .A(n13430), .ZN(n13431) );
  OAI21_X1 U16682 ( .B1(n13715), .B2(n13432), .A(n13431), .ZN(P1_U3156) );
  INV_X1 U16683 ( .A(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13437) );
  INV_X1 U16684 ( .A(DATAI_31_), .ZN(n20918) );
  OAI22_X2 U16685 ( .A1(n20918), .A2(n13693), .B1(n19484), .B2(n13694), .ZN(
        n20728) );
  INV_X1 U16686 ( .A(n14457), .ZN(n13761) );
  NOR2_X2 U16687 ( .A1(n20298), .A2(n13761), .ZN(n20727) );
  NOR2_X2 U16688 ( .A1(n13690), .A2(n13433), .ZN(n20725) );
  AOI22_X1 U16689 ( .A1(n20727), .A2(n20740), .B1(n20725), .B2(n20742), .ZN(
        n13434) );
  OAI21_X1 U16690 ( .B1(n20733), .B2(n20295), .A(n13434), .ZN(n13435) );
  AOI21_X1 U16691 ( .B1(n20728), .B2(n20682), .A(n13435), .ZN(n13436) );
  OAI21_X1 U16692 ( .B1(n13715), .B2(n13437), .A(n13436), .ZN(P1_U3160) );
  INV_X1 U16693 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13442) );
  INV_X1 U16694 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16691) );
  INV_X1 U16695 ( .A(DATAI_24_), .ZN(n21008) );
  OAI22_X2 U16696 ( .A1(n16691), .A2(n13694), .B1(n21008), .B2(n13693), .ZN(
        n20688) );
  NOR2_X2 U16697 ( .A1(n13438), .A2(n20298), .ZN(n20679) );
  AOI22_X1 U16698 ( .A1(n20680), .A2(n20742), .B1(n20679), .B2(n20740), .ZN(
        n13439) );
  OAI21_X1 U16699 ( .B1(n20691), .B2(n20295), .A(n13439), .ZN(n13440) );
  AOI21_X1 U16700 ( .B1(n20688), .B2(n20682), .A(n13440), .ZN(n13441) );
  OAI21_X1 U16701 ( .B1(n13715), .B2(n13442), .A(n13441), .ZN(P1_U3153) );
  NOR2_X1 U16702 ( .A1(n13444), .A2(n13443), .ZN(n13445) );
  OR2_X1 U16703 ( .A1(n13458), .A2(n13445), .ZN(n15648) );
  INV_X1 U16704 ( .A(n13317), .ZN(n13447) );
  OAI211_X1 U16705 ( .C1(n13447), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n15109), .B(n13446), .ZN(n13449) );
  NAND2_X1 U16706 ( .A1(n15089), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n13448) );
  OAI211_X1 U16707 ( .C1(n15648), .C2(n15089), .A(n13449), .B(n13448), .ZN(
        P2_U2881) );
  INV_X1 U16708 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20242) );
  OAI222_X1 U16709 ( .A1(n13617), .A2(n14500), .B1(n14498), .B2(n20242), .C1(
        n14505), .C2(n13450), .ZN(P1_U2902) );
  INV_X1 U16710 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19399) );
  XNOR2_X1 U16711 ( .A(n16529), .B(n13451), .ZN(n19272) );
  OAI222_X1 U16712 ( .A1(n19357), .A2(n19399), .B1(n15133), .B2(n19389), .C1(
        n19272), .C2(n19355), .ZN(P2_U2907) );
  INV_X1 U16713 ( .A(n14383), .ZN(n13454) );
  AOI22_X1 U16714 ( .A1(n16194), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n16319), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n13452) );
  OAI21_X1 U16715 ( .B1(n14373), .B2(n16202), .A(n13452), .ZN(n13453) );
  AOI21_X1 U16716 ( .B1(n13454), .B2(n16205), .A(n13453), .ZN(n13455) );
  OAI21_X1 U16717 ( .B1(n20135), .B2(n13456), .A(n13455), .ZN(P1_U2996) );
  XOR2_X1 U16718 ( .A(n13446), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n13460)
         );
  OAI21_X1 U16719 ( .B1(n13458), .B2(n13457), .A(n13585), .ZN(n15640) );
  MUX2_X1 U16720 ( .A(n10585), .B(n15640), .S(n15116), .Z(n13459) );
  OAI21_X1 U16721 ( .B1(n13460), .B2(n15106), .A(n13459), .ZN(P2_U2880) );
  NAND2_X1 U16722 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13729) );
  OAI211_X1 U16723 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n13911), .B(n13729), .ZN(n13469) );
  INV_X1 U16724 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20772) );
  NOR2_X1 U16725 ( .A1(n14779), .A2(n20772), .ZN(n13607) );
  MUX2_X1 U16726 ( .A(n14188), .B(n13130), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n13463) );
  AND2_X1 U16727 ( .A1(n14163), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13462) );
  NOR2_X1 U16728 ( .A1(n13463), .A2(n13462), .ZN(n13465) );
  NOR2_X1 U16729 ( .A1(n13464), .A2(n13465), .ZN(n13724) );
  AOI21_X1 U16730 ( .B1(n13465), .B2(n13464), .A(n13724), .ZN(n13844) );
  INV_X1 U16731 ( .A(n13844), .ZN(n13677) );
  NOR2_X1 U16732 ( .A1(n16259), .A2(n13677), .ZN(n13466) );
  AOI211_X1 U16733 ( .C1(n13467), .C2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n13607), .B(n13466), .ZN(n13468) );
  OAI211_X1 U16734 ( .C1(n13611), .C2(n16260), .A(n13469), .B(n13468), .ZN(
        P1_U3027) );
  INV_X1 U16735 ( .A(n20680), .ZN(n13474) );
  OR2_X1 U16736 ( .A1(n13068), .A2(n13470), .ZN(n20413) );
  OR2_X1 U16737 ( .A1(n20413), .A2(n13471), .ZN(n13473) );
  AOI22_X1 U16738 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n13478), .B1(n13691), 
        .B2(n20596), .ZN(n13472) );
  INV_X1 U16739 ( .A(n20679), .ZN(n20613) );
  OAI22_X1 U16740 ( .A1(n13474), .A2(n13625), .B1(n13624), .B2(n20613), .ZN(
        n13475) );
  AOI21_X1 U16741 ( .B1(n13790), .B2(n20688), .A(n13475), .ZN(n13481) );
  INV_X1 U16742 ( .A(n13476), .ZN(n20647) );
  NOR2_X1 U16743 ( .A1(n13477), .A2(n20647), .ZN(n13479) );
  NAND2_X1 U16744 ( .A1(n13699), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n13480) );
  OAI211_X1 U16745 ( .C1(n20691), .C2(n13697), .A(n13481), .B(n13480), .ZN(
        P1_U3089) );
  AOI22_X1 U16746 ( .A1(DATAI_17_), .A2(n13686), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n13687), .ZN(n20695) );
  INV_X1 U16747 ( .A(DATAI_25_), .ZN(n20876) );
  INV_X1 U16748 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16689) );
  OAI22_X2 U16749 ( .A1(n20876), .A2(n13693), .B1(n16689), .B2(n13694), .ZN(
        n20692) );
  NOR2_X2 U16750 ( .A1(n13690), .A2(n13482), .ZN(n20735) );
  INV_X1 U16751 ( .A(n20735), .ZN(n13483) );
  NOR2_X2 U16752 ( .A1(n14480), .A2(n20298), .ZN(n20734) );
  INV_X1 U16753 ( .A(n20734), .ZN(n20616) );
  OAI22_X1 U16754 ( .A1(n13483), .A2(n13625), .B1(n13624), .B2(n20616), .ZN(
        n13484) );
  AOI21_X1 U16755 ( .B1(n13790), .B2(n20692), .A(n13484), .ZN(n13486) );
  NAND2_X1 U16756 ( .A1(n13699), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n13485) );
  OAI211_X1 U16757 ( .C1(n20695), .C2(n13697), .A(n13486), .B(n13485), .ZN(
        P1_U3090) );
  INV_X1 U16758 ( .A(n20701), .ZN(n13487) );
  INV_X1 U16759 ( .A(n20700), .ZN(n20622) );
  OAI22_X1 U16760 ( .A1(n13487), .A2(n13625), .B1(n13624), .B2(n20622), .ZN(
        n13488) );
  AOI21_X1 U16761 ( .B1(n13790), .B2(n20702), .A(n13488), .ZN(n13490) );
  NAND2_X1 U16762 ( .A1(n13699), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n13489) );
  OAI211_X1 U16763 ( .C1(n9829), .C2(n13697), .A(n13490), .B(n13489), .ZN(
        P1_U3092) );
  INV_X1 U16764 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19414) );
  NOR2_X1 U16765 ( .A1(n19361), .A2(n15230), .ZN(n13507) );
  NAND2_X1 U16766 ( .A1(n13492), .A2(n13491), .ZN(n13495) );
  INV_X1 U16767 ( .A(n13493), .ZN(n13494) );
  AND2_X1 U16768 ( .A1(n13495), .A2(n13494), .ZN(n20069) );
  XNOR2_X1 U16769 ( .A(n19727), .B(n20069), .ZN(n19367) );
  XNOR2_X1 U16770 ( .A(n19440), .B(n20077), .ZN(n19373) );
  XNOR2_X1 U16771 ( .A(n15724), .B(n20086), .ZN(n19377) );
  XNOR2_X1 U16772 ( .A(n13497), .B(n13496), .ZN(n19386) );
  NAND2_X1 U16773 ( .A1(n20093), .A2(n19386), .ZN(n19384) );
  AOI22_X1 U16774 ( .A1(n19377), .A2(n19384), .B1(n15724), .B2(n13498), .ZN(
        n19372) );
  OAI22_X1 U16775 ( .A1(n19373), .A2(n19372), .B1(n19440), .B2(n20077), .ZN(
        n19368) );
  NAND2_X1 U16776 ( .A1(n19367), .A2(n19368), .ZN(n19366) );
  OAI21_X1 U16777 ( .B1(n20070), .B2(n20069), .A(n19366), .ZN(n13500) );
  OAI21_X1 U16778 ( .B1(n13493), .B2(n13499), .A(n13503), .ZN(n19359) );
  NAND2_X1 U16779 ( .A1(n13500), .A2(n19359), .ZN(n19362) );
  INV_X1 U16780 ( .A(n13501), .ZN(n13502) );
  NAND2_X1 U16781 ( .A1(n13503), .A2(n13502), .ZN(n13504) );
  NAND2_X1 U16782 ( .A1(n13505), .A2(n13504), .ZN(n15662) );
  INV_X1 U16783 ( .A(n15662), .ZN(n13506) );
  AOI21_X1 U16784 ( .B1(n13507), .B2(n19362), .A(n13506), .ZN(n13508) );
  OAI222_X1 U16785 ( .A1(n19357), .A2(n19414), .B1(n19474), .B2(n19389), .C1(
        n19355), .C2(n13508), .ZN(P2_U2914) );
  NAND3_X1 U16786 ( .A1(n12755), .A2(n20100), .A3(n13509), .ZN(n13582) );
  NOR2_X1 U16787 ( .A1(n13510), .A2(n19591), .ZN(n20110) );
  NAND2_X1 U16788 ( .A1(n13512), .A2(n13511), .ZN(n13513) );
  NOR2_X1 U16789 ( .A1(n13514), .A2(n13513), .ZN(n13519) );
  NAND2_X1 U16790 ( .A1(n14916), .A2(n13515), .ZN(n13516) );
  OR2_X1 U16791 ( .A1(n13517), .A2(n13516), .ZN(n13518) );
  INV_X1 U16792 ( .A(n13559), .ZN(n13541) );
  INV_X1 U16793 ( .A(n13520), .ZN(n13567) );
  NAND2_X1 U16794 ( .A1(n13563), .A2(n13567), .ZN(n13550) );
  INV_X1 U16795 ( .A(n13521), .ZN(n13523) );
  NAND2_X1 U16796 ( .A1(n13523), .A2(n13522), .ZN(n13552) );
  NAND2_X1 U16797 ( .A1(n13524), .A2(n13552), .ZN(n13530) );
  NOR2_X1 U16798 ( .A1(n13526), .A2(n13525), .ZN(n13553) );
  INV_X1 U16799 ( .A(n12741), .ZN(n13527) );
  NAND2_X1 U16800 ( .A1(n13549), .A2(n13527), .ZN(n13554) );
  NOR2_X1 U16801 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13528) );
  OAI22_X1 U16802 ( .A1(n13553), .A2(n13530), .B1(n13554), .B2(n13528), .ZN(
        n13529) );
  AOI21_X1 U16803 ( .B1(n13550), .B2(n13530), .A(n13529), .ZN(n13531) );
  OAI21_X1 U16804 ( .B1(n12429), .B2(n13541), .A(n13531), .ZN(n15695) );
  NAND2_X1 U16805 ( .A1(n15685), .A2(n13522), .ZN(n13533) );
  OAI21_X1 U16806 ( .B1(n15695), .B2(n15685), .A(n13533), .ZN(n13576) );
  INV_X1 U16807 ( .A(n13576), .ZN(n13548) );
  NOR2_X1 U16808 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19554) );
  INV_X1 U16809 ( .A(n19554), .ZN(n19525) );
  INV_X1 U16810 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13539) );
  INV_X1 U16811 ( .A(n12409), .ZN(n13534) );
  NAND2_X1 U16812 ( .A1(n13535), .A2(n13534), .ZN(n13542) );
  INV_X1 U16813 ( .A(n13536), .ZN(n13537) );
  OAI21_X1 U16814 ( .B1(n15690), .B2(n13539), .A(n13537), .ZN(n13538) );
  AOI22_X1 U16815 ( .A1(n13539), .A2(n13549), .B1(n13542), .B2(n13538), .ZN(
        n13540) );
  OAI21_X1 U16816 ( .B1(n14958), .B2(n13541), .A(n13540), .ZN(n20060) );
  MUX2_X1 U16817 ( .A(n13542), .B(n13549), .S(n15690), .Z(n13543) );
  AOI21_X1 U16818 ( .B1(n16591), .B2(n13559), .A(n13543), .ZN(n15683) );
  NAND2_X1 U16819 ( .A1(n15683), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13544) );
  OR2_X1 U16820 ( .A1(n20060), .A2(n13544), .ZN(n13545) );
  AOI22_X1 U16821 ( .A1(n13545), .A2(n20088), .B1(n20060), .B2(n13544), .ZN(
        n13546) );
  OAI22_X1 U16822 ( .A1(n13576), .A2(n19525), .B1(n15685), .B2(n13546), .ZN(
        n13547) );
  OAI21_X1 U16823 ( .B1(n13548), .B2(n20079), .A(n13547), .ZN(n13561) );
  AOI22_X1 U16824 ( .A1(n13550), .A2(n13552), .B1(n12741), .B2(n13549), .ZN(
        n13551) );
  INV_X1 U16825 ( .A(n13551), .ZN(n13557) );
  AND2_X1 U16826 ( .A1(n13553), .A2(n13552), .ZN(n13555) );
  OAI21_X1 U16827 ( .B1(n13555), .B2(n12287), .A(n13554), .ZN(n13556) );
  MUX2_X1 U16828 ( .A(n13557), .B(n13556), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13558) );
  AOI211_X1 U16829 ( .C1(n13270), .C2(n13559), .A(n10806), .B(n13558), .ZN(
        n15698) );
  MUX2_X1 U16830 ( .A(n15698), .B(n10489), .S(n15685), .Z(n13577) );
  OR2_X1 U16831 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13577), .ZN(
        n13560) );
  AOI221_X1 U16832 ( .B1(n13561), .B2(n13560), .C1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n13577), .A(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n13579) );
  OR2_X1 U16833 ( .A1(n13562), .A2(n10456), .ZN(n13566) );
  INV_X1 U16834 ( .A(n13563), .ZN(n13564) );
  NAND2_X1 U16835 ( .A1(n13568), .A2(n13564), .ZN(n13565) );
  OAI211_X1 U16836 ( .C1(n13568), .C2(n13567), .A(n13566), .B(n13565), .ZN(
        n20104) );
  OAI21_X1 U16837 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n13569), .ZN(n13573) );
  INV_X1 U16838 ( .A(n15856), .ZN(n13570) );
  NAND3_X1 U16839 ( .A1(n14916), .A2(n13571), .A3(n13570), .ZN(n13572) );
  OAI211_X1 U16840 ( .C1(n20115), .C2(n20106), .A(n13573), .B(n13572), .ZN(
        n13574) );
  NOR2_X1 U16841 ( .A1(n20104), .A2(n13574), .ZN(n13575) );
  OAI21_X1 U16842 ( .B1(n13577), .B2(n13576), .A(n13575), .ZN(n13578) );
  AOI211_X1 U16843 ( .C1(n15685), .C2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n13579), .B(n13578), .ZN(n16606) );
  INV_X1 U16844 ( .A(n16606), .ZN(n13580) );
  OAI21_X1 U16845 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(n13580), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n13581) );
  OAI21_X1 U16846 ( .B1(n19976), .B2(n19974), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n13584) );
  NAND2_X1 U16847 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13583), .ZN(n16119) );
  NAND2_X1 U16848 ( .A1(n13584), .A2(n16119), .ZN(P2_U3593) );
  AOI21_X1 U16849 ( .B1(n13586), .B2(n13585), .A(n13599), .ZN(n19296) );
  INV_X1 U16850 ( .A(n19296), .ZN(n13592) );
  OAI211_X1 U16851 ( .C1(n13587), .C2(n13589), .A(n13588), .B(n15109), .ZN(
        n13591) );
  NAND2_X1 U16852 ( .A1(n15089), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13590) );
  OAI211_X1 U16853 ( .C1(n13592), .C2(n15089), .A(n13591), .B(n13590), .ZN(
        P2_U2879) );
  INV_X1 U16854 ( .A(n13624), .ZN(n13692) );
  AOI22_X1 U16855 ( .A1(n20727), .A2(n13692), .B1(n20725), .B2(n13691), .ZN(
        n13594) );
  NAND2_X1 U16856 ( .A1(n13790), .A2(n20728), .ZN(n13593) );
  OAI211_X1 U16857 ( .C1(n13697), .C2(n20733), .A(n13594), .B(n13593), .ZN(
        n13595) );
  AOI21_X1 U16858 ( .B1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n13699), .A(
        n13595), .ZN(n13596) );
  INV_X1 U16859 ( .A(n13596), .ZN(P1_U3096) );
  XNOR2_X1 U16860 ( .A(n13588), .B(n13597), .ZN(n13604) );
  INV_X1 U16861 ( .A(n13598), .ZN(n13601) );
  INV_X1 U16862 ( .A(n13599), .ZN(n13600) );
  NAND2_X1 U16863 ( .A1(n13601), .A2(n13600), .ZN(n13602) );
  AND2_X1 U16864 ( .A1(n13602), .A2(n14871), .ZN(n16493) );
  INV_X1 U16865 ( .A(n16493), .ZN(n15626) );
  MUX2_X1 U16866 ( .A(n10119), .B(n15626), .S(n15116), .Z(n13603) );
  OAI21_X1 U16867 ( .B1(n13604), .B2(n15106), .A(n13603), .ZN(P2_U2878) );
  AOI21_X1 U16868 ( .B1(n13606), .B2(n13368), .A(n13605), .ZN(n13851) );
  AOI21_X1 U16869 ( .B1(n16194), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n13607), .ZN(n13608) );
  OAI21_X1 U16870 ( .B1(n13842), .B2(n16202), .A(n13608), .ZN(n13609) );
  AOI21_X1 U16871 ( .B1(n13851), .B2(n16205), .A(n13609), .ZN(n13610) );
  OAI21_X1 U16872 ( .B1(n20135), .B2(n13611), .A(n13610), .ZN(P1_U2995) );
  INV_X1 U16873 ( .A(n13851), .ZN(n13675) );
  INV_X1 U16874 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20238) );
  OAI222_X1 U16875 ( .A1(n13675), .A2(n14505), .B1(n14500), .B2(n13623), .C1(
        n20238), .C2(n14498), .ZN(P1_U2900) );
  AOI22_X1 U16876 ( .A1(DATAI_21_), .A2(n13686), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n13687), .ZN(n20717) );
  INV_X1 U16877 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n19473) );
  INV_X1 U16878 ( .A(DATAI_29_), .ZN(n20891) );
  OAI22_X2 U16879 ( .A1(n19473), .A2(n13694), .B1(n20891), .B2(n13693), .ZN(
        n20714) );
  NOR2_X2 U16880 ( .A1(n13690), .A2(n14432), .ZN(n20713) );
  INV_X1 U16881 ( .A(n20713), .ZN(n13612) );
  NOR2_X2 U16882 ( .A1(n13720), .A2(n20298), .ZN(n20712) );
  INV_X1 U16883 ( .A(n20712), .ZN(n20629) );
  OAI22_X1 U16884 ( .A1(n13612), .A2(n13625), .B1(n13624), .B2(n20629), .ZN(
        n13613) );
  AOI21_X1 U16885 ( .B1(n13790), .B2(n20714), .A(n13613), .ZN(n13615) );
  NAND2_X1 U16886 ( .A1(n13699), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n13614) );
  OAI211_X1 U16887 ( .C1(n9831), .C2(n13697), .A(n13615), .B(n13614), .ZN(
        P1_U3094) );
  AOI22_X1 U16888 ( .A1(DATAI_18_), .A2(n13686), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n13687), .ZN(n20699) );
  INV_X1 U16889 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n19457) );
  INV_X1 U16890 ( .A(DATAI_26_), .ZN(n20931) );
  OAI22_X2 U16891 ( .A1(n19457), .A2(n13694), .B1(n20931), .B2(n13693), .ZN(
        n20696) );
  NOR2_X2 U16892 ( .A1(n13690), .A2(n13616), .ZN(n20743) );
  INV_X1 U16893 ( .A(n20743), .ZN(n13618) );
  NOR2_X2 U16894 ( .A1(n13617), .A2(n20298), .ZN(n20741) );
  INV_X1 U16895 ( .A(n20741), .ZN(n20619) );
  OAI22_X1 U16896 ( .A1(n13618), .A2(n13625), .B1(n13624), .B2(n20619), .ZN(
        n13619) );
  AOI21_X1 U16897 ( .B1(n13790), .B2(n20696), .A(n13619), .ZN(n13621) );
  NAND2_X1 U16898 ( .A1(n13699), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n13620) );
  OAI211_X1 U16899 ( .C1(n20699), .C2(n13697), .A(n13621), .B(n13620), .ZN(
        P1_U3091) );
  AOI22_X1 U16900 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n13687), .B1(DATAI_20_), 
        .B2(n13686), .ZN(n20711) );
  INV_X1 U16901 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16685) );
  INV_X1 U16902 ( .A(DATAI_28_), .ZN(n20995) );
  OAI22_X2 U16903 ( .A1(n16685), .A2(n13694), .B1(n20995), .B2(n13693), .ZN(
        n20708) );
  NOR2_X2 U16904 ( .A1(n13690), .A2(n13622), .ZN(n20707) );
  INV_X1 U16905 ( .A(n20707), .ZN(n13626) );
  NOR2_X2 U16906 ( .A1(n13623), .A2(n20298), .ZN(n20706) );
  INV_X1 U16907 ( .A(n20706), .ZN(n20626) );
  OAI22_X1 U16908 ( .A1(n13626), .A2(n13625), .B1(n13624), .B2(n20626), .ZN(
        n13627) );
  AOI21_X1 U16909 ( .B1(n13790), .B2(n20708), .A(n13627), .ZN(n13629) );
  NAND2_X1 U16910 ( .A1(n13699), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n13628) );
  OAI211_X1 U16911 ( .C1(n20711), .C2(n13697), .A(n13629), .B(n13628), .ZN(
        P1_U3093) );
  NOR2_X1 U16912 ( .A1(n13630), .A2(n13631), .ZN(n13716) );
  INV_X1 U16913 ( .A(n13632), .ZN(n13634) );
  INV_X1 U16914 ( .A(n13633), .ZN(n13748) );
  OAI21_X1 U16915 ( .B1(n13716), .B2(n13634), .A(n13748), .ZN(n20179) );
  INV_X1 U16916 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20215) );
  NAND2_X1 U16917 ( .A1(n14154), .A2(n20215), .ZN(n13638) );
  NAND2_X1 U16918 ( .A1(n14140), .A2(n20215), .ZN(n13635) );
  OAI211_X1 U16919 ( .C1(n14188), .C2(n13636), .A(n13635), .B(n13292), .ZN(
        n13637) );
  AND2_X1 U16920 ( .A1(n13638), .A2(n13637), .ZN(n13723) );
  MUX2_X1 U16921 ( .A(n14166), .B(n13292), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n13640) );
  NAND2_X1 U16922 ( .A1(n14163), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13639) );
  NAND2_X1 U16923 ( .A1(n13640), .A2(n13639), .ZN(n13755) );
  XNOR2_X1 U16924 ( .A(n13758), .B(n13755), .ZN(n20182) );
  AOI22_X1 U16925 ( .A1(n20182), .A2(n14430), .B1(n14429), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n13641) );
  OAI21_X1 U16926 ( .B1(n20179), .B2(n14420), .A(n13641), .ZN(P1_U2866) );
  INV_X1 U16927 ( .A(n14460), .ZN(n13688) );
  OAI222_X1 U16928 ( .A1(n20179), .A2(n14505), .B1(n14500), .B2(n13688), .C1(
        n14498), .C2(n11329), .ZN(P1_U2898) );
  INV_X1 U16929 ( .A(n20845), .ZN(n16096) );
  NAND2_X1 U16930 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n16096), .ZN(n16093) );
  OAI21_X1 U16931 ( .B1(n20846), .B2(n16093), .A(n14779), .ZN(n13642) );
  INV_X1 U16932 ( .A(n13642), .ZN(n13646) );
  NAND2_X1 U16933 ( .A1(n13644), .A2(n13643), .ZN(n13645) );
  NAND2_X1 U16934 ( .A1(n13646), .A2(n13645), .ZN(n13647) );
  NAND2_X1 U16935 ( .A1(n13649), .A2(n13663), .ZN(n13650) );
  NAND2_X1 U16936 ( .A1(n20178), .A2(n13650), .ZN(n20199) );
  INV_X1 U16937 ( .A(n20199), .ZN(n14384) );
  INV_X1 U16938 ( .A(n13652), .ZN(n20674) );
  INV_X1 U16939 ( .A(n13663), .ZN(n13653) );
  OR2_X1 U16940 ( .A1(n13654), .A2(n13653), .ZN(n13847) );
  INV_X1 U16941 ( .A(n13847), .ZN(n14381) );
  INV_X1 U16942 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14385) );
  NAND2_X1 U16943 ( .A1(n13660), .A2(n14385), .ZN(n13655) );
  NAND2_X1 U16944 ( .A1(n13656), .A2(n13655), .ZN(n13659) );
  AND2_X1 U16945 ( .A1(n20850), .A2(n20841), .ZN(n16086) );
  OAI21_X1 U16946 ( .B1(n9666), .B2(n13657), .A(n16086), .ZN(n13662) );
  AND3_X2 U16947 ( .A1(n13659), .A2(n13663), .A3(n13662), .ZN(n20175) );
  NAND2_X1 U16948 ( .A1(n13660), .A2(n13663), .ZN(n13661) );
  AOI22_X1 U16949 ( .A1(n20175), .A2(P1_EBX_REG_1__SCAN_IN), .B1(n13763), .B2(
        n20832), .ZN(n13668) );
  INV_X1 U16950 ( .A(n16086), .ZN(n13664) );
  AND3_X1 U16951 ( .A1(n13664), .A2(P1_EBX_REG_31__SCAN_IN), .A3(n13663), .ZN(
        n13665) );
  NAND2_X1 U16952 ( .A1(n13666), .A2(n20183), .ZN(n13667) );
  OAI211_X1 U16953 ( .C1(n13734), .C2(n20832), .A(n13668), .B(n13667), .ZN(
        n13672) );
  NOR2_X1 U16954 ( .A1(n13669), .A2(n16345), .ZN(n13670) );
  MUX2_X1 U16955 ( .A(n20197), .B(n20196), .S(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n13671) );
  AOI211_X1 U16956 ( .C1(n20674), .C2(n14381), .A(n13672), .B(n13671), .ZN(
        n13673) );
  OAI21_X1 U16957 ( .B1(n13674), .B2(n14384), .A(n13673), .ZN(P1_U2839) );
  INV_X1 U16958 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13676) );
  OAI222_X1 U16959 ( .A1(n13677), .A2(n20209), .B1(n20216), .B2(n13676), .C1(
        n14420), .C2(n13675), .ZN(P1_U2868) );
  INV_X1 U16960 ( .A(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13681) );
  AOI22_X1 U16961 ( .A1(n20713), .A2(n20742), .B1(n20712), .B2(n20740), .ZN(
        n13678) );
  OAI21_X1 U16962 ( .B1(n9831), .B2(n20295), .A(n13678), .ZN(n13679) );
  AOI21_X1 U16963 ( .B1(n20714), .B2(n20682), .A(n13679), .ZN(n13680) );
  OAI21_X1 U16964 ( .B1(n13715), .B2(n13681), .A(n13680), .ZN(P1_U3158) );
  INV_X1 U16965 ( .A(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13685) );
  AOI22_X1 U16966 ( .A1(n20707), .A2(n20742), .B1(n20706), .B2(n20740), .ZN(
        n13682) );
  OAI21_X1 U16967 ( .B1(n20711), .B2(n20295), .A(n13682), .ZN(n13683) );
  AOI21_X1 U16968 ( .B1(n20708), .B2(n20682), .A(n13683), .ZN(n13684) );
  OAI21_X1 U16969 ( .B1(n13715), .B2(n13685), .A(n13684), .ZN(P1_U3157) );
  AOI22_X1 U16970 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n13687), .B1(DATAI_22_), 
        .B2(n13686), .ZN(n20723) );
  NOR2_X2 U16971 ( .A1(n20298), .A2(n13688), .ZN(n20719) );
  NOR2_X2 U16972 ( .A1(n13690), .A2(n13689), .ZN(n20718) );
  AOI22_X1 U16973 ( .A1(n20719), .A2(n13692), .B1(n20718), .B2(n13691), .ZN(
        n13696) );
  INV_X1 U16974 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16682) );
  INV_X1 U16975 ( .A(DATAI_30_), .ZN(n21009) );
  OAI22_X2 U16976 ( .A1(n16682), .A2(n13694), .B1(n21009), .B2(n13693), .ZN(
        n20720) );
  NAND2_X1 U16977 ( .A1(n13790), .A2(n20720), .ZN(n13695) );
  OAI211_X1 U16978 ( .C1(n13697), .C2(n20723), .A(n13696), .B(n13695), .ZN(
        n13698) );
  AOI21_X1 U16979 ( .B1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B2(n13699), .A(
        n13698), .ZN(n13700) );
  INV_X1 U16980 ( .A(n13700), .ZN(P1_U3095) );
  XNOR2_X1 U16981 ( .A(n13702), .B(n13701), .ZN(n16576) );
  XNOR2_X1 U16982 ( .A(n13703), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13704) );
  XNOR2_X1 U16983 ( .A(n13705), .B(n13704), .ZN(n16579) );
  NAND2_X1 U16984 ( .A1(n16579), .A2(n16495), .ZN(n13710) );
  OAI22_X1 U16985 ( .A1(n19438), .A2(n13706), .B1(n10684), .B2(n19300), .ZN(
        n13708) );
  NOR2_X1 U16986 ( .A1(n16491), .A2(n14930), .ZN(n13707) );
  AOI211_X1 U16987 ( .C1(n13270), .C2(n19435), .A(n13708), .B(n13707), .ZN(
        n13709) );
  OAI211_X1 U16988 ( .C1(n16576), .C2(n19429), .A(n13710), .B(n13709), .ZN(
        P2_U3011) );
  INV_X1 U16989 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13714) );
  AOI22_X1 U16990 ( .A1(n20719), .A2(n20740), .B1(n20718), .B2(n20742), .ZN(
        n13711) );
  OAI21_X1 U16991 ( .B1(n20723), .B2(n20295), .A(n13711), .ZN(n13712) );
  AOI21_X1 U16992 ( .B1(n20720), .B2(n20682), .A(n13712), .ZN(n13713) );
  OAI21_X1 U16993 ( .B1(n13715), .B2(n13714), .A(n13713), .ZN(P1_U3159) );
  INV_X1 U16994 ( .A(n13716), .ZN(n13718) );
  NAND2_X1 U16995 ( .A1(n13631), .A2(n13630), .ZN(n13717) );
  AND2_X1 U16996 ( .A1(n13718), .A2(n13717), .ZN(n20213) );
  INV_X1 U16997 ( .A(n20213), .ZN(n13719) );
  OAI222_X1 U16998 ( .A1(n14500), .A2(n13720), .B1(n14498), .B2(n11310), .C1(
        n14505), .C2(n13719), .ZN(P1_U2899) );
  XOR2_X1 U16999 ( .A(n13722), .B(n13721), .Z(n16206) );
  OR2_X1 U17000 ( .A1(n13724), .A2(n13723), .ZN(n13725) );
  NAND2_X1 U17001 ( .A1(n13758), .A2(n13725), .ZN(n20210) );
  INV_X1 U17002 ( .A(n13729), .ZN(n13728) );
  NAND2_X1 U17003 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13728), .ZN(
        n13923) );
  INV_X1 U17004 ( .A(n13923), .ZN(n13912) );
  NAND2_X1 U17005 ( .A1(n13912), .A2(n13726), .ZN(n14642) );
  AOI21_X1 U17006 ( .B1(n14765), .B2(n14642), .A(n14652), .ZN(n14766) );
  OAI211_X1 U17007 ( .C1(n16284), .C2(n13728), .A(n14766), .B(n13727), .ZN(
        n16309) );
  NOR2_X1 U17008 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13729), .ZN(
        n16310) );
  AOI22_X1 U17009 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n16309), .B1(
        n16310), .B2(n13911), .ZN(n13730) );
  NAND2_X1 U17010 ( .A1(n16319), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n16207) );
  OAI211_X1 U17011 ( .C1(n16259), .C2(n20210), .A(n13730), .B(n16207), .ZN(
        n13731) );
  AOI21_X1 U17012 ( .B1(n16206), .B2(n20285), .A(n13731), .ZN(n13732) );
  INV_X1 U17013 ( .A(n13732), .ZN(P1_U3026) );
  NAND2_X1 U17014 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n13733) );
  NOR2_X1 U17015 ( .A1(n13768), .A2(n13733), .ZN(n14378) );
  INV_X1 U17016 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n13735) );
  OAI21_X1 U17017 ( .B1(n13736), .B2(n20832), .A(n13735), .ZN(n13737) );
  NAND2_X1 U17018 ( .A1(n20185), .A2(n13737), .ZN(n13746) );
  NAND2_X1 U17019 ( .A1(n13738), .A2(n20199), .ZN(n13745) );
  INV_X1 U17020 ( .A(n13068), .ZN(n20297) );
  AOI22_X1 U17021 ( .A1(n20196), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20175), .B2(P1_EBX_REG_2__SCAN_IN), .ZN(n13741) );
  NAND2_X1 U17022 ( .A1(n13739), .A2(n20183), .ZN(n13740) );
  OAI211_X1 U17023 ( .C1(n20189), .C2(n13742), .A(n13741), .B(n13740), .ZN(
        n13743) );
  AOI21_X1 U17024 ( .B1(n20297), .B2(n14381), .A(n13743), .ZN(n13744) );
  OAI211_X1 U17025 ( .C1(n14378), .C2(n13746), .A(n13745), .B(n13744), .ZN(
        P1_U2838) );
  INV_X1 U17026 ( .A(n13747), .ZN(n13749) );
  AOI21_X1 U17027 ( .B1(n13749), .B2(n13748), .A(n9704), .ZN(n16199) );
  INV_X1 U17028 ( .A(n16199), .ZN(n20169) );
  INV_X1 U17029 ( .A(n13758), .ZN(n13754) );
  INV_X1 U17030 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n13750) );
  NAND2_X1 U17031 ( .A1(n14154), .A2(n13750), .ZN(n13753) );
  INV_X1 U17032 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16324) );
  NAND2_X1 U17033 ( .A1(n14140), .A2(n13750), .ZN(n13751) );
  OAI211_X1 U17034 ( .C1(n14188), .C2(n16324), .A(n13751), .B(n13292), .ZN(
        n13752) );
  AND2_X1 U17035 ( .A1(n13753), .A2(n13752), .ZN(n13756) );
  AOI21_X1 U17036 ( .B1(n13754), .B2(n13755), .A(n13756), .ZN(n13759) );
  NAND2_X1 U17037 ( .A1(n13756), .A2(n13755), .ZN(n13757) );
  NOR2_X1 U17038 ( .A1(n13759), .A2(n9800), .ZN(n20165) );
  AOI22_X1 U17039 ( .A1(n20165), .A2(n14430), .B1(n14429), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n13760) );
  OAI21_X1 U17040 ( .B1(n20169), .B2(n14420), .A(n13760), .ZN(P1_U2865) );
  OAI222_X1 U17041 ( .A1(n20169), .A2(n14505), .B1(n14500), .B2(n13761), .C1(
        n14498), .C2(n11386), .ZN(P1_U2897) );
  OAI21_X1 U17042 ( .B1(n9704), .B2(n10277), .A(n13762), .ZN(n13866) );
  NAND2_X1 U17043 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .ZN(n13764) );
  NAND3_X1 U17044 ( .A1(n20190), .A2(P1_REIP_REG_6__SCAN_IN), .A3(
        P1_REIP_REG_5__SCAN_IN), .ZN(n20173) );
  NOR2_X1 U17045 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20173), .ZN(n13776) );
  MUX2_X1 U17046 ( .A(n14166), .B(n13292), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n13766) );
  NAND2_X1 U17047 ( .A1(n14163), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13765) );
  NAND2_X1 U17048 ( .A1(n13766), .A2(n13765), .ZN(n16294) );
  XNOR2_X1 U17049 ( .A(n9800), .B(n16294), .ZN(n16305) );
  NAND2_X1 U17050 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n13767) );
  NAND3_X1 U17051 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(n14378), .ZN(n20184) );
  NOR2_X1 U17052 ( .A1(n13767), .A2(n20184), .ZN(n20162) );
  NAND3_X1 U17053 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .A3(n20162), .ZN(n13870) );
  AND2_X1 U17054 ( .A1(n20185), .A2(n13870), .ZN(n20157) );
  NOR2_X1 U17055 ( .A1(n13769), .A2(n13768), .ZN(n16156) );
  INV_X1 U17056 ( .A(n16156), .ZN(n20191) );
  INV_X1 U17057 ( .A(n20191), .ZN(n20174) );
  AOI21_X1 U17058 ( .B1(n20175), .B2(P1_EBX_REG_8__SCAN_IN), .A(n20174), .ZN(
        n13772) );
  INV_X1 U17059 ( .A(n13862), .ZN(n13770) );
  NAND2_X1 U17060 ( .A1(n20197), .A2(n13770), .ZN(n13771) );
  OAI211_X1 U17061 ( .C1(n20177), .C2(n11400), .A(n13772), .B(n13771), .ZN(
        n13773) );
  AOI21_X1 U17062 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(n20157), .A(n13773), .ZN(
        n13774) );
  OAI21_X1 U17063 ( .B1(n16305), .B2(n20193), .A(n13774), .ZN(n13775) );
  AOI21_X1 U17064 ( .B1(n13776), .B2(P1_REIP_REG_7__SCAN_IN), .A(n13775), .ZN(
        n13777) );
  OAI21_X1 U17065 ( .B1(n13866), .B2(n20178), .A(n13777), .ZN(P1_U2832) );
  INV_X1 U17066 ( .A(DATAI_8_), .ZN(n20930) );
  NAND2_X1 U17067 ( .A1(n14438), .A2(BUF1_REG_8__SCAN_IN), .ZN(n13778) );
  OAI21_X1 U17068 ( .B1(n14438), .B2(n20930), .A(n13778), .ZN(n20248) );
  AOI22_X1 U17069 ( .A1(n14503), .A2(n20248), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n14502), .ZN(n13779) );
  OAI21_X1 U17070 ( .B1(n13866), .B2(n14505), .A(n13779), .ZN(P1_U2896) );
  NOR2_X1 U17071 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13780), .ZN(
        n13819) );
  NOR2_X1 U17072 ( .A1(n13786), .A2(n20753), .ZN(n20530) );
  NOR3_X1 U17073 ( .A1(n13790), .A2(n20678), .A3(n20461), .ZN(n13782) );
  NOR2_X1 U17074 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n20678), .ZN(n20526) );
  NOR2_X1 U17075 ( .A1(n13782), .A2(n20526), .ZN(n13789) );
  INV_X1 U17076 ( .A(n13789), .ZN(n13783) );
  OR2_X1 U17077 ( .A1(n20413), .A2(n13652), .ZN(n13788) );
  OR2_X1 U17078 ( .A1(n20529), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20356) );
  AND2_X1 U17079 ( .A1(n20356), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20352) );
  AOI21_X1 U17080 ( .B1(n13783), .B2(n13788), .A(n20352), .ZN(n13784) );
  OAI211_X1 U17081 ( .C1(n13819), .C2(n20609), .A(n20686), .B(n13784), .ZN(
        n13785) );
  INV_X1 U17082 ( .A(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13794) );
  INV_X1 U17083 ( .A(n13786), .ZN(n13787) );
  NOR2_X1 U17084 ( .A1(n13787), .A2(n20753), .ZN(n20601) );
  INV_X1 U17085 ( .A(n20601), .ZN(n20676) );
  OAI22_X1 U17086 ( .A1(n13789), .A2(n13788), .B1(n20676), .B2(n20356), .ZN(
        n13823) );
  INV_X1 U17087 ( .A(n13790), .ZN(n13821) );
  AOI22_X1 U17088 ( .A1(n20461), .A2(n20728), .B1(n20725), .B2(n13819), .ZN(
        n13791) );
  OAI21_X1 U17089 ( .B1(n13821), .B2(n20733), .A(n13791), .ZN(n13792) );
  AOI21_X1 U17090 ( .B1(n13823), .B2(n20727), .A(n13792), .ZN(n13793) );
  OAI21_X1 U17091 ( .B1(n13826), .B2(n13794), .A(n13793), .ZN(P1_U3088) );
  INV_X1 U17092 ( .A(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13798) );
  AOI22_X1 U17093 ( .A1(n20461), .A2(n20692), .B1(n20735), .B2(n13819), .ZN(
        n13795) );
  OAI21_X1 U17094 ( .B1(n13821), .B2(n20695), .A(n13795), .ZN(n13796) );
  AOI21_X1 U17095 ( .B1(n13823), .B2(n20734), .A(n13796), .ZN(n13797) );
  OAI21_X1 U17096 ( .B1(n13826), .B2(n13798), .A(n13797), .ZN(P1_U3082) );
  INV_X1 U17097 ( .A(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13802) );
  AOI22_X1 U17098 ( .A1(n20461), .A2(n20714), .B1(n20713), .B2(n13819), .ZN(
        n13799) );
  OAI21_X1 U17099 ( .B1(n13821), .B2(n9831), .A(n13799), .ZN(n13800) );
  AOI21_X1 U17100 ( .B1(n13823), .B2(n20712), .A(n13800), .ZN(n13801) );
  OAI21_X1 U17101 ( .B1(n13826), .B2(n13802), .A(n13801), .ZN(P1_U3086) );
  INV_X1 U17102 ( .A(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13806) );
  AOI22_X1 U17103 ( .A1(n20461), .A2(n20708), .B1(n20707), .B2(n13819), .ZN(
        n13803) );
  OAI21_X1 U17104 ( .B1(n13821), .B2(n20711), .A(n13803), .ZN(n13804) );
  AOI21_X1 U17105 ( .B1(n13823), .B2(n20706), .A(n13804), .ZN(n13805) );
  OAI21_X1 U17106 ( .B1(n13826), .B2(n13806), .A(n13805), .ZN(P1_U3085) );
  INV_X1 U17107 ( .A(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13810) );
  AOI22_X1 U17108 ( .A1(n20461), .A2(n20720), .B1(n20718), .B2(n13819), .ZN(
        n13807) );
  OAI21_X1 U17109 ( .B1(n13821), .B2(n20723), .A(n13807), .ZN(n13808) );
  AOI21_X1 U17110 ( .B1(n13823), .B2(n20719), .A(n13808), .ZN(n13809) );
  OAI21_X1 U17111 ( .B1(n13826), .B2(n13810), .A(n13809), .ZN(P1_U3087) );
  INV_X1 U17112 ( .A(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13814) );
  AOI22_X1 U17113 ( .A1(n20461), .A2(n20702), .B1(n20701), .B2(n13819), .ZN(
        n13811) );
  OAI21_X1 U17114 ( .B1(n13821), .B2(n9829), .A(n13811), .ZN(n13812) );
  AOI21_X1 U17115 ( .B1(n13823), .B2(n20700), .A(n13812), .ZN(n13813) );
  OAI21_X1 U17116 ( .B1(n13826), .B2(n13814), .A(n13813), .ZN(P1_U3084) );
  INV_X1 U17117 ( .A(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13818) );
  AOI22_X1 U17118 ( .A1(n20461), .A2(n20696), .B1(n20743), .B2(n13819), .ZN(
        n13815) );
  OAI21_X1 U17119 ( .B1(n13821), .B2(n20699), .A(n13815), .ZN(n13816) );
  AOI21_X1 U17120 ( .B1(n13823), .B2(n20741), .A(n13816), .ZN(n13817) );
  OAI21_X1 U17121 ( .B1(n13826), .B2(n13818), .A(n13817), .ZN(P1_U3083) );
  INV_X1 U17122 ( .A(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13825) );
  AOI22_X1 U17123 ( .A1(n20461), .A2(n20688), .B1(n20680), .B2(n13819), .ZN(
        n13820) );
  OAI21_X1 U17124 ( .B1(n20691), .B2(n13821), .A(n13820), .ZN(n13822) );
  AOI21_X1 U17125 ( .B1(n13823), .B2(n20679), .A(n13822), .ZN(n13824) );
  OAI21_X1 U17126 ( .B1(n13826), .B2(n13825), .A(n13824), .ZN(P1_U3081) );
  OAI22_X1 U17127 ( .A1(n20278), .A2(n20193), .B1(n13827), .B2(n20192), .ZN(
        n13830) );
  AOI21_X1 U17128 ( .B1(n20177), .B2(n20189), .A(n13828), .ZN(n13829) );
  AOI211_X1 U17129 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(n20185), .A(n13830), .B(
        n13829), .ZN(n13832) );
  NAND2_X1 U17130 ( .A1(n11347), .A2(n14381), .ZN(n13831) );
  OAI211_X1 U17131 ( .C1(n13833), .C2(n14384), .A(n13832), .B(n13831), .ZN(
        P1_U2840) );
  XOR2_X1 U17132 ( .A(n13834), .B(n13835), .Z(n16330) );
  NAND2_X1 U17133 ( .A1(n16330), .A2(n11980), .ZN(n13838) );
  INV_X1 U17134 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20777) );
  NOR2_X1 U17135 ( .A1(n14779), .A2(n20777), .ZN(n16326) );
  NOR2_X1 U17136 ( .A1(n16202), .A2(n20188), .ZN(n13836) );
  AOI211_X1 U17137 ( .C1(n16194), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16326), .B(n13836), .ZN(n13837) );
  OAI211_X1 U17138 ( .C1(n14551), .C2(n20179), .A(n13838), .B(n13837), .ZN(
        P1_U2993) );
  INV_X1 U17139 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13839) );
  OAI222_X1 U17140 ( .A1(n13866), .A2(n14420), .B1(n20209), .B2(n16305), .C1(
        n20216), .C2(n13839), .ZN(P1_U2864) );
  NOR3_X1 U17141 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n14372), .A3(n20771), .ZN(
        n13850) );
  INV_X1 U17142 ( .A(n16337), .ZN(n13848) );
  NAND3_X1 U17143 ( .A1(n20184), .A2(n20185), .A3(P1_REIP_REG_4__SCAN_IN), 
        .ZN(n13846) );
  AOI21_X1 U17144 ( .B1(n20175), .B2(P1_EBX_REG_4__SCAN_IN), .A(n16156), .ZN(
        n13841) );
  NAND2_X1 U17145 ( .A1(n20196), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13840) );
  OAI211_X1 U17146 ( .C1(n20189), .C2(n13842), .A(n13841), .B(n13840), .ZN(
        n13843) );
  AOI21_X1 U17147 ( .B1(n20183), .B2(n13844), .A(n13843), .ZN(n13845) );
  OAI211_X1 U17148 ( .C1(n13848), .C2(n13847), .A(n13846), .B(n13845), .ZN(
        n13849) );
  AOI211_X1 U17149 ( .C1(n13851), .C2(n20199), .A(n13850), .B(n13849), .ZN(
        n13852) );
  INV_X1 U17150 ( .A(n13852), .ZN(P1_U2836) );
  AND2_X1 U17151 ( .A1(n13762), .A2(n13853), .ZN(n13855) );
  OR2_X1 U17152 ( .A1(n13855), .A2(n13854), .ZN(n20205) );
  INV_X1 U17153 ( .A(DATAI_9_), .ZN(n20915) );
  NAND2_X1 U17154 ( .A1(n14438), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13856) );
  OAI21_X1 U17155 ( .B1(n14438), .B2(n20915), .A(n13856), .ZN(n20250) );
  AOI22_X1 U17156 ( .A1(n14503), .A2(n20250), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n14502), .ZN(n13857) );
  OAI21_X1 U17157 ( .B1(n20205), .B2(n14505), .A(n13857), .ZN(P1_U2895) );
  XNOR2_X1 U17158 ( .A(n13858), .B(n16314), .ZN(n13859) );
  XNOR2_X1 U17159 ( .A(n13860), .B(n13859), .ZN(n16313) );
  NAND2_X1 U17160 ( .A1(n16313), .A2(n11980), .ZN(n13865) );
  INV_X1 U17161 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n13861) );
  NOR2_X1 U17162 ( .A1(n14779), .A2(n13861), .ZN(n16306) );
  NOR2_X1 U17163 ( .A1(n16202), .A2(n13862), .ZN(n13863) );
  AOI211_X1 U17164 ( .C1(n16194), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16306), .B(n13863), .ZN(n13864) );
  OAI211_X1 U17165 ( .C1(n14551), .C2(n13866), .A(n13865), .B(n13864), .ZN(
        P1_U2991) );
  XOR2_X1 U17166 ( .A(n13867), .B(n13854), .Z(n14636) );
  INV_X1 U17167 ( .A(n14636), .ZN(n13884) );
  AOI22_X1 U17168 ( .A1(n14503), .A2(n14448), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n14502), .ZN(n13868) );
  OAI21_X1 U17169 ( .B1(n13884), .B2(n14505), .A(n13868), .ZN(P1_U2894) );
  NAND2_X1 U17170 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .ZN(n13869) );
  NAND2_X1 U17171 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n13871) );
  NOR2_X1 U17172 ( .A1(n13871), .A2(n13870), .ZN(n14075) );
  OAI221_X1 U17173 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(P1_REIP_REG_9__SCAN_IN), 
        .C1(P1_REIP_REG_10__SCAN_IN), .C2(n20158), .A(n10269), .ZN(n13883) );
  INV_X1 U17174 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n20208) );
  NAND2_X1 U17175 ( .A1(n14154), .A2(n20208), .ZN(n13874) );
  INV_X1 U17176 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16303) );
  NAND2_X1 U17177 ( .A1(n14140), .A2(n20208), .ZN(n13872) );
  OAI211_X1 U17178 ( .C1(n14188), .C2(n16303), .A(n13872), .B(n13292), .ZN(
        n13873) );
  AND2_X1 U17179 ( .A1(n13874), .A2(n13873), .ZN(n16293) );
  MUX2_X1 U17180 ( .A(n14166), .B(n13292), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n13876) );
  NAND2_X1 U17181 ( .A1(n14163), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13875) );
  NAND2_X1 U17182 ( .A1(n13876), .A2(n13875), .ZN(n13877) );
  OR2_X1 U17183 ( .A1(n16295), .A2(n13877), .ZN(n13878) );
  AND2_X1 U17184 ( .A1(n13900), .A2(n13878), .ZN(n16288) );
  AOI21_X1 U17185 ( .B1(n20175), .B2(P1_EBX_REG_10__SCAN_IN), .A(n16156), .ZN(
        n13880) );
  NAND2_X1 U17186 ( .A1(n20196), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13879) );
  OAI211_X1 U17187 ( .C1(n20189), .C2(n14634), .A(n13880), .B(n13879), .ZN(
        n13881) );
  AOI21_X1 U17188 ( .B1(n16288), .B2(n20183), .A(n13881), .ZN(n13882) );
  OAI211_X1 U17189 ( .C1(n13884), .C2(n20178), .A(n13883), .B(n13882), .ZN(
        P1_U2830) );
  INV_X1 U17190 ( .A(n16288), .ZN(n13886) );
  INV_X1 U17191 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n13885) );
  OAI222_X1 U17192 ( .A1(n13886), .A2(n20209), .B1(n20216), .B2(n13885), .C1(
        n14420), .C2(n13884), .ZN(P1_U2862) );
  XNOR2_X1 U17193 ( .A(n16174), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13887) );
  XNOR2_X1 U17194 ( .A(n13888), .B(n13887), .ZN(n16300) );
  NAND2_X1 U17195 ( .A1(n16300), .A2(n11980), .ZN(n13892) );
  INV_X1 U17196 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n13889) );
  OR2_X1 U17197 ( .A1(n14779), .A2(n13889), .ZN(n16297) );
  OAI21_X1 U17198 ( .B1(n16209), .B2(n20155), .A(n16297), .ZN(n13890) );
  AOI21_X1 U17199 ( .B1(n16204), .B2(n20150), .A(n13890), .ZN(n13891) );
  OAI211_X1 U17200 ( .C1(n14551), .C2(n20205), .A(n13892), .B(n13891), .ZN(
        P1_U2990) );
  INV_X1 U17201 ( .A(n13893), .ZN(n13894) );
  AOI21_X1 U17202 ( .B1(n13896), .B2(n13895), .A(n13894), .ZN(n16190) );
  INV_X1 U17203 ( .A(n16190), .ZN(n13905) );
  MUX2_X1 U17204 ( .A(n14151), .B(n14166), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n13898) );
  NAND2_X1 U17205 ( .A1(n14164), .A2(n11911), .ZN(n13897) );
  NAND2_X1 U17206 ( .A1(n13898), .A2(n13897), .ZN(n13901) );
  INV_X1 U17207 ( .A(n13918), .ZN(n13899) );
  AOI21_X1 U17208 ( .B1(n13901), .B2(n13900), .A(n13899), .ZN(n16275) );
  AOI22_X1 U17209 ( .A1(n16275), .A2(n14430), .B1(n14429), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n13902) );
  OAI21_X1 U17210 ( .B1(n13905), .B2(n14420), .A(n13902), .ZN(P1_U2861) );
  INV_X1 U17211 ( .A(DATAI_11_), .ZN(n20892) );
  NAND2_X1 U17212 ( .A1(n14438), .A2(BUF1_REG_11__SCAN_IN), .ZN(n13903) );
  OAI21_X1 U17213 ( .B1(n14438), .B2(n20892), .A(n13903), .ZN(n20252) );
  AOI22_X1 U17214 ( .A1(n14503), .A2(n20252), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n14502), .ZN(n13904) );
  OAI21_X1 U17215 ( .B1(n13905), .B2(n14505), .A(n13904), .ZN(P1_U2893) );
  NAND2_X1 U17216 ( .A1(n13907), .A2(n13906), .ZN(n13910) );
  OAI21_X1 U17217 ( .B1(n16186), .B2(n14617), .A(n13908), .ZN(n13909) );
  XOR2_X1 U17218 ( .A(n13910), .B(n13909), .Z(n16185) );
  NAND3_X1 U17219 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16290) );
  NOR3_X1 U17220 ( .A1(n14627), .A2(n16303), .A3(n16290), .ZN(n16276) );
  NAND2_X1 U17221 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16276), .ZN(
        n14639) );
  NAND2_X1 U17222 ( .A1(n13912), .A2(n13911), .ZN(n16328) );
  NOR2_X1 U17223 ( .A1(n14639), .A2(n16328), .ZN(n13921) );
  INV_X1 U17224 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14640) );
  NAND2_X1 U17225 ( .A1(n13292), .A2(n14640), .ZN(n13914) );
  INV_X1 U17226 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n14076) );
  NAND2_X1 U17227 ( .A1(n14140), .A2(n14076), .ZN(n13913) );
  NAND3_X1 U17228 ( .A1(n13914), .A2(n14166), .A3(n13913), .ZN(n13916) );
  NAND2_X1 U17229 ( .A1(n13129), .A2(n14076), .ZN(n13915) );
  AND2_X1 U17230 ( .A1(n13916), .A2(n13915), .ZN(n13917) );
  AND2_X1 U17231 ( .A1(n13918), .A2(n13917), .ZN(n13919) );
  NOR2_X1 U17232 ( .A1(n14363), .A2(n13919), .ZN(n13931) );
  INV_X1 U17233 ( .A(n13931), .ZN(n14080) );
  INV_X1 U17234 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n20786) );
  OAI22_X1 U17235 ( .A1(n14080), .A2(n16259), .B1(n20786), .B2(n14779), .ZN(
        n13920) );
  AOI21_X1 U17236 ( .B1(n13921), .B2(n14640), .A(n13920), .ZN(n13927) );
  NOR2_X1 U17237 ( .A1(n13923), .A2(n13922), .ZN(n16283) );
  AOI21_X1 U17238 ( .B1(n16276), .B2(n16283), .A(n16284), .ZN(n13924) );
  INV_X1 U17239 ( .A(n14766), .ZN(n16285) );
  AOI211_X1 U17240 ( .C1(n14765), .C2(n14639), .A(n13924), .B(n16285), .ZN(
        n16281) );
  OAI21_X1 U17241 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16308), .A(
        n16281), .ZN(n13925) );
  NAND2_X1 U17242 ( .A1(n13925), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13926) );
  OAI211_X1 U17243 ( .C1(n16185), .C2(n16260), .A(n13927), .B(n13926), .ZN(
        P1_U3019) );
  OAI21_X1 U17244 ( .B1(n13928), .B2(n13930), .A(n13929), .ZN(n14084) );
  INV_X1 U17245 ( .A(n14084), .ZN(n16182) );
  NAND2_X1 U17246 ( .A1(n16182), .A2(n20212), .ZN(n13933) );
  NAND2_X1 U17247 ( .A1(n13931), .A2(n14430), .ZN(n13932) );
  OAI211_X1 U17248 ( .C1(n14076), .C2(n20216), .A(n13933), .B(n13932), .ZN(
        P1_U2860) );
  NOR2_X1 U17249 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19111) );
  INV_X1 U17250 ( .A(n19111), .ZN(n19146) );
  AOI22_X1 U17251 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13937) );
  AOI22_X1 U17252 ( .A1(n17407), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n15929), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13936) );
  AOI22_X1 U17253 ( .A1(n15864), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13935) );
  AOI22_X1 U17254 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13934) );
  NAND4_X1 U17255 ( .A1(n13937), .A2(n13936), .A3(n13935), .A4(n13934), .ZN(
        n13947) );
  NOR2_X2 U17256 ( .A1(n19092), .A2(n13938), .ZN(n17455) );
  AOI22_X1 U17257 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13945) );
  AOI22_X1 U17258 ( .A1(n17380), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17432), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13944) );
  AOI22_X1 U17259 ( .A1(n9656), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13943) );
  INV_X2 U17260 ( .A(n13974), .ZN(n17395) );
  AOI22_X1 U17261 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n9658), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13942) );
  NAND4_X1 U17262 ( .A1(n13945), .A2(n13944), .A3(n13943), .A4(n13942), .ZN(
        n13946) );
  AOI22_X1 U17263 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17432), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13952) );
  AOI22_X1 U17264 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13951) );
  AOI22_X1 U17265 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13950) );
  AOI22_X1 U17266 ( .A1(n17407), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n15929), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13949) );
  NAND4_X1 U17267 ( .A1(n13952), .A2(n13951), .A3(n13950), .A4(n13949), .ZN(
        n13958) );
  AOI22_X1 U17268 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13956) );
  AOI22_X1 U17269 ( .A1(n15864), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13955) );
  AOI22_X1 U17270 ( .A1(n17380), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9656), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13954) );
  AOI22_X1 U17271 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(n9658), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13953) );
  NAND4_X1 U17272 ( .A1(n13956), .A2(n13955), .A3(n13954), .A4(n13953), .ZN(
        n13957) );
  AOI22_X1 U17273 ( .A1(n17456), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n15929), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13963) );
  AOI22_X1 U17274 ( .A1(n17380), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9656), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13962) );
  AOI22_X1 U17275 ( .A1(n17447), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13961) );
  AOI22_X1 U17276 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13960) );
  NAND4_X1 U17277 ( .A1(n13963), .A2(n13962), .A3(n13961), .A4(n13960), .ZN(
        n13970) );
  AOI22_X1 U17278 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13968) );
  AOI22_X1 U17279 ( .A1(n15864), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13964), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13967) );
  AOI22_X1 U17280 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13966) );
  AOI22_X1 U17281 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(n9658), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13965) );
  NAND4_X1 U17282 ( .A1(n13968), .A2(n13967), .A3(n13966), .A4(n13965), .ZN(
        n13969) );
  AOI22_X1 U17283 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13983) );
  AOI22_X1 U17284 ( .A1(n17432), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17407), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13982) );
  INV_X1 U17285 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13973) );
  AOI22_X1 U17286 ( .A1(n15929), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13972) );
  OAI21_X1 U17287 ( .B1(n13959), .B2(n13973), .A(n13972), .ZN(n13980) );
  AOI22_X1 U17288 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13978) );
  AOI22_X1 U17289 ( .A1(n9656), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13977) );
  AOI22_X1 U17290 ( .A1(n17380), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13976) );
  AOI22_X1 U17291 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(n9658), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13975) );
  NAND4_X1 U17292 ( .A1(n13978), .A2(n13977), .A3(n13976), .A4(n13975), .ZN(
        n13979) );
  NOR2_X1 U17293 ( .A1(n18512), .A2(n17661), .ZN(n14031) );
  AOI22_X1 U17294 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13987) );
  AOI22_X1 U17295 ( .A1(n17380), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13986) );
  AOI22_X1 U17296 ( .A1(n15864), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9656), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13985) );
  AOI22_X1 U17297 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n15929), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13984) );
  NAND4_X1 U17298 ( .A1(n13987), .A2(n13986), .A3(n13985), .A4(n13984), .ZN(
        n13993) );
  AOI22_X1 U17299 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13991) );
  AOI22_X1 U17300 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13990) );
  AOI22_X1 U17301 ( .A1(n17407), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13989) );
  AOI22_X1 U17302 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n9658), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13988) );
  NAND4_X1 U17303 ( .A1(n13991), .A2(n13990), .A3(n13989), .A4(n13988), .ZN(
        n13992) );
  AOI22_X1 U17304 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n15929), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13997) );
  AOI22_X1 U17305 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17407), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13996) );
  AOI22_X1 U17306 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13995) );
  AOI22_X1 U17307 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9656), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13994) );
  NAND4_X1 U17308 ( .A1(n13997), .A2(n13996), .A3(n13995), .A4(n13994), .ZN(
        n14003) );
  AOI22_X1 U17309 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14001) );
  AOI22_X1 U17310 ( .A1(n17432), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14000) );
  AOI22_X1 U17311 ( .A1(n15864), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17380), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13999) );
  AOI22_X1 U17312 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n9658), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13998) );
  NAND4_X1 U17313 ( .A1(n14001), .A2(n14000), .A3(n13999), .A4(n13998), .ZN(
        n14002) );
  NOR2_X1 U17314 ( .A1(n18506), .A2(n18501), .ZN(n15878) );
  NAND4_X1 U17315 ( .A1(n18497), .A2(n18493), .A3(n14031), .A4(n15878), .ZN(
        n14033) );
  NAND2_X1 U17316 ( .A1(n15877), .A2(n18506), .ZN(n18935) );
  AOI22_X1 U17317 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n15929), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14013) );
  AOI22_X1 U17318 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17432), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14012) );
  INV_X1 U17319 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17493) );
  AOI22_X1 U17320 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14004) );
  OAI21_X1 U17321 ( .B1(n13959), .B2(n17493), .A(n14004), .ZN(n14010) );
  AOI22_X1 U17322 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14008) );
  AOI22_X1 U17323 ( .A1(n15864), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9656), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14007) );
  AOI22_X1 U17324 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17407), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14006) );
  AOI22_X1 U17325 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(n9658), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14005) );
  NAND4_X1 U17326 ( .A1(n14008), .A2(n14007), .A3(n14006), .A4(n14005), .ZN(
        n14009) );
  AOI211_X1 U17327 ( .C1(n17380), .C2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A(
        n14010), .B(n14009), .ZN(n14011) );
  NAND3_X1 U17328 ( .A1(n14013), .A2(n14012), .A3(n14011), .ZN(n15883) );
  NAND2_X1 U17329 ( .A1(n18935), .A2(n18489), .ZN(n14032) );
  INV_X1 U17330 ( .A(n18506), .ZN(n17503) );
  NAND2_X1 U17331 ( .A1(n18501), .A2(n17503), .ZN(n14030) );
  INV_X1 U17332 ( .A(n14030), .ZN(n14059) );
  NOR2_X1 U17333 ( .A1(n14032), .A2(n14059), .ZN(n14028) );
  NOR2_X1 U17334 ( .A1(n15883), .A2(n18501), .ZN(n15886) );
  INV_X1 U17335 ( .A(n14048), .ZN(n14029) );
  AOI22_X1 U17336 ( .A1(n17380), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14017) );
  AOI22_X1 U17337 ( .A1(n15864), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13964), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14016) );
  AOI22_X1 U17338 ( .A1(n17432), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14015) );
  AOI22_X1 U17339 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9656), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14014) );
  NAND4_X1 U17340 ( .A1(n14017), .A2(n14016), .A3(n14015), .A4(n14014), .ZN(
        n14023) );
  AOI22_X1 U17341 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14021) );
  AOI22_X1 U17342 ( .A1(n17407), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14020) );
  AOI22_X1 U17343 ( .A1(n15929), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14019) );
  AOI22_X1 U17344 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(n9658), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14018) );
  NAND4_X1 U17345 ( .A1(n14021), .A2(n14020), .A3(n14019), .A4(n14018), .ZN(
        n14022) );
  NOR2_X4 U17346 ( .A1(n14023), .A2(n14022), .ZN(n19136) );
  NAND2_X1 U17347 ( .A1(n18506), .A2(n17511), .ZN(n14056) );
  NAND2_X1 U17348 ( .A1(n17489), .A2(n14056), .ZN(n16125) );
  NAND3_X1 U17349 ( .A1(n19136), .A2(n17661), .A3(n16125), .ZN(n14060) );
  INV_X1 U17350 ( .A(n18493), .ZN(n14024) );
  OAI22_X1 U17351 ( .A1(n14031), .A2(n14024), .B1(n15877), .B2(n14056), .ZN(
        n14027) );
  NOR2_X1 U17352 ( .A1(n18512), .A2(n15878), .ZN(n14025) );
  AOI21_X1 U17353 ( .B1(n18482), .B2(n16806), .A(n15883), .ZN(n14057) );
  OAI22_X1 U17354 ( .A1(n18497), .A2(n14025), .B1(n15878), .B2(n14057), .ZN(
        n14026) );
  AOI211_X1 U17355 ( .C1(n18482), .C2(n14028), .A(n14027), .B(n14026), .ZN(
        n14061) );
  OAI211_X1 U17356 ( .C1(n18493), .C2(n14029), .A(n14060), .B(n14061), .ZN(
        n15985) );
  NOR2_X2 U17357 ( .A1(n14033), .A2(n15985), .ZN(n18929) );
  NAND2_X1 U17358 ( .A1(n18493), .A2(n18489), .ZN(n18934) );
  NAND3_X1 U17359 ( .A1(n14031), .A2(n15831), .A3(n19136), .ZN(n14034) );
  NAND2_X1 U17360 ( .A1(n18506), .A2(n15984), .ZN(n14047) );
  NOR2_X1 U17361 ( .A1(n18489), .A2(n14033), .ZN(n14062) );
  NOR2_X1 U17362 ( .A1(n18976), .A2(n14062), .ZN(n16786) );
  INV_X1 U17363 ( .A(n18976), .ZN(n17700) );
  INV_X1 U17364 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18926) );
  OAI21_X1 U17365 ( .B1(n14035), .B2(n19108), .A(n18926), .ZN(n14067) );
  NAND2_X1 U17366 ( .A1(n18943), .A2(n14067), .ZN(n18925) );
  NOR2_X1 U17367 ( .A1(n19146), .A2(n18925), .ZN(n14066) );
  NAND2_X1 U17368 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19095), .ZN(n16802) );
  NAND2_X1 U17369 ( .A1(n18957), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14049) );
  AOI22_X1 U17370 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n18959), .B2(n19108), .ZN(
        n14053) );
  XNOR2_X1 U17371 ( .A(n14049), .B(n14053), .ZN(n14045) );
  AOI22_X1 U17372 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18964), .B1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n19102), .ZN(n14040) );
  OR2_X1 U17373 ( .A1(n14053), .A2(n14049), .ZN(n14036) );
  NAND2_X1 U17374 ( .A1(n14040), .A2(n14041), .ZN(n14037) );
  OAI21_X1 U17375 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n19102), .A(
        n14037), .ZN(n14038) );
  OAI22_X1 U17376 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18968), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n14038), .ZN(n14042) );
  NOR2_X1 U17377 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18968), .ZN(
        n14039) );
  NAND2_X1 U17378 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n14038), .ZN(
        n14043) );
  AOI22_X1 U17379 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n14042), .B1(
        n14039), .B2(n14043), .ZN(n14050) );
  XOR2_X1 U17380 ( .A(n14041), .B(n14040), .Z(n15876) );
  NAND2_X1 U17381 ( .A1(n14050), .A2(n15876), .ZN(n14051) );
  AOI21_X1 U17382 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n14043), .A(
        n14042), .ZN(n14044) );
  NAND2_X1 U17383 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n19137) );
  NAND2_X1 U17384 ( .A1(n16780), .A2(n19137), .ZN(n14064) );
  NAND2_X2 U17385 ( .A1(n19127), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19072) );
  INV_X1 U17386 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18997) );
  NAND2_X1 U17387 ( .A1(n18997), .A2(n19009), .ZN(n16784) );
  NAND3_X1 U17388 ( .A1(n19007), .A2(n19072), .A3(n16784), .ZN(n19134) );
  INV_X1 U17389 ( .A(n19134), .ZN(n16803) );
  NAND2_X1 U17390 ( .A1(n14046), .A2(n16803), .ZN(n17660) );
  OAI211_X1 U17391 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n18957), .A(
        n14050), .B(n14049), .ZN(n15874) );
  OAI211_X1 U17392 ( .C1(n14053), .C2(n15874), .A(n14052), .B(n14051), .ZN(
        n16608) );
  INV_X1 U17393 ( .A(n16608), .ZN(n18922) );
  OAI211_X1 U17394 ( .C1(n14054), .C2(n18943), .A(n19137), .B(n16780), .ZN(
        n14055) );
  INV_X1 U17395 ( .A(n14055), .ZN(n16124) );
  INV_X1 U17396 ( .A(n14056), .ZN(n18952) );
  OAI211_X1 U17397 ( .C1(n18497), .C2(n18952), .A(n15984), .B(n14057), .ZN(
        n14058) );
  NOR2_X1 U17398 ( .A1(n14059), .A2(n14058), .ZN(n15873) );
  OAI211_X1 U17399 ( .C1(n14062), .C2(n15873), .A(n14061), .B(n14060), .ZN(
        n15880) );
  AOI211_X1 U17400 ( .C1(n15983), .C2(n18922), .A(n16124), .B(n15880), .ZN(
        n14063) );
  NOR2_X1 U17401 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19086), .ZN(n18481) );
  INV_X1 U17402 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18470) );
  NAND3_X1 U17403 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n19084)
         );
  NOR2_X1 U17404 ( .A1(n18470), .A2(n19084), .ZN(n14065) );
  MUX2_X1 U17405 ( .A(n14066), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n19116), .Z(P3_U3284) );
  OR2_X1 U17406 ( .A1(n14067), .A2(n15860), .ZN(n18469) );
  NOR2_X1 U17407 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18469), .ZN(n14068) );
  NAND2_X1 U17408 ( .A1(n19095), .A2(n18978), .ZN(n18143) );
  NAND2_X1 U17409 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18468) );
  INV_X1 U17410 ( .A(n18766), .ZN(n18558) );
  OAI21_X1 U17411 ( .B1(n14068), .B2(n19084), .A(n18558), .ZN(n18475) );
  INV_X1 U17412 ( .A(n18475), .ZN(n14069) );
  NAND2_X1 U17413 ( .A1(n18978), .A2(n19086), .ZN(n16782) );
  NAND2_X1 U17414 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18045) );
  INV_X1 U17415 ( .A(n18045), .ZN(n18103) );
  NOR2_X1 U17416 ( .A1(n19130), .A2(n18103), .ZN(n15853) );
  AOI21_X1 U17417 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n15853), .ZN(n15854) );
  NOR2_X1 U17418 ( .A1(n14069), .A2(n15854), .ZN(n14071) );
  INV_X1 U17419 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n19135) );
  NOR3_X1 U17420 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n19135), .ZN(n18535) );
  NOR2_X1 U17421 ( .A1(n19086), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18516) );
  OR2_X1 U17422 ( .A1(n18516), .A2(n14069), .ZN(n15852) );
  OR2_X1 U17423 ( .A1(n18535), .A2(n15852), .ZN(n14070) );
  MUX2_X1 U17424 ( .A(n14071), .B(n14070), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  INV_X1 U17425 ( .A(DATAI_12_), .ZN(n14073) );
  NAND2_X1 U17426 ( .A1(n14438), .A2(BUF1_REG_12__SCAN_IN), .ZN(n14072) );
  OAI21_X1 U17427 ( .B1(n14438), .B2(n14073), .A(n14072), .ZN(n20254) );
  AOI22_X1 U17428 ( .A1(n14503), .A2(n20254), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n14502), .ZN(n14074) );
  OAI21_X1 U17429 ( .B1(n14084), .B2(n14505), .A(n14074), .ZN(P1_U2892) );
  NAND3_X1 U17430 ( .A1(n20158), .A2(P1_REIP_REG_10__SCAN_IN), .A3(
        P1_REIP_REG_9__SCAN_IN), .ZN(n16159) );
  INV_X1 U17431 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20785) );
  OAI21_X1 U17432 ( .B1(n16159), .B2(n20785), .A(n20786), .ZN(n14082) );
  NAND3_X1 U17433 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .A3(n14075), .ZN(n14169) );
  AND2_X1 U17434 ( .A1(n20185), .A2(n14169), .ZN(n14361) );
  NOR2_X1 U17435 ( .A1(n20192), .A2(n14076), .ZN(n14077) );
  AOI211_X1 U17436 ( .C1(n20197), .C2(n16181), .A(n14077), .B(n16156), .ZN(
        n14079) );
  NAND2_X1 U17437 ( .A1(n20196), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14078) );
  OAI211_X1 U17438 ( .C1(n14080), .C2(n20193), .A(n14079), .B(n14078), .ZN(
        n14081) );
  AOI21_X1 U17439 ( .B1(n14082), .B2(n14361), .A(n14081), .ZN(n14083) );
  OAI21_X1 U17440 ( .B1(n14084), .B2(n20178), .A(n14083), .ZN(P1_U2828) );
  INV_X1 U17441 ( .A(n15245), .ZN(n14085) );
  NOR2_X1 U17442 ( .A1(n9732), .A2(n14085), .ZN(n14086) );
  NAND2_X1 U17443 ( .A1(n14088), .A2(n10861), .ZN(n14089) );
  XNOR2_X1 U17444 ( .A(n14089), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14090) );
  XNOR2_X1 U17445 ( .A(n14091), .B(n14090), .ZN(n14114) );
  XNOR2_X1 U17446 ( .A(n14094), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14103) );
  OR2_X1 U17447 ( .A1(n14103), .A2(n19429), .ZN(n14101) );
  NOR2_X1 U17448 ( .A1(n19300), .A2(n20042), .ZN(n14106) );
  AOI21_X1 U17449 ( .B1(n16477), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14106), .ZN(n14095) );
  OAI21_X1 U17450 ( .B1(n16491), .B2(n14096), .A(n14095), .ZN(n14097) );
  INV_X1 U17451 ( .A(n14097), .ZN(n14098) );
  OAI21_X1 U17452 ( .B1(n14114), .B2(n19431), .A(n14102), .ZN(P2_U2983) );
  NOR3_X1 U17453 ( .A1(n15431), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14104), .ZN(n14105) );
  AOI211_X1 U17454 ( .C1(n15117), .C2(n16582), .A(n14106), .B(n14105), .ZN(
        n14110) );
  INV_X1 U17455 ( .A(n14107), .ZN(n14108) );
  AOI22_X1 U17456 ( .A1(n14964), .A2(n16592), .B1(n14108), .B2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14109) );
  OAI21_X1 U17457 ( .B1(n14114), .B2(n16570), .A(n14113), .ZN(P2_U3015) );
  AOI22_X1 U17458 ( .A1(n14153), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n14163), .ZN(n14168) );
  AND2_X1 U17459 ( .A1(n14163), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14115) );
  AOI21_X1 U17460 ( .B1(n14153), .B2(P1_EBX_REG_30__SCAN_IN), .A(n14115), .ZN(
        n14190) );
  MUX2_X1 U17461 ( .A(n14154), .B(n14188), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n14117) );
  NOR2_X1 U17462 ( .A1(n14153), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14116) );
  NOR2_X1 U17463 ( .A1(n14117), .A2(n14116), .ZN(n14362) );
  INV_X1 U17464 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16266) );
  NAND2_X1 U17465 ( .A1(n13292), .A2(n16266), .ZN(n14119) );
  INV_X1 U17466 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n16148) );
  NAND2_X1 U17467 ( .A1(n14140), .A2(n16148), .ZN(n14118) );
  NAND3_X1 U17468 ( .A1(n14119), .A2(n14166), .A3(n14118), .ZN(n14121) );
  NAND2_X1 U17469 ( .A1(n13129), .A2(n16148), .ZN(n14120) );
  NAND2_X1 U17470 ( .A1(n14121), .A2(n14120), .ZN(n14423) );
  MUX2_X1 U17471 ( .A(n14151), .B(n14166), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n14123) );
  INV_X1 U17472 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14781) );
  NAND2_X1 U17473 ( .A1(n14164), .A2(n14781), .ZN(n14122) );
  NAND2_X1 U17474 ( .A1(n14123), .A2(n14122), .ZN(n14415) );
  NAND2_X1 U17475 ( .A1(n13292), .A2(n14124), .ZN(n14126) );
  INV_X1 U17476 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14127) );
  NAND2_X1 U17477 ( .A1(n14140), .A2(n14127), .ZN(n14125) );
  NAND3_X1 U17478 ( .A1(n14126), .A2(n14166), .A3(n14125), .ZN(n14129) );
  NAND2_X1 U17479 ( .A1(n14188), .A2(n14127), .ZN(n14128) );
  AND2_X1 U17480 ( .A1(n14129), .A2(n14128), .ZN(n14413) );
  MUX2_X1 U17481 ( .A(n14151), .B(n14166), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n14131) );
  NAND2_X1 U17482 ( .A1(n14164), .A2(n11909), .ZN(n14130) );
  NAND2_X1 U17483 ( .A1(n14131), .A2(n14130), .ZN(n14352) );
  NAND2_X1 U17484 ( .A1(n13292), .A2(n16248), .ZN(n14133) );
  INV_X1 U17485 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14403) );
  NAND2_X1 U17486 ( .A1(n14140), .A2(n14403), .ZN(n14132) );
  NAND3_X1 U17487 ( .A1(n14133), .A2(n14166), .A3(n14132), .ZN(n14135) );
  NAND2_X1 U17488 ( .A1(n13129), .A2(n14403), .ZN(n14134) );
  NAND2_X1 U17489 ( .A1(n14135), .A2(n14134), .ZN(n14336) );
  MUX2_X1 U17490 ( .A(n14151), .B(n14166), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n14137) );
  NAND2_X1 U17491 ( .A1(n14164), .A2(n14746), .ZN(n14136) );
  NAND2_X1 U17492 ( .A1(n14137), .A2(n14136), .ZN(n14323) );
  MUX2_X1 U17493 ( .A(n14188), .B(n13130), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n14139) );
  AND2_X1 U17494 ( .A1(n14163), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14138) );
  NOR2_X1 U17495 ( .A1(n14139), .A2(n14138), .ZN(n14311) );
  INV_X1 U17496 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14399) );
  NAND2_X1 U17497 ( .A1(n14154), .A2(n14399), .ZN(n14143) );
  INV_X1 U17498 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14740) );
  NAND2_X1 U17499 ( .A1(n14140), .A2(n14399), .ZN(n14141) );
  OAI211_X1 U17500 ( .C1(n13129), .C2(n14740), .A(n14141), .B(n13292), .ZN(
        n14142) );
  AND2_X1 U17501 ( .A1(n14143), .A2(n14142), .ZN(n14298) );
  INV_X1 U17502 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14729) );
  NAND2_X1 U17503 ( .A1(n13292), .A2(n14729), .ZN(n14144) );
  OAI211_X1 U17504 ( .C1(P1_EBX_REG_22__SCAN_IN), .C2(n14163), .A(n14144), .B(
        n14166), .ZN(n14147) );
  INV_X1 U17505 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14145) );
  NAND2_X1 U17506 ( .A1(n14188), .A2(n14145), .ZN(n14146) );
  AND2_X1 U17507 ( .A1(n14147), .A2(n14146), .ZN(n14283) );
  MUX2_X1 U17508 ( .A(n14151), .B(n14166), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n14148) );
  OAI21_X1 U17509 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n14153), .A(
        n14148), .ZN(n14271) );
  AOI21_X1 U17510 ( .B1(n14539), .B2(n13292), .A(n13129), .ZN(n14149) );
  OAI21_X1 U17511 ( .B1(P1_EBX_REG_24__SCAN_IN), .B2(n14163), .A(n14149), .ZN(
        n14150) );
  OAI21_X1 U17512 ( .B1(P1_EBX_REG_24__SCAN_IN), .B2(n14166), .A(n14150), .ZN(
        n14262) );
  MUX2_X1 U17513 ( .A(n14151), .B(n14166), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n14152) );
  OAI21_X1 U17514 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n14153), .A(
        n14152), .ZN(n14247) );
  MUX2_X1 U17515 ( .A(n14154), .B(n14188), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n14155) );
  AOI21_X1 U17516 ( .B1(n14164), .B2(n14156), .A(n14155), .ZN(n14223) );
  MUX2_X1 U17517 ( .A(n14166), .B(n13292), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n14158) );
  NAND2_X1 U17518 ( .A1(n14163), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14157) );
  NAND2_X1 U17519 ( .A1(n14158), .A2(n14157), .ZN(n14237) );
  INV_X1 U17520 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14162) );
  NOR2_X1 U17521 ( .A1(n14163), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n14159) );
  AOI211_X1 U17522 ( .C1(n14160), .C2(n13292), .A(n13129), .B(n14159), .ZN(
        n14161) );
  AOI21_X1 U17523 ( .B1(n14188), .B2(n14162), .A(n14161), .ZN(n14213) );
  NOR2_X1 U17524 ( .A1(n14163), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n14165) );
  AOI21_X1 U17525 ( .B1(n14164), .B2(n14682), .A(n14165), .ZN(n14187) );
  MUX2_X1 U17526 ( .A(n14187), .B(n14165), .S(n13129), .Z(n14204) );
  NAND2_X1 U17527 ( .A1(n14212), .A2(n14204), .ZN(n14203) );
  MUX2_X1 U17528 ( .A(n14190), .B(n14166), .S(n14203), .Z(n14167) );
  XOR2_X1 U17529 ( .A(n14168), .B(n14167), .Z(n14666) );
  NAND2_X1 U17530 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n14174) );
  AND2_X1 U17531 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(P1_REIP_REG_21__SCAN_IN), 
        .ZN(n14181) );
  NAND2_X1 U17532 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .ZN(n14170) );
  NOR2_X1 U17533 ( .A1(n14170), .A2(n14169), .ZN(n16134) );
  NAND4_X1 U17534 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .A4(n16134), .ZN(n14321) );
  NAND2_X1 U17535 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n14171) );
  NOR2_X1 U17536 ( .A1(n14321), .A2(n14171), .ZN(n14172) );
  NAND2_X1 U17537 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n14183) );
  INV_X1 U17538 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20873) );
  NOR2_X1 U17539 ( .A1(n14183), .A2(n20873), .ZN(n14173) );
  NAND3_X1 U17540 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .A3(n14227), .ZN(n14205) );
  OAI21_X1 U17541 ( .B1(n14174), .B2(n14205), .A(n20185), .ZN(n14197) );
  AOI22_X1 U17542 ( .A1(n20196), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B1(
        P1_EBX_REG_31__SCAN_IN), .B2(n20175), .ZN(n14175) );
  OAI21_X1 U17543 ( .B1(n21036), .B2(n14197), .A(n14175), .ZN(n14176) );
  AOI21_X1 U17544 ( .B1(n14666), .B2(n20183), .A(n14176), .ZN(n14185) );
  NAND2_X1 U17545 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n14177) );
  NAND3_X1 U17546 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n14322) );
  INV_X1 U17547 ( .A(n14322), .ZN(n14178) );
  NAND2_X1 U17548 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n14178), .ZN(n14179) );
  AND2_X1 U17549 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n14180) );
  AND2_X1 U17550 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n14182) );
  NAND4_X1 U17551 ( .A1(n14210), .A2(P1_REIP_REG_29__SCAN_IN), .A3(
        P1_REIP_REG_30__SCAN_IN), .A4(n21036), .ZN(n14184) );
  AOI21_X1 U17552 ( .B1(n14210), .B2(P1_REIP_REG_29__SCAN_IN), .A(
        P1_REIP_REG_30__SCAN_IN), .ZN(n14198) );
  NAND2_X1 U17553 ( .A1(n14387), .A2(n20151), .ZN(n14196) );
  AOI22_X1 U17554 ( .A1(n14203), .A2(n14188), .B1(n14187), .B2(n14212), .ZN(
        n14189) );
  XOR2_X1 U17555 ( .A(n14190), .B(n14189), .Z(n14675) );
  INV_X1 U17556 ( .A(n14191), .ZN(n14193) );
  AOI22_X1 U17557 ( .A1(n20196), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(n20175), .ZN(n14192) );
  OAI21_X1 U17558 ( .B1(n20189), .B2(n14193), .A(n14192), .ZN(n14194) );
  AOI21_X1 U17559 ( .B1(n14675), .B2(n20183), .A(n14194), .ZN(n14195) );
  OAI211_X1 U17560 ( .C1(n14198), .C2(n14197), .A(n14196), .B(n14195), .ZN(
        P1_U2810) );
  INV_X1 U17561 ( .A(n14199), .ZN(n14201) );
  INV_X1 U17562 ( .A(n14202), .ZN(n14510) );
  INV_X1 U17563 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20917) );
  OAI21_X1 U17564 ( .B1(n14212), .B2(n14204), .A(n14203), .ZN(n14678) );
  NOR2_X1 U17565 ( .A1(n14678), .A2(n20193), .ZN(n14209) );
  NAND2_X1 U17566 ( .A1(n20185), .A2(n14205), .ZN(n14218) );
  AOI22_X1 U17567 ( .A1(n20196), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B1(
        n20175), .B2(P1_EBX_REG_29__SCAN_IN), .ZN(n14207) );
  NAND2_X1 U17568 ( .A1(n20197), .A2(n14513), .ZN(n14206) );
  OAI211_X1 U17569 ( .C1(n14218), .C2(n20917), .A(n14207), .B(n14206), .ZN(
        n14208) );
  AOI211_X1 U17570 ( .C1(n14210), .C2(n20917), .A(n14209), .B(n14208), .ZN(
        n14211) );
  OAI21_X1 U17571 ( .B1(n14202), .B2(n20178), .A(n14211), .ZN(P1_U2811) );
  AOI21_X1 U17572 ( .B1(n14213), .B2(n14222), .A(n14212), .ZN(n14693) );
  AOI22_X1 U17573 ( .A1(n20196), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B1(
        n20175), .B2(P1_EBX_REG_28__SCAN_IN), .ZN(n14217) );
  INV_X1 U17574 ( .A(n14214), .ZN(n14215) );
  NAND2_X1 U17575 ( .A1(n20197), .A2(n14215), .ZN(n14216) );
  OAI211_X1 U17576 ( .C1(n14218), .C2(n21005), .A(n14217), .B(n14216), .ZN(
        n14220) );
  NOR3_X1 U17577 ( .A1(n14231), .A2(P1_REIP_REG_28__SCAN_IN), .A3(n20887), 
        .ZN(n14219) );
  AOI211_X1 U17578 ( .C1(n14693), .C2(n20183), .A(n14220), .B(n14219), .ZN(
        n14221) );
  OAI21_X1 U17579 ( .B1(n14444), .B2(n20178), .A(n14221), .ZN(P1_U2812) );
  INV_X1 U17580 ( .A(n14222), .ZN(n14225) );
  AOI21_X1 U17581 ( .B1(n9690), .B2(n14237), .A(n14223), .ZN(n14224) );
  NOR2_X1 U17582 ( .A1(n14225), .A2(n14224), .ZN(n14702) );
  INV_X1 U17583 ( .A(n14226), .ZN(n14230) );
  NOR2_X1 U17584 ( .A1(n20161), .A2(n14227), .ZN(n14238) );
  NAND2_X1 U17585 ( .A1(n14238), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14229) );
  AOI22_X1 U17586 ( .A1(n20196), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B1(
        n20175), .B2(P1_EBX_REG_27__SCAN_IN), .ZN(n14228) );
  OAI211_X1 U17587 ( .C1(n20189), .C2(n14230), .A(n14229), .B(n14228), .ZN(
        n14233) );
  NOR2_X1 U17588 ( .A1(n14231), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14232) );
  AOI211_X1 U17589 ( .C1(n20183), .C2(n14702), .A(n14233), .B(n14232), .ZN(
        n14234) );
  OAI21_X1 U17590 ( .B1(n14447), .B2(n20178), .A(n14234), .ZN(P1_U2813) );
  AOI21_X1 U17591 ( .B1(n14236), .B2(n14235), .A(n9686), .ZN(n14523) );
  INV_X1 U17592 ( .A(n14523), .ZN(n14451) );
  XNOR2_X1 U17593 ( .A(n9690), .B(n14237), .ZN(n14392) );
  INV_X1 U17594 ( .A(n14392), .ZN(n16214) );
  NAND2_X1 U17595 ( .A1(n14238), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14240) );
  AOI22_X1 U17596 ( .A1(n20196), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(
        n20175), .B2(P1_EBX_REG_26__SCAN_IN), .ZN(n14239) );
  OAI211_X1 U17597 ( .C1(n20189), .C2(n14519), .A(n14240), .B(n14239), .ZN(
        n14242) );
  INV_X1 U17598 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20809) );
  NOR3_X1 U17599 ( .A1(n14250), .A2(P1_REIP_REG_26__SCAN_IN), .A3(n20809), 
        .ZN(n14241) );
  AOI211_X1 U17600 ( .C1(n20183), .C2(n16214), .A(n14242), .B(n14241), .ZN(
        n14243) );
  OAI21_X1 U17601 ( .B1(n14451), .B2(n20178), .A(n14243), .ZN(P1_U2814) );
  INV_X1 U17602 ( .A(n14235), .ZN(n14245) );
  AOI21_X1 U17603 ( .B1(n14246), .B2(n14244), .A(n14245), .ZN(n14530) );
  INV_X1 U17604 ( .A(n14530), .ZN(n14454) );
  AOI21_X1 U17605 ( .B1(n14247), .B2(n14261), .A(n9690), .ZN(n14711) );
  INV_X1 U17606 ( .A(n14533), .ZN(n14249) );
  AOI22_X1 U17607 ( .A1(n20196), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B1(
        n20175), .B2(P1_EBX_REG_25__SCAN_IN), .ZN(n14248) );
  OAI21_X1 U17608 ( .B1(n20189), .B2(n14249), .A(n14248), .ZN(n14252) );
  NOR2_X1 U17609 ( .A1(n14250), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14251) );
  AOI211_X1 U17610 ( .C1(n14711), .C2(n20183), .A(n14252), .B(n14251), .ZN(
        n14257) );
  INV_X1 U17611 ( .A(n14277), .ZN(n14253) );
  INV_X1 U17612 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20806) );
  NOR3_X1 U17613 ( .A1(n14253), .A2(P1_REIP_REG_24__SCAN_IN), .A3(n20806), 
        .ZN(n14265) );
  INV_X1 U17614 ( .A(n14254), .ZN(n14255) );
  AND2_X1 U17615 ( .A1(n20185), .A2(n14255), .ZN(n14276) );
  OAI21_X1 U17616 ( .B1(n14265), .B2(n14276), .A(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n14256) );
  OAI211_X1 U17617 ( .C1(n14454), .C2(n20178), .A(n14257), .B(n14256), .ZN(
        P1_U2815) );
  BUF_X1 U17618 ( .A(n14258), .Z(n14259) );
  OAI21_X1 U17619 ( .B1(n14259), .B2(n14260), .A(n14244), .ZN(n14541) );
  OAI21_X1 U17620 ( .B1(n14272), .B2(n14262), .A(n14261), .ZN(n14395) );
  INV_X1 U17621 ( .A(n14395), .ZN(n14722) );
  AOI22_X1 U17622 ( .A1(n20196), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        n20175), .B2(P1_EBX_REG_24__SCAN_IN), .ZN(n14264) );
  NAND2_X1 U17623 ( .A1(n14276), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14263) );
  OAI211_X1 U17624 ( .C1(n20189), .C2(n14542), .A(n14264), .B(n14263), .ZN(
        n14266) );
  AOI211_X1 U17625 ( .C1(n14722), .C2(n20183), .A(n14266), .B(n14265), .ZN(
        n14267) );
  OAI21_X1 U17626 ( .B1(n14541), .B2(n20178), .A(n14267), .ZN(P1_U2816) );
  INV_X1 U17627 ( .A(n14259), .ZN(n14269) );
  OAI21_X1 U17628 ( .B1(n14270), .B2(n14268), .A(n14269), .ZN(n14552) );
  INV_X1 U17629 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14397) );
  OAI22_X1 U17630 ( .A1(n20177), .A2(n14550), .B1(n20192), .B2(n14397), .ZN(
        n14275) );
  AND2_X1 U17631 ( .A1(n14285), .A2(n14271), .ZN(n14273) );
  OR2_X1 U17632 ( .A1(n14273), .A2(n14272), .ZN(n16224) );
  NOR2_X1 U17633 ( .A1(n16224), .A2(n20193), .ZN(n14274) );
  AOI211_X1 U17634 ( .C1(n20197), .C2(n14555), .A(n14275), .B(n14274), .ZN(
        n14279) );
  OAI21_X1 U17635 ( .B1(n14277), .B2(P1_REIP_REG_23__SCAN_IN), .A(n14276), 
        .ZN(n14278) );
  OAI211_X1 U17636 ( .C1(n14552), .C2(n20178), .A(n14279), .B(n14278), .ZN(
        P1_U2817) );
  INV_X1 U17637 ( .A(n14305), .ZN(n14294) );
  XNOR2_X1 U17638 ( .A(P1_REIP_REG_22__SCAN_IN), .B(P1_REIP_REG_21__SCAN_IN), 
        .ZN(n14293) );
  AOI21_X1 U17639 ( .B1(n14282), .B2(n14281), .A(n14268), .ZN(n14560) );
  NAND2_X1 U17640 ( .A1(n14560), .A2(n20151), .ZN(n14292) );
  NAND2_X1 U17641 ( .A1(n14300), .A2(n14283), .ZN(n14284) );
  AND2_X1 U17642 ( .A1(n14285), .A2(n14284), .ZN(n14726) );
  INV_X1 U17643 ( .A(n14286), .ZN(n14287) );
  NAND2_X1 U17644 ( .A1(n20185), .A2(n14287), .ZN(n14317) );
  INV_X1 U17645 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20859) );
  AOI22_X1 U17646 ( .A1(n20196), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n20175), .B2(P1_EBX_REG_22__SCAN_IN), .ZN(n14289) );
  NAND2_X1 U17647 ( .A1(n20197), .A2(n14563), .ZN(n14288) );
  OAI211_X1 U17648 ( .C1(n14317), .C2(n20859), .A(n14289), .B(n14288), .ZN(
        n14290) );
  AOI21_X1 U17649 ( .B1(n14726), .B2(n20183), .A(n14290), .ZN(n14291) );
  OAI211_X1 U17650 ( .C1(n14294), .C2(n14293), .A(n14292), .B(n14291), .ZN(
        P1_U2818) );
  INV_X1 U17651 ( .A(n14281), .ZN(n14296) );
  AOI21_X1 U17652 ( .B1(n14297), .B2(n14295), .A(n14296), .ZN(n14573) );
  INV_X1 U17653 ( .A(n14573), .ZN(n14467) );
  INV_X1 U17654 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20802) );
  OR2_X1 U17655 ( .A1(n9770), .A2(n14298), .ZN(n14299) );
  NAND2_X1 U17656 ( .A1(n14300), .A2(n14299), .ZN(n14738) );
  AOI22_X1 U17657 ( .A1(n20196), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n20175), .B2(P1_EBX_REG_21__SCAN_IN), .ZN(n14301) );
  OAI21_X1 U17658 ( .B1(n20802), .B2(n14317), .A(n14301), .ZN(n14302) );
  AOI21_X1 U17659 ( .B1(n20197), .B2(n14569), .A(n14302), .ZN(n14303) );
  OAI21_X1 U17660 ( .B1(n14738), .B2(n20193), .A(n14303), .ZN(n14304) );
  AOI21_X1 U17661 ( .B1(n14305), .B2(n20802), .A(n14304), .ZN(n14306) );
  OAI21_X1 U17662 ( .B1(n14467), .B2(n20178), .A(n14306), .ZN(P1_U2819) );
  AOI21_X1 U17663 ( .B1(n14331), .B2(P1_REIP_REG_19__SCAN_IN), .A(
        P1_REIP_REG_20__SCAN_IN), .ZN(n14318) );
  INV_X1 U17664 ( .A(n14295), .ZN(n14308) );
  AOI21_X1 U17665 ( .B1(n14309), .B2(n14307), .A(n14308), .ZN(n14578) );
  NAND2_X1 U17666 ( .A1(n14578), .A2(n20151), .ZN(n14316) );
  INV_X1 U17667 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n14579) );
  INV_X1 U17668 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14310) );
  OAI22_X1 U17669 ( .A1(n20177), .A2(n14579), .B1(n14310), .B2(n20192), .ZN(
        n14314) );
  AND2_X1 U17670 ( .A1(n14325), .A2(n14311), .ZN(n14312) );
  OR2_X1 U17671 ( .A1(n14312), .A2(n9770), .ZN(n14744) );
  NOR2_X1 U17672 ( .A1(n14744), .A2(n20193), .ZN(n14313) );
  AOI211_X1 U17673 ( .C1(n20197), .C2(n14581), .A(n14314), .B(n14313), .ZN(
        n14315) );
  OAI211_X1 U17674 ( .C1(n14318), .C2(n14317), .A(n14316), .B(n14315), .ZN(
        P1_U2820) );
  OAI21_X1 U17675 ( .B1(n14319), .B2(n14320), .A(n14307), .ZN(n14586) );
  NAND2_X1 U17676 ( .A1(n20185), .A2(n14321), .ZN(n14355) );
  OR3_X1 U17677 ( .A1(n16146), .A2(n14322), .A3(P1_REIP_REG_18__SCAN_IN), .ZN(
        n14345) );
  INV_X1 U17678 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20800) );
  AOI21_X1 U17679 ( .B1(n14355), .B2(n14345), .A(n20800), .ZN(n14330) );
  NAND2_X1 U17680 ( .A1(n14337), .A2(n14323), .ZN(n14324) );
  NAND2_X1 U17681 ( .A1(n14325), .A2(n14324), .ZN(n16232) );
  INV_X1 U17682 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14402) );
  OAI22_X1 U17683 ( .A1(n16232), .A2(n20193), .B1(n20192), .B2(n14402), .ZN(
        n14326) );
  INV_X1 U17684 ( .A(n14326), .ZN(n14327) );
  OAI211_X1 U17685 ( .C1(n20177), .C2(n14328), .A(n14327), .B(n20191), .ZN(
        n14329) );
  AOI211_X1 U17686 ( .C1(n20197), .C2(n14587), .A(n14330), .B(n14329), .ZN(
        n14333) );
  NAND2_X1 U17687 ( .A1(n14331), .A2(n20800), .ZN(n14332) );
  OAI211_X1 U17688 ( .C1(n14586), .C2(n20178), .A(n14333), .B(n14332), .ZN(
        P1_U2821) );
  AOI21_X1 U17689 ( .B1(n14335), .B2(n14334), .A(n14319), .ZN(n14601) );
  INV_X1 U17690 ( .A(n14601), .ZN(n14478) );
  OR2_X1 U17691 ( .A1(n14351), .A2(n14336), .ZN(n14338) );
  AND2_X1 U17692 ( .A1(n14338), .A2(n14337), .ZN(n16241) );
  INV_X1 U17693 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20798) );
  NAND2_X1 U17694 ( .A1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n20196), .ZN(
        n14339) );
  NAND2_X1 U17695 ( .A1(n20191), .A2(n14339), .ZN(n14340) );
  AOI21_X1 U17696 ( .B1(n20175), .B2(P1_EBX_REG_18__SCAN_IN), .A(n14340), .ZN(
        n14343) );
  INV_X1 U17697 ( .A(n14596), .ZN(n14341) );
  NAND2_X1 U17698 ( .A1(n20197), .A2(n14341), .ZN(n14342) );
  OAI211_X1 U17699 ( .C1(n14355), .C2(n20798), .A(n14343), .B(n14342), .ZN(
        n14344) );
  AOI21_X1 U17700 ( .B1(n16241), .B2(n20183), .A(n14344), .ZN(n14346) );
  OAI211_X1 U17701 ( .C1(n14478), .C2(n20178), .A(n14346), .B(n14345), .ZN(
        P1_U2822) );
  NAND2_X1 U17702 ( .A1(n14348), .A2(n14349), .ZN(n14350) );
  AND2_X1 U17703 ( .A1(n14334), .A2(n14350), .ZN(n14613) );
  AOI21_X1 U17704 ( .B1(n14352), .B2(n14411), .A(n14351), .ZN(n16251) );
  AOI21_X1 U17705 ( .B1(n20175), .B2(P1_EBX_REG_17__SCAN_IN), .A(n20174), .ZN(
        n14354) );
  NAND2_X1 U17706 ( .A1(n20196), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14353) );
  OAI211_X1 U17707 ( .C1(n20189), .C2(n14611), .A(n14354), .B(n14353), .ZN(
        n14357) );
  INV_X1 U17708 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20795) );
  NAND2_X1 U17709 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n16128) );
  AOI221_X1 U17710 ( .B1(n16146), .B2(n20795), .C1(n16128), .C2(n20795), .A(
        n14355), .ZN(n14356) );
  AOI211_X1 U17711 ( .C1(n16251), .C2(n20183), .A(n14357), .B(n14356), .ZN(
        n14358) );
  OAI21_X1 U17712 ( .B1(n14487), .B2(n20178), .A(n14358), .ZN(P1_U2823) );
  AOI21_X1 U17713 ( .B1(n14360), .B2(n13929), .A(n14359), .ZN(n14624) );
  INV_X1 U17714 ( .A(n14624), .ZN(n14506) );
  INV_X1 U17715 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20789) );
  AOI22_X1 U17716 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n14361), .B1(n16147), 
        .B2(n20789), .ZN(n14370) );
  INV_X1 U17717 ( .A(n14362), .ZN(n14365) );
  INV_X1 U17718 ( .A(n14363), .ZN(n14364) );
  AOI21_X1 U17719 ( .B1(n14365), .B2(n14364), .A(n14424), .ZN(n16269) );
  NOR2_X1 U17720 ( .A1(n20177), .A2(n14621), .ZN(n14366) );
  AOI211_X1 U17721 ( .C1(n20175), .C2(P1_EBX_REG_13__SCAN_IN), .A(n20174), .B(
        n14366), .ZN(n14367) );
  OAI21_X1 U17722 ( .B1(n14620), .B2(n20189), .A(n14367), .ZN(n14368) );
  AOI21_X1 U17723 ( .B1(n16269), .B2(n20183), .A(n14368), .ZN(n14369) );
  OAI211_X1 U17724 ( .C1(n14506), .C2(n20178), .A(n14370), .B(n14369), .ZN(
        P1_U2827) );
  OAI22_X1 U17725 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n14372), .B1(n20192), 
        .B2(n14371), .ZN(n14375) );
  NOR2_X1 U17726 ( .A1(n20189), .A2(n14373), .ZN(n14374) );
  AOI211_X1 U17727 ( .C1(n20196), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n14375), .B(n14374), .ZN(n14376) );
  OAI21_X1 U17728 ( .B1(n20193), .B2(n14377), .A(n14376), .ZN(n14380) );
  NOR3_X1 U17729 ( .A1(n14378), .A2(n20161), .A3(n20771), .ZN(n14379) );
  AOI211_X1 U17730 ( .C1(n14381), .C2(n20467), .A(n14380), .B(n14379), .ZN(
        n14382) );
  OAI21_X1 U17731 ( .B1(n14384), .B2(n14383), .A(n14382), .ZN(P1_U2837) );
  INV_X1 U17732 ( .A(n14666), .ZN(n14386) );
  OAI22_X1 U17733 ( .A1(n14386), .A2(n20209), .B1(n14385), .B2(n20216), .ZN(
        P1_U2841) );
  INV_X1 U17734 ( .A(n14387), .ZN(n14436) );
  AOI22_X1 U17735 ( .A1(n14675), .A2(n14430), .B1(P1_EBX_REG_30__SCAN_IN), 
        .B2(n14429), .ZN(n14388) );
  OAI21_X1 U17736 ( .B1(n14436), .B2(n14420), .A(n14388), .ZN(P1_U2842) );
  INV_X1 U17737 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14389) );
  OAI222_X1 U17738 ( .A1(n14389), .A2(n20216), .B1(n20209), .B2(n14678), .C1(
        n14202), .C2(n14420), .ZN(P1_U2843) );
  AOI22_X1 U17739 ( .A1(n14693), .A2(n14430), .B1(n14429), .B2(
        P1_EBX_REG_28__SCAN_IN), .ZN(n14390) );
  OAI21_X1 U17740 ( .B1(n14444), .B2(n14420), .A(n14390), .ZN(P1_U2844) );
  AOI22_X1 U17741 ( .A1(n14702), .A2(n14430), .B1(n14429), .B2(
        P1_EBX_REG_27__SCAN_IN), .ZN(n14391) );
  OAI21_X1 U17742 ( .B1(n14447), .B2(n14420), .A(n14391), .ZN(P1_U2845) );
  INV_X1 U17743 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14393) );
  OAI222_X1 U17744 ( .A1(n14393), .A2(n20216), .B1(n20209), .B2(n14392), .C1(
        n14420), .C2(n14451), .ZN(P1_U2846) );
  AOI22_X1 U17745 ( .A1(n14711), .A2(n14430), .B1(n14429), .B2(
        P1_EBX_REG_25__SCAN_IN), .ZN(n14394) );
  OAI21_X1 U17746 ( .B1(n14454), .B2(n14420), .A(n14394), .ZN(P1_U2847) );
  INV_X1 U17747 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14396) );
  OAI222_X1 U17748 ( .A1(n14396), .A2(n20216), .B1(n20209), .B2(n14395), .C1(
        n14541), .C2(n14420), .ZN(P1_U2848) );
  OAI222_X1 U17749 ( .A1(n16224), .A2(n20209), .B1(n14397), .B2(n20216), .C1(
        n14552), .C2(n14420), .ZN(P1_U2849) );
  INV_X1 U17750 ( .A(n14560), .ZN(n14463) );
  AOI22_X1 U17751 ( .A1(n14726), .A2(n14430), .B1(n14429), .B2(
        P1_EBX_REG_22__SCAN_IN), .ZN(n14398) );
  OAI21_X1 U17752 ( .B1(n14463), .B2(n14420), .A(n14398), .ZN(P1_U2850) );
  OAI22_X1 U17753 ( .A1(n14738), .A2(n20209), .B1(n14399), .B2(n20216), .ZN(
        n14400) );
  AOI21_X1 U17754 ( .B1(n14573), .B2(n20212), .A(n14400), .ZN(n14401) );
  INV_X1 U17755 ( .A(n14401), .ZN(P1_U2851) );
  INV_X1 U17756 ( .A(n14578), .ZN(n14471) );
  OAI222_X1 U17757 ( .A1(n14744), .A2(n20209), .B1(n20216), .B2(n14310), .C1(
        n14420), .C2(n14471), .ZN(P1_U2852) );
  OAI222_X1 U17758 ( .A1(n16232), .A2(n20209), .B1(n14402), .B2(n20216), .C1(
        n14586), .C2(n14420), .ZN(P1_U2853) );
  NOR2_X1 U17759 ( .A1(n20216), .A2(n14403), .ZN(n14404) );
  AOI21_X1 U17760 ( .B1(n16241), .B2(n14430), .A(n14404), .ZN(n14405) );
  OAI21_X1 U17761 ( .B1(n14478), .B2(n14420), .A(n14405), .ZN(P1_U2854) );
  AOI22_X1 U17762 ( .A1(n16251), .A2(n14430), .B1(n14429), .B2(
        P1_EBX_REG_17__SCAN_IN), .ZN(n14406) );
  OAI21_X1 U17763 ( .B1(n14487), .B2(n14420), .A(n14406), .ZN(P1_U2855) );
  INV_X1 U17764 ( .A(n14418), .ZN(n14408) );
  NAND2_X1 U17765 ( .A1(n14407), .A2(n14408), .ZN(n14409) );
  AOI21_X1 U17766 ( .B1(n14410), .B2(n14409), .A(n11548), .ZN(n16161) );
  INV_X1 U17767 ( .A(n16161), .ZN(n14494) );
  INV_X1 U17768 ( .A(n14411), .ZN(n14412) );
  AOI21_X1 U17769 ( .B1(n14413), .B2(n14417), .A(n14412), .ZN(n16133) );
  AOI22_X1 U17770 ( .A1(n16133), .A2(n14430), .B1(n14429), .B2(
        P1_EBX_REG_16__SCAN_IN), .ZN(n14414) );
  OAI21_X1 U17771 ( .B1(n14494), .B2(n14420), .A(n14414), .ZN(P1_U2856) );
  NAND2_X1 U17772 ( .A1(n14426), .A2(n14415), .ZN(n14416) );
  NAND2_X1 U17773 ( .A1(n14417), .A2(n14416), .ZN(n16138) );
  XNOR2_X1 U17774 ( .A(n14407), .B(n14418), .ZN(n16166) );
  INV_X1 U17775 ( .A(n16166), .ZN(n14497) );
  INV_X1 U17776 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14419) );
  OAI222_X1 U17777 ( .A1(n16138), .A2(n20209), .B1(n14420), .B2(n14497), .C1(
        n20216), .C2(n14419), .ZN(P1_U2857) );
  INV_X1 U17778 ( .A(n14359), .ZN(n14422) );
  AOI21_X1 U17779 ( .B1(n10258), .B2(n14422), .A(n14407), .ZN(n16178) );
  OR2_X1 U17780 ( .A1(n14424), .A2(n14423), .ZN(n14425) );
  NAND2_X1 U17781 ( .A1(n14426), .A2(n14425), .ZN(n16258) );
  OAI22_X1 U17782 ( .A1(n16258), .A2(n20209), .B1(n16148), .B2(n20216), .ZN(
        n14427) );
  AOI21_X1 U17783 ( .B1(n16178), .B2(n20212), .A(n14427), .ZN(n14428) );
  INV_X1 U17784 ( .A(n14428), .ZN(P1_U2858) );
  AOI22_X1 U17785 ( .A1(n16269), .A2(n14430), .B1(n14429), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14431) );
  OAI21_X1 U17786 ( .B1(n14506), .B2(n14420), .A(n14431), .ZN(P1_U2859) );
  NOR2_X1 U17787 ( .A1(n14437), .A2(n16682), .ZN(n14434) );
  INV_X1 U17788 ( .A(n14491), .ZN(n14483) );
  INV_X1 U17789 ( .A(DATAI_14_), .ZN(n21034) );
  MUX2_X1 U17790 ( .A(n21034), .B(n16708), .S(n14438), .Z(n20258) );
  NAND3_X1 U17791 ( .A1(n14498), .A2(n14432), .A3(n11306), .ZN(n14481) );
  OAI22_X1 U17792 ( .A1(n14483), .A2(n21009), .B1(n20258), .B2(n14481), .ZN(
        n14433) );
  AOI211_X1 U17793 ( .C1(n14502), .C2(P1_EAX_REG_30__SCAN_IN), .A(n14434), .B(
        n14433), .ZN(n14435) );
  OAI21_X1 U17794 ( .B1(n14436), .B2(n14505), .A(n14435), .ZN(P1_U2874) );
  AOI22_X1 U17795 ( .A1(n14488), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n14502), .ZN(n14441) );
  INV_X1 U17796 ( .A(DATAI_13_), .ZN(n20989) );
  NAND2_X1 U17797 ( .A1(n14438), .A2(BUF1_REG_13__SCAN_IN), .ZN(n14439) );
  OAI21_X1 U17798 ( .B1(n14438), .B2(n20989), .A(n14439), .ZN(n20256) );
  AOI22_X1 U17799 ( .A1(n14491), .A2(DATAI_29_), .B1(n14490), .B2(n20256), 
        .ZN(n14440) );
  OAI211_X1 U17800 ( .C1(n14202), .C2(n14505), .A(n14441), .B(n14440), .ZN(
        P1_U2875) );
  AOI22_X1 U17801 ( .A1(n14488), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n14502), .ZN(n14443) );
  AOI22_X1 U17802 ( .A1(n14491), .A2(DATAI_28_), .B1(n14490), .B2(n20254), 
        .ZN(n14442) );
  OAI211_X1 U17803 ( .C1(n14444), .C2(n14505), .A(n14443), .B(n14442), .ZN(
        P1_U2876) );
  AOI22_X1 U17804 ( .A1(n14488), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n14502), .ZN(n14446) );
  AOI22_X1 U17805 ( .A1(n14491), .A2(DATAI_27_), .B1(n14490), .B2(n20252), 
        .ZN(n14445) );
  OAI211_X1 U17806 ( .C1(n14447), .C2(n14505), .A(n14446), .B(n14445), .ZN(
        P1_U2877) );
  AOI22_X1 U17807 ( .A1(n14488), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n14502), .ZN(n14450) );
  AOI22_X1 U17808 ( .A1(n14491), .A2(DATAI_26_), .B1(n14490), .B2(n14448), 
        .ZN(n14449) );
  OAI211_X1 U17809 ( .C1(n14451), .C2(n14505), .A(n14450), .B(n14449), .ZN(
        P1_U2878) );
  AOI22_X1 U17810 ( .A1(n14488), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n14502), .ZN(n14453) );
  AOI22_X1 U17811 ( .A1(n14491), .A2(DATAI_25_), .B1(n14490), .B2(n20250), 
        .ZN(n14452) );
  OAI211_X1 U17812 ( .C1(n14454), .C2(n14505), .A(n14453), .B(n14452), .ZN(
        P1_U2879) );
  AOI22_X1 U17813 ( .A1(n14488), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n14502), .ZN(n14456) );
  AOI22_X1 U17814 ( .A1(n14491), .A2(DATAI_24_), .B1(n14490), .B2(n20248), 
        .ZN(n14455) );
  OAI211_X1 U17815 ( .C1(n14541), .C2(n14505), .A(n14456), .B(n14455), .ZN(
        P1_U2880) );
  AOI22_X1 U17816 ( .A1(n14488), .A2(BUF1_REG_23__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n14502), .ZN(n14459) );
  AOI22_X1 U17817 ( .A1(n14491), .A2(DATAI_23_), .B1(n14490), .B2(n14457), 
        .ZN(n14458) );
  OAI211_X1 U17818 ( .C1(n14552), .C2(n14505), .A(n14459), .B(n14458), .ZN(
        P1_U2881) );
  AOI22_X1 U17819 ( .A1(n14488), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n14502), .ZN(n14462) );
  AOI22_X1 U17820 ( .A1(n14491), .A2(DATAI_22_), .B1(n14490), .B2(n14460), 
        .ZN(n14461) );
  OAI211_X1 U17821 ( .C1(n14463), .C2(n14505), .A(n14462), .B(n14461), .ZN(
        P1_U2882) );
  AOI22_X1 U17822 ( .A1(n14488), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n14502), .ZN(n14466) );
  AOI22_X1 U17823 ( .A1(n14491), .A2(DATAI_21_), .B1(n14490), .B2(n14464), 
        .ZN(n14465) );
  OAI211_X1 U17824 ( .C1(n14467), .C2(n14505), .A(n14466), .B(n14465), .ZN(
        P1_U2883) );
  AOI22_X1 U17825 ( .A1(n14488), .A2(BUF1_REG_20__SCAN_IN), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(n14502), .ZN(n14470) );
  AOI22_X1 U17826 ( .A1(n14491), .A2(DATAI_20_), .B1(n14490), .B2(n14468), 
        .ZN(n14469) );
  OAI211_X1 U17827 ( .C1(n14471), .C2(n14505), .A(n14470), .B(n14469), .ZN(
        P1_U2884) );
  AOI22_X1 U17828 ( .A1(n14488), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n14502), .ZN(n14474) );
  AOI22_X1 U17829 ( .A1(n14491), .A2(DATAI_19_), .B1(n14490), .B2(n14472), 
        .ZN(n14473) );
  OAI211_X1 U17830 ( .C1(n14586), .C2(n14505), .A(n14474), .B(n14473), .ZN(
        P1_U2885) );
  AOI22_X1 U17831 ( .A1(n14488), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n14502), .ZN(n14477) );
  AOI22_X1 U17832 ( .A1(n14491), .A2(DATAI_18_), .B1(n14490), .B2(n14475), 
        .ZN(n14476) );
  OAI211_X1 U17833 ( .C1(n14478), .C2(n14505), .A(n14477), .B(n14476), .ZN(
        P1_U2886) );
  NOR2_X1 U17834 ( .A1(n14498), .A2(n14479), .ZN(n14485) );
  INV_X1 U17835 ( .A(DATAI_17_), .ZN(n14482) );
  OAI22_X1 U17836 ( .A1(n14483), .A2(n14482), .B1(n14481), .B2(n14480), .ZN(
        n14484) );
  AOI211_X1 U17837 ( .C1(BUF1_REG_17__SCAN_IN), .C2(n14488), .A(n14485), .B(
        n14484), .ZN(n14486) );
  OAI21_X1 U17838 ( .B1(n14487), .B2(n14505), .A(n14486), .ZN(P1_U2887) );
  AOI22_X1 U17839 ( .A1(n14488), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n14502), .ZN(n14493) );
  AOI22_X1 U17840 ( .A1(n14491), .A2(DATAI_16_), .B1(n14490), .B2(n14489), 
        .ZN(n14492) );
  OAI211_X1 U17841 ( .C1(n14494), .C2(n14505), .A(n14493), .B(n14492), .ZN(
        P1_U2888) );
  OAI222_X1 U17842 ( .A1(n14505), .A2(n14497), .B1(n14500), .B2(n14496), .C1(
        n14498), .C2(n14495), .ZN(P1_U2889) );
  INV_X1 U17843 ( .A(n16178), .ZN(n14501) );
  INV_X1 U17844 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14499) );
  OAI222_X1 U17845 ( .A1(n14501), .A2(n14505), .B1(n14500), .B2(n20258), .C1(
        n14499), .C2(n14498), .ZN(P1_U2890) );
  AOI22_X1 U17846 ( .A1(n14503), .A2(n20256), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n14502), .ZN(n14504) );
  OAI21_X1 U17847 ( .B1(n14506), .B2(n14505), .A(n14504), .ZN(P1_U2891) );
  MUX2_X1 U17848 ( .A(n14508), .B(n16173), .S(n14507), .Z(n14509) );
  XNOR2_X1 U17849 ( .A(n14509), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14687) );
  NAND2_X1 U17850 ( .A1(n14510), .A2(n16205), .ZN(n14515) );
  OR2_X1 U17851 ( .A1(n14779), .A2(n20917), .ZN(n14681) );
  OAI21_X1 U17852 ( .B1(n16209), .B2(n14511), .A(n14681), .ZN(n14512) );
  AOI21_X1 U17853 ( .B1(n16204), .B2(n14513), .A(n14512), .ZN(n14514) );
  OAI211_X1 U17854 ( .C1(n20135), .C2(n14687), .A(n14515), .B(n14514), .ZN(
        P1_U2970) );
  OAI21_X1 U17855 ( .B1(n14536), .B2(n14647), .A(n16173), .ZN(n14516) );
  NAND2_X1 U17856 ( .A1(n14517), .A2(n14516), .ZN(n14518) );
  XOR2_X1 U17857 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n14518), .Z(
        n16213) );
  NOR2_X1 U17858 ( .A1(n16202), .A2(n14519), .ZN(n14522) );
  INV_X1 U17859 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20811) );
  OAI22_X1 U17860 ( .A1(n16209), .A2(n14520), .B1(n14779), .B2(n20811), .ZN(
        n14521) );
  AOI211_X1 U17861 ( .C1(n14523), .C2(n16205), .A(n14522), .B(n14521), .ZN(
        n14524) );
  OAI21_X1 U17862 ( .B1(n20135), .B2(n16213), .A(n14524), .ZN(P1_U2973) );
  MUX2_X1 U17863 ( .A(n14539), .B(n14525), .S(n16174), .Z(n14528) );
  NAND2_X1 U17864 ( .A1(n14526), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14537) );
  AND2_X1 U17865 ( .A1(n14537), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14527) );
  NOR2_X1 U17866 ( .A1(n14528), .A2(n14527), .ZN(n14529) );
  XNOR2_X1 U17867 ( .A(n14529), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14713) );
  NAND2_X1 U17868 ( .A1(n14530), .A2(n16205), .ZN(n14535) );
  OR2_X1 U17869 ( .A1(n14779), .A2(n20809), .ZN(n14708) );
  OAI21_X1 U17870 ( .B1(n16209), .B2(n14531), .A(n14708), .ZN(n14532) );
  AOI21_X1 U17871 ( .B1(n16204), .B2(n14533), .A(n14532), .ZN(n14534) );
  OAI211_X1 U17872 ( .C1(n14713), .C2(n20135), .A(n14535), .B(n14534), .ZN(
        P1_U2974) );
  NAND2_X1 U17873 ( .A1(n14536), .A2(n16174), .ZN(n14538) );
  MUX2_X1 U17874 ( .A(n16174), .B(n14538), .S(n14537), .Z(n14540) );
  XNOR2_X1 U17875 ( .A(n14540), .B(n14539), .ZN(n14724) );
  INV_X1 U17876 ( .A(n14541), .ZN(n14546) );
  NOR2_X1 U17877 ( .A1(n16202), .A2(n14542), .ZN(n14545) );
  OR2_X1 U17878 ( .A1(n14779), .A2(n20873), .ZN(n14719) );
  OAI21_X1 U17879 ( .B1(n16209), .B2(n14543), .A(n14719), .ZN(n14544) );
  OAI21_X1 U17880 ( .B1(n14724), .B2(n20135), .A(n14547), .ZN(P1_U2975) );
  XNOR2_X1 U17881 ( .A(n16174), .B(n11915), .ZN(n14548) );
  XNOR2_X1 U17882 ( .A(n14549), .B(n14548), .ZN(n16223) );
  OAI22_X1 U17883 ( .A1(n16209), .A2(n14550), .B1(n14779), .B2(n20806), .ZN(
        n14554) );
  NOR2_X1 U17884 ( .A1(n14552), .A2(n14551), .ZN(n14553) );
  OAI21_X1 U17885 ( .B1(n16223), .B2(n20135), .A(n14556), .ZN(P1_U2976) );
  NAND2_X1 U17886 ( .A1(n14558), .A2(n14557), .ZN(n14559) );
  XNOR2_X1 U17887 ( .A(n14559), .B(n14729), .ZN(n14734) );
  NAND2_X1 U17888 ( .A1(n14560), .A2(n16205), .ZN(n14565) );
  OR2_X1 U17889 ( .A1(n14779), .A2(n20859), .ZN(n14727) );
  OAI21_X1 U17890 ( .B1(n16209), .B2(n14561), .A(n14727), .ZN(n14562) );
  AOI21_X1 U17891 ( .B1(n16204), .B2(n14563), .A(n14562), .ZN(n14564) );
  OAI211_X1 U17892 ( .C1(n14734), .C2(n20135), .A(n14565), .B(n14564), .ZN(
        P1_U2977) );
  NOR3_X1 U17893 ( .A1(n14593), .A2(n16174), .A3(n14746), .ZN(n14576) );
  NOR3_X1 U17894 ( .A1(n14595), .A2(n16173), .A3(n14566), .ZN(n14575) );
  INV_X1 U17895 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14567) );
  AOI22_X1 U17896 ( .A1(n14576), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n14575), .B2(n14567), .ZN(n14568) );
  XOR2_X1 U17897 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n14568), .Z(
        n14743) );
  NAND2_X1 U17898 ( .A1(n16204), .A2(n14569), .ZN(n14570) );
  NAND2_X1 U17899 ( .A1(n16319), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14737) );
  OAI211_X1 U17900 ( .C1(n16209), .C2(n14571), .A(n14570), .B(n14737), .ZN(
        n14572) );
  AOI21_X1 U17901 ( .B1(n14573), .B2(n16205), .A(n14572), .ZN(n14574) );
  OAI21_X1 U17902 ( .B1(n14743), .B2(n20135), .A(n14574), .ZN(P1_U2978) );
  NOR2_X1 U17903 ( .A1(n14576), .A2(n14575), .ZN(n14577) );
  XOR2_X1 U17904 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n14577), .Z(
        n14754) );
  NAND2_X1 U17905 ( .A1(n14578), .A2(n16205), .ZN(n14583) );
  INV_X1 U17906 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20877) );
  OR2_X1 U17907 ( .A1(n14779), .A2(n20877), .ZN(n14745) );
  OAI21_X1 U17908 ( .B1(n16209), .B2(n14579), .A(n14745), .ZN(n14580) );
  AOI21_X1 U17909 ( .B1(n16204), .B2(n14581), .A(n14580), .ZN(n14582) );
  OAI211_X1 U17910 ( .C1(n14754), .C2(n20135), .A(n14583), .B(n14582), .ZN(
        P1_U2979) );
  OAI21_X1 U17911 ( .B1(n16173), .B2(n16248), .A(n14593), .ZN(n14585) );
  XNOR2_X1 U17912 ( .A(n16174), .B(n14746), .ZN(n14584) );
  XNOR2_X1 U17913 ( .A(n14585), .B(n14584), .ZN(n16231) );
  INV_X1 U17914 ( .A(n14586), .ZN(n14591) );
  INV_X1 U17915 ( .A(n14587), .ZN(n14589) );
  AOI22_X1 U17916 ( .A1(n16194), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n16319), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n14588) );
  OAI21_X1 U17917 ( .B1(n14589), .B2(n16202), .A(n14588), .ZN(n14590) );
  AOI21_X1 U17918 ( .B1(n14591), .B2(n16205), .A(n14590), .ZN(n14592) );
  OAI21_X1 U17919 ( .B1(n16231), .B2(n20135), .A(n14592), .ZN(P1_U2980) );
  OAI21_X1 U17920 ( .B1(n14595), .B2(n14594), .A(n14593), .ZN(n16243) );
  NOR2_X1 U17921 ( .A1(n16202), .A2(n14596), .ZN(n14600) );
  INV_X1 U17922 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14598) );
  NOR2_X1 U17923 ( .A1(n14779), .A2(n20798), .ZN(n16246) );
  INV_X1 U17924 ( .A(n16246), .ZN(n14597) );
  OAI21_X1 U17925 ( .B1(n16209), .B2(n14598), .A(n14597), .ZN(n14599) );
  AOI211_X1 U17926 ( .C1(n14601), .C2(n16205), .A(n14600), .B(n14599), .ZN(
        n14602) );
  OAI21_X1 U17927 ( .B1(n20135), .B2(n16243), .A(n14602), .ZN(P1_U2981) );
  INV_X1 U17928 ( .A(n16186), .ZN(n14758) );
  INV_X1 U17929 ( .A(n14603), .ZN(n14755) );
  NOR2_X1 U17930 ( .A1(n14758), .A2(n14755), .ZN(n16172) );
  AOI21_X1 U17931 ( .B1(n16172), .B2(n14605), .A(n14604), .ZN(n14608) );
  NOR2_X1 U17932 ( .A1(n16173), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14607) );
  NAND2_X1 U17933 ( .A1(n14608), .A2(n16174), .ZN(n14606) );
  OAI21_X1 U17934 ( .B1(n14608), .B2(n14607), .A(n14606), .ZN(n14609) );
  XNOR2_X1 U17935 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B(n14609), .ZN(
        n16252) );
  INV_X1 U17936 ( .A(n16252), .ZN(n14615) );
  AOI22_X1 U17937 ( .A1(n16194), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n16319), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n14610) );
  OAI21_X1 U17938 ( .B1(n14611), .B2(n16202), .A(n14610), .ZN(n14612) );
  AOI21_X1 U17939 ( .B1(n14613), .B2(n16205), .A(n14612), .ZN(n14614) );
  OAI21_X1 U17940 ( .B1(n14615), .B2(n20135), .A(n14614), .ZN(P1_U2982) );
  NOR3_X1 U17941 ( .A1(n16172), .A2(n14617), .A3(n14616), .ZN(n14618) );
  XOR2_X1 U17942 ( .A(n14619), .B(n14618), .Z(n16268) );
  NOR2_X1 U17943 ( .A1(n16202), .A2(n14620), .ZN(n14623) );
  OAI22_X1 U17944 ( .A1(n16209), .A2(n14621), .B1(n14779), .B2(n20789), .ZN(
        n14622) );
  AOI211_X1 U17945 ( .C1(n14624), .C2(n16205), .A(n14623), .B(n14622), .ZN(
        n14625) );
  OAI21_X1 U17946 ( .B1(n16268), .B2(n20135), .A(n14625), .ZN(P1_U2986) );
  NAND2_X1 U17947 ( .A1(n14626), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14630) );
  XNOR2_X1 U17948 ( .A(n16186), .B(n14627), .ZN(n14629) );
  MUX2_X1 U17949 ( .A(n14630), .B(n14629), .S(n14628), .Z(n14632) );
  NOR3_X1 U17950 ( .A1(n14626), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n16173), .ZN(n16187) );
  INV_X1 U17951 ( .A(n16187), .ZN(n14631) );
  NAND2_X1 U17952 ( .A1(n14632), .A2(n14631), .ZN(n16289) );
  INV_X1 U17953 ( .A(n16289), .ZN(n14638) );
  AOI22_X1 U17954 ( .A1(n16194), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n16319), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14633) );
  OAI21_X1 U17955 ( .B1(n14634), .B2(n16202), .A(n14633), .ZN(n14635) );
  AOI21_X1 U17956 ( .B1(n14636), .B2(n16205), .A(n14635), .ZN(n14637) );
  OAI21_X1 U17957 ( .B1(n14638), .B2(n20135), .A(n14637), .ZN(P1_U2989) );
  NOR2_X1 U17958 ( .A1(n14740), .A2(n14729), .ZN(n14725) );
  INV_X1 U17959 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16273) );
  NAND4_X1 U17960 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16240) );
  NOR3_X1 U17961 ( .A1(n16248), .A2(n16273), .A3(n16240), .ZN(n14651) );
  NOR2_X1 U17962 ( .A1(n14640), .A2(n14639), .ZN(n14763) );
  NAND2_X1 U17963 ( .A1(n14763), .A2(n16283), .ZN(n14650) );
  INV_X1 U17964 ( .A(n14763), .ZN(n14641) );
  NOR2_X1 U17965 ( .A1(n14642), .A2(n14641), .ZN(n14649) );
  INV_X1 U17966 ( .A(n14643), .ZN(n14645) );
  NOR2_X1 U17967 ( .A1(n10128), .A2(n14650), .ZN(n14644) );
  AOI22_X1 U17968 ( .A1(n14765), .A2(n14649), .B1(n14645), .B2(n14644), .ZN(
        n14750) );
  OAI21_X1 U17969 ( .B1(n20287), .B2(n14650), .A(n14750), .ZN(n16267) );
  NAND2_X1 U17970 ( .A1(n14651), .A2(n16267), .ZN(n16237) );
  NOR2_X1 U17971 ( .A1(n14646), .A2(n16237), .ZN(n14741) );
  NAND2_X1 U17972 ( .A1(n14725), .A2(n14741), .ZN(n14714) );
  NOR2_X1 U17973 ( .A1(n14647), .A2(n14714), .ZN(n16212) );
  NAND2_X1 U17974 ( .A1(n16212), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14700) );
  INV_X1 U17975 ( .A(n14689), .ZN(n14660) );
  OR3_X1 U17976 ( .A1(n14700), .A2(n14660), .A3(n14682), .ZN(n14672) );
  NAND2_X1 U17977 ( .A1(n11923), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14664) );
  INV_X1 U17978 ( .A(n14725), .ZN(n14658) );
  NAND2_X1 U17979 ( .A1(n16312), .A2(n14648), .ZN(n14661) );
  AOI21_X1 U17980 ( .B1(n14649), .B2(n14651), .A(n14715), .ZN(n14654) );
  INV_X1 U17981 ( .A(n14650), .ZN(n14767) );
  AOI21_X1 U17982 ( .B1(n14651), .B2(n14767), .A(n16284), .ZN(n14653) );
  INV_X1 U17983 ( .A(n16230), .ZN(n14655) );
  NAND2_X1 U17984 ( .A1(n14656), .A2(n14655), .ZN(n14657) );
  AOI21_X1 U17985 ( .B1(n16287), .B2(n14658), .A(n14735), .ZN(n16229) );
  NAND2_X1 U17986 ( .A1(n16229), .A2(n14705), .ZN(n14717) );
  NAND2_X1 U17987 ( .A1(n14717), .A2(n14661), .ZN(n16216) );
  INV_X1 U17988 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16211) );
  OAI21_X1 U17989 ( .B1(n16211), .B2(n14709), .A(n16287), .ZN(n14659) );
  NAND2_X1 U17990 ( .A1(n16216), .A2(n14659), .ZN(n14697) );
  AOI21_X1 U17991 ( .B1(n14660), .B2(n16287), .A(n14697), .ZN(n14683) );
  OAI211_X1 U17992 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16312), .A(
        n14683), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14670) );
  NAND3_X1 U17993 ( .A1(n14670), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14661), .ZN(n14663) );
  OAI211_X1 U17994 ( .C1(n14672), .C2(n14664), .A(n14663), .B(n14662), .ZN(
        n14665) );
  AOI21_X1 U17995 ( .B1(n14666), .B2(n20282), .A(n14665), .ZN(n14667) );
  OAI21_X1 U17996 ( .B1(n14668), .B2(n16260), .A(n14667), .ZN(P1_U3000) );
  INV_X1 U17997 ( .A(n14669), .ZN(n14674) );
  INV_X1 U17998 ( .A(n14670), .ZN(n14671) );
  AOI21_X1 U17999 ( .B1(n11919), .B2(n14672), .A(n14671), .ZN(n14673) );
  AOI211_X1 U18000 ( .C1(n14675), .C2(n20282), .A(n14674), .B(n14673), .ZN(
        n14676) );
  OAI21_X1 U18001 ( .B1(n14677), .B2(n16260), .A(n14676), .ZN(P1_U3001) );
  INV_X1 U18002 ( .A(n14678), .ZN(n14685) );
  INV_X1 U18003 ( .A(n14700), .ZN(n14679) );
  NAND3_X1 U18004 ( .A1(n14679), .A2(n14689), .A3(n14682), .ZN(n14680) );
  OAI211_X1 U18005 ( .C1(n14683), .C2(n14682), .A(n14681), .B(n14680), .ZN(
        n14684) );
  AOI21_X1 U18006 ( .B1(n14685), .B2(n20282), .A(n14684), .ZN(n14686) );
  OAI21_X1 U18007 ( .B1(n14687), .B2(n16260), .A(n14686), .ZN(P1_U3002) );
  INV_X1 U18008 ( .A(n14688), .ZN(n14692) );
  NOR3_X1 U18009 ( .A1(n14700), .A2(n14690), .A3(n14689), .ZN(n14691) );
  AOI211_X1 U18010 ( .C1(n14697), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14692), .B(n14691), .ZN(n14695) );
  NAND2_X1 U18011 ( .A1(n14693), .A2(n20282), .ZN(n14694) );
  OAI211_X1 U18012 ( .C1(n14696), .C2(n16260), .A(n14695), .B(n14694), .ZN(
        P1_U3003) );
  NAND2_X1 U18013 ( .A1(n14697), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14699) );
  OAI211_X1 U18014 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n14700), .A(
        n14699), .B(n14698), .ZN(n14701) );
  AOI21_X1 U18015 ( .B1(n14702), .B2(n20282), .A(n14701), .ZN(n14703) );
  OAI21_X1 U18016 ( .B1(n14704), .B2(n16260), .A(n14703), .ZN(P1_U3004) );
  INV_X1 U18017 ( .A(n14714), .ZN(n16222) );
  NAND2_X1 U18018 ( .A1(n16222), .A2(n14705), .ZN(n14706) );
  NOR2_X1 U18019 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n14706), .ZN(
        n16217) );
  INV_X1 U18020 ( .A(n16217), .ZN(n14707) );
  OAI211_X1 U18021 ( .C1(n16216), .C2(n14709), .A(n14708), .B(n14707), .ZN(
        n14710) );
  AOI21_X1 U18022 ( .B1(n14711), .B2(n20282), .A(n14710), .ZN(n14712) );
  OAI21_X1 U18023 ( .B1(n14713), .B2(n16260), .A(n14712), .ZN(P1_U3006) );
  NOR2_X1 U18024 ( .A1(n11915), .A2(n14714), .ZN(n14718) );
  NAND3_X1 U18025 ( .A1(n16229), .A2(n14715), .A3(n16308), .ZN(n14716) );
  OAI211_X1 U18026 ( .C1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n14718), .A(
        n14717), .B(n14716), .ZN(n14720) );
  NAND2_X1 U18027 ( .A1(n14720), .A2(n14719), .ZN(n14721) );
  AOI21_X1 U18028 ( .B1(n14722), .B2(n20282), .A(n14721), .ZN(n14723) );
  OAI21_X1 U18029 ( .B1(n14724), .B2(n16260), .A(n14723), .ZN(P1_U3007) );
  AOI21_X1 U18030 ( .B1(n14740), .B2(n14729), .A(n14725), .ZN(n14732) );
  INV_X1 U18031 ( .A(n14735), .ZN(n14730) );
  NAND2_X1 U18032 ( .A1(n14726), .A2(n20282), .ZN(n14728) );
  OAI211_X1 U18033 ( .C1(n14730), .C2(n14729), .A(n14728), .B(n14727), .ZN(
        n14731) );
  AOI21_X1 U18034 ( .B1(n14741), .B2(n14732), .A(n14731), .ZN(n14733) );
  OAI21_X1 U18035 ( .B1(n14734), .B2(n16260), .A(n14733), .ZN(P1_U3009) );
  NAND2_X1 U18036 ( .A1(n14735), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14736) );
  OAI211_X1 U18037 ( .C1(n14738), .C2(n16259), .A(n14737), .B(n14736), .ZN(
        n14739) );
  AOI21_X1 U18038 ( .B1(n14741), .B2(n14740), .A(n14739), .ZN(n14742) );
  OAI21_X1 U18039 ( .B1(n14743), .B2(n16260), .A(n14742), .ZN(P1_U3010) );
  INV_X1 U18040 ( .A(n14744), .ZN(n14749) );
  INV_X1 U18041 ( .A(n14745), .ZN(n14748) );
  NOR3_X1 U18042 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n14746), .A3(
        n16237), .ZN(n14747) );
  AOI211_X1 U18043 ( .C1(n20282), .C2(n14749), .A(n14748), .B(n14747), .ZN(
        n14753) );
  AOI21_X1 U18044 ( .B1(n14750), .B2(n20287), .A(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14751) );
  OAI21_X1 U18045 ( .B1(n16230), .B2(n14751), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14752) );
  OAI211_X1 U18046 ( .C1(n14754), .C2(n16260), .A(n14753), .B(n14752), .ZN(
        P1_U3011) );
  AOI211_X1 U18047 ( .C1(n14758), .C2(n14757), .A(n14756), .B(n14755), .ZN(
        n14775) );
  NOR2_X1 U18048 ( .A1(n14760), .A2(n14759), .ZN(n14774) );
  AND2_X1 U18049 ( .A1(n14775), .A2(n14774), .ZN(n14776) );
  NOR2_X1 U18050 ( .A1(n14760), .A2(n14776), .ZN(n14762) );
  XOR2_X1 U18051 ( .A(n14762), .B(n14761), .Z(n16160) );
  NAND2_X1 U18052 ( .A1(n16160), .A2(n20285), .ZN(n14773) );
  AOI22_X1 U18053 ( .A1(n16133), .A2(n20282), .B1(n16319), .B2(
        P1_REIP_REG_16__SCAN_IN), .ZN(n14772) );
  NAND2_X1 U18054 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14763), .ZN(
        n16257) );
  AOI21_X1 U18055 ( .B1(n14765), .B2(n16257), .A(n14764), .ZN(n14768) );
  OAI221_X1 U18056 ( .B1(n14768), .B2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), 
        .C1(n14768), .C2(n14767), .A(n14766), .ZN(n16238) );
  INV_X1 U18057 ( .A(n16238), .ZN(n16274) );
  OAI21_X1 U18058 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16312), .A(
        n16274), .ZN(n14782) );
  NAND2_X1 U18059 ( .A1(n14782), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14771) );
  NAND2_X1 U18060 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n16267), .ZN(
        n16239) );
  NOR2_X1 U18061 ( .A1(n16266), .A2(n16239), .ZN(n16249) );
  NOR2_X1 U18062 ( .A1(n14781), .A2(n14124), .ZN(n16250) );
  AOI21_X1 U18063 ( .B1(n14781), .B2(n14124), .A(n16250), .ZN(n14769) );
  NAND2_X1 U18064 ( .A1(n16249), .A2(n14769), .ZN(n14770) );
  NAND4_X1 U18065 ( .A1(n14773), .A2(n14772), .A3(n14771), .A4(n14770), .ZN(
        P1_U3015) );
  NOR2_X1 U18066 ( .A1(n14775), .A2(n14774), .ZN(n14777) );
  NOR2_X1 U18067 ( .A1(n14777), .A2(n14776), .ZN(n16169) );
  INV_X1 U18068 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n14778) );
  OAI22_X1 U18069 ( .A1(n16138), .A2(n16259), .B1(n14779), .B2(n14778), .ZN(
        n14780) );
  AOI21_X1 U18070 ( .B1(n16249), .B2(n14781), .A(n14780), .ZN(n14784) );
  NAND2_X1 U18071 ( .A1(n14782), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14783) );
  OAI211_X1 U18072 ( .C1(n16169), .C2(n16260), .A(n14784), .B(n14783), .ZN(
        P1_U3016) );
  OAI21_X1 U18073 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n9673), .A(n20568), 
        .ZN(n14785) );
  OAI21_X1 U18074 ( .B1(n14786), .B2(n13652), .A(n14785), .ZN(n14787) );
  MUX2_X1 U18075 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n14787), .S(
        n20293), .Z(P1_U3477) );
  NOR3_X1 U18076 ( .A1(n14788), .A2(n13346), .A3(n14795), .ZN(n14791) );
  NOR2_X1 U18077 ( .A1(n13652), .A2(n14789), .ZN(n14790) );
  AOI211_X1 U18078 ( .C1(n14793), .C2(n14792), .A(n14791), .B(n14790), .ZN(
        n16068) );
  INV_X1 U18079 ( .A(n14794), .ZN(n14798) );
  NOR3_X1 U18080 ( .A1(n13346), .A2(n14795), .A3(n14802), .ZN(n14796) );
  AOI21_X1 U18081 ( .B1(n14798), .B2(n14797), .A(n14796), .ZN(n14799) );
  OAI21_X1 U18082 ( .B1(n16068), .B2(n14804), .A(n14799), .ZN(n14800) );
  MUX2_X1 U18083 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14800), .S(
        n16340), .Z(P1_U3473) );
  INV_X1 U18084 ( .A(n16061), .ZN(n14805) );
  INV_X1 U18085 ( .A(n14801), .ZN(n14803) );
  OAI22_X1 U18086 ( .A1(n14805), .A2(n14804), .B1(n14803), .B2(n14802), .ZN(
        n14806) );
  MUX2_X1 U18087 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14806), .S(
        n16340), .Z(P1_U3469) );
  INV_X1 U18088 ( .A(n14807), .ZN(n14821) );
  OAI22_X1 U18089 ( .A1(n10158), .A2(n19334), .B1(n20040), .B2(n19301), .ZN(
        n14817) );
  INV_X1 U18090 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n14814) );
  NOR2_X1 U18091 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n14810), .ZN(n14811) );
  NAND2_X1 U18092 ( .A1(n19153), .A2(n14811), .ZN(n14812) );
  OAI22_X1 U18093 ( .A1(n14815), .A2(n19320), .B1(n14814), .B2(n19303), .ZN(
        n14816) );
  AOI211_X1 U18094 ( .C1(n14818), .C2(n19324), .A(n14817), .B(n14816), .ZN(
        n14819) );
  OAI211_X1 U18095 ( .C1(n14821), .C2(n19321), .A(n14820), .B(n14819), .ZN(
        P2_U2825) );
  OAI211_X1 U18096 ( .C1(n14823), .C2(n15313), .A(n19315), .B(n14822), .ZN(
        n14836) );
  NOR2_X1 U18097 ( .A1(n15025), .A2(n14824), .ZN(n14825) );
  OR2_X1 U18098 ( .A1(n15009), .A2(n14825), .ZN(n15498) );
  NOR2_X1 U18099 ( .A1(n9727), .A2(n14827), .ZN(n14828) );
  OR2_X1 U18100 ( .A1(n14826), .A2(n14828), .ZN(n15503) );
  INV_X1 U18101 ( .A(n15503), .ZN(n16420) );
  OAI22_X1 U18102 ( .A1(n14829), .A2(n19334), .B1(n20026), .B2(n19301), .ZN(
        n14830) );
  AOI21_X1 U18103 ( .B1(n19327), .B2(n16420), .A(n14830), .ZN(n14832) );
  NAND2_X1 U18104 ( .A1(n19326), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n14831) );
  OAI211_X1 U18105 ( .C1(n15498), .C2(n19321), .A(n14832), .B(n14831), .ZN(
        n14833) );
  AOI21_X1 U18106 ( .B1(n14834), .B2(n19324), .A(n14833), .ZN(n14835) );
  NAND2_X1 U18107 ( .A1(n14836), .A2(n14835), .ZN(P2_U2832) );
  XOR2_X1 U18108 ( .A(n14837), .B(n15038), .Z(n15533) );
  NAND2_X1 U18109 ( .A1(n15533), .A2(n19314), .ZN(n14843) );
  NAND2_X1 U18110 ( .A1(n15192), .A2(n14838), .ZN(n14839) );
  AND2_X1 U18111 ( .A1(n15173), .A2(n14839), .ZN(n15526) );
  OAI22_X1 U18112 ( .A1(n14840), .A2(n19334), .B1(n20022), .B2(n19301), .ZN(
        n14841) );
  AOI21_X1 U18113 ( .B1(n19327), .B2(n15526), .A(n14841), .ZN(n14842) );
  OAI211_X1 U18114 ( .C1(n19303), .C2(n14844), .A(n14843), .B(n14842), .ZN(
        n14848) );
  INV_X1 U18115 ( .A(n19179), .ZN(n14845) );
  AOI221_X1 U18116 ( .B1(n14846), .B2(n14845), .C1(n15336), .C2(n19179), .A(
        n19977), .ZN(n14847) );
  AOI211_X1 U18117 ( .C1(n19324), .C2(n14849), .A(n14848), .B(n14847), .ZN(
        n14850) );
  INV_X1 U18118 ( .A(n14850), .ZN(P2_U2834) );
  NOR2_X1 U18119 ( .A1(n19244), .A2(n14851), .ZN(n14853) );
  XNOR2_X1 U18120 ( .A(n14853), .B(n14852), .ZN(n14854) );
  NAND2_X1 U18121 ( .A1(n14854), .A2(n19315), .ZN(n14865) );
  INV_X1 U18122 ( .A(n14855), .ZN(n15098) );
  NAND2_X1 U18123 ( .A1(n15098), .A2(n14856), .ZN(n14857) );
  AND2_X1 U18124 ( .A1(n15081), .A2(n14857), .ZN(n16455) );
  INV_X1 U18125 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n20011) );
  OAI21_X1 U18126 ( .B1(n20011), .B2(n19301), .A(n19300), .ZN(n14863) );
  AOI21_X1 U18127 ( .B1(n14860), .B2(n14859), .A(n14858), .ZN(n19344) );
  AOI22_X1 U18128 ( .A1(n19327), .A2(n19344), .B1(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n19308), .ZN(n14861) );
  OAI21_X1 U18129 ( .B1(n19303), .B2(n10725), .A(n14861), .ZN(n14862) );
  AOI211_X1 U18130 ( .C1(n16455), .C2(n19314), .A(n14863), .B(n14862), .ZN(
        n14864) );
  OAI211_X1 U18131 ( .C1(n19304), .C2(n14866), .A(n14865), .B(n14864), .ZN(
        P2_U2842) );
  NAND2_X1 U18132 ( .A1(n19310), .A2(n14867), .ZN(n14868) );
  XNOR2_X1 U18133 ( .A(n14869), .B(n14868), .ZN(n14881) );
  AND2_X1 U18134 ( .A1(n14871), .A2(n14870), .ZN(n14872) );
  OR2_X1 U18135 ( .A1(n14872), .A2(n15103), .ZN(n16547) );
  INV_X1 U18136 ( .A(n16547), .ZN(n16487) );
  NAND2_X1 U18137 ( .A1(n16487), .A2(n19314), .ZN(n14879) );
  OAI22_X1 U18138 ( .A1(n14874), .A2(n19304), .B1(n14873), .B2(n19334), .ZN(
        n14875) );
  INV_X1 U18139 ( .A(n14875), .ZN(n14876) );
  OAI21_X1 U18140 ( .B1(n19303), .B2(n15115), .A(n14876), .ZN(n14877) );
  AOI211_X1 U18141 ( .C1(n19325), .C2(P2_REIP_REG_10__SCAN_IN), .A(n19427), 
        .B(n14877), .ZN(n14878) );
  OAI211_X1 U18142 ( .C1(n16548), .C2(n19320), .A(n14879), .B(n14878), .ZN(
        n14880) );
  AOI21_X1 U18143 ( .B1(n14881), .B2(n19315), .A(n14880), .ZN(n14882) );
  INV_X1 U18144 ( .A(n14882), .ZN(P2_U2845) );
  INV_X1 U18145 ( .A(n14883), .ZN(n14894) );
  NOR2_X1 U18146 ( .A1(n19244), .A2(n14884), .ZN(n14886) );
  XNOR2_X1 U18147 ( .A(n14886), .B(n14885), .ZN(n14887) );
  NAND2_X1 U18148 ( .A1(n14887), .A2(n19315), .ZN(n14893) );
  OAI21_X1 U18149 ( .B1(n16500), .B2(n19334), .A(n19300), .ZN(n14889) );
  NOR2_X1 U18150 ( .A1(n19320), .A2(n15627), .ZN(n14888) );
  AOI211_X1 U18151 ( .C1(n19325), .C2(P2_REIP_REG_9__SCAN_IN), .A(n14889), .B(
        n14888), .ZN(n14890) );
  OAI21_X1 U18152 ( .B1(n15626), .B2(n19321), .A(n14890), .ZN(n14891) );
  AOI21_X1 U18153 ( .B1(P2_EBX_REG_9__SCAN_IN), .B2(n19326), .A(n14891), .ZN(
        n14892) );
  OAI211_X1 U18154 ( .C1(n19304), .C2(n14894), .A(n14893), .B(n14892), .ZN(
        P2_U2846) );
  NOR2_X1 U18155 ( .A1(n19244), .A2(n14895), .ZN(n14896) );
  XNOR2_X1 U18156 ( .A(n14896), .B(n15401), .ZN(n14897) );
  NAND2_X1 U18157 ( .A1(n14897), .A2(n19315), .ZN(n14905) );
  AOI22_X1 U18158 ( .A1(n14898), .A2(n19324), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n19326), .ZN(n14899) );
  OAI21_X1 U18159 ( .B1(n10706), .B2(n19334), .A(n14899), .ZN(n14902) );
  AOI21_X1 U18160 ( .B1(n19325), .B2(P2_REIP_REG_7__SCAN_IN), .A(n19427), .ZN(
        n14900) );
  OAI21_X1 U18161 ( .B1(n15640), .B2(n19321), .A(n14900), .ZN(n14901) );
  AOI211_X1 U18162 ( .C1(n14903), .C2(n19327), .A(n14902), .B(n14901), .ZN(
        n14904) );
  NAND2_X1 U18163 ( .A1(n14905), .A2(n14904), .ZN(P2_U2848) );
  NOR2_X1 U18164 ( .A1(n19244), .A2(n14906), .ZN(n14907) );
  XNOR2_X1 U18165 ( .A(n14907), .B(n15424), .ZN(n14908) );
  NAND2_X1 U18166 ( .A1(n14908), .A2(n19315), .ZN(n14915) );
  NOR2_X1 U18167 ( .A1(n14909), .A2(n19304), .ZN(n14913) );
  NAND2_X1 U18168 ( .A1(n15425), .A2(n19314), .ZN(n14911) );
  AOI21_X1 U18169 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n19308), .A(
        n19427), .ZN(n14910) );
  OAI211_X1 U18170 ( .C1(n19301), .C2(n15426), .A(n14911), .B(n14910), .ZN(
        n14912) );
  AOI211_X1 U18171 ( .C1(P2_EBX_REG_5__SCAN_IN), .C2(n19326), .A(n14913), .B(
        n14912), .ZN(n14914) );
  OAI211_X1 U18172 ( .C1(n15662), .C2(n19320), .A(n14915), .B(n14914), .ZN(
        P2_U2850) );
  NAND2_X1 U18173 ( .A1(n14917), .A2(n14916), .ZN(n19154) );
  AND2_X1 U18174 ( .A1(n19310), .A2(n14918), .ZN(n14920) );
  AOI21_X1 U18175 ( .B1(n19425), .B2(n14920), .A(n19977), .ZN(n14919) );
  OAI21_X1 U18176 ( .B1(n19425), .B2(n14920), .A(n14919), .ZN(n14928) );
  INV_X1 U18177 ( .A(n19359), .ZN(n14921) );
  AOI22_X1 U18178 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n19326), .B1(n19327), .B2(
        n14921), .ZN(n14922) );
  OAI211_X1 U18179 ( .C1(n19439), .C2(n19334), .A(n19300), .B(n14922), .ZN(
        n14923) );
  AOI21_X1 U18180 ( .B1(n19325), .B2(P2_REIP_REG_4__SCAN_IN), .A(n14923), .ZN(
        n14924) );
  OAI21_X1 U18181 ( .B1(n14925), .B2(n19304), .A(n14924), .ZN(n14926) );
  AOI21_X1 U18182 ( .B1(n19434), .B2(n19314), .A(n14926), .ZN(n14927) );
  OAI211_X1 U18183 ( .C1(n19154), .C2(n19361), .A(n14928), .B(n14927), .ZN(
        P2_U2851) );
  NOR2_X1 U18184 ( .A1(n19244), .A2(n14929), .ZN(n14931) );
  XNOR2_X1 U18185 ( .A(n14931), .B(n14930), .ZN(n14932) );
  NAND2_X1 U18186 ( .A1(n14932), .A2(n19315), .ZN(n14939) );
  AOI22_X1 U18187 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n19308), .B1(
        n19327), .B2(n20069), .ZN(n14933) );
  OAI21_X1 U18188 ( .B1(n19301), .B2(n10684), .A(n14933), .ZN(n14934) );
  AOI21_X1 U18189 ( .B1(n19326), .B2(P2_EBX_REG_3__SCAN_IN), .A(n14934), .ZN(
        n14935) );
  OAI21_X1 U18190 ( .B1(n14936), .B2(n19304), .A(n14935), .ZN(n14937) );
  AOI21_X1 U18191 ( .B1(n13270), .B2(n19314), .A(n14937), .ZN(n14938) );
  OAI211_X1 U18192 ( .C1(n19154), .C2(n19727), .A(n14939), .B(n14938), .ZN(
        P2_U2852) );
  NAND2_X1 U18193 ( .A1(n19310), .A2(n14959), .ZN(n14940) );
  XNOR2_X1 U18194 ( .A(n14941), .B(n14940), .ZN(n14950) );
  OAI22_X1 U18195 ( .A1(n19304), .A2(n14942), .B1(n20000), .B2(n19301), .ZN(
        n14946) );
  OAI22_X1 U18196 ( .A1(n19303), .A2(n14944), .B1(n14943), .B2(n19334), .ZN(
        n14945) );
  AOI211_X1 U18197 ( .C1(n19327), .C2(n20077), .A(n14946), .B(n14945), .ZN(
        n14948) );
  INV_X1 U18198 ( .A(n19154), .ZN(n19337) );
  NAND2_X1 U18199 ( .A1(n19440), .A2(n19337), .ZN(n14947) );
  OAI211_X1 U18200 ( .C1(n19321), .C2(n12429), .A(n14948), .B(n14947), .ZN(
        n14949) );
  AOI21_X1 U18201 ( .B1(n14950), .B2(n19315), .A(n14949), .ZN(n14951) );
  INV_X1 U18202 ( .A(n14951), .ZN(P2_U2853) );
  OAI22_X1 U18203 ( .A1(n19303), .A2(n14953), .B1(n19304), .B2(n14952), .ZN(
        n14956) );
  OAI22_X1 U18204 ( .A1(n14954), .A2(n19334), .B1(n10624), .B2(n19301), .ZN(
        n14955) );
  AOI211_X1 U18205 ( .C1(n19327), .C2(n20086), .A(n14956), .B(n14955), .ZN(
        n14957) );
  OAI21_X1 U18206 ( .B1(n14958), .B2(n19321), .A(n14957), .ZN(n14962) );
  NAND2_X1 U18207 ( .A1(n19244), .A2(n19315), .ZN(n19333) );
  OAI211_X1 U18208 ( .C1(n19340), .C2(n14960), .A(n19310), .B(n14959), .ZN(
        n15691) );
  OAI22_X1 U18209 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19333), .B1(
        n15691), .B2(n19977), .ZN(n14961) );
  AOI211_X1 U18210 ( .C1(n19337), .C2(n20082), .A(n14962), .B(n14961), .ZN(
        n14963) );
  INV_X1 U18211 ( .A(n14963), .ZN(P2_U2854) );
  MUX2_X1 U18212 ( .A(P2_EBX_REG_31__SCAN_IN), .B(n14964), .S(n15116), .Z(
        P2_U2856) );
  OR2_X1 U18213 ( .A1(n14967), .A2(n14966), .ZN(n15120) );
  NAND3_X1 U18214 ( .A1(n15120), .A2(n14968), .A3(n15109), .ZN(n14970) );
  NAND2_X1 U18215 ( .A1(n15089), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14969) );
  OAI211_X1 U18216 ( .C1(n15089), .C2(n16348), .A(n14970), .B(n14969), .ZN(
        P2_U2858) );
  INV_X1 U18217 ( .A(n14971), .ZN(n14972) );
  NAND2_X1 U18218 ( .A1(n14973), .A2(n14972), .ZN(n14975) );
  XNOR2_X1 U18219 ( .A(n14975), .B(n14974), .ZN(n15138) );
  NAND2_X1 U18220 ( .A1(n15089), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n14978) );
  AOI21_X1 U18221 ( .B1(n14976), .B2(n14984), .A(n9685), .ZN(n16363) );
  NAND2_X1 U18222 ( .A1(n16363), .A2(n15116), .ZN(n14977) );
  OAI211_X1 U18223 ( .C1(n15138), .C2(n15106), .A(n14978), .B(n14977), .ZN(
        P2_U2859) );
  OAI21_X1 U18224 ( .B1(n9758), .B2(n14981), .A(n14980), .ZN(n15144) );
  OR2_X1 U18225 ( .A1(n14991), .A2(n14982), .ZN(n14983) );
  NAND2_X1 U18226 ( .A1(n14984), .A2(n14983), .ZN(n16374) );
  NOR2_X1 U18227 ( .A1(n16374), .A2(n15089), .ZN(n14985) );
  AOI21_X1 U18228 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n15089), .A(n14985), .ZN(
        n14986) );
  OAI21_X1 U18229 ( .B1(n15144), .B2(n15106), .A(n14986), .ZN(P2_U2860) );
  OAI21_X1 U18230 ( .B1(n14987), .B2(n14989), .A(n14988), .ZN(n15154) );
  AND2_X1 U18231 ( .A1(n15000), .A2(n14990), .ZN(n14992) );
  OR2_X1 U18232 ( .A1(n14992), .A2(n14991), .ZN(n16384) );
  NOR2_X1 U18233 ( .A1(n16384), .A2(n15089), .ZN(n14993) );
  AOI21_X1 U18234 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n15089), .A(n14993), .ZN(
        n14994) );
  OAI21_X1 U18235 ( .B1(n15154), .B2(n15106), .A(n14994), .ZN(P2_U2861) );
  OAI21_X1 U18236 ( .B1(n14995), .B2(n14997), .A(n14996), .ZN(n15164) );
  NAND2_X1 U18237 ( .A1(n15011), .A2(n14998), .ZN(n14999) );
  NAND2_X1 U18238 ( .A1(n15000), .A2(n14999), .ZN(n16396) );
  NOR2_X1 U18239 ( .A1(n16396), .A2(n15089), .ZN(n15001) );
  AOI21_X1 U18240 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n15089), .A(n15001), .ZN(
        n15002) );
  OAI21_X1 U18241 ( .B1(n15164), .B2(n15106), .A(n15002), .ZN(P2_U2862) );
  AOI21_X1 U18242 ( .B1(n15003), .B2(n15005), .A(n15004), .ZN(n15006) );
  XOR2_X1 U18243 ( .A(n15007), .B(n15006), .Z(n15171) );
  OR2_X1 U18244 ( .A1(n15009), .A2(n15008), .ZN(n15010) );
  NAND2_X1 U18245 ( .A1(n15011), .A2(n15010), .ZN(n16407) );
  NOR2_X1 U18246 ( .A1(n16407), .A2(n15089), .ZN(n15012) );
  AOI21_X1 U18247 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n15089), .A(n15012), .ZN(
        n15013) );
  OAI21_X1 U18248 ( .B1(n15171), .B2(n15106), .A(n15013), .ZN(P2_U2863) );
  AOI21_X1 U18249 ( .B1(n15014), .B2(n15016), .A(n15015), .ZN(n16421) );
  NAND2_X1 U18250 ( .A1(n16421), .A2(n15109), .ZN(n15018) );
  NAND2_X1 U18251 ( .A1(n15089), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n15017) );
  OAI211_X1 U18252 ( .C1(n15498), .C2(n15089), .A(n15018), .B(n15017), .ZN(
        P2_U2864) );
  INV_X1 U18253 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n15028) );
  AOI21_X1 U18254 ( .B1(n15021), .B2(n15020), .A(n12166), .ZN(n15179) );
  NAND2_X1 U18255 ( .A1(n15179), .A2(n15109), .ZN(n15027) );
  AND2_X1 U18256 ( .A1(n15023), .A2(n15022), .ZN(n15024) );
  NOR2_X1 U18257 ( .A1(n15025), .A2(n15024), .ZN(n16048) );
  NAND2_X1 U18258 ( .A1(n16048), .A2(n15116), .ZN(n15026) );
  OAI211_X1 U18259 ( .C1(n15116), .C2(n15028), .A(n15027), .B(n15026), .ZN(
        P2_U2865) );
  OAI21_X1 U18260 ( .B1(n15029), .B2(n15030), .A(n15020), .ZN(n15189) );
  NAND2_X1 U18261 ( .A1(n15089), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n15032) );
  NAND2_X1 U18262 ( .A1(n15533), .A2(n15116), .ZN(n15031) );
  OAI211_X1 U18263 ( .C1(n15189), .C2(n15106), .A(n15032), .B(n15031), .ZN(
        P2_U2866) );
  AOI21_X1 U18264 ( .B1(n15035), .B2(n15034), .A(n15029), .ZN(n15197) );
  NAND2_X1 U18265 ( .A1(n15197), .A2(n15109), .ZN(n15041) );
  OR2_X1 U18266 ( .A1(n15046), .A2(n15036), .ZN(n15037) );
  NAND2_X1 U18267 ( .A1(n15038), .A2(n15037), .ZN(n19189) );
  INV_X1 U18268 ( .A(n19189), .ZN(n15039) );
  NAND2_X1 U18269 ( .A1(n15039), .A2(n15116), .ZN(n15040) );
  OAI211_X1 U18270 ( .C1(n15116), .C2(n19181), .A(n15041), .B(n15040), .ZN(
        P2_U2867) );
  OAI21_X1 U18271 ( .B1(n15042), .B2(n15043), .A(n15034), .ZN(n15212) );
  NOR2_X1 U18272 ( .A1(n15053), .A2(n15044), .ZN(n15045) );
  OR2_X1 U18273 ( .A1(n15046), .A2(n15045), .ZN(n19201) );
  NOR2_X1 U18274 ( .A1(n19201), .A2(n15089), .ZN(n15047) );
  AOI21_X1 U18275 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n15089), .A(n15047), .ZN(
        n15048) );
  OAI21_X1 U18276 ( .B1(n15212), .B2(n15106), .A(n15048), .ZN(P2_U2868) );
  AOI21_X1 U18277 ( .B1(n15050), .B2(n15049), .A(n15042), .ZN(n15219) );
  NAND2_X1 U18278 ( .A1(n15219), .A2(n15109), .ZN(n15055) );
  AND2_X1 U18279 ( .A1(n15061), .A2(n15051), .ZN(n15052) );
  NOR2_X1 U18280 ( .A1(n15053), .A2(n15052), .ZN(n19215) );
  NAND2_X1 U18281 ( .A1(n19215), .A2(n15116), .ZN(n15054) );
  OAI211_X1 U18282 ( .C1(n15116), .C2(n19208), .A(n15055), .B(n15054), .ZN(
        P2_U2869) );
  AND2_X1 U18283 ( .A1(n15056), .A2(n15057), .ZN(n15064) );
  OAI21_X1 U18284 ( .B1(n15064), .B2(n15058), .A(n15049), .ZN(n15231) );
  NAND2_X1 U18285 ( .A1(n15068), .A2(n15059), .ZN(n15060) );
  NAND2_X1 U18286 ( .A1(n15061), .A2(n15060), .ZN(n19227) );
  NOR2_X1 U18287 ( .A1(n19227), .A2(n15089), .ZN(n15062) );
  AOI21_X1 U18288 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n15089), .A(n15062), .ZN(
        n15063) );
  OAI21_X1 U18289 ( .B1(n15231), .B2(n15106), .A(n15063), .ZN(P2_U2870) );
  OR2_X1 U18290 ( .A1(n15083), .A2(n15073), .ZN(n15065) );
  AOI21_X1 U18291 ( .B1(n15066), .B2(n15065), .A(n15064), .ZN(n15238) );
  NAND2_X1 U18292 ( .A1(n15238), .A2(n15109), .ZN(n15071) );
  OR2_X1 U18293 ( .A1(n15076), .A2(n15067), .ZN(n15069) );
  NAND2_X1 U18294 ( .A1(n19238), .A2(n15116), .ZN(n15070) );
  OAI211_X1 U18295 ( .C1(n15116), .C2(n15072), .A(n15071), .B(n15070), .ZN(
        P2_U2871) );
  XNOR2_X1 U18296 ( .A(n15083), .B(n15073), .ZN(n15079) );
  NOR2_X1 U18297 ( .A1(n9766), .A2(n15074), .ZN(n15075) );
  OR2_X1 U18298 ( .A1(n15076), .A2(n15075), .ZN(n16508) );
  INV_X1 U18299 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n15077) );
  MUX2_X1 U18300 ( .A(n16508), .B(n15077), .S(n15089), .Z(n15078) );
  OAI21_X1 U18301 ( .B1(n15079), .B2(n15106), .A(n15078), .ZN(P2_U2872) );
  AND2_X1 U18302 ( .A1(n15081), .A2(n15080), .ZN(n15082) );
  OR2_X1 U18303 ( .A1(n15082), .A2(n9766), .ZN(n15603) );
  AND2_X1 U18304 ( .A1(n9703), .A2(n15088), .ZN(n15085) );
  OAI211_X1 U18305 ( .C1(n15085), .C2(n15084), .A(n15109), .B(n15083), .ZN(
        n15087) );
  NAND2_X1 U18306 ( .A1(n15089), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n15086) );
  OAI211_X1 U18307 ( .C1(n15603), .C2(n15089), .A(n15087), .B(n15086), .ZN(
        P2_U2873) );
  XNOR2_X1 U18308 ( .A(n9703), .B(n15088), .ZN(n15091) );
  INV_X1 U18309 ( .A(n16455), .ZN(n16519) );
  MUX2_X1 U18310 ( .A(n16519), .B(n10725), .S(n15089), .Z(n15090) );
  OAI21_X1 U18311 ( .B1(n15091), .B2(n15106), .A(n15090), .ZN(P2_U2874) );
  AOI21_X1 U18312 ( .B1(n15092), .B2(n15101), .A(n15093), .ZN(n15094) );
  OR3_X1 U18313 ( .A1(n9703), .A2(n15094), .A3(n15106), .ZN(n15100) );
  NAND2_X1 U18314 ( .A1(n15095), .A2(n15096), .ZN(n15097) );
  NAND2_X1 U18315 ( .A1(n19274), .A2(n15116), .ZN(n15099) );
  OAI211_X1 U18316 ( .C1(n15116), .C2(n10722), .A(n15100), .B(n15099), .ZN(
        P2_U2875) );
  XNOR2_X1 U18317 ( .A(n15092), .B(n15101), .ZN(n15107) );
  OAI21_X1 U18318 ( .B1(n15103), .B2(n15102), .A(n15095), .ZN(n19281) );
  MUX2_X1 U18319 ( .A(n15104), .B(n19281), .S(n15116), .Z(n15105) );
  OAI21_X1 U18320 ( .B1(n15107), .B2(n15106), .A(n15105), .ZN(P2_U2876) );
  INV_X1 U18321 ( .A(n15108), .ZN(n15112) );
  INV_X1 U18322 ( .A(n15092), .ZN(n15110) );
  OAI211_X1 U18323 ( .C1(n15112), .C2(n15111), .A(n15110), .B(n15109), .ZN(
        n15114) );
  NAND2_X1 U18324 ( .A1(n16487), .A2(n15116), .ZN(n15113) );
  OAI211_X1 U18325 ( .C1(n15116), .C2(n15115), .A(n15114), .B(n15113), .ZN(
        P2_U2877) );
  INV_X1 U18326 ( .A(n16419), .ZN(n15206) );
  AOI22_X1 U18327 ( .A1(n15117), .A2(n19383), .B1(P2_EAX_REG_31__SCAN_IN), 
        .B2(n19382), .ZN(n15119) );
  NAND2_X1 U18328 ( .A1(n16418), .A2(BUF2_REG_31__SCAN_IN), .ZN(n15118) );
  OAI211_X1 U18329 ( .C1(n15206), .C2(n19484), .A(n15119), .B(n15118), .ZN(
        P2_U2888) );
  NAND3_X1 U18330 ( .A1(n15120), .A2(n14968), .A3(n19385), .ZN(n15127) );
  INV_X1 U18331 ( .A(n15121), .ZN(n15122) );
  AOI21_X1 U18332 ( .B1(n15123), .B2(n15131), .A(n15122), .ZN(n16349) );
  AOI22_X1 U18333 ( .A1(n16349), .A2(n19383), .B1(P2_EAX_REG_29__SCAN_IN), 
        .B2(n19382), .ZN(n15126) );
  AOI22_X1 U18334 ( .A1(n16418), .A2(BUF2_REG_29__SCAN_IN), .B1(n16419), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n15125) );
  NAND2_X1 U18335 ( .A1(n16417), .A2(n19345), .ZN(n15124) );
  NAND4_X1 U18336 ( .A1(n15127), .A2(n15126), .A3(n15125), .A4(n15124), .ZN(
        P2_U2890) );
  OR2_X1 U18337 ( .A1(n15128), .A2(n15129), .ZN(n15130) );
  NAND2_X1 U18338 ( .A1(n15131), .A2(n15130), .ZN(n16369) );
  INV_X1 U18339 ( .A(n16369), .ZN(n15440) );
  OAI22_X1 U18340 ( .A1(n15134), .A2(n15133), .B1(n19357), .B2(n15132), .ZN(
        n15135) );
  AOI21_X1 U18341 ( .B1(n19383), .B2(n15440), .A(n15135), .ZN(n15137) );
  AOI22_X1 U18342 ( .A1(n16418), .A2(BUF2_REG_28__SCAN_IN), .B1(n16419), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n15136) );
  OAI211_X1 U18343 ( .C1(n15138), .C2(n15230), .A(n15137), .B(n15136), .ZN(
        P2_U2891) );
  NOR2_X1 U18344 ( .A1(n15147), .A2(n15139), .ZN(n15140) );
  OR2_X1 U18345 ( .A1(n15128), .A2(n15140), .ZN(n16373) );
  OAI22_X1 U18346 ( .A1(n19358), .A2(n16373), .B1(n19357), .B2(n13018), .ZN(
        n15141) );
  AOI21_X1 U18347 ( .B1(n16417), .B2(n19348), .A(n15141), .ZN(n15143) );
  AOI22_X1 U18348 ( .A1(n16418), .A2(BUF2_REG_27__SCAN_IN), .B1(n16419), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n15142) );
  OAI211_X1 U18349 ( .C1(n15144), .C2(n15230), .A(n15143), .B(n15142), .ZN(
        P2_U2892) );
  AND2_X1 U18350 ( .A1(n15158), .A2(n15145), .ZN(n15146) );
  NOR2_X1 U18351 ( .A1(n15147), .A2(n15146), .ZN(n16385) );
  INV_X1 U18352 ( .A(n16385), .ZN(n15149) );
  OAI22_X1 U18353 ( .A1(n19358), .A2(n15149), .B1(n19357), .B2(n15148), .ZN(
        n15150) );
  AOI21_X1 U18354 ( .B1(n16417), .B2(n15151), .A(n15150), .ZN(n15153) );
  AOI22_X1 U18355 ( .A1(n16418), .A2(BUF2_REG_26__SCAN_IN), .B1(n16419), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n15152) );
  OAI211_X1 U18356 ( .C1(n15154), .C2(n15230), .A(n15153), .B(n15152), .ZN(
        P2_U2893) );
  NAND2_X1 U18357 ( .A1(n15156), .A2(n15155), .ZN(n15157) );
  AND2_X1 U18358 ( .A1(n15158), .A2(n15157), .ZN(n15478) );
  INV_X1 U18359 ( .A(n15478), .ZN(n16395) );
  OAI22_X1 U18360 ( .A1(n19358), .A2(n16395), .B1(n19357), .B2(n15159), .ZN(
        n15160) );
  AOI21_X1 U18361 ( .B1(n16417), .B2(n15161), .A(n15160), .ZN(n15163) );
  AOI22_X1 U18362 ( .A1(n16418), .A2(BUF2_REG_25__SCAN_IN), .B1(n16419), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n15162) );
  OAI211_X1 U18363 ( .C1(n15164), .C2(n15230), .A(n15163), .B(n15162), .ZN(
        P2_U2894) );
  INV_X1 U18364 ( .A(n15165), .ZN(n15166) );
  XNOR2_X1 U18365 ( .A(n14826), .B(n15166), .ZN(n15490) );
  INV_X1 U18366 ( .A(n15490), .ZN(n16406) );
  OAI22_X1 U18367 ( .A1(n19358), .A2(n16406), .B1(n19357), .B2(n15167), .ZN(
        n15168) );
  AOI21_X1 U18368 ( .B1(n16417), .B2(n19351), .A(n15168), .ZN(n15170) );
  AOI22_X1 U18369 ( .A1(n16418), .A2(BUF2_REG_24__SCAN_IN), .B1(n16419), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n15169) );
  OAI211_X1 U18370 ( .C1(n15171), .C2(n15230), .A(n15170), .B(n15169), .ZN(
        P2_U2895) );
  AND2_X1 U18371 ( .A1(n15173), .A2(n15172), .ZN(n15174) );
  OR2_X1 U18372 ( .A1(n15174), .A2(n9727), .ZN(n16060) );
  AOI22_X1 U18373 ( .A1(n16418), .A2(BUF2_REG_22__SCAN_IN), .B1(n16419), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n15177) );
  AOI22_X1 U18374 ( .A1(n16417), .A2(n15175), .B1(n19382), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n15176) );
  OAI211_X1 U18375 ( .C1(n19358), .C2(n16060), .A(n15177), .B(n15176), .ZN(
        n15178) );
  AOI21_X1 U18376 ( .B1(n15179), .B2(n19385), .A(n15178), .ZN(n15180) );
  INV_X1 U18377 ( .A(n15180), .ZN(P2_U2897) );
  NAND2_X1 U18378 ( .A1(n16417), .A2(n15181), .ZN(n15182) );
  OAI21_X1 U18379 ( .B1(n19357), .B2(n15183), .A(n15182), .ZN(n15187) );
  INV_X1 U18380 ( .A(n16418), .ZN(n15208) );
  INV_X1 U18381 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n15185) );
  INV_X1 U18382 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n15184) );
  OAI22_X1 U18383 ( .A1(n15208), .A2(n15185), .B1(n15206), .B2(n15184), .ZN(
        n15186) );
  AOI211_X1 U18384 ( .C1(n19383), .C2(n15526), .A(n15187), .B(n15186), .ZN(
        n15188) );
  OAI21_X1 U18385 ( .B1(n15189), .B2(n15230), .A(n15188), .ZN(P2_U2898) );
  OR2_X1 U18386 ( .A1(n15190), .A2(n15200), .ZN(n15191) );
  NAND2_X1 U18387 ( .A1(n15192), .A2(n15191), .ZN(n19193) );
  AOI22_X1 U18388 ( .A1(n16418), .A2(BUF2_REG_20__SCAN_IN), .B1(n16419), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n15195) );
  AOI22_X1 U18389 ( .A1(n16417), .A2(n15193), .B1(n19382), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n15194) );
  OAI211_X1 U18390 ( .C1(n19358), .C2(n19193), .A(n15195), .B(n15194), .ZN(
        n15196) );
  AOI21_X1 U18391 ( .B1(n15197), .B2(n19385), .A(n15196), .ZN(n15198) );
  INV_X1 U18392 ( .A(n15198), .ZN(P2_U2899) );
  AOI21_X1 U18393 ( .B1(n15201), .B2(n15199), .A(n15200), .ZN(n19202) );
  NAND2_X1 U18394 ( .A1(n16417), .A2(n15202), .ZN(n15203) );
  OAI21_X1 U18395 ( .B1(n19357), .B2(n15204), .A(n15203), .ZN(n15210) );
  INV_X1 U18396 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n15207) );
  INV_X1 U18397 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n15205) );
  OAI22_X1 U18398 ( .A1(n15208), .A2(n15207), .B1(n15206), .B2(n15205), .ZN(
        n15209) );
  AOI211_X1 U18399 ( .C1(n19383), .C2(n19202), .A(n15210), .B(n15209), .ZN(
        n15211) );
  OAI21_X1 U18400 ( .B1(n15212), .B2(n15230), .A(n15211), .ZN(P2_U2900) );
  OR2_X1 U18401 ( .A1(n15224), .A2(n15213), .ZN(n15214) );
  NAND2_X1 U18402 ( .A1(n15214), .A2(n15199), .ZN(n19219) );
  AOI22_X1 U18403 ( .A1(n16418), .A2(BUF2_REG_18__SCAN_IN), .B1(n16419), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n15217) );
  AOI22_X1 U18404 ( .A1(n16417), .A2(n15215), .B1(n19382), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n15216) );
  OAI211_X1 U18405 ( .C1(n19358), .C2(n19219), .A(n15217), .B(n15216), .ZN(
        n15218) );
  AOI21_X1 U18406 ( .B1(n15219), .B2(n19385), .A(n15218), .ZN(n15220) );
  INV_X1 U18407 ( .A(n15220), .ZN(P2_U2901) );
  NOR2_X1 U18408 ( .A1(n15221), .A2(n15222), .ZN(n15223) );
  OR2_X1 U18409 ( .A1(n15224), .A2(n15223), .ZN(n19226) );
  AOI22_X1 U18410 ( .A1(n16418), .A2(BUF2_REG_17__SCAN_IN), .B1(n16419), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n15227) );
  AOI22_X1 U18411 ( .A1(n16417), .A2(n15225), .B1(n19382), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n15226) );
  OAI211_X1 U18412 ( .C1(n19358), .C2(n19226), .A(n15227), .B(n15226), .ZN(
        n15228) );
  INV_X1 U18413 ( .A(n15228), .ZN(n15229) );
  OAI21_X1 U18414 ( .B1(n15231), .B2(n15230), .A(n15229), .ZN(P2_U2902) );
  NOR2_X1 U18415 ( .A1(n15232), .A2(n15241), .ZN(n15233) );
  OR2_X1 U18416 ( .A1(n15221), .A2(n15233), .ZN(n19242) );
  AOI22_X1 U18417 ( .A1(n16418), .A2(BUF2_REG_16__SCAN_IN), .B1(n16419), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n15236) );
  AOI22_X1 U18418 ( .A1(n16417), .A2(n15234), .B1(n19382), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n15235) );
  OAI211_X1 U18419 ( .C1(n19358), .C2(n19242), .A(n15236), .B(n15235), .ZN(
        n15237) );
  AOI21_X1 U18420 ( .B1(n15238), .B2(n19385), .A(n15237), .ZN(n15239) );
  INV_X1 U18421 ( .A(n15239), .ZN(P2_U2903) );
  AOI21_X1 U18422 ( .B1(n15242), .B2(n15240), .A(n15241), .ZN(n19251) );
  INV_X1 U18423 ( .A(n19251), .ZN(n15244) );
  INV_X1 U18424 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19393) );
  OAI222_X1 U18425 ( .A1(n15244), .A2(n19355), .B1(n19357), .B2(n19393), .C1(
        n15243), .C2(n19389), .ZN(P2_U2904) );
  NAND2_X1 U18426 ( .A1(n15246), .A2(n15245), .ZN(n15248) );
  XOR2_X1 U18427 ( .A(n15248), .B(n15247), .Z(n15437) );
  INV_X1 U18428 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n15249) );
  NOR2_X1 U18429 ( .A1(n19300), .A2(n15249), .ZN(n15433) );
  AOI21_X1 U18430 ( .B1(n16477), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15433), .ZN(n15252) );
  NAND2_X1 U18431 ( .A1(n19426), .A2(n15250), .ZN(n15251) );
  OAI211_X1 U18432 ( .C1(n16348), .C2(n16433), .A(n15252), .B(n15251), .ZN(
        n15253) );
  AOI21_X1 U18433 ( .B1(n15436), .B2(n16496), .A(n15253), .ZN(n15254) );
  OAI21_X1 U18434 ( .B1(n15437), .B2(n19431), .A(n15254), .ZN(P2_U2985) );
  AOI21_X1 U18435 ( .B1(n15259), .B2(n15258), .A(n15257), .ZN(n15260) );
  XOR2_X1 U18436 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n15261), .Z(
        n15262) );
  XNOR2_X1 U18437 ( .A(n15263), .B(n15262), .ZN(n15449) );
  INV_X1 U18438 ( .A(n15438), .ZN(n15268) );
  NOR2_X1 U18439 ( .A1(n19300), .A2(n20036), .ZN(n15439) );
  AOI21_X1 U18440 ( .B1(n16477), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15439), .ZN(n15264) );
  OAI21_X1 U18441 ( .B1(n16491), .B2(n16366), .A(n15264), .ZN(n15265) );
  INV_X1 U18442 ( .A(n15266), .ZN(n15267) );
  OAI21_X1 U18443 ( .B1(n15449), .B2(n19431), .A(n15269), .ZN(P2_U2986) );
  NAND2_X1 U18444 ( .A1(n15450), .A2(n16495), .ZN(n15277) );
  INV_X1 U18445 ( .A(n16374), .ZN(n15276) );
  NAND2_X1 U18446 ( .A1(n19426), .A2(n15271), .ZN(n15272) );
  NAND2_X1 U18447 ( .A1(n19427), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15456) );
  OAI211_X1 U18448 ( .C1(n19438), .C2(n15273), .A(n15272), .B(n15456), .ZN(
        n15275) );
  INV_X1 U18449 ( .A(n15274), .ZN(n15285) );
  NOR2_X1 U18450 ( .A1(n15278), .A2(n15291), .ZN(n15280) );
  MUX2_X1 U18451 ( .A(n15280), .B(n15291), .S(n15279), .Z(n15282) );
  AOI21_X1 U18452 ( .B1(n15283), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15284) );
  NOR2_X1 U18453 ( .A1(n15285), .A2(n15284), .ZN(n15471) );
  INV_X1 U18454 ( .A(n16389), .ZN(n15287) );
  NAND2_X1 U18455 ( .A1(n19427), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15464) );
  OAI21_X1 U18456 ( .B1(n19438), .B2(n10168), .A(n15464), .ZN(n15286) );
  AOI21_X1 U18457 ( .B1(n19426), .B2(n15287), .A(n15286), .ZN(n15288) );
  OAI21_X1 U18458 ( .B1(n16384), .B2(n16433), .A(n15288), .ZN(n15289) );
  AOI21_X1 U18459 ( .B1(n15471), .B2(n16496), .A(n15289), .ZN(n15290) );
  OAI21_X1 U18460 ( .B1(n19431), .B2(n15473), .A(n15290), .ZN(P2_U2988) );
  XNOR2_X1 U18461 ( .A(n15283), .B(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15485) );
  NOR2_X1 U18462 ( .A1(n15292), .A2(n15291), .ZN(n15293) );
  XNOR2_X1 U18463 ( .A(n15294), .B(n15293), .ZN(n15483) );
  NAND2_X1 U18464 ( .A1(n19427), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15474) );
  OAI21_X1 U18465 ( .B1(n19438), .B2(n15295), .A(n15474), .ZN(n15296) );
  AOI21_X1 U18466 ( .B1(n19426), .B2(n15297), .A(n15296), .ZN(n15298) );
  OAI21_X1 U18467 ( .B1(n16396), .B2(n16433), .A(n15298), .ZN(n15299) );
  AOI21_X1 U18468 ( .B1(n15483), .B2(n16495), .A(n15299), .ZN(n15300) );
  OAI21_X1 U18469 ( .B1(n15485), .B2(n19429), .A(n15300), .ZN(P2_U2989) );
  INV_X1 U18470 ( .A(n15283), .ZN(n15302) );
  OAI21_X1 U18471 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15301), .A(
        n15302), .ZN(n15497) );
  XNOR2_X1 U18472 ( .A(n15304), .B(n10218), .ZN(n15305) );
  XNOR2_X1 U18473 ( .A(n15303), .B(n15305), .ZN(n15495) );
  NOR2_X1 U18474 ( .A1(n16407), .A2(n16433), .ZN(n15308) );
  NAND2_X1 U18475 ( .A1(n19427), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n15487) );
  NAND2_X1 U18476 ( .A1(n16477), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15306) );
  OAI211_X1 U18477 ( .C1(n16491), .C2(n16411), .A(n15487), .B(n15306), .ZN(
        n15307) );
  AOI211_X1 U18478 ( .C1(n15495), .C2(n16495), .A(n15308), .B(n15307), .ZN(
        n15309) );
  OAI21_X1 U18479 ( .B1(n15497), .B2(n19429), .A(n15309), .ZN(P2_U2990) );
  OAI21_X1 U18480 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n9753), .A(
        n10142), .ZN(n15511) );
  XOR2_X1 U18481 ( .A(n15311), .B(n15310), .Z(n15509) );
  NOR2_X1 U18482 ( .A1(n15498), .A2(n16433), .ZN(n15315) );
  NAND2_X1 U18483 ( .A1(n19427), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n15502) );
  NAND2_X1 U18484 ( .A1(n16477), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15312) );
  OAI211_X1 U18485 ( .C1(n16491), .C2(n15313), .A(n15502), .B(n15312), .ZN(
        n15314) );
  AOI211_X1 U18486 ( .C1(n15509), .C2(n16495), .A(n15315), .B(n15314), .ZN(
        n15316) );
  OAI21_X1 U18487 ( .B1(n15511), .B2(n19429), .A(n15316), .ZN(P2_U2991) );
  NAND2_X1 U18488 ( .A1(n15318), .A2(n15317), .ZN(n15320) );
  XOR2_X1 U18489 ( .A(n15320), .B(n15319), .Z(n15522) );
  AOI21_X1 U18490 ( .B1(n15515), .B2(n15321), .A(n9753), .ZN(n15512) );
  NAND2_X1 U18491 ( .A1(n15512), .A2(n16496), .ZN(n15325) );
  NOR2_X1 U18492 ( .A1(n19300), .A2(n20024), .ZN(n15514) );
  AOI21_X1 U18493 ( .B1(n16477), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15514), .ZN(n15322) );
  OAI21_X1 U18494 ( .B1(n16491), .B2(n16057), .A(n15322), .ZN(n15323) );
  AOI21_X1 U18495 ( .B1(n16048), .B2(n19435), .A(n15323), .ZN(n15324) );
  OAI211_X1 U18496 ( .C1(n15522), .C2(n19431), .A(n15325), .B(n15324), .ZN(
        P2_U2992) );
  NAND2_X1 U18497 ( .A1(n15327), .A2(n15326), .ZN(n15334) );
  NAND2_X1 U18498 ( .A1(n15329), .A2(n16451), .ZN(n15597) );
  INV_X1 U18499 ( .A(n15594), .ZN(n15330) );
  AOI21_X1 U18500 ( .B1(n15597), .B2(n15595), .A(n15330), .ZN(n16437) );
  INV_X1 U18501 ( .A(n15331), .ZN(n15332) );
  NOR2_X1 U18502 ( .A1(n19300), .A2(n20022), .ZN(n15525) );
  AOI21_X1 U18503 ( .B1(n16477), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15525), .ZN(n15335) );
  OAI21_X1 U18504 ( .B1(n16491), .B2(n15336), .A(n15335), .ZN(n15339) );
  OAI21_X1 U18505 ( .B1(n15337), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15321), .ZN(n15530) );
  NOR2_X1 U18506 ( .A1(n15530), .A2(n19429), .ZN(n15338) );
  AOI211_X1 U18507 ( .C1(n19435), .C2(n15533), .A(n15339), .B(n15338), .ZN(
        n15340) );
  OAI21_X1 U18508 ( .B1(n15535), .B2(n19431), .A(n15340), .ZN(P2_U2993) );
  AND2_X1 U18509 ( .A1(n15342), .A2(n15341), .ZN(n15343) );
  OAI22_X1 U18510 ( .A1(n15344), .A2(n10039), .B1(n9722), .B2(n15343), .ZN(
        n15544) );
  NAND2_X1 U18511 ( .A1(n9653), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15360) );
  AOI21_X1 U18512 ( .B1(n15346), .B2(n15360), .A(n15337), .ZN(n15541) );
  NOR2_X1 U18513 ( .A1(n19189), .A2(n16433), .ZN(n15350) );
  NAND2_X1 U18514 ( .A1(n19427), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n15538) );
  NAND2_X1 U18515 ( .A1(n16477), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15347) );
  OAI211_X1 U18516 ( .C1(n16491), .C2(n15348), .A(n15538), .B(n15347), .ZN(
        n15349) );
  AOI211_X1 U18517 ( .C1(n15541), .C2(n16496), .A(n15350), .B(n15349), .ZN(
        n15351) );
  OAI21_X1 U18518 ( .B1(n15544), .B2(n19431), .A(n15351), .ZN(P2_U2994) );
  INV_X1 U18519 ( .A(n15364), .ZN(n15352) );
  AOI21_X1 U18520 ( .B1(n15365), .B2(n15363), .A(n15352), .ZN(n15356) );
  NAND2_X1 U18521 ( .A1(n15354), .A2(n15353), .ZN(n15355) );
  XNOR2_X1 U18522 ( .A(n15356), .B(n15355), .ZN(n15555) );
  OAI22_X1 U18523 ( .A1(n19438), .A2(n19197), .B1(n15357), .B2(n19300), .ZN(
        n15359) );
  NOR2_X1 U18524 ( .A1(n19201), .A2(n16433), .ZN(n15358) );
  AOI211_X1 U18525 ( .C1(n19426), .C2(n19196), .A(n15359), .B(n15358), .ZN(
        n15362) );
  OAI21_X1 U18526 ( .B1(n9653), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15360), .ZN(n15550) );
  OR2_X1 U18527 ( .A1(n15550), .A2(n19429), .ZN(n15361) );
  OAI211_X1 U18528 ( .C1(n15555), .C2(n19431), .A(n15362), .B(n15361), .ZN(
        P2_U2995) );
  NAND2_X1 U18529 ( .A1(n15364), .A2(n15363), .ZN(n15366) );
  XOR2_X1 U18530 ( .A(n15366), .B(n15365), .Z(n15565) );
  OAI21_X1 U18531 ( .B1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n9752), .A(
        n15345), .ZN(n15561) );
  INV_X1 U18532 ( .A(n15561), .ZN(n15371) );
  OAI22_X1 U18533 ( .A1(n20017), .A2(n19300), .B1(n16491), .B2(n15367), .ZN(
        n15370) );
  INV_X1 U18534 ( .A(n19215), .ZN(n15368) );
  OAI22_X1 U18535 ( .A1(n15368), .A2(n16433), .B1(n10163), .B2(n19438), .ZN(
        n15369) );
  AOI211_X1 U18536 ( .C1(n15371), .C2(n16496), .A(n15370), .B(n15369), .ZN(
        n15372) );
  OAI21_X1 U18537 ( .B1(n15565), .B2(n19431), .A(n15372), .ZN(P2_U2996) );
  XNOR2_X1 U18538 ( .A(n9701), .B(n15373), .ZN(n15591) );
  NOR2_X1 U18539 ( .A1(n15584), .A2(n19300), .ZN(n15376) );
  OAI22_X1 U18540 ( .A1(n10162), .A2(n19438), .B1(n16491), .B2(n15374), .ZN(
        n15375) );
  AOI211_X1 U18541 ( .C1(n19435), .C2(n19238), .A(n15376), .B(n15375), .ZN(
        n15380) );
  NOR2_X1 U18542 ( .A1(n15377), .A2(n16505), .ZN(n15566) );
  XNOR2_X1 U18543 ( .A(n15566), .B(n15577), .ZN(n15378) );
  NAND2_X1 U18544 ( .A1(n15378), .A2(n16496), .ZN(n15379) );
  OAI211_X1 U18545 ( .C1(n15591), .C2(n19431), .A(n15380), .B(n15379), .ZN(
        P2_U2998) );
  AOI21_X1 U18546 ( .B1(n15382), .B2(n15381), .A(n9748), .ZN(n16567) );
  NAND2_X1 U18547 ( .A1(n15383), .A2(n15398), .ZN(n15384) );
  NAND2_X1 U18548 ( .A1(n15384), .A2(n15399), .ZN(n15388) );
  AND2_X1 U18549 ( .A1(n15386), .A2(n15385), .ZN(n15387) );
  XNOR2_X1 U18550 ( .A(n15388), .B(n15387), .ZN(n16571) );
  AOI22_X1 U18551 ( .A1(n19435), .A2(n19296), .B1(n16477), .B2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n15392) );
  OAI22_X1 U18552 ( .A1(n10710), .A2(n19300), .B1(n16491), .B2(n15389), .ZN(
        n15390) );
  INV_X1 U18553 ( .A(n15390), .ZN(n15391) );
  OAI211_X1 U18554 ( .C1(n16571), .C2(n19431), .A(n15392), .B(n15391), .ZN(
        n15393) );
  AOI21_X1 U18555 ( .B1(n16567), .B2(n16496), .A(n15393), .ZN(n15394) );
  INV_X1 U18556 ( .A(n15394), .ZN(P2_U3006) );
  XNOR2_X1 U18557 ( .A(n15396), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15397) );
  XNOR2_X1 U18558 ( .A(n15395), .B(n15397), .ZN(n15646) );
  NAND2_X1 U18559 ( .A1(n15399), .A2(n15398), .ZN(n15400) );
  XNOR2_X1 U18560 ( .A(n15383), .B(n15400), .ZN(n15644) );
  OAI22_X1 U18561 ( .A1(n10706), .A2(n19438), .B1(n16491), .B2(n15401), .ZN(
        n15404) );
  OAI22_X1 U18562 ( .A1(n16433), .A2(n15640), .B1(n19300), .B2(n15402), .ZN(
        n15403) );
  AOI211_X1 U18563 ( .C1(n15644), .C2(n16495), .A(n15404), .B(n15403), .ZN(
        n15405) );
  OAI21_X1 U18564 ( .B1(n15646), .B2(n19429), .A(n15405), .ZN(P2_U3007) );
  OAI21_X1 U18565 ( .B1(n15407), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n15406), .ZN(n15655) );
  XOR2_X1 U18566 ( .A(n15408), .B(n15410), .Z(n15653) );
  OAI22_X1 U18567 ( .A1(n15411), .A2(n19438), .B1(n10860), .B2(n19300), .ZN(
        n15414) );
  INV_X1 U18568 ( .A(n19312), .ZN(n15412) );
  OAI22_X1 U18569 ( .A1(n16433), .A2(n15648), .B1(n16491), .B2(n15412), .ZN(
        n15413) );
  AOI211_X1 U18570 ( .C1(n15653), .C2(n16495), .A(n15414), .B(n15413), .ZN(
        n15415) );
  OAI21_X1 U18571 ( .B1(n15655), .B2(n19429), .A(n15415), .ZN(P2_U3008) );
  XNOR2_X1 U18572 ( .A(n15417), .B(n15416), .ZN(n15667) );
  OR2_X1 U18573 ( .A1(n15419), .A2(n15418), .ZN(n15420) );
  AOI22_X1 U18574 ( .A1(n15423), .A2(n15422), .B1(n15421), .B2(n15420), .ZN(
        n15665) );
  OAI22_X1 U18575 ( .A1(n10699), .A2(n19438), .B1(n16491), .B2(n15424), .ZN(
        n15428) );
  INV_X1 U18576 ( .A(n15425), .ZN(n15661) );
  OAI22_X1 U18577 ( .A1(n16433), .A2(n15661), .B1(n19300), .B2(n15426), .ZN(
        n15427) );
  AOI211_X1 U18578 ( .C1(n15665), .C2(n16496), .A(n15428), .B(n15427), .ZN(
        n15429) );
  OAI21_X1 U18579 ( .B1(n19431), .B2(n15667), .A(n15429), .ZN(P2_U3009) );
  NOR2_X1 U18580 ( .A1(n16348), .A2(n16574), .ZN(n15435) );
  INV_X1 U18581 ( .A(n15431), .ZN(n15454) );
  NOR3_X1 U18582 ( .A1(n15431), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15430), .ZN(n15432) );
  AOI21_X1 U18583 ( .B1(n15454), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15442) );
  AOI21_X1 U18584 ( .B1(n16582), .B2(n15440), .A(n15439), .ZN(n15441) );
  INV_X1 U18585 ( .A(n15444), .ZN(n15446) );
  NAND2_X1 U18586 ( .A1(n16363), .A2(n16592), .ZN(n15445) );
  NAND2_X1 U18587 ( .A1(n15446), .A2(n15445), .ZN(n15447) );
  OAI21_X1 U18588 ( .B1(n15449), .B2(n16570), .A(n15448), .ZN(P2_U3018) );
  NAND2_X1 U18589 ( .A1(n15450), .A2(n16584), .ZN(n15462) );
  OR3_X1 U18590 ( .A1(n15452), .A2(n15451), .A3(n16587), .ZN(n15461) );
  NAND2_X1 U18591 ( .A1(n15454), .A2(n15453), .ZN(n15455) );
  OAI211_X1 U18592 ( .C1(n16563), .C2(n16373), .A(n15456), .B(n15455), .ZN(
        n15458) );
  NOR2_X1 U18593 ( .A1(n16374), .A2(n16574), .ZN(n15457) );
  AOI211_X1 U18594 ( .C1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n15459), .A(
        n15458), .B(n15457), .ZN(n15460) );
  OAI211_X1 U18595 ( .C1(n15463), .C2(n15462), .A(n15461), .B(n15460), .ZN(
        P2_U3019) );
  NOR2_X1 U18596 ( .A1(n16384), .A2(n16574), .ZN(n15470) );
  INV_X1 U18597 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15468) );
  XNOR2_X1 U18598 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15465) );
  OAI21_X1 U18599 ( .B1(n15475), .B2(n15465), .A(n15464), .ZN(n15466) );
  AOI21_X1 U18600 ( .B1(n16582), .B2(n16385), .A(n15466), .ZN(n15467) );
  OAI21_X1 U18601 ( .B1(n15481), .B2(n15468), .A(n15467), .ZN(n15469) );
  AOI211_X1 U18602 ( .C1(n15471), .C2(n16566), .A(n15470), .B(n15469), .ZN(
        n15472) );
  OAI21_X1 U18603 ( .B1(n16570), .B2(n15473), .A(n15472), .ZN(P2_U3020) );
  OAI21_X1 U18604 ( .B1(n15475), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15474), .ZN(n15477) );
  NOR2_X1 U18605 ( .A1(n16396), .A2(n16574), .ZN(n15476) );
  AOI211_X1 U18606 ( .C1(n16582), .C2(n15478), .A(n15477), .B(n15476), .ZN(
        n15479) );
  OAI21_X1 U18607 ( .B1(n15481), .B2(n15480), .A(n15479), .ZN(n15482) );
  AOI21_X1 U18608 ( .B1(n15483), .B2(n16584), .A(n15482), .ZN(n15484) );
  OAI21_X1 U18609 ( .B1(n15485), .B2(n16587), .A(n15484), .ZN(P2_U3021) );
  NOR2_X1 U18610 ( .A1(n15486), .A2(n10218), .ZN(n15494) );
  INV_X1 U18611 ( .A(n15487), .ZN(n15488) );
  AOI21_X1 U18612 ( .B1(n15489), .B2(n10218), .A(n15488), .ZN(n15492) );
  NAND2_X1 U18613 ( .A1(n16582), .A2(n15490), .ZN(n15491) );
  OAI211_X1 U18614 ( .C1(n16407), .C2(n16574), .A(n15492), .B(n15491), .ZN(
        n15493) );
  AOI211_X1 U18615 ( .C1(n15495), .C2(n16584), .A(n15494), .B(n15493), .ZN(
        n15496) );
  OAI21_X1 U18616 ( .B1(n15497), .B2(n16587), .A(n15496), .ZN(P2_U3022) );
  INV_X1 U18617 ( .A(n15498), .ZN(n15505) );
  INV_X1 U18618 ( .A(n15499), .ZN(n15516) );
  OAI211_X1 U18619 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15516), .B(n15500), .ZN(
        n15501) );
  OAI211_X1 U18620 ( .C1(n16563), .C2(n15503), .A(n15502), .B(n15501), .ZN(
        n15504) );
  AOI21_X1 U18621 ( .B1(n15505), .B2(n16592), .A(n15504), .ZN(n15506) );
  OAI21_X1 U18622 ( .B1(n15507), .B2(n15513), .A(n15506), .ZN(n15508) );
  AOI21_X1 U18623 ( .B1(n15509), .B2(n16584), .A(n15508), .ZN(n15510) );
  OAI21_X1 U18624 ( .B1(n15511), .B2(n16587), .A(n15510), .ZN(P2_U3023) );
  NAND2_X1 U18625 ( .A1(n15512), .A2(n16566), .ZN(n15521) );
  NOR2_X1 U18626 ( .A1(n15513), .A2(n15515), .ZN(n15519) );
  AOI21_X1 U18627 ( .B1(n15516), .B2(n15515), .A(n15514), .ZN(n15517) );
  OAI21_X1 U18628 ( .B1(n16563), .B2(n16060), .A(n15517), .ZN(n15518) );
  AOI211_X1 U18629 ( .C1(n16048), .C2(n16592), .A(n15519), .B(n15518), .ZN(
        n15520) );
  OAI211_X1 U18630 ( .C1(n15522), .C2(n16570), .A(n15521), .B(n15520), .ZN(
        P2_U3024) );
  INV_X1 U18631 ( .A(n15523), .ZN(n15529) );
  AOI21_X1 U18632 ( .B1(n15545), .B2(n15524), .A(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15528) );
  AOI21_X1 U18633 ( .B1(n16582), .B2(n15526), .A(n15525), .ZN(n15527) );
  OAI21_X1 U18634 ( .B1(n15529), .B2(n15528), .A(n15527), .ZN(n15532) );
  NOR2_X1 U18635 ( .A1(n15530), .A2(n16587), .ZN(n15531) );
  AOI211_X1 U18636 ( .C1(n16592), .C2(n15533), .A(n15532), .B(n15531), .ZN(
        n15534) );
  OAI211_X1 U18637 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n15545), .B(n15536), .ZN(
        n15537) );
  OAI211_X1 U18638 ( .C1(n16563), .C2(n19193), .A(n15538), .B(n15537), .ZN(
        n15540) );
  NOR2_X1 U18639 ( .A1(n19189), .A2(n16574), .ZN(n15539) );
  AOI211_X1 U18640 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n15553), .A(
        n15540), .B(n15539), .ZN(n15543) );
  NAND2_X1 U18641 ( .A1(n15541), .A2(n16566), .ZN(n15542) );
  OAI211_X1 U18642 ( .C1(n15544), .C2(n16570), .A(n15543), .B(n15542), .ZN(
        P2_U3026) );
  INV_X1 U18643 ( .A(n15545), .ZN(n15547) );
  NAND2_X1 U18644 ( .A1(P2_REIP_REG_19__SCAN_IN), .A2(n19427), .ZN(n15546) );
  OAI21_X1 U18645 ( .B1(n15547), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15546), .ZN(n15548) );
  AOI21_X1 U18646 ( .B1(n16582), .B2(n19202), .A(n15548), .ZN(n15549) );
  OAI21_X1 U18647 ( .B1(n19201), .B2(n16574), .A(n15549), .ZN(n15552) );
  NOR2_X1 U18648 ( .A1(n15550), .A2(n16587), .ZN(n15551) );
  AOI211_X1 U18649 ( .C1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15553), .A(
        n15552), .B(n15551), .ZN(n15554) );
  OAI21_X1 U18650 ( .B1(n15555), .B2(n16570), .A(n15554), .ZN(P2_U3027) );
  NOR2_X1 U18651 ( .A1(n20017), .A2(n19300), .ZN(n15558) );
  NOR3_X1 U18652 ( .A1(n15556), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n16502), .ZN(n15557) );
  AOI211_X1 U18653 ( .C1(n15559), .C2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15558), .B(n15557), .ZN(n15560) );
  OAI21_X1 U18654 ( .B1(n16563), .B2(n19219), .A(n15560), .ZN(n15563) );
  NOR2_X1 U18655 ( .A1(n15561), .A2(n16587), .ZN(n15562) );
  AOI211_X1 U18656 ( .C1(n19215), .C2(n16592), .A(n15563), .B(n15562), .ZN(
        n15564) );
  OAI21_X1 U18657 ( .B1(n15565), .B2(n16570), .A(n15564), .ZN(P2_U3028) );
  NAND2_X1 U18658 ( .A1(n15566), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16425) );
  OAI21_X1 U18659 ( .B1(n16566), .B2(n15567), .A(n16425), .ZN(n15568) );
  OAI211_X1 U18660 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15569), .A(
        n15568), .B(n16506), .ZN(n15589) );
  AOI21_X1 U18661 ( .B1(n15577), .B2(n15570), .A(n15589), .ZN(n15583) );
  NAND2_X1 U18662 ( .A1(n15572), .A2(n15571), .ZN(n15574) );
  XOR2_X1 U18663 ( .A(n15574), .B(n15573), .Z(n16431) );
  NAND2_X1 U18664 ( .A1(n16431), .A2(n16584), .ZN(n15582) );
  INV_X1 U18665 ( .A(n19227), .ZN(n15580) );
  OAI22_X1 U18666 ( .A1(n16563), .A2(n19226), .B1(n15575), .B2(n19300), .ZN(
        n15579) );
  OAI21_X1 U18667 ( .B1(n15377), .B2(n16587), .A(n16502), .ZN(n15576) );
  NAND2_X1 U18668 ( .A1(n15576), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15587) );
  NOR3_X1 U18669 ( .A1(n15587), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15577), .ZN(n15578) );
  AOI211_X1 U18670 ( .C1(n16592), .C2(n15580), .A(n15579), .B(n15578), .ZN(
        n15581) );
  OAI211_X1 U18671 ( .C1(n15583), .C2(n16426), .A(n15582), .B(n15581), .ZN(
        P2_U3029) );
  OAI22_X1 U18672 ( .A1(n16563), .A2(n19242), .B1(n15584), .B2(n19300), .ZN(
        n15585) );
  AOI21_X1 U18673 ( .B1(n19238), .B2(n16592), .A(n15585), .ZN(n15586) );
  OAI21_X1 U18674 ( .B1(n15587), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n15586), .ZN(n15588) );
  AOI21_X1 U18675 ( .B1(n15589), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n15588), .ZN(n15590) );
  OAI21_X1 U18676 ( .B1(n15591), .B2(n16570), .A(n15590), .ZN(P2_U3030) );
  NOR2_X1 U18677 ( .A1(n15592), .A2(n16545), .ZN(n16479) );
  NAND2_X1 U18678 ( .A1(n16479), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16448) );
  INV_X1 U18679 ( .A(n15599), .ZN(n15593) );
  NOR2_X1 U18680 ( .A1(n16448), .A2(n15593), .ZN(n16449) );
  OAI21_X1 U18681 ( .B1(n16449), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n15377), .ZN(n16442) );
  AND2_X1 U18682 ( .A1(n15595), .A2(n15594), .ZN(n15596) );
  XNOR2_X1 U18683 ( .A(n15597), .B(n15596), .ZN(n16441) );
  INV_X1 U18684 ( .A(n16532), .ZN(n15598) );
  OR2_X1 U18685 ( .A1(n15598), .A2(n16546), .ZN(n16514) );
  OAI21_X1 U18686 ( .B1(n15598), .B2(n16525), .A(n16526), .ZN(n15612) );
  OAI21_X1 U18687 ( .B1(n15599), .B2(n16514), .A(n15612), .ZN(n16517) );
  NOR2_X1 U18688 ( .A1(n10947), .A2(n19300), .ZN(n15600) );
  AOI221_X1 U18689 ( .B1(n15602), .B2(n15601), .C1(n16517), .C2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(n15600), .ZN(n15608) );
  INV_X1 U18690 ( .A(n15603), .ZN(n19262) );
  OR2_X1 U18691 ( .A1(n15604), .A2(n14858), .ZN(n15605) );
  NAND2_X1 U18692 ( .A1(n15605), .A2(n15240), .ZN(n19343) );
  INV_X1 U18693 ( .A(n19343), .ZN(n15606) );
  AOI22_X1 U18694 ( .A1(n19262), .A2(n16592), .B1(n16582), .B2(n15606), .ZN(
        n15607) );
  OAI211_X1 U18695 ( .C1(n16441), .C2(n16570), .A(n15608), .B(n15607), .ZN(
        n15609) );
  INV_X1 U18696 ( .A(n15609), .ZN(n15610) );
  OAI21_X1 U18697 ( .B1(n16442), .B2(n16587), .A(n15610), .ZN(P2_U3032) );
  XNOR2_X1 U18698 ( .A(n16448), .B(n16515), .ZN(n16460) );
  NAND2_X1 U18699 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n19427), .ZN(n15611) );
  OAI221_X1 U18700 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16514), 
        .C1(n16515), .C2(n15612), .A(n15611), .ZN(n15615) );
  INV_X1 U18701 ( .A(n19274), .ZN(n15613) );
  OAI22_X1 U18702 ( .A1(n16574), .A2(n15613), .B1(n16563), .B2(n19272), .ZN(
        n15614) );
  NOR2_X1 U18703 ( .A1(n15615), .A2(n15614), .ZN(n15621) );
  NOR2_X1 U18704 ( .A1(n10067), .A2(n15618), .ZN(n15619) );
  XNOR2_X1 U18705 ( .A(n15616), .B(n15619), .ZN(n16459) );
  OR2_X1 U18706 ( .A1(n16459), .A2(n16570), .ZN(n15620) );
  OAI211_X1 U18707 ( .C1(n16460), .C2(n16587), .A(n15621), .B(n15620), .ZN(
        P2_U3034) );
  INV_X1 U18708 ( .A(n15592), .ZN(n15623) );
  AOI21_X1 U18709 ( .B1(n9912), .B2(n15624), .A(n15623), .ZN(n16497) );
  NAND2_X1 U18710 ( .A1(n16497), .A2(n16566), .ZN(n15638) );
  OAI22_X1 U18711 ( .A1(n16574), .A2(n15626), .B1(n15625), .B2(n19300), .ZN(
        n15629) );
  NOR2_X1 U18712 ( .A1(n16563), .A2(n15627), .ZN(n15628) );
  NOR2_X1 U18713 ( .A1(n15629), .A2(n15628), .ZN(n15637) );
  INV_X1 U18714 ( .A(n15631), .ZN(n16480) );
  NOR2_X1 U18715 ( .A1(n15632), .A2(n16480), .ZN(n15633) );
  XNOR2_X1 U18716 ( .A(n15630), .B(n15633), .ZN(n16494) );
  NAND2_X1 U18717 ( .A1(n16494), .A2(n16584), .ZN(n15636) );
  OAI21_X1 U18718 ( .B1(n15634), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n16525), .ZN(n15635) );
  NAND4_X1 U18719 ( .A1(n15638), .A2(n15637), .A3(n15636), .A4(n15635), .ZN(
        P2_U3037) );
  NAND2_X1 U18720 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19427), .ZN(n15639) );
  OAI221_X1 U18721 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16556), .C1(
        n16558), .C2(n16562), .A(n15639), .ZN(n15643) );
  OAI22_X1 U18722 ( .A1(n15641), .A2(n16563), .B1(n16574), .B2(n15640), .ZN(
        n15642) );
  AOI211_X1 U18723 ( .C1(n15644), .C2(n16584), .A(n15643), .B(n15642), .ZN(
        n15645) );
  OAI21_X1 U18724 ( .B1(n15646), .B2(n16587), .A(n15645), .ZN(P2_U3039) );
  NAND2_X1 U18725 ( .A1(n15647), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15650) );
  INV_X1 U18726 ( .A(n15648), .ZN(n19313) );
  AOI22_X1 U18727 ( .A1(n16592), .A2(n19313), .B1(n19427), .B2(
        P2_REIP_REG_6__SCAN_IN), .ZN(n15649) );
  OAI211_X1 U18728 ( .C1(n16563), .C2(n19319), .A(n15650), .B(n15649), .ZN(
        n15651) );
  AOI211_X1 U18729 ( .C1(n15653), .C2(n16584), .A(n15652), .B(n15651), .ZN(
        n15654) );
  OAI21_X1 U18730 ( .B1(n15655), .B2(n16587), .A(n15654), .ZN(P2_U3040) );
  NAND2_X1 U18731 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19427), .ZN(n15659) );
  INV_X1 U18732 ( .A(n15656), .ZN(n15657) );
  OAI211_X1 U18733 ( .C1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(n15677), .B(n15657), .ZN(n15658) );
  OAI211_X1 U18734 ( .C1(n15673), .C2(n15660), .A(n15659), .B(n15658), .ZN(
        n15664) );
  OAI22_X1 U18735 ( .A1(n15662), .A2(n16563), .B1(n16574), .B2(n15661), .ZN(
        n15663) );
  AOI211_X1 U18736 ( .C1(n15665), .C2(n16566), .A(n15664), .B(n15663), .ZN(
        n15666) );
  OAI21_X1 U18737 ( .B1(n16570), .B2(n15667), .A(n15666), .ZN(P2_U3041) );
  OAI21_X1 U18738 ( .B1(n15669), .B2(n15676), .A(n15668), .ZN(n15670) );
  INV_X1 U18739 ( .A(n15670), .ZN(n19430) );
  XOR2_X1 U18740 ( .A(n15671), .B(n15672), .Z(n19428) );
  INV_X1 U18741 ( .A(n15673), .ZN(n15675) );
  NOR2_X1 U18742 ( .A1(n10695), .A2(n19300), .ZN(n15674) );
  AOI221_X1 U18743 ( .B1(n15677), .B2(n15676), .C1(n15675), .C2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n15674), .ZN(n15679) );
  NAND2_X1 U18744 ( .A1(n19434), .A2(n16592), .ZN(n15678) );
  OAI211_X1 U18745 ( .C1(n19359), .C2(n16563), .A(n15679), .B(n15678), .ZN(
        n15680) );
  AOI21_X1 U18746 ( .B1(n19428), .B2(n16584), .A(n15680), .ZN(n15681) );
  OAI21_X1 U18747 ( .B1(n19430), .B2(n16587), .A(n15681), .ZN(P2_U3042) );
  OAI22_X1 U18748 ( .A1(n19310), .A2(n16585), .B1(n19340), .B2(n19244), .ZN(
        n15693) );
  OAI222_X1 U18749 ( .A1(n16602), .A2(n15684), .B1(n20065), .B2(n15683), .C1(
        n10677), .C2(n15693), .ZN(n15689) );
  NOR2_X1 U18750 ( .A1(n15685), .A2(n16605), .ZN(n15688) );
  INV_X1 U18751 ( .A(n16119), .ZN(n16115) );
  NAND2_X1 U18752 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(n16115), .ZN(n15686) );
  OAI21_X1 U18753 ( .B1(n20089), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n15686), 
        .ZN(n15687) );
  OR2_X1 U18754 ( .A1(n15688), .A2(n15687), .ZN(n20061) );
  MUX2_X1 U18755 ( .A(n15690), .B(n15689), .S(n20061), .Z(P2_U3601) );
  OAI21_X1 U18756 ( .B1(n19310), .B2(n15692), .A(n15691), .ZN(n20055) );
  INV_X1 U18757 ( .A(n15693), .ZN(n15694) );
  NOR2_X1 U18758 ( .A1(n15694), .A2(n10677), .ZN(n20056) );
  INV_X1 U18759 ( .A(n16602), .ZN(n20058) );
  AOI222_X1 U18760 ( .A1(n15695), .A2(n20059), .B1(n20055), .B2(n20056), .C1(
        n20058), .C2(n19440), .ZN(n15697) );
  INV_X1 U18761 ( .A(n20061), .ZN(n20063) );
  NAND2_X1 U18762 ( .A1(n20063), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15696) );
  OAI21_X1 U18763 ( .B1(n15697), .B2(n20063), .A(n15696), .ZN(P2_U3599) );
  OAI22_X1 U18764 ( .A1(n19727), .A2(n16602), .B1(n15698), .B2(n20065), .ZN(
        n15699) );
  MUX2_X1 U18765 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n15699), .S(
        n20061), .Z(P2_U3596) );
  NAND2_X1 U18766 ( .A1(n19727), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19671) );
  OAI21_X1 U18767 ( .B1(n19671), .B2(n19835), .A(n20068), .ZN(n15712) );
  INV_X1 U18768 ( .A(n15712), .ZN(n15705) );
  NAND3_X1 U18769 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n10331), .A3(
        n20088), .ZN(n19583) );
  AOI21_X1 U18770 ( .B1(n12531), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n15703) );
  NOR2_X1 U18771 ( .A1(n20096), .A2(n19583), .ZN(n19637) );
  NAND2_X1 U18772 ( .A1(n19591), .A2(n10677), .ZN(n19159) );
  NAND2_X1 U18773 ( .A1(n19974), .A2(n19159), .ZN(n20117) );
  INV_X1 U18774 ( .A(n20117), .ZN(n15700) );
  NAND2_X1 U18775 ( .A1(n15700), .A2(n16596), .ZN(n15701) );
  OAI21_X1 U18776 ( .B1(n15703), .B2(n19637), .A(n19919), .ZN(n15704) );
  INV_X1 U18777 ( .A(n19635), .ZN(n15706) );
  NAND2_X1 U18778 ( .A1(n15706), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n15716) );
  AOI22_X1 U18779 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19480), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19479), .ZN(n19924) );
  INV_X1 U18780 ( .A(n19924), .ZN(n19873) );
  NOR2_X2 U18781 ( .A1(n20115), .A2(n19468), .ZN(n19912) );
  AOI22_X1 U18782 ( .A1(n19662), .A2(n19873), .B1(n19912), .B2(n19637), .ZN(
        n15715) );
  INV_X1 U18783 ( .A(n12531), .ZN(n15710) );
  OAI21_X1 U18784 ( .B1(n15710), .B2(n19637), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15711) );
  OAI21_X1 U18785 ( .B1(n15712), .B2(n19583), .A(n15711), .ZN(n19631) );
  NOR2_X2 U18786 ( .A1(n19390), .A2(n19639), .ZN(n19913) );
  NAND2_X1 U18787 ( .A1(n19631), .A2(n19913), .ZN(n15714) );
  INV_X1 U18788 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n18476) );
  OAI22_X2 U18789 ( .A1(n16691), .A2(n19483), .B1(n18476), .B2(n19481), .ZN(
        n19921) );
  NAND2_X1 U18790 ( .A1(n19921), .A2(n19630), .ZN(n15713) );
  NAND4_X1 U18791 ( .A1(n15716), .A2(n15715), .A3(n15714), .A4(n15713), .ZN(
        P2_U3088) );
  NOR2_X2 U18792 ( .A1(n15717), .A2(n19639), .ZN(n19956) );
  AOI22_X1 U18793 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19480), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19479), .ZN(n19960) );
  AOI22_X1 U18794 ( .A1(n19662), .A2(n19898), .B1(n19637), .B2(n19955), .ZN(
        n15719) );
  INV_X1 U18795 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n17512) );
  NAND2_X1 U18796 ( .A1(n19957), .A2(n19630), .ZN(n15718) );
  OAI211_X1 U18797 ( .C1(n19635), .C2(n15720), .A(n15719), .B(n15718), .ZN(
        n15721) );
  AOI21_X1 U18798 ( .B1(n19956), .B2(n19631), .A(n15721), .ZN(n15722) );
  INV_X1 U18799 ( .A(n15722), .ZN(P2_U3094) );
  NAND2_X1 U18800 ( .A1(n20079), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19781) );
  NOR2_X1 U18801 ( .A1(n19495), .A2(n19781), .ZN(n19752) );
  INV_X1 U18802 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19726) );
  AOI21_X1 U18803 ( .B1(n19777), .B2(n19809), .A(n19726), .ZN(n15726) );
  NAND2_X1 U18804 ( .A1(n15728), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n15725) );
  OAI211_X1 U18805 ( .C1(n19752), .C2(n15726), .A(n15725), .B(n20089), .ZN(
        n15727) );
  NOR2_X1 U18806 ( .A1(n19523), .A2(n19781), .ZN(n19772) );
  INV_X1 U18807 ( .A(n19772), .ZN(n15732) );
  AOI21_X1 U18808 ( .B1(n15727), .B2(n15732), .A(n19639), .ZN(n19758) );
  INV_X1 U18809 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15736) );
  INV_X1 U18810 ( .A(n15728), .ZN(n15729) );
  OAI21_X1 U18811 ( .B1(n15729), .B2(n19772), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15730) );
  OAI21_X1 U18812 ( .B1(n19781), .B2(n19526), .A(n15730), .ZN(n19773) );
  INV_X1 U18813 ( .A(n19912), .ZN(n15733) );
  AOI22_X1 U18814 ( .A1(n19769), .A2(n19921), .B1(n19801), .B2(n19873), .ZN(
        n15731) );
  OAI21_X1 U18815 ( .B1(n15733), .B2(n15732), .A(n15731), .ZN(n15734) );
  AOI21_X1 U18816 ( .B1(n19773), .B2(n19913), .A(n15734), .ZN(n15735) );
  OAI21_X1 U18817 ( .B1(n19758), .B2(n15736), .A(n15735), .ZN(P2_U3128) );
  NAND3_X1 U18818 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20088), .ZN(n19831) );
  NOR2_X1 U18819 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19831), .ZN(
        n19821) );
  AOI21_X1 U18820 ( .B1(n12535), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n15742) );
  NOR2_X1 U18821 ( .A1(n15738), .A2(n15737), .ZN(n19586) );
  AOI21_X1 U18822 ( .B1(n19827), .B2(n19862), .A(n19726), .ZN(n15739) );
  AOI21_X1 U18823 ( .B1(n19586), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n15739), .ZN(n15740) );
  INV_X1 U18824 ( .A(n15740), .ZN(n15741) );
  OAI211_X1 U18825 ( .C1(n19821), .C2(n15742), .A(n15741), .B(n19919), .ZN(
        n19824) );
  INV_X1 U18826 ( .A(n19824), .ZN(n15755) );
  AOI22_X1 U18827 ( .A1(n19816), .A2(n19921), .B1(n19823), .B2(n19873), .ZN(
        n15749) );
  INV_X1 U18828 ( .A(n15743), .ZN(n15747) );
  INV_X1 U18829 ( .A(n19586), .ZN(n15746) );
  INV_X1 U18830 ( .A(n12535), .ZN(n15744) );
  OAI21_X1 U18831 ( .B1(n15744), .B2(n19821), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15745) );
  OAI21_X1 U18832 ( .B1(n15747), .B2(n15746), .A(n15745), .ZN(n19822) );
  AOI22_X1 U18833 ( .A1(n19822), .A2(n19913), .B1(n19912), .B2(n19821), .ZN(
        n15748) );
  OAI211_X1 U18834 ( .C1(n15755), .C2(n15750), .A(n15749), .B(n15748), .ZN(
        P2_U3144) );
  INV_X1 U18835 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n18485) );
  AOI22_X1 U18836 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19480), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19479), .ZN(n19930) );
  AOI22_X1 U18837 ( .A1(n19816), .A2(n19927), .B1(n19823), .B2(n19883), .ZN(
        n15753) );
  NOR2_X2 U18838 ( .A1(n19381), .A2(n19639), .ZN(n19926) );
  NOR2_X2 U18839 ( .A1(n15751), .A2(n19468), .ZN(n19925) );
  AOI22_X1 U18840 ( .A1(n19822), .A2(n19926), .B1(n19821), .B2(n19925), .ZN(
        n15752) );
  OAI211_X1 U18841 ( .C1(n15755), .C2(n15754), .A(n15753), .B(n15752), .ZN(
        P2_U3145) );
  AOI22_X1 U18842 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9656), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15760) );
  AOI22_X1 U18843 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15759) );
  AOI22_X1 U18844 ( .A1(n15864), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15758) );
  AOI22_X1 U18845 ( .A1(n17380), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15757) );
  NAND4_X1 U18846 ( .A1(n15760), .A2(n15759), .A3(n15758), .A4(n15757), .ZN(
        n15766) );
  AOI22_X1 U18847 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15764) );
  AOI22_X1 U18848 ( .A1(n17432), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15763) );
  AOI22_X1 U18849 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n15929), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15762) );
  AOI22_X1 U18850 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9658), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15761) );
  NAND4_X1 U18851 ( .A1(n15764), .A2(n15763), .A3(n15762), .A4(n15761), .ZN(
        n15765) );
  NOR2_X1 U18852 ( .A1(n15766), .A2(n15765), .ZN(n17240) );
  AOI22_X1 U18853 ( .A1(n17432), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15770) );
  AOI22_X1 U18854 ( .A1(n9656), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15769) );
  AOI22_X1 U18855 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n15929), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15768) );
  AOI22_X1 U18856 ( .A1(n15864), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17380), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15767) );
  NAND4_X1 U18857 ( .A1(n15770), .A2(n15769), .A3(n15768), .A4(n15767), .ZN(
        n15776) );
  AOI22_X1 U18858 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15774) );
  AOI22_X1 U18859 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17407), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15773) );
  AOI22_X1 U18860 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15772) );
  AOI22_X1 U18861 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9658), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15771) );
  NAND4_X1 U18862 ( .A1(n15774), .A2(n15773), .A3(n15772), .A4(n15771), .ZN(
        n15775) );
  NOR2_X1 U18863 ( .A1(n15776), .A2(n15775), .ZN(n17253) );
  AOI22_X1 U18864 ( .A1(n17380), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15780) );
  AOI22_X1 U18865 ( .A1(n17407), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15779) );
  AOI22_X1 U18866 ( .A1(n15864), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15929), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15778) );
  AOI22_X1 U18867 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9656), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15777) );
  NAND4_X1 U18868 ( .A1(n15780), .A2(n15779), .A3(n15778), .A4(n15777), .ZN(
        n15786) );
  AOI22_X1 U18869 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15784) );
  AOI22_X1 U18870 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15783) );
  AOI22_X1 U18871 ( .A1(n17432), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15782) );
  AOI22_X1 U18872 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9658), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15781) );
  NAND4_X1 U18873 ( .A1(n15784), .A2(n15783), .A3(n15782), .A4(n15781), .ZN(
        n15785) );
  NOR2_X1 U18874 ( .A1(n15786), .A2(n15785), .ZN(n17263) );
  AOI22_X1 U18875 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n15929), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15790) );
  AOI22_X1 U18876 ( .A1(n9656), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15789) );
  AOI22_X1 U18877 ( .A1(n17380), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17432), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15788) );
  AOI22_X1 U18878 ( .A1(n15864), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15787) );
  NAND4_X1 U18879 ( .A1(n15790), .A2(n15789), .A3(n15788), .A4(n15787), .ZN(
        n15796) );
  AOI22_X1 U18880 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15794) );
  AOI22_X1 U18881 ( .A1(n17407), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15793) );
  AOI22_X1 U18882 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15792) );
  AOI22_X1 U18883 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9658), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15791) );
  NAND4_X1 U18884 ( .A1(n15794), .A2(n15793), .A3(n15792), .A4(n15791), .ZN(
        n15795) );
  NOR2_X1 U18885 ( .A1(n15796), .A2(n15795), .ZN(n17264) );
  NOR2_X1 U18886 ( .A1(n17263), .A2(n17264), .ZN(n17262) );
  AOI22_X1 U18887 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15807) );
  INV_X1 U18888 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15799) );
  AOI22_X1 U18889 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n15929), .ZN(n15798) );
  AOI22_X1 U18890 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n9655), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15797) );
  OAI211_X1 U18891 ( .C1(n15799), .C2(n13974), .A(n15798), .B(n15797), .ZN(
        n15805) );
  AOI22_X1 U18892 ( .A1(n15864), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n17432), .ZN(n15803) );
  AOI22_X1 U18893 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17407), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n15802) );
  AOI22_X1 U18894 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n9656), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n17212), .ZN(n15801) );
  AOI22_X1 U18895 ( .A1(n17380), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17447), .ZN(n15800) );
  NAND4_X1 U18896 ( .A1(n15803), .A2(n15802), .A3(n15801), .A4(n15800), .ZN(
        n15804) );
  AOI211_X1 U18897 ( .C1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .C2(n9658), .A(
        n15805), .B(n15804), .ZN(n15806) );
  NAND2_X1 U18898 ( .A1(n15807), .A2(n15806), .ZN(n17258) );
  NAND2_X1 U18899 ( .A1(n17262), .A2(n17258), .ZN(n17257) );
  NOR2_X1 U18900 ( .A1(n17253), .A2(n17257), .ZN(n17252) );
  AOI22_X1 U18901 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15818) );
  INV_X1 U18902 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15810) );
  AOI22_X1 U18903 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17380), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15809) );
  AOI22_X1 U18904 ( .A1(n17407), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15929), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15808) );
  OAI211_X1 U18905 ( .C1(n13974), .C2(n15810), .A(n15809), .B(n15808), .ZN(
        n15816) );
  AOI22_X1 U18906 ( .A1(n17432), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15814) );
  AOI22_X1 U18907 ( .A1(n9656), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(n9655), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15813) );
  AOI22_X1 U18908 ( .A1(n15864), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15812) );
  AOI22_X1 U18909 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15811) );
  NAND4_X1 U18910 ( .A1(n15814), .A2(n15813), .A3(n15812), .A4(n15811), .ZN(
        n15815) );
  AOI211_X1 U18911 ( .C1(n9658), .C2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n15816), .B(n15815), .ZN(n15817) );
  NAND2_X1 U18912 ( .A1(n15818), .A2(n15817), .ZN(n17246) );
  NAND2_X1 U18913 ( .A1(n17252), .A2(n17246), .ZN(n17245) );
  NOR2_X1 U18914 ( .A1(n17240), .A2(n17245), .ZN(n17239) );
  AOI22_X1 U18915 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15828) );
  INV_X1 U18916 ( .A(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15838) );
  AOI22_X1 U18917 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15820) );
  AOI22_X1 U18918 ( .A1(n15864), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17432), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15819) );
  OAI211_X1 U18919 ( .C1(n13974), .C2(n15838), .A(n15820), .B(n15819), .ZN(
        n15826) );
  AOI22_X1 U18920 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n15929), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15824) );
  AOI22_X1 U18921 ( .A1(n9656), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15823) );
  AOI22_X1 U18922 ( .A1(n17407), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15822) );
  AOI22_X1 U18923 ( .A1(n17380), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15821) );
  NAND4_X1 U18924 ( .A1(n15824), .A2(n15823), .A3(n15822), .A4(n15821), .ZN(
        n15825) );
  AOI211_X1 U18925 ( .C1(n9658), .C2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A(
        n15826), .B(n15825), .ZN(n15827) );
  NAND2_X1 U18926 ( .A1(n15828), .A2(n15827), .ZN(n15829) );
  NAND2_X1 U18927 ( .A1(n17239), .A2(n15829), .ZN(n17234) );
  OAI21_X1 U18928 ( .B1(n17239), .B2(n15829), .A(n17234), .ZN(n17525) );
  NOR2_X1 U18929 ( .A1(n15877), .A2(n17489), .ZN(n15830) );
  AND2_X1 U18930 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n17232) );
  NAND2_X1 U18931 ( .A1(n18512), .A2(n17496), .ZN(n17502) );
  INV_X1 U18932 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n17199) );
  INV_X1 U18933 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16953) );
  INV_X1 U18934 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17345) );
  NAND2_X1 U18935 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17177) );
  INV_X1 U18936 ( .A(n17177), .ZN(n17490) );
  NAND2_X1 U18937 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n17490), .ZN(n17482) );
  INV_X1 U18938 ( .A(n17482), .ZN(n15832) );
  NAND3_X1 U18939 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n15832), .ZN(n17473) );
  INV_X1 U18940 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17469) );
  INV_X1 U18941 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17474) );
  NOR3_X1 U18942 ( .A1(n17102), .A2(n17469), .A3(n17474), .ZN(n17444) );
  NAND3_X1 U18943 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(P3_EBX_REG_8__SCAN_IN), 
        .A3(n17444), .ZN(n17427) );
  NAND4_X1 U18944 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .A3(P3_EBX_REG_11__SCAN_IN), .A4(P3_EBX_REG_10__SCAN_IN), .ZN(n15833)
         );
  NOR3_X1 U18945 ( .A1(n17473), .A2(n17427), .A3(n15833), .ZN(n15834) );
  NAND4_X1 U18946 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_15__SCAN_IN), 
        .A3(P3_EBX_REG_14__SCAN_IN), .A4(n15834), .ZN(n17346) );
  NOR3_X1 U18947 ( .A1(n17345), .A2(n17499), .A3(n17346), .ZN(n17320) );
  NAND2_X1 U18948 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17320), .ZN(n17306) );
  NAND2_X1 U18949 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17319), .ZN(n17290) );
  NOR2_X1 U18950 ( .A1(n17489), .A2(n17290), .ZN(n17292) );
  NAND2_X1 U18951 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17292), .ZN(n17279) );
  AND4_X1 U18952 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(P3_EBX_REG_24__SCAN_IN), .A4(P3_EBX_REG_23__SCAN_IN), .ZN(n17201)
         );
  NOR2_X1 U18953 ( .A1(n17500), .A2(n17241), .ZN(n17249) );
  INV_X1 U18954 ( .A(n17249), .ZN(n17243) );
  OAI21_X1 U18955 ( .B1(n17232), .B2(n17502), .A(n17243), .ZN(n17236) );
  INV_X1 U18956 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17244) );
  NOR2_X1 U18957 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17244), .ZN(n15835) );
  AOI22_X1 U18958 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17236), .B1(n17241), 
        .B2(n15835), .ZN(n15836) );
  OAI21_X1 U18959 ( .B1(n17525), .B2(n17494), .A(n15836), .ZN(P3_U2675) );
  AOI22_X1 U18960 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13971), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15848) );
  AOI22_X1 U18961 ( .A1(n15864), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17380), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15847) );
  AOI22_X1 U18962 ( .A1(n9656), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(n9655), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15837) );
  OAI21_X1 U18963 ( .B1(n15839), .B2(n15838), .A(n15837), .ZN(n15845) );
  AOI22_X1 U18964 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15843) );
  AOI22_X1 U18965 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15929), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15842) );
  AOI22_X1 U18966 ( .A1(n17432), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15841) );
  AOI22_X1 U18967 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9658), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15840) );
  NAND4_X1 U18968 ( .A1(n15843), .A2(n15842), .A3(n15841), .A4(n15840), .ZN(
        n15844) );
  AOI211_X1 U18969 ( .C1(n17334), .C2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n15845), .B(n15844), .ZN(n15846) );
  NAND3_X1 U18970 ( .A1(n15848), .A2(n15847), .A3(n15846), .ZN(n17601) );
  INV_X1 U18971 ( .A(n17601), .ZN(n15851) );
  INV_X1 U18972 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n17038) );
  INV_X1 U18973 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17431) );
  NOR3_X1 U18974 ( .A1(n17431), .A2(n17427), .A3(n17468), .ZN(n17415) );
  NAND2_X1 U18975 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n17415), .ZN(n17390) );
  NOR2_X1 U18976 ( .A1(n17038), .A2(n17390), .ZN(n15849) );
  NAND2_X1 U18977 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n15849), .ZN(n17372) );
  OAI21_X1 U18978 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n15849), .A(n17372), .ZN(
        n15850) );
  AOI22_X1 U18979 ( .A1(n17500), .A2(n15851), .B1(n15850), .B2(n17494), .ZN(
        P3_U2690) );
  NAND2_X1 U18980 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18647) );
  AOI221_X1 U18981 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18647), .C1(n15853), 
        .C2(n18647), .A(n15852), .ZN(n18474) );
  NOR2_X1 U18982 ( .A1(n15854), .A2(n18959), .ZN(n15855) );
  OAI21_X1 U18983 ( .B1(n15855), .B2(n18535), .A(n18475), .ZN(n18472) );
  AOI22_X1 U18984 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18474), .B1(
        n18472), .B2(n18964), .ZN(P3_U2865) );
  NOR4_X1 U18985 ( .A1(n12340), .A2(n15856), .A3(n20122), .A4(n20065), .ZN(
        n15857) );
  NAND2_X1 U18986 ( .A1(n20061), .A2(n15857), .ZN(n15858) );
  OAI21_X1 U18987 ( .B1(n20061), .B2(n15859), .A(n15858), .ZN(P2_U3595) );
  AOI22_X1 U18988 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15872) );
  INV_X1 U18989 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15863) );
  AOI22_X1 U18990 ( .A1(n17380), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15862) );
  AOI22_X1 U18991 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9656), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15861) );
  OAI211_X1 U18992 ( .C1(n13974), .C2(n15863), .A(n15862), .B(n15861), .ZN(
        n15870) );
  AOI22_X1 U18993 ( .A1(n15864), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15868) );
  AOI22_X1 U18994 ( .A1(n17432), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15867) );
  AOI22_X1 U18995 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15929), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15866) );
  AOI22_X1 U18996 ( .A1(n17407), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15865) );
  NAND4_X1 U18997 ( .A1(n15868), .A2(n15867), .A3(n15866), .A4(n15865), .ZN(
        n15869) );
  AOI211_X1 U18998 ( .C1(n9658), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n15870), .B(n15869), .ZN(n15871) );
  NAND2_X1 U18999 ( .A1(n18489), .A2(n16806), .ZN(n15884) );
  NOR2_X1 U19000 ( .A1(n18506), .A2(n15884), .ZN(n15882) );
  NAND2_X1 U19001 ( .A1(n15882), .A2(n15873), .ZN(n16668) );
  INV_X1 U19002 ( .A(n16668), .ZN(n18919) );
  INV_X1 U19003 ( .A(n15874), .ZN(n15875) );
  AOI21_X1 U19004 ( .B1(n15876), .B2(n15875), .A(n18917), .ZN(n16607) );
  OAI211_X1 U19005 ( .C1(n15878), .C2(n15877), .A(n18489), .B(n18922), .ZN(
        n15879) );
  INV_X1 U19006 ( .A(n15879), .ZN(n15881) );
  AOI21_X1 U19007 ( .B1(n19136), .B2(n15883), .A(n16803), .ZN(n15885) );
  INV_X1 U19008 ( .A(n19137), .ZN(n19002) );
  AOI21_X1 U19009 ( .B1(n15885), .B2(n15884), .A(n19002), .ZN(n16785) );
  INV_X1 U19010 ( .A(n15886), .ZN(n15887) );
  NAND3_X1 U19011 ( .A1(n16780), .A2(n16785), .A3(n15887), .ZN(n15888) );
  NAND2_X1 U19012 ( .A1(n18919), .A2(n18391), .ZN(n18467) );
  NOR2_X1 U19013 ( .A1(n16666), .A2(n18467), .ZN(n18384) );
  NAND2_X1 U19014 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16027) );
  NAND2_X1 U19015 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18158) );
  NOR2_X1 U19016 ( .A1(n18272), .A2(n17926), .ZN(n18247) );
  NAND2_X1 U19017 ( .A1(n18247), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18217) );
  INV_X1 U19018 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17880) );
  NOR2_X1 U19019 ( .A1(n18238), .A2(n17880), .ZN(n18219) );
  NAND2_X1 U19020 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18219), .ZN(
        n18205) );
  NOR2_X1 U19021 ( .A1(n18217), .A2(n18205), .ZN(n18151) );
  NAND2_X1 U19022 ( .A1(n18151), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18197) );
  NOR2_X1 U19023 ( .A1(n18190), .A2(n18197), .ZN(n17822) );
  INV_X1 U19024 ( .A(n17822), .ZN(n17832) );
  INV_X1 U19025 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17836) );
  NOR2_X1 U19026 ( .A1(n17832), .A2(n17836), .ZN(n18174) );
  INV_X1 U19027 ( .A(n18174), .ZN(n18172) );
  INV_X1 U19028 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18300) );
  NAND2_X1 U19029 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18334) );
  NOR2_X1 U19030 ( .A1(n18334), .A2(n17993), .ZN(n18322) );
  NAND2_X1 U19031 ( .A1(n18322), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18291) );
  INV_X1 U19032 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17983) );
  NOR2_X1 U19033 ( .A1(n18291), .A2(n17983), .ZN(n18297) );
  INV_X1 U19034 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18373) );
  AOI22_X1 U19035 ( .A1(n9656), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15929), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15893) );
  AOI22_X1 U19036 ( .A1(n17380), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15892) );
  AOI22_X1 U19037 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15891) );
  AOI22_X1 U19038 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17407), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15890) );
  NAND4_X1 U19039 ( .A1(n15893), .A2(n15892), .A3(n15891), .A4(n15890), .ZN(
        n15900) );
  AOI22_X1 U19040 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15898) );
  AOI22_X1 U19041 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15897) );
  AOI22_X1 U19042 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17432), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15896) );
  AOI22_X1 U19043 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9658), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15895) );
  NAND4_X1 U19044 ( .A1(n15898), .A2(n15897), .A3(n15896), .A4(n15895), .ZN(
        n15899) );
  AOI22_X1 U19045 ( .A1(n17432), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15904) );
  AOI22_X1 U19046 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15903) );
  AOI22_X1 U19047 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17380), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15902) );
  AOI22_X1 U19048 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17407), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15901) );
  NAND4_X1 U19049 ( .A1(n15904), .A2(n15903), .A3(n15902), .A4(n15901), .ZN(
        n15910) );
  AOI22_X1 U19050 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15908) );
  AOI22_X1 U19051 ( .A1(n9656), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15907) );
  AOI22_X1 U19052 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n15929), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15906) );
  AOI22_X1 U19053 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9658), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15905) );
  NAND4_X1 U19054 ( .A1(n15908), .A2(n15907), .A3(n15906), .A4(n15905), .ZN(
        n15909) );
  AOI22_X1 U19055 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n15911), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n17212), .ZN(n15917) );
  AOI22_X1 U19056 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n15912), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17447), .ZN(n15916) );
  AOI22_X1 U19057 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15915) );
  AOI22_X1 U19058 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n17395), .B1(
        n15913), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15914) );
  INV_X1 U19059 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17495) );
  AOI22_X1 U19060 ( .A1(n15940), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n15929), .ZN(n15918) );
  OAI21_X1 U19061 ( .B1(n17150), .B2(n17495), .A(n15918), .ZN(n15924) );
  AOI22_X1 U19062 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n9656), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17456), .ZN(n15919) );
  AOI22_X1 U19063 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n13948), .ZN(n15921) );
  AOI22_X1 U19064 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15936) );
  INV_X1 U19065 ( .A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15928) );
  AOI22_X1 U19066 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15927) );
  AOI22_X1 U19067 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9656), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15926) );
  OAI211_X1 U19068 ( .C1(n13974), .C2(n15928), .A(n15927), .B(n15926), .ZN(
        n15935) );
  AOI22_X1 U19069 ( .A1(n13964), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15933) );
  AOI22_X1 U19070 ( .A1(n17407), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15932) );
  AOI22_X1 U19071 ( .A1(n15940), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15931) );
  NAND4_X1 U19072 ( .A1(n15933), .A2(n15932), .A3(n15931), .A4(n15930), .ZN(
        n15934) );
  NAND2_X1 U19073 ( .A1(n17654), .A2(n15988), .ZN(n15969) );
  AOI22_X1 U19074 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15948) );
  INV_X1 U19075 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15939) );
  AOI22_X1 U19076 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15938) );
  AOI22_X1 U19077 ( .A1(n9656), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17432), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15937) );
  OAI211_X1 U19078 ( .C1(n13974), .C2(n15939), .A(n15938), .B(n15937), .ZN(
        n15946) );
  AOI22_X1 U19079 ( .A1(n17380), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15943) );
  AOI22_X1 U19080 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15942) );
  AOI22_X1 U19081 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17407), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15941) );
  NAND4_X1 U19082 ( .A1(n15944), .A2(n15943), .A3(n15942), .A4(n15941), .ZN(
        n15945) );
  AOI211_X1 U19083 ( .C1(n9658), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n15946), .B(n15945), .ZN(n15947) );
  NAND2_X1 U19084 ( .A1(n15948), .A2(n15947), .ZN(n16003) );
  NAND2_X1 U19085 ( .A1(n15973), .A2(n16003), .ZN(n15976) );
  AOI22_X1 U19086 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n15959) );
  INV_X1 U19087 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15951) );
  AOI22_X1 U19088 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n15950) );
  AOI22_X1 U19089 ( .A1(n17380), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n15929), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15949) );
  OAI211_X1 U19090 ( .C1(n13974), .C2(n15951), .A(n15950), .B(n15949), .ZN(
        n15957) );
  AOI22_X1 U19091 ( .A1(n9656), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n15955) );
  AOI22_X1 U19092 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n15954) );
  AOI22_X1 U19093 ( .A1(n17432), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n15953) );
  AOI22_X1 U19094 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17407), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15952) );
  NAND4_X1 U19095 ( .A1(n15955), .A2(n15954), .A3(n15953), .A4(n15952), .ZN(
        n15956) );
  AOI211_X1 U19096 ( .C1(n9658), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n15957), .B(n15956), .ZN(n15958) );
  NAND2_X1 U19097 ( .A1(n15959), .A2(n15958), .ZN(n16010) );
  OAI21_X1 U19098 ( .B1(n15960), .B2(n16666), .A(n18050), .ZN(n15980) );
  INV_X1 U19099 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19097) );
  NOR2_X1 U19100 ( .A1(n17654), .A2(n19097), .ZN(n15966) );
  XNOR2_X1 U19101 ( .A(n15995), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18134) );
  AOI22_X1 U19102 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15965) );
  INV_X1 U19103 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15962) );
  AOI22_X1 U19104 ( .A1(n13964), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15961) );
  AOI22_X1 U19105 ( .A1(n15940), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13948), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15964) );
  AOI22_X1 U19106 ( .A1(n17456), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15963) );
  NAND2_X1 U19107 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18142), .ZN(
        n18141) );
  NOR2_X1 U19108 ( .A1(n18134), .A2(n18141), .ZN(n18133) );
  NOR2_X1 U19109 ( .A1(n15966), .A2(n18133), .ZN(n18122) );
  NOR2_X1 U19110 ( .A1(n18122), .A2(n18121), .ZN(n18120) );
  NOR2_X1 U19111 ( .A1(n18436), .A2(n15967), .ZN(n15968) );
  INV_X1 U19112 ( .A(n17642), .ZN(n15989) );
  XOR2_X1 U19113 ( .A(n15989), .B(n15969), .Z(n15970) );
  XNOR2_X1 U19114 ( .A(n15971), .B(n15970), .ZN(n18114) );
  NOR2_X1 U19115 ( .A1(n18430), .A2(n18114), .ZN(n18113) );
  NOR2_X1 U19116 ( .A1(n15971), .A2(n15970), .ZN(n15972) );
  INV_X1 U19117 ( .A(n16003), .ZN(n17639) );
  XNOR2_X1 U19118 ( .A(n17639), .B(n15973), .ZN(n15974) );
  XNOR2_X1 U19119 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n15974), .ZN(
        n18099) );
  AND2_X1 U19120 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n15974), .ZN(
        n15975) );
  INV_X1 U19121 ( .A(n17635), .ZN(n15990) );
  XOR2_X1 U19122 ( .A(n15990), .B(n15976), .Z(n18085) );
  INV_X1 U19123 ( .A(n16010), .ZN(n17632) );
  XNOR2_X1 U19124 ( .A(n17632), .B(n15977), .ZN(n15978) );
  XNOR2_X1 U19125 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n15978), .ZN(
        n18073) );
  NAND2_X1 U19126 ( .A1(n18297), .A2(n18331), .ZN(n17970) );
  INV_X1 U19127 ( .A(n18154), .ZN(n16028) );
  NOR2_X1 U19128 ( .A1(n16027), .A2(n16028), .ZN(n16671) );
  NOR2_X1 U19129 ( .A1(n19136), .A2(n15984), .ZN(n15986) );
  AOI21_X1 U19130 ( .B1(n15986), .B2(n18915), .A(n15985), .ZN(n18933) );
  INV_X1 U19131 ( .A(n18463), .ZN(n18457) );
  NAND2_X1 U19132 ( .A1(n18142), .A2(n17654), .ZN(n15993) );
  NAND2_X1 U19133 ( .A1(n17647), .A2(n15993), .ZN(n15992) );
  NAND2_X1 U19134 ( .A1(n15992), .A2(n15989), .ZN(n16004) );
  NOR2_X1 U19135 ( .A1(n17639), .A2(n16004), .ZN(n15991) );
  NAND2_X1 U19136 ( .A1(n15991), .A2(n15990), .ZN(n16011) );
  NOR2_X1 U19137 ( .A1(n17632), .A2(n16011), .ZN(n16014) );
  NAND2_X1 U19138 ( .A1(n16014), .A2(n16666), .ZN(n16015) );
  XNOR2_X1 U19139 ( .A(n15991), .B(n17635), .ZN(n16008) );
  AND2_X1 U19140 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n16008), .ZN(
        n16009) );
  XOR2_X1 U19141 ( .A(n15992), .B(n17642), .Z(n16001) );
  NOR2_X1 U19142 ( .A1(n18430), .A2(n16001), .ZN(n16002) );
  NOR2_X1 U19143 ( .A1(n15994), .A2(n18436), .ZN(n16000) );
  INV_X1 U19144 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19112) );
  NOR2_X1 U19145 ( .A1(n15995), .A2(n19112), .ZN(n15998) );
  INV_X1 U19146 ( .A(n18142), .ZN(n15997) );
  NAND3_X1 U19147 ( .A1(n15997), .A2(n15995), .A3(n19112), .ZN(n15996) );
  OAI221_X1 U19148 ( .B1(n15998), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n15997), .C2(n15995), .A(n15996), .ZN(n18123) );
  NOR2_X1 U19149 ( .A1(n16000), .A2(n15999), .ZN(n18112) );
  XNOR2_X1 U19150 ( .A(n18430), .B(n16001), .ZN(n18111) );
  NOR2_X1 U19151 ( .A1(n18112), .A2(n18111), .ZN(n18110) );
  XOR2_X1 U19152 ( .A(n16004), .B(n16003), .Z(n16006) );
  NOR2_X1 U19153 ( .A1(n16005), .A2(n16006), .ZN(n16007) );
  INV_X1 U19154 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18097) );
  XNOR2_X1 U19155 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n16008), .ZN(
        n18088) );
  NOR2_X1 U19156 ( .A1(n18089), .A2(n18088), .ZN(n18087) );
  XOR2_X1 U19157 ( .A(n16011), .B(n16010), .Z(n16013) );
  INV_X1 U19158 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18374) );
  XNOR2_X1 U19159 ( .A(n16014), .B(n16666), .ZN(n16017) );
  NAND2_X1 U19160 ( .A1(n16016), .A2(n16017), .ZN(n18063) );
  NAND2_X1 U19161 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18063), .ZN(
        n16019) );
  NOR2_X1 U19162 ( .A1(n16015), .A2(n16019), .ZN(n16021) );
  INV_X1 U19163 ( .A(n16015), .ZN(n16020) );
  OR2_X1 U19164 ( .A1(n16017), .A2(n16016), .ZN(n18064) );
  OAI21_X1 U19165 ( .B1(n16020), .B2(n16019), .A(n18064), .ZN(n16018) );
  AOI21_X1 U19166 ( .B1(n16020), .B2(n16019), .A(n16018), .ZN(n18049) );
  NOR2_X2 U19167 ( .A1(n18049), .A2(n18380), .ZN(n18048) );
  INV_X1 U19168 ( .A(n18297), .ZN(n18292) );
  NAND2_X1 U19169 ( .A1(n17956), .A2(n18174), .ZN(n17818) );
  NAND3_X1 U19170 ( .A1(n18155), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16672) );
  NOR3_X1 U19171 ( .A1(n18190), .A2(n17836), .A3(n18158), .ZN(n16024) );
  INV_X1 U19172 ( .A(n16024), .ZN(n18160) );
  NOR2_X1 U19173 ( .A1(n18197), .A2(n18160), .ZN(n16026) );
  NAND2_X1 U19174 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n16026), .ZN(
        n16667) );
  INV_X1 U19175 ( .A(n16667), .ZN(n16022) );
  NAND2_X1 U19176 ( .A1(n18297), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n18274) );
  NAND3_X1 U19177 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18390) );
  INV_X1 U19178 ( .A(n18390), .ZN(n18241) );
  OAI21_X1 U19179 ( .B1(n19112), .B2(n19097), .A(n18436), .ZN(n18431) );
  NAND2_X1 U19180 ( .A1(n18241), .A2(n18431), .ZN(n18368) );
  NAND2_X1 U19181 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18367) );
  OR2_X1 U19182 ( .A1(n18380), .A2(n18367), .ZN(n18275) );
  NOR2_X1 U19183 ( .A1(n18368), .A2(n18275), .ZN(n18262) );
  NAND2_X1 U19184 ( .A1(n18243), .A2(n18262), .ZN(n18246) );
  NOR2_X1 U19185 ( .A1(n18436), .A2(n19097), .ZN(n18416) );
  NAND2_X1 U19186 ( .A1(n18241), .A2(n18416), .ZN(n18370) );
  OR2_X1 U19187 ( .A1(n18275), .A2(n18370), .ZN(n18311) );
  NOR2_X1 U19188 ( .A1(n9856), .A2(n18311), .ZN(n18206) );
  INV_X1 U19189 ( .A(n18206), .ZN(n18245) );
  INV_X1 U19190 ( .A(n18953), .ZN(n18312) );
  AOI21_X1 U19191 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18951), .A(
        n18312), .ZN(n18240) );
  OAI22_X1 U19192 ( .A1(n18949), .A2(n18246), .B1(n18245), .B2(n18240), .ZN(
        n18173) );
  NAND4_X1 U19193 ( .A1(n18391), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n16022), .A4(n18173), .ZN(n16655) );
  OAI21_X1 U19194 ( .B1(n18457), .B2(n16672), .A(n16655), .ZN(n16023) );
  AOI21_X1 U19195 ( .B1(n18384), .B2(n16671), .A(n16023), .ZN(n16103) );
  NOR2_X1 U19196 ( .A1(n19112), .A2(n18311), .ZN(n18336) );
  NAND2_X1 U19197 ( .A1(n18243), .A2(n18336), .ZN(n18261) );
  OAI21_X1 U19198 ( .B1(n18197), .B2(n18246), .A(n18931), .ZN(n18191) );
  OAI21_X1 U19199 ( .B1(n16024), .B2(n18949), .A(n18191), .ZN(n18157) );
  AOI221_X1 U19200 ( .B1(n18261), .B2(n18951), .C1(n16667), .C2(n18951), .A(
        n18157), .ZN(n16025) );
  OAI221_X1 U19201 ( .B1(n18953), .B2(n16026), .C1(n18953), .C2(n18206), .A(
        n16025), .ZN(n16105) );
  AOI21_X1 U19202 ( .B1(n18265), .B2(n10013), .A(n16105), .ZN(n16670) );
  NOR2_X1 U19203 ( .A1(n18267), .A2(n18459), .ZN(n18376) );
  INV_X1 U19204 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17776) );
  INV_X1 U19205 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18986) );
  INV_X1 U19206 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16651) );
  NOR2_X1 U19207 ( .A1(n16027), .A2(n16651), .ZN(n16635) );
  INV_X1 U19208 ( .A(n16635), .ZN(n16104) );
  NOR2_X1 U19209 ( .A1(n16104), .A2(n16028), .ZN(n16628) );
  INV_X1 U19210 ( .A(n18384), .ZN(n16030) );
  NAND2_X1 U19211 ( .A1(n18155), .A2(n16635), .ZN(n16629) );
  NAND2_X1 U19212 ( .A1(n18463), .A2(n16629), .ZN(n16029) );
  OAI21_X1 U19213 ( .B1(n16628), .B2(n16030), .A(n16029), .ZN(n16107) );
  AOI211_X1 U19214 ( .C1(n18376), .C2(n17776), .A(n18454), .B(n16107), .ZN(
        n16031) );
  OAI21_X1 U19215 ( .B1(n16670), .B2(n18459), .A(n16031), .ZN(n16046) );
  INV_X1 U19216 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18171) );
  INV_X1 U19217 ( .A(n16033), .ZN(n18017) );
  INV_X1 U19218 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18365) );
  INV_X1 U19219 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18338) );
  NAND2_X1 U19220 ( .A1(n18365), .A2(n18338), .ZN(n18027) );
  NOR2_X1 U19221 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18027), .ZN(
        n17950) );
  NOR2_X1 U19222 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17951) );
  NAND4_X1 U19223 ( .A1(n17950), .A2(n17951), .A3(n17983), .A4(n17957), .ZN(
        n16032) );
  NAND2_X1 U19224 ( .A1(n17927), .A2(n17926), .ZN(n17925) );
  NAND2_X1 U19225 ( .A1(n16035), .A2(n16034), .ZN(n17931) );
  NAND2_X1 U19226 ( .A1(n17931), .A2(n17822), .ZN(n16037) );
  NAND2_X1 U19227 ( .A1(n17914), .A2(n18238), .ZN(n16036) );
  NOR2_X1 U19228 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n16036), .ZN(
        n17875) );
  INV_X1 U19229 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17867) );
  NAND2_X1 U19230 ( .A1(n17875), .A2(n17867), .ZN(n17859) );
  NAND2_X1 U19231 ( .A1(n18247), .A2(n17931), .ZN(n17874) );
  INV_X1 U19232 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17907) );
  NOR2_X1 U19233 ( .A1(n17907), .A2(n18205), .ZN(n17860) );
  AND2_X1 U19234 ( .A1(n17860), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16039) );
  OR2_X1 U19235 ( .A1(n17952), .A2(n17830), .ZN(n17809) );
  OAI221_X1 U19236 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n18050), 
        .C1(n18171), .C2(n17810), .A(n17809), .ZN(n17799) );
  NOR2_X1 U19237 ( .A1(n17810), .A2(n18050), .ZN(n16041) );
  AND2_X1 U19238 ( .A1(n17952), .A2(n18158), .ZN(n16040) );
  NOR2_X1 U19239 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18050), .ZN(
        n16665) );
  AOI21_X1 U19240 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n18050), .A(
        n16665), .ZN(n17780) );
  AOI22_X1 U19241 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16046), .B1(
        n18362), .B2(n16645), .ZN(n16047) );
  NAND2_X1 U19242 ( .A1(n9652), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16642) );
  OAI211_X1 U19243 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16103), .A(
        n16047), .B(n16642), .ZN(P3_U2833) );
  NAND2_X1 U19244 ( .A1(n16048), .A2(n19314), .ZN(n16052) );
  OAI22_X1 U19245 ( .A1(n10752), .A2(n19334), .B1(n20024), .B2(n19301), .ZN(
        n16050) );
  AND2_X1 U19246 ( .A1(n19326), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n16049) );
  NOR2_X1 U19247 ( .A1(n16050), .A2(n16049), .ZN(n16051) );
  OAI211_X1 U19248 ( .C1(n19304), .C2(n16053), .A(n16052), .B(n16051), .ZN(
        n16054) );
  INV_X1 U19249 ( .A(n16054), .ZN(n16059) );
  OAI211_X1 U19250 ( .C1(n16057), .C2(n16056), .A(n19315), .B(n16055), .ZN(
        n16058) );
  OAI211_X1 U19251 ( .C1(n19320), .C2(n16060), .A(n16059), .B(n16058), .ZN(
        P2_U2833) );
  AND2_X1 U19252 ( .A1(n16062), .A2(n16061), .ZN(n16074) );
  NAND2_X1 U19253 ( .A1(n16062), .A2(n16063), .ZN(n16072) );
  NOR3_X1 U19254 ( .A1(n16065), .A2(n16064), .A3(n20643), .ZN(n16066) );
  NAND2_X1 U19255 ( .A1(n16066), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n16070) );
  OAI22_X1 U19256 ( .A1(n16068), .A2(n16067), .B1(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n16066), .ZN(n16069) );
  NAND2_X1 U19257 ( .A1(n16070), .A2(n16069), .ZN(n16071) );
  AOI222_X1 U19258 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n16072), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16071), .C1(n16072), 
        .C2(n16071), .ZN(n16073) );
  AOI222_X1 U19259 ( .A1(n20528), .A2(n16074), .B1(n20528), .B2(n16073), .C1(
        n16074), .C2(n16073), .ZN(n16075) );
  OR2_X1 U19260 ( .A1(n16075), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n16085) );
  AND2_X1 U19261 ( .A1(n21039), .A2(n21037), .ZN(n16078) );
  OAI211_X1 U19262 ( .C1(n16079), .C2(n16078), .A(n16077), .B(n16076), .ZN(
        n16080) );
  NOR2_X1 U19263 ( .A1(n16081), .A2(n16080), .ZN(n16082) );
  AND2_X1 U19264 ( .A1(n16083), .A2(n16082), .ZN(n16084) );
  INV_X1 U19265 ( .A(n16101), .ZN(n16092) );
  NAND2_X1 U19266 ( .A1(n16087), .A2(n16086), .ZN(n16090) );
  NOR3_X1 U19267 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20753), .A3(n20850), 
        .ZN(n16088) );
  OAI22_X1 U19268 ( .A1(n16091), .A2(n16090), .B1(n16089), .B2(n16088), .ZN(
        n16343) );
  AOI221_X1 U19269 ( .B1(n20846), .B2(n16345), .C1(n16092), .C2(n16345), .A(
        n16343), .ZN(n16094) );
  NOR2_X1 U19270 ( .A1(n16094), .A2(n20846), .ZN(n20752) );
  OAI211_X1 U19271 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20850), .A(n20752), 
        .B(n16093), .ZN(n16344) );
  AOI21_X1 U19272 ( .B1(n16096), .B2(n16095), .A(n16094), .ZN(n16097) );
  OAI22_X1 U19273 ( .A1(n16098), .A2(n16344), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n16097), .ZN(n16099) );
  OAI21_X1 U19274 ( .B1(n16101), .B2(n16100), .A(n16099), .ZN(P1_U3161) );
  NAND2_X1 U19275 ( .A1(n16635), .A2(n16669), .ZN(n16610) );
  OAI21_X1 U19276 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16102), .A(
        n16613), .ZN(n16638) );
  AOI22_X1 U19277 ( .A1(n18391), .A2(n16105), .B1(n18376), .B2(n16104), .ZN(
        n16106) );
  NAND2_X1 U19278 ( .A1(n16106), .A2(n18460), .ZN(n16653) );
  NOR2_X1 U19279 ( .A1(n16653), .A2(n16107), .ZN(n16108) );
  MUX2_X1 U19280 ( .A(n10288), .B(n16108), .S(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Z(n16109) );
  NAND2_X1 U19281 ( .A1(n9652), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16630) );
  OAI211_X1 U19282 ( .C1(n18388), .C2(n16638), .A(n16109), .B(n16630), .ZN(
        P3_U2832) );
  INV_X1 U19283 ( .A(HOLD), .ZN(n21016) );
  NOR2_X1 U19284 ( .A1(n20755), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20130) );
  INV_X1 U19285 ( .A(n20130), .ZN(n20760) );
  INV_X1 U19286 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21021) );
  NOR2_X1 U19287 ( .A1(n20129), .A2(n21021), .ZN(n16111) );
  NAND2_X1 U19288 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n16110) );
  AOI22_X1 U19289 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20840), .B1(n16111), 
        .B2(n16110), .ZN(n16113) );
  OAI211_X1 U19290 ( .C1(n21016), .C2(n20760), .A(n16113), .B(n16112), .ZN(
        P1_U3195) );
  AND2_X1 U19291 ( .A1(n16114), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR3_X1 U19292 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n16117) );
  INV_X1 U19293 ( .A(n19159), .ZN(n16116) );
  NOR3_X1 U19294 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19974), .A3(n20114), 
        .ZN(n16598) );
  NOR4_X1 U19295 ( .A1(n16117), .A2(n16116), .A3(n16598), .A4(n16115), .ZN(
        P2_U3178) );
  INV_X1 U19296 ( .A(n20102), .ZN(n16118) );
  OAI221_X1 U19297 ( .B1(n16120), .B2(n16119), .C1(n16118), .C2(n16119), .A(
        n19639), .ZN(n20094) );
  NOR2_X1 U19298 ( .A1(n16121), .A2(n20094), .ZN(P2_U3047) );
  NOR3_X1 U19299 ( .A1(n16122), .A2(n17661), .A3(n16806), .ZN(n16123) );
  INV_X1 U19300 ( .A(n17653), .ZN(n16127) );
  NAND2_X1 U19301 ( .A1(n18512), .A2(n16127), .ZN(n17652) );
  NOR2_X1 U19302 ( .A1(n16125), .A2(n17653), .ZN(n17656) );
  AOI22_X1 U19303 ( .A1(n17656), .A2(BUF2_REG_0__SCAN_IN), .B1(n17655), .B2(
        n18142), .ZN(n16126) );
  OAI221_X1 U19304 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17652), .C1(n17733), 
        .C2(n16127), .A(n16126), .ZN(P3_U2735) );
  OAI21_X1 U19305 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(P1_REIP_REG_15__SCAN_IN), 
        .A(n16128), .ZN(n16137) );
  INV_X1 U19306 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16129) );
  NOR2_X1 U19307 ( .A1(n20177), .A2(n16129), .ZN(n16130) );
  AOI211_X1 U19308 ( .C1(n20175), .C2(P1_EBX_REG_16__SCAN_IN), .A(n20174), .B(
        n16130), .ZN(n16131) );
  OAI21_X1 U19309 ( .B1(n16164), .B2(n20189), .A(n16131), .ZN(n16132) );
  AOI21_X1 U19310 ( .B1(n16133), .B2(n20183), .A(n16132), .ZN(n16136) );
  OR2_X1 U19311 ( .A1(n16134), .A2(n20161), .ZN(n16152) );
  INV_X1 U19312 ( .A(n16152), .ZN(n16143) );
  AOI22_X1 U19313 ( .A1(n16161), .A2(n20151), .B1(n16143), .B2(
        P1_REIP_REG_16__SCAN_IN), .ZN(n16135) );
  OAI211_X1 U19314 ( .C1(n16146), .C2(n16137), .A(n16136), .B(n16135), .ZN(
        P1_U2824) );
  INV_X1 U19315 ( .A(n16138), .ZN(n16139) );
  AOI22_X1 U19316 ( .A1(n16139), .A2(n20183), .B1(n20175), .B2(
        P1_EBX_REG_15__SCAN_IN), .ZN(n16140) );
  OAI211_X1 U19317 ( .C1(n20177), .C2(n16141), .A(n16140), .B(n20191), .ZN(
        n16142) );
  AOI21_X1 U19318 ( .B1(n16165), .B2(n20197), .A(n16142), .ZN(n16145) );
  AOI22_X1 U19319 ( .A1(n16166), .A2(n20151), .B1(P1_REIP_REG_15__SCAN_IN), 
        .B2(n16143), .ZN(n16144) );
  OAI211_X1 U19320 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n16146), .A(n16145), 
        .B(n16144), .ZN(P1_U2825) );
  AOI21_X1 U19321 ( .B1(n16147), .B2(P1_REIP_REG_13__SCAN_IN), .A(
        P1_REIP_REG_14__SCAN_IN), .ZN(n16153) );
  OAI22_X1 U19322 ( .A1(n16258), .A2(n20193), .B1(n16148), .B2(n20192), .ZN(
        n16149) );
  AOI211_X1 U19323 ( .C1(n20196), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16156), .B(n16149), .ZN(n16151) );
  AOI22_X1 U19324 ( .A1(n16178), .A2(n20151), .B1(n20197), .B2(n16177), .ZN(
        n16150) );
  OAI211_X1 U19325 ( .C1(n16153), .C2(n16152), .A(n16151), .B(n16150), .ZN(
        P1_U2826) );
  AOI22_X1 U19326 ( .A1(n16275), .A2(n20183), .B1(n20175), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n16154) );
  OAI21_X1 U19327 ( .B1(n16193), .B2(n20189), .A(n16154), .ZN(n16155) );
  AOI211_X1 U19328 ( .C1(n20196), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n16156), .B(n16155), .ZN(n16158) );
  AOI22_X1 U19329 ( .A1(n16190), .A2(n20151), .B1(P1_REIP_REG_11__SCAN_IN), 
        .B2(n10269), .ZN(n16157) );
  OAI211_X1 U19330 ( .C1(P1_REIP_REG_11__SCAN_IN), .C2(n16159), .A(n16158), 
        .B(n16157), .ZN(P1_U2829) );
  AOI22_X1 U19331 ( .A1(n16194), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n16319), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n16163) );
  AOI22_X1 U19332 ( .A1(n16161), .A2(n16205), .B1(n11980), .B2(n16160), .ZN(
        n16162) );
  OAI211_X1 U19333 ( .C1(n16202), .C2(n16164), .A(n16163), .B(n16162), .ZN(
        P1_U2983) );
  AOI22_X1 U19334 ( .A1(n16194), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n16319), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16168) );
  AOI22_X1 U19335 ( .A1(n16166), .A2(n16205), .B1(n16204), .B2(n16165), .ZN(
        n16167) );
  OAI211_X1 U19336 ( .C1(n16169), .C2(n20135), .A(n16168), .B(n16167), .ZN(
        P1_U2984) );
  INV_X1 U19337 ( .A(n16170), .ZN(n16171) );
  OAI21_X1 U19338 ( .B1(n16172), .B2(n16171), .A(n11906), .ZN(n16176) );
  AOI22_X1 U19339 ( .A1(n16174), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n16266), .B2(n16173), .ZN(n16175) );
  XNOR2_X1 U19340 ( .A(n16176), .B(n16175), .ZN(n16261) );
  AOI22_X1 U19341 ( .A1(n16194), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n16319), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16180) );
  AOI22_X1 U19342 ( .A1(n16178), .A2(n16205), .B1(n16204), .B2(n16177), .ZN(
        n16179) );
  OAI211_X1 U19343 ( .C1(n16261), .C2(n20135), .A(n16180), .B(n16179), .ZN(
        P1_U2985) );
  AOI22_X1 U19344 ( .A1(n16194), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n16319), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16184) );
  AOI22_X1 U19345 ( .A1(n16182), .A2(n16205), .B1(n16204), .B2(n16181), .ZN(
        n16183) );
  OAI211_X1 U19346 ( .C1(n16185), .C2(n20135), .A(n16184), .B(n16183), .ZN(
        P1_U2987) );
  AOI22_X1 U19347 ( .A1(n16194), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n16319), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16192) );
  NOR3_X1 U19348 ( .A1(n16186), .A2(n16174), .A3(n14627), .ZN(n16188) );
  NOR2_X1 U19349 ( .A1(n16188), .A2(n16187), .ZN(n16189) );
  XOR2_X1 U19350 ( .A(n11911), .B(n16189), .Z(n16278) );
  AOI22_X1 U19351 ( .A1(n16278), .A2(n11980), .B1(n16205), .B2(n16190), .ZN(
        n16191) );
  OAI211_X1 U19352 ( .C1(n16202), .C2(n16193), .A(n16192), .B(n16191), .ZN(
        P1_U2988) );
  AOI22_X1 U19353 ( .A1(n16194), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n16319), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16201) );
  NAND2_X1 U19354 ( .A1(n16197), .A2(n16196), .ZN(n16198) );
  XNOR2_X1 U19355 ( .A(n16195), .B(n16198), .ZN(n16321) );
  AOI22_X1 U19356 ( .A1(n16205), .A2(n16199), .B1(n16321), .B2(n11980), .ZN(
        n16200) );
  OAI211_X1 U19357 ( .C1(n16202), .C2(n20163), .A(n16201), .B(n16200), .ZN(
        P1_U2992) );
  INV_X1 U19358 ( .A(n16203), .ZN(n20198) );
  AOI222_X1 U19359 ( .A1(n16206), .A2(n11980), .B1(n16205), .B2(n20213), .C1(
        n20198), .C2(n16204), .ZN(n16208) );
  OAI211_X1 U19360 ( .C1(n16210), .C2(n16209), .A(n16208), .B(n16207), .ZN(
        P1_U2994) );
  AOI22_X1 U19361 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n16319), .B1(n16212), 
        .B2(n16211), .ZN(n16221) );
  INV_X1 U19362 ( .A(n16213), .ZN(n16215) );
  AOI22_X1 U19363 ( .A1(n16215), .A2(n20285), .B1(n20282), .B2(n16214), .ZN(
        n16220) );
  INV_X1 U19364 ( .A(n16216), .ZN(n16218) );
  OAI21_X1 U19365 ( .B1(n16218), .B2(n16217), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16219) );
  NAND3_X1 U19366 ( .A1(n16221), .A2(n16220), .A3(n16219), .ZN(P1_U3005) );
  AOI22_X1 U19367 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n16319), .B1(n16222), 
        .B2(n11915), .ZN(n16228) );
  INV_X1 U19368 ( .A(n16223), .ZN(n16226) );
  INV_X1 U19369 ( .A(n16224), .ZN(n16225) );
  AOI22_X1 U19370 ( .A1(n16226), .A2(n20285), .B1(n20282), .B2(n16225), .ZN(
        n16227) );
  OAI211_X1 U19371 ( .C1(n16229), .C2(n11915), .A(n16228), .B(n16227), .ZN(
        P1_U3008) );
  AOI22_X1 U19372 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n16230), .B1(
        n16319), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16236) );
  INV_X1 U19373 ( .A(n16231), .ZN(n16234) );
  INV_X1 U19374 ( .A(n16232), .ZN(n16233) );
  AOI22_X1 U19375 ( .A1(n16234), .A2(n20285), .B1(n20282), .B2(n16233), .ZN(
        n16235) );
  OAI211_X1 U19376 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n16237), .A(
        n16236), .B(n16235), .ZN(P1_U3012) );
  AOI21_X1 U19377 ( .B1(n16287), .B2(n16240), .A(n16238), .ZN(n16256) );
  NOR3_X1 U19378 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16240), .A3(
        n16239), .ZN(n16245) );
  INV_X1 U19379 ( .A(n16241), .ZN(n16242) );
  OAI22_X1 U19380 ( .A1(n16243), .A2(n16260), .B1(n16259), .B2(n16242), .ZN(
        n16244) );
  NOR3_X1 U19381 ( .A1(n16246), .A2(n16245), .A3(n16244), .ZN(n16247) );
  OAI21_X1 U19382 ( .B1(n16256), .B2(n16248), .A(n16247), .ZN(P1_U3013) );
  AOI21_X1 U19383 ( .B1(n16250), .B2(n16249), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16255) );
  AOI22_X1 U19384 ( .A1(n16252), .A2(n20285), .B1(n20282), .B2(n16251), .ZN(
        n16254) );
  NAND2_X1 U19385 ( .A1(n16319), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n16253) );
  OAI211_X1 U19386 ( .C1(n16256), .C2(n16255), .A(n16254), .B(n16253), .ZN(
        P1_U3014) );
  NOR3_X1 U19387 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16328), .A3(
        n16257), .ZN(n16263) );
  OAI22_X1 U19388 ( .A1(n16261), .A2(n16260), .B1(n16259), .B2(n16258), .ZN(
        n16262) );
  NOR2_X1 U19389 ( .A1(n16263), .A2(n16262), .ZN(n16265) );
  NAND2_X1 U19390 ( .A1(n16319), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n16264) );
  OAI211_X1 U19391 ( .C1(n16274), .C2(n16266), .A(n16265), .B(n16264), .ZN(
        P1_U3017) );
  AOI22_X1 U19392 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n16319), .B1(n16273), 
        .B2(n16267), .ZN(n16272) );
  INV_X1 U19393 ( .A(n16268), .ZN(n16270) );
  AOI22_X1 U19394 ( .A1(n16270), .A2(n20285), .B1(n20282), .B2(n16269), .ZN(
        n16271) );
  OAI211_X1 U19395 ( .C1(n16274), .C2(n16273), .A(n16272), .B(n16271), .ZN(
        P1_U3018) );
  AOI22_X1 U19396 ( .A1(n16275), .A2(n20282), .B1(n16319), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n16280) );
  NOR2_X1 U19397 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16328), .ZN(
        n16277) );
  AOI22_X1 U19398 ( .A1(n16278), .A2(n20285), .B1(n16277), .B2(n16276), .ZN(
        n16279) );
  OAI211_X1 U19399 ( .C1(n16281), .C2(n11911), .A(n16280), .B(n16279), .ZN(
        P1_U3020) );
  INV_X1 U19400 ( .A(n16290), .ZN(n16282) );
  OAI21_X1 U19401 ( .B1(n16284), .B2(n16283), .A(n16282), .ZN(n16286) );
  AOI21_X1 U19402 ( .B1(n16287), .B2(n16286), .A(n16285), .ZN(n16304) );
  AOI222_X1 U19403 ( .A1(n16289), .A2(n20285), .B1(n20282), .B2(n16288), .C1(
        P1_REIP_REG_10__SCAN_IN), .C2(n16319), .ZN(n16292) );
  NOR2_X1 U19404 ( .A1(n16290), .A2(n16328), .ZN(n16299) );
  OAI221_X1 U19405 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n14627), .C2(n16303), .A(
        n16299), .ZN(n16291) );
  OAI211_X1 U19406 ( .C1(n16304), .C2(n14627), .A(n16292), .B(n16291), .ZN(
        P1_U3021) );
  AOI21_X1 U19407 ( .B1(n9800), .B2(n16294), .A(n16293), .ZN(n16296) );
  OR2_X1 U19408 ( .A1(n16296), .A2(n16295), .ZN(n20204) );
  INV_X1 U19409 ( .A(n20204), .ZN(n20153) );
  INV_X1 U19410 ( .A(n16297), .ZN(n16298) );
  AOI21_X1 U19411 ( .B1(n20153), .B2(n20282), .A(n16298), .ZN(n16302) );
  AOI22_X1 U19412 ( .A1(n16300), .A2(n20285), .B1(n16299), .B2(n16303), .ZN(
        n16301) );
  OAI211_X1 U19413 ( .C1(n16304), .C2(n16303), .A(n16302), .B(n16301), .ZN(
        P1_U3022) );
  INV_X1 U19414 ( .A(n16305), .ZN(n16307) );
  AOI21_X1 U19415 ( .B1(n16307), .B2(n20282), .A(n16306), .ZN(n16317) );
  INV_X1 U19416 ( .A(n16308), .ZN(n16311) );
  AOI21_X1 U19417 ( .B1(n16311), .B2(n16310), .A(n16309), .ZN(n16333) );
  OAI21_X1 U19418 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16312), .A(
        n16333), .ZN(n16318) );
  AOI22_X1 U19419 ( .A1(n16313), .A2(n20285), .B1(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n16318), .ZN(n16316) );
  INV_X1 U19420 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16314) );
  NOR2_X1 U19421 ( .A1(n16332), .A2(n16328), .ZN(n16320) );
  OAI221_X1 U19422 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16314), .C2(n16324), .A(
        n16320), .ZN(n16315) );
  NAND3_X1 U19423 ( .A1(n16317), .A2(n16316), .A3(n16315), .ZN(P1_U3023) );
  INV_X1 U19424 ( .A(n16318), .ZN(n16325) );
  AOI22_X1 U19425 ( .A1(n20165), .A2(n20282), .B1(n16319), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16323) );
  AOI22_X1 U19426 ( .A1(n16321), .A2(n20285), .B1(n16320), .B2(n16324), .ZN(
        n16322) );
  OAI211_X1 U19427 ( .C1(n16325), .C2(n16324), .A(n16323), .B(n16322), .ZN(
        P1_U3024) );
  AOI21_X1 U19428 ( .B1(n20282), .B2(n20182), .A(n16326), .ZN(n16327) );
  OAI21_X1 U19429 ( .B1(n16328), .B2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n16327), .ZN(n16329) );
  AOI21_X1 U19430 ( .B1(n16330), .B2(n20285), .A(n16329), .ZN(n16331) );
  OAI21_X1 U19431 ( .B1(n16333), .B2(n16332), .A(n16331), .ZN(P1_U3025) );
  NAND4_X1 U19432 ( .A1(n16337), .A2(n16336), .A3(n16335), .A4(n16334), .ZN(
        n16338) );
  OAI21_X1 U19433 ( .B1(n16340), .B2(n16339), .A(n16338), .ZN(P1_U3468) );
  OAI221_X1 U19434 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(
        P1_STATEBS16_REG_SCAN_IN), .C1(n20846), .C2(n20850), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n20754) );
  NAND2_X1 U19435 ( .A1(n16341), .A2(n20754), .ZN(n16342) );
  AOI22_X1 U19436 ( .A1(n16345), .A2(n16344), .B1(n16343), .B2(n16342), .ZN(
        P1_U3162) );
  OAI21_X1 U19437 ( .B1(n20752), .B2(n20609), .A(n16346), .ZN(P1_U3466) );
  AOI22_X1 U19438 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19308), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n19325), .ZN(n16357) );
  AOI22_X1 U19439 ( .A1(n16347), .A2(n19324), .B1(P2_EBX_REG_29__SCAN_IN), 
        .B2(n19326), .ZN(n16356) );
  INV_X1 U19440 ( .A(n16348), .ZN(n16350) );
  AOI22_X1 U19441 ( .A1(n16350), .A2(n19314), .B1(n16349), .B2(n19327), .ZN(
        n16355) );
  OAI211_X1 U19442 ( .C1(n16353), .C2(n16352), .A(n19315), .B(n16351), .ZN(
        n16354) );
  NAND4_X1 U19443 ( .A1(n16357), .A2(n16356), .A3(n16355), .A4(n16354), .ZN(
        P2_U2826) );
  OAI22_X1 U19444 ( .A1(n10157), .A2(n19334), .B1(n20036), .B2(n19301), .ZN(
        n16359) );
  NOR2_X1 U19445 ( .A1(n19303), .A2(n10772), .ZN(n16358) );
  AOI211_X1 U19446 ( .C1(n16360), .C2(n19324), .A(n16359), .B(n16358), .ZN(
        n16361) );
  INV_X1 U19447 ( .A(n16361), .ZN(n16362) );
  AOI21_X1 U19448 ( .B1(n16363), .B2(n19314), .A(n16362), .ZN(n16368) );
  OAI211_X1 U19449 ( .C1(n16366), .C2(n16365), .A(n19315), .B(n16364), .ZN(
        n16367) );
  OAI211_X1 U19450 ( .C1(n19320), .C2(n16369), .A(n16368), .B(n16367), .ZN(
        P2_U2827) );
  AOI22_X1 U19451 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n19308), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n19325), .ZN(n16382) );
  INV_X1 U19452 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n16370) );
  OAI22_X1 U19453 ( .A1(n16371), .A2(n19304), .B1(n19303), .B2(n16370), .ZN(
        n16372) );
  INV_X1 U19454 ( .A(n16372), .ZN(n16381) );
  OAI22_X1 U19455 ( .A1(n16374), .A2(n19321), .B1(n16373), .B2(n19320), .ZN(
        n16375) );
  INV_X1 U19456 ( .A(n16375), .ZN(n16380) );
  OAI211_X1 U19457 ( .C1(n16378), .C2(n16377), .A(n19315), .B(n16376), .ZN(
        n16379) );
  NAND4_X1 U19458 ( .A1(n16382), .A2(n16381), .A3(n16380), .A4(n16379), .ZN(
        P2_U2828) );
  AOI22_X1 U19459 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19308), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n19325), .ZN(n16393) );
  AOI22_X1 U19460 ( .A1(n16383), .A2(n19324), .B1(P2_EBX_REG_26__SCAN_IN), 
        .B2(n19326), .ZN(n16392) );
  INV_X1 U19461 ( .A(n16384), .ZN(n16386) );
  AOI22_X1 U19462 ( .A1(n16386), .A2(n19314), .B1(n16385), .B2(n19327), .ZN(
        n16391) );
  OAI211_X1 U19463 ( .C1(n16389), .C2(n16388), .A(n19315), .B(n16387), .ZN(
        n16390) );
  NAND4_X1 U19464 ( .A1(n16393), .A2(n16392), .A3(n16391), .A4(n16390), .ZN(
        P2_U2829) );
  AOI22_X1 U19465 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19308), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19325), .ZN(n16404) );
  AOI22_X1 U19466 ( .A1(n16394), .A2(n19324), .B1(P2_EBX_REG_25__SCAN_IN), 
        .B2(n19326), .ZN(n16403) );
  OAI22_X1 U19467 ( .A1(n16396), .A2(n19321), .B1(n16395), .B2(n19320), .ZN(
        n16397) );
  INV_X1 U19468 ( .A(n16397), .ZN(n16402) );
  OAI211_X1 U19469 ( .C1(n16400), .C2(n16399), .A(n19315), .B(n16398), .ZN(
        n16401) );
  NAND4_X1 U19470 ( .A1(n16404), .A2(n16403), .A3(n16402), .A4(n16401), .ZN(
        P2_U2830) );
  AOI22_X1 U19471 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19308), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19325), .ZN(n16415) );
  AOI22_X1 U19472 ( .A1(n16405), .A2(n19324), .B1(P2_EBX_REG_24__SCAN_IN), 
        .B2(n19326), .ZN(n16414) );
  OAI22_X1 U19473 ( .A1(n16407), .A2(n19321), .B1(n16406), .B2(n19320), .ZN(
        n16408) );
  INV_X1 U19474 ( .A(n16408), .ZN(n16413) );
  OAI211_X1 U19475 ( .C1(n16411), .C2(n16410), .A(n19315), .B(n16409), .ZN(
        n16412) );
  NAND4_X1 U19476 ( .A1(n16415), .A2(n16414), .A3(n16413), .A4(n16412), .ZN(
        P2_U2831) );
  AOI22_X1 U19477 ( .A1(n16417), .A2(n16416), .B1(n19382), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n16424) );
  AOI22_X1 U19478 ( .A1(n16419), .A2(BUF1_REG_23__SCAN_IN), .B1(n16418), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n16423) );
  AOI22_X1 U19479 ( .A1(n16421), .A2(n19385), .B1(n19383), .B2(n16420), .ZN(
        n16422) );
  NAND3_X1 U19480 ( .A1(n16424), .A2(n16423), .A3(n16422), .ZN(P2_U2896) );
  AOI211_X1 U19481 ( .C1(n16426), .C2(n16425), .A(n19429), .B(n9752), .ZN(
        n16430) );
  AOI22_X1 U19482 ( .A1(P2_REIP_REG_17__SCAN_IN), .A2(n19427), .B1(n19426), 
        .B2(n19222), .ZN(n16427) );
  OAI21_X1 U19483 ( .B1(n16428), .B2(n19438), .A(n16427), .ZN(n16429) );
  AOI211_X1 U19484 ( .C1(n16431), .C2(n16495), .A(n16430), .B(n16429), .ZN(
        n16432) );
  OAI21_X1 U19485 ( .B1(n16433), .B2(n19227), .A(n16432), .ZN(P2_U2997) );
  AOI22_X1 U19486 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19427), .B1(n19426), 
        .B2(n19246), .ZN(n16440) );
  NAND2_X1 U19487 ( .A1(n16435), .A2(n16434), .ZN(n16436) );
  XNOR2_X1 U19488 ( .A(n16437), .B(n16436), .ZN(n16513) );
  INV_X1 U19489 ( .A(n16513), .ZN(n16438) );
  INV_X1 U19490 ( .A(n16508), .ZN(n19252) );
  XNOR2_X1 U19491 ( .A(n15377), .B(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16510) );
  AOI222_X1 U19492 ( .A1(n16438), .A2(n16495), .B1(n19435), .B2(n19252), .C1(
        n16496), .C2(n16510), .ZN(n16439) );
  OAI211_X1 U19493 ( .C1(n19249), .C2(n19438), .A(n16440), .B(n16439), .ZN(
        P2_U2999) );
  AOI22_X1 U19494 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n16477), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19427), .ZN(n16445) );
  OAI22_X1 U19495 ( .A1(n16442), .A2(n19429), .B1(n16441), .B2(n19431), .ZN(
        n16443) );
  AOI21_X1 U19496 ( .B1(n19435), .B2(n19262), .A(n16443), .ZN(n16444) );
  OAI211_X1 U19497 ( .C1(n16491), .C2(n16446), .A(n16445), .B(n16444), .ZN(
        P2_U3000) );
  AOI22_X1 U19498 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19427), .B1(n19426), 
        .B2(n16447), .ZN(n16457) );
  INV_X1 U19499 ( .A(n16448), .ZN(n16471) );
  NAND2_X1 U19500 ( .A1(n16471), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16450) );
  AOI21_X1 U19501 ( .B1(n12652), .B2(n16450), .A(n16449), .ZN(n16522) );
  NAND2_X1 U19502 ( .A1(n16452), .A2(n16451), .ZN(n16453) );
  XNOR2_X1 U19503 ( .A(n16454), .B(n16453), .ZN(n16518) );
  AOI222_X1 U19504 ( .A1(n16522), .A2(n16496), .B1(n16495), .B2(n16518), .C1(
        n19435), .C2(n16455), .ZN(n16456) );
  OAI211_X1 U19505 ( .C1(n16458), .C2(n19438), .A(n16457), .B(n16456), .ZN(
        P2_U3001) );
  AOI22_X1 U19506 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16477), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19427), .ZN(n16463) );
  OAI22_X1 U19507 ( .A1(n16460), .A2(n19429), .B1(n16459), .B2(n19431), .ZN(
        n16461) );
  AOI21_X1 U19508 ( .B1(n19435), .B2(n19274), .A(n16461), .ZN(n16462) );
  OAI211_X1 U19509 ( .C1(n16491), .C2(n19267), .A(n16463), .B(n16462), .ZN(
        P2_U3002) );
  AOI22_X1 U19510 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19427), .B1(n19426), 
        .B2(n16464), .ZN(n16475) );
  NOR2_X1 U19511 ( .A1(n10072), .A2(n16466), .ZN(n16470) );
  NOR2_X1 U19512 ( .A1(n16468), .A2(n16467), .ZN(n16469) );
  XNOR2_X1 U19513 ( .A(n16470), .B(n16469), .ZN(n16536) );
  INV_X1 U19514 ( .A(n19281), .ZN(n16473) );
  INV_X1 U19515 ( .A(n16479), .ZN(n16472) );
  AOI21_X1 U19516 ( .B1(n16542), .B2(n16472), .A(n16471), .ZN(n16539) );
  AOI222_X1 U19517 ( .A1(n16536), .A2(n16495), .B1(n19435), .B2(n16473), .C1(
        n16496), .C2(n16539), .ZN(n16474) );
  OAI211_X1 U19518 ( .C1(n16476), .C2(n19438), .A(n16475), .B(n16474), .ZN(
        P2_U3003) );
  AOI22_X1 U19519 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16477), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19427), .ZN(n16489) );
  AND2_X1 U19520 ( .A1(n15592), .A2(n16545), .ZN(n16478) );
  OR2_X1 U19521 ( .A1(n16479), .A2(n16478), .ZN(n16552) );
  NOR2_X1 U19522 ( .A1(n16481), .A2(n16480), .ZN(n16485) );
  NAND2_X1 U19523 ( .A1(n16483), .A2(n16482), .ZN(n16484) );
  XNOR2_X1 U19524 ( .A(n16485), .B(n16484), .ZN(n16555) );
  OAI22_X1 U19525 ( .A1(n16552), .A2(n19429), .B1(n16555), .B2(n19431), .ZN(
        n16486) );
  AOI21_X1 U19526 ( .B1(n19435), .B2(n16487), .A(n16486), .ZN(n16488) );
  OAI211_X1 U19527 ( .C1(n16491), .C2(n16490), .A(n16489), .B(n16488), .ZN(
        P2_U3004) );
  AOI22_X1 U19528 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19427), .B1(n19426), 
        .B2(n16492), .ZN(n16499) );
  AOI222_X1 U19529 ( .A1(n16497), .A2(n16496), .B1(n16495), .B2(n16494), .C1(
        n19435), .C2(n16493), .ZN(n16498) );
  OAI211_X1 U19530 ( .C1(n16500), .C2(n19438), .A(n16499), .B(n16498), .ZN(
        P2_U3005) );
  NAND2_X1 U19531 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19427), .ZN(n16501) );
  OAI21_X1 U19532 ( .B1(n16502), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n16501), .ZN(n16503) );
  AOI21_X1 U19533 ( .B1(n16582), .B2(n19251), .A(n16503), .ZN(n16504) );
  OAI21_X1 U19534 ( .B1(n16506), .B2(n16505), .A(n16504), .ZN(n16507) );
  INV_X1 U19535 ( .A(n16507), .ZN(n16512) );
  NOR2_X1 U19536 ( .A1(n16508), .A2(n16574), .ZN(n16509) );
  AOI21_X1 U19537 ( .B1(n16510), .B2(n16566), .A(n16509), .ZN(n16511) );
  OAI211_X1 U19538 ( .C1(n16513), .C2(n16570), .A(n16512), .B(n16511), .ZN(
        P2_U3031) );
  OAI21_X1 U19539 ( .B1(n16515), .B2(n16514), .A(n12652), .ZN(n16516) );
  AOI22_X1 U19540 ( .A1(n16517), .A2(n16516), .B1(n16582), .B2(n19344), .ZN(
        n16524) );
  INV_X1 U19541 ( .A(n16518), .ZN(n16520) );
  OAI22_X1 U19542 ( .A1(n16520), .A2(n16570), .B1(n16574), .B2(n16519), .ZN(
        n16521) );
  AOI21_X1 U19543 ( .B1(n16566), .B2(n16522), .A(n16521), .ZN(n16523) );
  OAI211_X1 U19544 ( .C1(n20011), .C2(n19300), .A(n16524), .B(n16523), .ZN(
        P2_U3033) );
  NAND2_X1 U19545 ( .A1(n16526), .A2(n16525), .ZN(n16544) );
  NAND2_X1 U19546 ( .A1(n16528), .A2(n16527), .ZN(n16531) );
  INV_X1 U19547 ( .A(n16529), .ZN(n16530) );
  NAND2_X1 U19548 ( .A1(n16531), .A2(n16530), .ZN(n19350) );
  AOI211_X1 U19549 ( .C1(n16545), .C2(n16542), .A(n16532), .B(n16546), .ZN(
        n16533) );
  AOI21_X1 U19550 ( .B1(n19427), .B2(P2_REIP_REG_11__SCAN_IN), .A(n16533), 
        .ZN(n16534) );
  OAI21_X1 U19551 ( .B1(n16563), .B2(n19350), .A(n16534), .ZN(n16535) );
  INV_X1 U19552 ( .A(n16535), .ZN(n16541) );
  INV_X1 U19553 ( .A(n16536), .ZN(n16537) );
  OAI22_X1 U19554 ( .A1(n16537), .A2(n16570), .B1(n16574), .B2(n19281), .ZN(
        n16538) );
  AOI21_X1 U19555 ( .B1(n16566), .B2(n16539), .A(n16538), .ZN(n16540) );
  OAI211_X1 U19556 ( .C1(n16542), .C2(n16544), .A(n16541), .B(n16540), .ZN(
        P2_U3035) );
  NAND2_X1 U19557 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n19427), .ZN(n16543) );
  OAI221_X1 U19558 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16546), 
        .C1(n16545), .C2(n16544), .A(n16543), .ZN(n16550) );
  OAI22_X1 U19559 ( .A1(n16548), .A2(n16563), .B1(n16574), .B2(n16547), .ZN(
        n16549) );
  NOR2_X1 U19560 ( .A1(n16550), .A2(n16549), .ZN(n16551) );
  OAI21_X1 U19561 ( .B1(n16552), .B2(n16587), .A(n16551), .ZN(n16553) );
  INV_X1 U19562 ( .A(n16553), .ZN(n16554) );
  OAI21_X1 U19563 ( .B1(n16555), .B2(n16570), .A(n16554), .ZN(P2_U3036) );
  AOI211_X1 U19564 ( .C1(n16558), .C2(n16561), .A(n16557), .B(n16556), .ZN(
        n16565) );
  OAI21_X1 U19565 ( .B1(n16560), .B2(n9774), .A(n16559), .ZN(n19354) );
  OAI22_X1 U19566 ( .A1(n16563), .A2(n19354), .B1(n16562), .B2(n16561), .ZN(
        n16564) );
  AOI211_X1 U19567 ( .C1(n19427), .C2(P2_REIP_REG_8__SCAN_IN), .A(n16565), .B(
        n16564), .ZN(n16569) );
  AOI22_X1 U19568 ( .A1(n16567), .A2(n16566), .B1(n16592), .B2(n19296), .ZN(
        n16568) );
  OAI211_X1 U19569 ( .C1(n16571), .C2(n16570), .A(n16569), .B(n16568), .ZN(
        P2_U3038) );
  AOI22_X1 U19570 ( .A1(n16572), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        n16582), .B2(n20069), .ZN(n16581) );
  INV_X1 U19571 ( .A(n13270), .ZN(n16573) );
  OAI22_X1 U19572 ( .A1(n16575), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        n16574), .B2(n16573), .ZN(n16578) );
  NOR2_X1 U19573 ( .A1(n16576), .A2(n16587), .ZN(n16577) );
  AOI211_X1 U19574 ( .C1(n16579), .C2(n16584), .A(n16578), .B(n16577), .ZN(
        n16580) );
  OAI211_X1 U19575 ( .C1(n10684), .C2(n19300), .A(n16581), .B(n16580), .ZN(
        P2_U3043) );
  AOI22_X1 U19576 ( .A1(n16584), .A2(n16583), .B1(n16582), .B2(n19386), .ZN(
        n16594) );
  OAI22_X1 U19577 ( .A1(n16588), .A2(n16587), .B1(n16586), .B2(n16585), .ZN(
        n16589) );
  AOI211_X1 U19578 ( .C1(n16592), .C2(n16591), .A(n16590), .B(n16589), .ZN(
        n16593) );
  OAI211_X1 U19579 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n16595), .A(
        n16594), .B(n16593), .ZN(P2_U3046) );
  NOR2_X1 U19580 ( .A1(n16597), .A2(n16596), .ZN(n20091) );
  OR2_X1 U19581 ( .A1(n19976), .A2(n20091), .ZN(n16600) );
  AOI211_X1 U19582 ( .C1(P2_STATE2_REG_0__SCAN_IN), .C2(n16600), .A(n16599), 
        .B(n16598), .ZN(n16604) );
  NAND2_X1 U19583 ( .A1(n19976), .A2(n20118), .ZN(n16601) );
  OAI211_X1 U19584 ( .C1(n19159), .C2(n16602), .A(n19974), .B(n16601), .ZN(
        n16603) );
  OAI211_X1 U19585 ( .C1(n16606), .C2(n16605), .A(n16604), .B(n16603), .ZN(
        P2_U3176) );
  INV_X1 U19586 ( .A(n16607), .ZN(n18918) );
  OAI22_X2 U19587 ( .A1(n16608), .A2(n18921), .B1(n18918), .B2(n16668), .ZN(
        n18974) );
  NOR2_X2 U19588 ( .A1(n19136), .A2(n16787), .ZN(n18136) );
  NOR2_X1 U19589 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17952), .ZN(
        n16611) );
  AOI21_X1 U19590 ( .B1(n17952), .B2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n16611), .ZN(n16617) );
  AND2_X1 U19591 ( .A1(n18050), .A2(n16609), .ZN(n16615) );
  INV_X1 U19592 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16654) );
  OAI21_X1 U19593 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n16654), .A(
        n16610), .ZN(n16612) );
  OAI22_X1 U19594 ( .A1(n16615), .A2(n16612), .B1(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16611), .ZN(n16616) );
  NAND2_X1 U19595 ( .A1(n16617), .A2(n16613), .ZN(n16614) );
  OAI22_X1 U19596 ( .A1(n16617), .A2(n16616), .B1(n16615), .B2(n16614), .ZN(
        n16664) );
  NAND2_X1 U19597 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17814) );
  NAND2_X1 U19598 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18102) );
  INV_X1 U19599 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18104) );
  NAND2_X1 U19600 ( .A1(n18083), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18075) );
  NAND2_X1 U19601 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18054) );
  INV_X1 U19602 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17081) );
  NAND2_X1 U19603 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17987) );
  NAND2_X1 U19604 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17935) );
  NAND2_X1 U19605 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n17919), .ZN(
        n17893) );
  NAND2_X1 U19606 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17894) );
  NAND2_X1 U19607 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17853) );
  NAND2_X1 U19608 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16639), .ZN(
        n16618) );
  XOR2_X2 U19609 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n16618), .Z(
        n17146) );
  INV_X1 U19610 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19069) );
  NOR2_X1 U19611 ( .A1(n19069), .A2(n18447), .ZN(n16659) );
  INV_X1 U19612 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17802) );
  NAND3_X1 U19613 ( .A1(n16619), .A2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17801) );
  NOR2_X1 U19614 ( .A1(n17802), .A2(n17801), .ZN(n17771) );
  NAND3_X1 U19615 ( .A1(n17771), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16643) );
  NOR2_X1 U19616 ( .A1(n16845), .A2(n16643), .ZN(n16620) );
  INV_X1 U19617 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18139) );
  NAND2_X1 U19618 ( .A1(n18986), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17977) );
  NAND2_X1 U19619 ( .A1(n16620), .A2(n17837), .ZN(n16632) );
  INV_X1 U19620 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16832) );
  XOR2_X1 U19621 ( .A(n16832), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16622) );
  NOR2_X1 U19622 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17881), .ZN(
        n16640) );
  INV_X1 U19623 ( .A(n16809), .ZN(n16621) );
  OR2_X1 U19624 ( .A1(n18819), .A2(n16620), .ZN(n16644) );
  OAI211_X1 U19625 ( .C1(n16621), .C2(n17977), .A(n18144), .B(n16644), .ZN(
        n16649) );
  NOR2_X1 U19626 ( .A1(n16640), .A2(n16649), .ZN(n16631) );
  OAI22_X1 U19627 ( .A1(n16632), .A2(n16622), .B1(n16631), .B2(n16832), .ZN(
        n16623) );
  AOI211_X1 U19628 ( .C1(n17980), .C2(n17133), .A(n16659), .B(n16623), .ZN(
        n16627) );
  INV_X1 U19629 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19096) );
  NAND3_X1 U19630 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n19096), .ZN(n16656) );
  OAI21_X1 U19631 ( .B1(n16629), .B2(n16654), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16624) );
  OAI21_X1 U19632 ( .B1(n16672), .B2(n16656), .A(n16624), .ZN(n16661) );
  INV_X1 U19633 ( .A(n18136), .ZN(n18148) );
  NOR2_X2 U19634 ( .A1(n16666), .A2(n18148), .ZN(n18012) );
  NAND2_X1 U19635 ( .A1(n16628), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16625) );
  XNOR2_X1 U19636 ( .A(n16625), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16660) );
  AOI22_X1 U19637 ( .A1(n18132), .A2(n16661), .B1(n18012), .B2(n16660), .ZN(
        n16626) );
  OAI211_X1 U19638 ( .C1(n18052), .C2(n16664), .A(n16627), .B(n16626), .ZN(
        P3_U2799) );
  XOR2_X1 U19639 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n16639), .Z(
        n16835) );
  INV_X1 U19640 ( .A(n18012), .ZN(n18051) );
  OR2_X1 U19641 ( .A1(n18051), .A2(n16628), .ZN(n16646) );
  NAND2_X1 U19642 ( .A1(n18132), .A2(n16629), .ZN(n16652) );
  AOI21_X1 U19643 ( .B1(n16646), .B2(n16652), .A(n16654), .ZN(n16634) );
  INV_X1 U19644 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16836) );
  OAI221_X1 U19645 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16632), .C1(
        n16836), .C2(n16631), .A(n16630), .ZN(n16633) );
  AOI211_X1 U19646 ( .C1(n17980), .C2(n16835), .A(n16634), .B(n16633), .ZN(
        n16637) );
  INV_X1 U19647 ( .A(n18309), .ZN(n18329) );
  NAND3_X1 U19648 ( .A1(n18151), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n17906), .ZN(n17844) );
  NOR2_X1 U19649 ( .A1(n18160), .A2(n17844), .ZN(n17795) );
  NAND3_X1 U19650 ( .A1(n16635), .A2(n17795), .A3(n16654), .ZN(n16636) );
  OAI211_X1 U19651 ( .C1(n16638), .C2(n18052), .A(n16637), .B(n16636), .ZN(
        P3_U2800) );
  AOI21_X1 U19652 ( .B1(n16845), .B2(n16809), .A(n16639), .ZN(n16844) );
  OAI21_X1 U19653 ( .B1(n16640), .B2(n17980), .A(n16844), .ZN(n16641) );
  OAI211_X1 U19654 ( .C1(n16644), .C2(n16643), .A(n16642), .B(n16641), .ZN(
        n16648) );
  NOR2_X1 U19655 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16671), .ZN(
        n16647) );
  OAI221_X1 U19656 ( .B1(n16652), .B2(n16651), .C1(n16652), .C2(n16672), .A(
        n16650), .ZN(P3_U2801) );
  AOI21_X1 U19657 ( .B1(n18376), .B2(n16654), .A(n16653), .ZN(n16657) );
  OAI22_X1 U19658 ( .A1(n16657), .A2(n19096), .B1(n16656), .B2(n16655), .ZN(
        n16658) );
  AOI211_X1 U19659 ( .C1(n16660), .C2(n18384), .A(n16659), .B(n16658), .ZN(
        n16663) );
  NAND2_X1 U19660 ( .A1(n18463), .A2(n16661), .ZN(n16662) );
  OAI211_X1 U19661 ( .C1(n16664), .C2(n18388), .A(n16663), .B(n16662), .ZN(
        P3_U2831) );
  NAND2_X1 U19662 ( .A1(n16665), .A2(n17779), .ZN(n16677) );
  INV_X1 U19663 ( .A(n16666), .ZN(n17628) );
  NAND2_X1 U19664 ( .A1(n18919), .A2(n17628), .ZN(n18330) );
  OAI22_X1 U19665 ( .A1(n18921), .A2(n18286), .B1(n18277), .B2(n18330), .ZN(
        n18242) );
  NOR2_X1 U19666 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n16667), .ZN(
        n17783) );
  OAI211_X1 U19667 ( .C1(n16671), .C2(n18330), .A(n18391), .B(n16670), .ZN(
        n16674) );
  INV_X1 U19668 ( .A(n18921), .ZN(n18317) );
  AND2_X1 U19669 ( .A1(n16672), .A2(n18317), .ZN(n16673) );
  INV_X1 U19670 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19065) );
  NOR2_X1 U19671 ( .A1(n18447), .A2(n19065), .ZN(n17774) );
  NAND3_X1 U19672 ( .A1(n17780), .A2(n17789), .A3(n18362), .ZN(n16675) );
  OAI211_X1 U19673 ( .C1(n16677), .C2(n18467), .A(n16676), .B(n16675), .ZN(
        P3_U2834) );
  NOR3_X1 U19674 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16679) );
  NOR4_X1 U19675 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16678) );
  NAND4_X1 U19676 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16679), .A3(n16678), .A4(
        U215), .ZN(U213) );
  INV_X1 U19677 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16774) );
  INV_X2 U19678 ( .A(U214), .ZN(n16736) );
  INV_X1 U19679 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16775) );
  OAI222_X1 U19680 ( .A1(U212), .A2(n16774), .B1(n16738), .B2(n19484), .C1(
        U214), .C2(n16775), .ZN(U216) );
  AOI22_X1 U19681 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16735), .ZN(n16681) );
  OAI21_X1 U19682 ( .B1(n16682), .B2(n16738), .A(n16681), .ZN(U217) );
  AOI22_X1 U19683 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16735), .ZN(n16683) );
  OAI21_X1 U19684 ( .B1(n19473), .B2(n16738), .A(n16683), .ZN(U218) );
  AOI22_X1 U19685 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16735), .ZN(n16684) );
  OAI21_X1 U19686 ( .B1(n16685), .B2(n16738), .A(n16684), .ZN(U219) );
  AOI22_X1 U19687 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16735), .ZN(n16686) );
  OAI21_X1 U19688 ( .B1(n19464), .B2(n16738), .A(n16686), .ZN(U220) );
  AOI22_X1 U19689 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16735), .ZN(n16687) );
  OAI21_X1 U19690 ( .B1(n19457), .B2(n16738), .A(n16687), .ZN(U221) );
  AOI22_X1 U19691 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16735), .ZN(n16688) );
  OAI21_X1 U19692 ( .B1(n16689), .B2(n16738), .A(n16688), .ZN(U222) );
  AOI22_X1 U19693 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16735), .ZN(n16690) );
  OAI21_X1 U19694 ( .B1(n16691), .B2(n16738), .A(n16690), .ZN(U223) );
  INV_X1 U19695 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16693) );
  AOI22_X1 U19696 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16735), .ZN(n16692) );
  OAI21_X1 U19697 ( .B1(n16693), .B2(n16738), .A(n16692), .ZN(U224) );
  INV_X1 U19698 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16695) );
  AOI22_X1 U19699 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16735), .ZN(n16694) );
  OAI21_X1 U19700 ( .B1(n16695), .B2(n16738), .A(n16694), .ZN(U225) );
  AOI22_X1 U19701 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16735), .ZN(n16696) );
  OAI21_X1 U19702 ( .B1(n15184), .B2(n16738), .A(n16696), .ZN(U226) );
  INV_X1 U19703 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16698) );
  AOI22_X1 U19704 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16735), .ZN(n16697) );
  OAI21_X1 U19705 ( .B1(n16698), .B2(n16738), .A(n16697), .ZN(U227) );
  AOI22_X1 U19706 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16735), .ZN(n16699) );
  OAI21_X1 U19707 ( .B1(n15205), .B2(n16738), .A(n16699), .ZN(U228) );
  INV_X1 U19708 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16701) );
  AOI22_X1 U19709 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16735), .ZN(n16700) );
  OAI21_X1 U19710 ( .B1(n16701), .B2(n16738), .A(n16700), .ZN(U229) );
  INV_X1 U19711 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16703) );
  AOI22_X1 U19712 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16735), .ZN(n16702) );
  OAI21_X1 U19713 ( .B1(n16703), .B2(n16738), .A(n16702), .ZN(U230) );
  INV_X1 U19714 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16705) );
  AOI22_X1 U19715 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16735), .ZN(n16704) );
  OAI21_X1 U19716 ( .B1(n16705), .B2(n16738), .A(n16704), .ZN(U231) );
  AOI22_X1 U19717 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16735), .ZN(n16706) );
  OAI21_X1 U19718 ( .B1(n13021), .B2(n16738), .A(n16706), .ZN(U232) );
  AOI22_X1 U19719 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16735), .ZN(n16707) );
  OAI21_X1 U19720 ( .B1(n16708), .B2(n16738), .A(n16707), .ZN(U233) );
  AOI22_X1 U19721 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16735), .ZN(n16709) );
  OAI21_X1 U19722 ( .B1(n16710), .B2(n16738), .A(n16709), .ZN(U234) );
  INV_X1 U19723 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16712) );
  AOI22_X1 U19724 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16735), .ZN(n16711) );
  OAI21_X1 U19725 ( .B1(n16712), .B2(n16738), .A(n16711), .ZN(U235) );
  AOI22_X1 U19726 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16735), .ZN(n16713) );
  OAI21_X1 U19727 ( .B1(n16714), .B2(n16738), .A(n16713), .ZN(U236) );
  AOI22_X1 U19728 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16735), .ZN(n16715) );
  OAI21_X1 U19729 ( .B1(n16716), .B2(n16738), .A(n16715), .ZN(U237) );
  AOI22_X1 U19730 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16735), .ZN(n16717) );
  OAI21_X1 U19731 ( .B1(n16718), .B2(n16738), .A(n16717), .ZN(U238) );
  AOI22_X1 U19732 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16735), .ZN(n16719) );
  OAI21_X1 U19733 ( .B1(n16720), .B2(n16738), .A(n16719), .ZN(U239) );
  INV_X1 U19734 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16722) );
  AOI22_X1 U19735 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16735), .ZN(n16721) );
  OAI21_X1 U19736 ( .B1(n16722), .B2(n16738), .A(n16721), .ZN(U240) );
  INV_X1 U19737 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16724) );
  AOI22_X1 U19738 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16735), .ZN(n16723) );
  OAI21_X1 U19739 ( .B1(n16724), .B2(n16738), .A(n16723), .ZN(U241) );
  AOI22_X1 U19740 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16735), .ZN(n16725) );
  OAI21_X1 U19741 ( .B1(n16726), .B2(n16738), .A(n16725), .ZN(U242) );
  INV_X1 U19742 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16728) );
  AOI22_X1 U19743 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16735), .ZN(n16727) );
  OAI21_X1 U19744 ( .B1(n16728), .B2(n16738), .A(n16727), .ZN(U243) );
  INV_X1 U19745 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16730) );
  AOI22_X1 U19746 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16735), .ZN(n16729) );
  OAI21_X1 U19747 ( .B1(n16730), .B2(n16738), .A(n16729), .ZN(U244) );
  AOI22_X1 U19748 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16735), .ZN(n16731) );
  OAI21_X1 U19749 ( .B1(n16732), .B2(n16738), .A(n16731), .ZN(U245) );
  AOI22_X1 U19750 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16735), .ZN(n16733) );
  OAI21_X1 U19751 ( .B1(n16734), .B2(n16738), .A(n16733), .ZN(U246) );
  AOI22_X1 U19752 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16736), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16735), .ZN(n16737) );
  OAI21_X1 U19753 ( .B1(n16739), .B2(n16738), .A(n16737), .ZN(U247) );
  OAI22_X1 U19754 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16772), .ZN(n16740) );
  INV_X1 U19755 ( .A(n16740), .ZN(U251) );
  OAI22_X1 U19756 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16772), .ZN(n16741) );
  INV_X1 U19757 ( .A(n16741), .ZN(U252) );
  INV_X1 U19758 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16742) );
  INV_X1 U19759 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18488) );
  AOI22_X1 U19760 ( .A1(n16768), .A2(n16742), .B1(n18488), .B2(U215), .ZN(U253) );
  INV_X1 U19761 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16743) );
  INV_X1 U19762 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18492) );
  AOI22_X1 U19763 ( .A1(n16772), .A2(n16743), .B1(n18492), .B2(U215), .ZN(U254) );
  INV_X1 U19764 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16744) );
  INV_X1 U19765 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18496) );
  AOI22_X1 U19766 ( .A1(n16772), .A2(n16744), .B1(n18496), .B2(U215), .ZN(U255) );
  INV_X1 U19767 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16745) );
  INV_X1 U19768 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18500) );
  AOI22_X1 U19769 ( .A1(n16768), .A2(n16745), .B1(n18500), .B2(U215), .ZN(U256) );
  INV_X1 U19770 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16746) );
  INV_X1 U19771 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18505) );
  AOI22_X1 U19772 ( .A1(n16772), .A2(n16746), .B1(n18505), .B2(U215), .ZN(U257) );
  INV_X1 U19773 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16747) );
  INV_X1 U19774 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18509) );
  AOI22_X1 U19775 ( .A1(n16768), .A2(n16747), .B1(n18509), .B2(U215), .ZN(U258) );
  INV_X1 U19776 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16748) );
  INV_X1 U19777 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17627) );
  AOI22_X1 U19778 ( .A1(n16768), .A2(n16748), .B1(n17627), .B2(U215), .ZN(U259) );
  INV_X1 U19779 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16749) );
  INV_X1 U19780 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17623) );
  AOI22_X1 U19781 ( .A1(n16772), .A2(n16749), .B1(n17623), .B2(U215), .ZN(U260) );
  OAI22_X1 U19782 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16768), .ZN(n16750) );
  INV_X1 U19783 ( .A(n16750), .ZN(U261) );
  INV_X1 U19784 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16751) );
  INV_X1 U19785 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17614) );
  AOI22_X1 U19786 ( .A1(n16772), .A2(n16751), .B1(n17614), .B2(U215), .ZN(U262) );
  INV_X1 U19787 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16752) );
  INV_X1 U19788 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17609) );
  AOI22_X1 U19789 ( .A1(n16768), .A2(n16752), .B1(n17609), .B2(U215), .ZN(U263) );
  OAI22_X1 U19790 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16768), .ZN(n16753) );
  INV_X1 U19791 ( .A(n16753), .ZN(U264) );
  OAI22_X1 U19792 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16768), .ZN(n16754) );
  INV_X1 U19793 ( .A(n16754), .ZN(U265) );
  OAI22_X1 U19794 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16772), .ZN(n16755) );
  INV_X1 U19795 ( .A(n16755), .ZN(U266) );
  OAI22_X1 U19796 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16772), .ZN(n16756) );
  INV_X1 U19797 ( .A(n16756), .ZN(U267) );
  OAI22_X1 U19798 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16772), .ZN(n16757) );
  INV_X1 U19799 ( .A(n16757), .ZN(U268) );
  OAI22_X1 U19800 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16772), .ZN(n16758) );
  INV_X1 U19801 ( .A(n16758), .ZN(U269) );
  OAI22_X1 U19802 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16772), .ZN(n16759) );
  INV_X1 U19803 ( .A(n16759), .ZN(U270) );
  OAI22_X1 U19804 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16772), .ZN(n16760) );
  INV_X1 U19805 ( .A(n16760), .ZN(U271) );
  OAI22_X1 U19806 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16772), .ZN(n16761) );
  INV_X1 U19807 ( .A(n16761), .ZN(U272) );
  INV_X1 U19808 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n16762) );
  INV_X1 U19809 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n18504) );
  AOI22_X1 U19810 ( .A1(n16772), .A2(n16762), .B1(n18504), .B2(U215), .ZN(U273) );
  OAI22_X1 U19811 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16772), .ZN(n16763) );
  INV_X1 U19812 ( .A(n16763), .ZN(U274) );
  INV_X1 U19813 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n16764) );
  AOI22_X1 U19814 ( .A1(n16772), .A2(n16764), .B1(n18476), .B2(U215), .ZN(U275) );
  INV_X1 U19815 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n16765) );
  AOI22_X1 U19816 ( .A1(n16768), .A2(n16765), .B1(n18485), .B2(U215), .ZN(U276) );
  INV_X1 U19817 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n16766) );
  INV_X1 U19818 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n19458) );
  AOI22_X1 U19819 ( .A1(n16772), .A2(n16766), .B1(n19458), .B2(U215), .ZN(U277) );
  INV_X1 U19820 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n16767) );
  INV_X1 U19821 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n19463) );
  AOI22_X1 U19822 ( .A1(n16768), .A2(n16767), .B1(n19463), .B2(U215), .ZN(U278) );
  OAI22_X1 U19823 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16772), .ZN(n16769) );
  INV_X1 U19824 ( .A(n16769), .ZN(U279) );
  INV_X1 U19825 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n16770) );
  INV_X1 U19826 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n19472) );
  AOI22_X1 U19827 ( .A1(n16772), .A2(n16770), .B1(n19472), .B2(U215), .ZN(U280) );
  INV_X1 U19828 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n16771) );
  AOI22_X1 U19829 ( .A1(n16772), .A2(n16771), .B1(n17512), .B2(U215), .ZN(U281) );
  INV_X1 U19830 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19482) );
  AOI22_X1 U19831 ( .A1(n16772), .A2(n16774), .B1(n19482), .B2(U215), .ZN(U282) );
  INV_X1 U19832 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16773) );
  AOI222_X1 U19833 ( .A1(n16775), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16774), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16773), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16776) );
  INV_X2 U19834 ( .A(n16778), .ZN(n16777) );
  INV_X1 U19835 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19029) );
  INV_X1 U19836 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20008) );
  AOI22_X1 U19837 ( .A1(n16777), .A2(n19029), .B1(n20008), .B2(n16778), .ZN(
        U347) );
  INV_X1 U19838 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19027) );
  INV_X1 U19839 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20007) );
  AOI22_X1 U19840 ( .A1(n16777), .A2(n19027), .B1(n20007), .B2(n16778), .ZN(
        U348) );
  INV_X1 U19841 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19025) );
  INV_X1 U19842 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20006) );
  AOI22_X1 U19843 ( .A1(n16777), .A2(n19025), .B1(n20006), .B2(n16778), .ZN(
        U349) );
  INV_X1 U19844 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19023) );
  INV_X1 U19845 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20005) );
  AOI22_X1 U19846 ( .A1(n16777), .A2(n19023), .B1(n20005), .B2(n16778), .ZN(
        U350) );
  INV_X1 U19847 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19021) );
  INV_X1 U19848 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20004) );
  AOI22_X1 U19849 ( .A1(n16777), .A2(n19021), .B1(n20004), .B2(n16778), .ZN(
        U351) );
  INV_X1 U19850 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19018) );
  INV_X1 U19851 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20003) );
  AOI22_X1 U19852 ( .A1(n16777), .A2(n19018), .B1(n20003), .B2(n16778), .ZN(
        U352) );
  INV_X1 U19853 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19017) );
  INV_X1 U19854 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20002) );
  AOI22_X1 U19855 ( .A1(n16777), .A2(n19017), .B1(n20002), .B2(n16778), .ZN(
        U353) );
  INV_X1 U19856 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19015) );
  AOI22_X1 U19857 ( .A1(n16777), .A2(n19015), .B1(n20001), .B2(n16778), .ZN(
        U354) );
  INV_X1 U19858 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19067) );
  INV_X1 U19859 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20039) );
  AOI22_X1 U19860 ( .A1(n16777), .A2(n19067), .B1(n20039), .B2(n16778), .ZN(
        U356) );
  INV_X1 U19861 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19064) );
  INV_X1 U19862 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20037) );
  AOI22_X1 U19863 ( .A1(n16777), .A2(n19064), .B1(n20037), .B2(n16778), .ZN(
        U357) );
  INV_X1 U19864 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19063) );
  INV_X1 U19865 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20035) );
  AOI22_X1 U19866 ( .A1(n16777), .A2(n19063), .B1(n20035), .B2(n16778), .ZN(
        U358) );
  INV_X1 U19867 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19061) );
  INV_X1 U19868 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20033) );
  AOI22_X1 U19869 ( .A1(n16777), .A2(n19061), .B1(n20033), .B2(n16778), .ZN(
        U359) );
  INV_X1 U19870 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19059) );
  INV_X1 U19871 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20031) );
  AOI22_X1 U19872 ( .A1(n16777), .A2(n19059), .B1(n20031), .B2(n16778), .ZN(
        U360) );
  INV_X1 U19873 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19057) );
  INV_X1 U19874 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20029) );
  AOI22_X1 U19875 ( .A1(n16777), .A2(n19057), .B1(n20029), .B2(n16778), .ZN(
        U361) );
  INV_X1 U19876 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19054) );
  INV_X1 U19877 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20027) );
  AOI22_X1 U19878 ( .A1(n16777), .A2(n19054), .B1(n20027), .B2(n16778), .ZN(
        U362) );
  INV_X1 U19879 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19053) );
  INV_X1 U19880 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20025) );
  AOI22_X1 U19881 ( .A1(n16777), .A2(n19053), .B1(n20025), .B2(n16778), .ZN(
        U363) );
  INV_X1 U19882 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19051) );
  INV_X1 U19883 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20023) );
  AOI22_X1 U19884 ( .A1(n16777), .A2(n19051), .B1(n20023), .B2(n16778), .ZN(
        U364) );
  INV_X1 U19885 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19013) );
  INV_X1 U19886 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19999) );
  AOI22_X1 U19887 ( .A1(n16777), .A2(n19013), .B1(n19999), .B2(n16778), .ZN(
        U365) );
  INV_X1 U19888 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19049) );
  INV_X1 U19889 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20021) );
  AOI22_X1 U19890 ( .A1(n16777), .A2(n19049), .B1(n20021), .B2(n16778), .ZN(
        U366) );
  INV_X1 U19891 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19047) );
  INV_X1 U19892 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20019) );
  AOI22_X1 U19893 ( .A1(n16777), .A2(n19047), .B1(n20019), .B2(n16778), .ZN(
        U367) );
  INV_X1 U19894 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19045) );
  INV_X1 U19895 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20018) );
  AOI22_X1 U19896 ( .A1(n16777), .A2(n19045), .B1(n20018), .B2(n16778), .ZN(
        U368) );
  INV_X1 U19897 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19042) );
  INV_X1 U19898 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20016) );
  AOI22_X1 U19899 ( .A1(n16777), .A2(n19042), .B1(n20016), .B2(n16778), .ZN(
        U369) );
  INV_X1 U19900 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19041) );
  INV_X1 U19901 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20015) );
  AOI22_X1 U19902 ( .A1(n16777), .A2(n19041), .B1(n20015), .B2(n16778), .ZN(
        U370) );
  INV_X1 U19903 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19039) );
  INV_X1 U19904 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20014) );
  AOI22_X1 U19905 ( .A1(n16777), .A2(n19039), .B1(n20014), .B2(n16778), .ZN(
        U371) );
  INV_X1 U19906 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19036) );
  INV_X1 U19907 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20013) );
  AOI22_X1 U19908 ( .A1(n16777), .A2(n19036), .B1(n20013), .B2(n16778), .ZN(
        U372) );
  INV_X1 U19909 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19035) );
  INV_X1 U19910 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20012) );
  AOI22_X1 U19911 ( .A1(n16777), .A2(n19035), .B1(n20012), .B2(n16778), .ZN(
        U373) );
  INV_X1 U19912 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19033) );
  INV_X1 U19913 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20010) );
  AOI22_X1 U19914 ( .A1(n16777), .A2(n19033), .B1(n20010), .B2(n16778), .ZN(
        U374) );
  INV_X1 U19915 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19031) );
  INV_X1 U19916 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20009) );
  AOI22_X1 U19917 ( .A1(n16777), .A2(n19031), .B1(n20009), .B2(n16778), .ZN(
        U375) );
  INV_X1 U19918 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19010) );
  INV_X1 U19919 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19998) );
  AOI22_X1 U19920 ( .A1(n16777), .A2(n19010), .B1(n19998), .B2(n16778), .ZN(
        U376) );
  INV_X1 U19921 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16779) );
  NAND2_X1 U19922 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n19009), .ZN(n18996) );
  AOI22_X1 U19923 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18996), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n19007), .ZN(n19083) );
  OAI21_X1 U19924 ( .B1(n19007), .B2(n16779), .A(n19080), .ZN(P3_U2633) );
  OAI21_X1 U19925 ( .B1(n16786), .B2(n17699), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16781) );
  OAI21_X1 U19926 ( .B1(n16782), .B2(n16802), .A(n16781), .ZN(P3_U2634) );
  AOI21_X1 U19927 ( .B1(n19007), .B2(n19009), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16783) );
  AOI22_X1 U19928 ( .A1(n19127), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16783), 
        .B2(n19144), .ZN(P3_U2635) );
  INV_X1 U19929 ( .A(BS16), .ZN(n20920) );
  AOI21_X1 U19930 ( .B1(n16784), .B2(n20920), .A(n19080), .ZN(n19079) );
  INV_X1 U19931 ( .A(n19079), .ZN(n19081) );
  OAI21_X1 U19932 ( .B1(n19083), .B2(n19135), .A(n19081), .ZN(P3_U2636) );
  NOR3_X1 U19933 ( .A1(n16786), .A2(n16785), .A3(n18917), .ZN(n18923) );
  NOR2_X1 U19934 ( .A1(n18923), .A2(n18983), .ZN(n19128) );
  OAI21_X1 U19935 ( .B1(n19128), .B2(n18470), .A(n16787), .ZN(P3_U2637) );
  NOR4_X1 U19936 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16791) );
  NOR4_X1 U19937 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16790) );
  NOR4_X1 U19938 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16789) );
  NOR4_X1 U19939 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16788) );
  NAND4_X1 U19940 ( .A1(n16791), .A2(n16790), .A3(n16789), .A4(n16788), .ZN(
        n16797) );
  NOR4_X1 U19941 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16795) );
  AOI211_X1 U19942 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16794) );
  NOR4_X1 U19943 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16793) );
  NOR4_X1 U19944 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16792) );
  NAND4_X1 U19945 ( .A1(n16795), .A2(n16794), .A3(n16793), .A4(n16792), .ZN(
        n16796) );
  NOR2_X1 U19946 ( .A1(n16797), .A2(n16796), .ZN(n19125) );
  INV_X1 U19947 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19077) );
  NOR3_X1 U19948 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16799) );
  OAI21_X1 U19949 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16799), .A(n19125), .ZN(
        n16798) );
  OAI21_X1 U19950 ( .B1(n19125), .B2(n19077), .A(n16798), .ZN(P3_U2638) );
  INV_X1 U19951 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19074) );
  NOR2_X1 U19952 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19119) );
  OAI21_X1 U19953 ( .B1(n16799), .B2(n19119), .A(n19125), .ZN(n16800) );
  OAI21_X1 U19954 ( .B1(n19125), .B2(n19074), .A(n16800), .ZN(P3_U2639) );
  NOR3_X1 U19955 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .ZN(n18991) );
  INV_X1 U19956 ( .A(n17137), .ZN(n16801) );
  INV_X1 U19957 ( .A(n16802), .ZN(n18145) );
  NOR2_X2 U19958 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n19086), .ZN(n18852) );
  NAND2_X1 U19959 ( .A1(n18145), .A2(n18852), .ZN(n18979) );
  OAI211_X1 U19960 ( .C1(n16803), .C2(n16806), .A(n19137), .B(n19135), .ZN(
        n16804) );
  INV_X1 U19961 ( .A(n16804), .ZN(n18975) );
  NAND2_X1 U19962 ( .A1(n17130), .A2(n17661), .ZN(n16808) );
  AOI211_X4 U19963 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n16806), .A(n18975), .B(
        n16808), .ZN(n17196) );
  INV_X1 U19964 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19071) );
  INV_X1 U19965 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19062) );
  INV_X1 U19966 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19060) );
  INV_X1 U19967 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19056) );
  INV_X1 U19968 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n19052) );
  INV_X1 U19969 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19048) );
  INV_X1 U19970 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19032) );
  INV_X1 U19971 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19028) );
  INV_X1 U19972 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n19019) );
  INV_X1 U19973 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19016) );
  NAND2_X1 U19974 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17167) );
  INV_X1 U19975 ( .A(n17167), .ZN(n17144) );
  NAND2_X1 U19976 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n17144), .ZN(n17136) );
  NOR3_X1 U19977 ( .A1(n19019), .A2(n19016), .A3(n17136), .ZN(n17096) );
  INV_X1 U19978 ( .A(n17096), .ZN(n17058) );
  NAND3_X1 U19979 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(P3_REIP_REG_7__SCAN_IN), 
        .A3(P3_REIP_REG_6__SCAN_IN), .ZN(n17059) );
  NOR2_X1 U19980 ( .A1(n17058), .A2(n17059), .ZN(n17060) );
  NAND2_X1 U19981 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n17060), .ZN(n17056) );
  NOR2_X1 U19982 ( .A1(n19028), .A2(n17056), .ZN(n17043) );
  NAND2_X1 U19983 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n17043), .ZN(n17037) );
  NOR2_X1 U19984 ( .A1(n19032), .A2(n17037), .ZN(n17013) );
  NAND3_X1 U19985 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .A3(n17013), .ZN(n16998) );
  NAND2_X1 U19986 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16986) );
  NOR2_X1 U19987 ( .A1(n16998), .A2(n16986), .ZN(n16976) );
  NAND2_X1 U19988 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n16976), .ZN(n16954) );
  NAND2_X1 U19989 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n16955) );
  NOR3_X1 U19990 ( .A1(n19048), .A2(n16954), .A3(n16955), .ZN(n16918) );
  NAND2_X1 U19991 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n16918), .ZN(n16921) );
  NOR2_X1 U19992 ( .A1(n19052), .A2(n16921), .ZN(n16915) );
  NAND2_X1 U19993 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16915), .ZN(n16884) );
  NOR2_X1 U19994 ( .A1(n19056), .A2(n16884), .ZN(n16891) );
  NAND2_X1 U19995 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16891), .ZN(n16883) );
  NOR2_X1 U19996 ( .A1(n19060), .A2(n16883), .ZN(n16824) );
  NAND2_X1 U19997 ( .A1(n17168), .A2(n16824), .ZN(n16867) );
  NOR3_X1 U19998 ( .A1(n19065), .A2(n19062), .A3(n16867), .ZN(n16848) );
  NAND2_X1 U19999 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16848), .ZN(n16826) );
  NOR3_X1 U20000 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n19071), .A3(n16826), 
        .ZN(n16805) );
  AOI21_X1 U20001 ( .B1(n17196), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16805), .ZN(
        n16831) );
  NAND2_X1 U20002 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n16806), .ZN(n16807) );
  AOI211_X4 U20003 ( .C1(n19135), .C2(n19137), .A(n16808), .B(n16807), .ZN(
        n17195) );
  NOR3_X1 U20004 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17169) );
  INV_X1 U20005 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17152) );
  NAND2_X1 U20006 ( .A1(n17169), .A2(n17152), .ZN(n17151) );
  NOR2_X1 U20007 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17151), .ZN(n17129) );
  NAND2_X1 U20008 ( .A1(n17129), .A2(n17474), .ZN(n17124) );
  NAND2_X1 U20009 ( .A1(n17106), .A2(n17102), .ZN(n17099) );
  INV_X1 U20010 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17078) );
  NAND2_X1 U20011 ( .A1(n17086), .A2(n17078), .ZN(n17077) );
  INV_X1 U20012 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17052) );
  NAND2_X1 U20013 ( .A1(n17061), .A2(n17052), .ZN(n17051) );
  INV_X1 U20014 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17027) );
  NAND2_X1 U20015 ( .A1(n17032), .A2(n17027), .ZN(n17026) );
  INV_X1 U20016 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16996) );
  NAND2_X1 U20017 ( .A1(n17006), .A2(n16996), .ZN(n16994) );
  NAND2_X1 U20018 ( .A1(n16984), .A2(n17345), .ZN(n16981) );
  NAND2_X1 U20019 ( .A1(n16959), .A2(n16953), .ZN(n16952) );
  INV_X1 U20020 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17291) );
  NAND2_X1 U20021 ( .A1(n16939), .A2(n17291), .ZN(n16930) );
  INV_X1 U20022 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16906) );
  NAND2_X1 U20023 ( .A1(n16919), .A2(n16906), .ZN(n16913) );
  INV_X1 U20024 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17247) );
  NAND2_X1 U20025 ( .A1(n16898), .A2(n17247), .ZN(n16890) );
  NAND2_X1 U20026 ( .A1(n16874), .A2(n17244), .ZN(n16870) );
  NOR2_X1 U20027 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16870), .ZN(n16856) );
  INV_X1 U20028 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16851) );
  NAND2_X1 U20029 ( .A1(n16856), .A2(n16851), .ZN(n16833) );
  NOR2_X1 U20030 ( .A1(n17188), .A2(n16833), .ZN(n16840) );
  INV_X1 U20031 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17205) );
  OAI21_X1 U20032 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16820), .A(
        n16809), .ZN(n17786) );
  INV_X1 U20033 ( .A(n17786), .ZN(n16858) );
  OAI21_X1 U20034 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17769), .A(
        n16821), .ZN(n17803) );
  INV_X1 U20035 ( .A(n17803), .ZN(n16876) );
  INV_X1 U20036 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16905) );
  NOR2_X1 U20037 ( .A1(n16905), .A2(n16816), .ZN(n16819) );
  AOI21_X1 U20038 ( .B1(n16905), .B2(n16816), .A(n16819), .ZN(n17824) );
  INV_X1 U20039 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17855) );
  NAND2_X1 U20040 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17882), .ZN(
        n16946) );
  NAND2_X1 U20041 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17850), .ZN(
        n16813) );
  INV_X1 U20042 ( .A(n16813), .ZN(n16814) );
  NAND2_X1 U20043 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16814), .ZN(
        n16810) );
  NOR2_X1 U20044 ( .A1(n17853), .A2(n16813), .ZN(n17812) );
  AOI21_X1 U20045 ( .B1(n17855), .B2(n16810), .A(n17812), .ZN(n17858) );
  OAI21_X1 U20046 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17850), .A(
        n16813), .ZN(n16811) );
  INV_X1 U20047 ( .A(n16811), .ZN(n17886) );
  INV_X1 U20048 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17191) );
  AND2_X1 U20049 ( .A1(n17850), .A2(n17191), .ZN(n16812) );
  NOR2_X1 U20050 ( .A1(n17886), .A2(n16937), .ZN(n16938) );
  INV_X1 U20051 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17872) );
  AOI22_X1 U20052 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16814), .B1(
        n16813), .B2(n17872), .ZN(n17868) );
  INV_X1 U20053 ( .A(n17868), .ZN(n16815) );
  OR2_X1 U20054 ( .A1(n16920), .A2(n9985), .ZN(n16908) );
  OAI21_X1 U20055 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17812), .A(
        n16816), .ZN(n16817) );
  INV_X1 U20056 ( .A(n16817), .ZN(n17847) );
  NOR2_X1 U20057 ( .A1(n16909), .A2(n17146), .ZN(n16900) );
  NOR2_X1 U20058 ( .A1(n17824), .A2(n16900), .ZN(n16899) );
  OR2_X1 U20059 ( .A1(n16899), .A2(n17146), .ZN(n16885) );
  INV_X1 U20060 ( .A(n17769), .ZN(n16818) );
  OAI21_X1 U20061 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16819), .A(
        n16818), .ZN(n17816) );
  INV_X1 U20062 ( .A(n17816), .ZN(n16888) );
  AOI21_X1 U20063 ( .B1(n17773), .B2(n16821), .A(n16820), .ZN(n17787) );
  INV_X1 U20064 ( .A(n16844), .ZN(n16823) );
  NOR2_X1 U20065 ( .A1(n16843), .A2(n9985), .ZN(n16834) );
  NAND2_X1 U20066 ( .A1(n17133), .A2(n16801), .ZN(n17181) );
  NOR3_X1 U20067 ( .A1(n16835), .A2(n16834), .A3(n17181), .ZN(n16829) );
  INV_X1 U20068 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19066) );
  NAND2_X1 U20069 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16825) );
  OR2_X1 U20070 ( .A1(n17190), .A2(n16824), .ZN(n16882) );
  NAND2_X1 U20071 ( .A1(n17189), .A2(n16882), .ZN(n16879) );
  AOI221_X1 U20072 ( .B1(n19066), .B2(n17168), .C1(n16825), .C2(n17168), .A(
        n16879), .ZN(n16854) );
  NOR2_X1 U20073 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16826), .ZN(n16838) );
  INV_X1 U20074 ( .A(n16838), .ZN(n16827) );
  AOI21_X1 U20075 ( .B1(n16854), .B2(n16827), .A(n19069), .ZN(n16828) );
  AOI211_X1 U20076 ( .C1(n16840), .C2(n17205), .A(n16829), .B(n16828), .ZN(
        n16830) );
  OAI211_X1 U20077 ( .C1(n16832), .C2(n17180), .A(n16831), .B(n16830), .ZN(
        P3_U2640) );
  NAND2_X1 U20078 ( .A1(n17195), .A2(n16833), .ZN(n16849) );
  XOR2_X1 U20079 ( .A(n16835), .B(n16834), .Z(n16839) );
  OAI22_X1 U20080 ( .A1(n16854), .A2(n19071), .B1(n16836), .B2(n17180), .ZN(
        n16837) );
  AOI211_X1 U20081 ( .C1(n16839), .C2(n16801), .A(n16838), .B(n16837), .ZN(
        n16842) );
  OAI21_X1 U20082 ( .B1(n17196), .B2(n16840), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16841) );
  AOI211_X1 U20083 ( .C1(n16844), .C2(n9772), .A(n16843), .B(n17137), .ZN(
        n16847) );
  OAI22_X1 U20084 ( .A1(n16845), .A2(n17180), .B1(n17182), .B2(n16851), .ZN(
        n16846) );
  AOI211_X1 U20085 ( .C1(n16848), .C2(n19066), .A(n16847), .B(n16846), .ZN(
        n16853) );
  INV_X1 U20086 ( .A(n16849), .ZN(n16850) );
  OAI21_X1 U20087 ( .B1(n16856), .B2(n16851), .A(n16850), .ZN(n16852) );
  OAI211_X1 U20088 ( .C1(n16854), .C2(n19066), .A(n16853), .B(n16852), .ZN(
        P3_U2642) );
  INV_X1 U20089 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17772) );
  NOR3_X1 U20090 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n19062), .A3(n16867), 
        .ZN(n16855) );
  AOI21_X1 U20091 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17196), .A(n16855), .ZN(
        n16863) );
  INV_X1 U20092 ( .A(n16879), .ZN(n16873) );
  OAI21_X1 U20093 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n16867), .A(n16873), 
        .ZN(n16861) );
  AOI211_X1 U20094 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16870), .A(n16856), .B(
        n17188), .ZN(n16860) );
  AOI211_X1 U20095 ( .C1(n16858), .C2(n16857), .A(n9790), .B(n17137), .ZN(
        n16859) );
  AOI211_X1 U20096 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16861), .A(n16860), 
        .B(n16859), .ZN(n16862) );
  OAI211_X1 U20097 ( .C1(n17772), .C2(n17180), .A(n16863), .B(n16862), .ZN(
        P3_U2643) );
  INV_X1 U20098 ( .A(n16864), .ZN(n16866) );
  AOI211_X1 U20099 ( .C1(n17787), .C2(n16866), .A(n16865), .B(n17137), .ZN(
        n16869) );
  OAI22_X1 U20100 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16867), .B1(n17773), 
        .B2(n17180), .ZN(n16868) );
  AOI211_X1 U20101 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n17196), .A(n16869), .B(
        n16868), .ZN(n16872) );
  OAI211_X1 U20102 ( .C1(n16874), .C2(n17244), .A(n17195), .B(n16870), .ZN(
        n16871) );
  OAI211_X1 U20103 ( .C1(n16873), .C2(n19062), .A(n16872), .B(n16871), .ZN(
        P3_U2644) );
  AOI22_X1 U20104 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17145), .B1(
        n17196), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16881) );
  AOI211_X1 U20105 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16890), .A(n16874), .B(
        n17188), .ZN(n16878) );
  AOI211_X1 U20106 ( .C1(n16876), .C2(n9773), .A(n16875), .B(n17137), .ZN(
        n16877) );
  AOI211_X1 U20107 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n16879), .A(n16878), 
        .B(n16877), .ZN(n16880) );
  OAI211_X1 U20108 ( .C1(n16883), .C2(n16882), .A(n16881), .B(n16880), .ZN(
        P3_U2645) );
  AOI22_X1 U20109 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17145), .B1(
        n17196), .B2(P3_EBX_REG_25__SCAN_IN), .ZN(n16895) );
  NOR2_X1 U20110 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17190), .ZN(n16896) );
  INV_X1 U20111 ( .A(n16884), .ZN(n16897) );
  OAI21_X1 U20112 ( .B1(n16897), .B2(n17190), .A(n17189), .ZN(n16914) );
  INV_X1 U20113 ( .A(n16885), .ZN(n16887) );
  AOI211_X1 U20114 ( .C1(n16888), .C2(n16887), .A(n16886), .B(n17137), .ZN(
        n16889) );
  AOI221_X1 U20115 ( .B1(n16896), .B2(P3_REIP_REG_25__SCAN_IN), .C1(n16914), 
        .C2(P3_REIP_REG_25__SCAN_IN), .A(n16889), .ZN(n16894) );
  OAI211_X1 U20116 ( .C1(n16898), .C2(n17247), .A(n17195), .B(n16890), .ZN(
        n16893) );
  INV_X1 U20117 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19058) );
  NAND3_X1 U20118 ( .A1(n17168), .A2(n16891), .A3(n19058), .ZN(n16892) );
  NAND4_X1 U20119 ( .A1(n16895), .A2(n16894), .A3(n16893), .A4(n16892), .ZN(
        P3_U2646) );
  AOI22_X1 U20120 ( .A1(n17196), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16897), 
        .B2(n16896), .ZN(n16904) );
  AOI211_X1 U20121 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16913), .A(n16898), .B(
        n17188), .ZN(n16902) );
  AOI211_X1 U20122 ( .C1(n17824), .C2(n16900), .A(n16899), .B(n17137), .ZN(
        n16901) );
  AOI211_X1 U20123 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16914), .A(n16902), 
        .B(n16901), .ZN(n16903) );
  OAI211_X1 U20124 ( .C1(n16905), .C2(n17180), .A(n16904), .B(n16903), .ZN(
        P3_U2647) );
  NOR2_X1 U20125 ( .A1(n16919), .A2(n16906), .ZN(n16907) );
  OAI22_X1 U20126 ( .A1(n17188), .A2(n16907), .B1(n17182), .B2(n16906), .ZN(
        n16912) );
  INV_X1 U20127 ( .A(n16908), .ZN(n16910) );
  AOI211_X1 U20128 ( .C1(n17847), .C2(n16910), .A(n16909), .B(n17137), .ZN(
        n16911) );
  AOI21_X1 U20129 ( .B1(n16913), .B2(n16912), .A(n16911), .ZN(n16917) );
  OAI221_X1 U20130 ( .B1(P3_REIP_REG_23__SCAN_IN), .B2(n17168), .C1(
        P3_REIP_REG_23__SCAN_IN), .C2(n16915), .A(n16914), .ZN(n16916) );
  OAI211_X1 U20131 ( .C1(n17180), .C2(n17839), .A(n16917), .B(n16916), .ZN(
        P3_U2648) );
  OAI21_X1 U20132 ( .B1(n17190), .B2(n16918), .A(n17189), .ZN(n16934) );
  INV_X1 U20133 ( .A(n16934), .ZN(n16945) );
  INV_X1 U20134 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19050) );
  NAND3_X1 U20135 ( .A1(n17168), .A2(n16918), .A3(n19050), .ZN(n16935) );
  AOI211_X1 U20136 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16930), .A(n16919), .B(
        n17188), .ZN(n16925) );
  AOI211_X1 U20137 ( .C1(n17858), .C2(n9814), .A(n16920), .B(n17137), .ZN(
        n16924) );
  NOR3_X1 U20138 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n17190), .A3(n16921), 
        .ZN(n16923) );
  OAI22_X1 U20139 ( .A1(n17855), .A2(n17180), .B1(n17182), .B2(n17199), .ZN(
        n16922) );
  NOR4_X1 U20140 ( .A1(n16925), .A2(n16924), .A3(n16923), .A4(n16922), .ZN(
        n16926) );
  OAI221_X1 U20141 ( .B1(n19052), .B2(n16945), .C1(n19052), .C2(n16935), .A(
        n16926), .ZN(P3_U2649) );
  INV_X1 U20142 ( .A(n16927), .ZN(n16929) );
  AOI211_X1 U20143 ( .C1(n17868), .C2(n16929), .A(n16928), .B(n17137), .ZN(
        n16933) );
  OAI211_X1 U20144 ( .C1(n16939), .C2(n17291), .A(n17195), .B(n16930), .ZN(
        n16931) );
  OAI21_X1 U20145 ( .B1(n17180), .B2(n17872), .A(n16931), .ZN(n16932) );
  AOI211_X1 U20146 ( .C1(n16934), .C2(P3_REIP_REG_21__SCAN_IN), .A(n16933), 
        .B(n16932), .ZN(n16936) );
  OAI211_X1 U20147 ( .C1(n17291), .C2(n17182), .A(n16936), .B(n16935), .ZN(
        P3_U2650) );
  AOI22_X1 U20148 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17145), .B1(
        n17196), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n16944) );
  AOI211_X1 U20149 ( .C1(n17886), .C2(n16937), .A(n16938), .B(n17137), .ZN(
        n16942) );
  NOR4_X1 U20150 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n17190), .A3(n16954), 
        .A4(n16955), .ZN(n16941) );
  AOI211_X1 U20151 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16952), .A(n16939), .B(
        n17188), .ZN(n16940) );
  NOR3_X1 U20152 ( .A1(n16942), .A2(n16941), .A3(n16940), .ZN(n16943) );
  OAI211_X1 U20153 ( .C1(n19048), .C2(n16945), .A(n16944), .B(n16943), .ZN(
        P3_U2651) );
  NAND2_X1 U20154 ( .A1(n17168), .A2(n16954), .ZN(n16974) );
  NAND2_X1 U20155 ( .A1(n17189), .A2(n16974), .ZN(n16980) );
  INV_X1 U20156 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17912) );
  NOR2_X1 U20157 ( .A1(n18139), .A2(n17893), .ZN(n17892) );
  INV_X1 U20158 ( .A(n17892), .ZN(n16969) );
  NOR2_X1 U20159 ( .A1(n17912), .A2(n16969), .ZN(n16963) );
  OAI21_X1 U20160 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16963), .A(
        n16946), .ZN(n17897) );
  INV_X1 U20161 ( .A(n17897), .ZN(n16948) );
  INV_X1 U20162 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17946) );
  NAND3_X1 U20163 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17964), .A3(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17009) );
  NOR2_X1 U20164 ( .A1(n17946), .A2(n17009), .ZN(n16972) );
  INV_X1 U20165 ( .A(n16972), .ZN(n16993) );
  OAI21_X1 U20166 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16993), .A(
        n17133), .ZN(n16999) );
  OAI21_X1 U20167 ( .B1(n16963), .B2(n17146), .A(n16999), .ZN(n16964) );
  INV_X1 U20168 ( .A(n16937), .ZN(n16947) );
  AOI221_X1 U20169 ( .B1(n16948), .B2(n16964), .C1(n17897), .C2(n16947), .A(
        n17137), .ZN(n16951) );
  AOI22_X1 U20170 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17145), .B1(
        n17196), .B2(P3_EBX_REG_19__SCAN_IN), .ZN(n16949) );
  INV_X1 U20171 ( .A(n16949), .ZN(n16950) );
  AOI211_X1 U20172 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(n16980), .A(n16951), 
        .B(n16950), .ZN(n16958) );
  OAI211_X1 U20173 ( .C1(n16959), .C2(n16953), .A(n17195), .B(n16952), .ZN(
        n16957) );
  NOR2_X1 U20174 ( .A1(n17190), .A2(n16954), .ZN(n16962) );
  OAI211_X1 U20175 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(P3_REIP_REG_18__SCAN_IN), .A(n16962), .B(n16955), .ZN(n16956) );
  NAND4_X1 U20176 ( .A1(n16958), .A2(n18447), .A3(n16957), .A4(n16956), .ZN(
        P3_U2652) );
  AOI211_X1 U20177 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16981), .A(n16959), .B(
        n17188), .ZN(n16960) );
  AOI21_X1 U20178 ( .B1(n17145), .B2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16960), .ZN(n16968) );
  INV_X1 U20179 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19044) );
  INV_X1 U20180 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17331) );
  OAI21_X1 U20181 ( .B1(n17182), .B2(n17331), .A(n18447), .ZN(n16961) );
  AOI221_X1 U20182 ( .B1(n16962), .B2(n19044), .C1(n16980), .C2(
        P3_REIP_REG_18__SCAN_IN), .A(n16961), .ZN(n16967) );
  NOR2_X1 U20183 ( .A1(n17133), .A2(n17137), .ZN(n17068) );
  AOI21_X1 U20184 ( .B1(n17912), .B2(n16969), .A(n16963), .ZN(n17908) );
  AOI221_X1 U20185 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17908), .C1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n17908), .A(n17137), .ZN(n16965) );
  OAI22_X1 U20186 ( .A1(n17068), .A2(n16965), .B1(n17908), .B2(n16964), .ZN(
        n16966) );
  NAND3_X1 U20187 ( .A1(n16968), .A2(n16967), .A3(n16966), .ZN(P3_U2653) );
  NOR2_X1 U20188 ( .A1(n17935), .A2(n17009), .ZN(n16970) );
  OAI21_X1 U20189 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16970), .A(
        n16969), .ZN(n17921) );
  INV_X1 U20190 ( .A(n16970), .ZN(n16971) );
  OAI21_X1 U20191 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16972), .A(
        n16971), .ZN(n17938) );
  NAND2_X1 U20192 ( .A1(n17938), .A2(n16999), .ZN(n16988) );
  NAND2_X1 U20193 ( .A1(n17133), .A2(n16988), .ZN(n16973) );
  XNOR2_X1 U20194 ( .A(n17921), .B(n16973), .ZN(n16978) );
  INV_X1 U20195 ( .A(n16974), .ZN(n16975) );
  AOI22_X1 U20196 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n17145), .B1(
        n16976), .B2(n16975), .ZN(n16977) );
  OAI211_X1 U20197 ( .C1(n17137), .C2(n16978), .A(n16977), .B(n18447), .ZN(
        n16979) );
  AOI21_X1 U20198 ( .B1(P3_REIP_REG_17__SCAN_IN), .B2(n16980), .A(n16979), 
        .ZN(n16983) );
  OAI211_X1 U20199 ( .C1(n16984), .C2(n17345), .A(n17195), .B(n16981), .ZN(
        n16982) );
  OAI211_X1 U20200 ( .C1(n17345), .C2(n17182), .A(n16983), .B(n16982), .ZN(
        P3_U2654) );
  AOI22_X1 U20201 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17145), .B1(
        n17196), .B2(P3_EBX_REG_16__SCAN_IN), .ZN(n16992) );
  INV_X1 U20202 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19040) );
  INV_X1 U20203 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19038) );
  AOI211_X1 U20204 ( .C1(n19040), .C2(n19038), .A(n16998), .B(n17190), .ZN(
        n16987) );
  AOI211_X1 U20205 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16994), .A(n16984), .B(
        n17188), .ZN(n16985) );
  AOI211_X1 U20206 ( .C1(n16987), .C2(n16986), .A(n9652), .B(n16985), .ZN(
        n16991) );
  INV_X1 U20207 ( .A(n16998), .ZN(n17014) );
  OAI21_X1 U20208 ( .B1(n17014), .B2(n17190), .A(n17189), .ZN(n17010) );
  NAND2_X1 U20209 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n17010), .ZN(n16990) );
  OAI211_X1 U20210 ( .C1(n17938), .C2(n16999), .A(n16801), .B(n16988), .ZN(
        n16989) );
  NAND4_X1 U20211 ( .A1(n16992), .A2(n16991), .A3(n16990), .A4(n16989), .ZN(
        P3_U2655) );
  INV_X1 U20212 ( .A(n17009), .ZN(n17933) );
  OAI21_X1 U20213 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17933), .A(
        n16993), .ZN(n17943) );
  AOI21_X1 U20214 ( .B1(n17133), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n17137), .ZN(n17185) );
  OAI21_X1 U20215 ( .B1(n17068), .B2(n17946), .A(n17185), .ZN(n17005) );
  OAI211_X1 U20216 ( .C1(n17006), .C2(n16996), .A(n17195), .B(n16994), .ZN(
        n16995) );
  OAI211_X1 U20217 ( .C1(n17182), .C2(n16996), .A(n18447), .B(n16995), .ZN(
        n16997) );
  AOI21_X1 U20218 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17145), .A(
        n16997), .ZN(n17004) );
  NOR2_X1 U20219 ( .A1(n17190), .A2(n16998), .ZN(n17002) );
  INV_X1 U20220 ( .A(n17943), .ZN(n17000) );
  NOR3_X1 U20221 ( .A1(n17000), .A2(n17137), .A3(n16999), .ZN(n17001) );
  AOI221_X1 U20222 ( .B1(n17010), .B2(P3_REIP_REG_15__SCAN_IN), .C1(n17002), 
        .C2(n19038), .A(n17001), .ZN(n17003) );
  OAI211_X1 U20223 ( .C1(n17943), .C2(n17005), .A(n17004), .B(n17003), .ZN(
        P3_U2656) );
  AOI211_X1 U20224 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17026), .A(n17006), .B(
        n17188), .ZN(n17008) );
  INV_X1 U20225 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17373) );
  OAI21_X1 U20226 ( .B1(n17182), .B2(n17373), .A(n18447), .ZN(n17007) );
  AOI211_X1 U20227 ( .C1(n17145), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n17008), .B(n17007), .ZN(n17017) );
  NAND2_X1 U20228 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17191), .ZN(
        n17132) );
  NOR3_X1 U20229 ( .A1(n17985), .A2(n17987), .A3(n17132), .ZN(n17012) );
  NOR2_X1 U20230 ( .A1(n17012), .A2(n17181), .ZN(n17021) );
  AND2_X1 U20231 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17964), .ZN(
        n17019) );
  OAI21_X1 U20232 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n17019), .A(
        n17009), .ZN(n17965) );
  AOI22_X1 U20233 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n17010), .B1(n17021), 
        .B2(n17965), .ZN(n17016) );
  INV_X1 U20234 ( .A(n17965), .ZN(n17011) );
  OAI211_X1 U20235 ( .C1(n17012), .C2(n17146), .A(n16801), .B(n17011), .ZN(
        n17015) );
  NAND2_X1 U20236 ( .A1(n17168), .A2(n17013), .ZN(n17022) );
  INV_X1 U20237 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n19034) );
  NAND4_X1 U20238 ( .A1(n17017), .A2(n17016), .A3(n17015), .A4(n10284), .ZN(
        P3_U2657) );
  INV_X1 U20239 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17025) );
  NAND2_X1 U20240 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18046), .ZN(
        n17069) );
  INV_X1 U20241 ( .A(n17069), .ZN(n17109) );
  NAND2_X1 U20242 ( .A1(n17018), .A2(n17109), .ZN(n17045) );
  INV_X1 U20243 ( .A(n17045), .ZN(n17978) );
  NAND2_X1 U20244 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17978), .ZN(
        n17034) );
  AOI21_X1 U20245 ( .B1(n17025), .B2(n17034), .A(n17019), .ZN(n17979) );
  INV_X1 U20246 ( .A(n17979), .ZN(n17020) );
  AOI22_X1 U20247 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17145), .B1(
        n17021), .B2(n17020), .ZN(n17031) );
  INV_X1 U20248 ( .A(n17189), .ZN(n17192) );
  AOI21_X1 U20249 ( .B1(n17168), .B2(n17037), .A(n17192), .ZN(n17048) );
  OAI21_X1 U20250 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n17190), .A(n17048), 
        .ZN(n17024) );
  OAI22_X1 U20251 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n17022), .B1(n17182), 
        .B2(n17027), .ZN(n17023) );
  AOI211_X1 U20252 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n17024), .A(n9652), .B(
        n17023), .ZN(n17030) );
  OAI211_X1 U20253 ( .C1(n17068), .C2(n17025), .A(n17979), .B(n17185), .ZN(
        n17029) );
  OAI211_X1 U20254 ( .C1(n17032), .C2(n17027), .A(n17195), .B(n17026), .ZN(
        n17028) );
  NAND4_X1 U20255 ( .A1(n17031), .A2(n17030), .A3(n17029), .A4(n17028), .ZN(
        P3_U2658) );
  AOI211_X1 U20256 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17051), .A(n17032), .B(
        n17188), .ZN(n17033) );
  AOI21_X1 U20257 ( .B1(n17145), .B2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n17033), .ZN(n17042) );
  OAI21_X1 U20258 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17978), .A(
        n17034), .ZN(n17995) );
  OAI21_X1 U20259 ( .B1(n17985), .B2(n17132), .A(n17133), .ZN(n17035) );
  XOR2_X1 U20260 ( .A(n17995), .B(n17035), .Z(n17040) );
  NAND2_X1 U20261 ( .A1(n17168), .A2(n19032), .ZN(n17036) );
  OAI22_X1 U20262 ( .A1(n17182), .A2(n17038), .B1(n17037), .B2(n17036), .ZN(
        n17039) );
  AOI211_X1 U20263 ( .C1(n16801), .C2(n17040), .A(n9652), .B(n17039), .ZN(
        n17041) );
  OAI211_X1 U20264 ( .C1(n19032), .C2(n17048), .A(n17042), .B(n17041), .ZN(
        P3_U2659) );
  AOI21_X1 U20265 ( .B1(n17168), .B2(n17043), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n17049) );
  NOR2_X1 U20266 ( .A1(n18054), .A2(n17069), .ZN(n17083) );
  NAND2_X1 U20267 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17083), .ZN(
        n17067) );
  NOR2_X1 U20268 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17067), .ZN(
        n17044) );
  AOI21_X1 U20269 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17044), .A(
        n17146), .ZN(n17046) );
  NOR2_X1 U20270 ( .A1(n18022), .A2(n17067), .ZN(n17055) );
  OAI21_X1 U20271 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17055), .A(
        n17045), .ZN(n18007) );
  XOR2_X1 U20272 ( .A(n17046), .B(n18007), .Z(n17047) );
  OAI22_X1 U20273 ( .A1(n17049), .A2(n17048), .B1(n17137), .B2(n17047), .ZN(
        n17050) );
  AOI211_X1 U20274 ( .C1(n17196), .C2(P3_EBX_REG_11__SCAN_IN), .A(n9652), .B(
        n17050), .ZN(n17054) );
  OAI211_X1 U20275 ( .C1(n17061), .C2(n17052), .A(n17195), .B(n17051), .ZN(
        n17053) );
  OAI211_X1 U20276 ( .C1(n17180), .C2(n18009), .A(n17054), .B(n17053), .ZN(
        P3_U2660) );
  AOI21_X1 U20277 ( .B1(n18022), .B2(n17067), .A(n17055), .ZN(n18025) );
  OAI21_X1 U20278 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17067), .A(
        n17133), .ZN(n17072) );
  XOR2_X1 U20279 ( .A(n18025), .B(n17072), .Z(n17066) );
  NOR3_X1 U20280 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n17190), .A3(n17056), 
        .ZN(n17057) );
  AOI211_X1 U20281 ( .C1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n17145), .A(
        n9652), .B(n17057), .ZN(n17065) );
  AOI221_X1 U20282 ( .B1(n17059), .B2(n17168), .C1(n17058), .C2(n17168), .A(
        n17192), .ZN(n17091) );
  INV_X1 U20283 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19026) );
  NAND3_X1 U20284 ( .A1(n17168), .A2(n17060), .A3(n19026), .ZN(n17073) );
  AOI21_X1 U20285 ( .B1(n17091), .B2(n17073), .A(n19028), .ZN(n17063) );
  AOI211_X1 U20286 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17077), .A(n17061), .B(
        n17188), .ZN(n17062) );
  AOI211_X1 U20287 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17196), .A(n17063), .B(
        n17062), .ZN(n17064) );
  OAI211_X1 U20288 ( .C1(n17137), .C2(n17066), .A(n17065), .B(n17064), .ZN(
        P3_U2661) );
  INV_X1 U20289 ( .A(n17091), .ZN(n17076) );
  OAI21_X1 U20290 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17083), .A(
        n17067), .ZN(n18037) );
  INV_X1 U20291 ( .A(n17068), .ZN(n17162) );
  INV_X1 U20292 ( .A(n18054), .ZN(n17070) );
  NOR2_X1 U20293 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17069), .ZN(
        n17111) );
  OAI221_X1 U20294 ( .B1(n18037), .B2(n17070), .C1(n18037), .C2(n17111), .A(
        n16801), .ZN(n17071) );
  AOI22_X1 U20295 ( .A1(n18037), .A2(n17072), .B1(n17162), .B2(n17071), .ZN(
        n17075) );
  OAI211_X1 U20296 ( .C1(n17182), .C2(n17078), .A(n18447), .B(n17073), .ZN(
        n17074) );
  AOI211_X1 U20297 ( .C1(n17076), .C2(P3_REIP_REG_9__SCAN_IN), .A(n17075), .B(
        n17074), .ZN(n17080) );
  OAI211_X1 U20298 ( .C1(n17086), .C2(n17078), .A(n17195), .B(n17077), .ZN(
        n17079) );
  OAI211_X1 U20299 ( .C1(n17180), .C2(n17081), .A(n17080), .B(n17079), .ZN(
        P3_U2662) );
  INV_X1 U20300 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19024) );
  INV_X1 U20301 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19022) );
  INV_X1 U20302 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19020) );
  NAND2_X1 U20303 ( .A1(n17168), .A2(n17096), .ZN(n17097) );
  NOR4_X1 U20304 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n19022), .A3(n19020), .A4(
        n17097), .ZN(n17082) );
  AOI211_X1 U20305 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17145), .A(
        n9652), .B(n17082), .ZN(n17090) );
  INV_X1 U20306 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17084) );
  NAND2_X1 U20307 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17109), .ZN(
        n17093) );
  AOI21_X1 U20308 ( .B1(n17084), .B2(n17093), .A(n17083), .ZN(n18047) );
  INV_X1 U20309 ( .A(n18046), .ZN(n18059) );
  INV_X1 U20310 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18061) );
  NOR2_X1 U20311 ( .A1(n18059), .A2(n18061), .ZN(n18055) );
  INV_X1 U20312 ( .A(n17132), .ZN(n17166) );
  AOI21_X1 U20313 ( .B1(n18055), .B2(n17166), .A(n17146), .ZN(n17092) );
  OAI21_X1 U20314 ( .B1(n18047), .B2(n17092), .A(n16801), .ZN(n17085) );
  AOI21_X1 U20315 ( .B1(n18047), .B2(n17092), .A(n17085), .ZN(n17088) );
  AOI211_X1 U20316 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17099), .A(n17086), .B(
        n17188), .ZN(n17087) );
  AOI211_X1 U20317 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17196), .A(n17088), .B(
        n17087), .ZN(n17089) );
  OAI211_X1 U20318 ( .C1(n19024), .C2(n17091), .A(n17090), .B(n17089), .ZN(
        P3_U2663) );
  NOR2_X1 U20319 ( .A1(n17111), .A2(n17146), .ZN(n17095) );
  INV_X1 U20320 ( .A(n17092), .ZN(n17094) );
  OAI21_X1 U20321 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17109), .A(
        n17093), .ZN(n18070) );
  MUX2_X1 U20322 ( .A(n17095), .B(n17094), .S(n18070), .Z(n17105) );
  OAI21_X1 U20323 ( .B1(n17096), .B2(n17190), .A(n17189), .ZN(n17117) );
  NOR2_X1 U20324 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n17097), .ZN(n17113) );
  NOR3_X1 U20325 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n19020), .A3(n17097), .ZN(
        n17098) );
  AOI211_X1 U20326 ( .C1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n17145), .A(
        n9652), .B(n17098), .ZN(n17101) );
  OAI211_X1 U20327 ( .C1(n17106), .C2(n17102), .A(n17195), .B(n17099), .ZN(
        n17100) );
  OAI211_X1 U20328 ( .C1(n17102), .C2(n17182), .A(n17101), .B(n17100), .ZN(
        n17103) );
  AOI221_X1 U20329 ( .B1(n17117), .B2(P3_REIP_REG_7__SCAN_IN), .C1(n17113), 
        .C2(P3_REIP_REG_7__SCAN_IN), .A(n17103), .ZN(n17104) );
  OAI21_X1 U20330 ( .B1(n17137), .B2(n17105), .A(n17104), .ZN(P3_U2664) );
  AOI211_X1 U20331 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17124), .A(n17106), .B(
        n17188), .ZN(n17108) );
  OAI22_X1 U20332 ( .A1(n18082), .A2(n17180), .B1(n17182), .B2(n17469), .ZN(
        n17107) );
  NOR3_X1 U20333 ( .A1(n9652), .A2(n17108), .A3(n17107), .ZN(n17116) );
  NOR2_X1 U20334 ( .A1(n18139), .A2(n18075), .ZN(n17118) );
  INV_X1 U20335 ( .A(n17118), .ZN(n17110) );
  AOI21_X1 U20336 ( .B1(n18082), .B2(n17110), .A(n17109), .ZN(n18079) );
  NOR3_X1 U20337 ( .A1(n18079), .A2(n17111), .A3(n17181), .ZN(n17112) );
  AOI211_X1 U20338 ( .C1(n17117), .C2(P3_REIP_REG_6__SCAN_IN), .A(n17113), .B(
        n17112), .ZN(n17115) );
  OAI211_X1 U20339 ( .C1(n17118), .C2(n17146), .A(n18079), .B(n17185), .ZN(
        n17114) );
  NAND3_X1 U20340 ( .A1(n17116), .A2(n17115), .A3(n17114), .ZN(P3_U2665) );
  INV_X1 U20341 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17127) );
  NOR2_X1 U20342 ( .A1(n17190), .A2(n17136), .ZN(n17128) );
  AOI21_X1 U20343 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n17128), .A(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17122) );
  INV_X1 U20344 ( .A(n17117), .ZN(n17121) );
  NAND2_X1 U20345 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18083), .ZN(
        n17131) );
  AOI21_X1 U20346 ( .B1(n17127), .B2(n17131), .A(n17118), .ZN(n18090) );
  INV_X1 U20347 ( .A(n17131), .ZN(n17119) );
  AOI21_X1 U20348 ( .B1(n17191), .B2(n17119), .A(n17146), .ZN(n17135) );
  XNOR2_X1 U20349 ( .A(n18090), .B(n17135), .ZN(n17120) );
  OAI22_X1 U20350 ( .A1(n17122), .A2(n17121), .B1(n17137), .B2(n17120), .ZN(
        n17123) );
  AOI211_X1 U20351 ( .C1(n17196), .C2(P3_EBX_REG_5__SCAN_IN), .A(n9652), .B(
        n17123), .ZN(n17126) );
  OAI211_X1 U20352 ( .C1(n17129), .C2(n17474), .A(n17195), .B(n17124), .ZN(
        n17125) );
  OAI211_X1 U20353 ( .C1(n17180), .C2(n17127), .A(n17126), .B(n17125), .ZN(
        P3_U2666) );
  AOI22_X1 U20354 ( .A1(n17196), .A2(P3_EBX_REG_4__SCAN_IN), .B1(n17128), .B2(
        n19016), .ZN(n17143) );
  AOI211_X1 U20355 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17151), .A(n17129), .B(
        n17188), .ZN(n17141) );
  NAND2_X1 U20356 ( .A1(n18482), .A2(n17130), .ZN(n19150) );
  AOI21_X1 U20357 ( .B1(n17150), .B2(n18926), .A(n19150), .ZN(n17140) );
  NOR2_X1 U20358 ( .A1(n18139), .A2(n18102), .ZN(n17148) );
  OAI21_X1 U20359 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17148), .A(
        n17131), .ZN(n18105) );
  OR2_X1 U20360 ( .A1(n18102), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18109) );
  OAI22_X1 U20361 ( .A1(n17133), .A2(n18105), .B1(n17132), .B2(n18109), .ZN(
        n17134) );
  AOI21_X1 U20362 ( .B1(n17135), .B2(n18105), .A(n17134), .ZN(n17138) );
  AOI21_X1 U20363 ( .B1(n17168), .B2(n17136), .A(n17192), .ZN(n17158) );
  OAI22_X1 U20364 ( .A1(n17138), .A2(n17137), .B1(n19016), .B2(n17158), .ZN(
        n17139) );
  NOR4_X1 U20365 ( .A1(n9652), .A2(n17141), .A3(n17140), .A4(n17139), .ZN(
        n17142) );
  OAI211_X1 U20366 ( .C1(n18104), .C2(n17180), .A(n17143), .B(n17142), .ZN(
        P3_U2667) );
  AOI21_X1 U20367 ( .B1(n17168), .B2(n17144), .A(P3_REIP_REG_3__SCAN_IN), .ZN(
        n17159) );
  AOI22_X1 U20368 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n17145), .B1(
        n17196), .B2(P3_EBX_REG_3__SCAN_IN), .ZN(n17157) );
  NAND2_X1 U20369 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17161) );
  INV_X1 U20370 ( .A(n17161), .ZN(n17147) );
  AOI21_X1 U20371 ( .B1(n17147), .B2(n17191), .A(n17146), .ZN(n17165) );
  INV_X1 U20372 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17149) );
  AOI21_X1 U20373 ( .B1(n17149), .B2(n17161), .A(n17148), .ZN(n18115) );
  XOR2_X1 U20374 ( .A(n17165), .B(n18115), .Z(n17155) );
  NOR2_X1 U20375 ( .A1(n19102), .A2(n19108), .ZN(n18937) );
  NAND2_X1 U20376 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18937), .ZN(
        n18939) );
  INV_X1 U20377 ( .A(n18939), .ZN(n17160) );
  OAI21_X1 U20378 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n17160), .A(
        n17150), .ZN(n19087) );
  OAI211_X1 U20379 ( .C1(n17169), .C2(n17152), .A(n17195), .B(n17151), .ZN(
        n17153) );
  OAI21_X1 U20380 ( .B1(n19150), .B2(n19087), .A(n17153), .ZN(n17154) );
  AOI21_X1 U20381 ( .B1(n17155), .B2(n16801), .A(n17154), .ZN(n17156) );
  OAI211_X1 U20382 ( .C1(n17159), .C2(n17158), .A(n17157), .B(n17156), .ZN(
        P3_U2668) );
  AOI21_X1 U20383 ( .B1(n9639), .B2(n18944), .A(n17160), .ZN(n19098) );
  INV_X1 U20384 ( .A(n19150), .ZN(n17179) );
  INV_X1 U20385 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18129) );
  INV_X1 U20386 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17171) );
  OAI22_X1 U20387 ( .A1(n18129), .A2(n17180), .B1(n17182), .B2(n17171), .ZN(
        n17164) );
  INV_X1 U20388 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n19012) );
  OAI21_X1 U20389 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n17161), .ZN(n18125) );
  OAI22_X1 U20390 ( .A1(n19012), .A2(n17189), .B1(n18125), .B2(n17162), .ZN(
        n17163) );
  AOI211_X1 U20391 ( .C1(n19098), .C2(n17179), .A(n17164), .B(n17163), .ZN(
        n17176) );
  OAI211_X1 U20392 ( .C1(n17166), .C2(n18125), .A(n16801), .B(n17165), .ZN(
        n17175) );
  OAI211_X1 U20393 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17168), .B(n17167), .ZN(n17174) );
  NOR2_X1 U20394 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17172) );
  INV_X1 U20395 ( .A(n17169), .ZN(n17170) );
  OAI211_X1 U20396 ( .C1(n17172), .C2(n17171), .A(n17195), .B(n17170), .ZN(
        n17173) );
  NAND4_X1 U20397 ( .A1(n17176), .A2(n17175), .A3(n17174), .A4(n17173), .ZN(
        P3_U2669) );
  OAI21_X1 U20398 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n17177), .ZN(n17498) );
  NAND2_X1 U20399 ( .A1(n18944), .A2(n17178), .ZN(n18955) );
  INV_X1 U20400 ( .A(n18955), .ZN(n19105) );
  AOI22_X1 U20401 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17192), .B1(n19105), 
        .B2(n17179), .ZN(n17187) );
  OAI21_X1 U20402 ( .B1(n17191), .B2(n17181), .A(n17180), .ZN(n17184) );
  INV_X1 U20403 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17497) );
  OAI22_X1 U20404 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17190), .B1(n17182), 
        .B2(n17497), .ZN(n17183) );
  AOI221_X1 U20405 ( .B1(n17185), .B2(n18139), .C1(n17184), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n17183), .ZN(n17186) );
  OAI211_X1 U20406 ( .C1(n17188), .C2(n17498), .A(n17187), .B(n17186), .ZN(
        P3_U2670) );
  NAND2_X1 U20407 ( .A1(n17190), .A2(n17189), .ZN(n17194) );
  NOR3_X1 U20408 ( .A1(n19111), .A2(n17192), .A3(n17191), .ZN(n17193) );
  AOI21_X1 U20409 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(n17194), .A(n17193), .ZN(
        n17198) );
  OAI21_X1 U20410 ( .B1(n17196), .B2(n17195), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n17197) );
  OAI211_X1 U20411 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n19150), .A(
        n17198), .B(n17197), .ZN(P3_U2671) );
  NOR3_X1 U20412 ( .A1(n17199), .A2(n17291), .A3(n17290), .ZN(n17200) );
  NAND4_X1 U20413 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17201), .A3(n17232), 
        .A4(n17200), .ZN(n17204) );
  NOR2_X1 U20414 ( .A1(n17205), .A2(n17204), .ZN(n17231) );
  NAND2_X1 U20415 ( .A1(n17494), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17203) );
  NAND2_X1 U20416 ( .A1(n17231), .A2(n18512), .ZN(n17202) );
  OAI22_X1 U20417 ( .A1(n17231), .A2(n17203), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17202), .ZN(P3_U2672) );
  NAND2_X1 U20418 ( .A1(n17205), .A2(n17204), .ZN(n17206) );
  NAND2_X1 U20419 ( .A1(n17206), .A2(n17494), .ZN(n17230) );
  AOI22_X1 U20420 ( .A1(n9656), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17432), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17210) );
  AOI22_X1 U20421 ( .A1(n17380), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17407), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17209) );
  AOI22_X1 U20422 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17208) );
  AOI22_X1 U20423 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17207) );
  NAND4_X1 U20424 ( .A1(n17210), .A2(n17209), .A3(n17208), .A4(n17207), .ZN(
        n17218) );
  AOI22_X1 U20425 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17216) );
  AOI22_X1 U20426 ( .A1(n15929), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17215) );
  AOI22_X1 U20427 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17214) );
  AOI22_X1 U20428 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9658), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17213) );
  NAND4_X1 U20429 ( .A1(n17216), .A2(n17215), .A3(n17214), .A4(n17213), .ZN(
        n17217) );
  NOR2_X1 U20430 ( .A1(n17218), .A2(n17217), .ZN(n17235) );
  NOR2_X1 U20431 ( .A1(n17235), .A2(n17234), .ZN(n17233) );
  AOI22_X1 U20432 ( .A1(n17380), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9656), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17222) );
  AOI22_X1 U20433 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17221) );
  AOI22_X1 U20434 ( .A1(n17456), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17219) );
  NAND4_X1 U20435 ( .A1(n17222), .A2(n17221), .A3(n17220), .A4(n17219), .ZN(
        n17228) );
  AOI22_X1 U20436 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17226) );
  AOI22_X1 U20437 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17225) );
  AOI22_X1 U20438 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17432), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17224) );
  AOI22_X1 U20439 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9658), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17223) );
  NAND4_X1 U20440 ( .A1(n17226), .A2(n17225), .A3(n17224), .A4(n17223), .ZN(
        n17227) );
  NOR2_X1 U20441 ( .A1(n17228), .A2(n17227), .ZN(n17229) );
  XOR2_X1 U20442 ( .A(n17233), .B(n17229), .Z(n17513) );
  OAI22_X1 U20443 ( .A1(n17231), .A2(n17230), .B1(n17513), .B2(n17494), .ZN(
        P3_U2673) );
  NAND2_X1 U20444 ( .A1(n17241), .A2(n17232), .ZN(n17238) );
  AOI21_X1 U20445 ( .B1(n17235), .B2(n17234), .A(n17233), .ZN(n17517) );
  AOI22_X1 U20446 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17236), .B1(n17517), 
        .B2(n17500), .ZN(n17237) );
  OAI21_X1 U20447 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n17238), .A(n17237), .ZN(
        P3_U2674) );
  AOI21_X1 U20448 ( .B1(n17240), .B2(n17245), .A(n17239), .ZN(n17526) );
  AOI22_X1 U20449 ( .A1(n17500), .A2(n17526), .B1(n17241), .B2(n17244), .ZN(
        n17242) );
  OAI21_X1 U20450 ( .B1(n17244), .B2(n17243), .A(n17242), .ZN(P3_U2676) );
  OAI21_X1 U20451 ( .B1(n17252), .B2(n17246), .A(n17245), .ZN(n17534) );
  NAND3_X1 U20452 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(n17261), .ZN(n17251) );
  NOR2_X1 U20453 ( .A1(n17247), .A2(n17251), .ZN(n17256) );
  INV_X1 U20454 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n17248) );
  AOI22_X1 U20455 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17249), .B1(n17256), 
        .B2(n17248), .ZN(n17250) );
  OAI21_X1 U20456 ( .B1(n17534), .B2(n17494), .A(n17250), .ZN(P3_U2677) );
  INV_X1 U20457 ( .A(n17251), .ZN(n17260) );
  AOI21_X1 U20458 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17494), .A(n17260), .ZN(
        n17255) );
  AOI21_X1 U20459 ( .B1(n17253), .B2(n17257), .A(n17252), .ZN(n17535) );
  INV_X1 U20460 ( .A(n17535), .ZN(n17254) );
  OAI22_X1 U20461 ( .A1(n17256), .A2(n17255), .B1(n17254), .B2(n17494), .ZN(
        P3_U2678) );
  AOI22_X1 U20462 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17494), .B1(
        P3_EBX_REG_23__SCAN_IN), .B2(n17261), .ZN(n17259) );
  OAI21_X1 U20463 ( .B1(n17262), .B2(n17258), .A(n17257), .ZN(n17545) );
  OAI22_X1 U20464 ( .A1(n17260), .A2(n17259), .B1(n17545), .B2(n17494), .ZN(
        P3_U2679) );
  AND2_X1 U20465 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n17261), .ZN(n17267) );
  AOI21_X1 U20466 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17494), .A(n17261), .ZN(
        n17266) );
  AOI21_X1 U20467 ( .B1(n17264), .B2(n17263), .A(n17262), .ZN(n17546) );
  INV_X1 U20468 ( .A(n17546), .ZN(n17265) );
  OAI22_X1 U20469 ( .A1(n17267), .A2(n17266), .B1(n17494), .B2(n17265), .ZN(
        P3_U2680) );
  AOI22_X1 U20470 ( .A1(n17380), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17271) );
  AOI22_X1 U20471 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17270) );
  AOI22_X1 U20472 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17269) );
  AOI22_X1 U20473 ( .A1(n17432), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17268) );
  NAND4_X1 U20474 ( .A1(n17271), .A2(n17270), .A3(n17269), .A4(n17268), .ZN(
        n17277) );
  AOI22_X1 U20475 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17275) );
  AOI22_X1 U20476 ( .A1(n9656), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17274) );
  AOI22_X1 U20477 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9658), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17272) );
  NAND4_X1 U20478 ( .A1(n17275), .A2(n17274), .A3(n17273), .A4(n17272), .ZN(
        n17276) );
  NOR2_X1 U20479 ( .A1(n17277), .A2(n17276), .ZN(n17554) );
  NAND3_X1 U20480 ( .A1(n17279), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17494), 
        .ZN(n17278) );
  OAI221_X1 U20481 ( .B1(n17279), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17494), 
        .C2(n17554), .A(n17278), .ZN(P3_U2681) );
  AOI22_X1 U20482 ( .A1(n17380), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9656), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17283) );
  AOI22_X1 U20483 ( .A1(n15929), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17282) );
  AOI22_X1 U20484 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17432), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17281) );
  AOI22_X1 U20485 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13971), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17280) );
  NAND4_X1 U20486 ( .A1(n17283), .A2(n17282), .A3(n17281), .A4(n17280), .ZN(
        n17289) );
  AOI22_X1 U20487 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17287) );
  AOI22_X1 U20488 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17286) );
  AOI22_X1 U20489 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17285) );
  AOI22_X1 U20490 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9658), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17284) );
  NAND4_X1 U20491 ( .A1(n17287), .A2(n17286), .A3(n17285), .A4(n17284), .ZN(
        n17288) );
  NOR2_X1 U20492 ( .A1(n17289), .A2(n17288), .ZN(n17561) );
  AND2_X1 U20493 ( .A1(n17494), .A2(n17290), .ZN(n17304) );
  AOI22_X1 U20494 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17304), .B1(n17292), 
        .B2(n17291), .ZN(n17293) );
  OAI21_X1 U20495 ( .B1(n17561), .B2(n17494), .A(n17293), .ZN(P3_U2682) );
  AOI22_X1 U20496 ( .A1(n17432), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17297) );
  AOI22_X1 U20497 ( .A1(n15864), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9656), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17296) );
  AOI22_X1 U20498 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17295) );
  AOI22_X1 U20499 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17380), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17294) );
  NAND4_X1 U20500 ( .A1(n17297), .A2(n17296), .A3(n17295), .A4(n17294), .ZN(
        n17303) );
  AOI22_X1 U20501 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17301) );
  AOI22_X1 U20502 ( .A1(n17456), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17300) );
  AOI22_X1 U20503 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9658), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17298) );
  NAND4_X1 U20504 ( .A1(n17301), .A2(n17300), .A3(n17299), .A4(n17298), .ZN(
        n17302) );
  NOR2_X1 U20505 ( .A1(n17303), .A2(n17302), .ZN(n17566) );
  OAI21_X1 U20506 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17319), .A(n17304), .ZN(
        n17305) );
  OAI21_X1 U20507 ( .B1(n17566), .B2(n17494), .A(n17305), .ZN(P3_U2683) );
  INV_X1 U20508 ( .A(n17306), .ZN(n17307) );
  OAI21_X1 U20509 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17307), .A(n17494), .ZN(
        n17318) );
  AOI22_X1 U20510 ( .A1(n17432), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13971), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17311) );
  AOI22_X1 U20511 ( .A1(n17380), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17310) );
  AOI22_X1 U20512 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17309) );
  AOI22_X1 U20513 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9656), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17308) );
  NAND4_X1 U20514 ( .A1(n17311), .A2(n17310), .A3(n17309), .A4(n17308), .ZN(
        n17317) );
  AOI22_X1 U20515 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17315) );
  AOI22_X1 U20516 ( .A1(n15864), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17314) );
  AOI22_X1 U20517 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9658), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17312) );
  NAND4_X1 U20518 ( .A1(n17315), .A2(n17314), .A3(n17313), .A4(n17312), .ZN(
        n17316) );
  NOR2_X1 U20519 ( .A1(n17317), .A2(n17316), .ZN(n17571) );
  OAI22_X1 U20520 ( .A1(n17319), .A2(n17318), .B1(n17571), .B2(n17494), .ZN(
        P3_U2684) );
  OR2_X1 U20521 ( .A1(n17331), .A2(n17320), .ZN(n17333) );
  AOI22_X1 U20522 ( .A1(n15864), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17324) );
  AOI22_X1 U20523 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17323) );
  AOI22_X1 U20524 ( .A1(n17380), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17322) );
  NAND4_X1 U20525 ( .A1(n17324), .A2(n17323), .A3(n17322), .A4(n17321), .ZN(
        n17330) );
  AOI22_X1 U20526 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17328) );
  AOI22_X1 U20527 ( .A1(n17432), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17327) );
  AOI22_X1 U20528 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17326) );
  AOI22_X1 U20529 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9658), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17325) );
  NAND4_X1 U20530 ( .A1(n17328), .A2(n17327), .A3(n17326), .A4(n17325), .ZN(
        n17329) );
  NOR2_X1 U20531 ( .A1(n17330), .A2(n17329), .ZN(n17575) );
  NOR2_X1 U20532 ( .A1(n17489), .A2(n17372), .ZN(n17387) );
  NAND3_X1 U20533 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(n17387), .ZN(n17374) );
  INV_X1 U20534 ( .A(n17374), .ZN(n17349) );
  NAND3_X1 U20535 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17361), .A3(n17331), 
        .ZN(n17332) );
  OAI221_X1 U20536 ( .B1(n17500), .B2(n17333), .C1(n17494), .C2(n17575), .A(
        n17332), .ZN(P3_U2685) );
  AOI22_X1 U20537 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n15929), .ZN(n17338) );
  AOI22_X1 U20538 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n17380), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n9655), .ZN(n17337) );
  AOI22_X1 U20539 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n17334), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17447), .ZN(n17336) );
  AOI22_X1 U20540 ( .A1(n15864), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17335) );
  NAND4_X1 U20541 ( .A1(n17338), .A2(n17337), .A3(n17336), .A4(n17335), .ZN(
        n17344) );
  AOI22_X1 U20542 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17342) );
  AOI22_X1 U20543 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17456), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n9656), .ZN(n17341) );
  AOI22_X1 U20544 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17340) );
  AOI22_X1 U20545 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n9667), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n9658), .ZN(n17339) );
  NAND4_X1 U20546 ( .A1(n17342), .A2(n17341), .A3(n17340), .A4(n17339), .ZN(
        n17343) );
  NOR2_X1 U20547 ( .A1(n17344), .A2(n17343), .ZN(n17582) );
  NOR2_X1 U20548 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17361), .ZN(n17348) );
  AOI211_X1 U20549 ( .C1(n18512), .C2(n17346), .A(n17345), .B(n17499), .ZN(
        n17347) );
  OAI22_X1 U20550 ( .A1(n17582), .A2(n17494), .B1(n17348), .B2(n17347), .ZN(
        P3_U2686) );
  AOI21_X1 U20551 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17494), .A(n17349), .ZN(
        n17360) );
  AOI22_X1 U20552 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17353) );
  AOI22_X1 U20553 ( .A1(n15864), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17352) );
  AOI22_X1 U20554 ( .A1(n17432), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17350) );
  NAND4_X1 U20555 ( .A1(n17353), .A2(n17352), .A3(n17351), .A4(n17350), .ZN(
        n17359) );
  AOI22_X1 U20556 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17357) );
  AOI22_X1 U20557 ( .A1(n17380), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17356) );
  AOI22_X1 U20558 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9656), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17355) );
  AOI22_X1 U20559 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9658), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17354) );
  NAND4_X1 U20560 ( .A1(n17357), .A2(n17356), .A3(n17355), .A4(n17354), .ZN(
        n17358) );
  NOR2_X1 U20561 ( .A1(n17359), .A2(n17358), .ZN(n17589) );
  OAI22_X1 U20562 ( .A1(n17361), .A2(n17360), .B1(n17589), .B2(n17494), .ZN(
        P3_U2687) );
  AOI22_X1 U20563 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17365) );
  AOI22_X1 U20564 ( .A1(n15864), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17364) );
  AOI22_X1 U20565 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17362) );
  NAND4_X1 U20566 ( .A1(n17365), .A2(n17364), .A3(n17363), .A4(n17362), .ZN(
        n17371) );
  AOI22_X1 U20567 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17369) );
  AOI22_X1 U20568 ( .A1(n15756), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17368) );
  AOI22_X1 U20569 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17380), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17367) );
  AOI22_X1 U20570 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9658), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17366) );
  NAND4_X1 U20571 ( .A1(n17369), .A2(n17368), .A3(n17367), .A4(n17366), .ZN(
        n17370) );
  NOR2_X1 U20572 ( .A1(n17371), .A2(n17370), .ZN(n17593) );
  NOR2_X1 U20573 ( .A1(n17373), .A2(n17372), .ZN(n17389) );
  OAI21_X1 U20574 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17389), .A(n17374), .ZN(
        n17375) );
  AOI22_X1 U20575 ( .A1(n17500), .A2(n17593), .B1(n17375), .B2(n17494), .ZN(
        P3_U2688) );
  AOI22_X1 U20576 ( .A1(n17432), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17379) );
  AOI22_X1 U20577 ( .A1(n15864), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17378) );
  AOI22_X1 U20578 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13971), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17377) );
  AOI22_X1 U20579 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17376) );
  NAND4_X1 U20580 ( .A1(n17379), .A2(n17378), .A3(n17377), .A4(n17376), .ZN(
        n17386) );
  AOI22_X1 U20581 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17384) );
  AOI22_X1 U20582 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17380), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17383) );
  AOI22_X1 U20583 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9658), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17381) );
  NAND4_X1 U20584 ( .A1(n17384), .A2(n17383), .A3(n17382), .A4(n17381), .ZN(
        n17385) );
  NOR2_X1 U20585 ( .A1(n17386), .A2(n17385), .ZN(n17600) );
  OAI21_X1 U20586 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17387), .A(n17494), .ZN(
        n17388) );
  OAI22_X1 U20587 ( .A1(n17600), .A2(n17494), .B1(n17389), .B2(n17388), .ZN(
        P3_U2689) );
  OR2_X1 U20588 ( .A1(n17489), .A2(n17390), .ZN(n17414) );
  AOI22_X1 U20589 ( .A1(n17380), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17432), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17394) );
  AOI22_X1 U20590 ( .A1(n15864), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17393) );
  AOI22_X1 U20591 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17392) );
  AOI22_X1 U20592 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n15756), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17391) );
  NAND4_X1 U20593 ( .A1(n17394), .A2(n17393), .A3(n17392), .A4(n17391), .ZN(
        n17401) );
  AOI22_X1 U20594 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17399) );
  AOI22_X1 U20595 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n15929), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17398) );
  AOI22_X1 U20596 ( .A1(n17407), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17397) );
  AOI22_X1 U20597 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9658), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17396) );
  NAND4_X1 U20598 ( .A1(n17399), .A2(n17398), .A3(n17397), .A4(n17396), .ZN(
        n17400) );
  NOR2_X1 U20599 ( .A1(n17401), .A2(n17400), .ZN(n17606) );
  NAND3_X1 U20600 ( .A1(n17414), .A2(P3_EBX_REG_12__SCAN_IN), .A3(n17494), 
        .ZN(n17402) );
  OAI221_X1 U20601 ( .B1(n17414), .B2(P3_EBX_REG_12__SCAN_IN), .C1(n17494), 
        .C2(n17606), .A(n17402), .ZN(P3_U2691) );
  AOI22_X1 U20602 ( .A1(n15864), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n15756), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17406) );
  AOI22_X1 U20603 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17405) );
  AOI22_X1 U20604 ( .A1(n17380), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17404) );
  AOI22_X1 U20605 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17403) );
  NAND4_X1 U20606 ( .A1(n17406), .A2(n17405), .A3(n17404), .A4(n17403), .ZN(
        n17413) );
  AOI22_X1 U20607 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17411) );
  AOI22_X1 U20608 ( .A1(n17407), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17410) );
  AOI22_X1 U20609 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n15929), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17409) );
  AOI22_X1 U20610 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9658), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17408) );
  NAND4_X1 U20611 ( .A1(n17411), .A2(n17410), .A3(n17409), .A4(n17408), .ZN(
        n17412) );
  NOR2_X1 U20612 ( .A1(n17413), .A2(n17412), .ZN(n17611) );
  OAI211_X1 U20613 ( .C1(P3_EBX_REG_11__SCAN_IN), .C2(n17415), .A(n17414), .B(
        n17494), .ZN(n17416) );
  OAI21_X1 U20614 ( .B1(n17611), .B2(n17494), .A(n17416), .ZN(P3_U2692) );
  OAI21_X1 U20615 ( .B1(n17427), .B2(n17468), .A(n17494), .ZN(n17445) );
  AOI22_X1 U20616 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17420) );
  AOI22_X1 U20617 ( .A1(n15864), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17419) );
  AOI22_X1 U20618 ( .A1(n15756), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13971), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17418) );
  AOI22_X1 U20619 ( .A1(n17432), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17417) );
  NAND4_X1 U20620 ( .A1(n17420), .A2(n17419), .A3(n17418), .A4(n17417), .ZN(
        n17426) );
  AOI22_X1 U20621 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17424) );
  AOI22_X1 U20622 ( .A1(n17380), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17423) );
  AOI22_X1 U20623 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n15929), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17422) );
  AOI22_X1 U20624 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9658), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17421) );
  NAND4_X1 U20625 ( .A1(n17424), .A2(n17423), .A3(n17422), .A4(n17421), .ZN(
        n17425) );
  NOR2_X1 U20626 ( .A1(n17426), .A2(n17425), .ZN(n17618) );
  INV_X1 U20627 ( .A(n17618), .ZN(n17429) );
  NOR2_X1 U20628 ( .A1(n17473), .A2(n17502), .ZN(n17485) );
  NOR2_X1 U20629 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17427), .ZN(n17428) );
  AOI22_X1 U20630 ( .A1(n17500), .A2(n17429), .B1(n17485), .B2(n17428), .ZN(
        n17430) );
  OAI21_X1 U20631 ( .B1(n17431), .B2(n17445), .A(n17430), .ZN(P3_U2693) );
  AOI22_X1 U20632 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n17212), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17437) );
  AOI22_X1 U20633 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n9649), .B1(
        n17380), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17436) );
  AOI22_X1 U20634 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17435) );
  AOI22_X1 U20635 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n9655), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n17447), .ZN(n17434) );
  NAND4_X1 U20636 ( .A1(n17437), .A2(n17436), .A3(n17435), .A4(n17434), .ZN(
        n17443) );
  AOI22_X1 U20637 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n15860), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17441) );
  AOI22_X1 U20638 ( .A1(n9656), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n15929), .ZN(n17440) );
  AOI22_X1 U20639 ( .A1(n15864), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17456), .ZN(n17439) );
  AOI22_X1 U20640 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n9658), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n9667), .ZN(n17438) );
  NAND4_X1 U20641 ( .A1(n17441), .A2(n17440), .A3(n17439), .A4(n17438), .ZN(
        n17442) );
  NOR2_X1 U20642 ( .A1(n17443), .A2(n17442), .ZN(n17620) );
  NAND2_X1 U20643 ( .A1(n17444), .A2(n17478), .ZN(n17465) );
  INV_X1 U20644 ( .A(n17465), .ZN(n17463) );
  AOI21_X1 U20645 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17463), .A(
        P3_EBX_REG_9__SCAN_IN), .ZN(n17446) );
  OAI22_X1 U20646 ( .A1(n17620), .A2(n17494), .B1(n17446), .B2(n17445), .ZN(
        P3_U2694) );
  AOI22_X1 U20647 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17447), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17454) );
  AOI22_X1 U20648 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17432), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17452) );
  AOI22_X1 U20649 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17380), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17451) );
  NAND4_X1 U20650 ( .A1(n17454), .A2(n17453), .A3(n17452), .A4(n17451), .ZN(
        n17462) );
  AOI22_X1 U20651 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17460) );
  AOI22_X1 U20652 ( .A1(n15756), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17459) );
  AOI22_X1 U20653 ( .A1(n17456), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17458) );
  AOI22_X1 U20654 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9658), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17457) );
  NAND4_X1 U20655 ( .A1(n17460), .A2(n17459), .A3(n17458), .A4(n17457), .ZN(
        n17461) );
  NOR2_X1 U20656 ( .A1(n17462), .A2(n17461), .ZN(n17624) );
  INV_X1 U20657 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n17464) );
  OAI33_X1 U20658 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17489), .A3(n17465), .B1(
        n17464), .B2(n17500), .B3(n17463), .ZN(n17466) );
  INV_X1 U20659 ( .A(n17466), .ZN(n17467) );
  OAI21_X1 U20660 ( .B1(n17624), .B2(n17494), .A(n17467), .ZN(P3_U2695) );
  NOR3_X1 U20661 ( .A1(n17469), .A2(n17474), .A3(n17468), .ZN(n17470) );
  NAND2_X1 U20662 ( .A1(n18512), .A2(n17470), .ZN(n17472) );
  NOR2_X1 U20663 ( .A1(n17500), .A2(n17470), .ZN(n17475) );
  AOI22_X1 U20664 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17500), .B1(
        P3_EBX_REG_7__SCAN_IN), .B2(n17475), .ZN(n17471) );
  OAI21_X1 U20665 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17472), .A(n17471), .ZN(
        P3_U2696) );
  INV_X1 U20666 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17477) );
  NOR3_X1 U20667 ( .A1(n17474), .A2(n17473), .A3(n17502), .ZN(n17481) );
  OAI21_X1 U20668 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17481), .A(n17475), .ZN(
        n17476) );
  OAI21_X1 U20669 ( .B1(n17494), .B2(n17477), .A(n17476), .ZN(P3_U2697) );
  OAI21_X1 U20670 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17478), .A(n17494), .ZN(
        n17480) );
  INV_X1 U20671 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17479) );
  OAI22_X1 U20672 ( .A1(n17481), .A2(n17480), .B1(n17479), .B2(n17494), .ZN(
        P3_U2698) );
  NOR2_X1 U20673 ( .A1(n17482), .A2(n17502), .ZN(n17491) );
  AND2_X1 U20674 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17491), .ZN(n17488) );
  AOI21_X1 U20675 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17494), .A(n17488), .ZN(
        n17484) );
  INV_X1 U20676 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17483) );
  OAI22_X1 U20677 ( .A1(n17485), .A2(n17484), .B1(n17483), .B2(n17494), .ZN(
        P3_U2699) );
  AOI21_X1 U20678 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17494), .A(n17491), .ZN(
        n17487) );
  INV_X1 U20679 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17486) );
  OAI22_X1 U20680 ( .A1(n17488), .A2(n17487), .B1(n17486), .B2(n17494), .ZN(
        P3_U2700) );
  AOI221_X1 U20681 ( .B1(n17490), .B2(n17496), .C1(n17489), .C2(n17496), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n17492) );
  AOI211_X1 U20682 ( .C1(n17500), .C2(n17493), .A(n17492), .B(n17491), .ZN(
        P3_U2701) );
  OAI222_X1 U20683 ( .A1(n17498), .A2(n17502), .B1(n17497), .B2(n17496), .C1(
        n17495), .C2(n17494), .ZN(P3_U2702) );
  AOI22_X1 U20684 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17500), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17499), .ZN(n17501) );
  OAI21_X1 U20685 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17502), .A(n17501), .ZN(
        P3_U2703) );
  NAND2_X1 U20686 ( .A1(n17603), .A2(n17503), .ZN(n17553) );
  INV_X1 U20687 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17725) );
  INV_X1 U20688 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17721) );
  INV_X1 U20689 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17719) );
  INV_X1 U20690 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17717) );
  INV_X1 U20691 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17703) );
  INV_X1 U20692 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17735) );
  NAND4_X1 U20693 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17504) );
  NOR3_X1 U20694 ( .A1(n17735), .A2(n17733), .A3(n17504), .ZN(n17505) );
  NAND3_X1 U20695 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(n17505), .ZN(n17595) );
  NAND3_X1 U20696 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .A3(P3_EAX_REG_11__SCAN_IN), .ZN(n17596) );
  NAND4_X1 U20697 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_10__SCAN_IN), 
        .A3(P3_EAX_REG_9__SCAN_IN), .A4(P3_EAX_REG_8__SCAN_IN), .ZN(n17506) );
  NAND2_X1 U20698 ( .A1(P3_EAX_REG_15__SCAN_IN), .A2(n17594), .ZN(n17590) );
  INV_X1 U20699 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17715) );
  INV_X1 U20700 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17713) );
  INV_X1 U20701 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17707) );
  INV_X1 U20702 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17705) );
  NOR4_X1 U20703 ( .A1(n17715), .A2(n17713), .A3(n17707), .A4(n17705), .ZN(
        n17507) );
  NAND4_X1 U20704 ( .A1(n17585), .A2(P3_EAX_REG_20__SCAN_IN), .A3(
        P3_EAX_REG_19__SCAN_IN), .A4(n17507), .ZN(n17548) );
  NAND2_X1 U20705 ( .A1(n18512), .A2(n17547), .ZN(n17540) );
  NAND2_X1 U20706 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17536), .ZN(n17531) );
  NAND2_X1 U20707 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17527), .ZN(n17522) );
  NAND2_X1 U20708 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17519), .ZN(n17518) );
  NOR2_X1 U20709 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n17518), .ZN(n17509) );
  NAND2_X1 U20710 ( .A1(n17646), .A2(n17518), .ZN(n17516) );
  OAI21_X1 U20711 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17652), .A(n17516), .ZN(
        n17508) );
  AOI22_X1 U20712 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17509), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17508), .ZN(n17510) );
  OAI21_X1 U20713 ( .B1(n19482), .B2(n17553), .A(n17510), .ZN(P3_U2704) );
  INV_X1 U20714 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17731) );
  OAI22_X1 U20715 ( .A1(n17513), .A2(n17648), .B1(n17512), .B2(n17553), .ZN(
        n17514) );
  AOI21_X1 U20716 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17584), .A(n17514), .ZN(
        n17515) );
  OAI221_X1 U20717 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17518), .C1(n17731), 
        .C2(n17516), .A(n17515), .ZN(P3_U2705) );
  AOI22_X1 U20718 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17584), .B1(n17655), .B2(
        n17517), .ZN(n17521) );
  OAI211_X1 U20719 ( .C1(n17519), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17646), .B(
        n17518), .ZN(n17520) );
  OAI211_X1 U20720 ( .C1(n17553), .C2(n19472), .A(n17521), .B(n17520), .ZN(
        P3_U2706) );
  AOI22_X1 U20721 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17584), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17583), .ZN(n17524) );
  OAI211_X1 U20722 ( .C1(n17527), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17646), .B(
        n17522), .ZN(n17523) );
  OAI211_X1 U20723 ( .C1(n17525), .C2(n17648), .A(n17524), .B(n17523), .ZN(
        P3_U2707) );
  AOI22_X1 U20724 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17584), .B1(n17655), .B2(
        n17526), .ZN(n17530) );
  AOI211_X1 U20725 ( .C1(n17725), .C2(n17531), .A(n17527), .B(n17603), .ZN(
        n17528) );
  INV_X1 U20726 ( .A(n17528), .ZN(n17529) );
  OAI211_X1 U20727 ( .C1(n17553), .C2(n19463), .A(n17530), .B(n17529), .ZN(
        P3_U2708) );
  AOI22_X1 U20728 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17584), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17583), .ZN(n17533) );
  OAI211_X1 U20729 ( .C1(n17536), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17646), .B(
        n17531), .ZN(n17532) );
  OAI211_X1 U20730 ( .C1(n17534), .C2(n17648), .A(n17533), .B(n17532), .ZN(
        P3_U2709) );
  AOI22_X1 U20731 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17584), .B1(n17655), .B2(
        n17535), .ZN(n17539) );
  AOI211_X1 U20732 ( .C1(n17721), .C2(n17541), .A(n17536), .B(n17603), .ZN(
        n17537) );
  INV_X1 U20733 ( .A(n17537), .ZN(n17538) );
  OAI211_X1 U20734 ( .C1(n17553), .C2(n18485), .A(n17539), .B(n17538), .ZN(
        P3_U2710) );
  AOI22_X1 U20735 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17584), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17583), .ZN(n17544) );
  OAI21_X1 U20736 ( .B1(n17719), .B2(n17603), .A(n17540), .ZN(n17542) );
  NAND2_X1 U20737 ( .A1(n17542), .A2(n17541), .ZN(n17543) );
  OAI211_X1 U20738 ( .C1(n17545), .C2(n17648), .A(n17544), .B(n17543), .ZN(
        P3_U2711) );
  AOI22_X1 U20739 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n17583), .B1(n17655), .B2(
        n17546), .ZN(n17551) );
  AOI211_X1 U20740 ( .C1(n17717), .C2(n17548), .A(n17603), .B(n17547), .ZN(
        n17549) );
  AOI21_X1 U20741 ( .B1(n17584), .B2(BUF2_REG_7__SCAN_IN), .A(n17549), .ZN(
        n17550) );
  NAND2_X1 U20742 ( .A1(n17551), .A2(n17550), .ZN(P3_U2712) );
  NAND2_X1 U20743 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .ZN(n17552) );
  NAND2_X1 U20744 ( .A1(n18512), .A2(n17585), .ZN(n17576) );
  NAND2_X1 U20745 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17577), .ZN(n17572) );
  NAND2_X1 U20746 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17562), .ZN(n17558) );
  NAND2_X1 U20747 ( .A1(n17558), .A2(P3_EAX_REG_22__SCAN_IN), .ZN(n17557) );
  OAI22_X1 U20748 ( .A1(n17554), .A2(n17648), .B1(n18504), .B2(n17553), .ZN(
        n17555) );
  AOI21_X1 U20749 ( .B1(BUF2_REG_6__SCAN_IN), .B2(n17584), .A(n17555), .ZN(
        n17556) );
  OAI221_X1 U20750 ( .B1(n17558), .B2(P3_EAX_REG_22__SCAN_IN), .C1(n17557), 
        .C2(n17603), .A(n17556), .ZN(P3_U2713) );
  AOI22_X1 U20751 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17584), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n17583), .ZN(n17560) );
  OAI211_X1 U20752 ( .C1(n17562), .C2(P3_EAX_REG_21__SCAN_IN), .A(n17646), .B(
        n17558), .ZN(n17559) );
  OAI211_X1 U20753 ( .C1(n17561), .C2(n17648), .A(n17560), .B(n17559), .ZN(
        P3_U2714) );
  AOI22_X1 U20754 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17584), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17583), .ZN(n17565) );
  INV_X1 U20755 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17711) );
  INV_X1 U20756 ( .A(n17572), .ZN(n17568) );
  NAND2_X1 U20757 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17568), .ZN(n17567) );
  AOI211_X1 U20758 ( .C1(n17711), .C2(n17567), .A(n17562), .B(n17603), .ZN(
        n17563) );
  INV_X1 U20759 ( .A(n17563), .ZN(n17564) );
  OAI211_X1 U20760 ( .C1(n17566), .C2(n17648), .A(n17565), .B(n17564), .ZN(
        P3_U2715) );
  AOI22_X1 U20761 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17584), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17583), .ZN(n17570) );
  OAI211_X1 U20762 ( .C1(n17568), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17646), .B(
        n17567), .ZN(n17569) );
  OAI211_X1 U20763 ( .C1(n17571), .C2(n17648), .A(n17570), .B(n17569), .ZN(
        P3_U2716) );
  AOI22_X1 U20764 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17584), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17583), .ZN(n17574) );
  OAI211_X1 U20765 ( .C1(n17577), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17646), .B(
        n17572), .ZN(n17573) );
  OAI211_X1 U20766 ( .C1(n17575), .C2(n17648), .A(n17574), .B(n17573), .ZN(
        P3_U2717) );
  AOI22_X1 U20767 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17584), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17583), .ZN(n17581) );
  OAI21_X1 U20768 ( .B1(n17705), .B2(n17603), .A(n17576), .ZN(n17579) );
  INV_X1 U20769 ( .A(n17577), .ZN(n17578) );
  NAND2_X1 U20770 ( .A1(n17579), .A2(n17578), .ZN(n17580) );
  OAI211_X1 U20771 ( .C1(n17582), .C2(n17648), .A(n17581), .B(n17580), .ZN(
        P3_U2718) );
  AOI22_X1 U20772 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17584), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17583), .ZN(n17588) );
  AOI211_X1 U20773 ( .C1(n17703), .C2(n17590), .A(n17603), .B(n17585), .ZN(
        n17586) );
  INV_X1 U20774 ( .A(n17586), .ZN(n17587) );
  OAI211_X1 U20775 ( .C1(n17589), .C2(n17648), .A(n17588), .B(n17587), .ZN(
        P3_U2719) );
  OAI211_X1 U20776 ( .C1(P3_EAX_REG_15__SCAN_IN), .C2(n17594), .A(n17646), .B(
        n17590), .ZN(n17592) );
  NAND2_X1 U20777 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17656), .ZN(n17591) );
  OAI211_X1 U20778 ( .C1(n17593), .C2(n17648), .A(n17592), .B(n17591), .ZN(
        P3_U2720) );
  INV_X1 U20779 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17763) );
  NOR3_X1 U20780 ( .A1(n17603), .A2(n17594), .A3(n17763), .ZN(n17598) );
  INV_X1 U20781 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17751) );
  NOR2_X1 U20782 ( .A1(n17595), .A2(n17652), .ZN(n17630) );
  NAND2_X1 U20783 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17630), .ZN(n17619) );
  NAND2_X1 U20784 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17622), .ZN(n17615) );
  NOR3_X1 U20785 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17596), .A3(n17615), .ZN(
        n17597) );
  AOI211_X1 U20786 ( .C1(n17656), .C2(BUF2_REG_14__SCAN_IN), .A(n17598), .B(
        n17597), .ZN(n17599) );
  OAI21_X1 U20787 ( .B1(n17600), .B2(n17648), .A(n17599), .ZN(P3_U2721) );
  INV_X1 U20788 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17755) );
  NOR2_X1 U20789 ( .A1(n17755), .A2(n17615), .ZN(n17613) );
  NAND2_X1 U20790 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17613), .ZN(n17605) );
  NAND2_X1 U20791 ( .A1(n17605), .A2(P3_EAX_REG_13__SCAN_IN), .ZN(n17604) );
  AOI22_X1 U20792 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17656), .B1(n17655), .B2(
        n17601), .ZN(n17602) );
  OAI221_X1 U20793 ( .B1(n17605), .B2(P3_EAX_REG_13__SCAN_IN), .C1(n17604), 
        .C2(n17603), .A(n17602), .ZN(P3_U2722) );
  INV_X1 U20794 ( .A(n17605), .ZN(n17608) );
  AOI21_X1 U20795 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17646), .A(n17613), .ZN(
        n17607) );
  OAI222_X1 U20796 ( .A1(n17651), .A2(n17609), .B1(n17608), .B2(n17607), .C1(
        n17648), .C2(n17606), .ZN(P3_U2723) );
  INV_X1 U20797 ( .A(n17615), .ZN(n17610) );
  AOI21_X1 U20798 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17646), .A(n17610), .ZN(
        n17612) );
  OAI222_X1 U20799 ( .A1(n17651), .A2(n17614), .B1(n17613), .B2(n17612), .C1(
        n17648), .C2(n17611), .ZN(P3_U2724) );
  OAI211_X1 U20800 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n17622), .A(n17646), .B(
        n17615), .ZN(n17617) );
  NAND2_X1 U20801 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17656), .ZN(n17616) );
  OAI211_X1 U20802 ( .C1(n17618), .C2(n17648), .A(n17617), .B(n17616), .ZN(
        P3_U2725) );
  INV_X1 U20803 ( .A(n17619), .ZN(n17626) );
  AOI21_X1 U20804 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17646), .A(n17626), .ZN(
        n17621) );
  OAI222_X1 U20805 ( .A1(n17651), .A2(n17623), .B1(n17622), .B2(n17621), .C1(
        n17648), .C2(n17620), .ZN(P3_U2726) );
  AOI21_X1 U20806 ( .B1(P3_EAX_REG_8__SCAN_IN), .B2(n17646), .A(n17630), .ZN(
        n17625) );
  OAI222_X1 U20807 ( .A1(n17651), .A2(n17627), .B1(n17626), .B2(n17625), .C1(
        n17648), .C2(n17624), .ZN(P3_U2727) );
  INV_X1 U20808 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17745) );
  INV_X1 U20809 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17741) );
  INV_X1 U20810 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17737) );
  NOR4_X1 U20811 ( .A1(n17737), .A2(n17735), .A3(n17733), .A4(n17652), .ZN(
        n17650) );
  NAND2_X1 U20812 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17650), .ZN(n17638) );
  NOR2_X1 U20813 ( .A1(n17741), .A2(n17638), .ZN(n17641) );
  NAND2_X1 U20814 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17641), .ZN(n17631) );
  NOR2_X1 U20815 ( .A1(n17745), .A2(n17631), .ZN(n17634) );
  AOI21_X1 U20816 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17646), .A(n17634), .ZN(
        n17629) );
  OAI222_X1 U20817 ( .A1(n17651), .A2(n18509), .B1(n17630), .B2(n17629), .C1(
        n17648), .C2(n17628), .ZN(P3_U2728) );
  INV_X1 U20818 ( .A(n17631), .ZN(n17637) );
  AOI21_X1 U20819 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17646), .A(n17637), .ZN(
        n17633) );
  OAI222_X1 U20820 ( .A1(n18505), .A2(n17651), .B1(n17634), .B2(n17633), .C1(
        n17648), .C2(n17632), .ZN(P3_U2729) );
  AOI21_X1 U20821 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17646), .A(n17641), .ZN(
        n17636) );
  OAI222_X1 U20822 ( .A1(n18500), .A2(n17651), .B1(n17637), .B2(n17636), .C1(
        n17648), .C2(n17635), .ZN(P3_U2730) );
  INV_X1 U20823 ( .A(n17638), .ZN(n17644) );
  AOI21_X1 U20824 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17646), .A(n17644), .ZN(
        n17640) );
  OAI222_X1 U20825 ( .A1(n18496), .A2(n17651), .B1(n17641), .B2(n17640), .C1(
        n17648), .C2(n17639), .ZN(P3_U2731) );
  AOI21_X1 U20826 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17646), .A(n17650), .ZN(
        n17643) );
  OAI222_X1 U20827 ( .A1(n18492), .A2(n17651), .B1(n17644), .B2(n17643), .C1(
        n17648), .C2(n17642), .ZN(P3_U2732) );
  NOR3_X1 U20828 ( .A1(n17735), .A2(n17733), .A3(n17652), .ZN(n17645) );
  AOI21_X1 U20829 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17646), .A(n17645), .ZN(
        n17649) );
  OAI222_X1 U20830 ( .A1(n18488), .A2(n17651), .B1(n17650), .B2(n17649), .C1(
        n17648), .C2(n17647), .ZN(P3_U2733) );
  OR2_X1 U20831 ( .A1(n17733), .A2(n17652), .ZN(n17659) );
  AOI21_X1 U20832 ( .B1(n18512), .B2(n17733), .A(n17653), .ZN(n17658) );
  AOI22_X1 U20833 ( .A1(n17656), .A2(BUF2_REG_1__SCAN_IN), .B1(n17655), .B2(
        n17654), .ZN(n17657) );
  OAI221_X1 U20834 ( .B1(P3_EAX_REG_1__SCAN_IN), .B2(n17659), .C1(n17735), 
        .C2(n17658), .A(n17657), .ZN(P3_U2734) );
  AND2_X1 U20835 ( .A1(n17676), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U20836 ( .A1(n17679), .A2(n17661), .ZN(n17678) );
  AOI22_X1 U20837 ( .A1(n19133), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(n17695), .ZN(n17662) );
  OAI21_X1 U20838 ( .B1(n17731), .B2(n17678), .A(n17662), .ZN(P3_U2737) );
  INV_X1 U20839 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17729) );
  AOI22_X1 U20840 ( .A1(n19133), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17695), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17663) );
  OAI21_X1 U20841 ( .B1(n17729), .B2(n17678), .A(n17663), .ZN(P3_U2738) );
  INV_X1 U20842 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17727) );
  AOI22_X1 U20843 ( .A1(n19133), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17695), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17664) );
  OAI21_X1 U20844 ( .B1(n17727), .B2(n17678), .A(n17664), .ZN(P3_U2739) );
  AOI22_X1 U20845 ( .A1(n19133), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17676), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17665) );
  OAI21_X1 U20846 ( .B1(n17725), .B2(n17678), .A(n17665), .ZN(P3_U2740) );
  INV_X1 U20847 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17723) );
  AOI22_X1 U20848 ( .A1(n19133), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17695), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17666) );
  OAI21_X1 U20849 ( .B1(n17723), .B2(n17678), .A(n17666), .ZN(P3_U2741) );
  AOI22_X1 U20850 ( .A1(n19133), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17676), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17667) );
  OAI21_X1 U20851 ( .B1(n17721), .B2(n17678), .A(n17667), .ZN(P3_U2742) );
  AOI22_X1 U20852 ( .A1(n19133), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17676), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17668) );
  OAI21_X1 U20853 ( .B1(n17719), .B2(n17678), .A(n17668), .ZN(P3_U2743) );
  CLKBUF_X1 U20854 ( .A(n19133), .Z(n17696) );
  AOI22_X1 U20855 ( .A1(n17696), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17695), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17669) );
  OAI21_X1 U20856 ( .B1(n17717), .B2(n17678), .A(n17669), .ZN(P3_U2744) );
  AOI22_X1 U20857 ( .A1(n17696), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17676), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17670) );
  OAI21_X1 U20858 ( .B1(n17715), .B2(n17678), .A(n17670), .ZN(P3_U2745) );
  AOI22_X1 U20859 ( .A1(n17696), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17676), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17671) );
  OAI21_X1 U20860 ( .B1(n17713), .B2(n17678), .A(n17671), .ZN(P3_U2746) );
  AOI22_X1 U20861 ( .A1(n17696), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17676), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17672) );
  OAI21_X1 U20862 ( .B1(n17711), .B2(n17678), .A(n17672), .ZN(P3_U2747) );
  INV_X1 U20863 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17709) );
  AOI22_X1 U20864 ( .A1(n17696), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17676), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17673) );
  OAI21_X1 U20865 ( .B1(n17709), .B2(n17678), .A(n17673), .ZN(P3_U2748) );
  AOI22_X1 U20866 ( .A1(n17696), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17676), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17674) );
  OAI21_X1 U20867 ( .B1(n17707), .B2(n17678), .A(n17674), .ZN(P3_U2749) );
  AOI22_X1 U20868 ( .A1(n17696), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17676), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17675) );
  OAI21_X1 U20869 ( .B1(n17705), .B2(n17678), .A(n17675), .ZN(P3_U2750) );
  AOI22_X1 U20870 ( .A1(n17696), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17676), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17677) );
  OAI21_X1 U20871 ( .B1(n17703), .B2(n17678), .A(n17677), .ZN(P3_U2751) );
  INV_X1 U20872 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17768) );
  AOI22_X1 U20873 ( .A1(n17696), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17695), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17680) );
  OAI21_X1 U20874 ( .B1(n17768), .B2(n17698), .A(n17680), .ZN(P3_U2752) );
  AOI22_X1 U20875 ( .A1(n17696), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17695), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17681) );
  OAI21_X1 U20876 ( .B1(n17763), .B2(n17698), .A(n17681), .ZN(P3_U2753) );
  INV_X1 U20877 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17760) );
  AOI22_X1 U20878 ( .A1(n17696), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17695), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17682) );
  OAI21_X1 U20879 ( .B1(n17760), .B2(n17698), .A(n17682), .ZN(P3_U2754) );
  INV_X1 U20880 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17757) );
  AOI22_X1 U20881 ( .A1(n17696), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17695), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17683) );
  OAI21_X1 U20882 ( .B1(n17757), .B2(n17698), .A(n17683), .ZN(P3_U2755) );
  AOI22_X1 U20883 ( .A1(n17696), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17695), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17684) );
  OAI21_X1 U20884 ( .B1(n17755), .B2(n17698), .A(n17684), .ZN(P3_U2756) );
  INV_X1 U20885 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17753) );
  AOI22_X1 U20886 ( .A1(n17696), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17695), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17685) );
  OAI21_X1 U20887 ( .B1(n17753), .B2(n17698), .A(n17685), .ZN(P3_U2757) );
  AOI22_X1 U20888 ( .A1(n17696), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17695), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17686) );
  OAI21_X1 U20889 ( .B1(n17751), .B2(n17698), .A(n17686), .ZN(P3_U2758) );
  INV_X1 U20890 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17749) );
  AOI22_X1 U20891 ( .A1(n17696), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17695), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17687) );
  OAI21_X1 U20892 ( .B1(n17749), .B2(n17698), .A(n17687), .ZN(P3_U2759) );
  INV_X1 U20893 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17747) );
  AOI22_X1 U20894 ( .A1(n17696), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17695), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17688) );
  OAI21_X1 U20895 ( .B1(n17747), .B2(n17698), .A(n17688), .ZN(P3_U2760) );
  AOI22_X1 U20896 ( .A1(n17696), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17695), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17689) );
  OAI21_X1 U20897 ( .B1(n17745), .B2(n17698), .A(n17689), .ZN(P3_U2761) );
  INV_X1 U20898 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17743) );
  AOI22_X1 U20899 ( .A1(n17696), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17695), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17690) );
  OAI21_X1 U20900 ( .B1(n17743), .B2(n17698), .A(n17690), .ZN(P3_U2762) );
  AOI22_X1 U20901 ( .A1(n17696), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17695), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17691) );
  OAI21_X1 U20902 ( .B1(n17741), .B2(n17698), .A(n17691), .ZN(P3_U2763) );
  INV_X1 U20903 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17739) );
  AOI22_X1 U20904 ( .A1(n17696), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17695), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17692) );
  OAI21_X1 U20905 ( .B1(n17739), .B2(n17698), .A(n17692), .ZN(P3_U2764) );
  AOI22_X1 U20906 ( .A1(n17696), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17695), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17693) );
  OAI21_X1 U20907 ( .B1(n17737), .B2(n17698), .A(n17693), .ZN(P3_U2765) );
  AOI22_X1 U20908 ( .A1(n17696), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17695), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17694) );
  OAI21_X1 U20909 ( .B1(n17735), .B2(n17698), .A(n17694), .ZN(P3_U2766) );
  AOI22_X1 U20910 ( .A1(n17696), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17695), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17697) );
  OAI21_X1 U20911 ( .B1(n17733), .B2(n17698), .A(n17697), .ZN(P3_U2767) );
  AOI22_X1 U20912 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17765), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17764), .ZN(n17702) );
  OAI21_X1 U20913 ( .B1(n17703), .B2(n17767), .A(n17702), .ZN(P3_U2768) );
  AOI22_X1 U20914 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17765), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17764), .ZN(n17704) );
  OAI21_X1 U20915 ( .B1(n17705), .B2(n17767), .A(n17704), .ZN(P3_U2769) );
  AOI22_X1 U20916 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17765), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17764), .ZN(n17706) );
  OAI21_X1 U20917 ( .B1(n17707), .B2(n17767), .A(n17706), .ZN(P3_U2770) );
  AOI22_X1 U20918 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17765), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17764), .ZN(n17708) );
  OAI21_X1 U20919 ( .B1(n17709), .B2(n17767), .A(n17708), .ZN(P3_U2771) );
  AOI22_X1 U20920 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17761), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17764), .ZN(n17710) );
  OAI21_X1 U20921 ( .B1(n17711), .B2(n17767), .A(n17710), .ZN(P3_U2772) );
  AOI22_X1 U20922 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17761), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17764), .ZN(n17712) );
  OAI21_X1 U20923 ( .B1(n17713), .B2(n17767), .A(n17712), .ZN(P3_U2773) );
  AOI22_X1 U20924 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17761), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17764), .ZN(n17714) );
  OAI21_X1 U20925 ( .B1(n17715), .B2(n17767), .A(n17714), .ZN(P3_U2774) );
  AOI22_X1 U20926 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17761), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17764), .ZN(n17716) );
  OAI21_X1 U20927 ( .B1(n17717), .B2(n17767), .A(n17716), .ZN(P3_U2775) );
  AOI22_X1 U20928 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17761), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17764), .ZN(n17718) );
  OAI21_X1 U20929 ( .B1(n17719), .B2(n17767), .A(n17718), .ZN(P3_U2776) );
  AOI22_X1 U20930 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17761), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17764), .ZN(n17720) );
  OAI21_X1 U20931 ( .B1(n17721), .B2(n17767), .A(n17720), .ZN(P3_U2777) );
  AOI22_X1 U20932 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17761), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17764), .ZN(n17722) );
  OAI21_X1 U20933 ( .B1(n17723), .B2(n17767), .A(n17722), .ZN(P3_U2778) );
  AOI22_X1 U20934 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17761), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17764), .ZN(n17724) );
  OAI21_X1 U20935 ( .B1(n17725), .B2(n17767), .A(n17724), .ZN(P3_U2779) );
  AOI22_X1 U20936 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17765), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17764), .ZN(n17726) );
  OAI21_X1 U20937 ( .B1(n17727), .B2(n17767), .A(n17726), .ZN(P3_U2780) );
  AOI22_X1 U20938 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17765), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17764), .ZN(n17728) );
  OAI21_X1 U20939 ( .B1(n17729), .B2(n17767), .A(n17728), .ZN(P3_U2781) );
  AOI22_X1 U20940 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17765), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17764), .ZN(n17730) );
  OAI21_X1 U20941 ( .B1(n17731), .B2(n17767), .A(n17730), .ZN(P3_U2782) );
  AOI22_X1 U20942 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17765), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17764), .ZN(n17732) );
  OAI21_X1 U20943 ( .B1(n17733), .B2(n17767), .A(n17732), .ZN(P3_U2783) );
  AOI22_X1 U20944 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17765), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17764), .ZN(n17734) );
  OAI21_X1 U20945 ( .B1(n17735), .B2(n17767), .A(n17734), .ZN(P3_U2784) );
  AOI22_X1 U20946 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17765), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17764), .ZN(n17736) );
  OAI21_X1 U20947 ( .B1(n17737), .B2(n17767), .A(n17736), .ZN(P3_U2785) );
  AOI22_X1 U20948 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17765), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17764), .ZN(n17738) );
  OAI21_X1 U20949 ( .B1(n17739), .B2(n17767), .A(n17738), .ZN(P3_U2786) );
  AOI22_X1 U20950 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17765), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17758), .ZN(n17740) );
  OAI21_X1 U20951 ( .B1(n17741), .B2(n17767), .A(n17740), .ZN(P3_U2787) );
  AOI22_X1 U20952 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17765), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17758), .ZN(n17742) );
  OAI21_X1 U20953 ( .B1(n17743), .B2(n17767), .A(n17742), .ZN(P3_U2788) );
  AOI22_X1 U20954 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17765), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17758), .ZN(n17744) );
  OAI21_X1 U20955 ( .B1(n17745), .B2(n17767), .A(n17744), .ZN(P3_U2789) );
  AOI22_X1 U20956 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17765), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17758), .ZN(n17746) );
  OAI21_X1 U20957 ( .B1(n17747), .B2(n17767), .A(n17746), .ZN(P3_U2790) );
  AOI22_X1 U20958 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17765), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17758), .ZN(n17748) );
  OAI21_X1 U20959 ( .B1(n17749), .B2(n17767), .A(n17748), .ZN(P3_U2791) );
  AOI22_X1 U20960 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17761), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17758), .ZN(n17750) );
  OAI21_X1 U20961 ( .B1(n17751), .B2(n17767), .A(n17750), .ZN(P3_U2792) );
  AOI22_X1 U20962 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17765), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17758), .ZN(n17752) );
  OAI21_X1 U20963 ( .B1(n17753), .B2(n17767), .A(n17752), .ZN(P3_U2793) );
  AOI22_X1 U20964 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17761), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17758), .ZN(n17754) );
  OAI21_X1 U20965 ( .B1(n17755), .B2(n17767), .A(n17754), .ZN(P3_U2794) );
  AOI22_X1 U20966 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17765), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17758), .ZN(n17756) );
  OAI21_X1 U20967 ( .B1(n17757), .B2(n17767), .A(n17756), .ZN(P3_U2795) );
  AOI22_X1 U20968 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17765), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17758), .ZN(n17759) );
  OAI21_X1 U20969 ( .B1(n17760), .B2(n17767), .A(n17759), .ZN(P3_U2796) );
  AOI22_X1 U20970 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17761), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17764), .ZN(n17762) );
  OAI21_X1 U20971 ( .B1(n17763), .B2(n17767), .A(n17762), .ZN(P3_U2797) );
  AOI22_X1 U20972 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17765), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17764), .ZN(n17766) );
  OAI21_X1 U20973 ( .B1(n17768), .B2(n17767), .A(n17766), .ZN(P3_U2798) );
  OAI22_X1 U20974 ( .A1(n17771), .A2(n18045), .B1(n17769), .B2(n17977), .ZN(
        n17770) );
  NOR2_X1 U20975 ( .A1(n18101), .A2(n17770), .ZN(n17800) );
  OAI21_X1 U20976 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17881), .A(
        n17800), .ZN(n17788) );
  NAND2_X1 U20977 ( .A1(n17771), .A2(n17837), .ZN(n17793) );
  AOI221_X1 U20978 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C1(n17773), .C2(n17772), .A(
        n17793), .ZN(n17775) );
  AOI211_X1 U20979 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17788), .A(
        n17775), .B(n17774), .ZN(n17785) );
  NOR2_X1 U20980 ( .A1(n18132), .A2(n18012), .ZN(n17887) );
  INV_X1 U20981 ( .A(n18132), .ZN(n18149) );
  OAI22_X1 U20982 ( .A1(n18155), .A2(n18149), .B1(n18154), .B2(n18051), .ZN(
        n17806) );
  NOR2_X1 U20983 ( .A1(n10013), .A2(n17806), .ZN(n17777) );
  NOR3_X1 U20984 ( .A1(n17887), .A2(n17777), .A3(n17776), .ZN(n17782) );
  AOI211_X1 U20985 ( .C1(n17780), .C2(n17779), .A(n17778), .B(n18052), .ZN(
        n17781) );
  AOI211_X1 U20986 ( .C1(n17783), .C2(n17906), .A(n17782), .B(n17781), .ZN(
        n17784) );
  OAI211_X1 U20987 ( .C1(n17996), .C2(n17786), .A(n17785), .B(n17784), .ZN(
        P3_U2802) );
  AOI22_X1 U20988 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17788), .B1(
        n17980), .B2(n17787), .ZN(n17797) );
  INV_X1 U20989 ( .A(n17789), .ZN(n17790) );
  NAND2_X1 U20990 ( .A1(n17791), .A2(n17790), .ZN(n17792) );
  XNOR2_X1 U20991 ( .A(n17952), .B(n17792), .ZN(n18165) );
  OAI22_X1 U20992 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17793), .B1(
        n18165), .B2(n18052), .ZN(n17794) );
  AOI221_X1 U20993 ( .B1(n17795), .B2(n10013), .C1(n17806), .C2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n17794), .ZN(n17796) );
  OAI211_X1 U20994 ( .C1(n18447), .C2(n19062), .A(n17797), .B(n17796), .ZN(
        P3_U2803) );
  AOI21_X1 U20995 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17799), .A(
        n17798), .ZN(n18170) );
  AOI221_X1 U20996 ( .B1(n18819), .B2(n17802), .C1(n17801), .C2(n17802), .A(
        n17800), .ZN(n17805) );
  AOI21_X1 U20997 ( .B1(n17996), .B2(n17881), .A(n17803), .ZN(n17804) );
  AOI211_X1 U20998 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n9652), .A(n17805), .B(
        n17804), .ZN(n17808) );
  NOR3_X1 U20999 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18171), .A3(
        n18172), .ZN(n18166) );
  AOI22_X1 U21000 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17806), .B1(
        n17906), .B2(n18166), .ZN(n17807) );
  OAI211_X1 U21001 ( .C1(n18170), .C2(n18052), .A(n17808), .B(n17807), .ZN(
        P3_U2804) );
  OAI21_X1 U21002 ( .B1(n18050), .B2(n17810), .A(n17809), .ZN(n17811) );
  XNOR2_X1 U21003 ( .A(n17811), .B(n18171), .ZN(n18184) );
  OAI22_X1 U21004 ( .A1(n16619), .A2(n18819), .B1(n17812), .B2(n17977), .ZN(
        n17813) );
  NOR2_X1 U21005 ( .A1(n18101), .A2(n17813), .ZN(n17838) );
  OAI21_X1 U21006 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17977), .A(
        n17838), .ZN(n17829) );
  NOR2_X1 U21007 ( .A1(n18447), .A2(n19058), .ZN(n18179) );
  NAND2_X1 U21008 ( .A1(n16619), .A2(n17837), .ZN(n17826) );
  OAI21_X1 U21009 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17814), .ZN(n17815) );
  OAI22_X1 U21010 ( .A1(n17996), .A2(n17816), .B1(n17826), .B2(n17815), .ZN(
        n17817) );
  AOI211_X1 U21011 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17829), .A(
        n18179), .B(n17817), .ZN(n17821) );
  XNOR2_X1 U21012 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17818), .ZN(
        n18181) );
  XNOR2_X1 U21013 ( .A(n17819), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n18180) );
  AOI22_X1 U21014 ( .A1(n18132), .A2(n18181), .B1(n18012), .B2(n18180), .ZN(
        n17820) );
  OAI211_X1 U21015 ( .C1(n18052), .C2(n18184), .A(n17821), .B(n17820), .ZN(
        P3_U2805) );
  NAND2_X1 U21016 ( .A1(n17956), .A2(n17822), .ZN(n18187) );
  NOR2_X1 U21017 ( .A1(n17832), .A2(n18277), .ZN(n18189) );
  INV_X1 U21018 ( .A(n18189), .ZN(n17823) );
  AOI22_X1 U21019 ( .A1(n18132), .A2(n18187), .B1(n18012), .B2(n17823), .ZN(
        n17849) );
  NOR2_X1 U21020 ( .A1(n18447), .A2(n19056), .ZN(n17828) );
  INV_X1 U21021 ( .A(n17824), .ZN(n17825) );
  OAI22_X1 U21022 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17826), .B1(
        n17825), .B2(n17996), .ZN(n17827) );
  AOI211_X1 U21023 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(n17829), .A(
        n17828), .B(n17827), .ZN(n17835) );
  AOI21_X1 U21024 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17831), .A(
        n17830), .ZN(n18196) );
  INV_X1 U21025 ( .A(n18196), .ZN(n17833) );
  NOR2_X1 U21026 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17832), .ZN(
        n18185) );
  AOI22_X1 U21027 ( .A1(n18041), .A2(n17833), .B1(n17906), .B2(n18185), .ZN(
        n17834) );
  OAI211_X1 U21028 ( .C1(n17849), .C2(n17836), .A(n17835), .B(n17834), .ZN(
        P3_U2806) );
  NOR2_X1 U21029 ( .A1(n17986), .A2(n17852), .ZN(n17873) );
  NAND2_X1 U21030 ( .A1(n9993), .A2(n17873), .ZN(n17840) );
  NAND2_X1 U21031 ( .A1(n9652), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n18200) );
  OAI221_X1 U21032 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17840), .C1(
        n17839), .C2(n17838), .A(n18200), .ZN(n17846) );
  AOI22_X1 U21033 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18050), .B1(
        n17841), .B2(n17859), .ZN(n17842) );
  NAND2_X1 U21034 ( .A1(n17888), .A2(n17842), .ZN(n17843) );
  XNOR2_X1 U21035 ( .A(n17843), .B(n18190), .ZN(n18202) );
  OAI22_X1 U21036 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17844), .B1(
        n18202), .B2(n18052), .ZN(n17845) );
  AOI211_X1 U21037 ( .C1(n17980), .C2(n17847), .A(n17846), .B(n17845), .ZN(
        n17848) );
  OAI21_X1 U21038 ( .B1(n17849), .B2(n18190), .A(n17848), .ZN(P3_U2807) );
  NAND2_X1 U21039 ( .A1(n18151), .A2(n17906), .ZN(n17866) );
  NOR2_X1 U21040 ( .A1(n18447), .A2(n19052), .ZN(n17857) );
  OAI21_X1 U21041 ( .B1(n17850), .B2(n17977), .A(n18144), .ZN(n17851) );
  AOI21_X1 U21042 ( .B1(n18103), .B2(n17852), .A(n17851), .ZN(n17884) );
  OAI21_X1 U21043 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17881), .A(
        n17884), .ZN(n17871) );
  AOI22_X1 U21044 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17871), .B1(
        n17873), .B2(n17853), .ZN(n17854) );
  AOI21_X1 U21045 ( .B1(n17872), .B2(n17855), .A(n17854), .ZN(n17856) );
  AOI211_X1 U21046 ( .C1(n17858), .C2(n17980), .A(n17857), .B(n17856), .ZN(
        n17865) );
  AOI22_X1 U21047 ( .A1(n18132), .A2(n18286), .B1(n18012), .B2(n18277), .ZN(
        n17941) );
  OAI21_X1 U21048 ( .B1(n18151), .B2(n17887), .A(n17941), .ZN(n17877) );
  INV_X1 U21049 ( .A(n17859), .ZN(n17862) );
  INV_X1 U21050 ( .A(n17874), .ZN(n17861) );
  OAI221_X1 U21051 ( .B1(n17862), .B2(n17861), .C1(n17862), .C2(n17860), .A(
        n17888), .ZN(n17863) );
  XNOR2_X1 U21052 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17863), .ZN(
        n18203) );
  AOI22_X1 U21053 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17877), .B1(
        n18041), .B2(n18203), .ZN(n17864) );
  OAI211_X1 U21054 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n17866), .A(
        n17865), .B(n17864), .ZN(P3_U2808) );
  NAND2_X1 U21055 ( .A1(n18219), .A2(n17867), .ZN(n18223) );
  INV_X1 U21056 ( .A(n18217), .ZN(n18215) );
  NAND2_X1 U21057 ( .A1(n18215), .A2(n17906), .ZN(n17905) );
  AOI22_X1 U21058 ( .A1(n9652), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n17980), 
        .B2(n17868), .ZN(n17869) );
  INV_X1 U21059 ( .A(n17869), .ZN(n17870) );
  AOI221_X1 U21060 ( .B1(n17873), .B2(n17872), .C1(n17871), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17870), .ZN(n17879) );
  NOR3_X1 U21061 ( .A1(n17907), .A2(n18050), .A3(n17874), .ZN(n17899) );
  INV_X1 U21062 ( .A(n17915), .ZN(n17900) );
  AOI22_X1 U21063 ( .A1(n18219), .A2(n17899), .B1(n17900), .B2(n17875), .ZN(
        n17876) );
  XNOR2_X1 U21064 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17876), .ZN(
        n18216) );
  AOI22_X1 U21065 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17877), .B1(
        n18041), .B2(n18216), .ZN(n17878) );
  OAI211_X1 U21066 ( .C1(n18223), .C2(n17905), .A(n17879), .B(n17878), .ZN(
        P3_U2809) );
  NAND2_X1 U21067 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17880), .ZN(
        n18234) );
  AOI21_X1 U21068 ( .B1(n17882), .B2(n18858), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17883) );
  NAND2_X1 U21069 ( .A1(n9652), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n18232) );
  OAI21_X1 U21070 ( .B1(n17884), .B2(n17883), .A(n18232), .ZN(n17885) );
  AOI221_X1 U21071 ( .B1(n17980), .B2(n17886), .C1(n17920), .C2(n17886), .A(
        n17885), .ZN(n17891) );
  NOR2_X1 U21072 ( .A1(n18217), .A2(n18238), .ZN(n18227) );
  OAI21_X1 U21073 ( .B1(n17887), .B2(n18227), .A(n17941), .ZN(n17902) );
  OAI221_X1 U21074 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17914), 
        .C1(n18238), .C2(n17899), .A(n17888), .ZN(n17889) );
  XNOR2_X1 U21075 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17889), .ZN(
        n18230) );
  AOI22_X1 U21076 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17902), .B1(
        n18041), .B2(n18230), .ZN(n17890) );
  OAI211_X1 U21077 ( .C1(n18234), .C2(n17905), .A(n17891), .B(n17890), .ZN(
        P3_U2810) );
  AOI21_X1 U21078 ( .B1(n18103), .B2(n17893), .A(n18101), .ZN(n17922) );
  OAI21_X1 U21079 ( .B1(n17892), .B2(n17977), .A(n17922), .ZN(n17911) );
  NOR2_X1 U21080 ( .A1(n17986), .A2(n17893), .ZN(n17913) );
  OAI211_X1 U21081 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17913), .B(n17894), .ZN(n17896) );
  NAND2_X1 U21082 ( .A1(n9652), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17895) );
  OAI211_X1 U21083 ( .C1(n17996), .C2(n17897), .A(n17896), .B(n17895), .ZN(
        n17898) );
  AOI21_X1 U21084 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17911), .A(
        n17898), .ZN(n17904) );
  AOI21_X1 U21085 ( .B1(n17914), .B2(n17900), .A(n17899), .ZN(n17901) );
  XNOR2_X1 U21086 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n17901), .ZN(
        n18235) );
  AOI22_X1 U21087 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17902), .B1(
        n18041), .B2(n18235), .ZN(n17903) );
  OAI211_X1 U21088 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17905), .A(
        n17904), .B(n17903), .ZN(P3_U2811) );
  INV_X1 U21089 ( .A(n17906), .ZN(n17942) );
  NAND2_X1 U21090 ( .A1(n18247), .A2(n17907), .ZN(n18255) );
  INV_X1 U21091 ( .A(n17908), .ZN(n17909) );
  OAI22_X1 U21092 ( .A1(n18447), .A2(n19044), .B1(n17996), .B2(n17909), .ZN(
        n17910) );
  AOI221_X1 U21093 ( .B1(n17913), .B2(n17912), .C1(n17911), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17910), .ZN(n17918) );
  OAI21_X1 U21094 ( .B1(n18247), .B2(n17942), .A(n17941), .ZN(n17928) );
  AOI21_X1 U21095 ( .B1(n17952), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17914), .ZN(n17916) );
  XNOR2_X1 U21096 ( .A(n17916), .B(n17915), .ZN(n18244) );
  AOI22_X1 U21097 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17928), .B1(
        n18041), .B2(n18244), .ZN(n17917) );
  OAI211_X1 U21098 ( .C1(n17942), .C2(n18255), .A(n17918), .B(n17917), .ZN(
        P3_U2812) );
  NAND2_X1 U21099 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17926), .ZN(
        n18260) );
  AOI21_X1 U21100 ( .B1(n18858), .B2(n17919), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17923) );
  OAI22_X1 U21101 ( .A1(n17923), .A2(n17922), .B1(n18126), .B2(n17921), .ZN(
        n17924) );
  AOI21_X1 U21102 ( .B1(n9652), .B2(P3_REIP_REG_17__SCAN_IN), .A(n17924), .ZN(
        n17930) );
  OAI21_X1 U21103 ( .B1(n17927), .B2(n17926), .A(n17925), .ZN(n18256) );
  AOI22_X1 U21104 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17928), .B1(
        n18041), .B2(n18256), .ZN(n17929) );
  OAI211_X1 U21105 ( .C1(n17942), .C2(n18260), .A(n17930), .B(n17929), .ZN(
        P3_U2813) );
  NAND2_X1 U21106 ( .A1(n17952), .A2(n18331), .ZN(n18032) );
  OAI22_X1 U21107 ( .A1(n17952), .A2(n17931), .B1(n18032), .B2(n9856), .ZN(
        n17932) );
  XNOR2_X1 U21108 ( .A(n18272), .B(n17932), .ZN(n18269) );
  AOI21_X1 U21109 ( .B1(n18103), .B2(n17934), .A(n18101), .ZN(n17967) );
  OAI21_X1 U21110 ( .B1(n17933), .B2(n17977), .A(n17967), .ZN(n17945) );
  AOI22_X1 U21111 ( .A1(n9652), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17945), .ZN(n17937) );
  NOR2_X1 U21112 ( .A1(n17986), .A2(n17934), .ZN(n17947) );
  OAI211_X1 U21113 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17947), .B(n17935), .ZN(n17936) );
  OAI211_X1 U21114 ( .C1(n17996), .C2(n17938), .A(n17937), .B(n17936), .ZN(
        n17939) );
  AOI21_X1 U21115 ( .B1(n18041), .B2(n18269), .A(n17939), .ZN(n17940) );
  OAI221_X1 U21116 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17942), 
        .C1(n18272), .C2(n17941), .A(n17940), .ZN(P3_U2814) );
  NOR2_X1 U21117 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17969), .ZN(
        n18280) );
  NAND2_X1 U21118 ( .A1(n18012), .A2(n18277), .ZN(n17961) );
  OAI22_X1 U21119 ( .A1(n18447), .A2(n19038), .B1(n17996), .B2(n17943), .ZN(
        n17944) );
  AOI221_X1 U21120 ( .B1(n17947), .B2(n17946), .C1(n17945), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17944), .ZN(n17960) );
  NAND3_X1 U21121 ( .A1(n18322), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n17948), .ZN(n17954) );
  NAND2_X1 U21122 ( .A1(n18017), .A2(n18050), .ZN(n18033) );
  INV_X1 U21123 ( .A(n18033), .ZN(n17949) );
  NAND2_X1 U21124 ( .A1(n17950), .A2(n17949), .ZN(n17992) );
  AOI21_X1 U21125 ( .B1(n17952), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n17951), .ZN(n17953) );
  AOI221_X1 U21126 ( .B1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n17954), 
        .C1(n17983), .C2(n17992), .A(n17953), .ZN(n17955) );
  XNOR2_X1 U21127 ( .A(n17955), .B(n17957), .ZN(n18283) );
  NOR2_X1 U21128 ( .A1(n17956), .A2(n18149), .ZN(n17958) );
  NAND2_X1 U21129 ( .A1(n17962), .A2(n17957), .ZN(n18285) );
  AOI22_X1 U21130 ( .A1(n18041), .A2(n18283), .B1(n17958), .B2(n18285), .ZN(
        n17959) );
  OAI211_X1 U21131 ( .C1(n18280), .C2(n17961), .A(n17960), .B(n17959), .ZN(
        P3_U2815) );
  OAI21_X1 U21132 ( .B1(n17963), .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n17962), .ZN(n18306) );
  AOI21_X1 U21133 ( .B1(n17964), .B2(n18858), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17966) );
  OAI22_X1 U21134 ( .A1(n17967), .A2(n17966), .B1(n18126), .B2(n17965), .ZN(
        n17968) );
  AOI21_X1 U21135 ( .B1(n9652), .B2(P3_REIP_REG_14__SCAN_IN), .A(n17968), .ZN(
        n17975) );
  AOI21_X1 U21136 ( .B1(n18300), .B2(n17970), .A(n17969), .ZN(n18303) );
  NOR2_X1 U21137 ( .A1(n18291), .A2(n18032), .ZN(n17972) );
  NOR2_X1 U21138 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17992), .ZN(
        n17971) );
  AOI22_X1 U21139 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17972), .B1(
        n17971), .B2(n17983), .ZN(n17973) );
  XNOR2_X1 U21140 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n17973), .ZN(
        n18302) );
  AOI22_X1 U21141 ( .A1(n18012), .A2(n18303), .B1(n18041), .B2(n18302), .ZN(
        n17974) );
  OAI211_X1 U21142 ( .C1(n18149), .C2(n18306), .A(n17975), .B(n17974), .ZN(
        P3_U2816) );
  AOI21_X1 U21143 ( .B1(n18103), .B2(n17985), .A(n18101), .ZN(n17976) );
  OAI21_X1 U21144 ( .B1(n17978), .B2(n17977), .A(n17976), .ZN(n17998) );
  AOI22_X1 U21145 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17998), .B1(
        n17980), .B2(n17979), .ZN(n17991) );
  NOR2_X1 U21146 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18291), .ZN(
        n18310) );
  INV_X1 U21147 ( .A(n18044), .ZN(n18013) );
  OAI22_X1 U21148 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17992), .B1(
        n18032), .B2(n18291), .ZN(n17981) );
  XNOR2_X1 U21149 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17981), .ZN(
        n18321) );
  INV_X1 U21150 ( .A(n18291), .ZN(n18290) );
  NAND2_X1 U21151 ( .A1(n18290), .A2(n18329), .ZN(n18316) );
  NOR2_X1 U21152 ( .A1(n18291), .A2(n18011), .ZN(n18314) );
  INV_X1 U21153 ( .A(n18314), .ZN(n17982) );
  AOI22_X1 U21154 ( .A1(n18132), .A2(n18316), .B1(n18012), .B2(n17982), .ZN(
        n18001) );
  OAI22_X1 U21155 ( .A1(n18321), .A2(n18052), .B1(n18001), .B2(n17983), .ZN(
        n17984) );
  AOI21_X1 U21156 ( .B1(n18310), .B2(n18013), .A(n17984), .ZN(n17990) );
  NAND2_X1 U21157 ( .A1(n9652), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n17989) );
  NOR2_X1 U21158 ( .A1(n17986), .A2(n17985), .ZN(n18000) );
  OAI211_X1 U21159 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n18000), .B(n17987), .ZN(n17988) );
  NAND4_X1 U21160 ( .A1(n17991), .A2(n17990), .A3(n17989), .A4(n17988), .ZN(
        P3_U2817) );
  OR2_X1 U21161 ( .A1(n18334), .A2(n18032), .ZN(n18019) );
  OAI21_X1 U21162 ( .B1(n17993), .B2(n18019), .A(n17992), .ZN(n17994) );
  XNOR2_X1 U21163 ( .A(n17994), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18328) );
  INV_X1 U21164 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17999) );
  NAND2_X1 U21165 ( .A1(n9652), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18326) );
  OAI21_X1 U21166 ( .B1(n17996), .B2(n17995), .A(n18326), .ZN(n17997) );
  AOI221_X1 U21167 ( .B1(n18000), .B2(n17999), .C1(n17998), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n17997), .ZN(n18005) );
  NOR2_X1 U21168 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18044), .ZN(
        n18003) );
  INV_X1 U21169 ( .A(n18001), .ZN(n18002) );
  AOI22_X1 U21170 ( .A1(n18322), .A2(n18003), .B1(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18002), .ZN(n18004) );
  OAI211_X1 U21171 ( .C1(n18328), .C2(n18052), .A(n18005), .B(n18004), .ZN(
        P3_U2818) );
  OAI22_X1 U21172 ( .A1(n18334), .A2(n18032), .B1(n18027), .B2(n18033), .ZN(
        n18006) );
  XNOR2_X1 U21173 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18006), .ZN(
        n18344) );
  NOR3_X1 U21174 ( .A1(n18819), .A2(n18059), .A3(n18054), .ZN(n18036) );
  NAND2_X1 U21175 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n18036), .ZN(
        n18035) );
  NOR2_X1 U21176 ( .A1(n18022), .A2(n18035), .ZN(n18021) );
  NOR2_X1 U21177 ( .A1(n18009), .A2(n18021), .ZN(n18010) );
  NAND2_X1 U21178 ( .A1(n9652), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n18342) );
  OAI21_X1 U21179 ( .B1(n18126), .B2(n18007), .A(n18342), .ZN(n18008) );
  AOI221_X1 U21180 ( .B1(n18071), .B2(n18010), .C1(n18009), .C2(n18021), .A(
        n18008), .ZN(n18016) );
  INV_X1 U21181 ( .A(n18334), .ZN(n18026) );
  AOI22_X1 U21182 ( .A1(n18132), .A2(n18309), .B1(n18012), .B2(n18011), .ZN(
        n18043) );
  OAI21_X1 U21183 ( .B1(n18026), .B2(n18044), .A(n18043), .ZN(n18014) );
  NOR2_X1 U21184 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18334), .ZN(
        n18340) );
  AOI22_X1 U21185 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18014), .B1(
        n18340), .B2(n18013), .ZN(n18015) );
  OAI211_X1 U21186 ( .C1(n18344), .C2(n18052), .A(n18016), .B(n18015), .ZN(
        P3_U2819) );
  OAI221_X1 U21187 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18033), .C1(
        n18365), .C2(n18032), .A(n18338), .ZN(n18020) );
  NAND4_X1 U21188 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18017), .A3(
        n18365), .A4(n18050), .ZN(n18018) );
  NAND3_X1 U21189 ( .A1(n18020), .A2(n18019), .A3(n18018), .ZN(n18352) );
  INV_X1 U21190 ( .A(n18071), .ZN(n18140) );
  AOI211_X1 U21191 ( .C1(n18035), .C2(n18022), .A(n18140), .B(n18021), .ZN(
        n18024) );
  NOR2_X1 U21192 ( .A1(n18447), .A2(n19028), .ZN(n18023) );
  AOI211_X1 U21193 ( .C1(n18025), .C2(n18135), .A(n18024), .B(n18023), .ZN(
        n18031) );
  INV_X1 U21194 ( .A(n18043), .ZN(n18029) );
  NOR2_X1 U21195 ( .A1(n18026), .A2(n18044), .ZN(n18028) );
  AOI22_X1 U21196 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18029), .B1(
        n18028), .B2(n18027), .ZN(n18030) );
  OAI211_X1 U21197 ( .C1(n18052), .C2(n18352), .A(n18031), .B(n18030), .ZN(
        P3_U2820) );
  NAND2_X1 U21198 ( .A1(n18033), .A2(n18032), .ZN(n18034) );
  XNOR2_X1 U21199 ( .A(n18034), .B(n18365), .ZN(n18361) );
  NOR2_X1 U21200 ( .A1(n18447), .A2(n19026), .ZN(n18360) );
  INV_X1 U21201 ( .A(n18035), .ZN(n18039) );
  AOI21_X1 U21202 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18071), .A(
        n18036), .ZN(n18038) );
  OAI22_X1 U21203 ( .A1(n18039), .A2(n18038), .B1(n18126), .B2(n18037), .ZN(
        n18040) );
  AOI211_X1 U21204 ( .C1(n18041), .C2(n18361), .A(n18360), .B(n18040), .ZN(
        n18042) );
  OAI221_X1 U21205 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18044), .C1(
        n18365), .C2(n18043), .A(n18042), .ZN(P3_U2821) );
  OAI21_X1 U21206 ( .B1(n18046), .B2(n18045), .A(n18144), .ZN(n18060) );
  AOI22_X1 U21207 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18060), .B1(
        n18047), .B2(n18135), .ZN(n18058) );
  AOI21_X1 U21208 ( .B1(n18049), .B2(n18380), .A(n18048), .ZN(n18383) );
  AOI21_X1 U21209 ( .B1(n18050), .B2(n18382), .A(n9767), .ZN(n18389) );
  OAI22_X1 U21210 ( .A1(n18389), .A2(n18052), .B1(n18051), .B2(n18382), .ZN(
        n18053) );
  AOI21_X1 U21211 ( .B1(n18132), .B2(n18383), .A(n18053), .ZN(n18057) );
  NAND2_X1 U21212 ( .A1(n9652), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n18377) );
  OAI211_X1 U21213 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n18055), .A(
        n18858), .B(n18054), .ZN(n18056) );
  NAND4_X1 U21214 ( .A1(n18058), .A2(n18057), .A3(n18377), .A4(n18056), .ZN(
        P3_U2822) );
  NOR2_X1 U21215 ( .A1(n18819), .A2(n18059), .ZN(n18062) );
  NOR2_X1 U21216 ( .A1(n18447), .A2(n19022), .ZN(n18393) );
  AOI221_X1 U21217 ( .B1(n18062), .B2(n18061), .C1(n18060), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18393), .ZN(n18069) );
  NAND2_X1 U21218 ( .A1(n18064), .A2(n18063), .ZN(n18065) );
  XNOR2_X1 U21219 ( .A(n18065), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18395) );
  AOI21_X1 U21220 ( .B1(n18373), .B2(n18067), .A(n18066), .ZN(n18394) );
  AOI22_X1 U21221 ( .A1(n18132), .A2(n18395), .B1(n18136), .B2(n18394), .ZN(
        n18068) );
  OAI211_X1 U21222 ( .C1(n18126), .C2(n18070), .A(n18069), .B(n18068), .ZN(
        P3_U2823) );
  OAI21_X1 U21223 ( .B1(n18075), .B2(n18819), .A(n18071), .ZN(n18093) );
  AOI21_X1 U21224 ( .B1(n18074), .B2(n18073), .A(n18072), .ZN(n18403) );
  NOR2_X1 U21225 ( .A1(n18447), .A2(n19020), .ZN(n18402) );
  NOR3_X1 U21226 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18075), .A3(
        n18819), .ZN(n18076) );
  AOI211_X1 U21227 ( .C1(n18136), .C2(n18403), .A(n18402), .B(n18076), .ZN(
        n18081) );
  AOI21_X1 U21228 ( .B1(n18078), .B2(n18374), .A(n18077), .ZN(n18404) );
  AOI22_X1 U21229 ( .A1(n18132), .A2(n18404), .B1(n18079), .B2(n18135), .ZN(
        n18080) );
  OAI211_X1 U21230 ( .C1(n18082), .C2(n18093), .A(n18081), .B(n18080), .ZN(
        P3_U2824) );
  AOI21_X1 U21231 ( .B1(n18083), .B2(n18144), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18094) );
  OAI21_X1 U21232 ( .B1(n18085), .B2(n9805), .A(n18084), .ZN(n18086) );
  XNOR2_X1 U21233 ( .A(n18086), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18409) );
  AOI22_X1 U21234 ( .A1(n18136), .A2(n18409), .B1(n9652), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n18092) );
  AOI21_X1 U21235 ( .B1(n18089), .B2(n18088), .A(n18087), .ZN(n18408) );
  AOI22_X1 U21236 ( .A1(n18132), .A2(n18408), .B1(n18090), .B2(n18135), .ZN(
        n18091) );
  OAI211_X1 U21237 ( .C1(n18094), .C2(n18093), .A(n18092), .B(n18091), .ZN(
        P3_U2825) );
  AOI21_X1 U21238 ( .B1(n18097), .B2(n18096), .A(n18095), .ZN(n18418) );
  AOI22_X1 U21239 ( .A1(n18132), .A2(n18418), .B1(n9652), .B2(
        P3_REIP_REG_4__SCAN_IN), .ZN(n18108) );
  AOI21_X1 U21240 ( .B1(n18100), .B2(n18099), .A(n18098), .ZN(n18415) );
  AOI21_X1 U21241 ( .B1(n18103), .B2(n18102), .A(n18101), .ZN(n18119) );
  OAI22_X1 U21242 ( .A1(n18126), .A2(n18105), .B1(n18119), .B2(n18104), .ZN(
        n18106) );
  AOI21_X1 U21243 ( .B1(n18136), .B2(n18415), .A(n18106), .ZN(n18107) );
  OAI211_X1 U21244 ( .C1(n18819), .C2(n18109), .A(n18108), .B(n18107), .ZN(
        P3_U2826) );
  AOI21_X1 U21245 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18144), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18118) );
  AOI21_X1 U21246 ( .B1(n18112), .B2(n18111), .A(n18110), .ZN(n18427) );
  AOI22_X1 U21247 ( .A1(n18132), .A2(n18427), .B1(n9652), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n18117) );
  AOI21_X1 U21248 ( .B1(n18430), .B2(n18114), .A(n18113), .ZN(n18423) );
  AOI22_X1 U21249 ( .A1(n18136), .A2(n18423), .B1(n18115), .B2(n18135), .ZN(
        n18116) );
  OAI211_X1 U21250 ( .C1(n18119), .C2(n18118), .A(n18117), .B(n18116), .ZN(
        P3_U2827) );
  AOI21_X1 U21251 ( .B1(n18122), .B2(n18121), .A(n18120), .ZN(n18443) );
  NOR2_X1 U21252 ( .A1(n18447), .A2(n19012), .ZN(n18444) );
  XNOR2_X1 U21253 ( .A(n18124), .B(n18123), .ZN(n18440) );
  OAI22_X1 U21254 ( .A1(n18126), .A2(n18125), .B1(n18149), .B2(n18440), .ZN(
        n18127) );
  AOI211_X1 U21255 ( .C1(n18136), .C2(n18443), .A(n18444), .B(n18127), .ZN(
        n18128) );
  OAI221_X1 U21256 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18819), .C1(
        n18129), .C2(n18144), .A(n18128), .ZN(P3_U2828) );
  NOR2_X1 U21257 ( .A1(n18142), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18130) );
  XOR2_X1 U21258 ( .A(n18130), .B(n18134), .Z(n18458) );
  INV_X1 U21259 ( .A(n18458), .ZN(n18131) );
  AOI22_X1 U21260 ( .A1(n18132), .A2(n18131), .B1(n9652), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n18138) );
  AOI21_X1 U21261 ( .B1(n18134), .B2(n18141), .A(n18133), .ZN(n18452) );
  AOI22_X1 U21262 ( .A1(n18136), .A2(n18452), .B1(n18139), .B2(n18135), .ZN(
        n18137) );
  OAI211_X1 U21263 ( .C1(n18140), .C2(n18139), .A(n18138), .B(n18137), .ZN(
        P3_U2829) );
  OAI21_X1 U21264 ( .B1(n18142), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18141), .ZN(n18466) );
  INV_X1 U21265 ( .A(n18466), .ZN(n18150) );
  INV_X1 U21266 ( .A(n18143), .ZN(n19139) );
  OAI21_X1 U21267 ( .B1(n18145), .B2(n19139), .A(n18144), .ZN(n18146) );
  AOI22_X1 U21268 ( .A1(n9652), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18146), .ZN(n18147) );
  OAI221_X1 U21269 ( .B1(n18150), .B2(n18149), .C1(n18466), .C2(n18148), .A(
        n18147), .ZN(P3_U2830) );
  AOI22_X1 U21270 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18454), .B1(
        n9652), .B2(P3_REIP_REG_27__SCAN_IN), .ZN(n18164) );
  NAND2_X1 U21271 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18153) );
  INV_X1 U21272 ( .A(n18951), .ZN(n18928) );
  NAND2_X1 U21273 ( .A1(n18953), .A2(n18928), .ZN(n18369) );
  INV_X1 U21274 ( .A(n18369), .ZN(n18433) );
  INV_X1 U21275 ( .A(n18197), .ZN(n18152) );
  INV_X1 U21276 ( .A(n18151), .ZN(n18208) );
  OAI21_X1 U21277 ( .B1(n18208), .B2(n18261), .A(n18951), .ZN(n18209) );
  OAI221_X1 U21278 ( .B1(n18433), .B2(n18206), .C1(n18433), .C2(n18152), .A(
        n18209), .ZN(n18186) );
  AOI21_X1 U21279 ( .B1(n18153), .B2(n18369), .A(n18186), .ZN(n18177) );
  OAI22_X1 U21280 ( .A1(n18155), .A2(n18921), .B1(n18154), .B2(n18330), .ZN(
        n18156) );
  AOI211_X1 U21281 ( .C1(n18158), .C2(n18369), .A(n18157), .B(n18156), .ZN(
        n18159) );
  AOI21_X1 U21282 ( .B1(n18177), .B2(n18159), .A(n18459), .ZN(n18167) );
  NOR2_X1 U21283 ( .A1(n18459), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n18162) );
  NOR3_X1 U21284 ( .A1(n18204), .A2(n18160), .A3(n18197), .ZN(n18161) );
  OAI22_X1 U21285 ( .A1(n18167), .A2(n18162), .B1(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18161), .ZN(n18163) );
  OAI211_X1 U21286 ( .C1(n18165), .C2(n18388), .A(n18164), .B(n18163), .ZN(
        P3_U2835) );
  AOI22_X1 U21287 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18454), .B1(
        n9652), .B2(P3_REIP_REG_26__SCAN_IN), .ZN(n18169) );
  AOI22_X1 U21288 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18167), .B1(
        n18214), .B2(n18166), .ZN(n18168) );
  OAI211_X1 U21289 ( .C1(n18170), .C2(n18388), .A(n18169), .B(n18168), .ZN(
        P3_U2836) );
  AOI221_X1 U21290 ( .B1(n18172), .B2(n18931), .C1(n18246), .C2(n18931), .A(
        n18171), .ZN(n18176) );
  AOI21_X1 U21291 ( .B1(n18174), .B2(n18173), .A(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18175) );
  AOI211_X1 U21292 ( .C1(n18177), .C2(n18176), .A(n18175), .B(n18459), .ZN(
        n18178) );
  AOI211_X1 U21293 ( .C1(n18454), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n18179), .B(n18178), .ZN(n18183) );
  AOI22_X1 U21294 ( .A1(n18463), .A2(n18181), .B1(n18384), .B2(n18180), .ZN(
        n18182) );
  OAI211_X1 U21295 ( .C1(n18388), .C2(n18184), .A(n18183), .B(n18182), .ZN(
        P3_U2837) );
  AOI22_X1 U21296 ( .A1(n9652), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n18214), 
        .B2(n18185), .ZN(n18195) );
  INV_X1 U21297 ( .A(n18267), .ZN(n18375) );
  AOI211_X1 U21298 ( .C1(n18317), .C2(n18187), .A(n18454), .B(n18186), .ZN(
        n18188) );
  OAI21_X1 U21299 ( .B1(n18189), .B2(n18330), .A(n18188), .ZN(n18193) );
  NOR2_X1 U21300 ( .A1(n18190), .A2(n18193), .ZN(n18192) );
  AOI21_X1 U21301 ( .B1(n18192), .B2(n18191), .A(n9652), .ZN(n18198) );
  OAI211_X1 U21302 ( .C1(n18375), .C2(n18193), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n18198), .ZN(n18194) );
  OAI211_X1 U21303 ( .C1(n18196), .C2(n18388), .A(n18195), .B(n18194), .ZN(
        P3_U2838) );
  NOR2_X1 U21304 ( .A1(n18204), .A2(n18197), .ZN(n18199) );
  OAI221_X1 U21305 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18199), 
        .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n18460), .A(n18198), .ZN(
        n18201) );
  OAI211_X1 U21306 ( .C1(n18202), .C2(n18388), .A(n18201), .B(n18200), .ZN(
        P3_U2839) );
  AOI22_X1 U21307 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18454), .B1(
        n18362), .B2(n18203), .ZN(n18213) );
  NOR2_X1 U21308 ( .A1(n18204), .A2(n18208), .ZN(n18211) );
  INV_X1 U21309 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18210) );
  INV_X1 U21310 ( .A(n18265), .ZN(n18347) );
  NAND2_X1 U21311 ( .A1(n18921), .A2(n18330), .ZN(n18333) );
  INV_X1 U21312 ( .A(n18330), .ZN(n18278) );
  OAI221_X1 U21313 ( .B1(n18953), .B2(n18206), .C1(n18953), .C2(n18227), .A(
        n18266), .ZN(n18207) );
  OAI211_X1 U21314 ( .C1(n19052), .C2(n18447), .A(n18213), .B(n18212), .ZN(
        P3_U2840) );
  NAND2_X1 U21315 ( .A1(n18215), .A2(n18214), .ZN(n18239) );
  AOI22_X1 U21316 ( .A1(n9652), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18362), 
        .B2(n18216), .ZN(n18222) );
  NOR2_X1 U21317 ( .A1(n18931), .A2(n18951), .ZN(n18453) );
  OAI21_X1 U21318 ( .B1(n18217), .B2(n18261), .A(n18951), .ZN(n18224) );
  OAI211_X1 U21319 ( .C1(n18453), .C2(n18219), .A(n18224), .B(n18218), .ZN(
        n18220) );
  OAI211_X1 U21320 ( .C1(n18459), .C2(n18220), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18447), .ZN(n18221) );
  OAI211_X1 U21321 ( .C1(n18239), .C2(n18223), .A(n18222), .B(n18221), .ZN(
        P3_U2841) );
  NAND2_X1 U21322 ( .A1(n18238), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18229) );
  INV_X1 U21323 ( .A(n18333), .ZN(n18226) );
  OAI211_X1 U21324 ( .C1(n18227), .C2(n18226), .A(n18225), .B(n18224), .ZN(
        n18228) );
  OAI21_X1 U21325 ( .B1(n18459), .B2(n18228), .A(n18447), .ZN(n18237) );
  OAI21_X1 U21326 ( .B1(n18453), .B2(n18229), .A(n18237), .ZN(n18231) );
  AOI22_X1 U21327 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18231), .B1(
        n18362), .B2(n18230), .ZN(n18233) );
  OAI211_X1 U21328 ( .C1(n18239), .C2(n18234), .A(n18233), .B(n18232), .ZN(
        P3_U2842) );
  AOI22_X1 U21329 ( .A1(n9652), .A2(P3_REIP_REG_19__SCAN_IN), .B1(n18362), 
        .B2(n18235), .ZN(n18236) );
  OAI221_X1 U21330 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18239), 
        .C1(n18238), .C2(n18237), .A(n18236), .ZN(P3_U2843) );
  INV_X1 U21331 ( .A(n18240), .ZN(n18437) );
  AOI22_X1 U21332 ( .A1(n18931), .A2(n18431), .B1(n18416), .B2(n18437), .ZN(
        n18425) );
  NOR2_X1 U21333 ( .A1(n18425), .A2(n18459), .ZN(n18414) );
  NAND2_X1 U21334 ( .A1(n18241), .A2(n18414), .ZN(n18407) );
  NOR2_X1 U21335 ( .A1(n18275), .A2(n18407), .ZN(n18307) );
  AOI22_X1 U21336 ( .A1(n18243), .A2(n18307), .B1(n18391), .B2(n18242), .ZN(
        n18273) );
  AOI22_X1 U21337 ( .A1(n9652), .A2(P3_REIP_REG_18__SCAN_IN), .B1(n18362), 
        .B2(n18244), .ZN(n18254) );
  NOR2_X1 U21338 ( .A1(n18928), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18435) );
  NOR3_X1 U21339 ( .A1(n18435), .A2(n18245), .A3(n18272), .ZN(n18251) );
  AND2_X1 U21340 ( .A1(n18246), .A2(n18931), .ZN(n18249) );
  INV_X1 U21341 ( .A(n18247), .ZN(n18248) );
  OAI22_X1 U21342 ( .A1(n18931), .A2(n18333), .B1(n18249), .B2(n18248), .ZN(
        n18250) );
  OAI211_X1 U21343 ( .C1(n18433), .C2(n18251), .A(n18266), .B(n18250), .ZN(
        n18257) );
  OAI21_X1 U21344 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18433), .A(
        n18391), .ZN(n18252) );
  OAI211_X1 U21345 ( .C1(n18257), .C2(n18252), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B(n18447), .ZN(n18253) );
  OAI211_X1 U21346 ( .C1(n18273), .C2(n18255), .A(n18254), .B(n18253), .ZN(
        P3_U2844) );
  AOI22_X1 U21347 ( .A1(n9652), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n18362), 
        .B2(n18256), .ZN(n18259) );
  OAI221_X1 U21348 ( .B1(n18454), .B2(n18391), .C1(n18454), .C2(n18257), .A(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18258) );
  OAI211_X1 U21349 ( .C1(n18273), .C2(n18260), .A(n18259), .B(n18258), .ZN(
        P3_U2845) );
  NOR2_X1 U21350 ( .A1(n18953), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18355) );
  INV_X1 U21351 ( .A(n18261), .ZN(n18263) );
  NOR2_X1 U21352 ( .A1(n18262), .A2(n18949), .ZN(n18332) );
  AOI221_X1 U21353 ( .B1(n18367), .B2(n18312), .C1(n18370), .C2(n18312), .A(
        n18332), .ZN(n18357) );
  OAI211_X1 U21354 ( .C1(n18263), .C2(n18928), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n18357), .ZN(n18264) );
  AOI211_X1 U21355 ( .C1(n18265), .C2(n18274), .A(n18355), .B(n18264), .ZN(
        n18282) );
  OAI211_X1 U21356 ( .C1(n18267), .C2(n18282), .A(n18391), .B(n18266), .ZN(
        n18268) );
  NAND2_X1 U21357 ( .A1(n18447), .A2(n18268), .ZN(n18271) );
  AOI22_X1 U21358 ( .A1(n9652), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n18362), 
        .B2(n18269), .ZN(n18270) );
  OAI221_X1 U21359 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18273), 
        .C1(n18272), .C2(n18271), .A(n18270), .ZN(P3_U2846) );
  AOI22_X1 U21360 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18454), .B1(
        n9652), .B2(P3_REIP_REG_15__SCAN_IN), .ZN(n18289) );
  INV_X1 U21361 ( .A(n18274), .ZN(n18276) );
  NOR3_X1 U21362 ( .A1(n18425), .A2(n18275), .A3(n18390), .ZN(n18296) );
  AOI21_X1 U21363 ( .B1(n18276), .B2(n18296), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18281) );
  NAND2_X1 U21364 ( .A1(n18278), .A2(n18277), .ZN(n18279) );
  OAI22_X1 U21365 ( .A1(n18282), .A2(n18281), .B1(n18280), .B2(n18279), .ZN(
        n18284) );
  AOI22_X1 U21366 ( .A1(n18391), .A2(n18284), .B1(n18362), .B2(n18283), .ZN(
        n18288) );
  NAND3_X1 U21367 ( .A1(n18463), .A2(n18286), .A3(n18285), .ZN(n18287) );
  NAND3_X1 U21368 ( .A1(n18289), .A2(n18288), .A3(n18287), .ZN(P3_U2847) );
  OAI21_X1 U21369 ( .B1(n18290), .B2(n18949), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18295) );
  INV_X1 U21370 ( .A(n18336), .ZN(n18354) );
  AOI221_X1 U21371 ( .B1(n18291), .B2(n18951), .C1(n18354), .C2(n18951), .A(
        n18332), .ZN(n18313) );
  OAI21_X1 U21372 ( .B1(n18292), .B2(n18311), .A(n18312), .ZN(n18293) );
  OAI211_X1 U21373 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n18453), .A(
        n18313), .B(n18293), .ZN(n18294) );
  OAI21_X1 U21374 ( .B1(n18295), .B2(n18294), .A(n18391), .ZN(n18299) );
  NAND2_X1 U21375 ( .A1(n18297), .A2(n18296), .ZN(n18298) );
  AOI222_X1 U21376 ( .A1(n18300), .A2(n18299), .B1(n18300), .B2(n18298), .C1(
        n18299), .C2(n18460), .ZN(n18301) );
  AOI21_X1 U21377 ( .B1(n9652), .B2(P3_REIP_REG_14__SCAN_IN), .A(n18301), .ZN(
        n18305) );
  AOI22_X1 U21378 ( .A1(n18384), .A2(n18303), .B1(n18362), .B2(n18302), .ZN(
        n18304) );
  OAI211_X1 U21379 ( .C1(n18457), .C2(n18306), .A(n18305), .B(n18304), .ZN(
        P3_U2848) );
  AOI21_X1 U21380 ( .B1(n18384), .B2(n18331), .A(n18307), .ZN(n18308) );
  OAI21_X1 U21381 ( .B1(n18309), .B2(n18457), .A(n18308), .ZN(n18353) );
  AOI22_X1 U21382 ( .A1(n9652), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18310), 
        .B2(n18353), .ZN(n18320) );
  NAND2_X1 U21383 ( .A1(n18312), .A2(n18311), .ZN(n18346) );
  AOI21_X1 U21384 ( .B1(n18322), .B2(n18346), .A(n18347), .ZN(n18337) );
  OAI21_X1 U21385 ( .B1(n18314), .B2(n18330), .A(n18313), .ZN(n18315) );
  AOI211_X1 U21386 ( .C1(n18317), .C2(n18316), .A(n18337), .B(n18315), .ZN(
        n18324) );
  OAI211_X1 U21387 ( .C1(n18347), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18391), .B(n18324), .ZN(n18318) );
  NAND3_X1 U21388 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18447), .A3(
        n18318), .ZN(n18319) );
  OAI211_X1 U21389 ( .C1(n18321), .C2(n18388), .A(n18320), .B(n18319), .ZN(
        P3_U2849) );
  AOI22_X1 U21390 ( .A1(n18322), .A2(n18353), .B1(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18391), .ZN(n18323) );
  AOI21_X1 U21391 ( .B1(n18324), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18323), .ZN(n18325) );
  AOI21_X1 U21392 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18454), .A(
        n18325), .ZN(n18327) );
  OAI211_X1 U21393 ( .C1(n18328), .C2(n18388), .A(n18327), .B(n18326), .ZN(
        P3_U2850) );
  OAI22_X1 U21394 ( .A1(n18331), .A2(n18330), .B1(n18921), .B2(n18329), .ZN(
        n18359) );
  AOI211_X1 U21395 ( .C1(n18334), .C2(n18333), .A(n18332), .B(n18359), .ZN(
        n18335) );
  OAI221_X1 U21396 ( .B1(n18928), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(
        n18928), .C2(n18336), .A(n18335), .ZN(n18349) );
  AOI211_X1 U21397 ( .C1(n18951), .C2(n18338), .A(n18337), .B(n18349), .ZN(
        n18339) );
  OAI21_X1 U21398 ( .B1(n18339), .B2(n18459), .A(n18460), .ZN(n18341) );
  AOI22_X1 U21399 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18341), .B1(
        n18340), .B2(n18353), .ZN(n18343) );
  OAI211_X1 U21400 ( .C1(n18344), .C2(n18388), .A(n18343), .B(n18342), .ZN(
        P3_U2851) );
  NOR2_X1 U21401 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18365), .ZN(
        n18345) );
  AOI22_X1 U21402 ( .A1(n9652), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18345), 
        .B2(n18353), .ZN(n18351) );
  OAI211_X1 U21403 ( .C1(n18347), .C2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n18391), .B(n18346), .ZN(n18348) );
  OAI211_X1 U21404 ( .C1(n18349), .C2(n18348), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n18447), .ZN(n18350) );
  OAI211_X1 U21405 ( .C1(n18352), .C2(n18388), .A(n18351), .B(n18350), .ZN(
        P3_U2852) );
  INV_X1 U21406 ( .A(n18353), .ZN(n18366) );
  OAI21_X1 U21407 ( .B1(n18355), .B2(n18951), .A(n18354), .ZN(n18356) );
  NAND3_X1 U21408 ( .A1(n18357), .A2(n18460), .A3(n18356), .ZN(n18358) );
  OAI21_X1 U21409 ( .B1(n18359), .B2(n18358), .A(n18447), .ZN(n18364) );
  AOI21_X1 U21410 ( .B1(n18362), .B2(n18361), .A(n18360), .ZN(n18363) );
  OAI221_X1 U21411 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18366), .C1(
        n18365), .C2(n18364), .A(n18363), .ZN(P3_U2853) );
  NOR2_X1 U21412 ( .A1(n18367), .A2(n18407), .ZN(n18381) );
  INV_X1 U21413 ( .A(n18368), .ZN(n18372) );
  OAI21_X1 U21414 ( .B1(n18435), .B2(n18370), .A(n18369), .ZN(n18371) );
  OAI21_X1 U21415 ( .B1(n18372), .B2(n18949), .A(n18371), .ZN(n18400) );
  AOI211_X1 U21416 ( .C1(n18375), .C2(n18374), .A(n18373), .B(n18400), .ZN(
        n18399) );
  INV_X1 U21417 ( .A(n18376), .ZN(n18448) );
  OAI21_X1 U21418 ( .B1(n18399), .B2(n18448), .A(n18460), .ZN(n18379) );
  INV_X1 U21419 ( .A(n18377), .ZN(n18378) );
  AOI221_X1 U21420 ( .B1(n18381), .B2(n18380), .C1(n18379), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18378), .ZN(n18387) );
  INV_X1 U21421 ( .A(n18382), .ZN(n18385) );
  AOI22_X1 U21422 ( .A1(n18385), .A2(n18384), .B1(n18463), .B2(n18383), .ZN(
        n18386) );
  OAI211_X1 U21423 ( .C1(n18389), .C2(n18388), .A(n18387), .B(n18386), .ZN(
        P3_U2854) );
  NOR2_X1 U21424 ( .A1(n18425), .A2(n18390), .ZN(n18392) );
  OAI221_X1 U21425 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n18392), .A(n18391), .ZN(
        n18398) );
  AOI21_X1 U21426 ( .B1(n18454), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18393), .ZN(n18397) );
  INV_X1 U21427 ( .A(n18467), .ZN(n18451) );
  AOI22_X1 U21428 ( .A1(n18463), .A2(n18395), .B1(n18451), .B2(n18394), .ZN(
        n18396) );
  OAI211_X1 U21429 ( .C1(n18399), .C2(n18398), .A(n18397), .B(n18396), .ZN(
        P3_U2855) );
  INV_X1 U21430 ( .A(n18400), .ZN(n18401) );
  OAI21_X1 U21431 ( .B1(n18401), .B2(n18459), .A(n18460), .ZN(n18410) );
  AOI21_X1 U21432 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18410), .A(
        n18402), .ZN(n18406) );
  AOI22_X1 U21433 ( .A1(n18463), .A2(n18404), .B1(n18451), .B2(n18403), .ZN(
        n18405) );
  OAI211_X1 U21434 ( .C1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n18407), .A(
        n18406), .B(n18405), .ZN(P3_U2856) );
  AOI22_X1 U21435 ( .A1(n9652), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18463), .B2(
        n18408), .ZN(n18413) );
  AOI22_X1 U21436 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18410), .B1(
        n18451), .B2(n18409), .ZN(n18412) );
  NAND4_X1 U21437 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n18414), .A4(n10010), .ZN(
        n18411) );
  NAND3_X1 U21438 ( .A1(n18413), .A2(n18412), .A3(n18411), .ZN(P3_U2857) );
  NAND2_X1 U21439 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18414), .ZN(
        n18422) );
  AOI22_X1 U21440 ( .A1(n9652), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18451), .B2(
        n18415), .ZN(n18421) );
  OAI22_X1 U21441 ( .A1(n18416), .A2(n18433), .B1(n18949), .B2(n18431), .ZN(
        n18417) );
  NOR3_X1 U21442 ( .A1(n18435), .A2(n18430), .A3(n18417), .ZN(n18424) );
  OAI21_X1 U21443 ( .B1(n18424), .B2(n18448), .A(n18460), .ZN(n18419) );
  AOI22_X1 U21444 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18419), .B1(
        n18463), .B2(n18418), .ZN(n18420) );
  OAI211_X1 U21445 ( .C1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n18422), .A(
        n18421), .B(n18420), .ZN(P3_U2858) );
  AOI22_X1 U21446 ( .A1(n9652), .A2(P3_REIP_REG_3__SCAN_IN), .B1(n18451), .B2(
        n18423), .ZN(n18429) );
  AOI211_X1 U21447 ( .C1(n18425), .C2(n18430), .A(n18424), .B(n18459), .ZN(
        n18426) );
  AOI21_X1 U21448 ( .B1(n18427), .B2(n18463), .A(n18426), .ZN(n18428) );
  OAI211_X1 U21449 ( .C1(n18430), .C2(n18460), .A(n18429), .B(n18428), .ZN(
        P3_U2859) );
  NOR2_X1 U21450 ( .A1(n18949), .A2(n18431), .ZN(n18442) );
  NAND2_X1 U21451 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18432) );
  OAI22_X1 U21452 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18433), .B1(
        n18949), .B2(n18432), .ZN(n18434) );
  OAI21_X1 U21453 ( .B1(n18435), .B2(n18434), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18439) );
  NAND3_X1 U21454 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18437), .A3(
        n18436), .ZN(n18438) );
  OAI211_X1 U21455 ( .C1(n18440), .C2(n18921), .A(n18439), .B(n18438), .ZN(
        n18441) );
  AOI211_X1 U21456 ( .C1(n18443), .C2(n18919), .A(n18442), .B(n18441), .ZN(
        n18446) );
  AOI21_X1 U21457 ( .B1(n18454), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n18444), .ZN(n18445) );
  OAI21_X1 U21458 ( .B1(n18446), .B2(n18459), .A(n18445), .ZN(P3_U2860) );
  INV_X1 U21459 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19011) );
  NOR2_X1 U21460 ( .A1(n18447), .A2(n19011), .ZN(n18450) );
  AOI211_X1 U21461 ( .C1(n18953), .C2(n19112), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18448), .ZN(n18449) );
  AOI211_X1 U21462 ( .C1(n18452), .C2(n18451), .A(n18450), .B(n18449), .ZN(
        n18456) );
  NOR3_X1 U21463 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18453), .A3(
        n18459), .ZN(n18462) );
  OAI21_X1 U21464 ( .B1(n18454), .B2(n18462), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18455) );
  OAI211_X1 U21465 ( .C1(n18458), .C2(n18457), .A(n18456), .B(n18455), .ZN(
        P3_U2861) );
  AOI221_X1 U21466 ( .B1(n18953), .B2(n18460), .C1(n18459), .C2(n18460), .A(
        n19112), .ZN(n18461) );
  AOI211_X1 U21467 ( .C1(n18463), .C2(n18466), .A(n18462), .B(n18461), .ZN(
        n18465) );
  NAND2_X1 U21468 ( .A1(n9652), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n18464) );
  OAI211_X1 U21469 ( .C1(n18467), .C2(n18466), .A(n18465), .B(n18464), .ZN(
        P3_U2862) );
  AOI21_X1 U21470 ( .B1(n18470), .B2(n18469), .A(n18468), .ZN(n18980) );
  OAI21_X1 U21471 ( .B1(n18980), .B2(n18516), .A(n18475), .ZN(n18471) );
  OAI221_X1 U21472 ( .B1(n18957), .B2(n19130), .C1(n18957), .C2(n18475), .A(
        n18471), .ZN(P3_U2863) );
  INV_X1 U21473 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18967) );
  NOR2_X1 U21474 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18967), .ZN(
        n18717) );
  NOR2_X1 U21475 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18964), .ZN(
        n18649) );
  NOR2_X1 U21476 ( .A1(n18717), .A2(n18649), .ZN(n18473) );
  OAI22_X1 U21477 ( .A1(n18474), .A2(n18967), .B1(n18473), .B2(n18472), .ZN(
        P3_U2866) );
  NOR2_X1 U21478 ( .A1(n18968), .A2(n18475), .ZN(P3_U2867) );
  NAND2_X1 U21479 ( .A1(n18858), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18796) );
  NOR2_X1 U21480 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18959), .ZN(
        n18716) );
  NAND3_X1 U21481 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n18716), .ZN(n18825) );
  NAND3_X1 U21482 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n18959), .ZN(n18791) );
  NOR2_X2 U21483 ( .A1(n18957), .A2(n18791), .ZN(n18885) );
  NOR2_X2 U21484 ( .A1(n18476), .A2(n18819), .ZN(n18859) );
  AND2_X1 U21485 ( .A1(n18766), .A2(BUF2_REG_0__SCAN_IN), .ZN(n18853) );
  INV_X1 U21486 ( .A(n18647), .ZN(n18477) );
  NAND2_X1 U21487 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18477), .ZN(
        n18851) );
  NOR2_X2 U21488 ( .A1(n18957), .A2(n18851), .ZN(n18908) );
  NAND2_X1 U21489 ( .A1(n18959), .A2(n18957), .ZN(n18960) );
  NAND2_X1 U21490 ( .A1(n18964), .A2(n18967), .ZN(n18556) );
  NOR2_X2 U21491 ( .A1(n18960), .A2(n18556), .ZN(n18577) );
  NOR2_X1 U21492 ( .A1(n18908), .A2(n18577), .ZN(n18536) );
  NOR2_X1 U21493 ( .A1(n18852), .A2(n18536), .ZN(n18510) );
  AOI22_X1 U21494 ( .A1(n18885), .A2(n18859), .B1(n18853), .B2(n18510), .ZN(
        n18484) );
  INV_X1 U21495 ( .A(n18885), .ZN(n18913) );
  AOI21_X1 U21496 ( .B1(n18825), .B2(n18913), .A(n18558), .ZN(n18822) );
  AOI211_X1 U21497 ( .C1(P3_STATE2_REG_3__SCAN_IN), .C2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18536), .B(n18558), .ZN(
        n18478) );
  AOI21_X1 U21498 ( .B1(n18822), .B2(n18535), .A(n18478), .ZN(n18513) );
  INV_X1 U21499 ( .A(n18479), .ZN(n18480) );
  NAND2_X1 U21500 ( .A1(n18481), .A2(n18480), .ZN(n18511) );
  NOR2_X1 U21501 ( .A1(n18482), .A2(n18511), .ZN(n18793) );
  AOI22_X1 U21502 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18513), .B1(
        n18577), .B2(n18793), .ZN(n18483) );
  OAI211_X1 U21503 ( .C1(n18796), .C2(n18825), .A(n18484), .B(n18483), .ZN(
        P3_U2868) );
  NAND2_X1 U21504 ( .A1(n18858), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18869) );
  NOR2_X1 U21505 ( .A1(n18485), .A2(n18819), .ZN(n18865) );
  AND2_X1 U21506 ( .A1(n18766), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18864) );
  AOI22_X1 U21507 ( .A1(n18885), .A2(n18865), .B1(n18510), .B2(n18864), .ZN(
        n18487) );
  NOR2_X2 U21508 ( .A1(n19136), .A2(n18511), .ZN(n18866) );
  AOI22_X1 U21509 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18513), .B1(
        n18577), .B2(n18866), .ZN(n18486) );
  OAI211_X1 U21510 ( .C1(n18825), .C2(n18869), .A(n18487), .B(n18486), .ZN(
        P3_U2869) );
  NAND2_X1 U21511 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18858), .ZN(n18831) );
  NAND2_X1 U21512 ( .A1(n18858), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18875) );
  INV_X1 U21513 ( .A(n18875), .ZN(n18828) );
  NOR2_X2 U21514 ( .A1(n18558), .A2(n18488), .ZN(n18870) );
  AOI22_X1 U21515 ( .A1(n18847), .A2(n18828), .B1(n18510), .B2(n18870), .ZN(
        n18491) );
  NOR2_X2 U21516 ( .A1(n18489), .A2(n18511), .ZN(n18872) );
  AOI22_X1 U21517 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18513), .B1(
        n18577), .B2(n18872), .ZN(n18490) );
  OAI211_X1 U21518 ( .C1(n18913), .C2(n18831), .A(n18491), .B(n18490), .ZN(
        P3_U2870) );
  NAND2_X1 U21519 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18858), .ZN(n18776) );
  NAND2_X1 U21520 ( .A1(n18858), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18882) );
  INV_X1 U21521 ( .A(n18882), .ZN(n18773) );
  NOR2_X2 U21522 ( .A1(n18558), .A2(n18492), .ZN(n18876) );
  AOI22_X1 U21523 ( .A1(n18847), .A2(n18773), .B1(n18510), .B2(n18876), .ZN(
        n18495) );
  NOR2_X2 U21524 ( .A1(n18493), .A2(n18511), .ZN(n18879) );
  AOI22_X1 U21525 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18513), .B1(
        n18577), .B2(n18879), .ZN(n18494) );
  OAI211_X1 U21526 ( .C1(n18913), .C2(n18776), .A(n18495), .B(n18494), .ZN(
        P3_U2871) );
  NAND2_X1 U21527 ( .A1(n18858), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18809) );
  NAND2_X1 U21528 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18858), .ZN(n18890) );
  INV_X1 U21529 ( .A(n18890), .ZN(n18806) );
  NOR2_X2 U21530 ( .A1(n18558), .A2(n18496), .ZN(n18883) );
  AOI22_X1 U21531 ( .A1(n18885), .A2(n18806), .B1(n18510), .B2(n18883), .ZN(
        n18499) );
  NOR2_X2 U21532 ( .A1(n18497), .A2(n18511), .ZN(n18886) );
  AOI22_X1 U21533 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18513), .B1(
        n18577), .B2(n18886), .ZN(n18498) );
  OAI211_X1 U21534 ( .C1(n18825), .C2(n18809), .A(n18499), .B(n18498), .ZN(
        P3_U2872) );
  NAND2_X1 U21535 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18858), .ZN(n18839) );
  NAND2_X1 U21536 ( .A1(n18858), .A2(BUF2_REG_21__SCAN_IN), .ZN(n18896) );
  INV_X1 U21537 ( .A(n18896), .ZN(n18836) );
  NOR2_X2 U21538 ( .A1(n18558), .A2(n18500), .ZN(n18891) );
  AOI22_X1 U21539 ( .A1(n18847), .A2(n18836), .B1(n18510), .B2(n18891), .ZN(
        n18503) );
  NOR2_X2 U21540 ( .A1(n18501), .A2(n18511), .ZN(n18893) );
  AOI22_X1 U21541 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18513), .B1(
        n18577), .B2(n18893), .ZN(n18502) );
  OAI211_X1 U21542 ( .C1(n18913), .C2(n18839), .A(n18503), .B(n18502), .ZN(
        P3_U2873) );
  NAND2_X1 U21543 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18858), .ZN(n18844) );
  NOR2_X1 U21544 ( .A1(n18819), .A2(n18504), .ZN(n18840) );
  NOR2_X2 U21545 ( .A1(n18558), .A2(n18505), .ZN(n18897) );
  AOI22_X1 U21546 ( .A1(n18847), .A2(n18840), .B1(n18510), .B2(n18897), .ZN(
        n18508) );
  NOR2_X2 U21547 ( .A1(n18506), .A2(n18511), .ZN(n18899) );
  AOI22_X1 U21548 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18513), .B1(
        n18577), .B2(n18899), .ZN(n18507) );
  OAI211_X1 U21549 ( .C1(n18913), .C2(n18844), .A(n18508), .B(n18507), .ZN(
        P3_U2874) );
  NAND2_X1 U21550 ( .A1(n18858), .A2(BUF2_REG_31__SCAN_IN), .ZN(n18790) );
  NAND2_X1 U21551 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18858), .ZN(n18912) );
  INV_X1 U21552 ( .A(n18912), .ZN(n18786) );
  NOR2_X2 U21553 ( .A1(n18509), .A2(n18558), .ZN(n18904) );
  AOI22_X1 U21554 ( .A1(n18847), .A2(n18786), .B1(n18510), .B2(n18904), .ZN(
        n18515) );
  NOR2_X2 U21555 ( .A1(n18512), .A2(n18511), .ZN(n18907) );
  AOI22_X1 U21556 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18513), .B1(
        n18577), .B2(n18907), .ZN(n18514) );
  OAI211_X1 U21557 ( .C1(n18913), .C2(n18790), .A(n18515), .B(n18514), .ZN(
        P3_U2875) );
  INV_X1 U21558 ( .A(n18908), .ZN(n18863) );
  AOI22_X1 U21559 ( .A1(n18847), .A2(n18859), .B1(n18853), .B2(n18531), .ZN(
        n18518) );
  INV_X1 U21560 ( .A(n18851), .ZN(n18856) );
  INV_X1 U21561 ( .A(n18556), .ZN(n18559) );
  NOR2_X1 U21562 ( .A1(n18558), .A2(n18516), .ZN(n18855) );
  AND2_X1 U21563 ( .A1(n18959), .A2(n18855), .ZN(n18602) );
  AOI22_X1 U21564 ( .A1(n18858), .A2(n18856), .B1(n18559), .B2(n18602), .ZN(
        n18532) );
  NAND2_X1 U21565 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18959), .ZN(
        n18695) );
  NOR2_X2 U21566 ( .A1(n18556), .A2(n18695), .ZN(n18598) );
  AOI22_X1 U21567 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18532), .B1(
        n18793), .B2(n18598), .ZN(n18517) );
  OAI211_X1 U21568 ( .C1(n18796), .C2(n18863), .A(n18518), .B(n18517), .ZN(
        P3_U2876) );
  AOI22_X1 U21569 ( .A1(n18847), .A2(n18865), .B1(n18864), .B2(n18531), .ZN(
        n18520) );
  AOI22_X1 U21570 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18532), .B1(
        n18866), .B2(n18598), .ZN(n18519) );
  OAI211_X1 U21571 ( .C1(n18863), .C2(n18869), .A(n18520), .B(n18519), .ZN(
        P3_U2877) );
  AOI22_X1 U21572 ( .A1(n18908), .A2(n18828), .B1(n18870), .B2(n18531), .ZN(
        n18522) );
  AOI22_X1 U21573 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18532), .B1(
        n18872), .B2(n18598), .ZN(n18521) );
  OAI211_X1 U21574 ( .C1(n18825), .C2(n18831), .A(n18522), .B(n18521), .ZN(
        P3_U2878) );
  AOI22_X1 U21575 ( .A1(n18908), .A2(n18773), .B1(n18876), .B2(n18531), .ZN(
        n18524) );
  AOI22_X1 U21576 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18532), .B1(
        n18879), .B2(n18598), .ZN(n18523) );
  OAI211_X1 U21577 ( .C1(n18825), .C2(n18776), .A(n18524), .B(n18523), .ZN(
        P3_U2879) );
  INV_X1 U21578 ( .A(n18809), .ZN(n18884) );
  AOI22_X1 U21579 ( .A1(n18908), .A2(n18884), .B1(n18883), .B2(n18531), .ZN(
        n18526) );
  AOI22_X1 U21580 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18532), .B1(
        n18886), .B2(n18598), .ZN(n18525) );
  OAI211_X1 U21581 ( .C1(n18825), .C2(n18890), .A(n18526), .B(n18525), .ZN(
        P3_U2880) );
  INV_X1 U21582 ( .A(n18839), .ZN(n18892) );
  AOI22_X1 U21583 ( .A1(n18847), .A2(n18892), .B1(n18891), .B2(n18531), .ZN(
        n18528) );
  AOI22_X1 U21584 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18532), .B1(
        n18893), .B2(n18598), .ZN(n18527) );
  OAI211_X1 U21585 ( .C1(n18863), .C2(n18896), .A(n18528), .B(n18527), .ZN(
        P3_U2881) );
  INV_X1 U21586 ( .A(n18844), .ZN(n18898) );
  AOI22_X1 U21587 ( .A1(n18847), .A2(n18898), .B1(n18897), .B2(n18531), .ZN(
        n18530) );
  AOI22_X1 U21588 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18532), .B1(
        n18899), .B2(n18598), .ZN(n18529) );
  OAI211_X1 U21589 ( .C1(n18863), .C2(n18902), .A(n18530), .B(n18529), .ZN(
        P3_U2882) );
  AOI22_X1 U21590 ( .A1(n18847), .A2(n18906), .B1(n18904), .B2(n18531), .ZN(
        n18534) );
  AOI22_X1 U21591 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18532), .B1(
        n18907), .B2(n18598), .ZN(n18533) );
  OAI211_X1 U21592 ( .C1(n18863), .C2(n18912), .A(n18534), .B(n18533), .ZN(
        P3_U2883) );
  NAND2_X1 U21593 ( .A1(n18716), .A2(n18559), .ZN(n18617) );
  INV_X1 U21594 ( .A(n18796), .ZN(n18854) );
  NOR2_X1 U21595 ( .A1(n18598), .A2(n18621), .ZN(n18580) );
  NOR2_X1 U21596 ( .A1(n18852), .A2(n18580), .ZN(n18552) );
  AOI22_X1 U21597 ( .A1(n18854), .A2(n18577), .B1(n18853), .B2(n18552), .ZN(
        n18539) );
  INV_X1 U21598 ( .A(n18535), .ZN(n18763) );
  OAI21_X1 U21599 ( .B1(n18536), .B2(n18763), .A(n18580), .ZN(n18537) );
  OAI211_X1 U21600 ( .C1(n18621), .C2(n19086), .A(n18766), .B(n18537), .ZN(
        n18553) );
  AOI22_X1 U21601 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18553), .B1(
        n18908), .B2(n18859), .ZN(n18538) );
  OAI211_X1 U21602 ( .C1(n18862), .C2(n18617), .A(n18539), .B(n18538), .ZN(
        P3_U2884) );
  INV_X1 U21603 ( .A(n18577), .ZN(n18572) );
  AOI22_X1 U21604 ( .A1(n18908), .A2(n18865), .B1(n18864), .B2(n18552), .ZN(
        n18541) );
  AOI22_X1 U21605 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18553), .B1(
        n18866), .B2(n18621), .ZN(n18540) );
  OAI211_X1 U21606 ( .C1(n18572), .C2(n18869), .A(n18541), .B(n18540), .ZN(
        P3_U2885) );
  INV_X1 U21607 ( .A(n18831), .ZN(n18871) );
  AOI22_X1 U21608 ( .A1(n18908), .A2(n18871), .B1(n18870), .B2(n18552), .ZN(
        n18543) );
  AOI22_X1 U21609 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18553), .B1(
        n18872), .B2(n18621), .ZN(n18542) );
  OAI211_X1 U21610 ( .C1(n18572), .C2(n18875), .A(n18543), .B(n18542), .ZN(
        P3_U2886) );
  INV_X1 U21611 ( .A(n18776), .ZN(n18878) );
  AOI22_X1 U21612 ( .A1(n18908), .A2(n18878), .B1(n18876), .B2(n18552), .ZN(
        n18545) );
  AOI22_X1 U21613 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18553), .B1(
        n18879), .B2(n18621), .ZN(n18544) );
  OAI211_X1 U21614 ( .C1(n18572), .C2(n18882), .A(n18545), .B(n18544), .ZN(
        P3_U2887) );
  AOI22_X1 U21615 ( .A1(n18577), .A2(n18884), .B1(n18883), .B2(n18552), .ZN(
        n18547) );
  AOI22_X1 U21616 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18553), .B1(
        n18886), .B2(n18621), .ZN(n18546) );
  OAI211_X1 U21617 ( .C1(n18863), .C2(n18890), .A(n18547), .B(n18546), .ZN(
        P3_U2888) );
  AOI22_X1 U21618 ( .A1(n18577), .A2(n18836), .B1(n18891), .B2(n18552), .ZN(
        n18549) );
  AOI22_X1 U21619 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18553), .B1(
        n18893), .B2(n18621), .ZN(n18548) );
  OAI211_X1 U21620 ( .C1(n18863), .C2(n18839), .A(n18549), .B(n18548), .ZN(
        P3_U2889) );
  AOI22_X1 U21621 ( .A1(n18577), .A2(n18840), .B1(n18897), .B2(n18552), .ZN(
        n18551) );
  AOI22_X1 U21622 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18553), .B1(
        n18899), .B2(n18621), .ZN(n18550) );
  OAI211_X1 U21623 ( .C1(n18863), .C2(n18844), .A(n18551), .B(n18550), .ZN(
        P3_U2890) );
  AOI22_X1 U21624 ( .A1(n18577), .A2(n18786), .B1(n18904), .B2(n18552), .ZN(
        n18555) );
  AOI22_X1 U21625 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18553), .B1(
        n18907), .B2(n18621), .ZN(n18554) );
  OAI211_X1 U21626 ( .C1(n18863), .C2(n18790), .A(n18555), .B(n18554), .ZN(
        P3_U2891) );
  NOR2_X1 U21627 ( .A1(n18959), .A2(n18556), .ZN(n18603) );
  NAND2_X1 U21628 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18603), .ZN(
        n18646) );
  INV_X1 U21629 ( .A(n18603), .ZN(n18557) );
  NOR2_X1 U21630 ( .A1(n18852), .A2(n18557), .ZN(n18575) );
  AOI22_X1 U21631 ( .A1(n18577), .A2(n18859), .B1(n18853), .B2(n18575), .ZN(
        n18561) );
  AOI21_X1 U21632 ( .B1(n18959), .B2(n18763), .A(n18558), .ZN(n18648) );
  OAI211_X1 U21633 ( .C1(n18635), .C2(n19086), .A(n18559), .B(n18648), .ZN(
        n18576) );
  AOI22_X1 U21634 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18576), .B1(
        n18854), .B2(n18598), .ZN(n18560) );
  OAI211_X1 U21635 ( .C1(n18862), .C2(n18646), .A(n18561), .B(n18560), .ZN(
        P3_U2892) );
  INV_X1 U21636 ( .A(n18598), .ZN(n18594) );
  AOI22_X1 U21637 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18576), .B1(
        n18864), .B2(n18575), .ZN(n18563) );
  AOI22_X1 U21638 ( .A1(n18577), .A2(n18865), .B1(n18866), .B2(n18635), .ZN(
        n18562) );
  OAI211_X1 U21639 ( .C1(n18869), .C2(n18594), .A(n18563), .B(n18562), .ZN(
        P3_U2893) );
  AOI22_X1 U21640 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18576), .B1(
        n18870), .B2(n18575), .ZN(n18565) );
  AOI22_X1 U21641 ( .A1(n18577), .A2(n18871), .B1(n18872), .B2(n18635), .ZN(
        n18564) );
  OAI211_X1 U21642 ( .C1(n18875), .C2(n18594), .A(n18565), .B(n18564), .ZN(
        P3_U2894) );
  AOI22_X1 U21643 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18576), .B1(
        n18876), .B2(n18575), .ZN(n18567) );
  AOI22_X1 U21644 ( .A1(n18879), .A2(n18635), .B1(n18773), .B2(n18598), .ZN(
        n18566) );
  OAI211_X1 U21645 ( .C1(n18572), .C2(n18776), .A(n18567), .B(n18566), .ZN(
        P3_U2895) );
  AOI22_X1 U21646 ( .A1(n18577), .A2(n18806), .B1(n18883), .B2(n18575), .ZN(
        n18569) );
  AOI22_X1 U21647 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18576), .B1(
        n18886), .B2(n18635), .ZN(n18568) );
  OAI211_X1 U21648 ( .C1(n18809), .C2(n18594), .A(n18569), .B(n18568), .ZN(
        P3_U2896) );
  AOI22_X1 U21649 ( .A1(n18836), .A2(n18598), .B1(n18891), .B2(n18575), .ZN(
        n18571) );
  AOI22_X1 U21650 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18576), .B1(
        n18893), .B2(n18635), .ZN(n18570) );
  OAI211_X1 U21651 ( .C1(n18572), .C2(n18839), .A(n18571), .B(n18570), .ZN(
        P3_U2897) );
  AOI22_X1 U21652 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18576), .B1(
        n18897), .B2(n18575), .ZN(n18574) );
  AOI22_X1 U21653 ( .A1(n18577), .A2(n18898), .B1(n18899), .B2(n18635), .ZN(
        n18573) );
  OAI211_X1 U21654 ( .C1(n18902), .C2(n18594), .A(n18574), .B(n18573), .ZN(
        P3_U2898) );
  AOI22_X1 U21655 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18576), .B1(
        n18904), .B2(n18575), .ZN(n18579) );
  AOI22_X1 U21656 ( .A1(n18577), .A2(n18906), .B1(n18907), .B2(n18635), .ZN(
        n18578) );
  OAI211_X1 U21657 ( .C1(n18912), .C2(n18594), .A(n18579), .B(n18578), .ZN(
        P3_U2899) );
  INV_X1 U21658 ( .A(n18960), .ZN(n18671) );
  NAND2_X1 U21659 ( .A1(n18671), .A2(n18649), .ZN(n18665) );
  AOI21_X1 U21660 ( .B1(n18646), .B2(n18665), .A(n18852), .ZN(n18597) );
  AOI22_X1 U21661 ( .A1(n18854), .A2(n18621), .B1(n18853), .B2(n18597), .ZN(
        n18583) );
  AOI221_X1 U21662 ( .B1(n18580), .B2(n18646), .C1(n18763), .C2(n18646), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18581) );
  OAI21_X1 U21663 ( .B1(n18667), .B2(n18581), .A(n18766), .ZN(n18599) );
  AOI22_X1 U21664 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18599), .B1(
        n18859), .B2(n18598), .ZN(n18582) );
  OAI211_X1 U21665 ( .C1(n18862), .C2(n18665), .A(n18583), .B(n18582), .ZN(
        P3_U2900) );
  INV_X1 U21666 ( .A(n18865), .ZN(n18800) );
  INV_X1 U21667 ( .A(n18869), .ZN(n18797) );
  AOI22_X1 U21668 ( .A1(n18797), .A2(n18621), .B1(n18864), .B2(n18597), .ZN(
        n18585) );
  AOI22_X1 U21669 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18599), .B1(
        n18866), .B2(n18667), .ZN(n18584) );
  OAI211_X1 U21670 ( .C1(n18800), .C2(n18594), .A(n18585), .B(n18584), .ZN(
        P3_U2901) );
  AOI22_X1 U21671 ( .A1(n18871), .A2(n18598), .B1(n18870), .B2(n18597), .ZN(
        n18587) );
  AOI22_X1 U21672 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18599), .B1(
        n18872), .B2(n18667), .ZN(n18586) );
  OAI211_X1 U21673 ( .C1(n18875), .C2(n18617), .A(n18587), .B(n18586), .ZN(
        P3_U2902) );
  AOI22_X1 U21674 ( .A1(n18773), .A2(n18621), .B1(n18876), .B2(n18597), .ZN(
        n18589) );
  AOI22_X1 U21675 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18599), .B1(
        n18879), .B2(n18667), .ZN(n18588) );
  OAI211_X1 U21676 ( .C1(n18776), .C2(n18594), .A(n18589), .B(n18588), .ZN(
        P3_U2903) );
  AOI22_X1 U21677 ( .A1(n18806), .A2(n18598), .B1(n18883), .B2(n18597), .ZN(
        n18591) );
  AOI22_X1 U21678 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18599), .B1(
        n18886), .B2(n18667), .ZN(n18590) );
  OAI211_X1 U21679 ( .C1(n18809), .C2(n18617), .A(n18591), .B(n18590), .ZN(
        P3_U2904) );
  AOI22_X1 U21680 ( .A1(n18836), .A2(n18621), .B1(n18891), .B2(n18597), .ZN(
        n18593) );
  AOI22_X1 U21681 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18599), .B1(
        n18893), .B2(n18667), .ZN(n18592) );
  OAI211_X1 U21682 ( .C1(n18839), .C2(n18594), .A(n18593), .B(n18592), .ZN(
        P3_U2905) );
  AOI22_X1 U21683 ( .A1(n18898), .A2(n18598), .B1(n18897), .B2(n18597), .ZN(
        n18596) );
  AOI22_X1 U21684 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18599), .B1(
        n18899), .B2(n18667), .ZN(n18595) );
  OAI211_X1 U21685 ( .C1(n18902), .C2(n18617), .A(n18596), .B(n18595), .ZN(
        P3_U2906) );
  AOI22_X1 U21686 ( .A1(n18906), .A2(n18598), .B1(n18904), .B2(n18597), .ZN(
        n18601) );
  AOI22_X1 U21687 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18599), .B1(
        n18907), .B2(n18667), .ZN(n18600) );
  OAI211_X1 U21688 ( .C1(n18912), .C2(n18617), .A(n18601), .B(n18600), .ZN(
        P3_U2907) );
  INV_X1 U21689 ( .A(n18649), .ZN(n18604) );
  AOI22_X1 U21690 ( .A1(n18859), .A2(n18621), .B1(n18853), .B2(n18620), .ZN(
        n18606) );
  AOI22_X1 U21691 ( .A1(n18858), .A2(n18603), .B1(n18649), .B2(n18602), .ZN(
        n18622) );
  NOR2_X2 U21692 ( .A1(n18604), .A2(n18695), .ZN(n18686) );
  AOI22_X1 U21693 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18622), .B1(
        n18793), .B2(n18686), .ZN(n18605) );
  OAI211_X1 U21694 ( .C1(n18796), .C2(n18646), .A(n18606), .B(n18605), .ZN(
        P3_U2908) );
  AOI22_X1 U21695 ( .A1(n18797), .A2(n18635), .B1(n18864), .B2(n18620), .ZN(
        n18608) );
  AOI22_X1 U21696 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18622), .B1(
        n18866), .B2(n18686), .ZN(n18607) );
  OAI211_X1 U21697 ( .C1(n18800), .C2(n18617), .A(n18608), .B(n18607), .ZN(
        P3_U2909) );
  AOI22_X1 U21698 ( .A1(n18828), .A2(n18635), .B1(n18870), .B2(n18620), .ZN(
        n18610) );
  AOI22_X1 U21699 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18622), .B1(
        n18872), .B2(n18686), .ZN(n18609) );
  OAI211_X1 U21700 ( .C1(n18831), .C2(n18617), .A(n18610), .B(n18609), .ZN(
        P3_U2910) );
  AOI22_X1 U21701 ( .A1(n18773), .A2(n18635), .B1(n18876), .B2(n18620), .ZN(
        n18612) );
  AOI22_X1 U21702 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18622), .B1(
        n18879), .B2(n18686), .ZN(n18611) );
  OAI211_X1 U21703 ( .C1(n18776), .C2(n18617), .A(n18612), .B(n18611), .ZN(
        P3_U2911) );
  AOI22_X1 U21704 ( .A1(n18884), .A2(n18635), .B1(n18883), .B2(n18620), .ZN(
        n18614) );
  AOI22_X1 U21705 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18622), .B1(
        n18886), .B2(n18686), .ZN(n18613) );
  OAI211_X1 U21706 ( .C1(n18890), .C2(n18617), .A(n18614), .B(n18613), .ZN(
        P3_U2912) );
  AOI22_X1 U21707 ( .A1(n18836), .A2(n18635), .B1(n18891), .B2(n18620), .ZN(
        n18616) );
  AOI22_X1 U21708 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18622), .B1(
        n18893), .B2(n18686), .ZN(n18615) );
  OAI211_X1 U21709 ( .C1(n18839), .C2(n18617), .A(n18616), .B(n18615), .ZN(
        P3_U2913) );
  AOI22_X1 U21710 ( .A1(n18898), .A2(n18621), .B1(n18897), .B2(n18620), .ZN(
        n18619) );
  AOI22_X1 U21711 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18622), .B1(
        n18899), .B2(n18686), .ZN(n18618) );
  OAI211_X1 U21712 ( .C1(n18902), .C2(n18646), .A(n18619), .B(n18618), .ZN(
        P3_U2914) );
  AOI22_X1 U21713 ( .A1(n18906), .A2(n18621), .B1(n18904), .B2(n18620), .ZN(
        n18624) );
  AOI22_X1 U21714 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18622), .B1(
        n18907), .B2(n18686), .ZN(n18623) );
  OAI211_X1 U21715 ( .C1(n18912), .C2(n18646), .A(n18624), .B(n18623), .ZN(
        P3_U2915) );
  NAND2_X1 U21716 ( .A1(n18649), .A2(n18716), .ZN(n18710) );
  INV_X1 U21717 ( .A(n18710), .ZN(n18712) );
  NOR2_X1 U21718 ( .A1(n18686), .A2(n18712), .ZN(n18672) );
  NOR2_X1 U21719 ( .A1(n18852), .A2(n18672), .ZN(n18642) );
  AOI22_X1 U21720 ( .A1(n18854), .A2(n18667), .B1(n18853), .B2(n18642), .ZN(
        n18628) );
  NOR2_X1 U21721 ( .A1(n18635), .A2(n18667), .ZN(n18625) );
  OAI21_X1 U21722 ( .B1(n18625), .B2(n18763), .A(n18672), .ZN(n18626) );
  OAI211_X1 U21723 ( .C1(n18712), .C2(n19086), .A(n18766), .B(n18626), .ZN(
        n18643) );
  AOI22_X1 U21724 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18643), .B1(
        n18859), .B2(n18635), .ZN(n18627) );
  OAI211_X1 U21725 ( .C1(n18862), .C2(n18710), .A(n18628), .B(n18627), .ZN(
        P3_U2916) );
  AOI22_X1 U21726 ( .A1(n18865), .A2(n18635), .B1(n18864), .B2(n18642), .ZN(
        n18630) );
  AOI22_X1 U21727 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18643), .B1(
        n18866), .B2(n18712), .ZN(n18629) );
  OAI211_X1 U21728 ( .C1(n18869), .C2(n18665), .A(n18630), .B(n18629), .ZN(
        P3_U2917) );
  AOI22_X1 U21729 ( .A1(n18828), .A2(n18667), .B1(n18870), .B2(n18642), .ZN(
        n18632) );
  AOI22_X1 U21730 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18643), .B1(
        n18872), .B2(n18712), .ZN(n18631) );
  OAI211_X1 U21731 ( .C1(n18831), .C2(n18646), .A(n18632), .B(n18631), .ZN(
        P3_U2918) );
  AOI22_X1 U21732 ( .A1(n18773), .A2(n18667), .B1(n18876), .B2(n18642), .ZN(
        n18634) );
  AOI22_X1 U21733 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18643), .B1(
        n18879), .B2(n18712), .ZN(n18633) );
  OAI211_X1 U21734 ( .C1(n18776), .C2(n18646), .A(n18634), .B(n18633), .ZN(
        P3_U2919) );
  AOI22_X1 U21735 ( .A1(n18806), .A2(n18635), .B1(n18883), .B2(n18642), .ZN(
        n18637) );
  AOI22_X1 U21736 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18643), .B1(
        n18886), .B2(n18712), .ZN(n18636) );
  OAI211_X1 U21737 ( .C1(n18809), .C2(n18665), .A(n18637), .B(n18636), .ZN(
        P3_U2920) );
  AOI22_X1 U21738 ( .A1(n18836), .A2(n18667), .B1(n18891), .B2(n18642), .ZN(
        n18639) );
  AOI22_X1 U21739 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18643), .B1(
        n18893), .B2(n18712), .ZN(n18638) );
  OAI211_X1 U21740 ( .C1(n18839), .C2(n18646), .A(n18639), .B(n18638), .ZN(
        P3_U2921) );
  AOI22_X1 U21741 ( .A1(n18840), .A2(n18667), .B1(n18897), .B2(n18642), .ZN(
        n18641) );
  AOI22_X1 U21742 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18643), .B1(
        n18899), .B2(n18712), .ZN(n18640) );
  OAI211_X1 U21743 ( .C1(n18844), .C2(n18646), .A(n18641), .B(n18640), .ZN(
        P3_U2922) );
  AOI22_X1 U21744 ( .A1(n18786), .A2(n18667), .B1(n18904), .B2(n18642), .ZN(
        n18645) );
  AOI22_X1 U21745 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18643), .B1(
        n18907), .B2(n18712), .ZN(n18644) );
  OAI211_X1 U21746 ( .C1(n18790), .C2(n18646), .A(n18645), .B(n18644), .ZN(
        P3_U2923) );
  NOR2_X1 U21747 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18647), .ZN(
        n18694) );
  NAND2_X1 U21748 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18694), .ZN(
        n18734) );
  OAI211_X1 U21749 ( .C1(n18736), .C2(n19086), .A(n18649), .B(n18648), .ZN(
        n18668) );
  INV_X1 U21750 ( .A(n18694), .ZN(n18650) );
  NOR2_X1 U21751 ( .A1(n18852), .A2(n18650), .ZN(n18666) );
  AOI22_X1 U21752 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18668), .B1(
        n18853), .B2(n18666), .ZN(n18652) );
  AOI22_X1 U21753 ( .A1(n18854), .A2(n18686), .B1(n18859), .B2(n18667), .ZN(
        n18651) );
  OAI211_X1 U21754 ( .C1(n18862), .C2(n18734), .A(n18652), .B(n18651), .ZN(
        P3_U2924) );
  AOI22_X1 U21755 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18668), .B1(
        n18864), .B2(n18666), .ZN(n18654) );
  AOI22_X1 U21756 ( .A1(n18797), .A2(n18686), .B1(n18866), .B2(n18736), .ZN(
        n18653) );
  OAI211_X1 U21757 ( .C1(n18800), .C2(n18665), .A(n18654), .B(n18653), .ZN(
        P3_U2925) );
  AOI22_X1 U21758 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18668), .B1(
        n18870), .B2(n18666), .ZN(n18656) );
  AOI22_X1 U21759 ( .A1(n18872), .A2(n18736), .B1(n18828), .B2(n18686), .ZN(
        n18655) );
  OAI211_X1 U21760 ( .C1(n18831), .C2(n18665), .A(n18656), .B(n18655), .ZN(
        P3_U2926) );
  INV_X1 U21761 ( .A(n18686), .ZN(n18693) );
  AOI22_X1 U21762 ( .A1(n18878), .A2(n18667), .B1(n18876), .B2(n18666), .ZN(
        n18658) );
  AOI22_X1 U21763 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18668), .B1(
        n18879), .B2(n18736), .ZN(n18657) );
  OAI211_X1 U21764 ( .C1(n18882), .C2(n18693), .A(n18658), .B(n18657), .ZN(
        P3_U2927) );
  AOI22_X1 U21765 ( .A1(n18806), .A2(n18667), .B1(n18883), .B2(n18666), .ZN(
        n18660) );
  AOI22_X1 U21766 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18668), .B1(
        n18886), .B2(n18736), .ZN(n18659) );
  OAI211_X1 U21767 ( .C1(n18809), .C2(n18693), .A(n18660), .B(n18659), .ZN(
        P3_U2928) );
  AOI22_X1 U21768 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18668), .B1(
        n18891), .B2(n18666), .ZN(n18662) );
  AOI22_X1 U21769 ( .A1(n18892), .A2(n18667), .B1(n18893), .B2(n18736), .ZN(
        n18661) );
  OAI211_X1 U21770 ( .C1(n18896), .C2(n18693), .A(n18662), .B(n18661), .ZN(
        P3_U2929) );
  AOI22_X1 U21771 ( .A1(n18840), .A2(n18686), .B1(n18897), .B2(n18666), .ZN(
        n18664) );
  AOI22_X1 U21772 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18668), .B1(
        n18899), .B2(n18736), .ZN(n18663) );
  OAI211_X1 U21773 ( .C1(n18844), .C2(n18665), .A(n18664), .B(n18663), .ZN(
        P3_U2930) );
  AOI22_X1 U21774 ( .A1(n18906), .A2(n18667), .B1(n18904), .B2(n18666), .ZN(
        n18670) );
  AOI22_X1 U21775 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18668), .B1(
        n18907), .B2(n18736), .ZN(n18669) );
  OAI211_X1 U21776 ( .C1(n18912), .C2(n18693), .A(n18670), .B(n18669), .ZN(
        P3_U2931) );
  NAND2_X1 U21777 ( .A1(n18671), .A2(n18717), .ZN(n18755) );
  NOR2_X1 U21778 ( .A1(n18736), .A2(n18759), .ZN(n18718) );
  NOR2_X1 U21779 ( .A1(n18852), .A2(n18718), .ZN(n18689) );
  AOI22_X1 U21780 ( .A1(n18854), .A2(n18712), .B1(n18853), .B2(n18689), .ZN(
        n18675) );
  OAI21_X1 U21781 ( .B1(n18672), .B2(n18763), .A(n18718), .ZN(n18673) );
  OAI211_X1 U21782 ( .C1(n18759), .C2(n19086), .A(n18766), .B(n18673), .ZN(
        n18690) );
  AOI22_X1 U21783 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18690), .B1(
        n18859), .B2(n18686), .ZN(n18674) );
  OAI211_X1 U21784 ( .C1(n18862), .C2(n18755), .A(n18675), .B(n18674), .ZN(
        P3_U2932) );
  AOI22_X1 U21785 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18690), .B1(
        n18864), .B2(n18689), .ZN(n18677) );
  AOI22_X1 U21786 ( .A1(n18797), .A2(n18712), .B1(n18866), .B2(n18759), .ZN(
        n18676) );
  OAI211_X1 U21787 ( .C1(n18800), .C2(n18693), .A(n18677), .B(n18676), .ZN(
        P3_U2933) );
  AOI22_X1 U21788 ( .A1(n18871), .A2(n18686), .B1(n18870), .B2(n18689), .ZN(
        n18679) );
  AOI22_X1 U21789 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18690), .B1(
        n18872), .B2(n18759), .ZN(n18678) );
  OAI211_X1 U21790 ( .C1(n18875), .C2(n18710), .A(n18679), .B(n18678), .ZN(
        P3_U2934) );
  AOI22_X1 U21791 ( .A1(n18773), .A2(n18712), .B1(n18876), .B2(n18689), .ZN(
        n18681) );
  AOI22_X1 U21792 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18690), .B1(
        n18879), .B2(n18759), .ZN(n18680) );
  OAI211_X1 U21793 ( .C1(n18776), .C2(n18693), .A(n18681), .B(n18680), .ZN(
        P3_U2935) );
  AOI22_X1 U21794 ( .A1(n18884), .A2(n18712), .B1(n18883), .B2(n18689), .ZN(
        n18683) );
  AOI22_X1 U21795 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18690), .B1(
        n18886), .B2(n18759), .ZN(n18682) );
  OAI211_X1 U21796 ( .C1(n18890), .C2(n18693), .A(n18683), .B(n18682), .ZN(
        P3_U2936) );
  AOI22_X1 U21797 ( .A1(n18892), .A2(n18686), .B1(n18891), .B2(n18689), .ZN(
        n18685) );
  AOI22_X1 U21798 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18690), .B1(
        n18893), .B2(n18759), .ZN(n18684) );
  OAI211_X1 U21799 ( .C1(n18896), .C2(n18710), .A(n18685), .B(n18684), .ZN(
        P3_U2937) );
  AOI22_X1 U21800 ( .A1(n18898), .A2(n18686), .B1(n18897), .B2(n18689), .ZN(
        n18688) );
  AOI22_X1 U21801 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18690), .B1(
        n18899), .B2(n18759), .ZN(n18687) );
  OAI211_X1 U21802 ( .C1(n18902), .C2(n18710), .A(n18688), .B(n18687), .ZN(
        P3_U2938) );
  AOI22_X1 U21803 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18690), .B1(
        n18904), .B2(n18689), .ZN(n18692) );
  AOI22_X1 U21804 ( .A1(n18907), .A2(n18759), .B1(n18786), .B2(n18712), .ZN(
        n18691) );
  OAI211_X1 U21805 ( .C1(n18790), .C2(n18693), .A(n18692), .B(n18691), .ZN(
        P3_U2939) );
  INV_X1 U21806 ( .A(n18717), .ZN(n18740) );
  AOI22_X1 U21807 ( .A1(n18859), .A2(n18712), .B1(n18853), .B2(n18711), .ZN(
        n18697) );
  NOR2_X1 U21808 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18740), .ZN(
        n18742) );
  AOI22_X1 U21809 ( .A1(n18858), .A2(n18694), .B1(n18855), .B2(n18742), .ZN(
        n18713) );
  NOR2_X2 U21810 ( .A1(n18740), .A2(n18695), .ZN(n18781) );
  AOI22_X1 U21811 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18713), .B1(
        n18793), .B2(n18781), .ZN(n18696) );
  OAI211_X1 U21812 ( .C1(n18796), .C2(n18734), .A(n18697), .B(n18696), .ZN(
        P3_U2940) );
  AOI22_X1 U21813 ( .A1(n18865), .A2(n18712), .B1(n18864), .B2(n18711), .ZN(
        n18699) );
  AOI22_X1 U21814 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18713), .B1(
        n18866), .B2(n18781), .ZN(n18698) );
  OAI211_X1 U21815 ( .C1(n18869), .C2(n18734), .A(n18699), .B(n18698), .ZN(
        P3_U2941) );
  AOI22_X1 U21816 ( .A1(n18828), .A2(n18736), .B1(n18870), .B2(n18711), .ZN(
        n18701) );
  AOI22_X1 U21817 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18713), .B1(
        n18872), .B2(n18781), .ZN(n18700) );
  OAI211_X1 U21818 ( .C1(n18831), .C2(n18710), .A(n18701), .B(n18700), .ZN(
        P3_U2942) );
  AOI22_X1 U21819 ( .A1(n18773), .A2(n18736), .B1(n18876), .B2(n18711), .ZN(
        n18703) );
  AOI22_X1 U21820 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18713), .B1(
        n18879), .B2(n18781), .ZN(n18702) );
  OAI211_X1 U21821 ( .C1(n18776), .C2(n18710), .A(n18703), .B(n18702), .ZN(
        P3_U2943) );
  AOI22_X1 U21822 ( .A1(n18884), .A2(n18736), .B1(n18883), .B2(n18711), .ZN(
        n18705) );
  AOI22_X1 U21823 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18713), .B1(
        n18886), .B2(n18781), .ZN(n18704) );
  OAI211_X1 U21824 ( .C1(n18890), .C2(n18710), .A(n18705), .B(n18704), .ZN(
        P3_U2944) );
  AOI22_X1 U21825 ( .A1(n18836), .A2(n18736), .B1(n18891), .B2(n18711), .ZN(
        n18707) );
  AOI22_X1 U21826 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18713), .B1(
        n18893), .B2(n18781), .ZN(n18706) );
  OAI211_X1 U21827 ( .C1(n18839), .C2(n18710), .A(n18707), .B(n18706), .ZN(
        P3_U2945) );
  AOI22_X1 U21828 ( .A1(n18840), .A2(n18736), .B1(n18897), .B2(n18711), .ZN(
        n18709) );
  AOI22_X1 U21829 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18713), .B1(
        n18899), .B2(n18781), .ZN(n18708) );
  OAI211_X1 U21830 ( .C1(n18844), .C2(n18710), .A(n18709), .B(n18708), .ZN(
        P3_U2946) );
  AOI22_X1 U21831 ( .A1(n18906), .A2(n18712), .B1(n18904), .B2(n18711), .ZN(
        n18715) );
  AOI22_X1 U21832 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18713), .B1(
        n18907), .B2(n18781), .ZN(n18714) );
  OAI211_X1 U21833 ( .C1(n18912), .C2(n18734), .A(n18715), .B(n18714), .ZN(
        P3_U2947) );
  NAND2_X1 U21834 ( .A1(n18717), .A2(n18716), .ZN(n18803) );
  NOR2_X1 U21835 ( .A1(n18781), .A2(n18815), .ZN(n18764) );
  NOR2_X1 U21836 ( .A1(n18852), .A2(n18764), .ZN(n18735) );
  AOI22_X1 U21837 ( .A1(n18854), .A2(n18759), .B1(n18853), .B2(n18735), .ZN(
        n18721) );
  OAI21_X1 U21838 ( .B1(n18718), .B2(n18763), .A(n18764), .ZN(n18719) );
  OAI211_X1 U21839 ( .C1(n18815), .C2(n19086), .A(n18766), .B(n18719), .ZN(
        n18737) );
  AOI22_X1 U21840 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18737), .B1(
        n18859), .B2(n18736), .ZN(n18720) );
  OAI211_X1 U21841 ( .C1(n18862), .C2(n18803), .A(n18721), .B(n18720), .ZN(
        P3_U2948) );
  AOI22_X1 U21842 ( .A1(n18865), .A2(n18736), .B1(n18864), .B2(n18735), .ZN(
        n18723) );
  AOI22_X1 U21843 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18737), .B1(
        n18866), .B2(n18815), .ZN(n18722) );
  OAI211_X1 U21844 ( .C1(n18869), .C2(n18755), .A(n18723), .B(n18722), .ZN(
        P3_U2949) );
  AOI22_X1 U21845 ( .A1(n18828), .A2(n18759), .B1(n18870), .B2(n18735), .ZN(
        n18725) );
  AOI22_X1 U21846 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18737), .B1(
        n18872), .B2(n18815), .ZN(n18724) );
  OAI211_X1 U21847 ( .C1(n18831), .C2(n18734), .A(n18725), .B(n18724), .ZN(
        P3_U2950) );
  AOI22_X1 U21848 ( .A1(n18773), .A2(n18759), .B1(n18876), .B2(n18735), .ZN(
        n18727) );
  AOI22_X1 U21849 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18737), .B1(
        n18879), .B2(n18815), .ZN(n18726) );
  OAI211_X1 U21850 ( .C1(n18776), .C2(n18734), .A(n18727), .B(n18726), .ZN(
        P3_U2951) );
  AOI22_X1 U21851 ( .A1(n18806), .A2(n18736), .B1(n18883), .B2(n18735), .ZN(
        n18729) );
  AOI22_X1 U21852 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18737), .B1(
        n18886), .B2(n18815), .ZN(n18728) );
  OAI211_X1 U21853 ( .C1(n18809), .C2(n18755), .A(n18729), .B(n18728), .ZN(
        P3_U2952) );
  AOI22_X1 U21854 ( .A1(n18892), .A2(n18736), .B1(n18891), .B2(n18735), .ZN(
        n18731) );
  AOI22_X1 U21855 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18737), .B1(
        n18893), .B2(n18815), .ZN(n18730) );
  OAI211_X1 U21856 ( .C1(n18896), .C2(n18755), .A(n18731), .B(n18730), .ZN(
        P3_U2953) );
  AOI22_X1 U21857 ( .A1(n18840), .A2(n18759), .B1(n18897), .B2(n18735), .ZN(
        n18733) );
  AOI22_X1 U21858 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18737), .B1(
        n18899), .B2(n18815), .ZN(n18732) );
  OAI211_X1 U21859 ( .C1(n18844), .C2(n18734), .A(n18733), .B(n18732), .ZN(
        P3_U2954) );
  AOI22_X1 U21860 ( .A1(n18906), .A2(n18736), .B1(n18904), .B2(n18735), .ZN(
        n18739) );
  AOI22_X1 U21861 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18737), .B1(
        n18907), .B2(n18815), .ZN(n18738) );
  OAI211_X1 U21862 ( .C1(n18912), .C2(n18755), .A(n18739), .B(n18738), .ZN(
        P3_U2955) );
  NOR2_X1 U21863 ( .A1(n18959), .A2(n18740), .ZN(n18792) );
  NAND2_X1 U21864 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18792), .ZN(
        n18843) );
  INV_X1 U21865 ( .A(n18792), .ZN(n18741) );
  NOR2_X1 U21866 ( .A1(n18852), .A2(n18741), .ZN(n18758) );
  AOI22_X1 U21867 ( .A1(n18854), .A2(n18781), .B1(n18853), .B2(n18758), .ZN(
        n18744) );
  AOI22_X1 U21868 ( .A1(n18858), .A2(n18742), .B1(n18855), .B2(n18792), .ZN(
        n18760) );
  AOI22_X1 U21869 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18760), .B1(
        n18859), .B2(n18759), .ZN(n18743) );
  OAI211_X1 U21870 ( .C1(n18862), .C2(n18843), .A(n18744), .B(n18743), .ZN(
        P3_U2956) );
  AOI22_X1 U21871 ( .A1(n18797), .A2(n18781), .B1(n18864), .B2(n18758), .ZN(
        n18746) );
  INV_X1 U21872 ( .A(n18843), .ZN(n18846) );
  AOI22_X1 U21873 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18760), .B1(
        n18866), .B2(n18846), .ZN(n18745) );
  OAI211_X1 U21874 ( .C1(n18800), .C2(n18755), .A(n18746), .B(n18745), .ZN(
        P3_U2957) );
  INV_X1 U21875 ( .A(n18781), .ZN(n18789) );
  AOI22_X1 U21876 ( .A1(n18871), .A2(n18759), .B1(n18870), .B2(n18758), .ZN(
        n18748) );
  AOI22_X1 U21877 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18760), .B1(
        n18872), .B2(n18846), .ZN(n18747) );
  OAI211_X1 U21878 ( .C1(n18875), .C2(n18789), .A(n18748), .B(n18747), .ZN(
        P3_U2958) );
  AOI22_X1 U21879 ( .A1(n18878), .A2(n18759), .B1(n18876), .B2(n18758), .ZN(
        n18750) );
  AOI22_X1 U21880 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18760), .B1(
        n18879), .B2(n18846), .ZN(n18749) );
  OAI211_X1 U21881 ( .C1(n18882), .C2(n18789), .A(n18750), .B(n18749), .ZN(
        P3_U2959) );
  AOI22_X1 U21882 ( .A1(n18884), .A2(n18781), .B1(n18883), .B2(n18758), .ZN(
        n18752) );
  AOI22_X1 U21883 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18760), .B1(
        n18886), .B2(n18846), .ZN(n18751) );
  OAI211_X1 U21884 ( .C1(n18890), .C2(n18755), .A(n18752), .B(n18751), .ZN(
        P3_U2960) );
  AOI22_X1 U21885 ( .A1(n18836), .A2(n18781), .B1(n18891), .B2(n18758), .ZN(
        n18754) );
  AOI22_X1 U21886 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18760), .B1(
        n18893), .B2(n18846), .ZN(n18753) );
  OAI211_X1 U21887 ( .C1(n18839), .C2(n18755), .A(n18754), .B(n18753), .ZN(
        P3_U2961) );
  AOI22_X1 U21888 ( .A1(n18898), .A2(n18759), .B1(n18897), .B2(n18758), .ZN(
        n18757) );
  AOI22_X1 U21889 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18760), .B1(
        n18899), .B2(n18846), .ZN(n18756) );
  OAI211_X1 U21890 ( .C1(n18902), .C2(n18789), .A(n18757), .B(n18756), .ZN(
        P3_U2962) );
  AOI22_X1 U21891 ( .A1(n18906), .A2(n18759), .B1(n18904), .B2(n18758), .ZN(
        n18762) );
  AOI22_X1 U21892 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18760), .B1(
        n18907), .B2(n18846), .ZN(n18761) );
  OAI211_X1 U21893 ( .C1(n18912), .C2(n18789), .A(n18762), .B(n18761), .ZN(
        P3_U2963) );
  NOR2_X1 U21894 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18791), .ZN(
        n18877) );
  CLKBUF_X1 U21895 ( .A(n18877), .Z(n18905) );
  NOR2_X1 U21896 ( .A1(n18846), .A2(n18905), .ZN(n18820) );
  NOR2_X1 U21897 ( .A1(n18852), .A2(n18820), .ZN(n18784) );
  AOI22_X1 U21898 ( .A1(n18859), .A2(n18781), .B1(n18853), .B2(n18784), .ZN(
        n18768) );
  OAI21_X1 U21899 ( .B1(n18764), .B2(n18763), .A(n18820), .ZN(n18765) );
  OAI211_X1 U21900 ( .C1(n18905), .C2(n19086), .A(n18766), .B(n18765), .ZN(
        n18785) );
  AOI22_X1 U21901 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18785), .B1(
        n18793), .B2(n18905), .ZN(n18767) );
  OAI211_X1 U21902 ( .C1(n18796), .C2(n18803), .A(n18768), .B(n18767), .ZN(
        P3_U2964) );
  AOI22_X1 U21903 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18785), .B1(
        n18864), .B2(n18784), .ZN(n18770) );
  AOI22_X1 U21904 ( .A1(n18866), .A2(n18877), .B1(n18865), .B2(n18781), .ZN(
        n18769) );
  OAI211_X1 U21905 ( .C1(n18869), .C2(n18803), .A(n18770), .B(n18769), .ZN(
        P3_U2965) );
  AOI22_X1 U21906 ( .A1(n18828), .A2(n18815), .B1(n18870), .B2(n18784), .ZN(
        n18772) );
  AOI22_X1 U21907 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18785), .B1(
        n18872), .B2(n18877), .ZN(n18771) );
  OAI211_X1 U21908 ( .C1(n18831), .C2(n18789), .A(n18772), .B(n18771), .ZN(
        P3_U2966) );
  AOI22_X1 U21909 ( .A1(n18773), .A2(n18815), .B1(n18876), .B2(n18784), .ZN(
        n18775) );
  AOI22_X1 U21910 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18785), .B1(
        n18879), .B2(n18877), .ZN(n18774) );
  OAI211_X1 U21911 ( .C1(n18776), .C2(n18789), .A(n18775), .B(n18774), .ZN(
        P3_U2967) );
  AOI22_X1 U21912 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18785), .B1(
        n18883), .B2(n18784), .ZN(n18778) );
  AOI22_X1 U21913 ( .A1(n18886), .A2(n18905), .B1(n18806), .B2(n18781), .ZN(
        n18777) );
  OAI211_X1 U21914 ( .C1(n18809), .C2(n18803), .A(n18778), .B(n18777), .ZN(
        P3_U2968) );
  AOI22_X1 U21915 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18785), .B1(
        n18891), .B2(n18784), .ZN(n18780) );
  AOI22_X1 U21916 ( .A1(n18893), .A2(n18877), .B1(n18836), .B2(n18815), .ZN(
        n18779) );
  OAI211_X1 U21917 ( .C1(n18839), .C2(n18789), .A(n18780), .B(n18779), .ZN(
        P3_U2969) );
  AOI22_X1 U21918 ( .A1(n18898), .A2(n18781), .B1(n18897), .B2(n18784), .ZN(
        n18783) );
  AOI22_X1 U21919 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18785), .B1(
        n18899), .B2(n18905), .ZN(n18782) );
  OAI211_X1 U21920 ( .C1(n18902), .C2(n18803), .A(n18783), .B(n18782), .ZN(
        P3_U2970) );
  AOI22_X1 U21921 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18785), .B1(
        n18904), .B2(n18784), .ZN(n18788) );
  AOI22_X1 U21922 ( .A1(n18907), .A2(n18905), .B1(n18786), .B2(n18815), .ZN(
        n18787) );
  OAI211_X1 U21923 ( .C1(n18790), .C2(n18789), .A(n18788), .B(n18787), .ZN(
        P3_U2971) );
  NOR2_X1 U21924 ( .A1(n18852), .A2(n18791), .ZN(n18814) );
  AOI22_X1 U21925 ( .A1(n18859), .A2(n18815), .B1(n18853), .B2(n18814), .ZN(
        n18795) );
  INV_X1 U21926 ( .A(n18791), .ZN(n18857) );
  AOI22_X1 U21927 ( .A1(n18858), .A2(n18792), .B1(n18857), .B2(n18855), .ZN(
        n18816) );
  AOI22_X1 U21928 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18816), .B1(
        n18885), .B2(n18793), .ZN(n18794) );
  OAI211_X1 U21929 ( .C1(n18796), .C2(n18843), .A(n18795), .B(n18794), .ZN(
        P3_U2972) );
  AOI22_X1 U21930 ( .A1(n18797), .A2(n18846), .B1(n18864), .B2(n18814), .ZN(
        n18799) );
  AOI22_X1 U21931 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18816), .B1(
        n18885), .B2(n18866), .ZN(n18798) );
  OAI211_X1 U21932 ( .C1(n18800), .C2(n18803), .A(n18799), .B(n18798), .ZN(
        P3_U2973) );
  AOI22_X1 U21933 ( .A1(n18828), .A2(n18846), .B1(n18870), .B2(n18814), .ZN(
        n18802) );
  AOI22_X1 U21934 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18816), .B1(
        n18885), .B2(n18872), .ZN(n18801) );
  OAI211_X1 U21935 ( .C1(n18831), .C2(n18803), .A(n18802), .B(n18801), .ZN(
        P3_U2974) );
  AOI22_X1 U21936 ( .A1(n18878), .A2(n18815), .B1(n18876), .B2(n18814), .ZN(
        n18805) );
  AOI22_X1 U21937 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18816), .B1(
        n18885), .B2(n18879), .ZN(n18804) );
  OAI211_X1 U21938 ( .C1(n18882), .C2(n18843), .A(n18805), .B(n18804), .ZN(
        P3_U2975) );
  AOI22_X1 U21939 ( .A1(n18806), .A2(n18815), .B1(n18883), .B2(n18814), .ZN(
        n18808) );
  AOI22_X1 U21940 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18816), .B1(
        n18885), .B2(n18886), .ZN(n18807) );
  OAI211_X1 U21941 ( .C1(n18809), .C2(n18843), .A(n18808), .B(n18807), .ZN(
        P3_U2976) );
  AOI22_X1 U21942 ( .A1(n18892), .A2(n18815), .B1(n18891), .B2(n18814), .ZN(
        n18811) );
  AOI22_X1 U21943 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18816), .B1(
        n18885), .B2(n18893), .ZN(n18810) );
  OAI211_X1 U21944 ( .C1(n18896), .C2(n18843), .A(n18811), .B(n18810), .ZN(
        P3_U2977) );
  AOI22_X1 U21945 ( .A1(n18898), .A2(n18815), .B1(n18897), .B2(n18814), .ZN(
        n18813) );
  AOI22_X1 U21946 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18816), .B1(
        n18885), .B2(n18899), .ZN(n18812) );
  OAI211_X1 U21947 ( .C1(n18902), .C2(n18843), .A(n18813), .B(n18812), .ZN(
        P3_U2978) );
  AOI22_X1 U21948 ( .A1(n18906), .A2(n18815), .B1(n18904), .B2(n18814), .ZN(
        n18818) );
  AOI22_X1 U21949 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18816), .B1(
        n18885), .B2(n18907), .ZN(n18817) );
  OAI211_X1 U21950 ( .C1(n18912), .C2(n18843), .A(n18818), .B(n18817), .ZN(
        P3_U2979) );
  AOI21_X1 U21951 ( .B1(n18825), .B2(n18913), .A(n18852), .ZN(n18845) );
  AOI22_X1 U21952 ( .A1(n18854), .A2(n18905), .B1(n18853), .B2(n18845), .ZN(
        n18824) );
  NOR2_X1 U21953 ( .A1(n18820), .A2(n18819), .ZN(n18821) );
  OAI22_X1 U21954 ( .A1(n18847), .A2(n19086), .B1(n18822), .B2(n18821), .ZN(
        n18848) );
  AOI22_X1 U21955 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18848), .B1(
        n18859), .B2(n18846), .ZN(n18823) );
  OAI211_X1 U21956 ( .C1(n18825), .C2(n18862), .A(n18824), .B(n18823), .ZN(
        P3_U2980) );
  INV_X1 U21957 ( .A(n18877), .ZN(n18889) );
  AOI22_X1 U21958 ( .A1(n18865), .A2(n18846), .B1(n18864), .B2(n18845), .ZN(
        n18827) );
  AOI22_X1 U21959 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18848), .B1(
        n18847), .B2(n18866), .ZN(n18826) );
  OAI211_X1 U21960 ( .C1(n18869), .C2(n18889), .A(n18827), .B(n18826), .ZN(
        P3_U2981) );
  AOI22_X1 U21961 ( .A1(n18828), .A2(n18905), .B1(n18870), .B2(n18845), .ZN(
        n18830) );
  AOI22_X1 U21962 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18848), .B1(
        n18847), .B2(n18872), .ZN(n18829) );
  OAI211_X1 U21963 ( .C1(n18831), .C2(n18843), .A(n18830), .B(n18829), .ZN(
        P3_U2982) );
  AOI22_X1 U21964 ( .A1(n18878), .A2(n18846), .B1(n18876), .B2(n18845), .ZN(
        n18833) );
  AOI22_X1 U21965 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18848), .B1(
        n18847), .B2(n18879), .ZN(n18832) );
  OAI211_X1 U21966 ( .C1(n18882), .C2(n18889), .A(n18833), .B(n18832), .ZN(
        P3_U2983) );
  AOI22_X1 U21967 ( .A1(n18884), .A2(n18877), .B1(n18883), .B2(n18845), .ZN(
        n18835) );
  AOI22_X1 U21968 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18848), .B1(
        n18847), .B2(n18886), .ZN(n18834) );
  OAI211_X1 U21969 ( .C1(n18890), .C2(n18843), .A(n18835), .B(n18834), .ZN(
        P3_U2984) );
  AOI22_X1 U21970 ( .A1(n18836), .A2(n18877), .B1(n18891), .B2(n18845), .ZN(
        n18838) );
  AOI22_X1 U21971 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18848), .B1(
        n18847), .B2(n18893), .ZN(n18837) );
  OAI211_X1 U21972 ( .C1(n18839), .C2(n18843), .A(n18838), .B(n18837), .ZN(
        P3_U2985) );
  AOI22_X1 U21973 ( .A1(n18840), .A2(n18877), .B1(n18897), .B2(n18845), .ZN(
        n18842) );
  AOI22_X1 U21974 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18848), .B1(
        n18847), .B2(n18899), .ZN(n18841) );
  OAI211_X1 U21975 ( .C1(n18844), .C2(n18843), .A(n18842), .B(n18841), .ZN(
        P3_U2986) );
  AOI22_X1 U21976 ( .A1(n18906), .A2(n18846), .B1(n18904), .B2(n18845), .ZN(
        n18850) );
  AOI22_X1 U21977 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18848), .B1(
        n18847), .B2(n18907), .ZN(n18849) );
  OAI211_X1 U21978 ( .C1(n18912), .C2(n18889), .A(n18850), .B(n18849), .ZN(
        P3_U2987) );
  NOR2_X1 U21979 ( .A1(n18852), .A2(n18851), .ZN(n18903) );
  AOI22_X1 U21980 ( .A1(n18854), .A2(n18885), .B1(n18853), .B2(n18903), .ZN(
        n18861) );
  AOI22_X1 U21981 ( .A1(n18858), .A2(n18857), .B1(n18856), .B2(n18855), .ZN(
        n18909) );
  AOI22_X1 U21982 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18909), .B1(
        n18859), .B2(n18877), .ZN(n18860) );
  OAI211_X1 U21983 ( .C1(n18863), .C2(n18862), .A(n18861), .B(n18860), .ZN(
        P3_U2988) );
  AOI22_X1 U21984 ( .A1(n18865), .A2(n18877), .B1(n18864), .B2(n18903), .ZN(
        n18868) );
  AOI22_X1 U21985 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18909), .B1(
        n18908), .B2(n18866), .ZN(n18867) );
  OAI211_X1 U21986 ( .C1(n18913), .C2(n18869), .A(n18868), .B(n18867), .ZN(
        P3_U2989) );
  AOI22_X1 U21987 ( .A1(n18871), .A2(n18905), .B1(n18870), .B2(n18903), .ZN(
        n18874) );
  AOI22_X1 U21988 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18909), .B1(
        n18908), .B2(n18872), .ZN(n18873) );
  OAI211_X1 U21989 ( .C1(n18913), .C2(n18875), .A(n18874), .B(n18873), .ZN(
        P3_U2990) );
  AOI22_X1 U21990 ( .A1(n18878), .A2(n18877), .B1(n18876), .B2(n18903), .ZN(
        n18881) );
  AOI22_X1 U21991 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18909), .B1(
        n18908), .B2(n18879), .ZN(n18880) );
  OAI211_X1 U21992 ( .C1(n18913), .C2(n18882), .A(n18881), .B(n18880), .ZN(
        P3_U2991) );
  AOI22_X1 U21993 ( .A1(n18885), .A2(n18884), .B1(n18883), .B2(n18903), .ZN(
        n18888) );
  AOI22_X1 U21994 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18909), .B1(
        n18908), .B2(n18886), .ZN(n18887) );
  OAI211_X1 U21995 ( .C1(n18890), .C2(n18889), .A(n18888), .B(n18887), .ZN(
        P3_U2992) );
  AOI22_X1 U21996 ( .A1(n18892), .A2(n18905), .B1(n18891), .B2(n18903), .ZN(
        n18895) );
  AOI22_X1 U21997 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18909), .B1(
        n18908), .B2(n18893), .ZN(n18894) );
  OAI211_X1 U21998 ( .C1(n18913), .C2(n18896), .A(n18895), .B(n18894), .ZN(
        P3_U2993) );
  AOI22_X1 U21999 ( .A1(n18898), .A2(n18905), .B1(n18897), .B2(n18903), .ZN(
        n18901) );
  AOI22_X1 U22000 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18909), .B1(
        n18908), .B2(n18899), .ZN(n18900) );
  OAI211_X1 U22001 ( .C1(n18913), .C2(n18902), .A(n18901), .B(n18900), .ZN(
        P3_U2994) );
  AOI22_X1 U22002 ( .A1(n18906), .A2(n18905), .B1(n18904), .B2(n18903), .ZN(
        n18911) );
  AOI22_X1 U22003 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18909), .B1(
        n18908), .B2(n18907), .ZN(n18910) );
  OAI211_X1 U22004 ( .C1(n18913), .C2(n18912), .A(n18911), .B(n18910), .ZN(
        P3_U2995) );
  NAND2_X1 U22005 ( .A1(n18915), .A2(n18914), .ZN(n18916) );
  AOI22_X1 U22006 ( .A1(n18919), .A2(n18918), .B1(n18917), .B2(n18916), .ZN(
        n18920) );
  OAI221_X1 U22007 ( .B1(n18922), .B2(n18949), .C1(n18922), .C2(n18921), .A(
        n18920), .ZN(n19129) );
  OAI21_X1 U22008 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18923), .ZN(n18924) );
  OAI211_X1 U22009 ( .C1(n18950), .C2(n18926), .A(n18925), .B(n18924), .ZN(
        n18973) );
  NAND2_X1 U22010 ( .A1(n19102), .A2(n18944), .ZN(n18936) );
  OAI21_X1 U22011 ( .B1(n19115), .B2(n18928), .A(n18927), .ZN(n18942) );
  NOR2_X1 U22012 ( .A1(n18942), .A2(n18929), .ZN(n18954) );
  INV_X1 U22013 ( .A(n18954), .ZN(n18930) );
  AOI22_X1 U22014 ( .A1(n18931), .A2(n18936), .B1(n18937), .B2(n18930), .ZN(
        n18932) );
  NOR2_X1 U22015 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18932), .ZN(
        n19089) );
  OAI21_X1 U22016 ( .B1(n18935), .B2(n18934), .A(n18933), .ZN(n18945) );
  OAI21_X1 U22017 ( .B1(n18953), .B2(n18937), .A(n18936), .ZN(n18938) );
  AOI21_X1 U22018 ( .B1(n18939), .B2(n18945), .A(n18938), .ZN(n19090) );
  NAND2_X1 U22019 ( .A1(n18950), .A2(n19090), .ZN(n18940) );
  AOI22_X1 U22020 ( .A1(n18950), .A2(n19089), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18940), .ZN(n18971) );
  NAND2_X1 U22021 ( .A1(n19108), .A2(n9639), .ZN(n18941) );
  OAI221_X1 U22022 ( .B1(n19108), .B2(n19102), .C1(n18943), .C2(n18942), .A(
        n18941), .ZN(n18948) );
  AND2_X1 U22023 ( .A1(n18944), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n18946) );
  NAND2_X1 U22024 ( .A1(n18946), .A2(n18945), .ZN(n18947) );
  OAI211_X1 U22025 ( .C1(n19098), .C2(n18949), .A(n18948), .B(n18947), .ZN(
        n19100) );
  MUX2_X1 U22026 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n19100), .S(
        n18950), .Z(n18966) );
  INV_X1 U22027 ( .A(n18950), .ZN(n18962) );
  NOR2_X1 U22028 ( .A1(n18952), .A2(n18951), .ZN(n18956) );
  AOI22_X1 U22029 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18953), .B1(
        n18956), .B2(n19115), .ZN(n19110) );
  OAI22_X1 U22030 ( .A1(n18956), .A2(n18955), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18954), .ZN(n19106) );
  OR3_X1 U22031 ( .A1(n19110), .A2(n18959), .A3(n18957), .ZN(n18958) );
  AOI22_X1 U22032 ( .A1(n19110), .A2(n18959), .B1(n19106), .B2(n18958), .ZN(
        n18961) );
  OAI21_X1 U22033 ( .B1(n18962), .B2(n18961), .A(n18960), .ZN(n18965) );
  AND2_X1 U22034 ( .A1(n18966), .A2(n18965), .ZN(n18963) );
  OAI221_X1 U22035 ( .B1(n18966), .B2(n18965), .C1(n18964), .C2(n18963), .A(
        n18968), .ZN(n18970) );
  AOI21_X1 U22036 ( .B1(n18968), .B2(n18967), .A(n18966), .ZN(n18969) );
  AOI222_X1 U22037 ( .A1(n18971), .A2(n18970), .B1(n18971), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18970), .C2(n18969), .ZN(
        n18972) );
  NOR4_X1 U22038 ( .A1(n18974), .A2(n19129), .A3(n18973), .A4(n18972), .ZN(
        n18984) );
  AOI22_X1 U22039 ( .A1(n19109), .A2(n19139), .B1(n19002), .B2(n19133), .ZN(
        n18981) );
  NAND3_X1 U22040 ( .A1(n19136), .A2(n18976), .A3(n18975), .ZN(n18977) );
  NAND3_X1 U22041 ( .A1(n18984), .A2(n19131), .A3(n18977), .ZN(n19085) );
  NAND2_X1 U22042 ( .A1(n19002), .A2(n18978), .ZN(n18985) );
  NAND4_X1 U22043 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19085), .A3(n18979), 
        .A4(n18985), .ZN(n18988) );
  OAI22_X1 U22044 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18981), .B1(n18980), 
        .B2(n18988), .ZN(n18982) );
  OAI21_X1 U22045 ( .B1(n18984), .B2(n18983), .A(n18982), .ZN(P3_U2996) );
  NOR3_X1 U22046 ( .A1(n19095), .A2(n18986), .A3(n18985), .ZN(n18990) );
  AOI211_X1 U22047 ( .C1(n19002), .C2(n19133), .A(n16801), .B(n18990), .ZN(
        n18987) );
  OAI21_X1 U22048 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(n18988), .A(n18987), 
        .ZN(P3_U2997) );
  INV_X1 U22049 ( .A(n19084), .ZN(n18989) );
  NOR4_X1 U22050 ( .A1(n19139), .A2(n18991), .A3(n18990), .A4(n18989), .ZN(
        P3_U2998) );
  AND2_X1 U22051 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n19080), .ZN(
        P3_U2999) );
  AND2_X1 U22052 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18992), .ZN(
        P3_U3000) );
  AND2_X1 U22053 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18992), .ZN(
        P3_U3001) );
  AND2_X1 U22054 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n19080), .ZN(
        P3_U3002) );
  AND2_X1 U22055 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n19080), .ZN(
        P3_U3003) );
  AND2_X1 U22056 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n19080), .ZN(
        P3_U3004) );
  AND2_X1 U22057 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n19080), .ZN(
        P3_U3005) );
  AND2_X1 U22058 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n19080), .ZN(
        P3_U3006) );
  AND2_X1 U22059 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18992), .ZN(
        P3_U3007) );
  AND2_X1 U22060 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18992), .ZN(
        P3_U3008) );
  AND2_X1 U22061 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18992), .ZN(
        P3_U3009) );
  AND2_X1 U22062 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18992), .ZN(
        P3_U3010) );
  AND2_X1 U22063 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18992), .ZN(
        P3_U3011) );
  AND2_X1 U22064 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18992), .ZN(
        P3_U3012) );
  AND2_X1 U22065 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18992), .ZN(
        P3_U3013) );
  AND2_X1 U22066 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18992), .ZN(
        P3_U3014) );
  AND2_X1 U22067 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18992), .ZN(
        P3_U3015) );
  AND2_X1 U22068 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18992), .ZN(
        P3_U3016) );
  AND2_X1 U22069 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n19080), .ZN(
        P3_U3017) );
  AND2_X1 U22070 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n19080), .ZN(
        P3_U3018) );
  AND2_X1 U22071 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n19080), .ZN(
        P3_U3019) );
  AND2_X1 U22072 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n19080), .ZN(
        P3_U3020) );
  AND2_X1 U22073 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18992), .ZN(P3_U3021) );
  AND2_X1 U22074 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n19080), .ZN(P3_U3022) );
  AND2_X1 U22075 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n19080), .ZN(P3_U3023) );
  AND2_X1 U22076 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n19080), .ZN(P3_U3024) );
  AND2_X1 U22077 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n19080), .ZN(P3_U3025) );
  AND2_X1 U22078 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n19080), .ZN(P3_U3026) );
  AND2_X1 U22079 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n19080), .ZN(P3_U3027) );
  AND2_X1 U22080 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n19080), .ZN(P3_U3028) );
  NOR2_X1 U22081 ( .A1(n19009), .A2(n21016), .ZN(n19005) );
  INV_X1 U22082 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18993) );
  NOR2_X1 U22083 ( .A1(n19005), .A2(n18993), .ZN(n18999) );
  OAI21_X1 U22084 ( .B1(n18997), .B2(n21016), .A(n18999), .ZN(n18994) );
  AOI22_X1 U22085 ( .A1(n19007), .A2(n19009), .B1(n19144), .B2(n18994), .ZN(
        n18995) );
  NAND3_X1 U22086 ( .A1(NA), .A2(n19007), .A3(n18997), .ZN(n19001) );
  OAI211_X1 U22087 ( .C1(n19137), .C2(n18996), .A(n18995), .B(n19001), .ZN(
        P3_U3029) );
  NOR2_X1 U22088 ( .A1(n18997), .A2(n21016), .ZN(n18998) );
  AOI22_X1 U22089 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18999), .B1(n18998), 
        .B2(n19009), .ZN(n19000) );
  NAND2_X1 U22090 ( .A1(n19002), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19003) );
  NAND3_X1 U22091 ( .A1(n19000), .A2(n19134), .A3(n19003), .ZN(P3_U3030) );
  AOI22_X1 U22092 ( .A1(n19002), .A2(P3_STATE_REG_1__SCAN_IN), .B1(n19007), 
        .B2(n19001), .ZN(n19008) );
  OAI22_X1 U22093 ( .A1(NA), .A2(n19003), .B1(P3_STATE_REG_1__SCAN_IN), .B2(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19004) );
  OAI22_X1 U22094 ( .A1(n19005), .A2(n19004), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n19006) );
  OAI22_X1 U22095 ( .A1(n19008), .A2(n19009), .B1(n19007), .B2(n19006), .ZN(
        P3_U3031) );
  NAND2_X2 U22096 ( .A1(n19127), .A2(n19009), .ZN(n19068) );
  OAI222_X1 U22097 ( .A1(n19011), .A2(n19072), .B1(n19010), .B2(n19127), .C1(
        n19012), .C2(n19068), .ZN(P3_U3032) );
  INV_X1 U22098 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19014) );
  OAI222_X1 U22099 ( .A1(n19068), .A2(n19014), .B1(n19013), .B2(n19127), .C1(
        n19012), .C2(n19072), .ZN(P3_U3033) );
  OAI222_X1 U22100 ( .A1(n19068), .A2(n19016), .B1(n19015), .B2(n19127), .C1(
        n19014), .C2(n19072), .ZN(P3_U3034) );
  OAI222_X1 U22101 ( .A1(n19068), .A2(n19019), .B1(n19017), .B2(n19127), .C1(
        n19016), .C2(n19072), .ZN(P3_U3035) );
  OAI222_X1 U22102 ( .A1(n19019), .A2(n19072), .B1(n19018), .B2(n19127), .C1(
        n19020), .C2(n19068), .ZN(P3_U3036) );
  OAI222_X1 U22103 ( .A1(n19068), .A2(n19022), .B1(n19021), .B2(n19127), .C1(
        n19020), .C2(n19072), .ZN(P3_U3037) );
  OAI222_X1 U22104 ( .A1(n19068), .A2(n19024), .B1(n19023), .B2(n19127), .C1(
        n19022), .C2(n19072), .ZN(P3_U3038) );
  OAI222_X1 U22105 ( .A1(n19068), .A2(n19026), .B1(n19025), .B2(n19127), .C1(
        n19024), .C2(n19072), .ZN(P3_U3039) );
  OAI222_X1 U22106 ( .A1(n19068), .A2(n19028), .B1(n19027), .B2(n19127), .C1(
        n19026), .C2(n19072), .ZN(P3_U3040) );
  INV_X1 U22107 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19030) );
  OAI222_X1 U22108 ( .A1(n19068), .A2(n19030), .B1(n19029), .B2(n19127), .C1(
        n19028), .C2(n19072), .ZN(P3_U3041) );
  OAI222_X1 U22109 ( .A1(n19068), .A2(n19032), .B1(n19031), .B2(n19127), .C1(
        n19030), .C2(n19072), .ZN(P3_U3042) );
  OAI222_X1 U22110 ( .A1(n19068), .A2(n19034), .B1(n19033), .B2(n19127), .C1(
        n19032), .C2(n19072), .ZN(P3_U3043) );
  INV_X1 U22111 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19037) );
  OAI222_X1 U22112 ( .A1(n19068), .A2(n19037), .B1(n19035), .B2(n19127), .C1(
        n19034), .C2(n19072), .ZN(P3_U3044) );
  OAI222_X1 U22113 ( .A1(n19037), .A2(n19072), .B1(n19036), .B2(n19127), .C1(
        n19038), .C2(n19068), .ZN(P3_U3045) );
  OAI222_X1 U22114 ( .A1(n19068), .A2(n19040), .B1(n19039), .B2(n19127), .C1(
        n19038), .C2(n19072), .ZN(P3_U3046) );
  INV_X1 U22115 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19043) );
  OAI222_X1 U22116 ( .A1(n19068), .A2(n19043), .B1(n19041), .B2(n19127), .C1(
        n19040), .C2(n19072), .ZN(P3_U3047) );
  OAI222_X1 U22117 ( .A1(n19043), .A2(n19072), .B1(n19042), .B2(n19127), .C1(
        n19044), .C2(n19068), .ZN(P3_U3048) );
  INV_X1 U22118 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19046) );
  OAI222_X1 U22119 ( .A1(n19068), .A2(n19046), .B1(n19045), .B2(n19127), .C1(
        n19044), .C2(n19072), .ZN(P3_U3049) );
  OAI222_X1 U22120 ( .A1(n19068), .A2(n19048), .B1(n19047), .B2(n19127), .C1(
        n19046), .C2(n19072), .ZN(P3_U3050) );
  OAI222_X1 U22121 ( .A1(n19068), .A2(n19050), .B1(n19049), .B2(n19127), .C1(
        n19048), .C2(n19072), .ZN(P3_U3051) );
  OAI222_X1 U22122 ( .A1(n19068), .A2(n19052), .B1(n19051), .B2(n19127), .C1(
        n19050), .C2(n19072), .ZN(P3_U3052) );
  INV_X1 U22123 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19055) );
  OAI222_X1 U22124 ( .A1(n19068), .A2(n19055), .B1(n19053), .B2(n19127), .C1(
        n19052), .C2(n19072), .ZN(P3_U3053) );
  OAI222_X1 U22125 ( .A1(n19055), .A2(n19072), .B1(n19054), .B2(n19127), .C1(
        n19056), .C2(n19068), .ZN(P3_U3054) );
  OAI222_X1 U22126 ( .A1(n19068), .A2(n19058), .B1(n19057), .B2(n19127), .C1(
        n19056), .C2(n19072), .ZN(P3_U3055) );
  OAI222_X1 U22127 ( .A1(n19068), .A2(n19060), .B1(n19059), .B2(n19127), .C1(
        n19058), .C2(n19072), .ZN(P3_U3056) );
  OAI222_X1 U22128 ( .A1(n19068), .A2(n19062), .B1(n19061), .B2(n19127), .C1(
        n19060), .C2(n19072), .ZN(P3_U3057) );
  OAI222_X1 U22129 ( .A1(n19068), .A2(n19065), .B1(n19063), .B2(n19127), .C1(
        n19062), .C2(n19072), .ZN(P3_U3058) );
  OAI222_X1 U22130 ( .A1(n19065), .A2(n19072), .B1(n19064), .B2(n19127), .C1(
        n19066), .C2(n19068), .ZN(P3_U3059) );
  OAI222_X1 U22131 ( .A1(n19068), .A2(n19071), .B1(n19067), .B2(n19127), .C1(
        n19066), .C2(n19072), .ZN(P3_U3060) );
  INV_X1 U22132 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19070) );
  OAI222_X1 U22133 ( .A1(n19072), .A2(n19071), .B1(n19070), .B2(n19127), .C1(
        n19069), .C2(n19068), .ZN(P3_U3061) );
  INV_X1 U22134 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n19073) );
  AOI22_X1 U22135 ( .A1(n19127), .A2(n19074), .B1(n19073), .B2(n19144), .ZN(
        P3_U3274) );
  INV_X1 U22136 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19120) );
  INV_X1 U22137 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n19075) );
  AOI22_X1 U22138 ( .A1(n19127), .A2(n19120), .B1(n19075), .B2(n19144), .ZN(
        P3_U3275) );
  INV_X1 U22139 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n19076) );
  AOI22_X1 U22140 ( .A1(n19127), .A2(n19077), .B1(n19076), .B2(n19144), .ZN(
        P3_U3276) );
  INV_X1 U22141 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19123) );
  INV_X1 U22142 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n19078) );
  AOI22_X1 U22143 ( .A1(n19127), .A2(n19123), .B1(n19078), .B2(n19144), .ZN(
        P3_U3277) );
  INV_X1 U22144 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19118) );
  AOI21_X1 U22145 ( .B1(n19080), .B2(n19118), .A(n19079), .ZN(P3_U3280) );
  INV_X1 U22146 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19082) );
  OAI21_X1 U22147 ( .B1(n19083), .B2(n19082), .A(n19081), .ZN(P3_U3281) );
  OAI221_X1 U22148 ( .B1(n19086), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n19086), 
        .C2(n19085), .A(n19084), .ZN(P3_U3282) );
  INV_X1 U22149 ( .A(n19087), .ZN(n19088) );
  AOI22_X1 U22150 ( .A1(n19111), .A2(n19089), .B1(n19109), .B2(n19088), .ZN(
        n19094) );
  INV_X1 U22151 ( .A(n19090), .ZN(n19091) );
  AOI21_X1 U22152 ( .B1(n19111), .B2(n19091), .A(n19116), .ZN(n19093) );
  OAI22_X1 U22153 ( .A1(n19116), .A2(n19094), .B1(n19093), .B2(n19092), .ZN(
        P3_U3285) );
  NOR2_X1 U22154 ( .A1(n19095), .A2(n19112), .ZN(n19103) );
  AOI22_X1 U22155 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n19097), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n19096), .ZN(n19104) );
  INV_X1 U22156 ( .A(n19104), .ZN(n19099) );
  AOI222_X1 U22157 ( .A1(n19100), .A2(n19111), .B1(n19103), .B2(n19099), .C1(
        n19109), .C2(n19098), .ZN(n19101) );
  INV_X1 U22158 ( .A(n19116), .ZN(n19113) );
  AOI22_X1 U22159 ( .A1(n19116), .A2(n9639), .B1(n19101), .B2(n19113), .ZN(
        P3_U3288) );
  AOI222_X1 U22160 ( .A1(n19106), .A2(n19111), .B1(n19109), .B2(n19105), .C1(
        n19104), .C2(n19103), .ZN(n19107) );
  AOI22_X1 U22161 ( .A1(n19116), .A2(n19108), .B1(n19107), .B2(n19113), .ZN(
        P3_U3289) );
  AOI222_X1 U22162 ( .A1(n19112), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n19111), 
        .B2(n19110), .C1(n19115), .C2(n19109), .ZN(n19114) );
  AOI22_X1 U22163 ( .A1(n19116), .A2(n19115), .B1(n19114), .B2(n19113), .ZN(
        P3_U3290) );
  NOR3_X1 U22164 ( .A1(n19118), .A2(P3_REIP_REG_0__SCAN_IN), .A3(
        P3_REIP_REG_1__SCAN_IN), .ZN(n19117) );
  AOI221_X1 U22165 ( .B1(n19119), .B2(n19118), .C1(P3_REIP_REG_1__SCAN_IN), 
        .C2(P3_REIP_REG_0__SCAN_IN), .A(n19117), .ZN(n19121) );
  INV_X1 U22166 ( .A(n19125), .ZN(n19122) );
  AOI22_X1 U22167 ( .A1(n19125), .A2(n19121), .B1(n19120), .B2(n19122), .ZN(
        P3_U3292) );
  NOR2_X1 U22168 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .ZN(n19124) );
  AOI22_X1 U22169 ( .A1(n19125), .A2(n19124), .B1(n19123), .B2(n19122), .ZN(
        P3_U3293) );
  INV_X1 U22170 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19126) );
  AOI22_X1 U22171 ( .A1(n19127), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19126), 
        .B2(n19144), .ZN(P3_U3294) );
  MUX2_X1 U22172 ( .A(P3_MORE_REG_SCAN_IN), .B(n19129), .S(n19128), .Z(
        P3_U3295) );
  OAI21_X1 U22173 ( .B1(n19131), .B2(n19130), .A(n19147), .ZN(n19132) );
  AOI21_X1 U22174 ( .B1(n19133), .B2(n19137), .A(n19132), .ZN(n19143) );
  AOI21_X1 U22175 ( .B1(n19136), .B2(n19135), .A(n19134), .ZN(n19138) );
  OAI211_X1 U22176 ( .C1(n19138), .C2(n19148), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n19137), .ZN(n19140) );
  AOI21_X1 U22177 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19140), .A(n19139), 
        .ZN(n19142) );
  NAND2_X1 U22178 ( .A1(n19143), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n19141) );
  OAI21_X1 U22179 ( .B1(n19143), .B2(n19142), .A(n19141), .ZN(P3_U3296) );
  OAI22_X1 U22180 ( .A1(n19144), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n19127), .ZN(n19145) );
  INV_X1 U22181 ( .A(n19145), .ZN(P3_U3297) );
  OAI21_X1 U22182 ( .B1(n19146), .B2(P3_STATE2_REG_2__SCAN_IN), .A(n19147), 
        .ZN(n19151) );
  OAI22_X1 U22183 ( .A1(n19148), .A2(n19147), .B1(n19151), .B2(
        P3_READREQUEST_REG_SCAN_IN), .ZN(n19149) );
  INV_X1 U22184 ( .A(n19149), .ZN(P3_U3298) );
  OAI21_X1 U22185 ( .B1(n19151), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n19150), 
        .ZN(n19152) );
  INV_X1 U22186 ( .A(n19152), .ZN(P3_U3299) );
  AOI21_X1 U22187 ( .B1(P2_MEMORYFETCH_REG_SCAN_IN), .B2(n19154), .A(n19153), 
        .ZN(n19155) );
  OAI21_X1 U22188 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(n19868), .A(n19155), 
        .ZN(P2_U2814) );
  INV_X1 U22189 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n19157) );
  NAND2_X1 U22190 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19997), .ZN(n19990) );
  NAND2_X1 U22191 ( .A1(n19986), .A2(n19156), .ZN(n19987) );
  OAI21_X1 U22192 ( .B1(n19986), .B2(n19990), .A(n19987), .ZN(n20054) );
  OAI21_X1 U22193 ( .B1(n19986), .B2(n19157), .A(n19981), .ZN(P2_U2815) );
  INV_X1 U22194 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n19160) );
  NAND2_X1 U22195 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20089), .ZN(n19158) );
  OAI22_X1 U22196 ( .A1(n20111), .A2(n19160), .B1(n19159), .B2(n19158), .ZN(
        P2_U2816) );
  NAND2_X1 U22197 ( .A1(n20098), .A2(n19991), .ZN(n19984) );
  AOI21_X1 U22198 ( .B1(n19986), .B2(n19984), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n19161) );
  AOI21_X1 U22199 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n20034), .A(n19161), 
        .ZN(P2_U2817) );
  AOI21_X1 U22200 ( .B1(n19991), .B2(n20920), .A(n19981), .ZN(n20050) );
  INV_X1 U22201 ( .A(n20050), .ZN(n20052) );
  OAI21_X1 U22202 ( .B1(n20054), .B2(n19726), .A(n20052), .ZN(P2_U2818) );
  NOR4_X1 U22203 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19165) );
  NOR4_X1 U22204 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19164) );
  NOR4_X1 U22205 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19163) );
  NOR4_X1 U22206 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19162) );
  NAND4_X1 U22207 ( .A1(n19165), .A2(n19164), .A3(n19163), .A4(n19162), .ZN(
        n19171) );
  NOR4_X1 U22208 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19169) );
  AOI211_X1 U22209 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19168) );
  NOR4_X1 U22210 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19167) );
  NOR4_X1 U22211 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19166) );
  NAND4_X1 U22212 ( .A1(n19169), .A2(n19168), .A3(n19167), .A4(n19166), .ZN(
        n19170) );
  NOR2_X1 U22213 ( .A1(n19171), .A2(n19170), .ZN(n19178) );
  INV_X1 U22214 ( .A(n19178), .ZN(n19177) );
  NOR2_X1 U22215 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19177), .ZN(n19172) );
  INV_X1 U22216 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20049) );
  AOI22_X1 U22217 ( .A1(n19172), .A2(n10658), .B1(n19177), .B2(n20049), .ZN(
        P2_U2820) );
  INV_X1 U22218 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20053) );
  INV_X1 U22219 ( .A(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20051) );
  NAND3_X1 U22220 ( .A1(n10658), .A2(n20053), .A3(n20051), .ZN(n19176) );
  INV_X1 U22221 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20047) );
  AOI22_X1 U22222 ( .A1(n19172), .A2(n19176), .B1(n19177), .B2(n20047), .ZN(
        P2_U2821) );
  NAND2_X1 U22223 ( .A1(n19172), .A2(n20053), .ZN(n19175) );
  OAI21_X1 U22224 ( .B1(n10658), .B2(n10624), .A(n19178), .ZN(n19173) );
  OAI21_X1 U22225 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19178), .A(n19173), 
        .ZN(n19174) );
  OAI221_X1 U22226 ( .B1(n19175), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19175), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19174), .ZN(P2_U2822) );
  INV_X1 U22227 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20045) );
  OAI221_X1 U22228 ( .B1(n19178), .B2(n20045), .C1(n19177), .C2(n19176), .A(
        n19175), .ZN(P2_U2823) );
  AOI211_X1 U22229 ( .C1(n19186), .C2(n19180), .A(n19977), .B(n19179), .ZN(
        n19183) );
  OAI22_X1 U22230 ( .A1(n19303), .A2(n19181), .B1(n20020), .B2(n19301), .ZN(
        n19182) );
  AOI211_X1 U22231 ( .C1(n19308), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n19183), .B(n19182), .ZN(n19192) );
  NAND2_X1 U22232 ( .A1(n19184), .A2(n19324), .ZN(n19188) );
  INV_X1 U22233 ( .A(n19333), .ZN(n19185) );
  NAND2_X1 U22234 ( .A1(n19186), .A2(n19185), .ZN(n19187) );
  OAI211_X1 U22235 ( .C1(n19321), .C2(n19189), .A(n19188), .B(n19187), .ZN(
        n19190) );
  INV_X1 U22236 ( .A(n19190), .ZN(n19191) );
  OAI211_X1 U22237 ( .C1(n19193), .C2(n19320), .A(n19192), .B(n19191), .ZN(
        P2_U2835) );
  NOR2_X1 U22238 ( .A1(n19244), .A2(n19194), .ZN(n19195) );
  XNOR2_X1 U22239 ( .A(n19196), .B(n19195), .ZN(n19206) );
  INV_X1 U22240 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n19198) );
  OAI222_X1 U22241 ( .A1(n19304), .A2(n19199), .B1(n19198), .B2(n19303), .C1(
        n19197), .C2(n19334), .ZN(n19200) );
  AOI211_X1 U22242 ( .C1(P2_REIP_REG_19__SCAN_IN), .C2(n19325), .A(n19427), 
        .B(n19200), .ZN(n19205) );
  INV_X1 U22243 ( .A(n19201), .ZN(n19203) );
  AOI22_X1 U22244 ( .A1(n19203), .A2(n19314), .B1(n19202), .B2(n19327), .ZN(
        n19204) );
  OAI211_X1 U22245 ( .C1(n19977), .C2(n19206), .A(n19205), .B(n19204), .ZN(
        P2_U2836) );
  OAI21_X1 U22246 ( .B1(n20017), .B2(n19301), .A(n19300), .ZN(n19211) );
  INV_X1 U22247 ( .A(n19207), .ZN(n19209) );
  OAI22_X1 U22248 ( .A1(n19209), .A2(n19304), .B1(n19208), .B2(n19303), .ZN(
        n19210) );
  AOI211_X1 U22249 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n19308), .A(
        n19211), .B(n19210), .ZN(n19218) );
  NAND2_X1 U22250 ( .A1(n19310), .A2(n19212), .ZN(n19213) );
  XNOR2_X1 U22251 ( .A(n19214), .B(n19213), .ZN(n19216) );
  AOI22_X1 U22252 ( .A1(n19216), .A2(n19315), .B1(n19215), .B2(n19314), .ZN(
        n19217) );
  OAI211_X1 U22253 ( .C1(n19219), .C2(n19320), .A(n19218), .B(n19217), .ZN(
        P2_U2837) );
  NOR2_X1 U22254 ( .A1(n19244), .A2(n19220), .ZN(n19221) );
  XNOR2_X1 U22255 ( .A(n19222), .B(n19221), .ZN(n19231) );
  INV_X1 U22256 ( .A(n19223), .ZN(n19224) );
  OAI222_X1 U22257 ( .A1(n19304), .A2(n19224), .B1(n10588), .B2(n19303), .C1(
        n16428), .C2(n19334), .ZN(n19225) );
  AOI211_X1 U22258 ( .C1(P2_REIP_REG_17__SCAN_IN), .C2(n19325), .A(n19427), 
        .B(n19225), .ZN(n19230) );
  OAI22_X1 U22259 ( .A1(n19227), .A2(n19321), .B1(n19226), .B2(n19320), .ZN(
        n19228) );
  INV_X1 U22260 ( .A(n19228), .ZN(n19229) );
  OAI211_X1 U22261 ( .C1(n19977), .C2(n19231), .A(n19230), .B(n19229), .ZN(
        P2_U2838) );
  AOI22_X1 U22262 ( .A1(n19232), .A2(n19324), .B1(P2_EBX_REG_16__SCAN_IN), 
        .B2(n19326), .ZN(n19233) );
  OAI211_X1 U22263 ( .C1(n15584), .C2(n19301), .A(n19233), .B(n19300), .ZN(
        n19234) );
  AOI21_X1 U22264 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n19308), .A(
        n19234), .ZN(n19241) );
  NAND2_X1 U22265 ( .A1(n19310), .A2(n19235), .ZN(n19236) );
  XNOR2_X1 U22266 ( .A(n19237), .B(n19236), .ZN(n19239) );
  AOI22_X1 U22267 ( .A1(n19239), .A2(n19315), .B1(n19238), .B2(n19314), .ZN(
        n19240) );
  OAI211_X1 U22268 ( .C1(n19242), .C2(n19320), .A(n19241), .B(n19240), .ZN(
        P2_U2839) );
  NOR2_X1 U22269 ( .A1(n19244), .A2(n19243), .ZN(n19245) );
  XNOR2_X1 U22270 ( .A(n19246), .B(n19245), .ZN(n19255) );
  AOI22_X1 U22271 ( .A1(n19247), .A2(n19324), .B1(P2_EBX_REG_15__SCAN_IN), 
        .B2(n19326), .ZN(n19248) );
  OAI21_X1 U22272 ( .B1(n19249), .B2(n19334), .A(n19248), .ZN(n19250) );
  AOI211_X1 U22273 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n19325), .A(n19427), 
        .B(n19250), .ZN(n19254) );
  AOI22_X1 U22274 ( .A1(n19252), .A2(n19314), .B1(n19327), .B2(n19251), .ZN(
        n19253) );
  OAI211_X1 U22275 ( .C1(n19977), .C2(n19255), .A(n19254), .B(n19253), .ZN(
        P2_U2840) );
  AOI22_X1 U22276 ( .A1(n19256), .A2(n19324), .B1(P2_EBX_REG_14__SCAN_IN), 
        .B2(n19326), .ZN(n19257) );
  OAI211_X1 U22277 ( .C1(n10947), .C2(n19301), .A(n19257), .B(n19300), .ZN(
        n19258) );
  AOI21_X1 U22278 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19308), .A(
        n19258), .ZN(n19265) );
  NAND2_X1 U22279 ( .A1(n19310), .A2(n19259), .ZN(n19260) );
  XNOR2_X1 U22280 ( .A(n19261), .B(n19260), .ZN(n19263) );
  AOI22_X1 U22281 ( .A1(n19263), .A2(n19315), .B1(n19262), .B2(n19314), .ZN(
        n19264) );
  OAI211_X1 U22282 ( .C1(n19343), .C2(n19320), .A(n19265), .B(n19264), .ZN(
        P2_U2841) );
  NAND2_X1 U22283 ( .A1(n19310), .A2(n19266), .ZN(n19284) );
  XNOR2_X1 U22284 ( .A(n19267), .B(n19284), .ZN(n19277) );
  INV_X1 U22285 ( .A(n19268), .ZN(n19269) );
  AOI22_X1 U22286 ( .A1(n19269), .A2(n19324), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19308), .ZN(n19270) );
  OAI21_X1 U22287 ( .B1(n19303), .B2(n10722), .A(n19270), .ZN(n19271) );
  AOI211_X1 U22288 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19325), .A(n19427), 
        .B(n19271), .ZN(n19276) );
  INV_X1 U22289 ( .A(n19272), .ZN(n19273) );
  AOI22_X1 U22290 ( .A1(n19274), .A2(n19314), .B1(n19327), .B2(n19273), .ZN(
        n19275) );
  OAI211_X1 U22291 ( .C1(n19977), .C2(n19277), .A(n19276), .B(n19275), .ZN(
        P2_U2843) );
  AOI22_X1 U22292 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n19308), .B1(
        P2_REIP_REG_11__SCAN_IN), .B2(n19325), .ZN(n19278) );
  OAI211_X1 U22293 ( .C1(n19320), .C2(n19350), .A(n19278), .B(n19300), .ZN(
        n19279) );
  AOI21_X1 U22294 ( .B1(n19326), .B2(P2_EBX_REG_11__SCAN_IN), .A(n19279), .ZN(
        n19280) );
  OAI21_X1 U22295 ( .B1(n19281), .B2(n19321), .A(n19280), .ZN(n19282) );
  AOI21_X1 U22296 ( .B1(n19283), .B2(n19324), .A(n19282), .ZN(n19288) );
  INV_X1 U22297 ( .A(n19284), .ZN(n19285) );
  OAI211_X1 U22298 ( .C1(n19286), .C2(n19289), .A(n19315), .B(n19285), .ZN(
        n19287) );
  OAI211_X1 U22299 ( .C1(n19333), .C2(n19289), .A(n19288), .B(n19287), .ZN(
        P2_U2844) );
  OAI222_X1 U22300 ( .A1(n10170), .A2(n19334), .B1(n19291), .B2(n19303), .C1(
        n19290), .C2(n19304), .ZN(n19292) );
  AOI211_X1 U22301 ( .C1(P2_REIP_REG_8__SCAN_IN), .C2(n19325), .A(n19427), .B(
        n19292), .ZN(n19299) );
  NAND2_X1 U22302 ( .A1(n19310), .A2(n19293), .ZN(n19294) );
  XNOR2_X1 U22303 ( .A(n19295), .B(n19294), .ZN(n19297) );
  AOI22_X1 U22304 ( .A1(n19297), .A2(n19315), .B1(n19314), .B2(n19296), .ZN(
        n19298) );
  OAI211_X1 U22305 ( .C1(n19354), .C2(n19320), .A(n19299), .B(n19298), .ZN(
        P2_U2847) );
  OAI21_X1 U22306 ( .B1(n10860), .B2(n19301), .A(n19300), .ZN(n19307) );
  INV_X1 U22307 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n19302) );
  OAI22_X1 U22308 ( .A1(n19305), .A2(n19304), .B1(n19303), .B2(n19302), .ZN(
        n19306) );
  AOI211_X1 U22309 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19308), .A(
        n19307), .B(n19306), .ZN(n19318) );
  NAND2_X1 U22310 ( .A1(n19310), .A2(n19309), .ZN(n19311) );
  XNOR2_X1 U22311 ( .A(n19312), .B(n19311), .ZN(n19316) );
  AOI22_X1 U22312 ( .A1(n19316), .A2(n19315), .B1(n19314), .B2(n19313), .ZN(
        n19317) );
  OAI211_X1 U22313 ( .C1(n19320), .C2(n19319), .A(n19318), .B(n19317), .ZN(
        P2_U2849) );
  OR2_X1 U22314 ( .A1(n19322), .A2(n19321), .ZN(n19331) );
  AOI22_X1 U22315 ( .A1(n19325), .A2(P2_REIP_REG_0__SCAN_IN), .B1(n19324), 
        .B2(n19323), .ZN(n19330) );
  NAND2_X1 U22316 ( .A1(n19326), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n19329) );
  NAND2_X1 U22317 ( .A1(n19327), .A2(n19386), .ZN(n19328) );
  NAND4_X1 U22318 ( .A1(n19331), .A2(n19330), .A3(n19329), .A4(n19328), .ZN(
        n19336) );
  INV_X1 U22319 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19332) );
  AOI21_X1 U22320 ( .B1(n19334), .B2(n19333), .A(n19332), .ZN(n19335) );
  AOI211_X1 U22321 ( .C1(n20093), .C2(n19337), .A(n19336), .B(n19335), .ZN(
        n19338) );
  OAI21_X1 U22322 ( .B1(n19340), .B2(n19339), .A(n19338), .ZN(P2_U2855) );
  INV_X1 U22323 ( .A(n19389), .ZN(n19352) );
  AOI22_X1 U22324 ( .A1(n19352), .A2(n19341), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n19382), .ZN(n19342) );
  OAI21_X1 U22325 ( .B1(n19355), .B2(n19343), .A(n19342), .ZN(P2_U2905) );
  INV_X1 U22326 ( .A(n19344), .ZN(n19347) );
  AOI22_X1 U22327 ( .A1(n19352), .A2(n19345), .B1(P2_EAX_REG_13__SCAN_IN), 
        .B2(n19382), .ZN(n19346) );
  OAI21_X1 U22328 ( .B1(n19355), .B2(n19347), .A(n19346), .ZN(P2_U2906) );
  AOI22_X1 U22329 ( .A1(n19352), .A2(n19348), .B1(P2_EAX_REG_11__SCAN_IN), 
        .B2(n19382), .ZN(n19349) );
  OAI21_X1 U22330 ( .B1(n19355), .B2(n19350), .A(n19349), .ZN(P2_U2908) );
  AOI22_X1 U22331 ( .A1(n19352), .A2(n19351), .B1(P2_EAX_REG_8__SCAN_IN), .B2(
        n19382), .ZN(n19353) );
  OAI21_X1 U22332 ( .B1(n19355), .B2(n19354), .A(n19353), .ZN(P2_U2911) );
  INV_X1 U22333 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19356) );
  OAI22_X1 U22334 ( .A1(n19359), .A2(n19358), .B1(n19357), .B2(n19356), .ZN(
        n19360) );
  INV_X1 U22335 ( .A(n19360), .ZN(n19365) );
  XNOR2_X1 U22336 ( .A(n19362), .B(n19361), .ZN(n19363) );
  NAND2_X1 U22337 ( .A1(n19363), .A2(n19385), .ZN(n19364) );
  OAI211_X1 U22338 ( .C1(n19469), .C2(n19389), .A(n19365), .B(n19364), .ZN(
        P2_U2915) );
  AOI22_X1 U22339 ( .A1(n19383), .A2(n20069), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19382), .ZN(n19371) );
  OAI21_X1 U22340 ( .B1(n19368), .B2(n19367), .A(n19366), .ZN(n19369) );
  NAND2_X1 U22341 ( .A1(n19369), .A2(n19385), .ZN(n19370) );
  OAI211_X1 U22342 ( .C1(n19465), .C2(n19389), .A(n19371), .B(n19370), .ZN(
        P2_U2916) );
  AOI22_X1 U22343 ( .A1(n19383), .A2(n20077), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19382), .ZN(n19376) );
  XNOR2_X1 U22344 ( .A(n19373), .B(n19372), .ZN(n19374) );
  NAND2_X1 U22345 ( .A1(n19374), .A2(n19385), .ZN(n19375) );
  OAI211_X1 U22346 ( .C1(n19460), .C2(n19389), .A(n19376), .B(n19375), .ZN(
        P2_U2917) );
  AOI22_X1 U22347 ( .A1(n19383), .A2(n20086), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19382), .ZN(n19380) );
  XNOR2_X1 U22348 ( .A(n19377), .B(n19384), .ZN(n19378) );
  NAND2_X1 U22349 ( .A1(n19378), .A2(n19385), .ZN(n19379) );
  OAI211_X1 U22350 ( .C1(n19381), .C2(n19389), .A(n19380), .B(n19379), .ZN(
        P2_U2918) );
  AOI22_X1 U22351 ( .A1(n19383), .A2(n19386), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n19382), .ZN(n19388) );
  OAI211_X1 U22352 ( .C1(n20093), .C2(n19386), .A(n19385), .B(n19384), .ZN(
        n19387) );
  OAI211_X1 U22353 ( .C1(n19390), .C2(n19389), .A(n19388), .B(n19387), .ZN(
        P2_U2919) );
  AND2_X1 U22354 ( .A1(n19410), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  AOI22_X1 U22355 ( .A1(n20113), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19392) );
  OAI21_X1 U22356 ( .B1(n19393), .B2(n19423), .A(n19392), .ZN(P2_U2936) );
  AOI22_X1 U22357 ( .A1(n20113), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19394) );
  OAI21_X1 U22358 ( .B1(n19395), .B2(n19423), .A(n19394), .ZN(P2_U2937) );
  AOI22_X1 U22359 ( .A1(n20113), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19396) );
  OAI21_X1 U22360 ( .B1(n19397), .B2(n19423), .A(n19396), .ZN(P2_U2938) );
  AOI22_X1 U22361 ( .A1(n20113), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19398) );
  OAI21_X1 U22362 ( .B1(n19399), .B2(n19423), .A(n19398), .ZN(P2_U2939) );
  AOI22_X1 U22363 ( .A1(n20113), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19400) );
  OAI21_X1 U22364 ( .B1(n19401), .B2(n19423), .A(n19400), .ZN(P2_U2940) );
  AOI22_X1 U22365 ( .A1(n20113), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19402) );
  OAI21_X1 U22366 ( .B1(n19403), .B2(n19423), .A(n19402), .ZN(P2_U2941) );
  AOI22_X1 U22367 ( .A1(n20113), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19404) );
  OAI21_X1 U22368 ( .B1(n19405), .B2(n19423), .A(n19404), .ZN(P2_U2942) );
  AOI22_X1 U22369 ( .A1(n20113), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19406) );
  OAI21_X1 U22370 ( .B1(n19407), .B2(n19423), .A(n19406), .ZN(P2_U2943) );
  AOI22_X1 U22371 ( .A1(n20113), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19408) );
  OAI21_X1 U22372 ( .B1(n19409), .B2(n19423), .A(n19408), .ZN(P2_U2944) );
  AOI22_X1 U22373 ( .A1(n20113), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19411) );
  OAI21_X1 U22374 ( .B1(n19412), .B2(n19423), .A(n19411), .ZN(P2_U2945) );
  AOI22_X1 U22375 ( .A1(n20113), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19413) );
  OAI21_X1 U22376 ( .B1(n19414), .B2(n19423), .A(n19413), .ZN(P2_U2946) );
  AOI22_X1 U22377 ( .A1(n20113), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19415) );
  OAI21_X1 U22378 ( .B1(n19356), .B2(n19423), .A(n19415), .ZN(P2_U2947) );
  INV_X1 U22379 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19417) );
  AOI22_X1 U22380 ( .A1(n20113), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19416) );
  OAI21_X1 U22381 ( .B1(n19417), .B2(n19423), .A(n19416), .ZN(P2_U2948) );
  INV_X1 U22382 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19419) );
  AOI22_X1 U22383 ( .A1(n20113), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19418) );
  OAI21_X1 U22384 ( .B1(n19419), .B2(n19423), .A(n19418), .ZN(P2_U2949) );
  INV_X1 U22385 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19421) );
  AOI22_X1 U22386 ( .A1(n20113), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19420) );
  OAI21_X1 U22387 ( .B1(n19421), .B2(n19423), .A(n19420), .ZN(P2_U2950) );
  INV_X1 U22388 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19424) );
  AOI22_X1 U22389 ( .A1(n20113), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19410), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19422) );
  OAI21_X1 U22390 ( .B1(n19424), .B2(n19423), .A(n19422), .ZN(P2_U2951) );
  AOI22_X1 U22391 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19427), .B1(n19426), 
        .B2(n19425), .ZN(n19437) );
  INV_X1 U22392 ( .A(n19428), .ZN(n19432) );
  OAI22_X1 U22393 ( .A1(n19432), .A2(n19431), .B1(n19430), .B2(n19429), .ZN(
        n19433) );
  AOI21_X1 U22394 ( .B1(n19435), .B2(n19434), .A(n19433), .ZN(n19436) );
  OAI211_X1 U22395 ( .C1(n19439), .C2(n19438), .A(n19437), .B(n19436), .ZN(
        P2_U3010) );
  INV_X1 U22396 ( .A(n19836), .ZN(n19441) );
  INV_X1 U22397 ( .A(n19864), .ZN(n19914) );
  NAND2_X1 U22398 ( .A1(n19554), .A2(n20088), .ZN(n19500) );
  NOR2_X1 U22399 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19500), .ZN(
        n19487) );
  AOI22_X1 U22400 ( .A1(n19488), .A2(n19921), .B1(n19912), .B2(n19487), .ZN(
        n19454) );
  INV_X1 U22401 ( .A(n19522), .ZN(n19442) );
  NOR2_X1 U22402 ( .A1(n19488), .A2(n19442), .ZN(n19443) );
  OAI21_X1 U22403 ( .B1(n19443), .B2(n19726), .A(n20068), .ZN(n19452) );
  NOR2_X1 U22404 ( .A1(n19444), .A2(n10331), .ZN(n19961) );
  NOR2_X1 U22405 ( .A1(n19961), .A2(n19487), .ZN(n19451) );
  INV_X1 U22406 ( .A(n19451), .ZN(n19447) );
  INV_X1 U22407 ( .A(n19487), .ZN(n19445) );
  OAI211_X1 U22408 ( .C1(n19448), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19868), 
        .B(n19445), .ZN(n19446) );
  OAI211_X1 U22409 ( .C1(n19452), .C2(n19447), .A(n19919), .B(n19446), .ZN(
        n19491) );
  INV_X1 U22410 ( .A(n19448), .ZN(n19449) );
  OAI21_X1 U22411 ( .B1(n19449), .B2(n19487), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19450) );
  AOI22_X1 U22412 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19491), .B1(
        n19913), .B2(n19490), .ZN(n19453) );
  OAI211_X1 U22413 ( .C1(n19924), .C2(n19522), .A(n19454), .B(n19453), .ZN(
        P2_U3048) );
  AOI22_X1 U22414 ( .A1(n19488), .A2(n19927), .B1(n19925), .B2(n19487), .ZN(
        n19456) );
  AOI22_X1 U22415 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19491), .B1(
        n19926), .B2(n19490), .ZN(n19455) );
  OAI211_X1 U22416 ( .C1(n19930), .C2(n19522), .A(n19456), .B(n19455), .ZN(
        P2_U3049) );
  AOI22_X1 U22417 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19480), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19479), .ZN(n19936) );
  OAI22_X2 U22418 ( .A1(n19458), .A2(n19481), .B1(n19457), .B2(n19483), .ZN(
        n19933) );
  AOI22_X1 U22419 ( .A1(n19488), .A2(n19933), .B1(n19931), .B2(n19487), .ZN(
        n19462) );
  NOR2_X2 U22420 ( .A1(n19460), .A2(n19639), .ZN(n19932) );
  AOI22_X1 U22421 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19491), .B1(
        n19932), .B2(n19490), .ZN(n19461) );
  OAI211_X1 U22422 ( .C1(n19936), .C2(n19522), .A(n19462), .B(n19461), .ZN(
        P2_U3050) );
  AOI22_X1 U22423 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19480), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19479), .ZN(n19942) );
  NOR2_X2 U22424 ( .A1(n10640), .A2(n19468), .ZN(n19937) );
  AOI22_X1 U22425 ( .A1(n19488), .A2(n19939), .B1(n19937), .B2(n19487), .ZN(
        n19467) );
  NOR2_X2 U22426 ( .A1(n19465), .A2(n19639), .ZN(n19938) );
  AOI22_X1 U22427 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19491), .B1(
        n19938), .B2(n19490), .ZN(n19466) );
  OAI211_X1 U22428 ( .C1(n19942), .C2(n19522), .A(n19467), .B(n19466), .ZN(
        P2_U3051) );
  AOI22_X1 U22429 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19480), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19479), .ZN(n19948) );
  AOI22_X1 U22430 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19480), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19479), .ZN(n19851) );
  INV_X1 U22431 ( .A(n19851), .ZN(n19945) );
  NOR2_X2 U22432 ( .A1(n10647), .A2(n19468), .ZN(n19943) );
  AOI22_X1 U22433 ( .A1(n19488), .A2(n19945), .B1(n19943), .B2(n19487), .ZN(
        n19471) );
  NOR2_X2 U22434 ( .A1(n19469), .A2(n19639), .ZN(n19944) );
  AOI22_X1 U22435 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19491), .B1(
        n19944), .B2(n19490), .ZN(n19470) );
  OAI211_X1 U22436 ( .C1(n19948), .C2(n19522), .A(n19471), .B(n19470), .ZN(
        P2_U3052) );
  AOI22_X1 U22437 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19480), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19479), .ZN(n19954) );
  AOI22_X1 U22438 ( .A1(n19488), .A2(n19951), .B1(n19949), .B2(n19487), .ZN(
        n19476) );
  NOR2_X2 U22439 ( .A1(n19474), .A2(n19639), .ZN(n19950) );
  AOI22_X1 U22440 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19491), .B1(
        n19950), .B2(n19490), .ZN(n19475) );
  OAI211_X1 U22441 ( .C1(n19954), .C2(n19522), .A(n19476), .B(n19475), .ZN(
        P2_U3053) );
  AOI22_X1 U22442 ( .A1(n19488), .A2(n19957), .B1(n19955), .B2(n19487), .ZN(
        n19478) );
  AOI22_X1 U22443 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19491), .B1(
        n19956), .B2(n19490), .ZN(n19477) );
  OAI211_X1 U22444 ( .C1(n19960), .C2(n19522), .A(n19478), .B(n19477), .ZN(
        P2_U3054) );
  AOI22_X1 U22445 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19480), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19479), .ZN(n19971) );
  AOI22_X1 U22446 ( .A1(n19488), .A2(n19965), .B1(n19962), .B2(n19487), .ZN(
        n19493) );
  NOR2_X2 U22447 ( .A1(n19489), .A2(n19639), .ZN(n19963) );
  AOI22_X1 U22448 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19491), .B1(
        n19963), .B2(n19490), .ZN(n19492) );
  OAI211_X1 U22449 ( .C1(n19971), .C2(n19522), .A(n19493), .B(n19492), .ZN(
        P2_U3055) );
  INV_X1 U22450 ( .A(n19921), .ZN(n19839) );
  INV_X1 U22451 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19591) );
  INV_X1 U22452 ( .A(n19972), .ZN(n19497) );
  INV_X1 U22453 ( .A(n19494), .ZN(n19496) );
  NOR2_X1 U22454 ( .A1(n19495), .A2(n19525), .ZN(n19517) );
  NOR3_X1 U22455 ( .A1(n19496), .A2(n19517), .A3(n19591), .ZN(n19499) );
  AOI211_X2 U22456 ( .C1(n19500), .C2(n19591), .A(n19497), .B(n19499), .ZN(
        n19518) );
  AOI22_X1 U22457 ( .A1(n19518), .A2(n19913), .B1(n19912), .B2(n19517), .ZN(
        n19504) );
  INV_X1 U22458 ( .A(n19671), .ZN(n19498) );
  INV_X1 U22459 ( .A(n19728), .ZN(n19694) );
  NAND2_X1 U22460 ( .A1(n19498), .A2(n19694), .ZN(n19501) );
  AOI21_X1 U22461 ( .B1(n19501), .B2(n19500), .A(n19499), .ZN(n19502) );
  OAI211_X1 U22462 ( .C1(n19517), .C2(n20089), .A(n19502), .B(n19919), .ZN(
        n19519) );
  NOR2_X2 U22463 ( .A1(n19728), .A2(n19667), .ZN(n19549) );
  AOI22_X1 U22464 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19519), .B1(
        n19549), .B2(n19873), .ZN(n19503) );
  OAI211_X1 U22465 ( .C1(n19839), .C2(n19522), .A(n19504), .B(n19503), .ZN(
        P2_U3056) );
  AOI22_X1 U22466 ( .A1(n19518), .A2(n19926), .B1(n19925), .B2(n19517), .ZN(
        n19506) );
  AOI22_X1 U22467 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19519), .B1(
        n19549), .B2(n19883), .ZN(n19505) );
  OAI211_X1 U22468 ( .C1(n19842), .C2(n19522), .A(n19506), .B(n19505), .ZN(
        P2_U3057) );
  INV_X1 U22469 ( .A(n19933), .ZN(n19845) );
  AOI22_X1 U22470 ( .A1(n19518), .A2(n19932), .B1(n19931), .B2(n19517), .ZN(
        n19508) );
  INV_X1 U22471 ( .A(n19936), .ZN(n19886) );
  AOI22_X1 U22472 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19519), .B1(
        n19549), .B2(n19886), .ZN(n19507) );
  OAI211_X1 U22473 ( .C1(n19845), .C2(n19522), .A(n19508), .B(n19507), .ZN(
        P2_U3058) );
  INV_X1 U22474 ( .A(n19939), .ZN(n19848) );
  AOI22_X1 U22475 ( .A1(n19518), .A2(n19938), .B1(n19937), .B2(n19517), .ZN(
        n19510) );
  AOI22_X1 U22476 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19519), .B1(
        n19549), .B2(n19889), .ZN(n19509) );
  OAI211_X1 U22477 ( .C1(n19848), .C2(n19522), .A(n19510), .B(n19509), .ZN(
        P2_U3059) );
  AOI22_X1 U22478 ( .A1(n19518), .A2(n19944), .B1(n19943), .B2(n19517), .ZN(
        n19512) );
  AOI22_X1 U22479 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19519), .B1(
        n19549), .B2(n19892), .ZN(n19511) );
  OAI211_X1 U22480 ( .C1(n19851), .C2(n19522), .A(n19512), .B(n19511), .ZN(
        P2_U3060) );
  INV_X1 U22481 ( .A(n19951), .ZN(n19854) );
  AOI22_X1 U22482 ( .A1(n19518), .A2(n19950), .B1(n19949), .B2(n19517), .ZN(
        n19514) );
  AOI22_X1 U22483 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19519), .B1(
        n19549), .B2(n19895), .ZN(n19513) );
  OAI211_X1 U22484 ( .C1(n19854), .C2(n19522), .A(n19514), .B(n19513), .ZN(
        P2_U3061) );
  AOI22_X1 U22485 ( .A1(n19518), .A2(n19956), .B1(n19955), .B2(n19517), .ZN(
        n19516) );
  AOI22_X1 U22486 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19519), .B1(
        n19549), .B2(n19898), .ZN(n19515) );
  OAI211_X1 U22487 ( .C1(n19857), .C2(n19522), .A(n19516), .B(n19515), .ZN(
        P2_U3062) );
  INV_X1 U22488 ( .A(n19965), .ZN(n19863) );
  AOI22_X1 U22489 ( .A1(n19518), .A2(n19963), .B1(n19962), .B2(n19517), .ZN(
        n19521) );
  AOI22_X1 U22490 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19519), .B1(
        n19549), .B2(n19903), .ZN(n19520) );
  OAI211_X1 U22491 ( .C1(n19863), .C2(n19522), .A(n19521), .B(n19520), .ZN(
        P2_U3063) );
  INV_X1 U22492 ( .A(n19528), .ZN(n19524) );
  NOR2_X1 U22493 ( .A1(n19523), .A2(n19525), .ZN(n19547) );
  OAI21_X1 U22494 ( .B1(n19524), .B2(n19547), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19527) );
  OR2_X1 U22495 ( .A1(n19526), .A2(n19525), .ZN(n19529) );
  NAND2_X1 U22496 ( .A1(n19527), .A2(n19529), .ZN(n19548) );
  AOI22_X1 U22497 ( .A1(n19548), .A2(n19913), .B1(n19912), .B2(n19547), .ZN(
        n19534) );
  AOI21_X1 U22498 ( .B1(n19528), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19532) );
  OAI21_X1 U22499 ( .B1(n19578), .B2(n19549), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19530) );
  NAND3_X1 U22500 ( .A1(n19530), .A2(n20068), .A3(n19529), .ZN(n19531) );
  OAI211_X1 U22501 ( .C1(n19547), .C2(n19532), .A(n19531), .B(n19919), .ZN(
        n19550) );
  AOI22_X1 U22502 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19550), .B1(
        n19549), .B2(n19921), .ZN(n19533) );
  OAI211_X1 U22503 ( .C1(n19924), .C2(n19576), .A(n19534), .B(n19533), .ZN(
        P2_U3064) );
  AOI22_X1 U22504 ( .A1(n19548), .A2(n19926), .B1(n19925), .B2(n19547), .ZN(
        n19536) );
  AOI22_X1 U22505 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19550), .B1(
        n19549), .B2(n19927), .ZN(n19535) );
  OAI211_X1 U22506 ( .C1(n19930), .C2(n19576), .A(n19536), .B(n19535), .ZN(
        P2_U3065) );
  AOI22_X1 U22507 ( .A1(n19548), .A2(n19932), .B1(n19931), .B2(n19547), .ZN(
        n19538) );
  AOI22_X1 U22508 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19550), .B1(
        n19549), .B2(n19933), .ZN(n19537) );
  OAI211_X1 U22509 ( .C1(n19936), .C2(n19576), .A(n19538), .B(n19537), .ZN(
        P2_U3066) );
  AOI22_X1 U22510 ( .A1(n19548), .A2(n19938), .B1(n19937), .B2(n19547), .ZN(
        n19540) );
  AOI22_X1 U22511 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19550), .B1(
        n19549), .B2(n19939), .ZN(n19539) );
  OAI211_X1 U22512 ( .C1(n19942), .C2(n19576), .A(n19540), .B(n19539), .ZN(
        P2_U3067) );
  AOI22_X1 U22513 ( .A1(n19548), .A2(n19944), .B1(n19943), .B2(n19547), .ZN(
        n19542) );
  AOI22_X1 U22514 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19550), .B1(
        n19549), .B2(n19945), .ZN(n19541) );
  OAI211_X1 U22515 ( .C1(n19948), .C2(n19576), .A(n19542), .B(n19541), .ZN(
        P2_U3068) );
  AOI22_X1 U22516 ( .A1(n19548), .A2(n19950), .B1(n19949), .B2(n19547), .ZN(
        n19544) );
  AOI22_X1 U22517 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19550), .B1(
        n19549), .B2(n19951), .ZN(n19543) );
  OAI211_X1 U22518 ( .C1(n19954), .C2(n19576), .A(n19544), .B(n19543), .ZN(
        P2_U3069) );
  AOI22_X1 U22519 ( .A1(n19548), .A2(n19956), .B1(n19955), .B2(n19547), .ZN(
        n19546) );
  AOI22_X1 U22520 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19550), .B1(
        n19549), .B2(n19957), .ZN(n19545) );
  OAI211_X1 U22521 ( .C1(n19960), .C2(n19576), .A(n19546), .B(n19545), .ZN(
        P2_U3070) );
  AOI22_X1 U22522 ( .A1(n19548), .A2(n19963), .B1(n19962), .B2(n19547), .ZN(
        n19552) );
  AOI22_X1 U22523 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19550), .B1(
        n19549), .B2(n19965), .ZN(n19551) );
  OAI211_X1 U22524 ( .C1(n19971), .C2(n19576), .A(n19552), .B(n19551), .ZN(
        P2_U3071) );
  AND2_X1 U22525 ( .A1(n19779), .A2(n19554), .ZN(n19577) );
  AOI22_X1 U22526 ( .A1(n19921), .A2(n19578), .B1(n19912), .B2(n19577), .ZN(
        n19563) );
  OAI21_X1 U22527 ( .B1(n19553), .B2(n19671), .A(n20068), .ZN(n19561) );
  NAND2_X1 U22528 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19554), .ZN(
        n19560) );
  INV_X1 U22529 ( .A(n19560), .ZN(n19557) );
  INV_X1 U22530 ( .A(n19577), .ZN(n19555) );
  OAI211_X1 U22531 ( .C1(n12532), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19555), 
        .B(n19868), .ZN(n19556) );
  OAI211_X1 U22532 ( .C1(n19561), .C2(n19557), .A(n19919), .B(n19556), .ZN(
        n19580) );
  INV_X1 U22533 ( .A(n12532), .ZN(n19558) );
  OAI21_X1 U22534 ( .B1(n19558), .B2(n19577), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19559) );
  OAI21_X1 U22535 ( .B1(n19561), .B2(n19560), .A(n19559), .ZN(n19579) );
  AOI22_X1 U22536 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19580), .B1(
        n19913), .B2(n19579), .ZN(n19562) );
  OAI211_X1 U22537 ( .C1(n19924), .C2(n19617), .A(n19563), .B(n19562), .ZN(
        P2_U3072) );
  AOI22_X1 U22538 ( .A1(n19595), .A2(n19883), .B1(n19925), .B2(n19577), .ZN(
        n19565) );
  AOI22_X1 U22539 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19580), .B1(
        n19926), .B2(n19579), .ZN(n19564) );
  OAI211_X1 U22540 ( .C1(n19842), .C2(n19576), .A(n19565), .B(n19564), .ZN(
        P2_U3073) );
  AOI22_X1 U22541 ( .A1(n19933), .A2(n19578), .B1(n19577), .B2(n19931), .ZN(
        n19567) );
  AOI22_X1 U22542 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19580), .B1(
        n19932), .B2(n19579), .ZN(n19566) );
  OAI211_X1 U22543 ( .C1(n19936), .C2(n19617), .A(n19567), .B(n19566), .ZN(
        P2_U3074) );
  AOI22_X1 U22544 ( .A1(n19595), .A2(n19889), .B1(n19577), .B2(n19937), .ZN(
        n19569) );
  AOI22_X1 U22545 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19580), .B1(
        n19938), .B2(n19579), .ZN(n19568) );
  OAI211_X1 U22546 ( .C1(n19848), .C2(n19576), .A(n19569), .B(n19568), .ZN(
        P2_U3075) );
  AOI22_X1 U22547 ( .A1(n19578), .A2(n19945), .B1(n19577), .B2(n19943), .ZN(
        n19571) );
  AOI22_X1 U22548 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19580), .B1(
        n19944), .B2(n19579), .ZN(n19570) );
  OAI211_X1 U22549 ( .C1(n19948), .C2(n19617), .A(n19571), .B(n19570), .ZN(
        P2_U3076) );
  AOI22_X1 U22550 ( .A1(n19595), .A2(n19895), .B1(n19577), .B2(n19949), .ZN(
        n19573) );
  AOI22_X1 U22551 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19580), .B1(
        n19950), .B2(n19579), .ZN(n19572) );
  OAI211_X1 U22552 ( .C1(n19854), .C2(n19576), .A(n19573), .B(n19572), .ZN(
        P2_U3077) );
  AOI22_X1 U22553 ( .A1(n19595), .A2(n19898), .B1(n19955), .B2(n19577), .ZN(
        n19575) );
  AOI22_X1 U22554 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19580), .B1(
        n19956), .B2(n19579), .ZN(n19574) );
  OAI211_X1 U22555 ( .C1(n19857), .C2(n19576), .A(n19575), .B(n19574), .ZN(
        P2_U3078) );
  AOI22_X1 U22556 ( .A1(n19965), .A2(n19578), .B1(n19577), .B2(n19962), .ZN(
        n19582) );
  AOI22_X1 U22557 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19580), .B1(
        n19963), .B2(n19579), .ZN(n19581) );
  OAI211_X1 U22558 ( .C1(n19971), .C2(n19617), .A(n19582), .B(n19581), .ZN(
        P2_U3079) );
  NOR2_X1 U22559 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19583), .ZN(
        n19612) );
  INV_X1 U22560 ( .A(n19612), .ZN(n19588) );
  AND2_X1 U22561 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19588), .ZN(n19584) );
  NAND2_X1 U22562 ( .A1(n19585), .A2(n19584), .ZN(n19594) );
  OAI21_X1 U22563 ( .B1(n19595), .B2(n19630), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19587) );
  NAND2_X1 U22564 ( .A1(n19586), .A2(n10331), .ZN(n19592) );
  AOI22_X1 U22565 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19588), .B1(n19587), 
        .B2(n19592), .ZN(n19589) );
  AND2_X1 U22566 ( .A1(n19919), .A2(n19589), .ZN(n19590) );
  OAI21_X1 U22567 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19592), .A(n19591), 
        .ZN(n19593) );
  AND2_X1 U22568 ( .A1(n19594), .A2(n19593), .ZN(n19613) );
  AOI22_X1 U22569 ( .A1(n19613), .A2(n19913), .B1(n19912), .B2(n19612), .ZN(
        n19597) );
  AOI22_X1 U22570 ( .A1(n19595), .A2(n19921), .B1(n19630), .B2(n19873), .ZN(
        n19596) );
  OAI211_X1 U22571 ( .C1(n19599), .C2(n19598), .A(n19597), .B(n19596), .ZN(
        P2_U3080) );
  AOI22_X1 U22572 ( .A1(n19613), .A2(n19926), .B1(n19925), .B2(n19612), .ZN(
        n19601) );
  AOI22_X1 U22573 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19614), .B1(
        n19630), .B2(n19883), .ZN(n19600) );
  OAI211_X1 U22574 ( .C1(n19842), .C2(n19617), .A(n19601), .B(n19600), .ZN(
        P2_U3081) );
  AOI22_X1 U22575 ( .A1(n19613), .A2(n19932), .B1(n19931), .B2(n19612), .ZN(
        n19603) );
  AOI22_X1 U22576 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19614), .B1(
        n19630), .B2(n19886), .ZN(n19602) );
  OAI211_X1 U22577 ( .C1(n19845), .C2(n19617), .A(n19603), .B(n19602), .ZN(
        P2_U3082) );
  AOI22_X1 U22578 ( .A1(n19613), .A2(n19938), .B1(n19937), .B2(n19612), .ZN(
        n19605) );
  AOI22_X1 U22579 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19614), .B1(
        n19630), .B2(n19889), .ZN(n19604) );
  OAI211_X1 U22580 ( .C1(n19848), .C2(n19617), .A(n19605), .B(n19604), .ZN(
        P2_U3083) );
  AOI22_X1 U22581 ( .A1(n19613), .A2(n19944), .B1(n19943), .B2(n19612), .ZN(
        n19607) );
  AOI22_X1 U22582 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19614), .B1(
        n19630), .B2(n19892), .ZN(n19606) );
  OAI211_X1 U22583 ( .C1(n19851), .C2(n19617), .A(n19607), .B(n19606), .ZN(
        P2_U3084) );
  AOI22_X1 U22584 ( .A1(n19613), .A2(n19950), .B1(n19949), .B2(n19612), .ZN(
        n19609) );
  AOI22_X1 U22585 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19614), .B1(
        n19630), .B2(n19895), .ZN(n19608) );
  OAI211_X1 U22586 ( .C1(n19854), .C2(n19617), .A(n19609), .B(n19608), .ZN(
        P2_U3085) );
  AOI22_X1 U22587 ( .A1(n19613), .A2(n19956), .B1(n19955), .B2(n19612), .ZN(
        n19611) );
  AOI22_X1 U22588 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19614), .B1(
        n19630), .B2(n19898), .ZN(n19610) );
  OAI211_X1 U22589 ( .C1(n19857), .C2(n19617), .A(n19611), .B(n19610), .ZN(
        P2_U3086) );
  AOI22_X1 U22590 ( .A1(n19613), .A2(n19963), .B1(n19962), .B2(n19612), .ZN(
        n19616) );
  AOI22_X1 U22591 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19614), .B1(
        n19630), .B2(n19903), .ZN(n19615) );
  OAI211_X1 U22592 ( .C1(n19863), .C2(n19617), .A(n19616), .B(n19615), .ZN(
        P2_U3087) );
  AOI22_X1 U22593 ( .A1(n19662), .A2(n19883), .B1(n19925), .B2(n19637), .ZN(
        n19619) );
  AOI22_X1 U22594 ( .A1(n19926), .A2(n19631), .B1(n19630), .B2(n19927), .ZN(
        n19618) );
  OAI211_X1 U22595 ( .C1(n19635), .C2(n12447), .A(n19619), .B(n19618), .ZN(
        P2_U3089) );
  INV_X1 U22596 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n19622) );
  AOI22_X1 U22597 ( .A1(n19933), .A2(n19630), .B1(n19637), .B2(n19931), .ZN(
        n19621) );
  AOI22_X1 U22598 ( .A1(n19932), .A2(n19631), .B1(n19662), .B2(n19886), .ZN(
        n19620) );
  OAI211_X1 U22599 ( .C1(n19635), .C2(n19622), .A(n19621), .B(n19620), .ZN(
        P2_U3090) );
  AOI22_X1 U22600 ( .A1(n19662), .A2(n19889), .B1(n19637), .B2(n19937), .ZN(
        n19624) );
  AOI22_X1 U22601 ( .A1(n19938), .A2(n19631), .B1(n19630), .B2(n19939), .ZN(
        n19623) );
  OAI211_X1 U22602 ( .C1(n19635), .C2(n12483), .A(n19624), .B(n19623), .ZN(
        P2_U3091) );
  INV_X1 U22603 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n19627) );
  AOI22_X1 U22604 ( .A1(n19630), .A2(n19945), .B1(n19637), .B2(n19943), .ZN(
        n19626) );
  AOI22_X1 U22605 ( .A1(n19944), .A2(n19631), .B1(n19662), .B2(n19892), .ZN(
        n19625) );
  OAI211_X1 U22606 ( .C1(n19635), .C2(n19627), .A(n19626), .B(n19625), .ZN(
        P2_U3092) );
  AOI22_X1 U22607 ( .A1(n19951), .A2(n19630), .B1(n19637), .B2(n19949), .ZN(
        n19629) );
  AOI22_X1 U22608 ( .A1(n19950), .A2(n19631), .B1(n19662), .B2(n19895), .ZN(
        n19628) );
  OAI211_X1 U22609 ( .C1(n19635), .C2(n12534), .A(n19629), .B(n19628), .ZN(
        P2_U3093) );
  AOI22_X1 U22610 ( .A1(n19965), .A2(n19630), .B1(n19637), .B2(n19962), .ZN(
        n19633) );
  AOI22_X1 U22611 ( .A1(n19963), .A2(n19631), .B1(n19662), .B2(n19903), .ZN(
        n19632) );
  OAI211_X1 U22612 ( .C1(n19635), .C2(n19634), .A(n19633), .B(n19632), .ZN(
        P2_U3095) );
  NOR2_X2 U22613 ( .A1(n19636), .A2(n19864), .ZN(n19690) );
  OAI21_X1 U22614 ( .B1(n19662), .B2(n19690), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19640) );
  NOR2_X1 U22615 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19670), .ZN(
        n19660) );
  NOR2_X1 U22616 ( .A1(n19637), .A2(n19660), .ZN(n19643) );
  AOI211_X1 U22617 ( .C1(n19641), .C2(n20089), .A(n20068), .B(n19660), .ZN(
        n19638) );
  OAI21_X1 U22618 ( .B1(n19641), .B2(n19660), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19642) );
  AOI22_X1 U22619 ( .A1(n19661), .A2(n19913), .B1(n19912), .B2(n19660), .ZN(
        n19645) );
  AOI22_X1 U22620 ( .A1(n19662), .A2(n19921), .B1(n19690), .B2(n19873), .ZN(
        n19644) );
  OAI211_X1 U22621 ( .C1(n19666), .C2(n19646), .A(n19645), .B(n19644), .ZN(
        P2_U3096) );
  AOI22_X1 U22622 ( .A1(n19661), .A2(n19926), .B1(n19925), .B2(n19660), .ZN(
        n19648) );
  AOI22_X1 U22623 ( .A1(n19662), .A2(n19927), .B1(n19690), .B2(n19883), .ZN(
        n19647) );
  OAI211_X1 U22624 ( .C1(n19666), .C2(n12420), .A(n19648), .B(n19647), .ZN(
        P2_U3097) );
  AOI22_X1 U22625 ( .A1(n19661), .A2(n19932), .B1(n19931), .B2(n19660), .ZN(
        n19650) );
  AOI22_X1 U22626 ( .A1(n19662), .A2(n19933), .B1(n19690), .B2(n19886), .ZN(
        n19649) );
  OAI211_X1 U22627 ( .C1(n19666), .C2(n12191), .A(n19650), .B(n19649), .ZN(
        P2_U3098) );
  AOI22_X1 U22628 ( .A1(n19661), .A2(n19938), .B1(n19937), .B2(n19660), .ZN(
        n19652) );
  AOI22_X1 U22629 ( .A1(n19662), .A2(n19939), .B1(n19690), .B2(n19889), .ZN(
        n19651) );
  OAI211_X1 U22630 ( .C1(n19666), .C2(n12477), .A(n19652), .B(n19651), .ZN(
        P2_U3099) );
  AOI22_X1 U22631 ( .A1(n19661), .A2(n19944), .B1(n19943), .B2(n19660), .ZN(
        n19654) );
  AOI22_X1 U22632 ( .A1(n19662), .A2(n19945), .B1(n19690), .B2(n19892), .ZN(
        n19653) );
  OAI211_X1 U22633 ( .C1(n19666), .C2(n19655), .A(n19654), .B(n19653), .ZN(
        P2_U3100) );
  AOI22_X1 U22634 ( .A1(n19661), .A2(n19950), .B1(n19949), .B2(n19660), .ZN(
        n19657) );
  AOI22_X1 U22635 ( .A1(n19662), .A2(n19951), .B1(n19690), .B2(n19895), .ZN(
        n19656) );
  OAI211_X1 U22636 ( .C1(n19666), .C2(n12545), .A(n19657), .B(n19656), .ZN(
        P2_U3101) );
  AOI22_X1 U22637 ( .A1(n19661), .A2(n19956), .B1(n19955), .B2(n19660), .ZN(
        n19659) );
  AOI22_X1 U22638 ( .A1(n19662), .A2(n19957), .B1(n19690), .B2(n19898), .ZN(
        n19658) );
  OAI211_X1 U22639 ( .C1(n19666), .C2(n12582), .A(n19659), .B(n19658), .ZN(
        P2_U3102) );
  INV_X1 U22640 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n19665) );
  AOI22_X1 U22641 ( .A1(n19661), .A2(n19963), .B1(n19962), .B2(n19660), .ZN(
        n19664) );
  AOI22_X1 U22642 ( .A1(n19662), .A2(n19965), .B1(n19690), .B2(n19903), .ZN(
        n19663) );
  OAI211_X1 U22643 ( .C1(n19666), .C2(n19665), .A(n19664), .B(n19663), .ZN(
        P2_U3103) );
  INV_X1 U22644 ( .A(n19702), .ZN(n19688) );
  OAI21_X1 U22645 ( .B1(n19668), .B2(n19688), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19669) );
  OAI21_X1 U22646 ( .B1(n19670), .B2(n19868), .A(n19669), .ZN(n19689) );
  AOI22_X1 U22647 ( .A1(n19689), .A2(n19913), .B1(n19688), .B2(n19912), .ZN(
        n19675) );
  NOR2_X1 U22648 ( .A1(n19671), .A2(n19864), .ZN(n20067) );
  OAI211_X1 U22649 ( .C1(n12518), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19868), 
        .B(n19702), .ZN(n19672) );
  OAI211_X1 U22650 ( .C1(n20067), .C2(n19673), .A(n19919), .B(n19672), .ZN(
        n19691) );
  AOI22_X1 U22651 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19691), .B1(
        n19690), .B2(n19921), .ZN(n19674) );
  OAI211_X1 U22652 ( .C1(n19924), .C2(n19725), .A(n19675), .B(n19674), .ZN(
        P2_U3104) );
  AOI22_X1 U22653 ( .A1(n19689), .A2(n19926), .B1(n19688), .B2(n19925), .ZN(
        n19677) );
  AOI22_X1 U22654 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19691), .B1(
        n19690), .B2(n19927), .ZN(n19676) );
  OAI211_X1 U22655 ( .C1(n19930), .C2(n19725), .A(n19677), .B(n19676), .ZN(
        P2_U3105) );
  AOI22_X1 U22656 ( .A1(n19689), .A2(n19932), .B1(n19688), .B2(n19931), .ZN(
        n19679) );
  AOI22_X1 U22657 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19691), .B1(
        n19690), .B2(n19933), .ZN(n19678) );
  OAI211_X1 U22658 ( .C1(n19936), .C2(n19725), .A(n19679), .B(n19678), .ZN(
        P2_U3106) );
  AOI22_X1 U22659 ( .A1(n19689), .A2(n19938), .B1(n19688), .B2(n19937), .ZN(
        n19681) );
  AOI22_X1 U22660 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19691), .B1(
        n19690), .B2(n19939), .ZN(n19680) );
  OAI211_X1 U22661 ( .C1(n19942), .C2(n19725), .A(n19681), .B(n19680), .ZN(
        P2_U3107) );
  AOI22_X1 U22662 ( .A1(n19689), .A2(n19944), .B1(n19688), .B2(n19943), .ZN(
        n19683) );
  AOI22_X1 U22663 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19691), .B1(
        n19690), .B2(n19945), .ZN(n19682) );
  OAI211_X1 U22664 ( .C1(n19948), .C2(n19725), .A(n19683), .B(n19682), .ZN(
        P2_U3108) );
  AOI22_X1 U22665 ( .A1(n19689), .A2(n19950), .B1(n19688), .B2(n19949), .ZN(
        n19685) );
  AOI22_X1 U22666 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19691), .B1(
        n19690), .B2(n19951), .ZN(n19684) );
  OAI211_X1 U22667 ( .C1(n19954), .C2(n19725), .A(n19685), .B(n19684), .ZN(
        P2_U3109) );
  AOI22_X1 U22668 ( .A1(n19689), .A2(n19956), .B1(n19688), .B2(n19955), .ZN(
        n19687) );
  AOI22_X1 U22669 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19691), .B1(
        n19690), .B2(n19957), .ZN(n19686) );
  OAI211_X1 U22670 ( .C1(n19960), .C2(n19725), .A(n19687), .B(n19686), .ZN(
        P2_U3110) );
  AOI22_X1 U22671 ( .A1(n19689), .A2(n19963), .B1(n19688), .B2(n19962), .ZN(
        n19693) );
  AOI22_X1 U22672 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19691), .B1(
        n19690), .B2(n19965), .ZN(n19692) );
  OAI211_X1 U22673 ( .C1(n19971), .C2(n19725), .A(n19693), .B(n19692), .ZN(
        P2_U3111) );
  INV_X1 U22674 ( .A(n19865), .ZN(n19695) );
  NOR2_X1 U22675 ( .A1(n19781), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19729) );
  INV_X1 U22676 ( .A(n19729), .ZN(n19735) );
  NOR2_X1 U22677 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19735), .ZN(
        n19720) );
  AOI22_X1 U22678 ( .A1(n19743), .A2(n19873), .B1(n19912), .B2(n19720), .ZN(
        n19707) );
  AOI21_X1 U22679 ( .B1(n19757), .B2(n19725), .A(n19726), .ZN(n19696) );
  NOR2_X1 U22680 ( .A1(n19696), .A2(n19868), .ZN(n19700) );
  INV_X1 U22681 ( .A(n19697), .ZN(n19701) );
  AOI21_X1 U22682 ( .B1(n19701), .B2(n20089), .A(n20068), .ZN(n19698) );
  AOI21_X1 U22683 ( .B1(n19700), .B2(n19702), .A(n19698), .ZN(n19699) );
  OAI21_X1 U22684 ( .B1(n19699), .B2(n19720), .A(n19919), .ZN(n19722) );
  INV_X1 U22685 ( .A(n19700), .ZN(n19705) );
  OAI21_X1 U22686 ( .B1(n19701), .B2(n19720), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19704) );
  NOR2_X1 U22687 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19720), .ZN(n19703) );
  AOI22_X1 U22688 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19722), .B1(
        n19913), .B2(n19721), .ZN(n19706) );
  OAI211_X1 U22689 ( .C1(n19839), .C2(n19725), .A(n19707), .B(n19706), .ZN(
        P2_U3112) );
  AOI22_X1 U22690 ( .A1(n19743), .A2(n19883), .B1(n19925), .B2(n19720), .ZN(
        n19709) );
  AOI22_X1 U22691 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19722), .B1(
        n19926), .B2(n19721), .ZN(n19708) );
  OAI211_X1 U22692 ( .C1(n19842), .C2(n19725), .A(n19709), .B(n19708), .ZN(
        P2_U3113) );
  AOI22_X1 U22693 ( .A1(n19743), .A2(n19886), .B1(n19931), .B2(n19720), .ZN(
        n19711) );
  AOI22_X1 U22694 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19722), .B1(
        n19932), .B2(n19721), .ZN(n19710) );
  OAI211_X1 U22695 ( .C1(n19845), .C2(n19725), .A(n19711), .B(n19710), .ZN(
        P2_U3114) );
  AOI22_X1 U22696 ( .A1(n19743), .A2(n19889), .B1(n19937), .B2(n19720), .ZN(
        n19713) );
  AOI22_X1 U22697 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19722), .B1(
        n19938), .B2(n19721), .ZN(n19712) );
  OAI211_X1 U22698 ( .C1(n19848), .C2(n19725), .A(n19713), .B(n19712), .ZN(
        P2_U3115) );
  AOI22_X1 U22699 ( .A1(n19743), .A2(n19892), .B1(n19943), .B2(n19720), .ZN(
        n19715) );
  AOI22_X1 U22700 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19722), .B1(
        n19944), .B2(n19721), .ZN(n19714) );
  OAI211_X1 U22701 ( .C1(n19851), .C2(n19725), .A(n19715), .B(n19714), .ZN(
        P2_U3116) );
  AOI22_X1 U22702 ( .A1(n19743), .A2(n19895), .B1(n19949), .B2(n19720), .ZN(
        n19717) );
  AOI22_X1 U22703 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19722), .B1(
        n19950), .B2(n19721), .ZN(n19716) );
  OAI211_X1 U22704 ( .C1(n19854), .C2(n19725), .A(n19717), .B(n19716), .ZN(
        P2_U3117) );
  AOI22_X1 U22705 ( .A1(n19743), .A2(n19898), .B1(n19955), .B2(n19720), .ZN(
        n19719) );
  AOI22_X1 U22706 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19722), .B1(
        n19956), .B2(n19721), .ZN(n19718) );
  OAI211_X1 U22707 ( .C1(n19857), .C2(n19725), .A(n19719), .B(n19718), .ZN(
        P2_U3118) );
  AOI22_X1 U22708 ( .A1(n19743), .A2(n19903), .B1(n19962), .B2(n19720), .ZN(
        n19724) );
  AOI22_X1 U22709 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19722), .B1(
        n19963), .B2(n19721), .ZN(n19723) );
  OAI211_X1 U22710 ( .C1(n19863), .C2(n19725), .A(n19724), .B(n19723), .ZN(
        P2_U3119) );
  AOI22_X1 U22711 ( .A1(n19743), .A2(n19921), .B1(n19912), .B2(n19752), .ZN(
        n19738) );
  NOR2_X1 U22712 ( .A1(n19727), .A2(n19726), .ZN(n19915) );
  INV_X1 U22713 ( .A(n19915), .ZN(n19832) );
  OAI21_X1 U22714 ( .B1(n19832), .B2(n19728), .A(n20068), .ZN(n19736) );
  NOR2_X1 U22715 ( .A1(n19736), .A2(n19729), .ZN(n19730) );
  AOI211_X1 U22716 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19732), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19730), .ZN(n19731) );
  OAI21_X1 U22717 ( .B1(n19731), .B2(n19752), .A(n19919), .ZN(n19754) );
  INV_X1 U22718 ( .A(n19732), .ZN(n19733) );
  OAI21_X1 U22719 ( .B1(n19733), .B2(n19752), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19734) );
  AOI22_X1 U22720 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19754), .B1(
        n19913), .B2(n19753), .ZN(n19737) );
  OAI211_X1 U22721 ( .C1(n19924), .C2(n19777), .A(n19738), .B(n19737), .ZN(
        P2_U3120) );
  AOI22_X1 U22722 ( .A1(n19743), .A2(n19927), .B1(n19925), .B2(n19752), .ZN(
        n19740) );
  AOI22_X1 U22723 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19754), .B1(
        n19926), .B2(n19753), .ZN(n19739) );
  OAI211_X1 U22724 ( .C1(n19930), .C2(n19777), .A(n19740), .B(n19739), .ZN(
        P2_U3121) );
  AOI22_X1 U22725 ( .A1(n19743), .A2(n19933), .B1(n19931), .B2(n19752), .ZN(
        n19742) );
  AOI22_X1 U22726 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19754), .B1(
        n19932), .B2(n19753), .ZN(n19741) );
  OAI211_X1 U22727 ( .C1(n19936), .C2(n19777), .A(n19742), .B(n19741), .ZN(
        P2_U3122) );
  AOI22_X1 U22728 ( .A1(n19743), .A2(n19939), .B1(n19937), .B2(n19752), .ZN(
        n19745) );
  AOI22_X1 U22729 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19754), .B1(
        n19938), .B2(n19753), .ZN(n19744) );
  OAI211_X1 U22730 ( .C1(n19942), .C2(n19777), .A(n19745), .B(n19744), .ZN(
        P2_U3123) );
  AOI22_X1 U22731 ( .A1(n19769), .A2(n19892), .B1(n19943), .B2(n19752), .ZN(
        n19747) );
  AOI22_X1 U22732 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19754), .B1(
        n19944), .B2(n19753), .ZN(n19746) );
  OAI211_X1 U22733 ( .C1(n19851), .C2(n19757), .A(n19747), .B(n19746), .ZN(
        P2_U3124) );
  AOI22_X1 U22734 ( .A1(n19769), .A2(n19895), .B1(n19949), .B2(n19752), .ZN(
        n19749) );
  AOI22_X1 U22735 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19754), .B1(
        n19950), .B2(n19753), .ZN(n19748) );
  OAI211_X1 U22736 ( .C1(n19854), .C2(n19757), .A(n19749), .B(n19748), .ZN(
        P2_U3125) );
  AOI22_X1 U22737 ( .A1(n19769), .A2(n19898), .B1(n19955), .B2(n19752), .ZN(
        n19751) );
  AOI22_X1 U22738 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19754), .B1(
        n19956), .B2(n19753), .ZN(n19750) );
  OAI211_X1 U22739 ( .C1(n19857), .C2(n19757), .A(n19751), .B(n19750), .ZN(
        P2_U3126) );
  AOI22_X1 U22740 ( .A1(n19769), .A2(n19903), .B1(n19962), .B2(n19752), .ZN(
        n19756) );
  AOI22_X1 U22741 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19754), .B1(
        n19963), .B2(n19753), .ZN(n19755) );
  OAI211_X1 U22742 ( .C1(n19863), .C2(n19757), .A(n19756), .B(n19755), .ZN(
        P2_U3127) );
  AOI22_X1 U22743 ( .A1(n19773), .A2(n19926), .B1(n19925), .B2(n19772), .ZN(
        n19760) );
  AOI22_X1 U22744 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19774), .B1(
        n19801), .B2(n19883), .ZN(n19759) );
  OAI211_X1 U22745 ( .C1(n19842), .C2(n19777), .A(n19760), .B(n19759), .ZN(
        P2_U3129) );
  AOI22_X1 U22746 ( .A1(n19773), .A2(n19932), .B1(n19931), .B2(n19772), .ZN(
        n19762) );
  AOI22_X1 U22747 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19774), .B1(
        n19801), .B2(n19886), .ZN(n19761) );
  OAI211_X1 U22748 ( .C1(n19845), .C2(n19777), .A(n19762), .B(n19761), .ZN(
        P2_U3130) );
  AOI22_X1 U22749 ( .A1(n19773), .A2(n19938), .B1(n19937), .B2(n19772), .ZN(
        n19764) );
  AOI22_X1 U22750 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19774), .B1(
        n19801), .B2(n19889), .ZN(n19763) );
  OAI211_X1 U22751 ( .C1(n19848), .C2(n19777), .A(n19764), .B(n19763), .ZN(
        P2_U3131) );
  AOI22_X1 U22752 ( .A1(n19773), .A2(n19944), .B1(n19943), .B2(n19772), .ZN(
        n19766) );
  AOI22_X1 U22753 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19774), .B1(
        n19801), .B2(n19892), .ZN(n19765) );
  OAI211_X1 U22754 ( .C1(n19851), .C2(n19777), .A(n19766), .B(n19765), .ZN(
        P2_U3132) );
  AOI22_X1 U22755 ( .A1(n19773), .A2(n19950), .B1(n19949), .B2(n19772), .ZN(
        n19768) );
  AOI22_X1 U22756 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19774), .B1(
        n19801), .B2(n19895), .ZN(n19767) );
  OAI211_X1 U22757 ( .C1(n19854), .C2(n19777), .A(n19768), .B(n19767), .ZN(
        P2_U3133) );
  AOI22_X1 U22758 ( .A1(n19773), .A2(n19956), .B1(n19955), .B2(n19772), .ZN(
        n19771) );
  AOI22_X1 U22759 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19774), .B1(
        n19769), .B2(n19957), .ZN(n19770) );
  OAI211_X1 U22760 ( .C1(n19960), .C2(n19809), .A(n19771), .B(n19770), .ZN(
        P2_U3134) );
  AOI22_X1 U22761 ( .A1(n19773), .A2(n19963), .B1(n19962), .B2(n19772), .ZN(
        n19776) );
  AOI22_X1 U22762 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19774), .B1(
        n19801), .B2(n19903), .ZN(n19775) );
  OAI211_X1 U22763 ( .C1(n19863), .C2(n19777), .A(n19776), .B(n19775), .ZN(
        P2_U3135) );
  INV_X1 U22764 ( .A(n19781), .ZN(n19778) );
  NAND2_X1 U22765 ( .A1(n19779), .A2(n19778), .ZN(n19784) );
  AND2_X1 U22766 ( .A1(n19784), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19780) );
  NAND2_X1 U22767 ( .A1(n12540), .A2(n19780), .ZN(n19785) );
  NOR2_X1 U22768 ( .A1(n20088), .A2(n19781), .ZN(n19788) );
  INV_X1 U22769 ( .A(n19788), .ZN(n19782) );
  OAI21_X1 U22770 ( .B1(n19782), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19591), 
        .ZN(n19783) );
  INV_X1 U22771 ( .A(n19784), .ZN(n19804) );
  AOI22_X1 U22772 ( .A1(n19805), .A2(n19913), .B1(n19912), .B2(n19804), .ZN(
        n19790) );
  OAI211_X1 U22773 ( .C1(n19804), .C2(n20089), .A(n19785), .B(n19919), .ZN(
        n19786) );
  INV_X1 U22774 ( .A(n19786), .ZN(n19787) );
  OAI221_X1 U22775 ( .B1(n19788), .B2(n20064), .C1(n19788), .C2(n19915), .A(
        n19787), .ZN(n19806) );
  AOI22_X1 U22776 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19806), .B1(
        n19801), .B2(n19921), .ZN(n19789) );
  OAI211_X1 U22777 ( .C1(n19924), .C2(n19827), .A(n19790), .B(n19789), .ZN(
        P2_U3136) );
  AOI22_X1 U22778 ( .A1(n19805), .A2(n19926), .B1(n19925), .B2(n19804), .ZN(
        n19792) );
  AOI22_X1 U22779 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19806), .B1(
        n19816), .B2(n19883), .ZN(n19791) );
  OAI211_X1 U22780 ( .C1(n19842), .C2(n19809), .A(n19792), .B(n19791), .ZN(
        P2_U3137) );
  AOI22_X1 U22781 ( .A1(n19805), .A2(n19932), .B1(n19931), .B2(n19804), .ZN(
        n19794) );
  AOI22_X1 U22782 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19806), .B1(
        n19801), .B2(n19933), .ZN(n19793) );
  OAI211_X1 U22783 ( .C1(n19936), .C2(n19827), .A(n19794), .B(n19793), .ZN(
        P2_U3138) );
  AOI22_X1 U22784 ( .A1(n19805), .A2(n19938), .B1(n19937), .B2(n19804), .ZN(
        n19796) );
  AOI22_X1 U22785 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19806), .B1(
        n19816), .B2(n19889), .ZN(n19795) );
  OAI211_X1 U22786 ( .C1(n19848), .C2(n19809), .A(n19796), .B(n19795), .ZN(
        P2_U3139) );
  AOI22_X1 U22787 ( .A1(n19805), .A2(n19944), .B1(n19943), .B2(n19804), .ZN(
        n19798) );
  AOI22_X1 U22788 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19806), .B1(
        n19816), .B2(n19892), .ZN(n19797) );
  OAI211_X1 U22789 ( .C1(n19851), .C2(n19809), .A(n19798), .B(n19797), .ZN(
        P2_U3140) );
  AOI22_X1 U22790 ( .A1(n19805), .A2(n19950), .B1(n19949), .B2(n19804), .ZN(
        n19800) );
  AOI22_X1 U22791 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19806), .B1(
        n19816), .B2(n19895), .ZN(n19799) );
  OAI211_X1 U22792 ( .C1(n19854), .C2(n19809), .A(n19800), .B(n19799), .ZN(
        P2_U3141) );
  AOI22_X1 U22793 ( .A1(n19805), .A2(n19956), .B1(n19955), .B2(n19804), .ZN(
        n19803) );
  AOI22_X1 U22794 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19806), .B1(
        n19801), .B2(n19957), .ZN(n19802) );
  OAI211_X1 U22795 ( .C1(n19960), .C2(n19827), .A(n19803), .B(n19802), .ZN(
        P2_U3142) );
  AOI22_X1 U22796 ( .A1(n19805), .A2(n19963), .B1(n19962), .B2(n19804), .ZN(
        n19808) );
  AOI22_X1 U22797 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19806), .B1(
        n19816), .B2(n19903), .ZN(n19807) );
  OAI211_X1 U22798 ( .C1(n19863), .C2(n19809), .A(n19808), .B(n19807), .ZN(
        P2_U3143) );
  AOI22_X1 U22799 ( .A1(n19822), .A2(n19932), .B1(n19821), .B2(n19931), .ZN(
        n19811) );
  AOI22_X1 U22800 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19824), .B1(
        n19823), .B2(n19886), .ZN(n19810) );
  OAI211_X1 U22801 ( .C1(n19845), .C2(n19827), .A(n19811), .B(n19810), .ZN(
        P2_U3146) );
  AOI22_X1 U22802 ( .A1(n19822), .A2(n19938), .B1(n19821), .B2(n19937), .ZN(
        n19813) );
  AOI22_X1 U22803 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19824), .B1(
        n19816), .B2(n19939), .ZN(n19812) );
  OAI211_X1 U22804 ( .C1(n19942), .C2(n19862), .A(n19813), .B(n19812), .ZN(
        P2_U3147) );
  AOI22_X1 U22805 ( .A1(n19822), .A2(n19944), .B1(n19821), .B2(n19943), .ZN(
        n19815) );
  AOI22_X1 U22806 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19824), .B1(
        n19823), .B2(n19892), .ZN(n19814) );
  OAI211_X1 U22807 ( .C1(n19851), .C2(n19827), .A(n19815), .B(n19814), .ZN(
        P2_U3148) );
  AOI22_X1 U22808 ( .A1(n19822), .A2(n19950), .B1(n19821), .B2(n19949), .ZN(
        n19818) );
  AOI22_X1 U22809 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19824), .B1(
        n19816), .B2(n19951), .ZN(n19817) );
  OAI211_X1 U22810 ( .C1(n19954), .C2(n19862), .A(n19818), .B(n19817), .ZN(
        P2_U3149) );
  AOI22_X1 U22811 ( .A1(n19822), .A2(n19956), .B1(n19821), .B2(n19955), .ZN(
        n19820) );
  AOI22_X1 U22812 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19824), .B1(
        n19823), .B2(n19898), .ZN(n19819) );
  OAI211_X1 U22813 ( .C1(n19857), .C2(n19827), .A(n19820), .B(n19819), .ZN(
        P2_U3150) );
  AOI22_X1 U22814 ( .A1(n19822), .A2(n19963), .B1(n19821), .B2(n19962), .ZN(
        n19826) );
  AOI22_X1 U22815 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19824), .B1(
        n19823), .B2(n19903), .ZN(n19825) );
  OAI211_X1 U22816 ( .C1(n19863), .C2(n19827), .A(n19826), .B(n19825), .ZN(
        P2_U3151) );
  INV_X1 U22817 ( .A(n19830), .ZN(n19828) );
  NOR2_X1 U22818 ( .A1(n20096), .A2(n19831), .ZN(n19870) );
  OAI21_X1 U22819 ( .B1(n19828), .B2(n19870), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19829) );
  OAI21_X1 U22820 ( .B1(n19831), .B2(n19868), .A(n19829), .ZN(n19858) );
  AOI22_X1 U22821 ( .A1(n19858), .A2(n19913), .B1(n19912), .B2(n19870), .ZN(
        n19838) );
  AOI21_X1 U22822 ( .B1(n19830), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19834) );
  OAI21_X1 U22823 ( .B1(n19832), .B2(n19835), .A(n19831), .ZN(n19833) );
  OAI211_X1 U22824 ( .C1(n19870), .C2(n19834), .A(n19833), .B(n19919), .ZN(
        n19859) );
  AOI22_X1 U22825 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19859), .B1(
        n19902), .B2(n19873), .ZN(n19837) );
  OAI211_X1 U22826 ( .C1(n19839), .C2(n19862), .A(n19838), .B(n19837), .ZN(
        P2_U3152) );
  AOI22_X1 U22827 ( .A1(n19858), .A2(n19926), .B1(n19925), .B2(n19870), .ZN(
        n19841) );
  AOI22_X1 U22828 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19859), .B1(
        n19902), .B2(n19883), .ZN(n19840) );
  OAI211_X1 U22829 ( .C1(n19842), .C2(n19862), .A(n19841), .B(n19840), .ZN(
        P2_U3153) );
  AOI22_X1 U22830 ( .A1(n19858), .A2(n19932), .B1(n19931), .B2(n19870), .ZN(
        n19844) );
  AOI22_X1 U22831 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19859), .B1(
        n19902), .B2(n19886), .ZN(n19843) );
  OAI211_X1 U22832 ( .C1(n19845), .C2(n19862), .A(n19844), .B(n19843), .ZN(
        P2_U3154) );
  AOI22_X1 U22833 ( .A1(n19858), .A2(n19938), .B1(n19937), .B2(n19870), .ZN(
        n19847) );
  AOI22_X1 U22834 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19859), .B1(
        n19902), .B2(n19889), .ZN(n19846) );
  OAI211_X1 U22835 ( .C1(n19848), .C2(n19862), .A(n19847), .B(n19846), .ZN(
        P2_U3155) );
  AOI22_X1 U22836 ( .A1(n19858), .A2(n19944), .B1(n19943), .B2(n19870), .ZN(
        n19850) );
  AOI22_X1 U22837 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19859), .B1(
        n19902), .B2(n19892), .ZN(n19849) );
  OAI211_X1 U22838 ( .C1(n19851), .C2(n19862), .A(n19850), .B(n19849), .ZN(
        P2_U3156) );
  AOI22_X1 U22839 ( .A1(n19858), .A2(n19950), .B1(n19949), .B2(n19870), .ZN(
        n19853) );
  AOI22_X1 U22840 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19859), .B1(
        n19902), .B2(n19895), .ZN(n19852) );
  OAI211_X1 U22841 ( .C1(n19854), .C2(n19862), .A(n19853), .B(n19852), .ZN(
        P2_U3157) );
  AOI22_X1 U22842 ( .A1(n19858), .A2(n19956), .B1(n19955), .B2(n19870), .ZN(
        n19856) );
  AOI22_X1 U22843 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19859), .B1(
        n19902), .B2(n19898), .ZN(n19855) );
  OAI211_X1 U22844 ( .C1(n19857), .C2(n19862), .A(n19856), .B(n19855), .ZN(
        P2_U3158) );
  AOI22_X1 U22845 ( .A1(n19858), .A2(n19963), .B1(n19962), .B2(n19870), .ZN(
        n19861) );
  AOI22_X1 U22846 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19859), .B1(
        n19902), .B2(n19903), .ZN(n19860) );
  OAI211_X1 U22847 ( .C1(n19863), .C2(n19862), .A(n19861), .B(n19860), .ZN(
        P2_U3159) );
  INV_X1 U22848 ( .A(n19966), .ZN(n19867) );
  INV_X1 U22849 ( .A(n19902), .ZN(n19866) );
  NAND2_X1 U22850 ( .A1(n19867), .A2(n19866), .ZN(n19869) );
  AOI21_X1 U22851 ( .B1(n19869), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19868), 
        .ZN(n19874) );
  NAND3_X1 U22852 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19917) );
  NOR2_X1 U22853 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19917), .ZN(
        n19901) );
  NOR2_X1 U22854 ( .A1(n19901), .A2(n19870), .ZN(n19878) );
  AOI21_X1 U22855 ( .B1(n19875), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19871) );
  OAI21_X1 U22856 ( .B1(n19871), .B2(n19901), .A(n19919), .ZN(n19872) );
  AOI22_X1 U22857 ( .A1(n19966), .A2(n19873), .B1(n19912), .B2(n19901), .ZN(
        n19881) );
  INV_X1 U22858 ( .A(n19874), .ZN(n19879) );
  INV_X1 U22859 ( .A(n19875), .ZN(n19876) );
  OAI21_X1 U22860 ( .B1(n19876), .B2(n19901), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19877) );
  AOI22_X1 U22861 ( .A1(n19913), .A2(n19904), .B1(n19902), .B2(n19921), .ZN(
        n19880) );
  OAI211_X1 U22862 ( .C1(n19908), .C2(n19882), .A(n19881), .B(n19880), .ZN(
        P2_U3160) );
  AOI22_X1 U22863 ( .A1(n19927), .A2(n19902), .B1(n19925), .B2(n19901), .ZN(
        n19885) );
  AOI22_X1 U22864 ( .A1(n19926), .A2(n19904), .B1(n19966), .B2(n19883), .ZN(
        n19884) );
  OAI211_X1 U22865 ( .C1(n19908), .C2(n12425), .A(n19885), .B(n19884), .ZN(
        P2_U3161) );
  AOI22_X1 U22866 ( .A1(n19966), .A2(n19886), .B1(n19931), .B2(n19901), .ZN(
        n19888) );
  AOI22_X1 U22867 ( .A1(n19932), .A2(n19904), .B1(n19902), .B2(n19933), .ZN(
        n19887) );
  OAI211_X1 U22868 ( .C1(n19908), .C2(n12200), .A(n19888), .B(n19887), .ZN(
        P2_U3162) );
  AOI22_X1 U22869 ( .A1(n19966), .A2(n19889), .B1(n19937), .B2(n19901), .ZN(
        n19891) );
  AOI22_X1 U22870 ( .A1(n19938), .A2(n19904), .B1(n19902), .B2(n19939), .ZN(
        n19890) );
  OAI211_X1 U22871 ( .C1(n19908), .C2(n12474), .A(n19891), .B(n19890), .ZN(
        P2_U3163) );
  AOI22_X1 U22872 ( .A1(n19966), .A2(n19892), .B1(n19943), .B2(n19901), .ZN(
        n19894) );
  AOI22_X1 U22873 ( .A1(n19944), .A2(n19904), .B1(n19902), .B2(n19945), .ZN(
        n19893) );
  OAI211_X1 U22874 ( .C1(n19908), .C2(n12245), .A(n19894), .B(n19893), .ZN(
        P2_U3164) );
  AOI22_X1 U22875 ( .A1(n19951), .A2(n19902), .B1(n19949), .B2(n19901), .ZN(
        n19897) );
  AOI22_X1 U22876 ( .A1(n19950), .A2(n19904), .B1(n19966), .B2(n19895), .ZN(
        n19896) );
  OAI211_X1 U22877 ( .C1(n19908), .C2(n12527), .A(n19897), .B(n19896), .ZN(
        P2_U3165) );
  AOI22_X1 U22878 ( .A1(n19966), .A2(n19898), .B1(n19955), .B2(n19901), .ZN(
        n19900) );
  AOI22_X1 U22879 ( .A1(n19956), .A2(n19904), .B1(n19902), .B2(n19957), .ZN(
        n19899) );
  OAI211_X1 U22880 ( .C1(n19908), .C2(n12571), .A(n19900), .B(n19899), .ZN(
        P2_U3166) );
  INV_X1 U22881 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n19907) );
  AOI22_X1 U22882 ( .A1(n19965), .A2(n19902), .B1(n19962), .B2(n19901), .ZN(
        n19906) );
  AOI22_X1 U22883 ( .A1(n19963), .A2(n19904), .B1(n19966), .B2(n19903), .ZN(
        n19905) );
  OAI211_X1 U22884 ( .C1(n19908), .C2(n19907), .A(n19906), .B(n19905), .ZN(
        P2_U3167) );
  INV_X1 U22885 ( .A(n12521), .ZN(n19909) );
  NOR3_X1 U22886 ( .A1(n19909), .A2(n19961), .A3(n19591), .ZN(n19916) );
  INV_X1 U22887 ( .A(n19917), .ZN(n19910) );
  AOI21_X1 U22888 ( .B1(n20089), .B2(n19910), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19911) );
  NOR2_X1 U22889 ( .A1(n19916), .A2(n19911), .ZN(n19964) );
  AOI22_X1 U22890 ( .A1(n19964), .A2(n19913), .B1(n19912), .B2(n19961), .ZN(
        n19923) );
  NAND2_X1 U22891 ( .A1(n19915), .A2(n19914), .ZN(n19918) );
  AOI21_X1 U22892 ( .B1(n19918), .B2(n19917), .A(n19916), .ZN(n19920) );
  OAI211_X1 U22893 ( .C1(n19961), .C2(n20089), .A(n19920), .B(n19919), .ZN(
        n19967) );
  AOI22_X1 U22894 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19967), .B1(
        n19966), .B2(n19921), .ZN(n19922) );
  OAI211_X1 U22895 ( .C1(n19924), .C2(n19970), .A(n19923), .B(n19922), .ZN(
        P2_U3168) );
  AOI22_X1 U22896 ( .A1(n19964), .A2(n19926), .B1(n19925), .B2(n19961), .ZN(
        n19929) );
  AOI22_X1 U22897 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19967), .B1(
        n19966), .B2(n19927), .ZN(n19928) );
  OAI211_X1 U22898 ( .C1(n19930), .C2(n19970), .A(n19929), .B(n19928), .ZN(
        P2_U3169) );
  AOI22_X1 U22899 ( .A1(n19964), .A2(n19932), .B1(n19931), .B2(n19961), .ZN(
        n19935) );
  AOI22_X1 U22900 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19967), .B1(
        n19966), .B2(n19933), .ZN(n19934) );
  OAI211_X1 U22901 ( .C1(n19936), .C2(n19970), .A(n19935), .B(n19934), .ZN(
        P2_U3170) );
  AOI22_X1 U22902 ( .A1(n19964), .A2(n19938), .B1(n19937), .B2(n19961), .ZN(
        n19941) );
  AOI22_X1 U22903 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19967), .B1(
        n19966), .B2(n19939), .ZN(n19940) );
  OAI211_X1 U22904 ( .C1(n19942), .C2(n19970), .A(n19941), .B(n19940), .ZN(
        P2_U3171) );
  AOI22_X1 U22905 ( .A1(n19964), .A2(n19944), .B1(n19943), .B2(n19961), .ZN(
        n19947) );
  AOI22_X1 U22906 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19967), .B1(
        n19966), .B2(n19945), .ZN(n19946) );
  OAI211_X1 U22907 ( .C1(n19948), .C2(n19970), .A(n19947), .B(n19946), .ZN(
        P2_U3172) );
  AOI22_X1 U22908 ( .A1(n19964), .A2(n19950), .B1(n19949), .B2(n19961), .ZN(
        n19953) );
  AOI22_X1 U22909 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19967), .B1(
        n19966), .B2(n19951), .ZN(n19952) );
  OAI211_X1 U22910 ( .C1(n19954), .C2(n19970), .A(n19953), .B(n19952), .ZN(
        P2_U3173) );
  AOI22_X1 U22911 ( .A1(n19964), .A2(n19956), .B1(n19955), .B2(n19961), .ZN(
        n19959) );
  AOI22_X1 U22912 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19967), .B1(
        n19966), .B2(n19957), .ZN(n19958) );
  OAI211_X1 U22913 ( .C1(n19960), .C2(n19970), .A(n19959), .B(n19958), .ZN(
        P2_U3174) );
  AOI22_X1 U22914 ( .A1(n19964), .A2(n19963), .B1(n19962), .B2(n19961), .ZN(
        n19969) );
  AOI22_X1 U22915 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19967), .B1(
        n19966), .B2(n19965), .ZN(n19968) );
  OAI211_X1 U22916 ( .C1(n19971), .C2(n19970), .A(n19969), .B(n19968), .ZN(
        P2_U3175) );
  INV_X1 U22917 ( .A(n19976), .ZN(n19973) );
  OAI211_X1 U22918 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n20114), .A(n19973), 
        .B(n19972), .ZN(n19979) );
  NOR2_X1 U22919 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19974), .ZN(n19975) );
  OAI211_X1 U22920 ( .C1(n19976), .C2(n19975), .A(P2_STATE2_REG_1__SCAN_IN), 
        .B(n20118), .ZN(n19978) );
  OAI211_X1 U22921 ( .C1(n19980), .C2(n19979), .A(n19978), .B(n19977), .ZN(
        P2_U3177) );
  AND2_X1 U22922 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n9638), .ZN(P2_U3179) );
  AND2_X1 U22923 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19981), .ZN(
        P2_U3180) );
  AND2_X1 U22924 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n9638), .ZN(P2_U3181) );
  AND2_X1 U22925 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n9638), .ZN(P2_U3182) );
  AND2_X1 U22926 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n9638), .ZN(P2_U3183) );
  AND2_X1 U22927 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n9638), .ZN(P2_U3184) );
  AND2_X1 U22928 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n9638), .ZN(P2_U3185) );
  AND2_X1 U22929 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n9638), .ZN(P2_U3186) );
  AND2_X1 U22930 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19981), .ZN(
        P2_U3187) );
  AND2_X1 U22931 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n9638), .ZN(P2_U3188) );
  AND2_X1 U22932 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19981), .ZN(
        P2_U3189) );
  AND2_X1 U22933 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n9638), .ZN(P2_U3190) );
  AND2_X1 U22934 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19981), .ZN(
        P2_U3191) );
  AND2_X1 U22935 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n9638), .ZN(P2_U3192) );
  AND2_X1 U22936 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19981), .ZN(
        P2_U3193) );
  AND2_X1 U22937 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n9638), .ZN(P2_U3194) );
  AND2_X1 U22938 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19981), .ZN(
        P2_U3195) );
  AND2_X1 U22939 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n9638), .ZN(P2_U3196) );
  AND2_X1 U22940 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n9638), .ZN(P2_U3197) );
  AND2_X1 U22941 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n9638), .ZN(P2_U3198) );
  AND2_X1 U22942 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n9638), .ZN(P2_U3199) );
  AND2_X1 U22943 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19981), .ZN(
        P2_U3200) );
  AND2_X1 U22944 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19981), .ZN(P2_U3201) );
  AND2_X1 U22945 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n9638), .ZN(P2_U3202)
         );
  AND2_X1 U22946 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19981), .ZN(P2_U3203) );
  AND2_X1 U22947 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n9638), .ZN(P2_U3204)
         );
  AND2_X1 U22948 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19981), .ZN(P2_U3205) );
  AND2_X1 U22949 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n9638), .ZN(P2_U3206)
         );
  AND2_X1 U22950 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19981), .ZN(P2_U3207) );
  AND2_X1 U22951 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n9638), .ZN(P2_U3208)
         );
  NAND2_X1 U22952 ( .A1(n20118), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19994) );
  NAND3_X1 U22953 ( .A1(n19994), .A2(P2_STATE_REG_0__SCAN_IN), .A3(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19982) );
  INV_X1 U22954 ( .A(NA), .ZN(n20762) );
  OAI21_X1 U22955 ( .B1(n20762), .B2(n19987), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19996) );
  NAND2_X1 U22956 ( .A1(n19982), .A2(n19996), .ZN(n19983) );
  OAI221_X1 U22957 ( .B1(n19984), .B2(P2_REQUESTPENDING_REG_SCAN_IN), .C1(
        n19984), .C2(n21016), .A(n19983), .ZN(P2_U3209) );
  AND2_X1 U22958 ( .A1(n19985), .A2(n19994), .ZN(n19989) );
  NOR2_X1 U22959 ( .A1(HOLD), .A2(n19986), .ZN(n19995) );
  OAI211_X1 U22960 ( .C1(n19995), .C2(n19997), .A(
        P2_REQUESTPENDING_REG_SCAN_IN), .B(n19987), .ZN(n19988) );
  OAI211_X1 U22961 ( .C1(n19990), .C2(n21016), .A(n19989), .B(n19988), .ZN(
        P2_U3210) );
  OAI22_X1 U22962 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19991), .B1(NA), 
        .B2(n19994), .ZN(n19992) );
  OAI211_X1 U22963 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19992), .ZN(n19993) );
  OAI221_X1 U22964 ( .B1(n19996), .B2(n19995), .C1(n19996), .C2(n19994), .A(
        n19993), .ZN(P2_U3211) );
  OAI222_X1 U22965 ( .A1(n20043), .A2(n20000), .B1(n19998), .B2(n20034), .C1(
        n10624), .C2(n20038), .ZN(P2_U3212) );
  OAI222_X1 U22966 ( .A1(n20038), .A2(n20000), .B1(n19999), .B2(n20034), .C1(
        n10684), .C2(n20043), .ZN(P2_U3213) );
  OAI222_X1 U22967 ( .A1(n20038), .A2(n10684), .B1(n20001), .B2(n20034), .C1(
        n10695), .C2(n20043), .ZN(P2_U3214) );
  OAI222_X1 U22968 ( .A1(n20043), .A2(n15426), .B1(n20002), .B2(n20034), .C1(
        n10695), .C2(n20038), .ZN(P2_U3215) );
  OAI222_X1 U22969 ( .A1(n20043), .A2(n10860), .B1(n20003), .B2(n20034), .C1(
        n15426), .C2(n20038), .ZN(P2_U3216) );
  OAI222_X1 U22970 ( .A1(n20043), .A2(n15402), .B1(n20004), .B2(n20034), .C1(
        n10860), .C2(n20038), .ZN(P2_U3217) );
  OAI222_X1 U22971 ( .A1(n20043), .A2(n10710), .B1(n20005), .B2(n20034), .C1(
        n15402), .C2(n20038), .ZN(P2_U3218) );
  OAI222_X1 U22972 ( .A1(n20043), .A2(n15625), .B1(n20006), .B2(n20034), .C1(
        n10710), .C2(n20038), .ZN(P2_U3219) );
  OAI222_X1 U22973 ( .A1(n20043), .A2(n10905), .B1(n20007), .B2(n20034), .C1(
        n15625), .C2(n20038), .ZN(P2_U3220) );
  OAI222_X1 U22974 ( .A1(n20043), .A2(n10717), .B1(n20008), .B2(n20034), .C1(
        n10905), .C2(n20038), .ZN(P2_U3221) );
  OAI222_X1 U22975 ( .A1(n20043), .A2(n10920), .B1(n20009), .B2(n20034), .C1(
        n10717), .C2(n20038), .ZN(P2_U3222) );
  OAI222_X1 U22976 ( .A1(n20043), .A2(n20011), .B1(n20010), .B2(n20034), .C1(
        n10920), .C2(n20038), .ZN(P2_U3223) );
  OAI222_X1 U22977 ( .A1(n20043), .A2(n10947), .B1(n20012), .B2(n20034), .C1(
        n20011), .C2(n20038), .ZN(P2_U3224) );
  OAI222_X1 U22978 ( .A1(n20043), .A2(n10731), .B1(n20013), .B2(n20034), .C1(
        n10947), .C2(n20038), .ZN(P2_U3225) );
  OAI222_X1 U22979 ( .A1(n20043), .A2(n15584), .B1(n20014), .B2(n20034), .C1(
        n10731), .C2(n20038), .ZN(P2_U3226) );
  OAI222_X1 U22980 ( .A1(n20043), .A2(n15575), .B1(n20015), .B2(n20034), .C1(
        n15584), .C2(n20038), .ZN(P2_U3227) );
  OAI222_X1 U22981 ( .A1(n20043), .A2(n20017), .B1(n20016), .B2(n20034), .C1(
        n15575), .C2(n20038), .ZN(P2_U3228) );
  OAI222_X1 U22982 ( .A1(n20043), .A2(n15357), .B1(n20018), .B2(n20034), .C1(
        n20017), .C2(n20038), .ZN(P2_U3229) );
  OAI222_X1 U22983 ( .A1(n20043), .A2(n20020), .B1(n20019), .B2(n20034), .C1(
        n15357), .C2(n20038), .ZN(P2_U3230) );
  OAI222_X1 U22984 ( .A1(n20043), .A2(n20022), .B1(n20021), .B2(n20034), .C1(
        n20020), .C2(n20038), .ZN(P2_U3231) );
  OAI222_X1 U22985 ( .A1(n20043), .A2(n20024), .B1(n20023), .B2(n20034), .C1(
        n20022), .C2(n20038), .ZN(P2_U3232) );
  OAI222_X1 U22986 ( .A1(n20043), .A2(n20026), .B1(n20025), .B2(n20034), .C1(
        n20024), .C2(n20038), .ZN(P2_U3233) );
  OAI222_X1 U22987 ( .A1(n20043), .A2(n20028), .B1(n20027), .B2(n20034), .C1(
        n20026), .C2(n20038), .ZN(P2_U3234) );
  OAI222_X1 U22988 ( .A1(n20043), .A2(n20030), .B1(n20029), .B2(n20034), .C1(
        n20028), .C2(n20038), .ZN(P2_U3235) );
  INV_X1 U22989 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20032) );
  OAI222_X1 U22990 ( .A1(n20043), .A2(n20032), .B1(n20031), .B2(n20034), .C1(
        n20030), .C2(n20038), .ZN(P2_U3236) );
  OAI222_X1 U22991 ( .A1(n20043), .A2(n10986), .B1(n20033), .B2(n20034), .C1(
        n20032), .C2(n20038), .ZN(P2_U3237) );
  OAI222_X1 U22992 ( .A1(n20038), .A2(n10986), .B1(n20035), .B2(n20034), .C1(
        n20036), .C2(n20043), .ZN(P2_U3238) );
  OAI222_X1 U22993 ( .A1(n20043), .A2(n15249), .B1(n20037), .B2(n20034), .C1(
        n20036), .C2(n20038), .ZN(P2_U3239) );
  OAI222_X1 U22994 ( .A1(n20043), .A2(n20040), .B1(n20039), .B2(n20034), .C1(
        n15249), .C2(n20038), .ZN(P2_U3240) );
  INV_X1 U22995 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20041) );
  OAI222_X1 U22996 ( .A1(n20043), .A2(n20042), .B1(n20041), .B2(n20034), .C1(
        n20040), .C2(n20038), .ZN(P2_U3241) );
  INV_X1 U22997 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n20044) );
  AOI22_X1 U22998 ( .A1(n20034), .A2(n20045), .B1(n20044), .B2(n20098), .ZN(
        P2_U3585) );
  MUX2_X1 U22999 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n20034), .Z(P2_U3586) );
  INV_X1 U23000 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n20046) );
  AOI22_X1 U23001 ( .A1(n20034), .A2(n20047), .B1(n20046), .B2(n20098), .ZN(
        P2_U3587) );
  INV_X1 U23002 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n20048) );
  AOI22_X1 U23003 ( .A1(n20034), .A2(n20049), .B1(n20048), .B2(n20098), .ZN(
        P2_U3588) );
  AOI21_X1 U23004 ( .B1(n9638), .B2(n20051), .A(n20050), .ZN(P2_U3591) );
  OAI21_X1 U23005 ( .B1(n20054), .B2(n20053), .A(n20052), .ZN(P2_U3592) );
  INV_X1 U23006 ( .A(n20055), .ZN(n20057) );
  AOI222_X1 U23007 ( .A1(n20060), .A2(n20059), .B1(n20082), .B2(n20058), .C1(
        n20057), .C2(n20056), .ZN(n20062) );
  AOI22_X1 U23008 ( .A1(n20063), .A2(n13539), .B1(n20062), .B2(n20061), .ZN(
        P2_U3600) );
  INV_X1 U23009 ( .A(n20094), .ZN(n20097) );
  AND2_X1 U23010 ( .A1(n20068), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20084) );
  NAND2_X1 U23011 ( .A1(n20064), .A2(n20084), .ZN(n20073) );
  NAND3_X1 U23012 ( .A1(n20082), .A2(n20065), .A3(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20066) );
  NAND2_X1 U23013 ( .A1(n20066), .A2(n20092), .ZN(n20074) );
  NAND2_X1 U23014 ( .A1(n20073), .A2(n20074), .ZN(n20071) );
  AOI222_X1 U23015 ( .A1(n20071), .A2(n20070), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20069), .C1(n20068), .C2(n20067), .ZN(n20072) );
  AOI22_X1 U23016 ( .A1(n20097), .A2(n10331), .B1(n20072), .B2(n20094), .ZN(
        P2_U3602) );
  OAI21_X1 U23017 ( .B1(n20075), .B2(n20074), .A(n20073), .ZN(n20076) );
  AOI21_X1 U23018 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20077), .A(n20076), 
        .ZN(n20078) );
  AOI22_X1 U23019 ( .A1(n20097), .A2(n20079), .B1(n20078), .B2(n20094), .ZN(
        P2_U3603) );
  INV_X1 U23020 ( .A(n20092), .ZN(n20081) );
  NOR2_X1 U23021 ( .A1(n20081), .A2(n20080), .ZN(n20083) );
  MUX2_X1 U23022 ( .A(n20084), .B(n20083), .S(n20082), .Z(n20085) );
  AOI21_X1 U23023 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20086), .A(n20085), 
        .ZN(n20087) );
  AOI22_X1 U23024 ( .A1(n20097), .A2(n20088), .B1(n20087), .B2(n20094), .ZN(
        P2_U3604) );
  NOR2_X1 U23025 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20089), .ZN(
        n20090) );
  AOI211_X1 U23026 ( .C1(n20093), .C2(n20092), .A(n20091), .B(n20090), .ZN(
        n20095) );
  AOI22_X1 U23027 ( .A1(n20097), .A2(n20096), .B1(n20095), .B2(n20094), .ZN(
        P2_U3605) );
  INV_X1 U23028 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20099) );
  AOI22_X1 U23029 ( .A1(n20034), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20099), 
        .B2(n20098), .ZN(P2_U3608) );
  AOI22_X1 U23030 ( .A1(n20103), .A2(n20102), .B1(n20101), .B2(n20100), .ZN(
        n20107) );
  INV_X1 U23031 ( .A(n20104), .ZN(n20105) );
  OAI21_X1 U23032 ( .B1(n20107), .B2(n20106), .A(n20105), .ZN(n20109) );
  MUX2_X1 U23033 ( .A(P2_MORE_REG_SCAN_IN), .B(n20109), .S(n20108), .Z(
        P2_U3609) );
  INV_X1 U23034 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20128) );
  NOR2_X1 U23035 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20110), .ZN(n20112) );
  AOI211_X1 U23036 ( .C1(n20114), .C2(n20113), .A(n20112), .B(n20111), .ZN(
        n20127) );
  NAND3_X1 U23037 ( .A1(n20116), .A2(n20115), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n20120) );
  OAI21_X1 U23038 ( .B1(n20118), .B2(n19591), .A(n20117), .ZN(n20119) );
  OAI21_X1 U23039 ( .B1(n20123), .B2(n20120), .A(n20119), .ZN(n20121) );
  INV_X1 U23040 ( .A(n20121), .ZN(n20126) );
  AOI211_X1 U23041 ( .C1(P2_STATEBS16_REG_SCAN_IN), .C2(n20123), .A(n20122), 
        .B(n10643), .ZN(n20124) );
  NOR2_X1 U23042 ( .A1(n20127), .A2(n20124), .ZN(n20125) );
  AOI22_X1 U23043 ( .A1(n20128), .A2(n20127), .B1(n20126), .B2(n20125), .ZN(
        P2_U3610) );
  MUX2_X1 U23044 ( .A(P2_M_IO_N_REG_SCAN_IN), .B(P2_MEMORYFETCH_REG_SCAN_IN), 
        .S(n20034), .Z(P2_U3611) );
  NOR2_X1 U23045 ( .A1(n20130), .A2(n20129), .ZN(n20132) );
  INV_X1 U23046 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20131) );
  INV_X1 U23047 ( .A(n20854), .ZN(n20855) );
  AOI21_X1 U23048 ( .B1(n20132), .B2(n20131), .A(n20855), .ZN(P1_U2802) );
  INV_X1 U23049 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n21024) );
  NOR2_X1 U23050 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20134) );
  NOR2_X1 U23051 ( .A1(n20855), .A2(n20134), .ZN(n20133) );
  AOI22_X1 U23052 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(n20855), .B1(n21024), 
        .B2(n20133), .ZN(P1_U2804) );
  AOI21_X1 U23053 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20760), .A(n20855), 
        .ZN(n20831) );
  OAI21_X1 U23054 ( .B1(BS16), .B2(n20134), .A(n20831), .ZN(n20829) );
  OAI21_X1 U23055 ( .B1(n20831), .B2(n20841), .A(n20829), .ZN(P1_U2805) );
  OAI21_X1 U23056 ( .B1(n20136), .B2(n21037), .A(n20135), .ZN(P1_U2806) );
  NOR4_X1 U23057 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20140) );
  NOR4_X1 U23058 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20139) );
  NOR4_X1 U23059 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20138) );
  NOR4_X1 U23060 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20137) );
  NAND4_X1 U23061 ( .A1(n20140), .A2(n20139), .A3(n20138), .A4(n20137), .ZN(
        n20146) );
  NOR4_X1 U23062 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20144) );
  AOI211_X1 U23063 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20143) );
  NOR4_X1 U23064 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20142) );
  NOR4_X1 U23065 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20141) );
  NAND4_X1 U23066 ( .A1(n20144), .A2(n20143), .A3(n20142), .A4(n20141), .ZN(
        n20145) );
  NOR2_X1 U23067 ( .A1(n20146), .A2(n20145), .ZN(n20838) );
  INV_X1 U23068 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20824) );
  NOR3_X1 U23069 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20148) );
  OAI21_X1 U23070 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20148), .A(n20838), .ZN(
        n20147) );
  OAI21_X1 U23071 ( .B1(n20838), .B2(n20824), .A(n20147), .ZN(P1_U2807) );
  INV_X1 U23072 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20830) );
  AOI21_X1 U23073 ( .B1(n20832), .B2(n20830), .A(n20148), .ZN(n20149) );
  INV_X1 U23074 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20821) );
  INV_X1 U23075 ( .A(n20838), .ZN(n20834) );
  AOI22_X1 U23076 ( .A1(n20838), .A2(n20149), .B1(n20821), .B2(n20834), .ZN(
        P1_U2808) );
  INV_X1 U23077 ( .A(n20205), .ZN(n20152) );
  AOI22_X1 U23078 ( .A1(n20152), .A2(n20151), .B1(n20197), .B2(n20150), .ZN(
        n20160) );
  AOI22_X1 U23079 ( .A1(n20153), .A2(n20183), .B1(n20175), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n20154) );
  OAI211_X1 U23080 ( .C1(n20177), .C2(n20155), .A(n20154), .B(n20191), .ZN(
        n20156) );
  AOI221_X1 U23081 ( .B1(n20158), .B2(n13889), .C1(n20157), .C2(
        P1_REIP_REG_9__SCAN_IN), .A(n20156), .ZN(n20159) );
  NAND2_X1 U23082 ( .A1(n20160), .A2(n20159), .ZN(P1_U2831) );
  INV_X1 U23083 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20168) );
  NOR2_X1 U23084 ( .A1(n20189), .A2(n20163), .ZN(n20164) );
  AOI211_X1 U23085 ( .C1(n20175), .C2(P1_EBX_REG_7__SCAN_IN), .A(n20174), .B(
        n20164), .ZN(n20167) );
  NAND2_X1 U23086 ( .A1(n20165), .A2(n20183), .ZN(n20166) );
  OAI211_X1 U23087 ( .C1(n20168), .C2(n20177), .A(n20167), .B(n20166), .ZN(
        n20171) );
  NOR2_X1 U23088 ( .A1(n20169), .A2(n20178), .ZN(n20170) );
  AOI211_X1 U23089 ( .C1(P1_REIP_REG_7__SCAN_IN), .C2(n10268), .A(n20171), .B(
        n20170), .ZN(n20172) );
  OAI21_X1 U23090 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(n20173), .A(n20172), .ZN(
        P1_U2833) );
  AOI21_X1 U23091 ( .B1(n20175), .B2(P1_EBX_REG_6__SCAN_IN), .A(n20174), .ZN(
        n20176) );
  OAI21_X1 U23092 ( .B1(n20177), .B2(n11325), .A(n20176), .ZN(n20181) );
  NOR2_X1 U23093 ( .A1(n20179), .A2(n20178), .ZN(n20180) );
  AOI211_X1 U23094 ( .C1(n20183), .C2(n20182), .A(n20181), .B(n20180), .ZN(
        n20187) );
  INV_X1 U23095 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20775) );
  AOI21_X1 U23096 ( .B1(n20185), .B2(n20184), .A(n20775), .ZN(n20203) );
  OAI21_X1 U23097 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(n20203), .A(n10268), .ZN(
        n20186) );
  OAI211_X1 U23098 ( .C1(n20189), .C2(n20188), .A(n20187), .B(n20186), .ZN(
        P1_U2834) );
  NOR2_X1 U23099 ( .A1(n20190), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n20202) );
  OAI21_X1 U23100 ( .B1(n20192), .B2(n20215), .A(n20191), .ZN(n20195) );
  NOR2_X1 U23101 ( .A1(n20210), .A2(n20193), .ZN(n20194) );
  AOI211_X1 U23102 ( .C1(n20196), .C2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n20195), .B(n20194), .ZN(n20201) );
  AOI22_X1 U23103 ( .A1(n20213), .A2(n20199), .B1(n20198), .B2(n20197), .ZN(
        n20200) );
  OAI211_X1 U23104 ( .C1(n20203), .C2(n20202), .A(n20201), .B(n20200), .ZN(
        P1_U2835) );
  OAI22_X1 U23105 ( .A1(n20205), .A2(n14420), .B1(n20209), .B2(n20204), .ZN(
        n20206) );
  INV_X1 U23106 ( .A(n20206), .ZN(n20207) );
  OAI21_X1 U23107 ( .B1(n20216), .B2(n20208), .A(n20207), .ZN(P1_U2863) );
  NOR2_X1 U23108 ( .A1(n20210), .A2(n20209), .ZN(n20211) );
  AOI21_X1 U23109 ( .B1(n20213), .B2(n20212), .A(n20211), .ZN(n20214) );
  OAI21_X1 U23110 ( .B1(n20216), .B2(n20215), .A(n20214), .ZN(P1_U2867) );
  AOI22_X1 U23111 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20220), .B1(n16114), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20217) );
  OAI21_X1 U23112 ( .B1(n20219), .B2(n20218), .A(n20217), .ZN(P1_U2921) );
  AOI22_X1 U23113 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20221) );
  OAI21_X1 U23114 ( .B1(n14499), .B2(n20246), .A(n20221), .ZN(P1_U2922) );
  INV_X1 U23115 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20223) );
  AOI22_X1 U23116 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20222) );
  OAI21_X1 U23117 ( .B1(n20223), .B2(n20246), .A(n20222), .ZN(P1_U2923) );
  INV_X1 U23118 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20225) );
  AOI22_X1 U23119 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20224) );
  OAI21_X1 U23120 ( .B1(n20225), .B2(n20246), .A(n20224), .ZN(P1_U2924) );
  INV_X1 U23121 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20227) );
  AOI22_X1 U23122 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20226) );
  OAI21_X1 U23123 ( .B1(n20227), .B2(n20246), .A(n20226), .ZN(P1_U2925) );
  INV_X1 U23124 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20229) );
  AOI22_X1 U23125 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20228) );
  OAI21_X1 U23126 ( .B1(n20229), .B2(n20246), .A(n20228), .ZN(P1_U2926) );
  INV_X1 U23127 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20231) );
  AOI22_X1 U23128 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20230) );
  OAI21_X1 U23129 ( .B1(n20231), .B2(n20246), .A(n20230), .ZN(P1_U2927) );
  INV_X1 U23130 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20233) );
  AOI22_X1 U23131 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20232) );
  OAI21_X1 U23132 ( .B1(n20233), .B2(n20246), .A(n20232), .ZN(P1_U2928) );
  AOI22_X1 U23133 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20234) );
  OAI21_X1 U23134 ( .B1(n11386), .B2(n20246), .A(n20234), .ZN(P1_U2929) );
  AOI22_X1 U23135 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20235) );
  OAI21_X1 U23136 ( .B1(n11329), .B2(n20246), .A(n20235), .ZN(P1_U2930) );
  AOI22_X1 U23137 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20236) );
  OAI21_X1 U23138 ( .B1(n11310), .B2(n20246), .A(n20236), .ZN(P1_U2931) );
  AOI22_X1 U23139 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20237) );
  OAI21_X1 U23140 ( .B1(n20238), .B2(n20246), .A(n20237), .ZN(P1_U2932) );
  AOI22_X1 U23141 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20239) );
  OAI21_X1 U23142 ( .B1(n20240), .B2(n20246), .A(n20239), .ZN(P1_U2933) );
  AOI22_X1 U23143 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20241) );
  OAI21_X1 U23144 ( .B1(n20242), .B2(n20246), .A(n20241), .ZN(P1_U2934) );
  AOI22_X1 U23145 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20243) );
  OAI21_X1 U23146 ( .B1(n20244), .B2(n20246), .A(n20243), .ZN(P1_U2935) );
  AOI22_X1 U23147 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20851), .B1(n16114), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20245) );
  OAI21_X1 U23148 ( .B1(n20247), .B2(n20246), .A(n20245), .ZN(P1_U2936) );
  AOI22_X1 U23149 ( .A1(n20275), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20274), .ZN(n20249) );
  NAND2_X1 U23150 ( .A1(n20260), .A2(n20248), .ZN(n20262) );
  NAND2_X1 U23151 ( .A1(n20249), .A2(n20262), .ZN(P1_U2945) );
  AOI22_X1 U23152 ( .A1(n20275), .A2(P1_EAX_REG_25__SCAN_IN), .B1(n20274), 
        .B2(P1_UWORD_REG_9__SCAN_IN), .ZN(n20251) );
  NAND2_X1 U23153 ( .A1(n20260), .A2(n20250), .ZN(n20264) );
  NAND2_X1 U23154 ( .A1(n20251), .A2(n20264), .ZN(P1_U2946) );
  AOI22_X1 U23155 ( .A1(n20275), .A2(P1_EAX_REG_27__SCAN_IN), .B1(n20274), 
        .B2(P1_UWORD_REG_11__SCAN_IN), .ZN(n20253) );
  NAND2_X1 U23156 ( .A1(n20260), .A2(n20252), .ZN(n20268) );
  NAND2_X1 U23157 ( .A1(n20253), .A2(n20268), .ZN(P1_U2948) );
  AOI22_X1 U23158 ( .A1(n20275), .A2(P1_EAX_REG_28__SCAN_IN), .B1(n20274), 
        .B2(P1_UWORD_REG_12__SCAN_IN), .ZN(n20255) );
  NAND2_X1 U23159 ( .A1(n20260), .A2(n20254), .ZN(n20270) );
  NAND2_X1 U23160 ( .A1(n20255), .A2(n20270), .ZN(P1_U2949) );
  AOI22_X1 U23161 ( .A1(n20275), .A2(P1_EAX_REG_29__SCAN_IN), .B1(n20274), 
        .B2(P1_UWORD_REG_13__SCAN_IN), .ZN(n20257) );
  NAND2_X1 U23162 ( .A1(n20260), .A2(n20256), .ZN(n20272) );
  NAND2_X1 U23163 ( .A1(n20257), .A2(n20272), .ZN(P1_U2950) );
  AOI22_X1 U23164 ( .A1(n20275), .A2(P1_EAX_REG_30__SCAN_IN), .B1(n20274), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n20261) );
  INV_X1 U23165 ( .A(n20258), .ZN(n20259) );
  NAND2_X1 U23166 ( .A1(n20260), .A2(n20259), .ZN(n20276) );
  NAND2_X1 U23167 ( .A1(n20261), .A2(n20276), .ZN(P1_U2951) );
  AOI22_X1 U23168 ( .A1(n20275), .A2(P1_EAX_REG_8__SCAN_IN), .B1(n20274), .B2(
        P1_LWORD_REG_8__SCAN_IN), .ZN(n20263) );
  NAND2_X1 U23169 ( .A1(n20263), .A2(n20262), .ZN(P1_U2960) );
  AOI22_X1 U23170 ( .A1(n20275), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n20274), .B2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n20265) );
  NAND2_X1 U23171 ( .A1(n20265), .A2(n20264), .ZN(P1_U2961) );
  AOI22_X1 U23172 ( .A1(n20275), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n20274), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n20267) );
  NAND2_X1 U23173 ( .A1(n20267), .A2(n20266), .ZN(P1_U2962) );
  AOI22_X1 U23174 ( .A1(n20275), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20274), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n20269) );
  NAND2_X1 U23175 ( .A1(n20269), .A2(n20268), .ZN(P1_U2963) );
  AOI22_X1 U23176 ( .A1(n20275), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n20274), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20271) );
  NAND2_X1 U23177 ( .A1(n20271), .A2(n20270), .ZN(P1_U2964) );
  AOI22_X1 U23178 ( .A1(n20275), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20274), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20273) );
  NAND2_X1 U23179 ( .A1(n20273), .A2(n20272), .ZN(P1_U2965) );
  AOI22_X1 U23180 ( .A1(n20275), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n20274), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20277) );
  NAND2_X1 U23181 ( .A1(n20277), .A2(n20276), .ZN(P1_U2966) );
  INV_X1 U23182 ( .A(n20278), .ZN(n20281) );
  INV_X1 U23183 ( .A(n20279), .ZN(n20280) );
  AOI21_X1 U23184 ( .B1(n20282), .B2(n20281), .A(n20280), .ZN(n20292) );
  AOI211_X1 U23185 ( .C1(n20286), .C2(n20285), .A(n20284), .B(n20283), .ZN(
        n20291) );
  INV_X1 U23186 ( .A(n20287), .ZN(n20288) );
  OAI21_X1 U23187 ( .B1(n20289), .B2(n20288), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20290) );
  NAND3_X1 U23188 ( .A1(n20292), .A2(n20291), .A3(n20290), .ZN(P1_U3031) );
  NOR2_X1 U23189 ( .A1(n20294), .A2(n20293), .ZN(P1_U3032) );
  NAND3_X1 U23190 ( .A1(n20528), .A2(n20532), .A3(n20602), .ZN(n20327) );
  NOR2_X1 U23191 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20327), .ZN(
        n20319) );
  AOI22_X1 U23192 ( .A1(n20745), .A2(n20688), .B1(n20680), .B2(n20319), .ZN(
        n20306) );
  OAI21_X1 U23193 ( .B1(n20347), .B2(n20745), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20296) );
  NAND2_X1 U23194 ( .A1(n20296), .A2(n20596), .ZN(n20304) );
  OR2_X1 U23195 ( .A1(n20467), .A2(n20297), .ZN(n20382) );
  NOR2_X1 U23196 ( .A1(n20382), .A2(n20674), .ZN(n20302) );
  INV_X1 U23197 ( .A(n20529), .ZN(n20299) );
  OR2_X1 U23198 ( .A1(n20299), .A2(n20468), .ZN(n20414) );
  INV_X1 U23199 ( .A(n20319), .ZN(n20300) );
  AOI22_X1 U23200 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20414), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n20300), .ZN(n20301) );
  OAI211_X1 U23201 ( .C1(n20304), .C2(n20302), .A(n20536), .B(n20301), .ZN(
        n20321) );
  INV_X1 U23202 ( .A(n20302), .ZN(n20303) );
  INV_X1 U23203 ( .A(n20530), .ZN(n20469) );
  AOI22_X1 U23204 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20321), .B1(
        n20679), .B2(n20320), .ZN(n20305) );
  OAI211_X1 U23205 ( .C1(n20691), .C2(n20324), .A(n20306), .B(n20305), .ZN(
        P1_U3033) );
  AOI22_X1 U23206 ( .A1(n20745), .A2(n20692), .B1(n20735), .B2(n20319), .ZN(
        n20308) );
  AOI22_X1 U23207 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20321), .B1(
        n20734), .B2(n20320), .ZN(n20307) );
  OAI211_X1 U23208 ( .C1(n20695), .C2(n20324), .A(n20308), .B(n20307), .ZN(
        P1_U3034) );
  AOI22_X1 U23209 ( .A1(n20745), .A2(n20696), .B1(n20743), .B2(n20319), .ZN(
        n20310) );
  AOI22_X1 U23210 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20321), .B1(
        n20741), .B2(n20320), .ZN(n20309) );
  OAI211_X1 U23211 ( .C1(n20699), .C2(n20324), .A(n20310), .B(n20309), .ZN(
        P1_U3035) );
  AOI22_X1 U23212 ( .A1(n20745), .A2(n20702), .B1(n20701), .B2(n20319), .ZN(
        n20312) );
  AOI22_X1 U23213 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20321), .B1(
        n20700), .B2(n20320), .ZN(n20311) );
  OAI211_X1 U23214 ( .C1(n9829), .C2(n20324), .A(n20312), .B(n20311), .ZN(
        P1_U3036) );
  AOI22_X1 U23215 ( .A1(n20745), .A2(n20708), .B1(n20707), .B2(n20319), .ZN(
        n20314) );
  AOI22_X1 U23216 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20321), .B1(
        n20706), .B2(n20320), .ZN(n20313) );
  OAI211_X1 U23217 ( .C1(n20711), .C2(n20324), .A(n20314), .B(n20313), .ZN(
        P1_U3037) );
  AOI22_X1 U23218 ( .A1(n20745), .A2(n20714), .B1(n20713), .B2(n20319), .ZN(
        n20316) );
  AOI22_X1 U23219 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20321), .B1(
        n20712), .B2(n20320), .ZN(n20315) );
  OAI211_X1 U23220 ( .C1(n9831), .C2(n20324), .A(n20316), .B(n20315), .ZN(
        P1_U3038) );
  AOI22_X1 U23221 ( .A1(n20745), .A2(n20720), .B1(n20718), .B2(n20319), .ZN(
        n20318) );
  AOI22_X1 U23222 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20321), .B1(
        n20719), .B2(n20320), .ZN(n20317) );
  OAI211_X1 U23223 ( .C1(n20723), .C2(n20324), .A(n20318), .B(n20317), .ZN(
        P1_U3039) );
  AOI22_X1 U23224 ( .A1(n20745), .A2(n20728), .B1(n20725), .B2(n20319), .ZN(
        n20323) );
  AOI22_X1 U23225 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20321), .B1(
        n20727), .B2(n20320), .ZN(n20322) );
  OAI211_X1 U23226 ( .C1(n20733), .C2(n20324), .A(n20323), .B(n20322), .ZN(
        P1_U3040) );
  NOR2_X1 U23227 ( .A1(n20643), .A2(n20327), .ZN(n20345) );
  INV_X1 U23228 ( .A(n20382), .ZN(n20326) );
  INV_X1 U23229 ( .A(n20325), .ZN(n20645) );
  AOI21_X1 U23230 ( .B1(n20326), .B2(n20645), .A(n20345), .ZN(n20328) );
  OAI22_X1 U23231 ( .A1(n20328), .A2(n20678), .B1(n20327), .B2(n20753), .ZN(
        n20346) );
  AOI22_X1 U23232 ( .A1(n20680), .A2(n20345), .B1(n20346), .B2(n20679), .ZN(
        n20332) );
  INV_X1 U23233 ( .A(n20327), .ZN(n20330) );
  OAI211_X1 U23234 ( .C1(n20386), .C2(n20841), .A(n20596), .B(n20328), .ZN(
        n20329) );
  OAI211_X1 U23235 ( .C1(n20596), .C2(n20330), .A(n20650), .B(n20329), .ZN(
        n20348) );
  AOI22_X1 U23236 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20348), .B1(
        n20347), .B2(n20688), .ZN(n20331) );
  OAI211_X1 U23237 ( .C1(n20691), .C2(n20373), .A(n20332), .B(n20331), .ZN(
        P1_U3041) );
  AOI22_X1 U23238 ( .A1(n20735), .A2(n20345), .B1(n20346), .B2(n20734), .ZN(
        n20334) );
  AOI22_X1 U23239 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20348), .B1(
        n20347), .B2(n20692), .ZN(n20333) );
  OAI211_X1 U23240 ( .C1(n20695), .C2(n20373), .A(n20334), .B(n20333), .ZN(
        P1_U3042) );
  AOI22_X1 U23241 ( .A1(n20743), .A2(n20345), .B1(n20346), .B2(n20741), .ZN(
        n20336) );
  AOI22_X1 U23242 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20348), .B1(
        n20347), .B2(n20696), .ZN(n20335) );
  OAI211_X1 U23243 ( .C1(n20699), .C2(n20373), .A(n20336), .B(n20335), .ZN(
        P1_U3043) );
  AOI22_X1 U23244 ( .A1(n20701), .A2(n20345), .B1(n20346), .B2(n20700), .ZN(
        n20338) );
  AOI22_X1 U23245 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20348), .B1(
        n20347), .B2(n20702), .ZN(n20337) );
  OAI211_X1 U23246 ( .C1(n9829), .C2(n20373), .A(n20338), .B(n20337), .ZN(
        P1_U3044) );
  AOI22_X1 U23247 ( .A1(n20707), .A2(n20345), .B1(n20346), .B2(n20706), .ZN(
        n20340) );
  AOI22_X1 U23248 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20348), .B1(
        n20347), .B2(n20708), .ZN(n20339) );
  OAI211_X1 U23249 ( .C1(n20711), .C2(n20373), .A(n20340), .B(n20339), .ZN(
        P1_U3045) );
  AOI22_X1 U23250 ( .A1(n20713), .A2(n20345), .B1(n20346), .B2(n20712), .ZN(
        n20342) );
  AOI22_X1 U23251 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20348), .B1(
        n20347), .B2(n20714), .ZN(n20341) );
  OAI211_X1 U23252 ( .C1(n9831), .C2(n20373), .A(n20342), .B(n20341), .ZN(
        P1_U3046) );
  AOI22_X1 U23253 ( .A1(n20719), .A2(n20346), .B1(n20718), .B2(n20345), .ZN(
        n20344) );
  AOI22_X1 U23254 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20348), .B1(
        n20347), .B2(n20720), .ZN(n20343) );
  OAI211_X1 U23255 ( .C1(n20723), .C2(n20373), .A(n20344), .B(n20343), .ZN(
        P1_U3047) );
  AOI22_X1 U23256 ( .A1(n20727), .A2(n20346), .B1(n20725), .B2(n20345), .ZN(
        n20350) );
  AOI22_X1 U23257 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20348), .B1(
        n20347), .B2(n20728), .ZN(n20349) );
  OAI211_X1 U23258 ( .C1(n20733), .C2(n20373), .A(n20350), .B(n20349), .ZN(
        P1_U3048) );
  NAND3_X1 U23259 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20528), .A3(
        n20532), .ZN(n20387) );
  NOR2_X1 U23260 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20387), .ZN(
        n20374) );
  AOI22_X1 U23261 ( .A1(n20375), .A2(n20688), .B1(n20680), .B2(n20374), .ZN(
        n20360) );
  OAI21_X1 U23262 ( .B1(n20406), .B2(n20375), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20351) );
  NAND2_X1 U23263 ( .A1(n20351), .A2(n20596), .ZN(n20358) );
  NOR2_X1 U23264 ( .A1(n20382), .A2(n13652), .ZN(n20355) );
  INV_X1 U23265 ( .A(n20374), .ZN(n20353) );
  AOI21_X1 U23266 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20353), .A(n20352), 
        .ZN(n20354) );
  OAI211_X1 U23267 ( .C1(n20358), .C2(n20355), .A(n20536), .B(n20354), .ZN(
        n20377) );
  INV_X1 U23268 ( .A(n20355), .ZN(n20357) );
  AOI22_X1 U23269 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20377), .B1(
        n20679), .B2(n20376), .ZN(n20359) );
  OAI211_X1 U23270 ( .C1(n20691), .C2(n20380), .A(n20360), .B(n20359), .ZN(
        P1_U3049) );
  AOI22_X1 U23271 ( .A1(n20375), .A2(n20692), .B1(n20735), .B2(n20374), .ZN(
        n20362) );
  AOI22_X1 U23272 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20377), .B1(
        n20734), .B2(n20376), .ZN(n20361) );
  OAI211_X1 U23273 ( .C1(n20695), .C2(n20380), .A(n20362), .B(n20361), .ZN(
        P1_U3050) );
  AOI22_X1 U23274 ( .A1(n20375), .A2(n20696), .B1(n20743), .B2(n20374), .ZN(
        n20364) );
  AOI22_X1 U23275 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20377), .B1(
        n20741), .B2(n20376), .ZN(n20363) );
  OAI211_X1 U23276 ( .C1(n20699), .C2(n20380), .A(n20364), .B(n20363), .ZN(
        P1_U3051) );
  AOI22_X1 U23277 ( .A1(n20375), .A2(n20702), .B1(n20701), .B2(n20374), .ZN(
        n20366) );
  AOI22_X1 U23278 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20377), .B1(
        n20700), .B2(n20376), .ZN(n20365) );
  OAI211_X1 U23279 ( .C1(n9829), .C2(n20380), .A(n20366), .B(n20365), .ZN(
        P1_U3052) );
  INV_X1 U23280 ( .A(n20708), .ZN(n20510) );
  INV_X1 U23281 ( .A(n20711), .ZN(n20623) );
  AOI22_X1 U23282 ( .A1(n20406), .A2(n20623), .B1(n20374), .B2(n20707), .ZN(
        n20368) );
  AOI22_X1 U23283 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20377), .B1(
        n20706), .B2(n20376), .ZN(n20367) );
  OAI211_X1 U23284 ( .C1(n20510), .C2(n20373), .A(n20368), .B(n20367), .ZN(
        P1_U3053) );
  AOI22_X1 U23285 ( .A1(n20375), .A2(n20714), .B1(n20713), .B2(n20374), .ZN(
        n20370) );
  AOI22_X1 U23286 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20377), .B1(
        n20712), .B2(n20376), .ZN(n20369) );
  OAI211_X1 U23287 ( .C1(n9831), .C2(n20380), .A(n20370), .B(n20369), .ZN(
        P1_U3054) );
  INV_X1 U23288 ( .A(n20720), .ZN(n20516) );
  INV_X1 U23289 ( .A(n20723), .ZN(n20630) );
  AOI22_X1 U23290 ( .A1(n20406), .A2(n20630), .B1(n20374), .B2(n20718), .ZN(
        n20372) );
  AOI22_X1 U23291 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20377), .B1(
        n20719), .B2(n20376), .ZN(n20371) );
  OAI211_X1 U23292 ( .C1(n20516), .C2(n20373), .A(n20372), .B(n20371), .ZN(
        P1_U3055) );
  AOI22_X1 U23293 ( .A1(n20375), .A2(n20728), .B1(n20725), .B2(n20374), .ZN(
        n20379) );
  AOI22_X1 U23294 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20377), .B1(
        n20727), .B2(n20376), .ZN(n20378) );
  OAI211_X1 U23295 ( .C1(n20733), .C2(n20380), .A(n20379), .B(n20378), .ZN(
        P1_U3056) );
  INV_X1 U23296 ( .A(n20387), .ZN(n20384) );
  NAND2_X1 U23297 ( .A1(n11347), .A2(n13425), .ZN(n20564) );
  NOR2_X1 U23298 ( .A1(n20562), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20405) );
  INV_X1 U23299 ( .A(n20405), .ZN(n20381) );
  OAI21_X1 U23300 ( .B1(n20382), .B2(n20564), .A(n20381), .ZN(n20389) );
  AOI21_X1 U23301 ( .B1(n20386), .B2(n20596), .A(n20568), .ZN(n20390) );
  INV_X1 U23302 ( .A(n20390), .ZN(n20383) );
  INV_X1 U23303 ( .A(n20691), .ZN(n20603) );
  AOI22_X1 U23304 ( .A1(n20435), .A2(n20603), .B1(n20405), .B2(n20680), .ZN(
        n20392) );
  NAND2_X1 U23305 ( .A1(n20678), .A2(n20387), .ZN(n20388) );
  OAI211_X1 U23306 ( .C1(n20390), .C2(n20389), .A(n20650), .B(n20388), .ZN(
        n20407) );
  AOI22_X1 U23307 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20407), .B1(
        n20406), .B2(n20688), .ZN(n20391) );
  OAI211_X1 U23308 ( .C1(n20410), .C2(n20613), .A(n20392), .B(n20391), .ZN(
        P1_U3057) );
  AOI22_X1 U23309 ( .A1(n20406), .A2(n20692), .B1(n20735), .B2(n20405), .ZN(
        n20394) );
  INV_X1 U23310 ( .A(n20695), .ZN(n20736) );
  AOI22_X1 U23311 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20407), .B1(
        n20435), .B2(n20736), .ZN(n20393) );
  OAI211_X1 U23312 ( .C1(n20410), .C2(n20616), .A(n20394), .B(n20393), .ZN(
        P1_U3058) );
  INV_X1 U23313 ( .A(n20699), .ZN(n20744) );
  AOI22_X1 U23314 ( .A1(n20435), .A2(n20744), .B1(n20405), .B2(n20743), .ZN(
        n20396) );
  AOI22_X1 U23315 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20407), .B1(
        n20406), .B2(n20696), .ZN(n20395) );
  OAI211_X1 U23316 ( .C1(n20410), .C2(n20619), .A(n20396), .B(n20395), .ZN(
        P1_U3059) );
  AOI22_X1 U23317 ( .A1(n20406), .A2(n20702), .B1(n20701), .B2(n20405), .ZN(
        n20398) );
  AOI22_X1 U23318 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20407), .B1(
        n20435), .B2(n9828), .ZN(n20397) );
  OAI211_X1 U23319 ( .C1(n20410), .C2(n20622), .A(n20398), .B(n20397), .ZN(
        P1_U3060) );
  AOI22_X1 U23320 ( .A1(n20406), .A2(n20708), .B1(n20707), .B2(n20405), .ZN(
        n20400) );
  AOI22_X1 U23321 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20407), .B1(
        n20435), .B2(n20623), .ZN(n20399) );
  OAI211_X1 U23322 ( .C1(n20410), .C2(n20626), .A(n20400), .B(n20399), .ZN(
        P1_U3061) );
  AOI22_X1 U23323 ( .A1(n20406), .A2(n20714), .B1(n20713), .B2(n20405), .ZN(
        n20402) );
  AOI22_X1 U23324 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20407), .B1(
        n20435), .B2(n9830), .ZN(n20401) );
  OAI211_X1 U23325 ( .C1(n20410), .C2(n20629), .A(n20402), .B(n20401), .ZN(
        P1_U3062) );
  INV_X1 U23326 ( .A(n20719), .ZN(n20633) );
  AOI22_X1 U23327 ( .A1(n20435), .A2(n20630), .B1(n20405), .B2(n20718), .ZN(
        n20404) );
  AOI22_X1 U23328 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20407), .B1(
        n20406), .B2(n20720), .ZN(n20403) );
  OAI211_X1 U23329 ( .C1(n20410), .C2(n20633), .A(n20404), .B(n20403), .ZN(
        P1_U3063) );
  INV_X1 U23330 ( .A(n20727), .ZN(n20640) );
  AOI22_X1 U23331 ( .A1(n20406), .A2(n20728), .B1(n20725), .B2(n20405), .ZN(
        n20409) );
  INV_X1 U23332 ( .A(n20733), .ZN(n20635) );
  AOI22_X1 U23333 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20407), .B1(
        n20435), .B2(n20635), .ZN(n20408) );
  OAI211_X1 U23334 ( .C1(n20410), .C2(n20640), .A(n20409), .B(n20408), .ZN(
        P1_U3064) );
  INV_X1 U23335 ( .A(n20442), .ZN(n20412) );
  NAND3_X1 U23336 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20528), .A3(
        n20602), .ZN(n20440) );
  NOR2_X1 U23337 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20440), .ZN(
        n20433) );
  INV_X1 U23338 ( .A(n20413), .ZN(n20439) );
  NAND2_X1 U23339 ( .A1(n20439), .A2(n13652), .ZN(n20416) );
  OAI22_X1 U23340 ( .A1(n20416), .A2(n20678), .B1(n20414), .B2(n20676), .ZN(
        n20434) );
  AOI22_X1 U23341 ( .A1(n20680), .A2(n20433), .B1(n20679), .B2(n20434), .ZN(
        n20420) );
  INV_X1 U23342 ( .A(n20465), .ZN(n20415) );
  OAI21_X1 U23343 ( .B1(n20435), .B2(n20415), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20417) );
  NAND2_X1 U23344 ( .A1(n20417), .A2(n20416), .ZN(n20418) );
  AOI22_X1 U23345 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20436), .B1(
        n20435), .B2(n20688), .ZN(n20419) );
  OAI211_X1 U23346 ( .C1(n20691), .C2(n20465), .A(n20420), .B(n20419), .ZN(
        P1_U3065) );
  AOI22_X1 U23347 ( .A1(n20735), .A2(n20433), .B1(n20734), .B2(n20434), .ZN(
        n20422) );
  AOI22_X1 U23348 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20436), .B1(
        n20435), .B2(n20692), .ZN(n20421) );
  OAI211_X1 U23349 ( .C1(n20695), .C2(n20465), .A(n20422), .B(n20421), .ZN(
        P1_U3066) );
  AOI22_X1 U23350 ( .A1(n20743), .A2(n20433), .B1(n20741), .B2(n20434), .ZN(
        n20424) );
  AOI22_X1 U23351 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20436), .B1(
        n20435), .B2(n20696), .ZN(n20423) );
  OAI211_X1 U23352 ( .C1(n20699), .C2(n20465), .A(n20424), .B(n20423), .ZN(
        P1_U3067) );
  AOI22_X1 U23353 ( .A1(n20701), .A2(n20433), .B1(n20700), .B2(n20434), .ZN(
        n20426) );
  AOI22_X1 U23354 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20436), .B1(
        n20435), .B2(n20702), .ZN(n20425) );
  OAI211_X1 U23355 ( .C1(n9829), .C2(n20465), .A(n20426), .B(n20425), .ZN(
        P1_U3068) );
  AOI22_X1 U23356 ( .A1(n20707), .A2(n20433), .B1(n20706), .B2(n20434), .ZN(
        n20428) );
  AOI22_X1 U23357 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20436), .B1(
        n20435), .B2(n20708), .ZN(n20427) );
  OAI211_X1 U23358 ( .C1(n20711), .C2(n20465), .A(n20428), .B(n20427), .ZN(
        P1_U3069) );
  AOI22_X1 U23359 ( .A1(n20713), .A2(n20433), .B1(n20712), .B2(n20434), .ZN(
        n20430) );
  AOI22_X1 U23360 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20436), .B1(
        n20435), .B2(n20714), .ZN(n20429) );
  OAI211_X1 U23361 ( .C1(n9831), .C2(n20465), .A(n20430), .B(n20429), .ZN(
        P1_U3070) );
  AOI22_X1 U23362 ( .A1(n20719), .A2(n20434), .B1(n20718), .B2(n20433), .ZN(
        n20432) );
  AOI22_X1 U23363 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20436), .B1(
        n20435), .B2(n20720), .ZN(n20431) );
  OAI211_X1 U23364 ( .C1(n20723), .C2(n20465), .A(n20432), .B(n20431), .ZN(
        P1_U3071) );
  AOI22_X1 U23365 ( .A1(n20727), .A2(n20434), .B1(n20725), .B2(n20433), .ZN(
        n20438) );
  AOI22_X1 U23366 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20436), .B1(
        n20435), .B2(n20728), .ZN(n20437) );
  OAI211_X1 U23367 ( .C1(n20733), .C2(n20465), .A(n20438), .B(n20437), .ZN(
        P1_U3072) );
  INV_X1 U23368 ( .A(n20688), .ZN(n20500) );
  NOR2_X1 U23369 ( .A1(n20643), .A2(n20440), .ZN(n20459) );
  AOI21_X1 U23370 ( .B1(n20439), .B2(n20645), .A(n20459), .ZN(n20441) );
  OAI22_X1 U23371 ( .A1(n20441), .A2(n20678), .B1(n20440), .B2(n20753), .ZN(
        n20460) );
  AOI22_X1 U23372 ( .A1(n20680), .A2(n20459), .B1(n20679), .B2(n20460), .ZN(
        n20446) );
  INV_X1 U23373 ( .A(n20440), .ZN(n20444) );
  OAI21_X1 U23374 ( .B1(n20442), .B2(n20841), .A(n20441), .ZN(n20443) );
  OAI221_X1 U23375 ( .B1(n20596), .B2(n20444), .C1(n20678), .C2(n20443), .A(
        n20650), .ZN(n20462) );
  AOI22_X1 U23376 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20462), .B1(
        n20461), .B2(n20603), .ZN(n20445) );
  OAI211_X1 U23377 ( .C1(n20500), .C2(n20465), .A(n20446), .B(n20445), .ZN(
        P1_U3073) );
  INV_X1 U23378 ( .A(n20692), .ZN(n20739) );
  AOI22_X1 U23379 ( .A1(n20735), .A2(n20459), .B1(n20734), .B2(n20460), .ZN(
        n20448) );
  AOI22_X1 U23380 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20462), .B1(
        n20461), .B2(n20736), .ZN(n20447) );
  OAI211_X1 U23381 ( .C1(n20739), .C2(n20465), .A(n20448), .B(n20447), .ZN(
        P1_U3074) );
  INV_X1 U23382 ( .A(n20696), .ZN(n20750) );
  AOI22_X1 U23383 ( .A1(n20743), .A2(n20459), .B1(n20741), .B2(n20460), .ZN(
        n20450) );
  AOI22_X1 U23384 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20462), .B1(
        n20461), .B2(n20744), .ZN(n20449) );
  OAI211_X1 U23385 ( .C1(n20750), .C2(n20465), .A(n20450), .B(n20449), .ZN(
        P1_U3075) );
  INV_X1 U23386 ( .A(n20702), .ZN(n20507) );
  AOI22_X1 U23387 ( .A1(n20701), .A2(n20459), .B1(n20700), .B2(n20460), .ZN(
        n20452) );
  AOI22_X1 U23388 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20462), .B1(
        n20461), .B2(n9828), .ZN(n20451) );
  OAI211_X1 U23389 ( .C1(n20507), .C2(n20465), .A(n20452), .B(n20451), .ZN(
        P1_U3076) );
  AOI22_X1 U23390 ( .A1(n20707), .A2(n20459), .B1(n20706), .B2(n20460), .ZN(
        n20454) );
  AOI22_X1 U23391 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20462), .B1(
        n20461), .B2(n20623), .ZN(n20453) );
  OAI211_X1 U23392 ( .C1(n20510), .C2(n20465), .A(n20454), .B(n20453), .ZN(
        P1_U3077) );
  INV_X1 U23393 ( .A(n20714), .ZN(n20513) );
  AOI22_X1 U23394 ( .A1(n20713), .A2(n20459), .B1(n20712), .B2(n20460), .ZN(
        n20456) );
  AOI22_X1 U23395 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20462), .B1(
        n20461), .B2(n9830), .ZN(n20455) );
  OAI211_X1 U23396 ( .C1(n20513), .C2(n20465), .A(n20456), .B(n20455), .ZN(
        P1_U3078) );
  AOI22_X1 U23397 ( .A1(n20719), .A2(n20460), .B1(n20718), .B2(n20459), .ZN(
        n20458) );
  AOI22_X1 U23398 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20462), .B1(
        n20461), .B2(n20630), .ZN(n20457) );
  OAI211_X1 U23399 ( .C1(n20516), .C2(n20465), .A(n20458), .B(n20457), .ZN(
        P1_U3079) );
  INV_X1 U23400 ( .A(n20728), .ZN(n20523) );
  AOI22_X1 U23401 ( .A1(n20727), .A2(n20460), .B1(n20725), .B2(n20459), .ZN(
        n20464) );
  AOI22_X1 U23402 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20462), .B1(
        n20461), .B2(n20635), .ZN(n20463) );
  OAI211_X1 U23403 ( .C1(n20523), .C2(n20465), .A(n20464), .B(n20463), .ZN(
        P1_U3080) );
  NAND3_X1 U23404 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20532), .A3(
        n20602), .ZN(n20494) );
  NOR2_X1 U23405 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20494), .ZN(
        n20488) );
  AND2_X1 U23406 ( .A1(n20467), .A2(n13068), .ZN(n20561) );
  AOI21_X1 U23407 ( .B1(n20561), .B2(n13652), .A(n20488), .ZN(n20471) );
  AND2_X1 U23408 ( .A1(n20468), .A2(n20529), .ZN(n20600) );
  INV_X1 U23409 ( .A(n20600), .ZN(n20605) );
  OAI22_X1 U23410 ( .A1(n20471), .A2(n20678), .B1(n20605), .B2(n20469), .ZN(
        n20489) );
  AOI22_X1 U23411 ( .A1(n20680), .A2(n20488), .B1(n20679), .B2(n20489), .ZN(
        n20475) );
  INV_X1 U23412 ( .A(n20522), .ZN(n20470) );
  OAI21_X1 U23413 ( .B1(n20470), .B2(n20490), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20472) );
  NAND2_X1 U23414 ( .A1(n20472), .A2(n20471), .ZN(n20473) );
  AOI22_X1 U23415 ( .A1(n20491), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n20688), .B2(n20490), .ZN(n20474) );
  OAI211_X1 U23416 ( .C1(n20691), .C2(n20522), .A(n20475), .B(n20474), .ZN(
        P1_U3097) );
  AOI22_X1 U23417 ( .A1(n20735), .A2(n20488), .B1(n20734), .B2(n20489), .ZN(
        n20477) );
  AOI22_X1 U23418 ( .A1(n20491), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n20692), .B2(n20490), .ZN(n20476) );
  OAI211_X1 U23419 ( .C1(n20695), .C2(n20522), .A(n20477), .B(n20476), .ZN(
        P1_U3098) );
  AOI22_X1 U23420 ( .A1(n20743), .A2(n20488), .B1(n20741), .B2(n20489), .ZN(
        n20479) );
  AOI22_X1 U23421 ( .A1(n20491), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n20696), .B2(n20490), .ZN(n20478) );
  OAI211_X1 U23422 ( .C1(n20699), .C2(n20522), .A(n20479), .B(n20478), .ZN(
        P1_U3099) );
  AOI22_X1 U23423 ( .A1(n20701), .A2(n20488), .B1(n20700), .B2(n20489), .ZN(
        n20481) );
  AOI22_X1 U23424 ( .A1(n20491), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n20702), .B2(n20490), .ZN(n20480) );
  OAI211_X1 U23425 ( .C1(n9829), .C2(n20522), .A(n20481), .B(n20480), .ZN(
        P1_U3100) );
  AOI22_X1 U23426 ( .A1(n20707), .A2(n20488), .B1(n20706), .B2(n20489), .ZN(
        n20483) );
  AOI22_X1 U23427 ( .A1(n20491), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n20708), .B2(n20490), .ZN(n20482) );
  OAI211_X1 U23428 ( .C1(n20711), .C2(n20522), .A(n20483), .B(n20482), .ZN(
        P1_U3101) );
  AOI22_X1 U23429 ( .A1(n20713), .A2(n20488), .B1(n20712), .B2(n20489), .ZN(
        n20485) );
  AOI22_X1 U23430 ( .A1(n20491), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n20714), .B2(n20490), .ZN(n20484) );
  OAI211_X1 U23431 ( .C1(n9831), .C2(n20522), .A(n20485), .B(n20484), .ZN(
        P1_U3102) );
  AOI22_X1 U23432 ( .A1(n20719), .A2(n20489), .B1(n20718), .B2(n20488), .ZN(
        n20487) );
  AOI22_X1 U23433 ( .A1(n20491), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n20720), .B2(n20490), .ZN(n20486) );
  OAI211_X1 U23434 ( .C1(n20723), .C2(n20522), .A(n20487), .B(n20486), .ZN(
        P1_U3103) );
  AOI22_X1 U23435 ( .A1(n20727), .A2(n20489), .B1(n20725), .B2(n20488), .ZN(
        n20493) );
  AOI22_X1 U23436 ( .A1(n20491), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n20728), .B2(n20490), .ZN(n20492) );
  OAI211_X1 U23437 ( .C1(n20733), .C2(n20522), .A(n20493), .B(n20492), .ZN(
        P1_U3104) );
  NOR2_X1 U23438 ( .A1(n20643), .A2(n20494), .ZN(n20517) );
  AOI21_X1 U23439 ( .B1(n20561), .B2(n20645), .A(n20517), .ZN(n20495) );
  OAI22_X1 U23440 ( .A1(n20495), .A2(n20678), .B1(n20494), .B2(n20753), .ZN(
        n20518) );
  AOI22_X1 U23441 ( .A1(n20680), .A2(n20517), .B1(n20679), .B2(n20518), .ZN(
        n20499) );
  INV_X1 U23442 ( .A(n20494), .ZN(n20497) );
  OAI211_X1 U23443 ( .C1(n20569), .C2(n20841), .A(n20596), .B(n20495), .ZN(
        n20496) );
  OAI211_X1 U23444 ( .C1(n20596), .C2(n20497), .A(n20650), .B(n20496), .ZN(
        n20519) );
  AOI22_X1 U23445 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20519), .B1(
        n20554), .B2(n20603), .ZN(n20498) );
  OAI211_X1 U23446 ( .C1(n20500), .C2(n20522), .A(n20499), .B(n20498), .ZN(
        P1_U3105) );
  AOI22_X1 U23447 ( .A1(n20735), .A2(n20517), .B1(n20734), .B2(n20518), .ZN(
        n20502) );
  AOI22_X1 U23448 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20519), .B1(
        n20554), .B2(n20736), .ZN(n20501) );
  OAI211_X1 U23449 ( .C1(n20739), .C2(n20522), .A(n20502), .B(n20501), .ZN(
        P1_U3106) );
  AOI22_X1 U23450 ( .A1(n20743), .A2(n20517), .B1(n20741), .B2(n20518), .ZN(
        n20504) );
  AOI22_X1 U23451 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20519), .B1(
        n20554), .B2(n20744), .ZN(n20503) );
  OAI211_X1 U23452 ( .C1(n20750), .C2(n20522), .A(n20504), .B(n20503), .ZN(
        P1_U3107) );
  AOI22_X1 U23453 ( .A1(n20701), .A2(n20517), .B1(n20700), .B2(n20518), .ZN(
        n20506) );
  AOI22_X1 U23454 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20519), .B1(
        n20554), .B2(n9828), .ZN(n20505) );
  OAI211_X1 U23455 ( .C1(n20507), .C2(n20522), .A(n20506), .B(n20505), .ZN(
        P1_U3108) );
  AOI22_X1 U23456 ( .A1(n20707), .A2(n20517), .B1(n20706), .B2(n20518), .ZN(
        n20509) );
  AOI22_X1 U23457 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20519), .B1(
        n20554), .B2(n20623), .ZN(n20508) );
  OAI211_X1 U23458 ( .C1(n20510), .C2(n20522), .A(n20509), .B(n20508), .ZN(
        P1_U3109) );
  AOI22_X1 U23459 ( .A1(n20713), .A2(n20517), .B1(n20712), .B2(n20518), .ZN(
        n20512) );
  AOI22_X1 U23460 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20519), .B1(
        n20554), .B2(n9830), .ZN(n20511) );
  OAI211_X1 U23461 ( .C1(n20513), .C2(n20522), .A(n20512), .B(n20511), .ZN(
        P1_U3110) );
  AOI22_X1 U23462 ( .A1(n20719), .A2(n20518), .B1(n20718), .B2(n20517), .ZN(
        n20515) );
  AOI22_X1 U23463 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20519), .B1(
        n20554), .B2(n20630), .ZN(n20514) );
  OAI211_X1 U23464 ( .C1(n20516), .C2(n20522), .A(n20515), .B(n20514), .ZN(
        P1_U3111) );
  AOI22_X1 U23465 ( .A1(n20727), .A2(n20518), .B1(n20725), .B2(n20517), .ZN(
        n20521) );
  AOI22_X1 U23466 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20519), .B1(
        n20554), .B2(n20635), .ZN(n20520) );
  OAI211_X1 U23467 ( .C1(n20523), .C2(n20522), .A(n20521), .B(n20520), .ZN(
        P1_U3112) );
  INV_X1 U23468 ( .A(n20554), .ZN(n20524) );
  NAND2_X1 U23469 ( .A1(n20524), .A2(n20596), .ZN(n20527) );
  INV_X1 U23470 ( .A(n20526), .ZN(n20598) );
  OAI21_X1 U23471 ( .B1(n20527), .B2(n20591), .A(n20598), .ZN(n20533) );
  AND2_X1 U23472 ( .A1(n20561), .A2(n20674), .ZN(n20537) );
  OR2_X1 U23473 ( .A1(n20529), .A2(n20528), .ZN(n20677) );
  INV_X1 U23474 ( .A(n20677), .ZN(n20531) );
  NAND3_X1 U23475 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n20532), .ZN(n20571) );
  NOR2_X1 U23476 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20571), .ZN(
        n20553) );
  AOI22_X1 U23477 ( .A1(n20591), .A2(n20603), .B1(n20553), .B2(n20680), .ZN(
        n20540) );
  INV_X1 U23478 ( .A(n20533), .ZN(n20538) );
  NAND2_X1 U23479 ( .A1(n20677), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20685) );
  OAI21_X1 U23480 ( .B1(n20609), .B2(n20553), .A(n20685), .ZN(n20534) );
  INV_X1 U23481 ( .A(n20534), .ZN(n20535) );
  AOI22_X1 U23482 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20555), .B1(
        n20554), .B2(n20688), .ZN(n20539) );
  OAI211_X1 U23483 ( .C1(n20558), .C2(n20613), .A(n20540), .B(n20539), .ZN(
        P1_U3113) );
  AOI22_X1 U23484 ( .A1(n20554), .A2(n20692), .B1(n20735), .B2(n20553), .ZN(
        n20542) );
  AOI22_X1 U23485 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20555), .B1(
        n20591), .B2(n20736), .ZN(n20541) );
  OAI211_X1 U23486 ( .C1(n20558), .C2(n20616), .A(n20542), .B(n20541), .ZN(
        P1_U3114) );
  AOI22_X1 U23487 ( .A1(n20554), .A2(n20696), .B1(n20743), .B2(n20553), .ZN(
        n20544) );
  AOI22_X1 U23488 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20555), .B1(
        n20591), .B2(n20744), .ZN(n20543) );
  OAI211_X1 U23489 ( .C1(n20558), .C2(n20619), .A(n20544), .B(n20543), .ZN(
        P1_U3115) );
  AOI22_X1 U23490 ( .A1(n20591), .A2(n9828), .B1(n20553), .B2(n20701), .ZN(
        n20546) );
  AOI22_X1 U23491 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20555), .B1(
        n20554), .B2(n20702), .ZN(n20545) );
  OAI211_X1 U23492 ( .C1(n20558), .C2(n20622), .A(n20546), .B(n20545), .ZN(
        P1_U3116) );
  AOI22_X1 U23493 ( .A1(n20591), .A2(n20623), .B1(n20553), .B2(n20707), .ZN(
        n20548) );
  AOI22_X1 U23494 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20555), .B1(
        n20554), .B2(n20708), .ZN(n20547) );
  OAI211_X1 U23495 ( .C1(n20558), .C2(n20626), .A(n20548), .B(n20547), .ZN(
        P1_U3117) );
  AOI22_X1 U23496 ( .A1(n20554), .A2(n20714), .B1(n20713), .B2(n20553), .ZN(
        n20550) );
  AOI22_X1 U23497 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20555), .B1(
        n20591), .B2(n9830), .ZN(n20549) );
  OAI211_X1 U23498 ( .C1(n20558), .C2(n20629), .A(n20550), .B(n20549), .ZN(
        P1_U3118) );
  AOI22_X1 U23499 ( .A1(n20554), .A2(n20720), .B1(n20718), .B2(n20553), .ZN(
        n20552) );
  AOI22_X1 U23500 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20555), .B1(
        n20591), .B2(n20630), .ZN(n20551) );
  OAI211_X1 U23501 ( .C1(n20558), .C2(n20633), .A(n20552), .B(n20551), .ZN(
        P1_U3119) );
  AOI22_X1 U23502 ( .A1(n20591), .A2(n20635), .B1(n20553), .B2(n20725), .ZN(
        n20557) );
  AOI22_X1 U23503 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20555), .B1(
        n20554), .B2(n20728), .ZN(n20556) );
  OAI211_X1 U23504 ( .C1(n20558), .C2(n20640), .A(n20557), .B(n20556), .ZN(
        P1_U3120) );
  INV_X1 U23505 ( .A(n20561), .ZN(n20565) );
  INV_X1 U23506 ( .A(n20562), .ZN(n20563) );
  NAND2_X1 U23507 ( .A1(n20563), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20567) );
  OAI21_X1 U23508 ( .B1(n20565), .B2(n20564), .A(n20567), .ZN(n20573) );
  INV_X1 U23509 ( .A(n20573), .ZN(n20566) );
  OAI22_X1 U23510 ( .A1(n20566), .A2(n20678), .B1(n20571), .B2(n20753), .ZN(
        n20590) );
  INV_X1 U23511 ( .A(n20567), .ZN(n20589) );
  AOI22_X1 U23512 ( .A1(n20590), .A2(n20679), .B1(n20680), .B2(n20589), .ZN(
        n20576) );
  AOI21_X1 U23513 ( .B1(n20569), .B2(n20596), .A(n20568), .ZN(n20574) );
  INV_X1 U23514 ( .A(n20650), .ZN(n20570) );
  AOI21_X1 U23515 ( .B1(n20678), .B2(n20571), .A(n20570), .ZN(n20572) );
  AOI22_X1 U23516 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20592), .B1(
        n20591), .B2(n20688), .ZN(n20575) );
  OAI211_X1 U23517 ( .C1(n20691), .C2(n20610), .A(n20576), .B(n20575), .ZN(
        P1_U3121) );
  AOI22_X1 U23518 ( .A1(n20590), .A2(n20734), .B1(n20735), .B2(n20589), .ZN(
        n20578) );
  AOI22_X1 U23519 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20592), .B1(
        n20591), .B2(n20692), .ZN(n20577) );
  OAI211_X1 U23520 ( .C1(n20695), .C2(n20610), .A(n20578), .B(n20577), .ZN(
        P1_U3122) );
  AOI22_X1 U23521 ( .A1(n20590), .A2(n20741), .B1(n20743), .B2(n20589), .ZN(
        n20580) );
  AOI22_X1 U23522 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20592), .B1(
        n20591), .B2(n20696), .ZN(n20579) );
  OAI211_X1 U23523 ( .C1(n20699), .C2(n20610), .A(n20580), .B(n20579), .ZN(
        P1_U3123) );
  AOI22_X1 U23524 ( .A1(n20590), .A2(n20700), .B1(n20701), .B2(n20589), .ZN(
        n20582) );
  AOI22_X1 U23525 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20592), .B1(
        n20591), .B2(n20702), .ZN(n20581) );
  OAI211_X1 U23526 ( .C1(n9829), .C2(n20610), .A(n20582), .B(n20581), .ZN(
        P1_U3124) );
  AOI22_X1 U23527 ( .A1(n20590), .A2(n20706), .B1(n20707), .B2(n20589), .ZN(
        n20584) );
  AOI22_X1 U23528 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20592), .B1(
        n20591), .B2(n20708), .ZN(n20583) );
  OAI211_X1 U23529 ( .C1(n20711), .C2(n20610), .A(n20584), .B(n20583), .ZN(
        P1_U3125) );
  AOI22_X1 U23530 ( .A1(n20590), .A2(n20712), .B1(n20713), .B2(n20589), .ZN(
        n20586) );
  AOI22_X1 U23531 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20592), .B1(
        n20591), .B2(n20714), .ZN(n20585) );
  OAI211_X1 U23532 ( .C1(n9831), .C2(n20610), .A(n20586), .B(n20585), .ZN(
        P1_U3126) );
  AOI22_X1 U23533 ( .A1(n20590), .A2(n20719), .B1(n20718), .B2(n20589), .ZN(
        n20588) );
  AOI22_X1 U23534 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20592), .B1(
        n20591), .B2(n20720), .ZN(n20587) );
  OAI211_X1 U23535 ( .C1(n20723), .C2(n20610), .A(n20588), .B(n20587), .ZN(
        P1_U3127) );
  AOI22_X1 U23536 ( .A1(n20590), .A2(n20727), .B1(n20725), .B2(n20589), .ZN(
        n20594) );
  AOI22_X1 U23537 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20592), .B1(
        n20591), .B2(n20728), .ZN(n20593) );
  OAI211_X1 U23538 ( .C1(n20733), .C2(n20610), .A(n20594), .B(n20593), .ZN(
        P1_U3128) );
  INV_X1 U23539 ( .A(n20669), .ZN(n20597) );
  NAND3_X1 U23540 ( .A1(n20597), .A2(n20596), .A3(n20610), .ZN(n20599) );
  NAND2_X1 U23541 ( .A1(n20599), .A2(n20598), .ZN(n20607) );
  NOR2_X1 U23542 ( .A1(n20644), .A2(n20674), .ZN(n20604) );
  NAND3_X1 U23543 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20602), .ZN(n20649) );
  NOR2_X1 U23544 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20649), .ZN(
        n20634) );
  AOI22_X1 U23545 ( .A1(n20669), .A2(n20603), .B1(n20634), .B2(n20680), .ZN(
        n20612) );
  INV_X1 U23546 ( .A(n20604), .ZN(n20606) );
  AOI22_X1 U23547 ( .A1(n20607), .A2(n20606), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20605), .ZN(n20608) );
  OAI211_X1 U23548 ( .C1(n20634), .C2(n20609), .A(n20686), .B(n20608), .ZN(
        n20637) );
  AOI22_X1 U23549 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20637), .B1(
        n20636), .B2(n20688), .ZN(n20611) );
  OAI211_X1 U23550 ( .C1(n20641), .C2(n20613), .A(n20612), .B(n20611), .ZN(
        P1_U3129) );
  AOI22_X1 U23551 ( .A1(n20669), .A2(n20736), .B1(n20634), .B2(n20735), .ZN(
        n20615) );
  AOI22_X1 U23552 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20637), .B1(
        n20636), .B2(n20692), .ZN(n20614) );
  OAI211_X1 U23553 ( .C1(n20641), .C2(n20616), .A(n20615), .B(n20614), .ZN(
        P1_U3130) );
  AOI22_X1 U23554 ( .A1(n20669), .A2(n20744), .B1(n20634), .B2(n20743), .ZN(
        n20618) );
  AOI22_X1 U23555 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20637), .B1(
        n20636), .B2(n20696), .ZN(n20617) );
  OAI211_X1 U23556 ( .C1(n20641), .C2(n20619), .A(n20618), .B(n20617), .ZN(
        P1_U3131) );
  AOI22_X1 U23557 ( .A1(n20669), .A2(n9828), .B1(n20634), .B2(n20701), .ZN(
        n20621) );
  AOI22_X1 U23558 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20637), .B1(
        n20636), .B2(n20702), .ZN(n20620) );
  OAI211_X1 U23559 ( .C1(n20641), .C2(n20622), .A(n20621), .B(n20620), .ZN(
        P1_U3132) );
  AOI22_X1 U23560 ( .A1(n20669), .A2(n20623), .B1(n20634), .B2(n20707), .ZN(
        n20625) );
  AOI22_X1 U23561 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20637), .B1(
        n20636), .B2(n20708), .ZN(n20624) );
  OAI211_X1 U23562 ( .C1(n20641), .C2(n20626), .A(n20625), .B(n20624), .ZN(
        P1_U3133) );
  AOI22_X1 U23563 ( .A1(n20669), .A2(n9830), .B1(n20634), .B2(n20713), .ZN(
        n20628) );
  AOI22_X1 U23564 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20637), .B1(
        n20636), .B2(n20714), .ZN(n20627) );
  OAI211_X1 U23565 ( .C1(n20641), .C2(n20629), .A(n20628), .B(n20627), .ZN(
        P1_U3134) );
  AOI22_X1 U23566 ( .A1(n20669), .A2(n20630), .B1(n20634), .B2(n20718), .ZN(
        n20632) );
  AOI22_X1 U23567 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20637), .B1(
        n20636), .B2(n20720), .ZN(n20631) );
  OAI211_X1 U23568 ( .C1(n20641), .C2(n20633), .A(n20632), .B(n20631), .ZN(
        P1_U3135) );
  AOI22_X1 U23569 ( .A1(n20669), .A2(n20635), .B1(n20634), .B2(n20725), .ZN(
        n20639) );
  AOI22_X1 U23570 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20637), .B1(
        n20636), .B2(n20728), .ZN(n20638) );
  OAI211_X1 U23571 ( .C1(n20641), .C2(n20640), .A(n20639), .B(n20638), .ZN(
        P1_U3136) );
  NOR2_X1 U23572 ( .A1(n20643), .A2(n20649), .ZN(n20667) );
  INV_X1 U23573 ( .A(n20644), .ZN(n20675) );
  AOI21_X1 U23574 ( .B1(n20675), .B2(n20645), .A(n20667), .ZN(n20646) );
  OAI22_X1 U23575 ( .A1(n20646), .A2(n20678), .B1(n20649), .B2(n20753), .ZN(
        n20668) );
  AOI22_X1 U23576 ( .A1(n20680), .A2(n20667), .B1(n20679), .B2(n20668), .ZN(
        n20654) );
  NOR2_X1 U23577 ( .A1(n20648), .A2(n20647), .ZN(n20652) );
  INV_X1 U23578 ( .A(n20649), .ZN(n20651) );
  OAI21_X1 U23579 ( .B1(n20652), .B2(n20651), .A(n20650), .ZN(n20670) );
  AOI22_X1 U23580 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20670), .B1(
        n20669), .B2(n20688), .ZN(n20653) );
  OAI211_X1 U23581 ( .C1(n20691), .C2(n20681), .A(n20654), .B(n20653), .ZN(
        P1_U3137) );
  AOI22_X1 U23582 ( .A1(n20735), .A2(n20667), .B1(n20734), .B2(n20668), .ZN(
        n20656) );
  AOI22_X1 U23583 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20670), .B1(
        n20669), .B2(n20692), .ZN(n20655) );
  OAI211_X1 U23584 ( .C1(n20695), .C2(n20681), .A(n20656), .B(n20655), .ZN(
        P1_U3138) );
  AOI22_X1 U23585 ( .A1(n20743), .A2(n20667), .B1(n20741), .B2(n20668), .ZN(
        n20658) );
  AOI22_X1 U23586 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20670), .B1(
        n20669), .B2(n20696), .ZN(n20657) );
  OAI211_X1 U23587 ( .C1(n20699), .C2(n20681), .A(n20658), .B(n20657), .ZN(
        P1_U3139) );
  AOI22_X1 U23588 ( .A1(n20701), .A2(n20667), .B1(n20700), .B2(n20668), .ZN(
        n20660) );
  AOI22_X1 U23589 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20670), .B1(
        n20669), .B2(n20702), .ZN(n20659) );
  OAI211_X1 U23590 ( .C1(n9829), .C2(n20681), .A(n20660), .B(n20659), .ZN(
        P1_U3140) );
  AOI22_X1 U23591 ( .A1(n20707), .A2(n20667), .B1(n20706), .B2(n20668), .ZN(
        n20662) );
  AOI22_X1 U23592 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20670), .B1(
        n20669), .B2(n20708), .ZN(n20661) );
  OAI211_X1 U23593 ( .C1(n20711), .C2(n20681), .A(n20662), .B(n20661), .ZN(
        P1_U3141) );
  AOI22_X1 U23594 ( .A1(n20713), .A2(n20667), .B1(n20712), .B2(n20668), .ZN(
        n20664) );
  AOI22_X1 U23595 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20670), .B1(
        n20669), .B2(n20714), .ZN(n20663) );
  OAI211_X1 U23596 ( .C1(n9831), .C2(n20681), .A(n20664), .B(n20663), .ZN(
        P1_U3142) );
  AOI22_X1 U23597 ( .A1(n20719), .A2(n20668), .B1(n20718), .B2(n20667), .ZN(
        n20666) );
  AOI22_X1 U23598 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20670), .B1(
        n20669), .B2(n20720), .ZN(n20665) );
  OAI211_X1 U23599 ( .C1(n20723), .C2(n20681), .A(n20666), .B(n20665), .ZN(
        P1_U3143) );
  AOI22_X1 U23600 ( .A1(n20727), .A2(n20668), .B1(n20725), .B2(n20667), .ZN(
        n20672) );
  AOI22_X1 U23601 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20670), .B1(
        n20669), .B2(n20728), .ZN(n20671) );
  OAI211_X1 U23602 ( .C1(n20733), .C2(n20681), .A(n20672), .B(n20671), .ZN(
        P1_U3144) );
  NOR2_X1 U23603 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20673), .ZN(
        n20724) );
  NAND2_X1 U23604 ( .A1(n20675), .A2(n20674), .ZN(n20683) );
  OAI22_X1 U23605 ( .A1(n20683), .A2(n20678), .B1(n20677), .B2(n20676), .ZN(
        n20726) );
  AOI22_X1 U23606 ( .A1(n20680), .A2(n20724), .B1(n20679), .B2(n20726), .ZN(
        n20690) );
  OAI21_X1 U23607 ( .B1(n20682), .B2(n20729), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20684) );
  AOI21_X1 U23608 ( .B1(n20684), .B2(n20683), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20687) );
  AOI22_X1 U23609 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20730), .B1(
        n20729), .B2(n20688), .ZN(n20689) );
  OAI211_X1 U23610 ( .C1(n20691), .C2(n20749), .A(n20690), .B(n20689), .ZN(
        P1_U3145) );
  AOI22_X1 U23611 ( .A1(n20735), .A2(n20724), .B1(n20734), .B2(n20726), .ZN(
        n20694) );
  AOI22_X1 U23612 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20730), .B1(
        n20729), .B2(n20692), .ZN(n20693) );
  OAI211_X1 U23613 ( .C1(n20695), .C2(n20749), .A(n20694), .B(n20693), .ZN(
        P1_U3146) );
  AOI22_X1 U23614 ( .A1(n20743), .A2(n20724), .B1(n20741), .B2(n20726), .ZN(
        n20698) );
  AOI22_X1 U23615 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20730), .B1(
        n20729), .B2(n20696), .ZN(n20697) );
  OAI211_X1 U23616 ( .C1(n20699), .C2(n20749), .A(n20698), .B(n20697), .ZN(
        P1_U3147) );
  AOI22_X1 U23617 ( .A1(n20701), .A2(n20724), .B1(n20700), .B2(n20726), .ZN(
        n20704) );
  AOI22_X1 U23618 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20730), .B1(
        n20729), .B2(n20702), .ZN(n20703) );
  OAI211_X1 U23619 ( .C1(n9829), .C2(n20749), .A(n20704), .B(n20703), .ZN(
        P1_U3148) );
  AOI22_X1 U23620 ( .A1(n20707), .A2(n20724), .B1(n20706), .B2(n20726), .ZN(
        n20710) );
  AOI22_X1 U23621 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20730), .B1(
        n20729), .B2(n20708), .ZN(n20709) );
  OAI211_X1 U23622 ( .C1(n20711), .C2(n20749), .A(n20710), .B(n20709), .ZN(
        P1_U3149) );
  AOI22_X1 U23623 ( .A1(n20713), .A2(n20724), .B1(n20712), .B2(n20726), .ZN(
        n20716) );
  AOI22_X1 U23624 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20730), .B1(
        n20729), .B2(n20714), .ZN(n20715) );
  OAI211_X1 U23625 ( .C1(n9831), .C2(n20749), .A(n20716), .B(n20715), .ZN(
        P1_U3150) );
  AOI22_X1 U23626 ( .A1(n20719), .A2(n20726), .B1(n20718), .B2(n20724), .ZN(
        n20722) );
  AOI22_X1 U23627 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20730), .B1(
        n20729), .B2(n20720), .ZN(n20721) );
  OAI211_X1 U23628 ( .C1(n20723), .C2(n20749), .A(n20722), .B(n20721), .ZN(
        P1_U3151) );
  AOI22_X1 U23629 ( .A1(n20727), .A2(n20726), .B1(n20725), .B2(n20724), .ZN(
        n20732) );
  AOI22_X1 U23630 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20730), .B1(
        n20729), .B2(n20728), .ZN(n20731) );
  OAI211_X1 U23631 ( .C1(n20733), .C2(n20749), .A(n20732), .B(n20731), .ZN(
        P1_U3152) );
  AOI22_X1 U23632 ( .A1(n20735), .A2(n20742), .B1(n20734), .B2(n20740), .ZN(
        n20738) );
  AOI22_X1 U23633 ( .A1(n20746), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n20745), .B2(n20736), .ZN(n20737) );
  OAI211_X1 U23634 ( .C1(n20739), .C2(n20749), .A(n20738), .B(n20737), .ZN(
        P1_U3154) );
  AOI22_X1 U23635 ( .A1(n20743), .A2(n20742), .B1(n20741), .B2(n20740), .ZN(
        n20748) );
  AOI22_X1 U23636 ( .A1(n20746), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n20745), .B2(n20744), .ZN(n20747) );
  OAI211_X1 U23637 ( .C1(n20750), .C2(n20749), .A(n20748), .B(n20747), .ZN(
        P1_U3155) );
  OAI221_X1 U23638 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20754), .C1(n20753), 
        .C2(n20752), .A(n20751), .ZN(P1_U3163) );
  AND2_X1 U23639 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20827), .ZN(
        P1_U3164) );
  AND2_X1 U23640 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20827), .ZN(
        P1_U3165) );
  AND2_X1 U23641 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20827), .ZN(
        P1_U3166) );
  AND2_X1 U23642 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20827), .ZN(
        P1_U3167) );
  AND2_X1 U23643 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20827), .ZN(
        P1_U3168) );
  AND2_X1 U23644 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20827), .ZN(
        P1_U3169) );
  AND2_X1 U23645 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20827), .ZN(
        P1_U3170) );
  AND2_X1 U23646 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20827), .ZN(
        P1_U3171) );
  AND2_X1 U23647 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20827), .ZN(
        P1_U3172) );
  AND2_X1 U23648 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20827), .ZN(
        P1_U3173) );
  AND2_X1 U23649 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20827), .ZN(
        P1_U3174) );
  AND2_X1 U23650 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20827), .ZN(
        P1_U3175) );
  AND2_X1 U23651 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20827), .ZN(
        P1_U3176) );
  AND2_X1 U23652 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20827), .ZN(
        P1_U3177) );
  AND2_X1 U23653 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20827), .ZN(
        P1_U3178) );
  AND2_X1 U23654 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20827), .ZN(
        P1_U3179) );
  AND2_X1 U23655 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20827), .ZN(
        P1_U3180) );
  AND2_X1 U23656 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20827), .ZN(
        P1_U3181) );
  AND2_X1 U23657 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20827), .ZN(
        P1_U3182) );
  AND2_X1 U23658 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20827), .ZN(
        P1_U3183) );
  AND2_X1 U23659 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20827), .ZN(
        P1_U3184) );
  AND2_X1 U23660 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20827), .ZN(
        P1_U3185) );
  AND2_X1 U23661 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20827), .ZN(P1_U3186) );
  AND2_X1 U23662 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20827), .ZN(P1_U3187) );
  AND2_X1 U23663 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20827), .ZN(P1_U3188) );
  AND2_X1 U23664 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20827), .ZN(P1_U3189) );
  AND2_X1 U23665 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20827), .ZN(P1_U3190) );
  AND2_X1 U23666 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20827), .ZN(P1_U3191) );
  AND2_X1 U23667 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20827), .ZN(P1_U3192) );
  AND2_X1 U23668 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20827), .ZN(P1_U3193) );
  OAI21_X1 U23669 ( .B1(n20755), .B2(n20850), .A(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20761) );
  INV_X1 U23670 ( .A(n20761), .ZN(n20759) );
  NOR2_X1 U23671 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20756) );
  OAI22_X1 U23672 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20762), .B1(n20756), 
        .B2(n21016), .ZN(n20757) );
  NOR2_X1 U23673 ( .A1(n21021), .A2(n20757), .ZN(n20758) );
  OAI22_X1 U23674 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20759), .B1(n20855), 
        .B2(n20758), .ZN(P1_U3194) );
  AOI21_X1 U23675 ( .B1(n20840), .B2(n20762), .A(n20760), .ZN(n20767) );
  OAI211_X1 U23676 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n21021), .A(
        P1_STATE_REG_0__SCAN_IN), .B(HOLD), .ZN(n20766) );
  OAI211_X1 U23677 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n20762), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n20761), .ZN(n20765) );
  NOR2_X1 U23678 ( .A1(NA), .A2(n20850), .ZN(n20763) );
  NAND4_X1 U23679 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .A3(P1_REQUESTPENDING_REG_SCAN_IN), .A4(n20763), .ZN(n20764) );
  OAI211_X1 U23680 ( .C1(n20767), .C2(n20766), .A(n20765), .B(n20764), .ZN(
        P1_U3196) );
  NAND2_X1 U23681 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20855), .ZN(n20810) );
  NOR2_X1 U23682 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20854), .ZN(n20791) );
  AOI22_X1 U23683 ( .A1(P1_ADDRESS_REG_0__SCAN_IN), .A2(n20854), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n20791), .ZN(n20768) );
  OAI21_X1 U23684 ( .B1(n20832), .B2(n20810), .A(n20768), .ZN(P1_U3197) );
  INV_X1 U23685 ( .A(n20810), .ZN(n20793) );
  AOI22_X1 U23686 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n20854), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n20793), .ZN(n20769) );
  OAI21_X1 U23687 ( .B1(n20771), .B2(n20816), .A(n20769), .ZN(P1_U3198) );
  INV_X1 U23688 ( .A(n20793), .ZN(n20819) );
  OAI222_X1 U23689 ( .A1(n20819), .A2(n20771), .B1(n20770), .B2(n20817), .C1(
        n20772), .C2(n20816), .ZN(P1_U3199) );
  INV_X1 U23690 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20773) );
  OAI222_X1 U23691 ( .A1(n20816), .A2(n20775), .B1(n20773), .B2(n20817), .C1(
        n20772), .C2(n20810), .ZN(P1_U3200) );
  INV_X1 U23692 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n20774) );
  OAI222_X1 U23693 ( .A1(n20810), .A2(n20775), .B1(n20774), .B2(n20817), .C1(
        n20777), .C2(n20816), .ZN(P1_U3201) );
  AOI22_X1 U23694 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n20854), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20791), .ZN(n20776) );
  OAI21_X1 U23695 ( .B1(n20777), .B2(n20810), .A(n20776), .ZN(P1_U3202) );
  INV_X1 U23696 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20779) );
  AOI22_X1 U23697 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n20854), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n20791), .ZN(n20778) );
  OAI21_X1 U23698 ( .B1(n20779), .B2(n20810), .A(n20778), .ZN(P1_U3203) );
  AOI22_X1 U23699 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(n20854), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n20793), .ZN(n20780) );
  OAI21_X1 U23700 ( .B1(n13889), .B2(n20816), .A(n20780), .ZN(P1_U3204) );
  INV_X1 U23701 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20781) );
  INV_X1 U23702 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20782) );
  OAI222_X1 U23703 ( .A1(n20819), .A2(n13889), .B1(n20781), .B2(n20817), .C1(
        n20782), .C2(n20816), .ZN(P1_U3205) );
  INV_X1 U23704 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20783) );
  OAI222_X1 U23705 ( .A1(n20816), .A2(n20785), .B1(n20783), .B2(n20817), .C1(
        n20782), .C2(n20810), .ZN(P1_U3206) );
  INV_X1 U23706 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n20784) );
  OAI222_X1 U23707 ( .A1(n20819), .A2(n20785), .B1(n20784), .B2(n20817), .C1(
        n20786), .C2(n20816), .ZN(P1_U3207) );
  INV_X1 U23708 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n20787) );
  OAI222_X1 U23709 ( .A1(n20816), .A2(n20789), .B1(n20787), .B2(n20855), .C1(
        n20786), .C2(n20810), .ZN(P1_U3208) );
  AOI22_X1 U23710 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n20854), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20791), .ZN(n20788) );
  OAI21_X1 U23711 ( .B1(n20789), .B2(n20810), .A(n20788), .ZN(P1_U3209) );
  AOI22_X1 U23712 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n20854), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20793), .ZN(n20790) );
  OAI21_X1 U23713 ( .B1(n14778), .B2(n20816), .A(n20790), .ZN(P1_U3210) );
  AOI22_X1 U23714 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(n20854), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n20791), .ZN(n20792) );
  OAI21_X1 U23715 ( .B1(n14778), .B2(n20810), .A(n20792), .ZN(P1_U3211) );
  AOI22_X1 U23716 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20854), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n20793), .ZN(n20794) );
  OAI21_X1 U23717 ( .B1(n20795), .B2(n20816), .A(n20794), .ZN(P1_U3212) );
  INV_X1 U23718 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n20796) );
  OAI222_X1 U23719 ( .A1(n20816), .A2(n20798), .B1(n20796), .B2(n20817), .C1(
        n20795), .C2(n20810), .ZN(P1_U3213) );
  INV_X1 U23720 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n20797) );
  OAI222_X1 U23721 ( .A1(n20819), .A2(n20798), .B1(n20797), .B2(n20817), .C1(
        n20800), .C2(n20816), .ZN(P1_U3214) );
  INV_X1 U23722 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n20799) );
  OAI222_X1 U23723 ( .A1(n20819), .A2(n20800), .B1(n20799), .B2(n20817), .C1(
        n20877), .C2(n20816), .ZN(P1_U3215) );
  INV_X1 U23724 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n20801) );
  OAI222_X1 U23725 ( .A1(n20816), .A2(n20802), .B1(n20801), .B2(n20855), .C1(
        n20877), .C2(n20810), .ZN(P1_U3216) );
  INV_X1 U23726 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20803) );
  OAI222_X1 U23727 ( .A1(n20816), .A2(n20859), .B1(n20803), .B2(n20855), .C1(
        n20802), .C2(n20819), .ZN(P1_U3217) );
  INV_X1 U23728 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n20804) );
  OAI222_X1 U23729 ( .A1(n20819), .A2(n20859), .B1(n20804), .B2(n20855), .C1(
        n20806), .C2(n20816), .ZN(P1_U3218) );
  INV_X1 U23730 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n20805) );
  OAI222_X1 U23731 ( .A1(n20819), .A2(n20806), .B1(n20805), .B2(n20855), .C1(
        n20873), .C2(n20816), .ZN(P1_U3219) );
  INV_X1 U23732 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20807) );
  OAI222_X1 U23733 ( .A1(n20816), .A2(n20809), .B1(n20807), .B2(n20855), .C1(
        n20873), .C2(n20810), .ZN(P1_U3220) );
  INV_X1 U23734 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20808) );
  OAI222_X1 U23735 ( .A1(n20819), .A2(n20809), .B1(n20808), .B2(n20855), .C1(
        n20811), .C2(n20816), .ZN(P1_U3221) );
  INV_X1 U23736 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20812) );
  OAI222_X1 U23737 ( .A1(n20816), .A2(n20887), .B1(n20812), .B2(n20855), .C1(
        n20811), .C2(n20810), .ZN(P1_U3222) );
  INV_X1 U23738 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n20813) );
  OAI222_X1 U23739 ( .A1(n20819), .A2(n20887), .B1(n20813), .B2(n20855), .C1(
        n21005), .C2(n20816), .ZN(P1_U3223) );
  INV_X1 U23740 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n20814) );
  OAI222_X1 U23741 ( .A1(n20819), .A2(n21005), .B1(n20814), .B2(n20855), .C1(
        n20917), .C2(n20816), .ZN(P1_U3224) );
  INV_X1 U23742 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n20815) );
  INV_X1 U23743 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n21006) );
  OAI222_X1 U23744 ( .A1(n20819), .A2(n20917), .B1(n20815), .B2(n20855), .C1(
        n21006), .C2(n20816), .ZN(P1_U3225) );
  INV_X1 U23745 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20818) );
  OAI222_X1 U23746 ( .A1(n20819), .A2(n21006), .B1(n20818), .B2(n20817), .C1(
        n21036), .C2(n20816), .ZN(P1_U3226) );
  INV_X1 U23747 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20820) );
  AOI22_X1 U23748 ( .A1(n20855), .A2(n20821), .B1(n20820), .B2(n20854), .ZN(
        P1_U3458) );
  INV_X1 U23749 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20884) );
  INV_X1 U23750 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20822) );
  AOI22_X1 U23751 ( .A1(n20855), .A2(n20884), .B1(n20822), .B2(n20854), .ZN(
        P1_U3459) );
  INV_X1 U23752 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20823) );
  AOI22_X1 U23753 ( .A1(n20855), .A2(n20824), .B1(n20823), .B2(n20854), .ZN(
        P1_U3460) );
  INV_X1 U23754 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20837) );
  INV_X1 U23755 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20825) );
  AOI22_X1 U23756 ( .A1(n20855), .A2(n20837), .B1(n20825), .B2(n20854), .ZN(
        P1_U3461) );
  INV_X1 U23757 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20828) );
  INV_X1 U23758 ( .A(n20829), .ZN(n20826) );
  AOI21_X1 U23759 ( .B1(n20828), .B2(n20827), .A(n20826), .ZN(P1_U3464) );
  OAI21_X1 U23760 ( .B1(n20831), .B2(n20830), .A(n20829), .ZN(P1_U3465) );
  AOI21_X1 U23761 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20833) );
  AOI22_X1 U23762 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20833), .B2(n20832), .ZN(n20835) );
  AOI22_X1 U23763 ( .A1(n20838), .A2(n20835), .B1(n20884), .B2(n20834), .ZN(
        P1_U3481) );
  OAI21_X1 U23764 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20838), .ZN(n20836) );
  OAI21_X1 U23765 ( .B1(n20838), .B2(n20837), .A(n20836), .ZN(P1_U3482) );
  INV_X1 U23766 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20839) );
  AOI22_X1 U23767 ( .A1(n20855), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20839), 
        .B2(n20854), .ZN(P1_U3483) );
  AOI211_X1 U23768 ( .C1(n20842), .C2(n20841), .A(n20753), .B(n20840), .ZN(
        n20844) );
  AND2_X1 U23769 ( .A1(n20844), .A2(n20843), .ZN(n20847) );
  OAI21_X1 U23770 ( .B1(n20847), .B2(n20846), .A(n20845), .ZN(n20853) );
  AOI211_X1 U23771 ( .C1(n20851), .C2(n20850), .A(n20849), .B(n20848), .ZN(
        n20852) );
  MUX2_X1 U23772 ( .A(n20853), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n20852), 
        .Z(P1_U3485) );
  AOI22_X1 U23773 ( .A1(n20855), .A2(n21033), .B1(n20992), .B2(n20854), .ZN(
        P1_U3486) );
  INV_X1 U23774 ( .A(DATAI_2_), .ZN(n20950) );
  INV_X1 U23775 ( .A(keyinput_f30), .ZN(n20949) );
  AOI22_X1 U23776 ( .A1(keyinput_f47), .A2(P1_W_R_N_REG_SCAN_IN), .B1(DATAI_5_), .B2(keyinput_f27), .ZN(n20856) );
  OAI221_X1 U23777 ( .B1(keyinput_f47), .B2(P1_W_R_N_REG_SCAN_IN), .C1(
        DATAI_5_), .C2(keyinput_f27), .A(n20856), .ZN(n20947) );
  AOI22_X1 U23778 ( .A1(DATAI_18_), .A2(keyinput_f14), .B1(DATAI_13_), .B2(
        keyinput_f19), .ZN(n20857) );
  OAI221_X1 U23779 ( .B1(DATAI_18_), .B2(keyinput_f14), .C1(DATAI_13_), .C2(
        keyinput_f19), .A(n20857), .ZN(n20946) );
  AOI22_X1 U23780 ( .A1(keyinput_f33), .A2(HOLD), .B1(n20859), .B2(
        keyinput_f61), .ZN(n20858) );
  OAI221_X1 U23781 ( .B1(keyinput_f33), .B2(HOLD), .C1(n20859), .C2(
        keyinput_f61), .A(n20858), .ZN(n20869) );
  OAI22_X1 U23782 ( .A1(DATAI_7_), .A2(keyinput_f25), .B1(keyinput_f41), .B2(
        P1_M_IO_N_REG_SCAN_IN), .ZN(n20860) );
  AOI221_X1 U23783 ( .B1(DATAI_7_), .B2(keyinput_f25), .C1(
        P1_M_IO_N_REG_SCAN_IN), .C2(keyinput_f41), .A(n20860), .ZN(n20867) );
  OAI22_X1 U23784 ( .A1(DATAI_21_), .A2(keyinput_f11), .B1(
        P1_ADS_N_REG_SCAN_IN), .B2(keyinput_f39), .ZN(n20861) );
  AOI221_X1 U23785 ( .B1(DATAI_21_), .B2(keyinput_f11), .C1(keyinput_f39), 
        .C2(P1_ADS_N_REG_SCAN_IN), .A(n20861), .ZN(n20866) );
  OAI22_X1 U23786 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(keyinput_f53), .B1(
        P1_REIP_REG_28__SCAN_IN), .B2(keyinput_f55), .ZN(n20862) );
  AOI221_X1 U23787 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(keyinput_f53), .C1(
        keyinput_f55), .C2(P1_REIP_REG_28__SCAN_IN), .A(n20862), .ZN(n20865)
         );
  OAI22_X1 U23788 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(keyinput_f60), .B1(
        keyinput_f28), .B2(DATAI_4_), .ZN(n20863) );
  AOI221_X1 U23789 ( .B1(P1_REIP_REG_23__SCAN_IN), .B2(keyinput_f60), .C1(
        DATAI_4_), .C2(keyinput_f28), .A(n20863), .ZN(n20864) );
  NAND4_X1 U23790 ( .A1(n20867), .A2(n20866), .A3(n20865), .A4(n20864), .ZN(
        n20868) );
  AOI211_X1 U23791 ( .C1(keyinput_f36), .C2(READY1), .A(n20869), .B(n20868), 
        .ZN(n20870) );
  OAI21_X1 U23792 ( .B1(keyinput_f36), .B2(READY1), .A(n20870), .ZN(n20945) );
  INV_X1 U23793 ( .A(DATAI_22_), .ZN(n20872) );
  AOI22_X1 U23794 ( .A1(n20873), .A2(keyinput_f59), .B1(keyinput_f10), .B2(
        n20872), .ZN(n20871) );
  OAI221_X1 U23795 ( .B1(n20873), .B2(keyinput_f59), .C1(n20872), .C2(
        keyinput_f10), .A(n20871), .ZN(n20882) );
  AOI22_X1 U23796 ( .A1(n21031), .A2(keyinput_f40), .B1(n21008), .B2(
        keyinput_f8), .ZN(n20874) );
  OAI221_X1 U23797 ( .B1(n21031), .B2(keyinput_f40), .C1(n21008), .C2(
        keyinput_f8), .A(n20874), .ZN(n20881) );
  AOI22_X1 U23798 ( .A1(n20877), .A2(keyinput_f63), .B1(keyinput_f7), .B2(
        n20876), .ZN(n20875) );
  OAI221_X1 U23799 ( .B1(n20877), .B2(keyinput_f63), .C1(n20876), .C2(
        keyinput_f7), .A(n20875), .ZN(n20880) );
  INV_X1 U23800 ( .A(DATAI_1_), .ZN(n21023) );
  AOI22_X1 U23801 ( .A1(n21023), .A2(keyinput_f31), .B1(keyinput_f46), .B2(
        n21037), .ZN(n20878) );
  OAI221_X1 U23802 ( .B1(n21023), .B2(keyinput_f31), .C1(n21037), .C2(
        keyinput_f46), .A(n20878), .ZN(n20879) );
  NOR4_X1 U23803 ( .A1(n20882), .A2(n20881), .A3(n20880), .A4(n20879), .ZN(
        n20943) );
  AOI22_X1 U23804 ( .A1(n20885), .A2(keyinput_f5), .B1(keyinput_f50), .B2(
        n20884), .ZN(n20883) );
  OAI221_X1 U23805 ( .B1(n20885), .B2(keyinput_f5), .C1(n20884), .C2(
        keyinput_f50), .A(n20883), .ZN(n20896) );
  AOI22_X1 U23806 ( .A1(n21036), .A2(keyinput_f52), .B1(keyinput_f56), .B2(
        n20887), .ZN(n20886) );
  OAI221_X1 U23807 ( .B1(n21036), .B2(keyinput_f52), .C1(n20887), .C2(
        keyinput_f56), .A(n20886), .ZN(n20895) );
  INV_X1 U23808 ( .A(READY2), .ZN(n20889) );
  AOI22_X1 U23809 ( .A1(n20889), .A2(keyinput_f37), .B1(keyinput_f0), .B2(
        n21033), .ZN(n20888) );
  OAI221_X1 U23810 ( .B1(n20889), .B2(keyinput_f37), .C1(n21033), .C2(
        keyinput_f0), .A(n20888), .ZN(n20894) );
  AOI22_X1 U23811 ( .A1(n20892), .A2(keyinput_f21), .B1(n20891), .B2(
        keyinput_f3), .ZN(n20890) );
  OAI221_X1 U23812 ( .B1(n20892), .B2(keyinput_f21), .C1(n20891), .C2(
        keyinput_f3), .A(n20890), .ZN(n20893) );
  NOR4_X1 U23813 ( .A1(n20896), .A2(n20895), .A3(n20894), .A4(n20893), .ZN(
        n20942) );
  OAI22_X1 U23814 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(keyinput_f57), .B1(
        DATAI_0_), .B2(keyinput_f32), .ZN(n20897) );
  AOI221_X1 U23815 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(keyinput_f57), .C1(
        keyinput_f32), .C2(DATAI_0_), .A(n20897), .ZN(n20904) );
  OAI22_X1 U23816 ( .A1(DATAI_19_), .A2(keyinput_f13), .B1(DATAI_16_), .B2(
        keyinput_f16), .ZN(n20898) );
  AOI221_X1 U23817 ( .B1(DATAI_19_), .B2(keyinput_f13), .C1(keyinput_f16), 
        .C2(DATAI_16_), .A(n20898), .ZN(n20903) );
  OAI22_X1 U23818 ( .A1(DATAI_15_), .A2(keyinput_f17), .B1(
        P1_BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_f51), .ZN(n20899) );
  AOI221_X1 U23819 ( .B1(DATAI_15_), .B2(keyinput_f17), .C1(keyinput_f51), 
        .C2(P1_BYTEENABLE_REG_3__SCAN_IN), .A(n20899), .ZN(n20902) );
  OAI22_X1 U23820 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(keyinput_f58), .B1(
        keyinput_f29), .B2(DATAI_3_), .ZN(n20900) );
  AOI221_X1 U23821 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(keyinput_f58), .C1(
        DATAI_3_), .C2(keyinput_f29), .A(n20900), .ZN(n20901) );
  NAND4_X1 U23822 ( .A1(n20904), .A2(n20903), .A3(n20902), .A4(n20901), .ZN(
        n20940) );
  OAI22_X1 U23823 ( .A1(DATAI_20_), .A2(keyinput_f12), .B1(keyinput_f34), .B2(
        NA), .ZN(n20905) );
  AOI221_X1 U23824 ( .B1(DATAI_20_), .B2(keyinput_f12), .C1(NA), .C2(
        keyinput_f34), .A(n20905), .ZN(n20912) );
  OAI22_X1 U23825 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(keyinput_f44), .B1(
        DATAI_12_), .B2(keyinput_f20), .ZN(n20906) );
  AOI221_X1 U23826 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_f44), .C1(
        keyinput_f20), .C2(DATAI_12_), .A(n20906), .ZN(n20911) );
  OAI22_X1 U23827 ( .A1(DATAI_30_), .A2(keyinput_f2), .B1(keyinput_f4), .B2(
        DATAI_28_), .ZN(n20907) );
  AOI221_X1 U23828 ( .B1(DATAI_30_), .B2(keyinput_f2), .C1(DATAI_28_), .C2(
        keyinput_f4), .A(n20907), .ZN(n20910) );
  OAI22_X1 U23829 ( .A1(DATAI_10_), .A2(keyinput_f22), .B1(
        P1_REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_f43), .ZN(n20908) );
  AOI221_X1 U23830 ( .B1(DATAI_10_), .B2(keyinput_f22), .C1(keyinput_f43), 
        .C2(P1_REQUESTPENDING_REG_SCAN_IN), .A(n20908), .ZN(n20909) );
  NAND4_X1 U23831 ( .A1(n20912), .A2(n20911), .A3(n20910), .A4(n20909), .ZN(
        n20939) );
  INV_X1 U23832 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n20914) );
  OAI22_X1 U23833 ( .A1(n20915), .A2(keyinput_f23), .B1(n20914), .B2(
        keyinput_f38), .ZN(n20913) );
  AOI221_X1 U23834 ( .B1(n20915), .B2(keyinput_f23), .C1(keyinput_f38), .C2(
        n20914), .A(n20913), .ZN(n20926) );
  OAI22_X1 U23835 ( .A1(n20918), .A2(keyinput_f1), .B1(n20917), .B2(
        keyinput_f54), .ZN(n20916) );
  AOI221_X1 U23836 ( .B1(n20918), .B2(keyinput_f1), .C1(keyinput_f54), .C2(
        n20917), .A(n20916), .ZN(n20925) );
  OAI22_X1 U23837 ( .A1(n21034), .A2(keyinput_f18), .B1(n20920), .B2(
        keyinput_f35), .ZN(n20919) );
  AOI221_X1 U23838 ( .B1(n21034), .B2(keyinput_f18), .C1(keyinput_f35), .C2(
        n20920), .A(n20919), .ZN(n20924) );
  INV_X1 U23839 ( .A(keyinput_f48), .ZN(n20922) );
  OAI22_X1 U23840 ( .A1(n21039), .A2(keyinput_f45), .B1(n20922), .B2(
        P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20921) );
  AOI221_X1 U23841 ( .B1(n21039), .B2(keyinput_f45), .C1(
        P1_BYTEENABLE_REG_0__SCAN_IN), .C2(n20922), .A(n20921), .ZN(n20923) );
  NAND4_X1 U23842 ( .A1(n20926), .A2(n20925), .A3(n20924), .A4(n20923), .ZN(
        n20938) );
  OAI22_X1 U23843 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(keyinput_f62), .B1(
        keyinput_f15), .B2(DATAI_17_), .ZN(n20927) );
  AOI221_X1 U23844 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(keyinput_f62), .C1(
        DATAI_17_), .C2(keyinput_f15), .A(n20927), .ZN(n20936) );
  OAI22_X1 U23845 ( .A1(DATAI_23_), .A2(keyinput_f9), .B1(
        P1_BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_f49), .ZN(n20928) );
  AOI221_X1 U23846 ( .B1(DATAI_23_), .B2(keyinput_f9), .C1(keyinput_f49), .C2(
        P1_BYTEENABLE_REG_1__SCAN_IN), .A(n20928), .ZN(n20935) );
  OAI22_X1 U23847 ( .A1(n20931), .A2(keyinput_f6), .B1(n20930), .B2(
        keyinput_f24), .ZN(n20929) );
  AOI221_X1 U23848 ( .B1(n20931), .B2(keyinput_f6), .C1(keyinput_f24), .C2(
        n20930), .A(n20929), .ZN(n20934) );
  OAI22_X1 U23849 ( .A1(n20960), .A2(keyinput_f26), .B1(P1_D_C_N_REG_SCAN_IN), 
        .B2(keyinput_f42), .ZN(n20932) );
  AOI221_X1 U23850 ( .B1(n20960), .B2(keyinput_f26), .C1(keyinput_f42), .C2(
        P1_D_C_N_REG_SCAN_IN), .A(n20932), .ZN(n20933) );
  NAND4_X1 U23851 ( .A1(n20936), .A2(n20935), .A3(n20934), .A4(n20933), .ZN(
        n20937) );
  NOR4_X1 U23852 ( .A1(n20940), .A2(n20939), .A3(n20938), .A4(n20937), .ZN(
        n20941) );
  NAND3_X1 U23853 ( .A1(n20943), .A2(n20942), .A3(n20941), .ZN(n20944) );
  NOR4_X1 U23854 ( .A1(n20947), .A2(n20946), .A3(n20945), .A4(n20944), .ZN(
        n20948) );
  AOI221_X1 U23855 ( .B1(DATAI_2_), .B2(keyinput_f30), .C1(n20950), .C2(n20949), .A(n20948), .ZN(n21052) );
  AOI22_X1 U23856 ( .A1(P1_BYTEENABLE_REG_2__SCAN_IN), .A2(keyinput_g50), .B1(
        DATAI_7_), .B2(keyinput_g25), .ZN(n20951) );
  OAI221_X1 U23857 ( .B1(P1_BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_g50), 
        .C1(DATAI_7_), .C2(keyinput_g25), .A(n20951), .ZN(n20958) );
  AOI22_X1 U23858 ( .A1(READY2), .A2(keyinput_g37), .B1(
        P1_REIP_REG_21__SCAN_IN), .B2(keyinput_g62), .ZN(n20952) );
  OAI221_X1 U23859 ( .B1(READY2), .B2(keyinput_g37), .C1(
        P1_REIP_REG_21__SCAN_IN), .C2(keyinput_g62), .A(n20952), .ZN(n20957)
         );
  AOI22_X1 U23860 ( .A1(P1_W_R_N_REG_SCAN_IN), .A2(keyinput_g47), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(keyinput_g63), .ZN(n20953) );
  OAI221_X1 U23861 ( .B1(P1_W_R_N_REG_SCAN_IN), .B2(keyinput_g47), .C1(
        P1_REIP_REG_20__SCAN_IN), .C2(keyinput_g63), .A(n20953), .ZN(n20956)
         );
  AOI22_X1 U23862 ( .A1(DATAI_9_), .A2(keyinput_g23), .B1(
        P1_REIP_REG_27__SCAN_IN), .B2(keyinput_g56), .ZN(n20954) );
  OAI221_X1 U23863 ( .B1(DATAI_9_), .B2(keyinput_g23), .C1(
        P1_REIP_REG_27__SCAN_IN), .C2(keyinput_g56), .A(n20954), .ZN(n20955)
         );
  NOR4_X1 U23864 ( .A1(n20958), .A2(n20957), .A3(n20956), .A4(n20955), .ZN(
        n20986) );
  XNOR2_X1 U23865 ( .A(NA), .B(keyinput_g34), .ZN(n20966) );
  AOI22_X1 U23866 ( .A1(BS16), .A2(keyinput_g35), .B1(n20960), .B2(
        keyinput_g26), .ZN(n20959) );
  OAI221_X1 U23867 ( .B1(BS16), .B2(keyinput_g35), .C1(n20960), .C2(
        keyinput_g26), .A(n20959), .ZN(n20965) );
  AOI22_X1 U23868 ( .A1(DATAI_8_), .A2(keyinput_g24), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(keyinput_g61), .ZN(n20961) );
  OAI221_X1 U23869 ( .B1(DATAI_8_), .B2(keyinput_g24), .C1(
        P1_REIP_REG_22__SCAN_IN), .C2(keyinput_g61), .A(n20961), .ZN(n20964)
         );
  AOI22_X1 U23870 ( .A1(P1_BYTEENABLE_REG_0__SCAN_IN), .A2(keyinput_g48), .B1(
        P1_BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_g51), .ZN(n20962) );
  OAI221_X1 U23871 ( .B1(P1_BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_g48), 
        .C1(P1_BYTEENABLE_REG_3__SCAN_IN), .C2(keyinput_g51), .A(n20962), .ZN(
        n20963) );
  NOR4_X1 U23872 ( .A1(n20966), .A2(n20965), .A3(n20964), .A4(n20963), .ZN(
        n20985) );
  AOI22_X1 U23873 ( .A1(DATAI_4_), .A2(keyinput_g28), .B1(DATAI_10_), .B2(
        keyinput_g22), .ZN(n20967) );
  OAI221_X1 U23874 ( .B1(DATAI_4_), .B2(keyinput_g28), .C1(DATAI_10_), .C2(
        keyinput_g22), .A(n20967), .ZN(n20974) );
  AOI22_X1 U23875 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(keyinput_g59), .B1(
        P1_REIP_REG_29__SCAN_IN), .B2(keyinput_g54), .ZN(n20968) );
  OAI221_X1 U23876 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(keyinput_g59), .C1(
        P1_REIP_REG_29__SCAN_IN), .C2(keyinput_g54), .A(n20968), .ZN(n20973)
         );
  AOI22_X1 U23877 ( .A1(DATAI_22_), .A2(keyinput_g10), .B1(DATAI_29_), .B2(
        keyinput_g3), .ZN(n20969) );
  OAI221_X1 U23878 ( .B1(DATAI_22_), .B2(keyinput_g10), .C1(DATAI_29_), .C2(
        keyinput_g3), .A(n20969), .ZN(n20972) );
  AOI22_X1 U23879 ( .A1(DATAI_26_), .A2(keyinput_g6), .B1(
        P1_REIP_REG_25__SCAN_IN), .B2(keyinput_g58), .ZN(n20970) );
  OAI221_X1 U23880 ( .B1(DATAI_26_), .B2(keyinput_g6), .C1(
        P1_REIP_REG_25__SCAN_IN), .C2(keyinput_g58), .A(n20970), .ZN(n20971)
         );
  NOR4_X1 U23881 ( .A1(n20974), .A2(n20973), .A3(n20972), .A4(n20971), .ZN(
        n20984) );
  AOI22_X1 U23882 ( .A1(DATAI_25_), .A2(keyinput_g7), .B1(DATAI_12_), .B2(
        keyinput_g20), .ZN(n20975) );
  OAI221_X1 U23883 ( .B1(DATAI_25_), .B2(keyinput_g7), .C1(DATAI_12_), .C2(
        keyinput_g20), .A(n20975), .ZN(n20982) );
  AOI22_X1 U23884 ( .A1(P1_BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput_g49), .B1(
        DATAI_3_), .B2(keyinput_g29), .ZN(n20976) );
  OAI221_X1 U23885 ( .B1(P1_BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_g49), 
        .C1(DATAI_3_), .C2(keyinput_g29), .A(n20976), .ZN(n20981) );
  AOI22_X1 U23886 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(keyinput_g39), .B1(
        P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_g44), .ZN(n20977) );
  OAI221_X1 U23887 ( .B1(P1_ADS_N_REG_SCAN_IN), .B2(keyinput_g39), .C1(
        P1_STATEBS16_REG_SCAN_IN), .C2(keyinput_g44), .A(n20977), .ZN(n20980)
         );
  AOI22_X1 U23888 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(keyinput_g57), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(keyinput_g60), .ZN(n20978) );
  OAI221_X1 U23889 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(keyinput_g57), .C1(
        P1_REIP_REG_23__SCAN_IN), .C2(keyinput_g60), .A(n20978), .ZN(n20979)
         );
  NOR4_X1 U23890 ( .A1(n20982), .A2(n20981), .A3(n20980), .A4(n20979), .ZN(
        n20983) );
  NAND4_X1 U23891 ( .A1(n20986), .A2(n20985), .A3(n20984), .A4(n20983), .ZN(
        n21050) );
  INV_X1 U23892 ( .A(DATAI_20_), .ZN(n20988) );
  AOI22_X1 U23893 ( .A1(n20989), .A2(keyinput_g19), .B1(keyinput_g12), .B2(
        n20988), .ZN(n20987) );
  OAI221_X1 U23894 ( .B1(n20989), .B2(keyinput_g19), .C1(n20988), .C2(
        keyinput_g12), .A(n20987), .ZN(n21001) );
  INV_X1 U23895 ( .A(DATAI_19_), .ZN(n20991) );
  AOI22_X1 U23896 ( .A1(n20992), .A2(keyinput_g41), .B1(n20991), .B2(
        keyinput_g13), .ZN(n20990) );
  OAI221_X1 U23897 ( .B1(n20992), .B2(keyinput_g41), .C1(n20991), .C2(
        keyinput_g13), .A(n20990), .ZN(n21000) );
  INV_X1 U23898 ( .A(READY1), .ZN(n20994) );
  AOI22_X1 U23899 ( .A1(n20995), .A2(keyinput_g4), .B1(n20994), .B2(
        keyinput_g36), .ZN(n20993) );
  OAI221_X1 U23900 ( .B1(n20995), .B2(keyinput_g4), .C1(n20994), .C2(
        keyinput_g36), .A(n20993), .ZN(n20999) );
  INV_X1 U23901 ( .A(DATAI_16_), .ZN(n20997) );
  AOI22_X1 U23902 ( .A1(n14482), .A2(keyinput_g15), .B1(keyinput_g16), .B2(
        n20997), .ZN(n20996) );
  OAI221_X1 U23903 ( .B1(n14482), .B2(keyinput_g15), .C1(n20997), .C2(
        keyinput_g16), .A(n20996), .ZN(n20998) );
  NOR4_X1 U23904 ( .A1(n21001), .A2(n21000), .A3(n20999), .A4(n20998), .ZN(
        n21048) );
  AOI22_X1 U23905 ( .A1(P1_READREQUEST_REG_SCAN_IN), .A2(keyinput_g38), .B1(
        DATAI_31_), .B2(keyinput_g1), .ZN(n21002) );
  OAI221_X1 U23906 ( .B1(P1_READREQUEST_REG_SCAN_IN), .B2(keyinput_g38), .C1(
        DATAI_31_), .C2(keyinput_g1), .A(n21002), .ZN(n21013) );
  AOI22_X1 U23907 ( .A1(DATAI_11_), .A2(keyinput_g21), .B1(DATAI_27_), .B2(
        keyinput_g5), .ZN(n21003) );
  OAI221_X1 U23908 ( .B1(DATAI_11_), .B2(keyinput_g21), .C1(DATAI_27_), .C2(
        keyinput_g5), .A(n21003), .ZN(n21012) );
  AOI22_X1 U23909 ( .A1(n21006), .A2(keyinput_g53), .B1(keyinput_g55), .B2(
        n21005), .ZN(n21004) );
  OAI221_X1 U23910 ( .B1(n21006), .B2(keyinput_g53), .C1(n21005), .C2(
        keyinput_g55), .A(n21004), .ZN(n21011) );
  AOI22_X1 U23911 ( .A1(n21009), .A2(keyinput_g2), .B1(keyinput_g8), .B2(
        n21008), .ZN(n21007) );
  OAI221_X1 U23912 ( .B1(n21009), .B2(keyinput_g2), .C1(n21008), .C2(
        keyinput_g8), .A(n21007), .ZN(n21010) );
  NOR4_X1 U23913 ( .A1(n21013), .A2(n21012), .A3(n21011), .A4(n21010), .ZN(
        n21047) );
  INV_X1 U23914 ( .A(DATAI_0_), .ZN(n21015) );
  AOI22_X1 U23915 ( .A1(n21016), .A2(keyinput_g33), .B1(n21015), .B2(
        keyinput_g32), .ZN(n21014) );
  OAI221_X1 U23916 ( .B1(n21016), .B2(keyinput_g33), .C1(n21015), .C2(
        keyinput_g32), .A(n21014), .ZN(n21028) );
  INV_X1 U23917 ( .A(DATAI_23_), .ZN(n21019) );
  INV_X1 U23918 ( .A(DATAI_18_), .ZN(n21018) );
  AOI22_X1 U23919 ( .A1(n21019), .A2(keyinput_g9), .B1(keyinput_g14), .B2(
        n21018), .ZN(n21017) );
  OAI221_X1 U23920 ( .B1(n21019), .B2(keyinput_g9), .C1(n21018), .C2(
        keyinput_g14), .A(n21017), .ZN(n21027) );
  AOI22_X1 U23921 ( .A1(n21021), .A2(keyinput_g43), .B1(n13022), .B2(
        keyinput_g17), .ZN(n21020) );
  OAI221_X1 U23922 ( .B1(n21021), .B2(keyinput_g43), .C1(n13022), .C2(
        keyinput_g17), .A(n21020), .ZN(n21026) );
  AOI22_X1 U23923 ( .A1(n21024), .A2(keyinput_g42), .B1(n21023), .B2(
        keyinput_g31), .ZN(n21022) );
  OAI221_X1 U23924 ( .B1(n21024), .B2(keyinput_g42), .C1(n21023), .C2(
        keyinput_g31), .A(n21022), .ZN(n21025) );
  NOR4_X1 U23925 ( .A1(n21028), .A2(n21027), .A3(n21026), .A4(n21025), .ZN(
        n21046) );
  INV_X1 U23926 ( .A(DATAI_5_), .ZN(n21030) );
  AOI22_X1 U23927 ( .A1(n21031), .A2(keyinput_g40), .B1(n21030), .B2(
        keyinput_g27), .ZN(n21029) );
  OAI221_X1 U23928 ( .B1(n21031), .B2(keyinput_g40), .C1(n21030), .C2(
        keyinput_g27), .A(n21029), .ZN(n21044) );
  AOI22_X1 U23929 ( .A1(n21034), .A2(keyinput_g18), .B1(keyinput_g0), .B2(
        n21033), .ZN(n21032) );
  OAI221_X1 U23930 ( .B1(n21034), .B2(keyinput_g18), .C1(n21033), .C2(
        keyinput_g0), .A(n21032), .ZN(n21043) );
  AOI22_X1 U23931 ( .A1(n21037), .A2(keyinput_g46), .B1(n21036), .B2(
        keyinput_g52), .ZN(n21035) );
  OAI221_X1 U23932 ( .B1(n21037), .B2(keyinput_g46), .C1(n21036), .C2(
        keyinput_g52), .A(n21035), .ZN(n21042) );
  INV_X1 U23933 ( .A(DATAI_21_), .ZN(n21040) );
  AOI22_X1 U23934 ( .A1(n21040), .A2(keyinput_g11), .B1(keyinput_g45), .B2(
        n21039), .ZN(n21038) );
  OAI221_X1 U23935 ( .B1(n21040), .B2(keyinput_g11), .C1(n21039), .C2(
        keyinput_g45), .A(n21038), .ZN(n21041) );
  NOR4_X1 U23936 ( .A1(n21044), .A2(n21043), .A3(n21042), .A4(n21041), .ZN(
        n21045) );
  NAND4_X1 U23937 ( .A1(n21048), .A2(n21047), .A3(n21046), .A4(n21045), .ZN(
        n21049) );
  OAI22_X1 U23938 ( .A1(DATAI_2_), .A2(keyinput_g30), .B1(n21050), .B2(n21049), 
        .ZN(n21051) );
  AOI211_X1 U23939 ( .C1(DATAI_2_), .C2(keyinput_g30), .A(n21052), .B(n21051), 
        .ZN(n21054) );
  AOI22_X1 U23940 ( .A1(n16776), .A2(P3_ADDRESS_REG_29__SCAN_IN), .B1(
        P2_ADDRESS_REG_29__SCAN_IN), .B2(n16778), .ZN(n21053) );
  XNOR2_X1 U23941 ( .A(n21054), .B(n21053), .ZN(U355) );
  AND2_X1 U14176 ( .A1(n11008), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11014) );
  AND2_X1 U11228 ( .A1(n11009), .A2(n13344), .ZN(n11112) );
  BUF_X2 U11103 ( .A(n11112), .Z(n11805) );
  XNOR2_X1 U11175 ( .A(n12023), .B(n10020), .ZN(n12421) );
  NAND2_X1 U15552 ( .A1(n12452), .A2(n12424), .ZN(n19875) );
  NAND2_X1 U15569 ( .A1(n12452), .A2(n12451), .ZN(n12535) );
  OR2_X1 U15563 ( .A1(n12439), .A2(n12450), .ZN(n19697) );
  INV_X1 U11444 ( .A(n12449), .ZN(n12452) );
  OR2_X1 U15557 ( .A1(n12439), .A2(n12448), .ZN(n12540) );
  OR2_X1 U15566 ( .A1(n12449), .A2(n12448), .ZN(n12521) );
  CLKBUF_X1 U11102 ( .A(n12421), .Z(n12980) );
  NAND3_X1 U11104 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13524) );
  CLKBUF_X1 U11106 ( .A(n12029), .Z(n12422) );
  CLKBUF_X1 U11112 ( .A(n10650), .Z(n13549) );
  CLKBUF_X1 U11126 ( .A(n17211), .Z(n9651) );
  CLKBUF_X1 U11128 ( .A(n13971), .Z(n17456) );
  AND2_X1 U11130 ( .A1(n11153), .A2(n11133), .ZN(n13071) );
  CLKBUF_X1 U11180 ( .A(n11155), .Z(n14788) );
  CLKBUF_X1 U11186 ( .A(n11153), .Z(n13622) );
  CLKBUF_X1 U11213 ( .A(n10608), .Z(n12765) );
  CLKBUF_X1 U11223 ( .A(n20116), .Z(n20122) );
  CLKBUF_X1 U11721 ( .A(n16768), .Z(n16772) );
  CLKBUF_X1 U11973 ( .A(n17761), .Z(n17765) );
endmodule

