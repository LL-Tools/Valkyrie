

module b14_C_SARLock_k_128_9 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910;

  INV_X2 U2400 ( .A(n2832), .ZN(n3001) );
  AND2_X4 U2401 ( .A1(n4686), .A2(n3031), .ZN(n2483) );
  NOR2_X1 U2402 ( .A1(n4686), .A2(n3031), .ZN(n2499) );
  NAND2_X1 U2403 ( .A1(n2423), .A2(IR_REG_31__SCAN_IN), .ZN(n2424) );
  INV_X1 U2404 ( .A(n3003), .ZN(n2558) );
  INV_X1 U2406 ( .A(IR_REG_31__SCAN_IN), .ZN(n2561) );
  AOI21_X1 U2407 ( .B1(n3693), .B2(n3690), .A(n3689), .ZN(n3767) );
  NOR2_X2 U2408 ( .A1(n2489), .A2(n2488), .ZN(n2908) );
  XNOR2_X2 U2409 ( .A(n2490), .B(IR_REG_2__SCAN_IN), .ZN(n4698) );
  XNOR2_X2 U2410 ( .A(n2424), .B(IR_REG_24__SCAN_IN), .ZN(n2852) );
  NAND2_X1 U2411 ( .A1(n3140), .A2(n2907), .ZN(n3245) );
  NAND2_X2 U2412 ( .A1(n3870), .A2(n3867), .ZN(n2943) );
  NAND4_X1 U2413 ( .A1(n2503), .A2(n2502), .A3(n2501), .A4(n2500), .ZN(n4238)
         );
  CLKBUF_X2 U2414 ( .A(n2158), .Z(n2533) );
  BUF_X2 U2415 ( .A(n2499), .Z(n2158) );
  BUF_X2 U2416 ( .A(n2171), .Z(n2700) );
  OAI21_X1 U2417 ( .B1(n3720), .B2(n3721), .A(n3718), .ZN(n3693) );
  AND2_X1 U2418 ( .A1(n2338), .A2(n2337), .ZN(n3720) );
  MUX2_X1 U2419 ( .A(REG1_REG_28__SCAN_IN), .B(n2996), .S(n4910), .Z(n2989) );
  MUX2_X1 U2420 ( .A(REG0_REG_28__SCAN_IN), .B(n2996), .S(n4902), .Z(n2997) );
  AND2_X1 U2421 ( .A1(n2376), .A2(n2184), .ZN(n4337) );
  NAND2_X1 U2422 ( .A1(n4514), .A2(n2931), .ZN(n4489) );
  NAND2_X1 U2423 ( .A1(n4513), .A2(n4515), .ZN(n4514) );
  NAND2_X1 U2424 ( .A1(n2317), .A2(n3492), .ZN(n3538) );
  NAND2_X1 U2425 ( .A1(n2290), .A2(n2173), .ZN(n3485) );
  AOI21_X1 U2426 ( .B1(n2309), .B2(n2311), .A(n2174), .ZN(n2306) );
  OAI21_X1 U2427 ( .B1(n2313), .B2(n2311), .A(n3307), .ZN(n2310) );
  OR2_X1 U2428 ( .A1(n2516), .A2(n3211), .ZN(n2517) );
  AOI21_X1 U2429 ( .B1(n2352), .B2(n2351), .A(n2162), .ZN(n2350) );
  NOR2_X2 U2430 ( .A1(n3047), .A2(n3048), .ZN(n4775) );
  INV_X1 U2431 ( .A(n3624), .ZN(n4237) );
  NAND2_X1 U2432 ( .A1(n2452), .A2(n2451), .ZN(n2944) );
  AND4_X1 U2433 ( .A1(n2537), .A2(n2536), .A3(n2535), .A4(n2534), .ZN(n3624)
         );
  AND4_X1 U2434 ( .A1(n2525), .A2(n2524), .A3(n2523), .A4(n2522), .ZN(n3238)
         );
  AOI21_X1 U2435 ( .B1(n4272), .B2(REG2_REG_4__SCAN_IN), .A(n2276), .ZN(n3122)
         );
  XNOR2_X1 U2436 ( .A(n2437), .B(n2436), .ZN(n3929) );
  XNOR2_X1 U2437 ( .A(n2439), .B(IR_REG_21__SCAN_IN), .ZN(n4689) );
  AOI21_X1 U2438 ( .B1(n2428), .B2(IR_REG_26__SCAN_IN), .A(n2427), .ZN(n2429)
         );
  NAND2_X1 U2439 ( .A1(n2389), .A2(IR_REG_31__SCAN_IN), .ZN(n2442) );
  INV_X1 U2440 ( .A(n2435), .ZN(n2421) );
  AND3_X1 U2441 ( .A1(n2214), .A2(n2212), .A3(n2384), .ZN(n2425) );
  INV_X1 U2442 ( .A(n2208), .ZN(n2441) );
  AND3_X1 U2443 ( .A1(n2539), .A2(n2400), .A3(n2401), .ZN(n2213) );
  AND2_X1 U2444 ( .A1(n2169), .A2(n2231), .ZN(n2210) );
  NOR2_X1 U2445 ( .A1(n2411), .A2(n2410), .ZN(n2412) );
  INV_X1 U2446 ( .A(IR_REG_2__SCAN_IN), .ZN(n2399) );
  INV_X1 U2447 ( .A(IR_REG_20__SCAN_IN), .ZN(n2436) );
  NOR2_X1 U2448 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2402)
         );
  NOR2_X1 U2449 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2403)
         );
  NOR2_X1 U2450 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2404)
         );
  NOR2_X1 U2451 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2405)
         );
  NAND2_X4 U2452 ( .A1(n2454), .A2(n2468), .ZN(n2477) );
  NAND2_X2 U2453 ( .A1(n2852), .A2(n2434), .ZN(n2454) );
  NOR2_X1 U2454 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2401)
         );
  AND4_X1 U2455 ( .A1(n2399), .A2(n2398), .A3(n2397), .A4(n2505), .ZN(n2564)
         );
  INV_X1 U2456 ( .A(IR_REG_6__SCAN_IN), .ZN(n2397) );
  NOR2_X1 U2457 ( .A1(n4235), .A2(n3414), .ZN(n2925) );
  AND2_X1 U2458 ( .A1(n2923), .A2(n2176), .ZN(n2381) );
  NAND2_X1 U2459 ( .A1(n2175), .A2(n2916), .ZN(n2353) );
  NAND2_X1 U2460 ( .A1(n3701), .A2(n2303), .ZN(n2302) );
  NAND2_X1 U2461 ( .A1(n2724), .A2(n3777), .ZN(n2303) );
  XNOR2_X1 U2462 ( .A(n2528), .B(n3001), .ZN(n2531) );
  OAI22_X1 U2463 ( .A1(n3238), .A2(n2749), .B1(n2477), .B2(n3615), .ZN(n2528)
         );
  NOR2_X1 U2464 ( .A1(n2866), .A2(n3026), .ZN(n2434) );
  NAND2_X1 U2465 ( .A1(n4789), .A2(n2275), .ZN(n4806) );
  OR2_X1 U2466 ( .A1(n4301), .A2(REG2_REG_17__SCAN_IN), .ZN(n2275) );
  NOR2_X1 U2467 ( .A1(n4806), .A2(n4807), .ZN(n4805) );
  INV_X1 U2468 ( .A(n2370), .ZN(n2368) );
  OR2_X1 U2469 ( .A1(n2182), .A2(n2375), .ZN(n2369) );
  NAND2_X1 U2470 ( .A1(n2370), .A2(n2367), .ZN(n2366) );
  AND2_X1 U2471 ( .A1(n2940), .A2(n2184), .ZN(n2375) );
  NOR2_X1 U2472 ( .A1(n2374), .A2(n2185), .ZN(n2372) );
  AOI22_X1 U2473 ( .A1(n4411), .A2(n2936), .B1(n3724), .B2(n4419), .ZN(n4391)
         );
  OR2_X1 U2474 ( .A1(n3939), .A2(n4524), .ZN(n2931) );
  NAND2_X1 U2475 ( .A1(n3197), .A2(n2912), .ZN(n2383) );
  AND2_X1 U2476 ( .A1(n2941), .A2(n3862), .ZN(n3150) );
  NOR2_X1 U2477 ( .A1(IR_REG_27__SCAN_IN), .A2(IR_REG_28__SCAN_IN), .ZN(n2440)
         );
  INV_X1 U2478 ( .A(IR_REG_23__SCAN_IN), .ZN(n2870) );
  INV_X1 U2479 ( .A(n3790), .ZN(n3757) );
  INV_X1 U2480 ( .A(IR_REG_22__SCAN_IN), .ZN(n2422) );
  NOR2_X1 U2481 ( .A1(n2609), .A2(n2406), .ZN(n2385) );
  INV_X1 U2482 ( .A(n3493), .ZN(n2322) );
  INV_X1 U2483 ( .A(n2325), .ZN(n2316) );
  NAND2_X1 U2484 ( .A1(n2327), .A2(n2326), .ZN(n2325) );
  INV_X1 U2485 ( .A(n3425), .ZN(n2326) );
  INV_X1 U2486 ( .A(n3424), .ZN(n2327) );
  NAND2_X1 U2487 ( .A1(n2280), .A2(n2279), .ZN(n2278) );
  NAND2_X1 U2488 ( .A1(n3076), .A2(n4697), .ZN(n2279) );
  NAND2_X1 U2489 ( .A1(n3100), .A2(REG2_REG_3__SCAN_IN), .ZN(n2280) );
  AOI21_X1 U2490 ( .B1(REG1_REG_9__SCAN_IN), .B2(n3467), .A(n4709), .ZN(n3469)
         );
  AOI21_X1 U2491 ( .B1(n4855), .B2(REG1_REG_11__SCAN_IN), .A(n4728), .ZN(n3471) );
  NOR2_X1 U2492 ( .A1(n4767), .A2(n2289), .ZN(n4299) );
  AND2_X1 U2493 ( .A1(n4298), .A2(REG2_REG_15__SCAN_IN), .ZN(n2289) );
  NOR2_X1 U2494 ( .A1(n2182), .A2(n2371), .ZN(n2370) );
  INV_X1 U2495 ( .A(n2372), .ZN(n2371) );
  NAND2_X1 U2496 ( .A1(n2206), .A2(n2967), .ZN(n2205) );
  INV_X1 U2497 ( .A(n3916), .ZN(n2206) );
  AND2_X1 U2498 ( .A1(n4326), .A2(n2992), .ZN(n4313) );
  OR2_X1 U2499 ( .A1(n4394), .A2(n2205), .ZN(n2203) );
  AOI21_X1 U2500 ( .B1(n4452), .B2(n3914), .A(n3814), .ZN(n4394) );
  INV_X1 U2501 ( .A(n2346), .ZN(n2344) );
  INV_X1 U2502 ( .A(n3809), .ZN(n2219) );
  NAND2_X1 U2503 ( .A1(n2905), .A2(n2904), .ZN(n3870) );
  NAND2_X1 U2504 ( .A1(n3871), .A2(n3874), .ZN(n2946) );
  AND2_X1 U2505 ( .A1(n3929), .A2(n4689), .ZN(n3191) );
  NOR2_X1 U2506 ( .A1(n3614), .A2(n3241), .ZN(n3228) );
  OR2_X1 U2507 ( .A1(n2441), .A2(n2561), .ZN(n3035) );
  AND2_X1 U2508 ( .A1(n2564), .A2(n2413), .ZN(n2211) );
  AND2_X1 U2509 ( .A1(n2412), .A2(n2210), .ZN(n2209) );
  NAND2_X1 U2510 ( .A1(n2421), .A2(n2328), .ZN(n2330) );
  AND2_X1 U2511 ( .A1(n2420), .A2(n2329), .ZN(n2328) );
  OR2_X1 U2512 ( .A1(n2705), .A2(IR_REG_14__SCAN_IN), .ZN(n2706) );
  OR2_X1 U2513 ( .A1(n3297), .A2(n3296), .ZN(n2313) );
  INV_X1 U2514 ( .A(n3538), .ZN(n2681) );
  INV_X1 U2515 ( .A(n3650), .ZN(n2339) );
  NAND2_X1 U2516 ( .A1(n2334), .A2(n3678), .ZN(n2333) );
  XNOR2_X1 U2517 ( .A(n2510), .B(n3001), .ZN(n2515) );
  NAND2_X1 U2518 ( .A1(n2947), .A2(n2846), .ZN(n2296) );
  INV_X1 U2519 ( .A(n2301), .ZN(n2300) );
  OAI21_X1 U2520 ( .B1(n2302), .B2(n2304), .A(n2727), .ZN(n2301) );
  NAND2_X1 U2521 ( .A1(n2305), .A2(n3700), .ZN(n2304) );
  INV_X1 U2522 ( .A(n3581), .ZN(n2696) );
  NOR2_X1 U2523 ( .A1(n2760), .A2(n3661), .ZN(n2761) );
  OR2_X1 U2524 ( .A1(n2757), .A2(n3660), .ZN(n2762) );
  AND2_X1 U2525 ( .A1(n2750), .A2(REG3_REG_19__SCAN_IN), .ZN(n2763) );
  NAND2_X1 U2526 ( .A1(n3424), .A2(n3425), .ZN(n2323) );
  NOR2_X1 U2527 ( .A1(n3744), .A2(n2335), .ZN(n2334) );
  INV_X1 U2528 ( .A(n3679), .ZN(n2335) );
  NOR2_X1 U2529 ( .A1(n2637), .A2(n2636), .ZN(n2646) );
  INV_X1 U2530 ( .A(n2483), .ZN(n2972) );
  INV_X1 U2531 ( .A(n2975), .ZN(n3793) );
  XNOR2_X1 U2532 ( .A(n2278), .B(n2277), .ZN(n4272) );
  INV_X1 U2533 ( .A(n4696), .ZN(n2277) );
  NAND2_X1 U2534 ( .A1(n3064), .A2(n3063), .ZN(n3066) );
  INV_X1 U2535 ( .A(IR_REG_5__SCAN_IN), .ZN(n2400) );
  NAND2_X1 U2536 ( .A1(n3088), .A2(n2270), .ZN(n2268) );
  NOR2_X1 U2537 ( .A1(n3159), .A2(n2271), .ZN(n2270) );
  OR2_X1 U2538 ( .A1(n2272), .A2(n3159), .ZN(n2267) );
  INV_X1 U2539 ( .A(n2250), .ZN(n2247) );
  NAND2_X1 U2540 ( .A1(n2159), .A2(n3095), .ZN(n2243) );
  NAND2_X1 U2541 ( .A1(n2251), .A2(n4692), .ZN(n2250) );
  INV_X1 U2542 ( .A(n3096), .ZN(n2251) );
  OR2_X1 U2543 ( .A1(n3155), .A2(n2244), .ZN(n2248) );
  NAND2_X1 U2544 ( .A1(n4692), .A2(n2245), .ZN(n2244) );
  INV_X1 U2545 ( .A(n3095), .ZN(n2245) );
  OR2_X1 U2546 ( .A1(n3155), .A2(n3095), .ZN(n2253) );
  NAND2_X1 U2547 ( .A1(n4732), .A2(n3458), .ZN(n3460) );
  OAI21_X1 U2548 ( .B1(n4294), .B2(n4293), .A(n2283), .ZN(n4295) );
  OR2_X1 U2549 ( .A1(n4292), .A2(REG2_REG_13__SCAN_IN), .ZN(n2283) );
  XNOR2_X1 U2550 ( .A(n4299), .B(n2720), .ZN(n4780) );
  NAND2_X1 U2551 ( .A1(n4780), .A2(n3596), .ZN(n4779) );
  NOR2_X1 U2552 ( .A1(n4762), .A2(n2240), .ZN(n4287) );
  AND2_X1 U2553 ( .A1(n4298), .A2(REG1_REG_15__SCAN_IN), .ZN(n2240) );
  OR2_X1 U2554 ( .A1(n2887), .A2(n3014), .ZN(n4311) );
  NOR2_X1 U2555 ( .A1(n4384), .A2(n2233), .ZN(n4570) );
  NAND2_X1 U2556 ( .A1(n2235), .A2(n2234), .ZN(n2233) );
  NOR2_X1 U2557 ( .A1(n4333), .A2(n2991), .ZN(n2234) );
  OR2_X1 U2558 ( .A1(n4423), .A2(n3746), .ZN(n2935) );
  AND2_X1 U2559 ( .A1(n2167), .A2(n2933), .ZN(n2346) );
  AND2_X1 U2560 ( .A1(n3940), .A2(n3714), .ZN(n2929) );
  AOI21_X1 U2561 ( .B1(n3516), .B2(n2926), .A(n2181), .ZN(n3548) );
  NAND2_X1 U2562 ( .A1(n3408), .A2(n2955), .ZN(n2926) );
  NAND2_X1 U2563 ( .A1(n3548), .A2(n3549), .ZN(n3547) );
  AOI21_X1 U2564 ( .B1(n2179), .B2(n2381), .A(n2163), .ZN(n2380) );
  NAND2_X1 U2565 ( .A1(n3368), .A2(n2381), .ZN(n2379) );
  INV_X1 U2566 ( .A(n2227), .ZN(n2226) );
  AOI21_X1 U2567 ( .B1(n2227), .B2(n2225), .A(n2224), .ZN(n2223) );
  OAI21_X1 U2568 ( .B1(n3327), .B2(n2951), .A(n3889), .ZN(n3315) );
  INV_X1 U2569 ( .A(n3827), .ZN(n2917) );
  OAI21_X1 U2570 ( .B1(n3618), .B2(n2949), .A(n3880), .ZN(n3221) );
  OR2_X1 U2571 ( .A1(n3613), .A2(n3622), .ZN(n3614) );
  AND2_X1 U2572 ( .A1(n3617), .A2(n2913), .ZN(n2382) );
  AND2_X1 U2573 ( .A1(n2970), .A2(n2969), .ZN(n4547) );
  INV_X1 U2574 ( .A(n2946), .ZN(n3829) );
  INV_X1 U2575 ( .A(n2235), .ZN(n2232) );
  NAND2_X1 U2576 ( .A1(n4479), .A2(n3255), .ZN(n4891) );
  AND2_X1 U2577 ( .A1(n3150), .A2(n3929), .ZN(n4636) );
  AND2_X1 U2578 ( .A1(n2854), .A2(n4687), .ZN(n3038) );
  AND2_X1 U2579 ( .A1(n2407), .A2(n2231), .ZN(n2214) );
  OR2_X1 U2580 ( .A1(n2445), .A2(n2388), .ZN(n2222) );
  NOR2_X1 U2581 ( .A1(n2443), .A2(n2221), .ZN(n2220) );
  CLKBUF_X1 U2582 ( .A(n2425), .Z(n2426) );
  INV_X1 U2583 ( .A(IR_REG_19__SCAN_IN), .ZN(n2464) );
  NAND2_X1 U2584 ( .A1(n3297), .A2(n3296), .ZN(n2312) );
  NAND2_X1 U2585 ( .A1(n3295), .A2(n2313), .ZN(n2308) );
  OR2_X1 U2586 ( .A1(n2839), .A2(n2817), .ZN(n4385) );
  INV_X1 U2587 ( .A(n3229), .ZN(n3241) );
  INV_X1 U2588 ( .A(n2293), .ZN(n2292) );
  OAI21_X1 U2589 ( .B1(n2529), .B2(n2294), .A(n3236), .ZN(n2293) );
  MUX2_X1 U2590 ( .A(n4698), .B(DATAI_2_), .S(n3794), .Z(n3257) );
  NAND2_X1 U2591 ( .A1(n2885), .A2(n4519), .ZN(n3784) );
  NAND2_X1 U2592 ( .A1(n2882), .A2(n3173), .ZN(n3787) );
  NAND2_X1 U2593 ( .A1(n2896), .A2(n2872), .ZN(n3790) );
  INV_X1 U2594 ( .A(n4691), .ZN(n4307) );
  NAND2_X1 U2595 ( .A1(n2829), .A2(n2828), .ZN(n4378) );
  XNOR2_X1 U2596 ( .A(n3066), .B(n4696), .ZN(n4271) );
  XNOR2_X1 U2597 ( .A(n3087), .B(n4694), .ZN(n3088) );
  NAND2_X1 U2598 ( .A1(n4733), .A2(n4734), .ZN(n4732) );
  XNOR2_X1 U2599 ( .A(n3460), .B(n4854), .ZN(n4745) );
  XNOR2_X1 U2600 ( .A(n2274), .B(n4304), .ZN(n4309) );
  NOR2_X1 U2601 ( .A1(n4805), .A2(n2198), .ZN(n2274) );
  AOI21_X1 U2602 ( .B1(n2164), .B2(n2364), .A(n2187), .ZN(n2363) );
  CLKBUF_X1 U2603 ( .A(n3190), .Z(n4557) );
  INV_X1 U2604 ( .A(IR_REG_18__SCAN_IN), .ZN(n2408) );
  INV_X1 U2605 ( .A(IR_REG_17__SCAN_IN), .ZN(n2386) );
  INV_X1 U2606 ( .A(n4347), .ZN(n2968) );
  INV_X1 U2607 ( .A(n2724), .ZN(n2305) );
  INV_X1 U2608 ( .A(n3933), .ZN(n2895) );
  AND2_X1 U2609 ( .A1(n4283), .A2(n4282), .ZN(n4284) );
  INV_X1 U2610 ( .A(n2939), .ZN(n2367) );
  NOR2_X1 U2611 ( .A1(n3920), .A2(n2202), .ZN(n2201) );
  INV_X1 U2612 ( .A(n4340), .ZN(n2202) );
  INV_X1 U2613 ( .A(n3892), .ZN(n2225) );
  INV_X1 U2614 ( .A(n3900), .ZN(n2224) );
  NAND2_X1 U2615 ( .A1(n3880), .A2(n3877), .ZN(n3617) );
  NOR2_X1 U2616 ( .A1(n2992), .A2(n4347), .ZN(n2235) );
  INV_X1 U2617 ( .A(n4365), .ZN(n2991) );
  AND2_X1 U2618 ( .A1(n2238), .A2(n4425), .ZN(n2237) );
  NOR2_X1 U2619 ( .A1(n4445), .A2(n2239), .ZN(n2238) );
  INV_X1 U2620 ( .A(n4459), .ZN(n2239) );
  NOR2_X1 U2621 ( .A1(n3441), .A2(n3435), .ZN(n2230) );
  INV_X1 U2622 ( .A(n3038), .ZN(n2986) );
  NAND2_X1 U2623 ( .A1(n2441), .A2(n2440), .ZN(n2444) );
  NOR2_X1 U2624 ( .A1(IR_REG_29__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2221)
         );
  NOR2_X1 U2625 ( .A1(n2320), .A2(n2170), .ZN(n2315) );
  NOR2_X1 U2626 ( .A1(n3492), .A2(n2321), .ZN(n2320) );
  INV_X1 U2627 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4098) );
  NAND2_X1 U2628 ( .A1(n3388), .A2(n3389), .ZN(n2290) );
  AND2_X1 U2629 ( .A1(n2759), .A2(n2758), .ZN(n3660) );
  INV_X1 U2630 ( .A(n2310), .ZN(n2309) );
  INV_X1 U2631 ( .A(n2312), .ZN(n2311) );
  AND2_X1 U2632 ( .A1(n2880), .A2(n2468), .ZN(n2832) );
  OR2_X1 U2633 ( .A1(n2774), .A2(n4039), .ZN(n2786) );
  OAI22_X1 U2634 ( .A1(n3408), .A2(n3003), .B1(n2792), .B2(n2955), .ZN(n3536)
         );
  INV_X1 U2635 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2661) );
  OR2_X1 U2636 ( .A1(n2662), .A2(n2661), .ZN(n2684) );
  OR2_X1 U2637 ( .A1(n3677), .A2(n3678), .ZN(n2336) );
  AND2_X1 U2638 ( .A1(n2896), .A2(n2895), .ZN(n2899) );
  OAI21_X1 U2639 ( .B1(n2300), .B2(n2299), .A(n2192), .ZN(n2297) );
  INV_X1 U2640 ( .A(n3711), .ZN(n2299) );
  NAND2_X1 U2641 ( .A1(n2725), .A2(n2724), .ZN(n3774) );
  NOR2_X1 U2642 ( .A1(n2725), .A2(n2724), .ZN(n3776) );
  OAI21_X1 U2643 ( .B1(n3035), .B2(n2415), .A(n2414), .ZN(n2417) );
  AND2_X1 U2644 ( .A1(n3184), .A2(n2994), .ZN(n2896) );
  INV_X1 U2645 ( .A(n4689), .ZN(n3862) );
  AND4_X1 U2646 ( .A1(n2716), .A2(n2715), .A3(n2714), .A4(n2713), .ZN(n3779)
         );
  NAND2_X1 U2647 ( .A1(n4699), .A2(REG2_REG_1__SCAN_IN), .ZN(n2284) );
  XNOR2_X1 U2648 ( .A(n3076), .B(n2281), .ZN(n3100) );
  AND2_X1 U2649 ( .A1(n2278), .A2(n4696), .ZN(n2276) );
  AND3_X1 U2650 ( .A1(n2268), .A2(n2191), .A3(n2267), .ZN(n3452) );
  XNOR2_X1 U2651 ( .A(n3469), .B(n3468), .ZN(n4720) );
  NOR2_X1 U2652 ( .A1(n4720), .A2(n2619), .ZN(n4719) );
  NOR2_X1 U2653 ( .A1(n4738), .A2(n3472), .ZN(n3476) );
  OR2_X1 U2654 ( .A1(n3476), .A2(n3475), .ZN(n4283) );
  XNOR2_X1 U2655 ( .A(n4284), .B(n2282), .ZN(n4749) );
  NOR2_X1 U2656 ( .A1(n4764), .A2(n4763), .ZN(n4762) );
  XNOR2_X1 U2657 ( .A(n4287), .B(n2720), .ZN(n4778) );
  NAND2_X1 U2658 ( .A1(n4778), .A2(n4777), .ZN(n4776) );
  NAND2_X1 U2659 ( .A1(n4779), .A2(n4300), .ZN(n4790) );
  AOI21_X1 U2660 ( .B1(n4798), .B2(n2260), .A(n2259), .ZN(n2258) );
  AND2_X1 U2661 ( .A1(n2194), .A2(n4289), .ZN(n2259) );
  AND2_X1 U2662 ( .A1(n2164), .A2(n3835), .ZN(n2362) );
  AND2_X1 U2663 ( .A1(n2368), .A2(n3835), .ZN(n2364) );
  NAND2_X1 U2664 ( .A1(n2200), .A2(n2199), .ZN(n4315) );
  AOI21_X1 U2665 ( .B1(n2201), .B2(n2205), .A(n3799), .ZN(n2199) );
  NAND2_X1 U2666 ( .A1(n4394), .A2(n2201), .ZN(n2200) );
  INV_X1 U2667 ( .A(n4361), .ZN(n3865) );
  AND2_X1 U2668 ( .A1(n4311), .A2(n2888), .ZN(n3634) );
  AND2_X1 U2669 ( .A1(n3794), .A2(DATAI_27_), .ZN(n4347) );
  AND2_X1 U2670 ( .A1(n2203), .A2(n2207), .ZN(n4339) );
  NAND2_X1 U2671 ( .A1(n2203), .A2(n2201), .ZN(n4338) );
  AND2_X1 U2672 ( .A1(n4355), .A2(n3840), .ZN(n4375) );
  AND2_X1 U2673 ( .A1(n2807), .A2(REG3_REG_24__SCAN_IN), .ZN(n2816) );
  OR2_X1 U2674 ( .A1(n2786), .A2(n3745), .ZN(n2796) );
  NOR2_X1 U2675 ( .A1(n2796), .A2(n4135), .ZN(n2807) );
  INV_X1 U2676 ( .A(n3746), .ZN(n4445) );
  AND3_X1 U2677 ( .A1(n2801), .A2(n2800), .A3(n2799), .ZN(n4440) );
  OAI22_X1 U2678 ( .A1(n4489), .A2(n2341), .B1(n2343), .B2(n2395), .ZN(n4433)
         );
  NAND2_X1 U2679 ( .A1(n2345), .A2(n2348), .ZN(n2341) );
  AOI21_X1 U2680 ( .B1(n2344), .B2(n2345), .A(n2186), .ZN(n2343) );
  NAND2_X1 U2681 ( .A1(n4433), .A2(n2934), .ZN(n4432) );
  NAND2_X1 U2682 ( .A1(n2963), .A2(n3811), .ZN(n4452) );
  OAI21_X1 U2683 ( .B1(n3599), .B2(n2218), .A(n2215), .ZN(n2963) );
  AND2_X1 U2684 ( .A1(n2216), .A2(n3907), .ZN(n2215) );
  NAND2_X1 U2685 ( .A1(n2217), .A2(n3591), .ZN(n2216) );
  NAND2_X1 U2686 ( .A1(n3598), .A2(n2217), .ZN(n4469) );
  AND2_X1 U2687 ( .A1(n2347), .A2(n2349), .ZN(n4467) );
  NAND2_X1 U2688 ( .A1(n4489), .A2(n2933), .ZN(n2347) );
  NOR2_X1 U2689 ( .A1(n2739), .A2(n2738), .ZN(n2750) );
  OR2_X1 U2690 ( .A1(n2711), .A2(n4139), .ZN(n2739) );
  AND4_X1 U2691 ( .A1(n2745), .A2(n2744), .A3(n2743), .A4(n2742), .ZN(n4542)
         );
  NAND2_X1 U2692 ( .A1(n3598), .A2(n3802), .ZN(n4540) );
  NAND2_X1 U2693 ( .A1(n3599), .A2(n3842), .ZN(n3598) );
  OR2_X1 U2694 ( .A1(n3567), .A2(n3785), .ZN(n3593) );
  OAI21_X1 U2695 ( .B1(n3548), .B2(n2358), .A(n2357), .ZN(n3592) );
  NAND2_X1 U2696 ( .A1(n2359), .A2(n2165), .ZN(n2357) );
  NAND2_X1 U2697 ( .A1(n2361), .A2(n2165), .ZN(n2358) );
  NAND2_X1 U2698 ( .A1(n3592), .A2(n3591), .ZN(n3590) );
  OR2_X1 U2699 ( .A1(n3561), .A2(n3559), .ZN(n3562) );
  AND4_X1 U2700 ( .A1(n2651), .A2(n2650), .A3(n2649), .A4(n2648), .ZN(n3539)
         );
  AND2_X1 U2701 ( .A1(n2380), .A2(n2378), .ZN(n2377) );
  INV_X1 U2702 ( .A(n3823), .ZN(n2378) );
  INV_X1 U2703 ( .A(n3364), .ZN(n3437) );
  AND4_X1 U2704 ( .A1(n2643), .A2(n2642), .A3(n2641), .A4(n2640), .ZN(n3409)
         );
  OR2_X1 U2705 ( .A1(n2620), .A2(n4036), .ZN(n2637) );
  NAND2_X1 U2706 ( .A1(n3315), .A2(n3893), .ZN(n2952) );
  INV_X1 U2707 ( .A(n2915), .ZN(n2351) );
  INV_X1 U2708 ( .A(n2353), .ZN(n2352) );
  AND4_X1 U2709 ( .A1(n2587), .A2(n2586), .A3(n2585), .A4(n2584), .ZN(n3390)
         );
  AND2_X1 U2710 ( .A1(n3887), .A2(n3889), .ZN(n3827) );
  NAND2_X1 U2711 ( .A1(n2950), .A2(n3886), .ZN(n3327) );
  AND4_X1 U2712 ( .A1(n2577), .A2(n2576), .A3(n2575), .A4(n2574), .ZN(n3300)
         );
  AOI21_X1 U2713 ( .B1(n3221), .B2(n3884), .A(n3220), .ZN(n3267) );
  OR2_X1 U2714 ( .A1(n2971), .A2(n4701), .ZN(n4528) );
  AND2_X1 U2715 ( .A1(n4701), .A2(n3045), .ZN(n4525) );
  NAND2_X1 U2716 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2551) );
  NAND2_X1 U2717 ( .A1(n2948), .A2(n3876), .ZN(n3618) );
  INV_X1 U2718 ( .A(n3617), .ZN(n3828) );
  INV_X1 U2719 ( .A(n2947), .ZN(n3214) );
  NAND2_X1 U2720 ( .A1(n3150), .A2(n4690), .ZN(n4565) );
  NOR2_X1 U2721 ( .A1(n4364), .A2(n4347), .ZN(n4346) );
  OR2_X1 U2722 ( .A1(n4384), .A2(n2991), .ZN(n4364) );
  NAND2_X1 U2723 ( .A1(n4401), .A2(n4382), .ZN(n4384) );
  AND2_X1 U2724 ( .A1(n4483), .A2(n2236), .ZN(n4401) );
  AND2_X1 U2725 ( .A1(n2237), .A2(n4403), .ZN(n2236) );
  NAND2_X1 U2726 ( .A1(n4483), .A2(n2237), .ZN(n4424) );
  NAND2_X1 U2727 ( .A1(n4483), .A2(n2238), .ZN(n4606) );
  NAND2_X1 U2728 ( .A1(n4483), .A2(n4459), .ZN(n4461) );
  AND2_X1 U2729 ( .A1(n4504), .A2(n4481), .ZN(n4483) );
  OR2_X1 U2730 ( .A1(n4552), .A2(n4524), .ZN(n4503) );
  NOR2_X1 U2731 ( .A1(n4503), .A2(n3665), .ZN(n4504) );
  NOR2_X1 U2732 ( .A1(n3593), .A2(n3594), .ZN(n4550) );
  INV_X1 U2733 ( .A(n4891), .ZN(n4638) );
  NAND2_X1 U2734 ( .A1(n3553), .A2(n3585), .ZN(n3567) );
  NOR2_X1 U2735 ( .A1(n3528), .A2(n3542), .ZN(n3553) );
  NAND2_X1 U2736 ( .A1(n2230), .A2(n3499), .ZN(n3528) );
  INV_X1 U2737 ( .A(n2230), .ZN(n3442) );
  AND2_X1 U2738 ( .A1(n3228), .A2(n2189), .ZN(n3383) );
  NAND2_X1 U2739 ( .A1(n3383), .A2(n3483), .ZN(n3441) );
  NAND2_X1 U2740 ( .A1(n3228), .A2(n2160), .ZN(n3334) );
  NAND2_X1 U2741 ( .A1(n3228), .A2(n2355), .ZN(n3333) );
  INV_X1 U2742 ( .A(n2994), .ZN(n3185) );
  NAND2_X1 U2743 ( .A1(n2454), .A2(n4843), .ZN(n3182) );
  INV_X1 U2744 ( .A(IR_REG_27__SCAN_IN), .ZN(n3034) );
  NAND2_X1 U2745 ( .A1(n2208), .A2(n2429), .ZN(n2866) );
  AND2_X1 U2746 ( .A1(n2561), .A2(n2413), .ZN(n2427) );
  NAND2_X1 U2747 ( .A1(n2460), .A2(n2459), .ZN(n2941) );
  NOR2_X1 U2748 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2420)
         );
  NOR2_X1 U2749 ( .A1(n2732), .A2(IR_REG_17__SCAN_IN), .ZN(n2746) );
  AND2_X1 U2750 ( .A1(n2717), .A2(n2709), .ZN(n4298) );
  AND2_X1 U2751 ( .A1(n2611), .A2(n2672), .ZN(n3467) );
  OR2_X1 U2752 ( .A1(n2565), .A2(n2578), .ZN(n3080) );
  AND2_X1 U2753 ( .A1(n2190), .A2(n2333), .ZN(n2332) );
  INV_X1 U2754 ( .A(n3377), .ZN(n3483) );
  CLKBUF_X1 U2755 ( .A(n3169), .Z(n3170) );
  XNOR2_X1 U2756 ( .A(n2515), .B(n2514), .ZN(n3211) );
  NAND2_X1 U2757 ( .A1(n3794), .A2(DATAI_1_), .ZN(n2475) );
  INV_X1 U2758 ( .A(REG3_REG_21__SCAN_IN), .ZN(n4039) );
  NAND2_X1 U2759 ( .A1(n2324), .A2(n2323), .ZN(n3496) );
  OAI21_X1 U2760 ( .B1(n3794), .B2(n2419), .A(n2418), .ZN(n3645) );
  NAND2_X1 U2761 ( .A1(n3794), .A2(DATAI_0_), .ZN(n2418) );
  NAND2_X1 U2762 ( .A1(n3794), .A2(DATAI_20_), .ZN(n4481) );
  NAND2_X1 U2763 ( .A1(n2324), .A2(n2318), .ZN(n2317) );
  NOR2_X1 U2764 ( .A1(n2319), .A2(n3493), .ZN(n2318) );
  INV_X1 U2765 ( .A(n2323), .ZN(n2319) );
  INV_X1 U2766 ( .A(n2955), .ZN(n3542) );
  AND2_X1 U2767 ( .A1(n2336), .A2(n2334), .ZN(n3742) );
  NAND2_X1 U2768 ( .A1(n2336), .A2(n3679), .ZN(n3743) );
  INV_X1 U2769 ( .A(n3780), .ZN(n3703) );
  INV_X1 U2770 ( .A(n3781), .ZN(n3725) );
  AND4_X1 U2771 ( .A1(n2731), .A2(n2730), .A3(n2729), .A4(n2728), .ZN(n4529)
         );
  INV_X1 U2772 ( .A(n3784), .ZN(n3769) );
  NAND2_X1 U2773 ( .A1(n3794), .A2(DATAI_26_), .ZN(n4365) );
  OAI211_X1 U2774 ( .C1(n4385), .C2(n2972), .A(n2819), .B(n2818), .ZN(n4398)
         );
  INV_X1 U2775 ( .A(n4440), .ZN(n3724) );
  INV_X1 U2776 ( .A(n4498), .ZN(n4455) );
  INV_X1 U2777 ( .A(n4542), .ZN(n3939) );
  INV_X1 U2778 ( .A(n4529), .ZN(n3940) );
  INV_X1 U2779 ( .A(n3408), .ZN(n3583) );
  INV_X1 U2780 ( .A(n3539), .ZN(n4235) );
  INV_X1 U2781 ( .A(n3300), .ZN(n4236) );
  OR2_X1 U2782 ( .A1(n2484), .A2(n2498), .ZN(n2503) );
  OR2_X1 U2783 ( .A1(n2484), .A2(n2455), .ZN(n2452) );
  OR2_X1 U2784 ( .A1(n2454), .A2(n3024), .ZN(n4240) );
  OAI21_X1 U2785 ( .B1(n4271), .B2(n3065), .A(n3067), .ZN(n3128) );
  AND2_X1 U2786 ( .A1(n2269), .A2(n2272), .ZN(n3160) );
  NAND2_X1 U2787 ( .A1(n2268), .A2(n2267), .ZN(n3158) );
  NAND2_X1 U2788 ( .A1(n3088), .A2(REG2_REG_6__SCAN_IN), .ZN(n2269) );
  NAND2_X1 U2789 ( .A1(n2241), .A2(n2248), .ZN(n3464) );
  NAND2_X1 U2790 ( .A1(n2246), .A2(n2243), .ZN(n2242) );
  NOR2_X1 U2791 ( .A1(n2247), .A2(n2583), .ZN(n2246) );
  NAND2_X1 U2792 ( .A1(n2253), .A2(n2159), .ZN(n2249) );
  OAI21_X1 U2793 ( .B1(n4720), .B2(n2265), .A(n2264), .ZN(n4728) );
  NAND2_X1 U2794 ( .A1(n2266), .A2(REG1_REG_10__SCAN_IN), .ZN(n2265) );
  NAND2_X1 U2795 ( .A1(n3470), .A2(n2266), .ZN(n2264) );
  INV_X1 U2796 ( .A(n4729), .ZN(n2266) );
  NAND2_X1 U2797 ( .A1(n4724), .A2(n3457), .ZN(n4733) );
  NAND2_X1 U2798 ( .A1(n4744), .A2(n3461), .ZN(n4294) );
  XNOR2_X1 U2799 ( .A(n4295), .B(n2282), .ZN(n4753) );
  NOR2_X1 U2800 ( .A1(n4753), .A2(n4754), .ZN(n4752) );
  NAND2_X1 U2801 ( .A1(n2262), .A2(n2258), .ZN(n2257) );
  OR2_X1 U2802 ( .A1(n4798), .A2(n2263), .ZN(n2262) );
  INV_X1 U2803 ( .A(n4289), .ZN(n2263) );
  OAI21_X1 U2804 ( .B1(n4372), .B2(n2368), .A(n2164), .ZN(n4328) );
  NAND2_X1 U2805 ( .A1(n2373), .A2(n2372), .ZN(n2376) );
  NAND2_X1 U2806 ( .A1(n2342), .A2(n2345), .ZN(n4450) );
  NAND2_X1 U2807 ( .A1(n4489), .A2(n2346), .ZN(n2342) );
  NAND2_X1 U2808 ( .A1(n3547), .A2(n2361), .ZN(n3560) );
  OAI21_X1 U2809 ( .B1(n3368), .B2(n2179), .A(n2923), .ZN(n3382) );
  NAND2_X1 U2810 ( .A1(n2354), .A2(n2916), .ZN(n3274) );
  NAND2_X1 U2811 ( .A1(n3225), .A2(n2915), .ZN(n2354) );
  AND2_X1 U2812 ( .A1(n3190), .A2(n3227), .ZN(n4331) );
  AND2_X1 U2813 ( .A1(n4535), .A2(n4636), .ZN(n4817) );
  INV_X1 U2814 ( .A(n4817), .ZN(n4555) );
  AND2_X1 U2815 ( .A1(n4557), .A2(n3192), .ZN(n4828) );
  INV_X1 U2816 ( .A(n4519), .ZN(n4826) );
  AND2_X2 U2817 ( .A1(n2995), .A2(n2994), .ZN(n4910) );
  INV_X1 U2818 ( .A(n4910), .ZN(n4908) );
  AOI21_X1 U2819 ( .B1(n4636), .B2(n4582), .A(n4581), .ZN(n4583) );
  AND2_X2 U2820 ( .A1(n3185), .A2(n2995), .ZN(n4902) );
  OR2_X1 U2821 ( .A1(n3038), .A2(n3182), .ZN(n4842) );
  AND2_X1 U2822 ( .A1(n2177), .A2(n2413), .ZN(n2387) );
  NAND2_X1 U2823 ( .A1(n2433), .A2(n2432), .ZN(n3026) );
  AND2_X1 U2824 ( .A1(n3044), .A2(STATE_REG_SCAN_IN), .ZN(n4843) );
  INV_X1 U2825 ( .A(n2941), .ZN(n4688) );
  AND2_X1 U2826 ( .A1(n2467), .A2(n2466), .ZN(n4691) );
  INV_X1 U2827 ( .A(n3467), .ZN(n4860) );
  XNOR2_X1 U2828 ( .A(n2589), .B(IR_REG_7__SCAN_IN), .ZN(n4693) );
  INV_X1 U2829 ( .A(n2539), .ZN(n2254) );
  NAND3_X1 U2830 ( .A1(n2287), .A2(n2285), .A3(n2286), .ZN(n4699) );
  NAND3_X1 U2831 ( .A1(n2288), .A2(IR_REG_31__SCAN_IN), .A3(IR_REG_0__SCAN_IN), 
        .ZN(n2286) );
  NAND2_X1 U2832 ( .A1(n2419), .A2(IR_REG_1__SCAN_IN), .ZN(n2285) );
  NAND2_X1 U2833 ( .A1(n2561), .A2(IR_REG_1__SCAN_IN), .ZN(n2287) );
  NAND2_X1 U2834 ( .A1(n2308), .A2(n2312), .ZN(n3308) );
  NAND2_X1 U2835 ( .A1(n3281), .A2(n2532), .ZN(n3237) );
  AOI21_X1 U2836 ( .B1(n4804), .B2(n2168), .A(n4803), .ZN(n4811) );
  NAND2_X1 U2837 ( .A1(n4794), .A2(n2257), .ZN(n2256) );
  NAND2_X1 U2838 ( .A1(n3280), .A2(n2529), .ZN(n3281) );
  OAI21_X1 U2839 ( .B1(n3794), .B2(n2476), .A(n2475), .ZN(n2904) );
  AND2_X1 U2840 ( .A1(n3096), .A2(n2252), .ZN(n2159) );
  INV_X1 U2841 ( .A(n3303), .ZN(n2355) );
  AND2_X1 U2842 ( .A1(n2355), .A2(n3326), .ZN(n2160) );
  AND2_X1 U2843 ( .A1(n2160), .A2(n3351), .ZN(n2161) );
  AND2_X1 U2844 ( .A1(n2356), .A2(n2355), .ZN(n2162) );
  NOR2_X1 U2845 ( .A1(n3437), .A2(n3483), .ZN(n2163) );
  AND2_X1 U2846 ( .A1(n2366), .A2(n2369), .ZN(n2164) );
  OR2_X1 U2847 ( .A1(n3941), .A2(n3785), .ZN(n2165) );
  NAND2_X1 U2848 ( .A1(n4398), .A2(n4377), .ZN(n2166) );
  NAND2_X1 U2849 ( .A1(n4455), .A2(n4472), .ZN(n2167) );
  INV_X1 U2850 ( .A(n2927), .ZN(n3585) );
  NAND2_X1 U2851 ( .A1(n2188), .A2(n2167), .ZN(n2345) );
  NOR2_X1 U2852 ( .A1(n3665), .A2(n4526), .ZN(n2932) );
  NAND2_X1 U2853 ( .A1(n2517), .A2(n2518), .ZN(n3280) );
  AND2_X1 U2854 ( .A1(n3078), .A2(n4318), .ZN(n4794) );
  INV_X1 U2855 ( .A(n2477), .ZN(n2847) );
  INV_X2 U2856 ( .A(n2749), .ZN(n2846) );
  OR2_X1 U2857 ( .A1(n4799), .A2(n4798), .ZN(n2168) );
  NAND2_X1 U2858 ( .A1(n2222), .A2(n2220), .ZN(n2447) );
  AND2_X1 U2859 ( .A1(n2408), .A2(n2386), .ZN(n2169) );
  AND2_X1 U2860 ( .A1(n3405), .A2(n3407), .ZN(n3823) );
  AND4_X1 U2861 ( .A1(n2474), .A2(n2473), .A3(n2472), .A4(n2471), .ZN(n2905)
         );
  NAND2_X1 U2862 ( .A1(n2446), .A2(n3031), .ZN(n2484) );
  INV_X1 U2863 ( .A(IR_REG_3__SCAN_IN), .ZN(n2505) );
  AND2_X1 U2864 ( .A1(n2539), .A2(n2400), .ZN(n2559) );
  AND2_X1 U2865 ( .A1(n2526), .A2(n2507), .ZN(n4697) );
  INV_X1 U2866 ( .A(n4697), .ZN(n2281) );
  AND3_X1 U2867 ( .A1(n2322), .A2(n2323), .A3(n3535), .ZN(n2170) );
  AND2_X1 U2868 ( .A1(n2447), .A2(n4686), .ZN(n2171) );
  INV_X1 U2869 ( .A(n3920), .ZN(n2207) );
  NAND2_X1 U2870 ( .A1(n3645), .A2(n2847), .ZN(n2172) );
  AND2_X1 U2871 ( .A1(n2630), .A2(n2618), .ZN(n2173) );
  AND2_X1 U2872 ( .A1(n2582), .A2(n2581), .ZN(n2174) );
  INV_X1 U2873 ( .A(n2406), .ZN(n2407) );
  INV_X1 U2874 ( .A(n2389), .ZN(n2443) );
  NAND2_X1 U2875 ( .A1(n2331), .A2(n2332), .ZN(n2338) );
  INV_X1 U2876 ( .A(n2204), .ZN(n4373) );
  OR2_X1 U2877 ( .A1(n4394), .A2(n3916), .ZN(n2204) );
  NAND2_X1 U2878 ( .A1(n3331), .A2(n3303), .ZN(n2175) );
  OR2_X1 U2879 ( .A1(n3364), .A2(n3377), .ZN(n2176) );
  AND2_X1 U2880 ( .A1(n2440), .A2(n2388), .ZN(n2177) );
  NOR2_X1 U2881 ( .A1(n2320), .A2(n2316), .ZN(n2178) );
  AND2_X1 U2882 ( .A1(n3481), .A2(n3392), .ZN(n2179) );
  INV_X1 U2883 ( .A(n2532), .ZN(n2294) );
  NAND2_X1 U2884 ( .A1(n2385), .A2(n2169), .ZN(n2435) );
  INV_X1 U2885 ( .A(IR_REG_21__SCAN_IN), .ZN(n2329) );
  INV_X1 U2886 ( .A(n3331), .ZN(n2356) );
  INV_X1 U2887 ( .A(n3535), .ZN(n2321) );
  OAI21_X1 U2888 ( .B1(n3756), .B2(n2762), .A(n2761), .ZN(n3681) );
  OR3_X1 U2889 ( .A1(n4384), .A2(n2991), .A3(n2232), .ZN(n2180) );
  INV_X1 U2890 ( .A(n2609), .ZN(n2212) );
  AND2_X1 U2891 ( .A1(n3583), .A2(n3542), .ZN(n2181) );
  NOR2_X1 U2892 ( .A1(n3865), .A2(n2968), .ZN(n2182) );
  AOI21_X1 U2893 ( .B1(n3420), .B2(n2392), .A(n2925), .ZN(n3516) );
  NOR2_X1 U2894 ( .A1(n4312), .A2(n4313), .ZN(n4327) );
  AND2_X1 U2895 ( .A1(n4498), .A2(n4481), .ZN(n2183) );
  OR2_X1 U2896 ( .A1(n4378), .A2(n2991), .ZN(n2184) );
  NAND2_X1 U2897 ( .A1(n2379), .A2(n2380), .ZN(n3433) );
  INV_X1 U2898 ( .A(n3351), .ZN(n2990) );
  MUX2_X1 U2899 ( .A(n4692), .B(n2593), .S(n3794), .Z(n3351) );
  AND2_X1 U2900 ( .A1(n4378), .A2(n2991), .ZN(n2185) );
  INV_X1 U2901 ( .A(IR_REG_4__SCAN_IN), .ZN(n2398) );
  INV_X1 U2902 ( .A(n3392), .ZN(n3369) );
  NOR2_X1 U2903 ( .A1(n3747), .A2(n4459), .ZN(n2186) );
  NOR2_X1 U2904 ( .A1(n4326), .A2(n4325), .ZN(n2187) );
  INV_X1 U2905 ( .A(n2395), .ZN(n2348) );
  INV_X1 U2906 ( .A(n2218), .ZN(n2217) );
  NAND2_X1 U2907 ( .A1(n2219), .A2(n3802), .ZN(n2218) );
  INV_X1 U2908 ( .A(n3782), .ZN(n3942) );
  AND4_X1 U2909 ( .A1(n2689), .A2(n2688), .A3(n2687), .A4(n2686), .ZN(n3782)
         );
  OAI21_X1 U2910 ( .B1(n3549), .B2(n2360), .A(n2928), .ZN(n2359) );
  INV_X1 U2911 ( .A(n2361), .ZN(n2360) );
  NAND2_X1 U2912 ( .A1(n3782), .A2(n3585), .ZN(n2361) );
  OR2_X1 U2913 ( .A1(n2932), .A2(n2183), .ZN(n2188) );
  AND2_X1 U2914 ( .A1(n2161), .A2(n3369), .ZN(n2189) );
  AND2_X1 U2915 ( .A1(n2340), .A2(n2339), .ZN(n2190) );
  INV_X1 U2916 ( .A(IR_REG_29__SCAN_IN), .ZN(n2388) );
  NAND2_X1 U2917 ( .A1(n4693), .A2(REG2_REG_7__SCAN_IN), .ZN(n2191) );
  INV_X1 U2918 ( .A(n2166), .ZN(n2374) );
  INV_X1 U2919 ( .A(n4757), .ZN(n2282) );
  NAND2_X1 U2920 ( .A1(n2922), .A2(n2921), .ZN(n3368) );
  NAND2_X1 U2921 ( .A1(n2307), .A2(n2306), .ZN(n3344) );
  INV_X1 U2922 ( .A(n3897), .ZN(n2228) );
  OR2_X1 U2923 ( .A1(n2736), .A2(n2735), .ZN(n2192) );
  NAND2_X1 U2924 ( .A1(n2290), .A2(n2618), .ZN(n3484) );
  NAND2_X1 U2925 ( .A1(n2909), .A2(n2946), .ZN(n3246) );
  INV_X1 U2926 ( .A(n2385), .ZN(n2732) );
  NAND2_X1 U2927 ( .A1(n2383), .A2(n2913), .ZN(n3620) );
  NOR2_X1 U2928 ( .A1(n4719), .A2(n3470), .ZN(n2193) );
  NAND2_X1 U2929 ( .A1(n3228), .A2(n2161), .ZN(n2229) );
  AND2_X1 U2930 ( .A1(n2965), .A2(n2964), .ZN(n4434) );
  INV_X1 U2931 ( .A(n4434), .ZN(n2934) );
  INV_X1 U2932 ( .A(n2932), .ZN(n2349) );
  XNOR2_X1 U2933 ( .A(n2719), .B(n2718), .ZN(n4850) );
  AND2_X1 U2934 ( .A1(n4302), .A2(REG1_REG_18__SCAN_IN), .ZN(n2194) );
  AND3_X1 U2935 ( .A1(n2249), .A2(n2248), .A3(n2250), .ZN(n2195) );
  INV_X1 U2936 ( .A(n2261), .ZN(n2260) );
  OR2_X1 U2937 ( .A1(n2194), .A2(n4289), .ZN(n2261) );
  NAND2_X1 U2938 ( .A1(n2258), .A2(n2261), .ZN(n2196) );
  AND2_X1 U2939 ( .A1(n3794), .A2(DATAI_23_), .ZN(n4419) );
  INV_X1 U2940 ( .A(n4419), .ZN(n4425) );
  INV_X1 U2941 ( .A(n4403), .ZN(n3726) );
  NAND2_X1 U2942 ( .A1(n3794), .A2(DATAI_24_), .ZN(n4403) );
  AND2_X1 U2943 ( .A1(n4794), .A2(n2196), .ZN(n2197) );
  INV_X1 U2944 ( .A(n4692), .ZN(n2252) );
  INV_X1 U2945 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2271) );
  INV_X1 U2946 ( .A(IR_REG_25__SCAN_IN), .ZN(n2231) );
  AND2_X1 U2947 ( .A1(n4302), .A2(REG2_REG_18__SCAN_IN), .ZN(n2198) );
  INV_X1 U2948 ( .A(IR_REG_28__SCAN_IN), .ZN(n2415) );
  NAND2_X1 U2949 ( .A1(n2213), .A2(n2564), .ZN(n2609) );
  AND2_X1 U2950 ( .A1(n2412), .A2(n2169), .ZN(n2384) );
  NAND4_X1 U2951 ( .A1(n2209), .A2(n2407), .A3(n2211), .A4(n2213), .ZN(n2208)
         );
  OAI21_X1 U2952 ( .B1(n3363), .B2(n2226), .A(n2223), .ZN(n3431) );
  OAI21_X1 U2953 ( .B1(n3363), .B2(n3362), .A(n3892), .ZN(n3376) );
  AOI21_X1 U2954 ( .B1(n3362), .B2(n3892), .A(n2228), .ZN(n2227) );
  AND2_X2 U2955 ( .A1(n2419), .A2(n2288), .ZN(n2539) );
  INV_X1 U2956 ( .A(n2229), .ZN(n3370) );
  NAND3_X1 U2957 ( .A1(n2407), .A2(n2212), .A3(n2384), .ZN(n2430) );
  AOI21_X1 U2958 ( .B1(n3155), .B2(n2159), .A(n2242), .ZN(n2241) );
  NAND2_X1 U2959 ( .A1(n2253), .A2(n3096), .ZN(n3465) );
  NAND2_X1 U2960 ( .A1(n2254), .A2(IR_REG_31__SCAN_IN), .ZN(n2490) );
  NAND2_X1 U2961 ( .A1(n4799), .A2(n2197), .ZN(n2255) );
  OAI211_X1 U2962 ( .C1(n4799), .C2(n2256), .A(n2255), .B(n4310), .ZN(U3259)
         );
  NOR2_X1 U2963 ( .A1(n4711), .A2(n4710), .ZN(n4709) );
  NOR2_X1 U2964 ( .A1(n4740), .A2(n4739), .ZN(n4738) );
  NOR2_X1 U2965 ( .A1(n4285), .A2(n4748), .ZN(n4764) );
  NAND2_X1 U2966 ( .A1(n4550), .A2(n4549), .ZN(n4552) );
  NAND2_X1 U2967 ( .A1(n2273), .A2(n4694), .ZN(n2272) );
  INV_X1 U2968 ( .A(n3087), .ZN(n2273) );
  INV_X1 U2969 ( .A(IR_REG_1__SCAN_IN), .ZN(n2288) );
  OAI21_X1 U2970 ( .B1(n4699), .B2(REG2_REG_1__SCAN_IN), .A(n2284), .ZN(n3072)
         );
  NAND3_X1 U2971 ( .A1(n2517), .A2(n2532), .A3(n2518), .ZN(n2291) );
  NAND2_X1 U2972 ( .A1(n2292), .A2(n2291), .ZN(n3235) );
  OR2_X4 U2973 ( .A1(n2477), .A2(n4636), .ZN(n3003) );
  AND2_X1 U2974 ( .A1(n2296), .A2(n2295), .ZN(n2514) );
  NAND2_X1 U2975 ( .A1(n4238), .A2(n2558), .ZN(n2295) );
  OAI21_X1 U2976 ( .B1(n2725), .B2(n2302), .A(n2300), .ZN(n3710) );
  NOR2_X2 U2977 ( .A1(n2298), .A2(n2297), .ZN(n3756) );
  NOR3_X2 U2978 ( .A1(n2725), .A2(n2302), .A3(n2299), .ZN(n2298) );
  NAND2_X1 U2979 ( .A1(n3295), .A2(n2309), .ZN(n2307) );
  NAND2_X1 U2980 ( .A1(n3423), .A2(n2325), .ZN(n2324) );
  INV_X1 U2981 ( .A(n2314), .ZN(n2680) );
  AOI21_X1 U2982 ( .B1(n3423), .B2(n2178), .A(n2315), .ZN(n2314) );
  NAND2_X1 U2983 ( .A1(n2421), .A2(n2420), .ZN(n2438) );
  INV_X1 U2984 ( .A(n2330), .ZN(n2457) );
  NAND2_X1 U2985 ( .A1(n2330), .A2(IR_REG_31__SCAN_IN), .ZN(n2458) );
  NAND2_X1 U2986 ( .A1(n3677), .A2(n2334), .ZN(n2331) );
  INV_X1 U2987 ( .A(n2338), .ZN(n3648) );
  NOR2_X1 U2988 ( .A1(n2814), .A2(n2815), .ZN(n2337) );
  INV_X1 U2989 ( .A(n3649), .ZN(n2340) );
  OAI21_X1 U2990 ( .B1(n3225), .B2(n2353), .A(n2350), .ZN(n3341) );
  INV_X1 U2991 ( .A(n3341), .ZN(n2918) );
  NAND2_X1 U2992 ( .A1(n4372), .A2(n2362), .ZN(n2365) );
  NAND2_X1 U2993 ( .A1(n4372), .A2(n2939), .ZN(n2373) );
  NAND2_X1 U2994 ( .A1(n2365), .A2(n2363), .ZN(n4330) );
  AND2_X1 U2995 ( .A1(n2373), .A2(n2166), .ZN(n4353) );
  NAND2_X1 U2996 ( .A1(n2379), .A2(n2377), .ZN(n3432) );
  NAND2_X1 U2997 ( .A1(n2383), .A2(n2382), .ZN(n3619) );
  NAND2_X1 U2998 ( .A1(n2425), .A2(n2387), .ZN(n2389) );
  AOI21_X2 U2999 ( .B1(n2697), .B2(n2696), .A(n2394), .ZN(n2725) );
  OR2_X1 U3000 ( .A1(n2484), .A2(n3057), .ZN(n2472) );
  INV_X1 U3001 ( .A(n2908), .ZN(n3672) );
  XNOR2_X1 U3002 ( .A(n4328), .B(n4327), .ZN(n3640) );
  OR2_X1 U3003 ( .A1(n3636), .A2(n4682), .ZN(n2390) );
  OR2_X1 U3004 ( .A1(n3636), .A2(n4629), .ZN(n2391) );
  NAND2_X1 U3005 ( .A1(n2459), .A2(IR_REG_31__SCAN_IN), .ZN(n2869) );
  AND4_X1 U3006 ( .A1(n2755), .A2(n2754), .A3(n2753), .A4(n2752), .ZN(n4475)
         );
  NAND4_X1 U3007 ( .A1(n2779), .A2(n2778), .A3(n2777), .A4(n2776), .ZN(n4473)
         );
  INV_X1 U3008 ( .A(n4473), .ZN(n3747) );
  AND4_X1 U3009 ( .A1(n2704), .A2(n2703), .A3(n2702), .A4(n2701), .ZN(n3603)
         );
  INV_X1 U3010 ( .A(n3603), .ZN(n3941) );
  OR2_X1 U3011 ( .A1(n3539), .A2(n3499), .ZN(n2392) );
  INV_X1 U3012 ( .A(n3785), .ZN(n3566) );
  AND3_X1 U3013 ( .A1(n3010), .A2(n3011), .A3(n3757), .ZN(n2393) );
  AND2_X1 U3014 ( .A1(n2695), .A2(n2694), .ZN(n2394) );
  AND2_X1 U3015 ( .A1(n3747), .A2(n4459), .ZN(n2395) );
  OR2_X1 U3016 ( .A1(n3779), .A2(n3705), .ZN(n2396) );
  INV_X1 U3017 ( .A(n3665), .ZN(n4506) );
  NAND2_X1 U3018 ( .A1(n3794), .A2(DATAI_21_), .ZN(n4459) );
  INV_X1 U3019 ( .A(n4699), .ZN(n2476) );
  INV_X2 U3020 ( .A(IR_REG_0__SCAN_IN), .ZN(n2419) );
  INV_X1 U3021 ( .A(IR_REG_24__SCAN_IN), .ZN(n2409) );
  NAND2_X1 U3022 ( .A1(n2464), .A2(n2870), .ZN(n2410) );
  AND2_X1 U3023 ( .A1(n3754), .A2(n3753), .ZN(n2757) );
  AND2_X1 U3024 ( .A1(n4468), .A2(n2962), .ZN(n3907) );
  INV_X1 U3025 ( .A(IR_REG_26__SCAN_IN), .ZN(n2413) );
  INV_X1 U3026 ( .A(n3487), .ZN(n2630) );
  INV_X1 U3027 ( .A(n3191), .ZN(n2468) );
  OR2_X1 U3028 ( .A1(n2484), .A2(n3261), .ZN(n2485) );
  NAND2_X1 U3029 ( .A1(n2908), .A2(n3257), .ZN(n3871) );
  NAND2_X1 U3030 ( .A1(n3235), .A2(n2547), .ZN(n3295) );
  INV_X1 U3031 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4036) );
  INV_X1 U3032 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2636) );
  INV_X1 U3033 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4139) );
  OR2_X1 U3034 ( .A1(n4427), .A2(n2972), .ZN(n2801) );
  AND2_X1 U3035 ( .A1(n2483), .A2(REG3_REG_2__SCAN_IN), .ZN(n2489) );
  INV_X1 U3036 ( .A(n4857), .ZN(n3468) );
  AND2_X1 U3037 ( .A1(n3794), .A2(DATAI_28_), .ZN(n2992) );
  INV_X1 U3038 ( .A(n3516), .ZN(n3517) );
  INV_X1 U3039 ( .A(n2992), .ZN(n4325) );
  INV_X1 U3040 ( .A(n3435), .ZN(n3443) );
  NOR2_X1 U3041 ( .A1(n2684), .A2(n4098), .ZN(n2698) );
  NAND2_X1 U3042 ( .A1(n2571), .A2(REG3_REG_7__SCAN_IN), .ZN(n2603) );
  INV_X1 U3043 ( .A(n3594), .ZN(n3705) );
  OR2_X1 U3044 ( .A1(n2603), .A2(n2602), .ZN(n2620) );
  NAND2_X1 U3045 ( .A1(n2763), .A2(REG3_REG_20__SCAN_IN), .ZN(n2774) );
  NAND2_X1 U3046 ( .A1(n3794), .A2(DATAI_22_), .ZN(n3746) );
  NAND2_X1 U3047 ( .A1(n2899), .A2(n4250), .ZN(n3781) );
  AND2_X1 U3048 ( .A1(n2894), .A2(n2893), .ZN(n4326) );
  AND4_X1 U3049 ( .A1(n2667), .A2(n2666), .A3(n2665), .A4(n2664), .ZN(n3408)
         );
  AND2_X1 U3050 ( .A1(n3794), .A2(n3046), .ZN(n3048) );
  AND2_X1 U3051 ( .A1(n3049), .A2(n3048), .ZN(n3078) );
  AND2_X1 U3052 ( .A1(n3839), .A2(n3838), .ZN(n4358) );
  INV_X1 U3053 ( .A(n4454), .ZN(n4423) );
  OR2_X1 U3054 ( .A1(n3182), .A2(n2884), .ZN(n4519) );
  OR2_X1 U3055 ( .A1(n2986), .A2(D_REG_0__SCAN_IN), .ZN(n2868) );
  NAND2_X1 U3056 ( .A1(n3794), .A2(DATAI_25_), .ZN(n4382) );
  INV_X1 U3057 ( .A(n3499), .ZN(n3414) );
  INV_X1 U3058 ( .A(n4525), .ZN(n4541) );
  AND2_X1 U3059 ( .A1(n2816), .A2(REG3_REG_25__SCAN_IN), .ZN(n2839) );
  NOR2_X1 U3060 ( .A1(n2551), .A2(n2550), .ZN(n2571) );
  OR3_X1 U3061 ( .A1(n2792), .A2(n3024), .A3(n2880), .ZN(n3933) );
  OR2_X1 U3062 ( .A1(n2873), .A2(n2972), .ZN(n2845) );
  AND4_X1 U3063 ( .A1(n2768), .A2(n2767), .A3(n2766), .A4(n2765), .ZN(n4498)
         );
  NAND2_X1 U3064 ( .A1(n4802), .A2(n4801), .ZN(n4803) );
  INV_X1 U3065 ( .A(n4565), .ZN(n4576) );
  INV_X1 U3066 ( .A(n4528), .ZN(n4545) );
  INV_X1 U3067 ( .A(n4547), .ZN(n4531) );
  INV_X1 U3068 ( .A(n3645), .ZN(n3152) );
  AND2_X1 U3069 ( .A1(n2868), .A2(n3039), .ZN(n2994) );
  AND2_X1 U3070 ( .A1(n2988), .A2(n2987), .ZN(n2995) );
  OR2_X1 U3071 ( .A1(n2578), .A2(n2561), .ZN(n2589) );
  OR2_X1 U3072 ( .A1(n3021), .A2(n3006), .ZN(n3023) );
  NAND2_X1 U3073 ( .A1(n2899), .A2(n4701), .ZN(n3780) );
  INV_X1 U3074 ( .A(n3787), .ZN(n3762) );
  NAND2_X1 U3075 ( .A1(n2845), .A2(n2844), .ZN(n4361) );
  OAI211_X1 U3076 ( .C1(n4405), .C2(n2972), .A(n2810), .B(n2809), .ZN(n4420)
         );
  INV_X1 U3077 ( .A(n4475), .ZN(n4526) );
  OR2_X1 U3078 ( .A1(n2677), .A2(n2676), .ZN(n3480) );
  INV_X1 U3079 ( .A(n4794), .ZN(n4797) );
  INV_X1 U3080 ( .A(n4331), .ZN(n4559) );
  NAND2_X1 U3081 ( .A1(n4910), .A2(n4636), .ZN(n4629) );
  NAND2_X1 U3082 ( .A1(n4902), .A2(n4636), .ZN(n4682) );
  INV_X1 U3083 ( .A(n4902), .ZN(n4900) );
  INV_X1 U3084 ( .A(n4842), .ZN(n4841) );
  XNOR2_X1 U3085 ( .A(n2898), .B(n2415), .ZN(n4701) );
  INV_X1 U3086 ( .A(n3459), .ZN(n4854) );
  INV_X1 U3087 ( .A(n3080), .ZN(n4694) );
  NAND4_X1 U3088 ( .A1(n2405), .A2(n2404), .A3(n2403), .A4(n2402), .ZN(n2406)
         );
  NAND4_X1 U3089 ( .A1(n2422), .A2(n2329), .A3(n2436), .A4(n2409), .ZN(n2411)
         );
  NAND2_X1 U3090 ( .A1(n3035), .A2(n3034), .ZN(n2414) );
  NAND2_X1 U3091 ( .A1(n3034), .A2(IR_REG_28__SCAN_IN), .ZN(n2416) );
  NAND2_X4 U3092 ( .A1(n2417), .A2(n2416), .ZN(n3794) );
  NAND2_X1 U3093 ( .A1(n2457), .A2(n2422), .ZN(n2459) );
  NAND2_X1 U3094 ( .A1(n2869), .A2(n2870), .ZN(n2423) );
  NOR2_X1 U3095 ( .A1(n2426), .A2(n2561), .ZN(n2428) );
  NAND2_X1 U3096 ( .A1(n2430), .A2(IR_REG_31__SCAN_IN), .ZN(n2431) );
  MUX2_X1 U3097 ( .A(IR_REG_31__SCAN_IN), .B(n2431), .S(IR_REG_25__SCAN_IN), 
        .Z(n2433) );
  INV_X1 U3098 ( .A(n2426), .ZN(n2432) );
  NAND2_X1 U3099 ( .A1(n2435), .A2(IR_REG_31__SCAN_IN), .ZN(n2465) );
  NAND2_X1 U3100 ( .A1(n2465), .A2(n2464), .ZN(n2467) );
  NAND2_X1 U3101 ( .A1(n2467), .A2(IR_REG_31__SCAN_IN), .ZN(n2437) );
  NAND2_X1 U3102 ( .A1(n2438), .A2(IR_REG_31__SCAN_IN), .ZN(n2439) );
  XNOR2_X2 U3103 ( .A(n2442), .B(IR_REG_30__SCAN_IN), .ZN(n4686) );
  INV_X1 U3104 ( .A(n4686), .ZN(n2446) );
  NAND2_X1 U3105 ( .A1(n2444), .A2(IR_REG_31__SCAN_IN), .ZN(n2445) );
  INV_X1 U3106 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2455) );
  INV_X1 U3107 ( .A(n2447), .ZN(n3031) );
  NAND2_X1 U3108 ( .A1(n2158), .A2(REG0_REG_0__SCAN_IN), .ZN(n2450) );
  NAND2_X1 U3109 ( .A1(n2171), .A2(REG2_REG_0__SCAN_IN), .ZN(n2449) );
  NAND2_X1 U3110 ( .A1(n2483), .A2(REG3_REG_0__SCAN_IN), .ZN(n2448) );
  AND3_X1 U3111 ( .A1(n2450), .A2(n2449), .A3(n2448), .ZN(n2451) );
  NAND2_X2 U3112 ( .A1(n2454), .A2(n3191), .ZN(n2749) );
  NAND2_X1 U3113 ( .A1(n2944), .A2(n2846), .ZN(n2453) );
  AND2_X1 U3114 ( .A1(n2172), .A2(n2453), .ZN(n2469) );
  OR2_X1 U3115 ( .A1(n2454), .A2(n2455), .ZN(n2456) );
  NAND2_X1 U3116 ( .A1(n2469), .A2(n2456), .ZN(n3642) );
  INV_X1 U3117 ( .A(n2944), .ZN(n2463) );
  MUX2_X1 U3118 ( .A(IR_REG_31__SCAN_IN), .B(n2458), .S(IR_REG_22__SCAN_IN), 
        .Z(n2460) );
  INV_X1 U3119 ( .A(n2454), .ZN(n2461) );
  AOI22_X1 U3120 ( .A1(n3645), .A2(n2846), .B1(IR_REG_0__SCAN_IN), .B2(n2461), 
        .ZN(n2462) );
  OAI21_X1 U3121 ( .B1(n2463), .B2(n3003), .A(n2462), .ZN(n3641) );
  NAND2_X1 U3122 ( .A1(n3642), .A2(n3641), .ZN(n3644) );
  OR2_X1 U3123 ( .A1(n2465), .A2(n2464), .ZN(n2466) );
  NAND2_X1 U3124 ( .A1(n4688), .A2(n4307), .ZN(n2880) );
  NAND2_X1 U3125 ( .A1(n2469), .A2(n2832), .ZN(n2470) );
  NAND2_X1 U3126 ( .A1(n3644), .A2(n2470), .ZN(n3670) );
  NAND2_X1 U3127 ( .A1(n2171), .A2(REG2_REG_1__SCAN_IN), .ZN(n2474) );
  NAND2_X1 U3128 ( .A1(n2483), .A2(REG3_REG_1__SCAN_IN), .ZN(n2473) );
  INV_X1 U3129 ( .A(REG1_REG_1__SCAN_IN), .ZN(n3057) );
  NAND2_X1 U3130 ( .A1(n2158), .A2(REG0_REG_1__SCAN_IN), .ZN(n2471) );
  INV_X1 U3131 ( .A(n2904), .ZN(n3147) );
  OAI22_X1 U3132 ( .A1(n2905), .A2(n2749), .B1(n2477), .B2(n3147), .ZN(n2478)
         );
  XNOR2_X1 U3133 ( .A(n2478), .B(n2832), .ZN(n2479) );
  OAI22_X1 U3134 ( .A1(n2905), .A2(n3003), .B1(n2749), .B2(n3147), .ZN(n2480)
         );
  XNOR2_X1 U3135 ( .A(n2479), .B(n2480), .ZN(n3669) );
  NAND2_X1 U3136 ( .A1(n3670), .A2(n3669), .ZN(n3671) );
  INV_X1 U3137 ( .A(n2479), .ZN(n2481) );
  NAND2_X1 U3138 ( .A1(n2481), .A2(n2480), .ZN(n2482) );
  NAND2_X1 U3139 ( .A1(n3671), .A2(n2482), .ZN(n3168) );
  INV_X1 U3140 ( .A(n3168), .ZN(n2493) );
  NAND2_X1 U3141 ( .A1(n2171), .A2(REG2_REG_2__SCAN_IN), .ZN(n2487) );
  NAND2_X1 U3142 ( .A1(n2158), .A2(REG0_REG_2__SCAN_IN), .ZN(n2486) );
  INV_X1 U3143 ( .A(REG1_REG_2__SCAN_IN), .ZN(n3261) );
  NAND3_X1 U3144 ( .A1(n2487), .A2(n2486), .A3(n2485), .ZN(n2488) );
  INV_X1 U3145 ( .A(n3257), .ZN(n2910) );
  OAI22_X1 U3146 ( .A1(n2908), .A2(n2749), .B1(n2910), .B2(n2477), .ZN(n2491)
         );
  XNOR2_X1 U3147 ( .A(n2491), .B(n3001), .ZN(n2494) );
  OAI22_X1 U31480 ( .A1(n2908), .A2(n3003), .B1(n2910), .B2(n2749), .ZN(n2495)
         );
  XNOR2_X1 U31490 ( .A(n2494), .B(n2495), .ZN(n3167) );
  INV_X1 U3150 ( .A(n3167), .ZN(n2492) );
  NAND2_X1 U3151 ( .A1(n2493), .A2(n2492), .ZN(n3169) );
  INV_X1 U3152 ( .A(n2494), .ZN(n2497) );
  INV_X1 U3153 ( .A(n2495), .ZN(n2496) );
  NAND2_X1 U3154 ( .A1(n2497), .A2(n2496), .ZN(n3212) );
  INV_X1 U3155 ( .A(n3212), .ZN(n2512) );
  INV_X1 U3156 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2498) );
  INV_X1 U3157 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2519) );
  NAND2_X1 U3158 ( .A1(n2483), .A2(n2519), .ZN(n2502) );
  NAND2_X1 U3159 ( .A1(n2533), .A2(REG0_REG_3__SCAN_IN), .ZN(n2501) );
  NAND2_X1 U3160 ( .A1(n2171), .A2(REG2_REG_3__SCAN_IN), .ZN(n2500) );
  NAND2_X1 U3161 ( .A1(n4238), .A2(n2846), .ZN(n2509) );
  NAND2_X1 U3162 ( .A1(n2539), .A2(n2399), .ZN(n2504) );
  NAND2_X1 U3163 ( .A1(n2504), .A2(IR_REG_31__SCAN_IN), .ZN(n2506) );
  NAND2_X1 U3164 ( .A1(n2506), .A2(n2505), .ZN(n2526) );
  OR2_X1 U3165 ( .A1(n2506), .A2(n2505), .ZN(n2507) );
  MUX2_X1 U3166 ( .A(n4697), .B(DATAI_3_), .S(n3794), .Z(n2947) );
  NAND2_X1 U3167 ( .A1(n2947), .A2(n2847), .ZN(n2508) );
  NAND2_X1 U3168 ( .A1(n2509), .A2(n2508), .ZN(n2510) );
  INV_X1 U3169 ( .A(n2515), .ZN(n2511) );
  AND2_X1 U3170 ( .A1(n2511), .A2(n2514), .ZN(n2516) );
  NOR2_X1 U3171 ( .A1(n2512), .A2(n2516), .ZN(n2513) );
  NAND2_X1 U3172 ( .A1(n3169), .A2(n2513), .ZN(n2518) );
  NAND2_X1 U3173 ( .A1(n2533), .A2(REG0_REG_4__SCAN_IN), .ZN(n2525) );
  INV_X1 U3174 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2520) );
  NAND2_X1 U3175 ( .A1(n2520), .A2(n2519), .ZN(n2521) );
  AND2_X1 U3176 ( .A1(n2521), .A2(n2551), .ZN(n3630) );
  NAND2_X1 U3177 ( .A1(n2483), .A2(n3630), .ZN(n2524) );
  NAND2_X1 U3178 ( .A1(n2171), .A2(REG2_REG_4__SCAN_IN), .ZN(n2523) );
  INV_X1 U3179 ( .A(REG1_REG_4__SCAN_IN), .ZN(n3065) );
  OR2_X1 U3180 ( .A1(n2484), .A2(n3065), .ZN(n2522) );
  NAND2_X1 U3181 ( .A1(n2526), .A2(IR_REG_31__SCAN_IN), .ZN(n2527) );
  XNOR2_X1 U3182 ( .A(n2527), .B(IR_REG_4__SCAN_IN), .ZN(n4696) );
  MUX2_X1 U3183 ( .A(n4696), .B(DATAI_4_), .S(n3794), .Z(n3622) );
  INV_X1 U3184 ( .A(n3622), .ZN(n3615) );
  OAI22_X1 U3185 ( .A1(n3238), .A2(n3003), .B1(n2749), .B2(n3615), .ZN(n2530)
         );
  XNOR2_X1 U3186 ( .A(n2531), .B(n2530), .ZN(n3279) );
  INV_X1 U3187 ( .A(n3279), .ZN(n2529) );
  NAND2_X1 U3188 ( .A1(n2531), .A2(n2530), .ZN(n2532) );
  NAND2_X1 U3189 ( .A1(n2533), .A2(REG0_REG_5__SCAN_IN), .ZN(n2537) );
  XNOR2_X1 U3190 ( .A(n2551), .B(REG3_REG_5__SCAN_IN), .ZN(n3231) );
  NAND2_X1 U3191 ( .A1(n2483), .A2(n3231), .ZN(n2536) );
  NAND2_X1 U3192 ( .A1(n2171), .A2(REG2_REG_5__SCAN_IN), .ZN(n2535) );
  INV_X1 U3193 ( .A(REG1_REG_5__SCAN_IN), .ZN(n3068) );
  OR2_X1 U3194 ( .A1(n2975), .A2(n3068), .ZN(n2534) );
  NAND2_X1 U3195 ( .A1(n2505), .A2(n2398), .ZN(n2538) );
  NOR2_X1 U3196 ( .A1(IR_REG_2__SCAN_IN), .A2(n2538), .ZN(n2560) );
  NAND2_X1 U3197 ( .A1(n2539), .A2(n2560), .ZN(n2540) );
  NAND2_X1 U3198 ( .A1(n2540), .A2(IR_REG_31__SCAN_IN), .ZN(n2541) );
  XNOR2_X1 U3199 ( .A(n2541), .B(n2400), .ZN(n3124) );
  INV_X1 U3200 ( .A(DATAI_5_), .ZN(n2542) );
  MUX2_X1 U3201 ( .A(n3124), .B(n2542), .S(n3794), .Z(n3229) );
  OAI22_X1 U3202 ( .A1(n3624), .A2(n2749), .B1(n2477), .B2(n3229), .ZN(n2543)
         );
  XNOR2_X1 U3203 ( .A(n2543), .B(n2832), .ZN(n2544) );
  OAI22_X1 U3204 ( .A1(n3624), .A2(n3003), .B1(n2749), .B2(n3229), .ZN(n2545)
         );
  XNOR2_X1 U3205 ( .A(n2544), .B(n2545), .ZN(n3236) );
  INV_X1 U3206 ( .A(n2544), .ZN(n2546) );
  NAND2_X1 U3207 ( .A1(n2546), .A2(n2545), .ZN(n2547) );
  INV_X1 U3208 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2548) );
  OR2_X1 U3209 ( .A1(n2975), .A2(n2548), .ZN(n2557) );
  NAND2_X1 U32100 ( .A1(n2533), .A2(REG0_REG_6__SCAN_IN), .ZN(n2556) );
  INV_X1 U32110 ( .A(n2551), .ZN(n2549) );
  AOI21_X1 U32120 ( .B1(n2549), .B2(REG3_REG_5__SCAN_IN), .A(
        REG3_REG_6__SCAN_IN), .ZN(n2552) );
  NAND2_X1 U32130 ( .A1(REG3_REG_5__SCAN_IN), .A2(REG3_REG_6__SCAN_IN), .ZN(
        n2550) );
  OR2_X1 U32140 ( .A1(n2552), .A2(n2571), .ZN(n3306) );
  INV_X1 U32150 ( .A(n3306), .ZN(n2553) );
  NAND2_X1 U32160 ( .A1(n2483), .A2(n2553), .ZN(n2555) );
  NAND2_X1 U32170 ( .A1(n2700), .A2(REG2_REG_6__SCAN_IN), .ZN(n2554) );
  NAND4_X1 U32180 ( .A1(n2557), .A2(n2556), .A3(n2555), .A4(n2554), .ZN(n3331)
         );
  NAND2_X1 U32190 ( .A1(n3331), .A2(n2558), .ZN(n2567) );
  AND2_X1 U32200 ( .A1(n2559), .A2(n2560), .ZN(n2562) );
  NOR2_X1 U32210 ( .A1(n2562), .A2(n2561), .ZN(n2563) );
  MUX2_X1 U32220 ( .A(n2561), .B(n2563), .S(IR_REG_6__SCAN_IN), .Z(n2565) );
  AND2_X1 U32230 ( .A1(n2564), .A2(n2559), .ZN(n2578) );
  MUX2_X1 U32240 ( .A(n4694), .B(DATAI_6_), .S(n3794), .Z(n3303) );
  NAND2_X1 U32250 ( .A1(n3303), .A2(n2846), .ZN(n2566) );
  NAND2_X1 U32260 ( .A1(n2567), .A2(n2566), .ZN(n3296) );
  NAND2_X1 U32270 ( .A1(n3331), .A2(n2846), .ZN(n2569) );
  NAND2_X1 U32280 ( .A1(n3303), .A2(n2847), .ZN(n2568) );
  NAND2_X1 U32290 ( .A1(n2569), .A2(n2568), .ZN(n2570) );
  XNOR2_X1 U32300 ( .A(n2570), .B(n3001), .ZN(n3297) );
  NAND2_X1 U32310 ( .A1(n2533), .A2(REG0_REG_7__SCAN_IN), .ZN(n2577) );
  OR2_X1 U32320 ( .A1(n2571), .A2(REG3_REG_7__SCAN_IN), .ZN(n2572) );
  AND2_X1 U32330 ( .A1(n2603), .A2(n2572), .ZN(n3336) );
  NAND2_X1 U32340 ( .A1(n2483), .A2(n3336), .ZN(n2576) );
  NAND2_X1 U32350 ( .A1(n2700), .A2(REG2_REG_7__SCAN_IN), .ZN(n2575) );
  INV_X1 U32360 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2573) );
  OR2_X1 U32370 ( .A1(n2975), .A2(n2573), .ZN(n2574) );
  MUX2_X1 U32380 ( .A(n4693), .B(DATAI_7_), .S(n3794), .Z(n3332) );
  INV_X1 U32390 ( .A(n3332), .ZN(n3326) );
  OAI22_X1 U32400 ( .A1(n3300), .A2(n2749), .B1(n2477), .B2(n3326), .ZN(n2579)
         );
  XNOR2_X1 U32410 ( .A(n2579), .B(n2832), .ZN(n2580) );
  OAI22_X1 U32420 ( .A1(n3300), .A2(n3003), .B1(n2749), .B2(n3326), .ZN(n2581)
         );
  XNOR2_X1 U32430 ( .A(n2580), .B(n2581), .ZN(n3307) );
  INV_X1 U32440 ( .A(n2580), .ZN(n2582) );
  NAND2_X1 U32450 ( .A1(n2533), .A2(REG0_REG_8__SCAN_IN), .ZN(n2587) );
  XNOR2_X1 U32460 ( .A(n2603), .B(REG3_REG_8__SCAN_IN), .ZN(n3353) );
  NAND2_X1 U32470 ( .A1(n2483), .A2(n3353), .ZN(n2586) );
  NAND2_X1 U32480 ( .A1(n2700), .A2(REG2_REG_8__SCAN_IN), .ZN(n2585) );
  INV_X1 U32490 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2583) );
  OR2_X1 U32500 ( .A1(n2975), .A2(n2583), .ZN(n2584) );
  INV_X1 U32510 ( .A(IR_REG_7__SCAN_IN), .ZN(n2588) );
  NAND2_X1 U32520 ( .A1(n2589), .A2(n2588), .ZN(n2590) );
  NAND2_X1 U32530 ( .A1(n2590), .A2(IR_REG_31__SCAN_IN), .ZN(n2592) );
  INV_X1 U32540 ( .A(IR_REG_8__SCAN_IN), .ZN(n2591) );
  XNOR2_X1 U32550 ( .A(n2592), .B(n2591), .ZN(n4692) );
  INV_X1 U32560 ( .A(DATAI_8_), .ZN(n2593) );
  OAI22_X1 U32570 ( .A1(n3390), .A2(n2792), .B1(n2477), .B2(n3351), .ZN(n2594)
         );
  XNOR2_X1 U32580 ( .A(n2594), .B(n3001), .ZN(n2595) );
  OAI22_X1 U32590 ( .A1(n3390), .A2(n3003), .B1(n2792), .B2(n3351), .ZN(n2596)
         );
  AND2_X1 U32600 ( .A1(n2595), .A2(n2596), .ZN(n3346) );
  INV_X1 U32610 ( .A(n2595), .ZN(n2598) );
  INV_X1 U32620 ( .A(n2596), .ZN(n2597) );
  NAND2_X1 U32630 ( .A1(n2598), .A2(n2597), .ZN(n3345) );
  OAI21_X1 U32640 ( .B1(n3344), .B2(n3346), .A(n3345), .ZN(n3388) );
  INV_X1 U32650 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2599) );
  OR2_X1 U32660 ( .A1(n2975), .A2(n2599), .ZN(n2608) );
  NAND2_X1 U32670 ( .A1(n2533), .A2(REG0_REG_9__SCAN_IN), .ZN(n2607) );
  INV_X1 U32680 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2601) );
  INV_X1 U32690 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2600) );
  OAI21_X1 U32700 ( .B1(n2603), .B2(n2601), .A(n2600), .ZN(n2604) );
  NAND2_X1 U32710 ( .A1(REG3_REG_8__SCAN_IN), .A2(REG3_REG_9__SCAN_IN), .ZN(
        n2602) );
  AND2_X1 U32720 ( .A1(n2604), .A2(n2620), .ZN(n3393) );
  NAND2_X1 U32730 ( .A1(n2483), .A2(n3393), .ZN(n2606) );
  NAND2_X1 U32740 ( .A1(n2700), .A2(REG2_REG_9__SCAN_IN), .ZN(n2605) );
  NAND4_X1 U32750 ( .A1(n2608), .A2(n2607), .A3(n2606), .A4(n2605), .ZN(n3481)
         );
  NAND2_X1 U32760 ( .A1(n3481), .A2(n2846), .ZN(n2613) );
  NAND2_X1 U32770 ( .A1(n2609), .A2(IR_REG_31__SCAN_IN), .ZN(n2610) );
  MUX2_X1 U32780 ( .A(IR_REG_31__SCAN_IN), .B(n2610), .S(IR_REG_9__SCAN_IN), 
        .Z(n2611) );
  OR2_X1 U32790 ( .A1(n2609), .A2(IR_REG_9__SCAN_IN), .ZN(n2672) );
  MUX2_X1 U32800 ( .A(n3467), .B(DATAI_9_), .S(n3794), .Z(n3392) );
  NAND2_X1 U32810 ( .A1(n3392), .A2(n2847), .ZN(n2612) );
  NAND2_X1 U32820 ( .A1(n2613), .A2(n2612), .ZN(n2614) );
  XNOR2_X1 U32830 ( .A(n2614), .B(n3001), .ZN(n2615) );
  AOI22_X1 U32840 ( .A1(n3481), .A2(n2558), .B1(n3392), .B2(n2846), .ZN(n2616)
         );
  XNOR2_X1 U32850 ( .A(n2615), .B(n2616), .ZN(n3389) );
  INV_X1 U32860 ( .A(n2615), .ZN(n2617) );
  NAND2_X1 U32870 ( .A1(n2617), .A2(n2616), .ZN(n2618) );
  INV_X1 U32880 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2619) );
  OR2_X1 U32890 ( .A1(n2975), .A2(n2619), .ZN(n2625) );
  NAND2_X1 U32900 ( .A1(n2533), .A2(REG0_REG_10__SCAN_IN), .ZN(n2624) );
  NAND2_X1 U32910 ( .A1(n2620), .A2(n4036), .ZN(n2621) );
  AND2_X1 U32920 ( .A1(n2637), .A2(n2621), .ZN(n3490) );
  NAND2_X1 U32930 ( .A1(n2483), .A2(n3490), .ZN(n2623) );
  NAND2_X1 U32940 ( .A1(n2700), .A2(REG2_REG_10__SCAN_IN), .ZN(n2622) );
  NAND4_X1 U32950 ( .A1(n2625), .A2(n2624), .A3(n2623), .A4(n2622), .ZN(n3364)
         );
  NAND2_X1 U32960 ( .A1(n3364), .A2(n2846), .ZN(n2628) );
  NAND2_X1 U32970 ( .A1(n2672), .A2(IR_REG_31__SCAN_IN), .ZN(n2626) );
  XNOR2_X1 U32980 ( .A(n2626), .B(IR_REG_10__SCAN_IN), .ZN(n4857) );
  MUX2_X1 U32990 ( .A(n4857), .B(DATAI_10_), .S(n3794), .Z(n3377) );
  NAND2_X1 U33000 ( .A1(n3377), .A2(n2847), .ZN(n2627) );
  NAND2_X1 U33010 ( .A1(n2628), .A2(n2627), .ZN(n2629) );
  XNOR2_X1 U33020 ( .A(n2629), .B(n2832), .ZN(n2631) );
  AOI22_X1 U33030 ( .A1(n3364), .A2(n2558), .B1(n2846), .B2(n3377), .ZN(n2632)
         );
  XNOR2_X1 U33040 ( .A(n2631), .B(n2632), .ZN(n3487) );
  INV_X1 U33050 ( .A(n2631), .ZN(n2634) );
  INV_X1 U33060 ( .A(n2632), .ZN(n2633) );
  NAND2_X1 U33070 ( .A1(n2634), .A2(n2633), .ZN(n2635) );
  NAND2_X1 U33080 ( .A1(n3485), .A2(n2635), .ZN(n3423) );
  NAND2_X1 U33090 ( .A1(n2533), .A2(REG0_REG_11__SCAN_IN), .ZN(n2643) );
  AND2_X1 U33100 ( .A1(n2637), .A2(n2636), .ZN(n2638) );
  NOR2_X1 U33110 ( .A1(n2646), .A2(n2638), .ZN(n3445) );
  NAND2_X1 U33120 ( .A1(n2483), .A2(n3445), .ZN(n2642) );
  NAND2_X1 U33130 ( .A1(n2700), .A2(REG2_REG_11__SCAN_IN), .ZN(n2641) );
  INV_X1 U33140 ( .A(REG1_REG_11__SCAN_IN), .ZN(n2639) );
  OR2_X1 U33150 ( .A1(n2975), .A2(n2639), .ZN(n2640) );
  OR2_X1 U33160 ( .A1(n2672), .A2(IR_REG_10__SCAN_IN), .ZN(n2644) );
  NAND2_X1 U33170 ( .A1(n2644), .A2(IR_REG_31__SCAN_IN), .ZN(n2652) );
  XNOR2_X1 U33180 ( .A(n2652), .B(IR_REG_11__SCAN_IN), .ZN(n4855) );
  MUX2_X1 U33190 ( .A(n4855), .B(DATAI_11_), .S(n3794), .Z(n3435) );
  OAI22_X1 U33200 ( .A1(n3409), .A2(n3003), .B1(n2792), .B2(n3443), .ZN(n3425)
         );
  INV_X2 U33210 ( .A(n2846), .ZN(n2792) );
  OAI22_X1 U33220 ( .A1(n3409), .A2(n2792), .B1(n2477), .B2(n3443), .ZN(n2645)
         );
  XNOR2_X1 U33230 ( .A(n2645), .B(n3001), .ZN(n3424) );
  NAND2_X1 U33240 ( .A1(n2158), .A2(REG0_REG_12__SCAN_IN), .ZN(n2651) );
  OR2_X1 U33250 ( .A1(n2646), .A2(REG3_REG_12__SCAN_IN), .ZN(n2647) );
  NAND2_X1 U33260 ( .A1(n2646), .A2(REG3_REG_12__SCAN_IN), .ZN(n2662) );
  AND2_X1 U33270 ( .A1(n2647), .A2(n2662), .ZN(n3501) );
  NAND2_X1 U33280 ( .A1(n2483), .A2(n3501), .ZN(n2650) );
  NAND2_X1 U33290 ( .A1(n2700), .A2(REG2_REG_12__SCAN_IN), .ZN(n2649) );
  INV_X1 U33300 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4740) );
  OR2_X1 U33310 ( .A1(n2975), .A2(n4740), .ZN(n2648) );
  INV_X1 U33320 ( .A(IR_REG_11__SCAN_IN), .ZN(n2669) );
  NAND2_X1 U33330 ( .A1(n2652), .A2(n2669), .ZN(n2653) );
  NAND2_X1 U33340 ( .A1(n2653), .A2(IR_REG_31__SCAN_IN), .ZN(n2654) );
  XNOR2_X1 U33350 ( .A(n2654), .B(IR_REG_12__SCAN_IN), .ZN(n3459) );
  INV_X1 U33360 ( .A(DATAI_12_), .ZN(n2655) );
  MUX2_X1 U33370 ( .A(n4854), .B(n2655), .S(n3794), .Z(n3499) );
  OAI22_X1 U33380 ( .A1(n3539), .A2(n2792), .B1(n2477), .B2(n3499), .ZN(n2656)
         );
  XNOR2_X1 U33390 ( .A(n2656), .B(n3001), .ZN(n2657) );
  OAI22_X1 U33400 ( .A1(n3539), .A2(n3003), .B1(n2792), .B2(n3499), .ZN(n2658)
         );
  AND2_X1 U33410 ( .A1(n2657), .A2(n2658), .ZN(n3493) );
  INV_X1 U33420 ( .A(n2657), .ZN(n2660) );
  INV_X1 U33430 ( .A(n2658), .ZN(n2659) );
  NAND2_X1 U33440 ( .A1(n2660), .A2(n2659), .ZN(n3492) );
  NAND2_X1 U33450 ( .A1(n2158), .A2(REG0_REG_13__SCAN_IN), .ZN(n2667) );
  NAND2_X1 U33460 ( .A1(n2662), .A2(n2661), .ZN(n2663) );
  AND2_X1 U33470 ( .A1(n2684), .A2(n2663), .ZN(n3543) );
  NAND2_X1 U33480 ( .A1(n2483), .A2(n3543), .ZN(n2666) );
  NAND2_X1 U33490 ( .A1(n2700), .A2(REG2_REG_13__SCAN_IN), .ZN(n2665) );
  INV_X1 U33500 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3577) );
  OR2_X1 U33510 ( .A1(n2975), .A2(n3577), .ZN(n2664) );
  INV_X1 U33520 ( .A(IR_REG_12__SCAN_IN), .ZN(n2670) );
  INV_X1 U3353 ( .A(IR_REG_10__SCAN_IN), .ZN(n2668) );
  NAND3_X1 U33540 ( .A1(n2670), .A2(n2669), .A3(n2668), .ZN(n2671) );
  NOR2_X1 U3355 ( .A1(n2672), .A2(n2671), .ZN(n2675) );
  NOR2_X1 U3356 ( .A1(n2675), .A2(n2561), .ZN(n2673) );
  MUX2_X1 U3357 ( .A(n2561), .B(n2673), .S(IR_REG_13__SCAN_IN), .Z(n2677) );
  INV_X1 U3358 ( .A(IR_REG_13__SCAN_IN), .ZN(n2674) );
  NAND2_X1 U3359 ( .A1(n2675), .A2(n2674), .ZN(n2705) );
  INV_X1 U3360 ( .A(n2705), .ZN(n2676) );
  INV_X1 U3361 ( .A(DATAI_13_), .ZN(n2678) );
  MUX2_X1 U3362 ( .A(n3480), .B(n2678), .S(n3794), .Z(n2955) );
  OAI22_X1 U3363 ( .A1(n3408), .A2(n2792), .B1(n2477), .B2(n2955), .ZN(n2679)
         );
  XNOR2_X1 U3364 ( .A(n2679), .B(n2832), .ZN(n3535) );
  NAND2_X1 U3365 ( .A1(n2680), .A2(n3536), .ZN(n2683) );
  NAND2_X1 U3366 ( .A1(n2681), .A2(n2321), .ZN(n2682) );
  NAND2_X1 U3367 ( .A1(n2683), .A2(n2682), .ZN(n3580) );
  INV_X1 U3368 ( .A(n3580), .ZN(n2697) );
  NAND2_X1 U3369 ( .A1(n2158), .A2(REG0_REG_14__SCAN_IN), .ZN(n2689) );
  AND2_X1 U3370 ( .A1(n2684), .A2(n4098), .ZN(n2685) );
  NOR2_X1 U3371 ( .A1(n2698), .A2(n2685), .ZN(n3587) );
  NAND2_X1 U3372 ( .A1(n2483), .A2(n3587), .ZN(n2688) );
  NAND2_X1 U3373 ( .A1(n2700), .A2(REG2_REG_14__SCAN_IN), .ZN(n2687) );
  INV_X1 U3374 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4750) );
  OR2_X1 U3375 ( .A1(n2975), .A2(n4750), .ZN(n2686) );
  NAND2_X1 U3376 ( .A1(n2705), .A2(IR_REG_31__SCAN_IN), .ZN(n2690) );
  XNOR2_X1 U3377 ( .A(n2690), .B(IR_REG_14__SCAN_IN), .ZN(n4757) );
  MUX2_X1 U3378 ( .A(n4757), .B(DATAI_14_), .S(n3794), .Z(n2927) );
  OAI22_X1 U3379 ( .A1(n3782), .A2(n2792), .B1(n3585), .B2(n2477), .ZN(n2691)
         );
  XNOR2_X1 U3380 ( .A(n2691), .B(n3001), .ZN(n2692) );
  OAI22_X1 U3381 ( .A1(n3782), .A2(n3003), .B1(n3585), .B2(n2792), .ZN(n2693)
         );
  AND2_X1 U3382 ( .A1(n2692), .A2(n2693), .ZN(n3581) );
  INV_X1 U3383 ( .A(n2692), .ZN(n2695) );
  INV_X1 U3384 ( .A(n2693), .ZN(n2694) );
  NAND2_X1 U3385 ( .A1(n2533), .A2(REG0_REG_15__SCAN_IN), .ZN(n2704) );
  NAND2_X1 U3386 ( .A1(n2698), .A2(REG3_REG_15__SCAN_IN), .ZN(n2711) );
  OR2_X1 U3387 ( .A1(n2698), .A2(REG3_REG_15__SCAN_IN), .ZN(n2699) );
  AND2_X1 U3388 ( .A1(n2711), .A2(n2699), .ZN(n3786) );
  NAND2_X1 U3389 ( .A1(n2483), .A2(n3786), .ZN(n2703) );
  NAND2_X1 U3390 ( .A1(n2700), .A2(REG2_REG_15__SCAN_IN), .ZN(n2702) );
  INV_X1 U3391 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4286) );
  OR2_X1 U3392 ( .A1(n2975), .A2(n4286), .ZN(n2701) );
  NAND2_X1 U3393 ( .A1(n2706), .A2(IR_REG_31__SCAN_IN), .ZN(n2708) );
  INV_X1 U3394 ( .A(IR_REG_15__SCAN_IN), .ZN(n2707) );
  NAND2_X1 U3395 ( .A1(n2708), .A2(n2707), .ZN(n2717) );
  OR2_X1 U3396 ( .A1(n2708), .A2(n2707), .ZN(n2709) );
  MUX2_X1 U3397 ( .A(n4298), .B(DATAI_15_), .S(n3794), .Z(n3785) );
  OAI22_X1 U3398 ( .A1(n3603), .A2(n2792), .B1(n2477), .B2(n3566), .ZN(n2710)
         );
  XNOR2_X1 U3399 ( .A(n2710), .B(n3001), .ZN(n2724) );
  OAI22_X1 U3400 ( .A1(n3603), .A2(n3003), .B1(n2792), .B2(n3566), .ZN(n3777)
         );
  INV_X1 U3401 ( .A(n3777), .ZN(n3700) );
  NAND2_X1 U3402 ( .A1(n2533), .A2(REG0_REG_16__SCAN_IN), .ZN(n2716) );
  NAND2_X1 U3403 ( .A1(n2711), .A2(n4139), .ZN(n2712) );
  AND2_X1 U3404 ( .A1(n2739), .A2(n2712), .ZN(n3707) );
  NAND2_X1 U3405 ( .A1(n2483), .A2(n3707), .ZN(n2715) );
  NAND2_X1 U3406 ( .A1(n2700), .A2(REG2_REG_16__SCAN_IN), .ZN(n2714) );
  INV_X1 U3407 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4777) );
  OR2_X1 U3408 ( .A1(n2975), .A2(n4777), .ZN(n2713) );
  NAND2_X1 U3409 ( .A1(n2717), .A2(IR_REG_31__SCAN_IN), .ZN(n2719) );
  INV_X1 U3410 ( .A(IR_REG_16__SCAN_IN), .ZN(n2718) );
  INV_X1 U3411 ( .A(n4850), .ZN(n2720) );
  MUX2_X1 U3412 ( .A(n2720), .B(DATAI_16_), .S(n3794), .Z(n3594) );
  OAI22_X1 U3413 ( .A1(n3779), .A2(n2792), .B1(n3705), .B2(n2477), .ZN(n2721)
         );
  XNOR2_X1 U3414 ( .A(n2721), .B(n3001), .ZN(n2723) );
  OAI22_X1 U3415 ( .A1(n3779), .A2(n3003), .B1(n3705), .B2(n2792), .ZN(n2722)
         );
  NOR2_X1 U3416 ( .A1(n2723), .A2(n2722), .ZN(n2726) );
  AOI21_X1 U3417 ( .B1(n2723), .B2(n2722), .A(n2726), .ZN(n3701) );
  INV_X1 U3418 ( .A(n2726), .ZN(n2727) );
  NAND2_X1 U3419 ( .A1(n2158), .A2(REG0_REG_17__SCAN_IN), .ZN(n2731) );
  XNOR2_X1 U3420 ( .A(n2739), .B(REG3_REG_17__SCAN_IN), .ZN(n4553) );
  NAND2_X1 U3421 ( .A1(n2483), .A2(n4553), .ZN(n2730) );
  NAND2_X1 U3422 ( .A1(n2700), .A2(REG2_REG_17__SCAN_IN), .ZN(n2729) );
  INV_X1 U3423 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4627) );
  OR2_X1 U3424 ( .A1(n2975), .A2(n4627), .ZN(n2728) );
  NAND2_X1 U3425 ( .A1(n2732), .A2(IR_REG_31__SCAN_IN), .ZN(n2733) );
  XNOR2_X1 U3426 ( .A(n2733), .B(IR_REG_17__SCAN_IN), .ZN(n4301) );
  INV_X1 U3427 ( .A(n4301), .ZN(n4848) );
  INV_X1 U3428 ( .A(DATAI_17_), .ZN(n4847) );
  MUX2_X1 U3429 ( .A(n4848), .B(n4847), .S(n3794), .Z(n4549) );
  OAI22_X1 U3430 ( .A1(n4529), .A2(n2792), .B1(n2477), .B2(n4549), .ZN(n2734)
         );
  XNOR2_X1 U3431 ( .A(n2734), .B(n3001), .ZN(n2736) );
  OAI22_X1 U3432 ( .A1(n4529), .A2(n3003), .B1(n2792), .B2(n4549), .ZN(n2735)
         );
  NAND2_X1 U3433 ( .A1(n2736), .A2(n2735), .ZN(n3711) );
  NAND2_X1 U3434 ( .A1(n2533), .A2(REG0_REG_18__SCAN_IN), .ZN(n2745) );
  INV_X1 U3435 ( .A(n2739), .ZN(n2737) );
  AOI21_X1 U3436 ( .B1(n2737), .B2(REG3_REG_17__SCAN_IN), .A(
        REG3_REG_18__SCAN_IN), .ZN(n2740) );
  NAND2_X1 U3437 ( .A1(REG3_REG_17__SCAN_IN), .A2(REG3_REG_18__SCAN_IN), .ZN(
        n2738) );
  OR2_X1 U3438 ( .A1(n2740), .A2(n2750), .ZN(n4520) );
  INV_X1 U3439 ( .A(n4520), .ZN(n2741) );
  NAND2_X1 U3440 ( .A1(n2483), .A2(n2741), .ZN(n2744) );
  NAND2_X1 U3441 ( .A1(n2700), .A2(REG2_REG_18__SCAN_IN), .ZN(n2743) );
  INV_X1 U3442 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4281) );
  OR2_X1 U3443 ( .A1(n2975), .A2(n4281), .ZN(n2742) );
  OR2_X1 U3444 ( .A1(n2746), .A2(n2561), .ZN(n2747) );
  XNOR2_X1 U3445 ( .A(n2747), .B(IR_REG_18__SCAN_IN), .ZN(n4302) );
  MUX2_X1 U3446 ( .A(n4302), .B(DATAI_18_), .S(n3794), .Z(n4524) );
  INV_X1 U3447 ( .A(n4524), .ZN(n4517) );
  OAI22_X1 U3448 ( .A1(n4542), .A2(n2792), .B1(n2477), .B2(n4517), .ZN(n2748)
         );
  XNOR2_X1 U3449 ( .A(n2748), .B(n3001), .ZN(n3754) );
  OAI22_X1 U3450 ( .A1(n4542), .A2(n3003), .B1(n2749), .B2(n4517), .ZN(n3753)
         );
  NAND2_X1 U3451 ( .A1(n2158), .A2(REG0_REG_19__SCAN_IN), .ZN(n2755) );
  NOR2_X1 U3452 ( .A1(n2750), .A2(REG3_REG_19__SCAN_IN), .ZN(n2751) );
  NOR2_X1 U3453 ( .A1(n2763), .A2(n2751), .ZN(n4508) );
  NAND2_X1 U3454 ( .A1(n2483), .A2(n4508), .ZN(n2754) );
  NAND2_X1 U3455 ( .A1(n2700), .A2(REG2_REG_19__SCAN_IN), .ZN(n2753) );
  INV_X1 U3456 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4620) );
  OR2_X1 U3457 ( .A1(n2975), .A2(n4620), .ZN(n2752) );
  MUX2_X1 U34580 ( .A(n4691), .B(DATAI_19_), .S(n3794), .Z(n3665) );
  OAI22_X1 U34590 ( .A1(n4475), .A2(n2792), .B1(n2477), .B2(n4506), .ZN(n2756)
         );
  XNOR2_X1 U3460 ( .A(n2756), .B(n3001), .ZN(n2759) );
  OAI22_X1 U3461 ( .A1(n4475), .A2(n3003), .B1(n2792), .B2(n4506), .ZN(n2758)
         );
  NOR3_X1 U3462 ( .A1(n3660), .A2(n3753), .A3(n3754), .ZN(n2760) );
  NOR2_X1 U3463 ( .A1(n2759), .A2(n2758), .ZN(n3661) );
  NAND2_X1 U3464 ( .A1(n2158), .A2(REG0_REG_20__SCAN_IN), .ZN(n2768) );
  OR2_X1 U3465 ( .A1(n2763), .A2(REG3_REG_20__SCAN_IN), .ZN(n2764) );
  AND2_X1 U3466 ( .A1(n2774), .A2(n2764), .ZN(n4484) );
  NAND2_X1 U34670 ( .A1(n2483), .A2(n4484), .ZN(n2767) );
  NAND2_X1 U3468 ( .A1(n2700), .A2(REG2_REG_20__SCAN_IN), .ZN(n2766) );
  INV_X1 U34690 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4616) );
  OR2_X1 U3470 ( .A1(n2975), .A2(n4616), .ZN(n2765) );
  OAI22_X1 U34710 ( .A1(n4498), .A2(n2792), .B1(n2477), .B2(n4481), .ZN(n2769)
         );
  XNOR2_X1 U3472 ( .A(n2769), .B(n3001), .ZN(n2770) );
  OAI22_X1 U34730 ( .A1(n4498), .A2(n3003), .B1(n2792), .B2(n4481), .ZN(n2771)
         );
  NAND2_X1 U3474 ( .A1(n2770), .A2(n2771), .ZN(n3733) );
  NAND2_X1 U34750 ( .A1(n3681), .A2(n3733), .ZN(n3732) );
  INV_X1 U3476 ( .A(n2770), .ZN(n2773) );
  INV_X1 U34770 ( .A(n2771), .ZN(n2772) );
  NAND2_X1 U3478 ( .A1(n2773), .A2(n2772), .ZN(n3735) );
  NAND2_X1 U34790 ( .A1(n3732), .A2(n3735), .ZN(n3677) );
  INV_X1 U3480 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4612) );
  OR2_X1 U34810 ( .A1(n2975), .A2(n4612), .ZN(n2779) );
  NAND2_X1 U3482 ( .A1(n2533), .A2(REG0_REG_21__SCAN_IN), .ZN(n2778) );
  NAND2_X1 U34830 ( .A1(n2774), .A2(n4039), .ZN(n2775) );
  AND2_X1 U3484 ( .A1(n2786), .A2(n2775), .ZN(n4462) );
  NAND2_X1 U34850 ( .A1(n2483), .A2(n4462), .ZN(n2777) );
  NAND2_X1 U3486 ( .A1(n2700), .A2(REG2_REG_21__SCAN_IN), .ZN(n2776) );
  NAND2_X1 U34870 ( .A1(n4473), .A2(n2846), .ZN(n2781) );
  OR2_X1 U3488 ( .A1(n4459), .A2(n2477), .ZN(n2780) );
  NAND2_X1 U34890 ( .A1(n2781), .A2(n2780), .ZN(n2782) );
  XNOR2_X1 U3490 ( .A(n2782), .B(n2832), .ZN(n2785) );
  NOR2_X1 U34910 ( .A1(n2792), .A2(n4459), .ZN(n2783) );
  AOI21_X1 U3492 ( .B1(n4473), .B2(n2558), .A(n2783), .ZN(n2784) );
  AND2_X1 U34930 ( .A1(n2785), .A2(n2784), .ZN(n3678) );
  OR2_X1 U3494 ( .A1(n2785), .A2(n2784), .ZN(n3679) );
  INV_X1 U34950 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4145) );
  OR2_X1 U3496 ( .A1(n2975), .A2(n4145), .ZN(n2791) );
  NAND2_X1 U34970 ( .A1(n2158), .A2(REG0_REG_22__SCAN_IN), .ZN(n2790) );
  INV_X1 U3498 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3745) );
  NAND2_X1 U34990 ( .A1(n2786), .A2(n3745), .ZN(n2787) );
  NAND2_X1 U3500 ( .A1(n2796), .A2(n2787), .ZN(n4443) );
  INV_X1 U35010 ( .A(n4443), .ZN(n3750) );
  NAND2_X1 U3502 ( .A1(n2483), .A2(n3750), .ZN(n2789) );
  NAND2_X1 U35030 ( .A1(n2700), .A2(REG2_REG_22__SCAN_IN), .ZN(n2788) );
  NAND4_X1 U3504 ( .A1(n2791), .A2(n2790), .A3(n2789), .A4(n2788), .ZN(n4454)
         );
  OAI22_X1 U35050 ( .A1(n4423), .A2(n2792), .B1(n3746), .B2(n2477), .ZN(n2793)
         );
  XNOR2_X1 U35060 ( .A(n2793), .B(n3001), .ZN(n2795) );
  OAI22_X1 U35070 ( .A1(n4423), .A2(n3003), .B1(n3746), .B2(n2792), .ZN(n2794)
         );
  XNOR2_X1 U35080 ( .A(n2795), .B(n2794), .ZN(n3744) );
  NOR2_X1 U35090 ( .A1(n2795), .A2(n2794), .ZN(n3650) );
  INV_X1 U35100 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4135) );
  INV_X1 U35110 ( .A(n2807), .ZN(n2798) );
  NAND2_X1 U35120 ( .A1(n2796), .A2(n4135), .ZN(n2797) );
  NAND2_X1 U35130 ( .A1(n2798), .A2(n2797), .ZN(n4427) );
  AOI22_X1 U35140 ( .A1(n3793), .A2(REG1_REG_23__SCAN_IN), .B1(n2158), .B2(
        REG0_REG_23__SCAN_IN), .ZN(n2800) );
  NAND2_X1 U35150 ( .A1(n2700), .A2(REG2_REG_23__SCAN_IN), .ZN(n2799) );
  OAI22_X1 U35160 ( .A1(n4440), .A2(n2792), .B1(n2477), .B2(n4425), .ZN(n2802)
         );
  XNOR2_X1 U35170 ( .A(n2802), .B(n3001), .ZN(n2803) );
  OAI22_X1 U35180 ( .A1(n4440), .A2(n3003), .B1(n2792), .B2(n4425), .ZN(n2804)
         );
  XNOR2_X1 U35190 ( .A(n2803), .B(n2804), .ZN(n3649) );
  INV_X1 U35200 ( .A(n2803), .ZN(n2806) );
  INV_X1 U35210 ( .A(n2804), .ZN(n2805) );
  NOR2_X1 U35220 ( .A1(n2806), .A2(n2805), .ZN(n2815) );
  NOR2_X1 U35230 ( .A1(n2807), .A2(REG3_REG_24__SCAN_IN), .ZN(n2808) );
  OR2_X1 U35240 ( .A1(n2816), .A2(n2808), .ZN(n4405) );
  AOI22_X1 U35250 ( .A1(n3793), .A2(REG1_REG_24__SCAN_IN), .B1(n2533), .B2(
        REG0_REG_24__SCAN_IN), .ZN(n2810) );
  NAND2_X1 U35260 ( .A1(n2700), .A2(REG2_REG_24__SCAN_IN), .ZN(n2809) );
  NAND2_X1 U35270 ( .A1(n4420), .A2(n2558), .ZN(n2812) );
  OR2_X1 U35280 ( .A1(n4403), .A2(n2792), .ZN(n2811) );
  NAND2_X1 U35290 ( .A1(n2812), .A2(n2811), .ZN(n2814) );
  AOI22_X1 U35300 ( .A1(n4420), .A2(n2846), .B1(n2847), .B2(n3726), .ZN(n2813)
         );
  XNOR2_X1 U35310 ( .A(n2813), .B(n3001), .ZN(n3721) );
  OAI21_X2 U35320 ( .B1(n3648), .B2(n2815), .A(n2814), .ZN(n3718) );
  NOR2_X1 U35330 ( .A1(n2816), .A2(REG3_REG_25__SCAN_IN), .ZN(n2817) );
  AOI22_X1 U35340 ( .A1(n3793), .A2(REG1_REG_25__SCAN_IN), .B1(n2158), .B2(
        REG0_REG_25__SCAN_IN), .ZN(n2819) );
  NAND2_X1 U35350 ( .A1(n2700), .A2(REG2_REG_25__SCAN_IN), .ZN(n2818) );
  NOR2_X1 U35360 ( .A1(n2477), .A2(n4382), .ZN(n2820) );
  AOI21_X1 U35370 ( .B1(n4398), .B2(n2846), .A(n2820), .ZN(n2821) );
  XNOR2_X1 U35380 ( .A(n2821), .B(n3001), .ZN(n2824) );
  NOR2_X1 U35390 ( .A1(n2792), .A2(n4382), .ZN(n2822) );
  AOI21_X1 U35400 ( .B1(n4398), .B2(n2558), .A(n2822), .ZN(n2823) );
  NAND2_X1 U35410 ( .A1(n2824), .A2(n2823), .ZN(n3690) );
  NOR2_X1 U35420 ( .A1(n2824), .A2(n2823), .ZN(n3689) );
  INV_X1 U35430 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3768) );
  XNOR2_X1 U35440 ( .A(n2839), .B(n3768), .ZN(n4367) );
  NAND2_X1 U35450 ( .A1(n4367), .A2(n2483), .ZN(n2829) );
  INV_X1 U35460 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4591) );
  NAND2_X1 U35470 ( .A1(n2700), .A2(REG2_REG_26__SCAN_IN), .ZN(n2826) );
  NAND2_X1 U35480 ( .A1(n2158), .A2(REG0_REG_26__SCAN_IN), .ZN(n2825) );
  OAI211_X1 U35490 ( .C1(n2975), .C2(n4591), .A(n2826), .B(n2825), .ZN(n2827)
         );
  INV_X1 U35500 ( .A(n2827), .ZN(n2828) );
  NAND2_X1 U35510 ( .A1(n4378), .A2(n2846), .ZN(n2831) );
  OR2_X1 U35520 ( .A1(n4365), .A2(n2477), .ZN(n2830) );
  NAND2_X1 U35530 ( .A1(n2831), .A2(n2830), .ZN(n2833) );
  XNOR2_X1 U35540 ( .A(n2833), .B(n2832), .ZN(n2836) );
  NOR2_X1 U35550 ( .A1(n2792), .A2(n4365), .ZN(n2834) );
  AOI21_X1 U35560 ( .B1(n4378), .B2(n2558), .A(n2834), .ZN(n2835) );
  OR2_X1 U35570 ( .A1(n2836), .A2(n2835), .ZN(n3764) );
  AND2_X1 U35580 ( .A1(n2836), .A2(n2835), .ZN(n3763) );
  AOI21_X1 U35590 ( .B1(n3767), .B2(n3764), .A(n3763), .ZN(n3000) );
  NAND2_X1 U35600 ( .A1(n2839), .A2(REG3_REG_26__SCAN_IN), .ZN(n2837) );
  INV_X1 U35610 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4035) );
  NAND2_X1 U35620 ( .A1(n2837), .A2(n4035), .ZN(n2840) );
  AND2_X1 U35630 ( .A1(REG3_REG_27__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2838) );
  NAND2_X1 U35640 ( .A1(n2839), .A2(n2838), .ZN(n2887) );
  NAND2_X1 U35650 ( .A1(n2840), .A2(n2887), .ZN(n2873) );
  INV_X1 U35660 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4030) );
  NAND2_X1 U35670 ( .A1(n2700), .A2(REG2_REG_27__SCAN_IN), .ZN(n2842) );
  NAND2_X1 U35680 ( .A1(n2158), .A2(REG0_REG_27__SCAN_IN), .ZN(n2841) );
  OAI211_X1 U35690 ( .C1(n2975), .C2(n4030), .A(n2842), .B(n2841), .ZN(n2843)
         );
  INV_X1 U35700 ( .A(n2843), .ZN(n2844) );
  NAND2_X1 U35710 ( .A1(n4361), .A2(n2846), .ZN(n2849) );
  NAND2_X1 U35720 ( .A1(n2847), .A2(n4347), .ZN(n2848) );
  NAND2_X1 U35730 ( .A1(n2849), .A2(n2848), .ZN(n2850) );
  XNOR2_X1 U35740 ( .A(n2850), .B(n3001), .ZN(n3009) );
  NOR2_X1 U35750 ( .A1(n2792), .A2(n2968), .ZN(n2851) );
  AOI21_X1 U35760 ( .B1(n4361), .B2(n2558), .A(n2851), .ZN(n3007) );
  XNOR2_X1 U35770 ( .A(n3009), .B(n3007), .ZN(n2999) );
  XNOR2_X1 U35780 ( .A(n3000), .B(n2999), .ZN(n2903) );
  NAND2_X1 U35790 ( .A1(n3026), .A2(B_REG_SCAN_IN), .ZN(n2853) );
  MUX2_X1 U35800 ( .A(n2853), .B(B_REG_SCAN_IN), .S(n2852), .Z(n2854) );
  INV_X1 U35810 ( .A(n2866), .ZN(n4687) );
  NOR4_X1 U3582 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_19__SCAN_IN), .ZN(n2858) );
  NOR4_X1 U3583 ( .A1(D_REG_12__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_7__SCAN_IN), .A4(D_REG_14__SCAN_IN), .ZN(n2857) );
  NOR4_X1 U3584 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2856) );
  NOR4_X1 U3585 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_22__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2855) );
  AND4_X1 U3586 ( .A1(n2858), .A2(n2857), .A3(n2856), .A4(n2855), .ZN(n2864)
         );
  NOR2_X1 U3587 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_5__SCAN_IN), .ZN(n2862) );
  NOR4_X1 U3588 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2861) );
  NOR4_X1 U3589 ( .A1(D_REG_3__SCAN_IN), .A2(D_REG_16__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_4__SCAN_IN), .ZN(n2860) );
  NOR4_X1 U3590 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_8__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2859) );
  AND4_X1 U3591 ( .A1(n2862), .A2(n2861), .A3(n2860), .A4(n2859), .ZN(n2863)
         );
  NAND2_X1 U3592 ( .A1(n2864), .A2(n2863), .ZN(n2984) );
  INV_X1 U3593 ( .A(D_REG_1__SCAN_IN), .ZN(n3042) );
  OR2_X1 U3594 ( .A1(n2984), .A2(n3042), .ZN(n2865) );
  NAND2_X1 U3595 ( .A1(n2866), .A2(n3026), .ZN(n2985) );
  INV_X1 U3596 ( .A(n2985), .ZN(n3041) );
  AOI21_X1 U3597 ( .B1(n3038), .B2(n2865), .A(n3041), .ZN(n3184) );
  INV_X1 U3598 ( .A(n2852), .ZN(n2867) );
  NAND2_X1 U3599 ( .A1(n2867), .A2(n2866), .ZN(n3039) );
  XNOR2_X1 U3600 ( .A(n2869), .B(n2870), .ZN(n3044) );
  NOR2_X1 U3601 ( .A1(n2941), .A2(n3862), .ZN(n3045) );
  INV_X1 U3602 ( .A(n3045), .ZN(n2971) );
  INV_X1 U3603 ( .A(n3929), .ZN(n4690) );
  NAND2_X1 U3604 ( .A1(n3150), .A2(n4691), .ZN(n2871) );
  NAND3_X1 U3605 ( .A1(n2971), .A2(n4565), .A3(n2871), .ZN(n2874) );
  NOR2_X1 U3606 ( .A1(n3182), .A2(n2874), .ZN(n2872) );
  INV_X1 U3607 ( .A(n2873), .ZN(n4348) );
  INV_X1 U3608 ( .A(n2896), .ZN(n2881) );
  NAND2_X1 U3609 ( .A1(n2874), .A2(n4565), .ZN(n2875) );
  NAND2_X1 U3610 ( .A1(n2881), .A2(n2875), .ZN(n2878) );
  NAND2_X1 U3611 ( .A1(n3929), .A2(n4307), .ZN(n2876) );
  AND2_X1 U3612 ( .A1(n3045), .A2(n2876), .ZN(n3181) );
  INV_X1 U3613 ( .A(n3181), .ZN(n2877) );
  NAND2_X1 U3614 ( .A1(n2878), .A2(n2877), .ZN(n3172) );
  NAND2_X1 U3615 ( .A1(n2454), .A2(n3044), .ZN(n2879) );
  OAI21_X1 U3616 ( .B1(n3172), .B2(n2879), .A(STATE_REG_SCAN_IN), .ZN(n2882)
         );
  INV_X1 U3617 ( .A(n4843), .ZN(n3024) );
  NAND2_X1 U3618 ( .A1(n2881), .A2(n2895), .ZN(n3173) );
  NOR2_X1 U3619 ( .A1(n3182), .A2(n4565), .ZN(n2883) );
  NAND2_X1 U3620 ( .A1(n2896), .A2(n2883), .ZN(n2885) );
  AND2_X1 U3621 ( .A1(n3929), .A2(n4691), .ZN(n4822) );
  NAND2_X1 U3622 ( .A1(n4822), .A2(n2941), .ZN(n3255) );
  NOR2_X1 U3623 ( .A1(n3255), .A2(n4689), .ZN(n2982) );
  INV_X1 U3624 ( .A(n2982), .ZN(n2884) );
  NAND2_X1 U3625 ( .A1(n3784), .A2(n4347), .ZN(n2886) );
  OAI21_X1 U3626 ( .B1(STATE_REG_SCAN_IN), .B2(n4035), .A(n2886), .ZN(n2901)
         );
  INV_X1 U3627 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3014) );
  NAND2_X1 U3628 ( .A1(n2887), .A2(n3014), .ZN(n2888) );
  NAND2_X1 U3629 ( .A1(n3634), .A2(n2483), .ZN(n2894) );
  INV_X1 U3630 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2891) );
  NAND2_X1 U3631 ( .A1(n2158), .A2(REG0_REG_28__SCAN_IN), .ZN(n2890) );
  NAND2_X1 U3632 ( .A1(n2700), .A2(REG2_REG_28__SCAN_IN), .ZN(n2889) );
  OAI211_X1 U3633 ( .C1(n2891), .C2(n2975), .A(n2890), .B(n2889), .ZN(n2892)
         );
  INV_X1 U3634 ( .A(n2892), .ZN(n2893) );
  NAND2_X1 U3635 ( .A1(n2441), .A2(n3034), .ZN(n2897) );
  NAND2_X1 U3636 ( .A1(n2897), .A2(IR_REG_31__SCAN_IN), .ZN(n2898) );
  INV_X1 U3637 ( .A(n4378), .ZN(n4345) );
  INV_X1 U3638 ( .A(n4701), .ZN(n4250) );
  OAI22_X1 U3639 ( .A1(n4326), .A2(n3780), .B1(n4345), .B2(n3781), .ZN(n2900)
         );
  AOI211_X1 U3640 ( .C1(n4348), .C2(n3787), .A(n2901), .B(n2900), .ZN(n2902)
         );
  OAI21_X1 U3641 ( .B1(n2903), .B2(n3790), .A(n2902), .ZN(U3211) );
  INV_X1 U3642 ( .A(n2905), .ZN(n2906) );
  NAND2_X1 U3643 ( .A1(n2906), .A2(n3147), .ZN(n3867) );
  AND2_X1 U3644 ( .A1(n2944), .A2(n3645), .ZN(n3138) );
  NAND2_X1 U3645 ( .A1(n2943), .A2(n3138), .ZN(n3140) );
  CLKBUF_X1 U3646 ( .A(n2906), .Z(n4239) );
  NAND2_X1 U3647 ( .A1(n4239), .A2(n2904), .ZN(n2907) );
  INV_X1 U3648 ( .A(n3245), .ZN(n2909) );
  NAND2_X1 U3649 ( .A1(n3672), .A2(n2910), .ZN(n3874) );
  NAND2_X1 U3650 ( .A1(n2908), .A2(n2910), .ZN(n2911) );
  NAND2_X1 U3651 ( .A1(n3246), .A2(n2911), .ZN(n3197) );
  NAND2_X1 U3652 ( .A1(n4238), .A2(n2947), .ZN(n2912) );
  INV_X1 U3653 ( .A(n4238), .ZN(n3251) );
  NAND2_X1 U3654 ( .A1(n3251), .A2(n3214), .ZN(n2913) );
  INV_X1 U3655 ( .A(n3238), .ZN(n3217) );
  NAND2_X1 U3656 ( .A1(n3217), .A2(n3615), .ZN(n3880) );
  NAND2_X1 U3657 ( .A1(n3238), .A2(n3622), .ZN(n3877) );
  NAND2_X1 U3658 ( .A1(n3217), .A2(n3622), .ZN(n2914) );
  NAND2_X1 U3659 ( .A1(n3619), .A2(n2914), .ZN(n3225) );
  NAND2_X1 U3660 ( .A1(n3624), .A2(n3229), .ZN(n2915) );
  NAND2_X1 U3661 ( .A1(n4237), .A2(n3241), .ZN(n2916) );
  NAND2_X1 U3662 ( .A1(n3300), .A2(n3332), .ZN(n3887) );
  NAND2_X1 U3663 ( .A1(n4236), .A2(n3326), .ZN(n3889) );
  NAND2_X1 U3664 ( .A1(n2918), .A2(n2917), .ZN(n3340) );
  NAND2_X1 U3665 ( .A1(n4236), .A2(n3332), .ZN(n2919) );
  NAND2_X1 U3666 ( .A1(n3340), .A2(n2919), .ZN(n3320) );
  NAND2_X1 U3667 ( .A1(n3390), .A2(n3351), .ZN(n2920) );
  NAND2_X1 U3668 ( .A1(n3320), .A2(n2920), .ZN(n2922) );
  INV_X1 U3669 ( .A(n3390), .ZN(n3309) );
  NAND2_X1 U3670 ( .A1(n3309), .A2(n2990), .ZN(n2921) );
  INV_X1 U3671 ( .A(n3481), .ZN(n3316) );
  NAND2_X1 U3672 ( .A1(n3316), .A2(n3369), .ZN(n2923) );
  NAND2_X1 U3673 ( .A1(n3409), .A2(n3435), .ZN(n3405) );
  INV_X1 U3674 ( .A(n3409), .ZN(n3497) );
  NAND2_X1 U3675 ( .A1(n3497), .A2(n3443), .ZN(n3407) );
  NAND2_X1 U3676 ( .A1(n3409), .A2(n3443), .ZN(n2924) );
  NAND2_X1 U3677 ( .A1(n3432), .A2(n2924), .ZN(n3420) );
  NAND2_X1 U3678 ( .A1(n3782), .A2(n2927), .ZN(n3800) );
  NAND2_X1 U3679 ( .A1(n3942), .A2(n3585), .ZN(n3808) );
  NAND2_X1 U3680 ( .A1(n3800), .A2(n3808), .ZN(n3549) );
  NAND2_X1 U3681 ( .A1(n3941), .A2(n3785), .ZN(n2928) );
  NAND2_X1 U3682 ( .A1(n3779), .A2(n3594), .ZN(n3906) );
  INV_X1 U3683 ( .A(n3779), .ZN(n4544) );
  NAND2_X1 U3684 ( .A1(n4544), .A2(n3705), .ZN(n3802) );
  NAND2_X1 U3685 ( .A1(n3906), .A2(n3802), .ZN(n3591) );
  NAND2_X1 U3686 ( .A1(n3590), .A2(n2396), .ZN(n4538) );
  NAND2_X1 U3687 ( .A1(n4529), .A2(n4549), .ZN(n2930) );
  INV_X1 U3688 ( .A(n4549), .ZN(n3714) );
  AOI21_X1 U3689 ( .B1(n4538), .B2(n2930), .A(n2929), .ZN(n4513) );
  NAND2_X1 U3690 ( .A1(n4542), .A2(n4524), .ZN(n4493) );
  NAND2_X1 U3691 ( .A1(n3939), .A2(n4517), .ZN(n4494) );
  NAND2_X1 U3692 ( .A1(n4493), .A2(n4494), .ZN(n4515) );
  NAND2_X1 U3693 ( .A1(n4526), .A2(n3665), .ZN(n2933) );
  INV_X1 U3694 ( .A(n4481), .ZN(n4472) );
  NAND2_X1 U3695 ( .A1(n4423), .A2(n4445), .ZN(n2965) );
  NAND2_X1 U3696 ( .A1(n4454), .A2(n3746), .ZN(n2964) );
  NAND2_X1 U3697 ( .A1(n4432), .A2(n2935), .ZN(n4411) );
  NAND2_X1 U3698 ( .A1(n4440), .A2(n4425), .ZN(n2936) );
  NAND2_X1 U3699 ( .A1(n4420), .A2(n3726), .ZN(n2938) );
  NOR2_X1 U3700 ( .A1(n4420), .A2(n3726), .ZN(n2937) );
  AOI21_X1 U3701 ( .B1(n4391), .B2(n2938), .A(n2937), .ZN(n4372) );
  INV_X1 U3702 ( .A(n4398), .ZN(n4359) );
  NAND2_X1 U3703 ( .A1(n4359), .A2(n4382), .ZN(n2939) );
  INV_X1 U3704 ( .A(n4382), .ZN(n4377) );
  NAND2_X1 U3705 ( .A1(n3865), .A2(n2968), .ZN(n2940) );
  NOR2_X1 U3706 ( .A1(n4326), .A2(n2992), .ZN(n4312) );
  XNOR2_X1 U3707 ( .A(n3191), .B(n2941), .ZN(n2942) );
  NAND2_X1 U3708 ( .A1(n2942), .A2(n4307), .ZN(n4479) );
  NAND2_X1 U3709 ( .A1(n2463), .A2(n3645), .ZN(n3866) );
  OR2_X1 U3710 ( .A1(n2943), .A2(n3866), .ZN(n2945) );
  NAND2_X1 U3711 ( .A1(n2945), .A2(n3870), .ZN(n3249) );
  NAND2_X1 U3712 ( .A1(n3249), .A2(n3829), .ZN(n3248) );
  NAND2_X1 U3713 ( .A1(n3248), .A2(n3871), .ZN(n3199) );
  NAND2_X1 U3714 ( .A1(n3251), .A2(n2947), .ZN(n3876) );
  NAND2_X1 U3715 ( .A1(n4238), .A2(n3214), .ZN(n3873) );
  AND2_X1 U3716 ( .A1(n3876), .A2(n3873), .ZN(n3831) );
  NAND2_X1 U3717 ( .A1(n3199), .A2(n3831), .ZN(n2948) );
  INV_X1 U3718 ( .A(n3877), .ZN(n2949) );
  NAND2_X1 U3719 ( .A1(n3624), .A2(n3241), .ZN(n3884) );
  AND2_X1 U3720 ( .A1(n4237), .A2(n3229), .ZN(n3220) );
  NAND2_X1 U3721 ( .A1(n3331), .A2(n2355), .ZN(n3882) );
  NAND2_X1 U3722 ( .A1(n3267), .A2(n3882), .ZN(n2950) );
  NAND2_X1 U3723 ( .A1(n2356), .A2(n3303), .ZN(n3886) );
  INV_X1 U3724 ( .A(n3887), .ZN(n2951) );
  NAND2_X1 U3725 ( .A1(n3390), .A2(n2990), .ZN(n3893) );
  NAND2_X1 U3726 ( .A1(n3309), .A2(n3351), .ZN(n3888) );
  NAND2_X1 U3727 ( .A1(n2952), .A2(n3888), .ZN(n3363) );
  AND2_X1 U3728 ( .A1(n3481), .A2(n3369), .ZN(n3362) );
  NAND2_X1 U3729 ( .A1(n3316), .A2(n3392), .ZN(n3892) );
  NAND2_X1 U3730 ( .A1(n3364), .A2(n3483), .ZN(n3897) );
  NAND2_X1 U3731 ( .A1(n3437), .A2(n3377), .ZN(n3900) );
  NAND2_X1 U3732 ( .A1(n4235), .A2(n3499), .ZN(n3518) );
  NAND2_X1 U3733 ( .A1(n3583), .A2(n2955), .ZN(n3513) );
  NAND2_X1 U3734 ( .A1(n3518), .A2(n3513), .ZN(n2954) );
  INV_X1 U3735 ( .A(n3407), .ZN(n2953) );
  NOR2_X1 U3736 ( .A1(n2954), .A2(n2953), .ZN(n3898) );
  NAND2_X1 U3737 ( .A1(n3431), .A2(n3898), .ZN(n2958) );
  NAND2_X1 U3738 ( .A1(n3539), .A2(n3414), .ZN(n3520) );
  NAND2_X1 U3739 ( .A1(n3405), .A2(n3520), .ZN(n2957) );
  INV_X1 U3740 ( .A(n2954), .ZN(n2956) );
  NOR2_X1 U3741 ( .A1(n3583), .A2(n2955), .ZN(n3514) );
  AOI21_X1 U3742 ( .B1(n2957), .B2(n2956), .A(n3514), .ZN(n3902) );
  NAND2_X1 U3743 ( .A1(n2958), .A2(n3902), .ZN(n3801) );
  INV_X1 U3744 ( .A(n3549), .ZN(n3824) );
  NAND2_X1 U3745 ( .A1(n3801), .A2(n3824), .ZN(n2959) );
  NAND2_X1 U3746 ( .A1(n2959), .A2(n3800), .ZN(n3561) );
  NAND2_X1 U3747 ( .A1(n3603), .A2(n3785), .ZN(n3804) );
  NAND2_X1 U3748 ( .A1(n3941), .A2(n3566), .ZN(n3807) );
  NAND2_X1 U3749 ( .A1(n3804), .A2(n3807), .ZN(n3559) );
  NAND2_X1 U3750 ( .A1(n3562), .A2(n3807), .ZN(n3599) );
  INV_X1 U3751 ( .A(n3591), .ZN(n3842) );
  NAND2_X1 U3752 ( .A1(n4526), .A2(n4506), .ZN(n3847) );
  AND2_X1 U3753 ( .A1(n4494), .A2(n3847), .ZN(n2960) );
  NAND2_X1 U3754 ( .A1(n3940), .A2(n4549), .ZN(n4490) );
  NAND2_X1 U3755 ( .A1(n2960), .A2(n4490), .ZN(n3809) );
  NAND2_X1 U3756 ( .A1(n4529), .A2(n3714), .ZN(n4491) );
  NAND2_X1 U3757 ( .A1(n4493), .A2(n4491), .ZN(n2961) );
  NOR2_X1 U3758 ( .A1(n4526), .A2(n4506), .ZN(n3848) );
  AOI21_X1 U3759 ( .B1(n2961), .B2(n2960), .A(n3848), .ZN(n4468) );
  NAND2_X1 U3760 ( .A1(n4498), .A2(n4472), .ZN(n2962) );
  NAND2_X1 U3761 ( .A1(n4455), .A2(n4481), .ZN(n3811) );
  INV_X1 U3762 ( .A(n2965), .ZN(n4415) );
  NOR2_X1 U3763 ( .A1(n4473), .A2(n4459), .ZN(n4412) );
  NOR2_X1 U3764 ( .A1(n4415), .A2(n4412), .ZN(n3914) );
  NAND2_X1 U3765 ( .A1(n3724), .A2(n4425), .ZN(n3845) );
  AND2_X1 U3766 ( .A1(n3845), .A2(n2964), .ZN(n3918) );
  AND2_X1 U3767 ( .A1(n4473), .A2(n4459), .ZN(n4414) );
  NAND2_X1 U3768 ( .A1(n2965), .A2(n4414), .ZN(n2966) );
  NAND2_X1 U3769 ( .A1(n3918), .A2(n2966), .ZN(n3814) );
  OR2_X1 U3770 ( .A1(n4420), .A2(n4403), .ZN(n3846) );
  NAND2_X1 U3771 ( .A1(n4440), .A2(n4419), .ZN(n4392) );
  NAND2_X1 U3772 ( .A1(n3846), .A2(n4392), .ZN(n3916) );
  OR2_X1 U3773 ( .A1(n4378), .A2(n4365), .ZN(n3839) );
  OR2_X1 U3774 ( .A1(n4398), .A2(n4382), .ZN(n4355) );
  NAND2_X1 U3775 ( .A1(n3839), .A2(n4355), .ZN(n3915) );
  INV_X1 U3776 ( .A(n3915), .ZN(n2967) );
  NAND2_X1 U3777 ( .A1(n4398), .A2(n4382), .ZN(n3840) );
  NAND2_X1 U3778 ( .A1(n4420), .A2(n4403), .ZN(n4374) );
  AND2_X1 U3779 ( .A1(n3840), .A2(n4374), .ZN(n4354) );
  NAND2_X1 U3780 ( .A1(n4378), .A2(n4365), .ZN(n3838) );
  OAI21_X1 U3781 ( .B1(n3915), .B2(n4354), .A(n3838), .ZN(n3920) );
  XNOR2_X1 U3782 ( .A(n4361), .B(n4347), .ZN(n4340) );
  NOR2_X1 U3783 ( .A1(n4361), .A2(n2968), .ZN(n3799) );
  XNOR2_X1 U3784 ( .A(n4315), .B(n4327), .ZN(n2981) );
  NAND2_X1 U3785 ( .A1(n4688), .A2(n4691), .ZN(n2970) );
  NAND2_X1 U3786 ( .A1(n4690), .A2(n4689), .ZN(n2969) );
  OR2_X1 U3787 ( .A1(n4311), .A2(n2972), .ZN(n2978) );
  INV_X1 U3788 ( .A(REG1_REG_29__SCAN_IN), .ZN(n4033) );
  NAND2_X1 U3789 ( .A1(n2700), .A2(REG2_REG_29__SCAN_IN), .ZN(n2974) );
  NAND2_X1 U3790 ( .A1(n2158), .A2(REG0_REG_29__SCAN_IN), .ZN(n2973) );
  OAI211_X1 U3791 ( .C1(n2975), .C2(n4033), .A(n2974), .B(n2973), .ZN(n2976)
         );
  INV_X1 U3792 ( .A(n2976), .ZN(n2977) );
  NAND2_X1 U3793 ( .A1(n2978), .A2(n2977), .ZN(n3859) );
  AOI22_X1 U3794 ( .A1(n3859), .A2(n4525), .B1(n4576), .B2(n2992), .ZN(n2979)
         );
  OAI21_X1 U3795 ( .B1(n3865), .B2(n4528), .A(n2979), .ZN(n2980) );
  AOI21_X1 U3796 ( .B1(n2981), .B2(n4531), .A(n2980), .ZN(n3633) );
  OAI21_X1 U3797 ( .B1(n3640), .B2(n4638), .A(n3633), .ZN(n2996) );
  OR3_X1 U3798 ( .A1(n3181), .A2(n3182), .A3(n2982), .ZN(n2983) );
  AOI21_X1 U3799 ( .B1(n3038), .B2(n2984), .A(n2983), .ZN(n2988) );
  OAI21_X1 U3800 ( .B1(n2986), .B2(D_REG_1__SCAN_IN), .A(n2985), .ZN(n2987) );
  INV_X1 U3801 ( .A(n2989), .ZN(n2993) );
  NAND2_X1 U3802 ( .A1(n3147), .A2(n3152), .ZN(n3258) );
  NOR2_X1 U3803 ( .A1(n3258), .A2(n3257), .ZN(n3256) );
  NAND2_X1 U3804 ( .A1(n3256), .A2(n3214), .ZN(n3613) );
  OAI21_X1 U3805 ( .B1(n4346), .B2(n4325), .A(n2180), .ZN(n3636) );
  NAND2_X1 U3806 ( .A1(n2993), .A2(n2391), .ZN(U3546) );
  INV_X1 U3807 ( .A(n2997), .ZN(n2998) );
  NAND2_X1 U3808 ( .A1(n2998), .A2(n2390), .ZN(U3514) );
  NAND2_X1 U3809 ( .A1(n3000), .A2(n2999), .ZN(n3021) );
  OAI22_X1 U3810 ( .A1(n4326), .A2(n2792), .B1(n4325), .B2(n2477), .ZN(n3002)
         );
  XNOR2_X1 U3811 ( .A(n3002), .B(n3001), .ZN(n3005) );
  OAI22_X1 U3812 ( .A1(n4326), .A2(n3003), .B1(n4325), .B2(n2792), .ZN(n3004)
         );
  XNOR2_X1 U3813 ( .A(n3005), .B(n3004), .ZN(n3013) );
  NAND2_X1 U3814 ( .A1(n3013), .A2(n3757), .ZN(n3006) );
  INV_X1 U3815 ( .A(n3013), .ZN(n3010) );
  INV_X1 U3816 ( .A(n3007), .ZN(n3008) );
  NAND2_X1 U3817 ( .A1(n3009), .A2(n3008), .ZN(n3011) );
  INV_X1 U3818 ( .A(n3011), .ZN(n3012) );
  NAND3_X1 U3819 ( .A1(n3013), .A2(n3757), .A3(n3012), .ZN(n3019) );
  OAI22_X1 U3820 ( .A1(n3769), .A2(n4325), .B1(STATE_REG_SCAN_IN), .B2(n3014), 
        .ZN(n3017) );
  INV_X1 U3821 ( .A(n3859), .ZN(n3015) );
  OAI22_X1 U3822 ( .A1(n3865), .A2(n3781), .B1(n3015), .B2(n3780), .ZN(n3016)
         );
  AOI211_X1 U3823 ( .C1(n3634), .C2(n3787), .A(n3017), .B(n3016), .ZN(n3018)
         );
  NAND2_X1 U3824 ( .A1(n3019), .A2(n3018), .ZN(n3020) );
  AOI21_X1 U3825 ( .B1(n3021), .B2(n2393), .A(n3020), .ZN(n3022) );
  NAND2_X1 U3826 ( .A1(n3023), .A2(n3022), .ZN(U3217) );
  INV_X2 U3827 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X2 U3828 ( .A(n4240), .ZN(U4043) );
  INV_X1 U3829 ( .A(n3480), .ZN(n4292) );
  NAND2_X1 U3830 ( .A1(n4292), .A2(STATE_REG_SCAN_IN), .ZN(n3025) );
  OAI21_X1 U3831 ( .B1(STATE_REG_SCAN_IN), .B2(n2678), .A(n3025), .ZN(U3339)
         );
  INV_X1 U3832 ( .A(DATAI_25_), .ZN(n4065) );
  INV_X1 U3833 ( .A(n3026), .ZN(n3027) );
  NAND2_X1 U3834 ( .A1(n3027), .A2(STATE_REG_SCAN_IN), .ZN(n3028) );
  OAI21_X1 U3835 ( .B1(STATE_REG_SCAN_IN), .B2(n4065), .A(n3028), .ZN(U3327)
         );
  INV_X1 U3836 ( .A(IR_REG_30__SCAN_IN), .ZN(n4032) );
  NAND3_X1 U3837 ( .A1(IR_REG_31__SCAN_IN), .A2(STATE_REG_SCAN_IN), .A3(n4032), 
        .ZN(n3030) );
  INV_X1 U3838 ( .A(DATAI_31_), .ZN(n3029) );
  OAI22_X1 U3839 ( .A1(n2389), .A2(n3030), .B1(STATE_REG_SCAN_IN), .B2(n3029), 
        .ZN(U3321) );
  INV_X1 U3840 ( .A(DATAI_29_), .ZN(n3033) );
  NAND2_X1 U3841 ( .A1(n3031), .A2(STATE_REG_SCAN_IN), .ZN(n3032) );
  OAI21_X1 U3842 ( .B1(STATE_REG_SCAN_IN), .B2(n3033), .A(n3032), .ZN(U3323)
         );
  INV_X1 U3843 ( .A(DATAI_27_), .ZN(n3037) );
  XNOR2_X1 U3844 ( .A(n3035), .B(n3034), .ZN(n4318) );
  INV_X1 U3845 ( .A(n4318), .ZN(n3050) );
  NAND2_X1 U3846 ( .A1(n3050), .A2(STATE_REG_SCAN_IN), .ZN(n3036) );
  OAI21_X1 U3847 ( .B1(STATE_REG_SCAN_IN), .B2(n3037), .A(n3036), .ZN(U3325)
         );
  INV_X1 U3848 ( .A(D_REG_0__SCAN_IN), .ZN(n4050) );
  INV_X1 U3849 ( .A(n3039), .ZN(n3040) );
  AOI22_X1 U3850 ( .A1(n4842), .A2(n4050), .B1(n3040), .B2(n4843), .ZN(U3458)
         );
  AOI22_X1 U3851 ( .A1(n4842), .A2(n3042), .B1(n3041), .B2(n4843), .ZN(U3459)
         );
  AOI222_X1 U3852 ( .A1(n2700), .A2(REG2_REG_30__SCAN_IN), .B1(n3793), .B2(
        REG1_REG_30__SCAN_IN), .C1(n2158), .C2(REG0_REG_30__SCAN_IN), .ZN(
        n4320) );
  NAND2_X1 U3853 ( .A1(n4240), .A2(DATAO_REG_30__SCAN_IN), .ZN(n3043) );
  OAI21_X1 U3854 ( .B1(n4320), .B2(n4240), .A(n3043), .ZN(U3580) );
  OR2_X1 U3855 ( .A1(n3044), .A2(U3149), .ZN(n3936) );
  NAND2_X1 U3856 ( .A1(n3182), .A2(n3936), .ZN(n3049) );
  INV_X1 U3857 ( .A(n3049), .ZN(n3047) );
  NAND2_X1 U3858 ( .A1(n3045), .A2(n3044), .ZN(n3046) );
  INV_X1 U3859 ( .A(n3078), .ZN(n3077) );
  OAI21_X1 U3860 ( .B1(n3050), .B2(REG1_REG_0__SCAN_IN), .A(n2419), .ZN(n3051)
         );
  OAI21_X1 U3861 ( .B1(REG2_REG_0__SCAN_IN), .B2(n4318), .A(n4250), .ZN(n4254)
         );
  MUX2_X1 U3862 ( .A(n3051), .B(n2419), .S(n4254), .Z(n3053) );
  INV_X1 U3863 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3052) );
  OAI22_X1 U3864 ( .A1(n3077), .A2(n3053), .B1(STATE_REG_SCAN_IN), .B2(n3052), 
        .ZN(n3055) );
  NOR3_X1 U3865 ( .A1(n4797), .A2(REG1_REG_0__SCAN_IN), .A3(n2419), .ZN(n3054)
         );
  AOI211_X1 U3866 ( .C1(n4775), .C2(ADDR_REG_0__SCAN_IN), .A(n3055), .B(n3054), 
        .ZN(n3056) );
  INV_X1 U3867 ( .A(n3056), .ZN(U3240) );
  XNOR2_X1 U3868 ( .A(n4698), .B(REG1_REG_2__SCAN_IN), .ZN(n4260) );
  INV_X1 U3869 ( .A(n4260), .ZN(n3059) );
  XNOR2_X1 U3870 ( .A(n4699), .B(n3057), .ZN(n4245) );
  AND2_X1 U3871 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n4244)
         );
  NAND2_X1 U3872 ( .A1(n4245), .A2(n4244), .ZN(n4243) );
  NAND2_X1 U3873 ( .A1(n4699), .A2(REG1_REG_1__SCAN_IN), .ZN(n3058) );
  NAND2_X1 U3874 ( .A1(n4243), .A2(n3058), .ZN(n4259) );
  NAND2_X1 U3875 ( .A1(n3059), .A2(n4259), .ZN(n3061) );
  NAND2_X1 U3876 ( .A1(n4698), .A2(REG1_REG_2__SCAN_IN), .ZN(n3060) );
  NAND2_X1 U3877 ( .A1(n3061), .A2(n3060), .ZN(n3062) );
  XNOR2_X1 U3878 ( .A(n3062), .B(n2281), .ZN(n3101) );
  NAND2_X1 U3879 ( .A1(n3101), .A2(REG1_REG_3__SCAN_IN), .ZN(n3064) );
  NAND2_X1 U3880 ( .A1(n3062), .A2(n4697), .ZN(n3063) );
  NAND2_X1 U3881 ( .A1(n3066), .A2(n4696), .ZN(n3067) );
  MUX2_X1 U3882 ( .A(n3068), .B(REG1_REG_5__SCAN_IN), .S(n3124), .Z(n3129) );
  NAND2_X1 U3883 ( .A1(n3128), .A2(n3129), .ZN(n3127) );
  OR2_X1 U3884 ( .A1(n3124), .A2(n3068), .ZN(n3069) );
  NAND2_X1 U3885 ( .A1(n3127), .A2(n3069), .ZN(n3092) );
  XNOR2_X1 U3886 ( .A(n3092), .B(n3080), .ZN(n3091) );
  XNOR2_X1 U3887 ( .A(n3091), .B(REG1_REG_6__SCAN_IN), .ZN(n3084) );
  INV_X1 U3888 ( .A(n3124), .ZN(n4695) );
  INV_X1 U3889 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3075) );
  INV_X1 U3890 ( .A(n4698), .ZN(n3074) );
  INV_X1 U3891 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3070) );
  INV_X1 U3892 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3071) );
  NOR3_X1 U3893 ( .A1(n3072), .A2(n3071), .A3(n2419), .ZN(n4241) );
  NOR2_X1 U3894 ( .A1(n2476), .A2(n3070), .ZN(n4262) );
  MUX2_X1 U3895 ( .A(REG2_REG_2__SCAN_IN), .B(n3075), .S(n4698), .Z(n3073) );
  OAI21_X1 U3896 ( .B1(n4241), .B2(n4262), .A(n3073), .ZN(n4267) );
  OAI21_X1 U3897 ( .B1(n3075), .B2(n3074), .A(n4267), .ZN(n3076) );
  INV_X1 U3898 ( .A(REG2_REG_5__SCAN_IN), .ZN(n4069) );
  MUX2_X1 U3899 ( .A(REG2_REG_5__SCAN_IN), .B(n4069), .S(n3124), .Z(n3121) );
  NOR2_X1 U3900 ( .A1(n3122), .A2(n3121), .ZN(n3120) );
  AOI21_X1 U3901 ( .B1(n4695), .B2(REG2_REG_5__SCAN_IN), .A(n3120), .ZN(n3087)
         );
  XOR2_X1 U3902 ( .A(REG2_REG_6__SCAN_IN), .B(n3088), .Z(n3082) );
  OR2_X1 U3903 ( .A1(n4701), .A2(n4318), .ZN(n4251) );
  NOR2_X2 U3904 ( .A1(n3077), .A2(n4251), .ZN(n4809) );
  AND2_X1 U3905 ( .A1(n3078), .A2(n4701), .ZN(n4758) );
  INV_X1 U3906 ( .A(n4758), .ZN(n4812) );
  INV_X1 U3907 ( .A(REG3_REG_6__SCAN_IN), .ZN(n4084) );
  NOR2_X1 U3908 ( .A1(STATE_REG_SCAN_IN), .A2(n4084), .ZN(n3302) );
  AOI21_X1 U3909 ( .B1(n4775), .B2(ADDR_REG_6__SCAN_IN), .A(n3302), .ZN(n3079)
         );
  OAI21_X1 U3910 ( .B1(n4812), .B2(n3080), .A(n3079), .ZN(n3081) );
  AOI21_X1 U3911 ( .B1(n3082), .B2(n4809), .A(n3081), .ZN(n3083) );
  OAI21_X1 U3912 ( .B1(n3084), .B2(n4797), .A(n3083), .ZN(U3246) );
  NOR2_X1 U3913 ( .A1(n4775), .A2(U4043), .ZN(U3148) );
  INV_X1 U3914 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n3086) );
  NAND2_X1 U3915 ( .A1(n3724), .A2(U4043), .ZN(n3085) );
  OAI21_X1 U3916 ( .B1(U4043), .B2(n3086), .A(n3085), .ZN(U3573) );
  INV_X1 U3917 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3955) );
  MUX2_X1 U3918 ( .A(n3955), .B(REG2_REG_7__SCAN_IN), .S(n4693), .Z(n3159) );
  XNOR2_X1 U3919 ( .A(n3452), .B(n4692), .ZN(n3454) );
  XOR2_X1 U3920 ( .A(REG2_REG_8__SCAN_IN), .B(n3454), .Z(n3099) );
  INV_X1 U3921 ( .A(n4809), .ZN(n4751) );
  NAND2_X1 U3922 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3349) );
  INV_X1 U3923 ( .A(n3349), .ZN(n3090) );
  NOR2_X1 U3924 ( .A1(n4812), .A2(n4692), .ZN(n3089) );
  AOI211_X1 U3925 ( .C1(n4775), .C2(ADDR_REG_8__SCAN_IN), .A(n3090), .B(n3089), 
        .ZN(n3098) );
  NAND2_X1 U3926 ( .A1(n3091), .A2(REG1_REG_6__SCAN_IN), .ZN(n3094) );
  NAND2_X1 U3927 ( .A1(n3092), .A2(n4694), .ZN(n3093) );
  NAND2_X1 U3928 ( .A1(n3094), .A2(n3093), .ZN(n3155) );
  AND2_X1 U3929 ( .A1(n4693), .A2(REG1_REG_7__SCAN_IN), .ZN(n3095) );
  OR2_X1 U3930 ( .A1(n4693), .A2(REG1_REG_7__SCAN_IN), .ZN(n3096) );
  OAI211_X1 U3931 ( .C1(n2195), .C2(REG1_REG_8__SCAN_IN), .A(n3464), .B(n4794), 
        .ZN(n3097) );
  OAI211_X1 U3932 ( .C1(n3099), .C2(n4751), .A(n3098), .B(n3097), .ZN(U3248)
         );
  INV_X1 U3933 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3206) );
  XNOR2_X1 U3934 ( .A(n3100), .B(n3206), .ZN(n3103) );
  XOR2_X1 U3935 ( .A(n3101), .B(REG1_REG_3__SCAN_IN), .Z(n3102) );
  AOI22_X1 U3936 ( .A1(n4809), .A2(n3103), .B1(n4794), .B2(n3102), .ZN(n3105)
         );
  AOI22_X1 U3937 ( .A1(n4775), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n3104) );
  OAI211_X1 U3938 ( .C1(n2281), .C2(n4812), .A(n3105), .B(n3104), .ZN(U3243)
         );
  INV_X1 U3939 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n3107) );
  NAND2_X1 U3940 ( .A1(n3364), .A2(U4043), .ZN(n3106) );
  OAI21_X1 U3941 ( .B1(U4043), .B2(n3107), .A(n3106), .ZN(U3560) );
  INV_X1 U3942 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n3109) );
  NAND2_X1 U3943 ( .A1(n3497), .A2(U4043), .ZN(n3108) );
  OAI21_X1 U3944 ( .B1(U4043), .B2(n3109), .A(n3108), .ZN(U3561) );
  INV_X1 U3945 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n3111) );
  NAND2_X1 U3946 ( .A1(n3331), .A2(U4043), .ZN(n3110) );
  OAI21_X1 U3947 ( .B1(U4043), .B2(n3111), .A(n3110), .ZN(U3556) );
  INV_X1 U3948 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n3113) );
  NAND2_X1 U3949 ( .A1(n3583), .A2(U4043), .ZN(n3112) );
  OAI21_X1 U3950 ( .B1(U4043), .B2(n3113), .A(n3112), .ZN(U3563) );
  INV_X1 U3951 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n3115) );
  NAND2_X1 U3952 ( .A1(n3309), .A2(U4043), .ZN(n3114) );
  OAI21_X1 U3953 ( .B1(U4043), .B2(n3115), .A(n3114), .ZN(U3558) );
  INV_X1 U3954 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n3117) );
  NAND2_X1 U3955 ( .A1(n3672), .A2(U4043), .ZN(n3116) );
  OAI21_X1 U3956 ( .B1(U4043), .B2(n3117), .A(n3116), .ZN(U3552) );
  INV_X1 U3957 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n3119) );
  NAND2_X1 U3958 ( .A1(n4378), .A2(U4043), .ZN(n3118) );
  OAI21_X1 U3959 ( .B1(U4043), .B2(n3119), .A(n3118), .ZN(U3576) );
  AOI211_X1 U3960 ( .C1(n3122), .C2(n3121), .A(n3120), .B(n4751), .ZN(n3126)
         );
  INV_X1 U3961 ( .A(REG3_REG_5__SCAN_IN), .ZN(n3958) );
  NOR2_X1 U3962 ( .A1(STATE_REG_SCAN_IN), .A2(n3958), .ZN(n3240) );
  AOI21_X1 U3963 ( .B1(n4775), .B2(ADDR_REG_5__SCAN_IN), .A(n3240), .ZN(n3123)
         );
  OAI21_X1 U3964 ( .B1(n4812), .B2(n3124), .A(n3123), .ZN(n3125) );
  NOR2_X1 U3965 ( .A1(n3126), .A2(n3125), .ZN(n3131) );
  OAI211_X1 U3966 ( .C1(n3129), .C2(n3128), .A(n4794), .B(n3127), .ZN(n3130)
         );
  NAND2_X1 U3967 ( .A1(n3131), .A2(n3130), .ZN(U3245) );
  INV_X1 U3968 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n3133) );
  NAND2_X1 U3969 ( .A1(n3217), .A2(U4043), .ZN(n3132) );
  OAI21_X1 U3970 ( .B1(U4043), .B2(n3133), .A(n3132), .ZN(U3554) );
  INV_X1 U3971 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n3135) );
  NAND2_X1 U3972 ( .A1(n3481), .A2(U4043), .ZN(n3134) );
  OAI21_X1 U3973 ( .B1(U4043), .B2(n3135), .A(n3134), .ZN(U3559) );
  INV_X1 U3974 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n3137) );
  NAND2_X1 U3975 ( .A1(n4398), .A2(U4043), .ZN(n3136) );
  OAI21_X1 U3976 ( .B1(U4043), .B2(n3137), .A(n3136), .ZN(U3575) );
  OR2_X1 U3977 ( .A1(n2943), .A2(n3138), .ZN(n3139) );
  NAND2_X1 U3978 ( .A1(n3140), .A2(n3139), .ZN(n3189) );
  NAND2_X1 U3979 ( .A1(n2904), .A2(n4576), .ZN(n3142) );
  NAND2_X1 U3980 ( .A1(n2944), .A2(n4545), .ZN(n3141) );
  OAI211_X1 U3981 ( .C1(n2908), .C2(n4541), .A(n3142), .B(n3141), .ZN(n3143)
         );
  INV_X1 U3982 ( .A(n3143), .ZN(n3146) );
  XNOR2_X1 U3983 ( .A(n2943), .B(n3866), .ZN(n3144) );
  NAND2_X1 U3984 ( .A1(n3144), .A2(n4531), .ZN(n3145) );
  OAI211_X1 U3985 ( .C1(n3189), .C2(n4479), .A(n3146), .B(n3145), .ZN(n3187)
         );
  INV_X1 U3986 ( .A(n4636), .ZN(n4894) );
  OAI21_X1 U3987 ( .B1(n3152), .B2(n3147), .A(n3258), .ZN(n3196) );
  OAI22_X1 U3988 ( .A1(n3189), .A2(n3255), .B1(n4894), .B2(n3196), .ZN(n3148)
         );
  NOR2_X1 U3989 ( .A1(n3187), .A2(n3148), .ZN(n4866) );
  NAND2_X1 U3990 ( .A1(n4908), .A2(REG1_REG_1__SCAN_IN), .ZN(n3149) );
  OAI21_X1 U3991 ( .B1(n4866), .B2(n4908), .A(n3149), .ZN(U3519) );
  INV_X1 U3992 ( .A(n3255), .ZN(n4899) );
  NAND2_X1 U3993 ( .A1(n2944), .A2(n3152), .ZN(n3868) );
  NAND2_X1 U3994 ( .A1(n3866), .A2(n3868), .ZN(n4827) );
  INV_X1 U3995 ( .A(n3150), .ZN(n3151) );
  NOR2_X1 U3996 ( .A1(n3152), .A2(n3151), .ZN(n4825) );
  INV_X1 U3997 ( .A(n4479), .ZN(n3626) );
  OAI21_X1 U3998 ( .B1(n3626), .B2(n4531), .A(n4827), .ZN(n3153) );
  OAI21_X1 U3999 ( .B1(n2905), .B2(n4541), .A(n3153), .ZN(n4823) );
  AOI211_X1 U4000 ( .C1(n4899), .C2(n4827), .A(n4825), .B(n4823), .ZN(n4864)
         );
  NAND2_X1 U4001 ( .A1(n4908), .A2(REG1_REG_0__SCAN_IN), .ZN(n3154) );
  OAI21_X1 U4002 ( .B1(n4864), .B2(n4908), .A(n3154), .ZN(U3518) );
  MUX2_X1 U4003 ( .A(n2573), .B(REG1_REG_7__SCAN_IN), .S(n4693), .Z(n3156) );
  XOR2_X1 U4004 ( .A(n3156), .B(n3155), .Z(n3164) );
  NAND2_X1 U4005 ( .A1(n4775), .A2(ADDR_REG_7__SCAN_IN), .ZN(n3157) );
  NAND2_X1 U4006 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3310) );
  NAND2_X1 U4007 ( .A1(n3157), .A2(n3310), .ZN(n3162) );
  AOI211_X1 U4008 ( .C1(n3160), .C2(n3159), .A(n4751), .B(n3158), .ZN(n3161)
         );
  AOI211_X1 U4009 ( .C1(n4758), .C2(n4693), .A(n3162), .B(n3161), .ZN(n3163)
         );
  OAI21_X1 U4010 ( .B1(n4797), .B2(n3164), .A(n3163), .ZN(U3247) );
  INV_X1 U4011 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n3166) );
  NAND2_X1 U4012 ( .A1(n3859), .A2(U4043), .ZN(n3165) );
  OAI21_X1 U4013 ( .B1(U4043), .B2(n3166), .A(n3165), .ZN(U3579) );
  INV_X1 U4014 ( .A(n3170), .ZN(n3171) );
  AOI21_X1 U4015 ( .B1(n3167), .B2(n3168), .A(n3171), .ZN(n3178) );
  AOI22_X1 U4016 ( .A1(n3725), .A2(n4239), .B1(n3257), .B2(n3784), .ZN(n3177)
         );
  INV_X1 U4017 ( .A(n3172), .ZN(n3175) );
  INV_X1 U4018 ( .A(n3182), .ZN(n3174) );
  NAND3_X1 U4019 ( .A1(n3175), .A2(n3174), .A3(n3173), .ZN(n3673) );
  AOI22_X1 U4020 ( .A1(REG3_REG_2__SCAN_IN), .A2(n3673), .B1(n3703), .B2(n4238), .ZN(n3176) );
  OAI211_X1 U4021 ( .C1(n3178), .C2(n3790), .A(n3177), .B(n3176), .ZN(U3234)
         );
  INV_X1 U4022 ( .A(DATAO_REG_28__SCAN_IN), .ZN(n3180) );
  INV_X1 U4023 ( .A(n4326), .ZN(n4342) );
  NAND2_X1 U4024 ( .A1(n4342), .A2(U4043), .ZN(n3179) );
  OAI21_X1 U4025 ( .B1(U4043), .B2(n3180), .A(n3179), .ZN(U3578) );
  NOR2_X1 U4026 ( .A1(n3182), .A2(n3181), .ZN(n3183) );
  NAND3_X1 U4027 ( .A1(n3185), .A2(n3184), .A3(n3183), .ZN(n3186) );
  NAND2_X1 U4028 ( .A1(n3186), .A2(n4519), .ZN(n3190) );
  AND2_X1 U4029 ( .A1(n3190), .A2(n4307), .ZN(n4535) );
  INV_X2 U4030 ( .A(n3190), .ZN(n4813) );
  MUX2_X1 U4031 ( .A(n3187), .B(REG2_REG_1__SCAN_IN), .S(n4813), .Z(n3188) );
  INV_X1 U4032 ( .A(n3188), .ZN(n3195) );
  INV_X1 U4033 ( .A(n3189), .ZN(n3193) );
  NAND2_X1 U4034 ( .A1(n3191), .A2(n4691), .ZN(n3226) );
  INV_X1 U4035 ( .A(n3226), .ZN(n3192) );
  AOI22_X1 U4036 ( .A1(n3193), .A2(n4828), .B1(REG3_REG_1__SCAN_IN), .B2(n4826), .ZN(n3194) );
  OAI211_X1 U4037 ( .C1(n4555), .C2(n3196), .A(n3195), .B(n3194), .ZN(U3289)
         );
  INV_X1 U4038 ( .A(n3831), .ZN(n3198) );
  XNOR2_X1 U4039 ( .A(n3197), .B(n3198), .ZN(n4869) );
  NAND2_X1 U4040 ( .A1(n4869), .A2(n3626), .ZN(n3205) );
  XNOR2_X1 U4041 ( .A(n3199), .B(n3831), .ZN(n3203) );
  OAI22_X1 U4042 ( .A1(n3238), .A2(n4541), .B1(n4565), .B2(n3214), .ZN(n3201)
         );
  NOR2_X1 U40430 ( .A1(n2908), .A2(n4528), .ZN(n3200) );
  OR2_X1 U4044 ( .A1(n3201), .A2(n3200), .ZN(n3202) );
  AOI21_X1 U4045 ( .B1(n3203), .B2(n4531), .A(n3202), .ZN(n3204) );
  AND2_X1 U4046 ( .A1(n3205), .A2(n3204), .ZN(n4871) );
  OAI22_X1 U4047 ( .A1(n4557), .A2(n3206), .B1(REG3_REG_3__SCAN_IN), .B2(n4519), .ZN(n3209) );
  OR2_X1 U4048 ( .A1(n3256), .A2(n3214), .ZN(n3207) );
  NAND2_X1 U4049 ( .A1(n3613), .A2(n3207), .ZN(n4867) );
  NOR2_X1 U4050 ( .A1(n4555), .A2(n4867), .ZN(n3208) );
  AOI211_X1 U4051 ( .C1(n4828), .C2(n4869), .A(n3209), .B(n3208), .ZN(n3210)
         );
  OAI21_X1 U4052 ( .B1(n4813), .B2(n4871), .A(n3210), .ZN(U3287) );
  NAND2_X1 U4053 ( .A1(n3170), .A2(n3212), .ZN(n3213) );
  XOR2_X1 U4054 ( .A(n3211), .B(n3213), .Z(n3219) );
  OAI22_X1 U4055 ( .A1(n3769), .A2(n3214), .B1(n3781), .B2(n2908), .ZN(n3216)
         );
  MUX2_X1 U4056 ( .A(n3787), .B(U3149), .S(REG3_REG_3__SCAN_IN), .Z(n3215) );
  AOI211_X1 U4057 ( .C1(n3703), .C2(n3217), .A(n3216), .B(n3215), .ZN(n3218)
         );
  OAI21_X1 U4058 ( .B1(n3219), .B2(n3790), .A(n3218), .ZN(U3215) );
  INV_X1 U4059 ( .A(n3220), .ZN(n3879) );
  AND2_X1 U4060 ( .A1(n3879), .A2(n3884), .ZN(n3825) );
  XOR2_X1 U4061 ( .A(n3825), .B(n3221), .Z(n3224) );
  AOI22_X1 U4062 ( .A1(n3331), .A2(n4525), .B1(n4576), .B2(n3241), .ZN(n3222)
         );
  OAI21_X1 U4063 ( .B1(n3238), .B2(n4528), .A(n3222), .ZN(n3223) );
  AOI21_X1 U4064 ( .B1(n3224), .B2(n4531), .A(n3223), .ZN(n4878) );
  XNOR2_X1 U4065 ( .A(n3225), .B(n3825), .ZN(n4881) );
  NAND2_X1 U4066 ( .A1(n4479), .A2(n3226), .ZN(n3227) );
  INV_X1 U4067 ( .A(n3614), .ZN(n3230) );
  INV_X1 U4068 ( .A(n3228), .ZN(n3272) );
  OAI21_X1 U4069 ( .B1(n3230), .B2(n3229), .A(n3272), .ZN(n4879) );
  NOR2_X1 U4070 ( .A1(n4555), .A2(n4879), .ZN(n3233) );
  INV_X1 U4071 ( .A(n3231), .ZN(n3244) );
  OAI22_X1 U4072 ( .A1(n3190), .A2(n4069), .B1(n3244), .B2(n4519), .ZN(n3232)
         );
  AOI211_X1 U4073 ( .C1(n4881), .C2(n4331), .A(n3233), .B(n3232), .ZN(n3234)
         );
  OAI21_X1 U4074 ( .B1(n4878), .B2(n4813), .A(n3234), .ZN(U3285) );
  OAI211_X1 U4075 ( .C1(n3237), .C2(n3236), .A(n3235), .B(n3757), .ZN(n3243)
         );
  OAI22_X1 U4076 ( .A1(n3238), .A2(n3781), .B1(n3780), .B2(n2356), .ZN(n3239)
         );
  AOI211_X1 U4077 ( .C1(n3241), .C2(n3784), .A(n3240), .B(n3239), .ZN(n3242)
         );
  OAI211_X1 U4078 ( .C1(n3762), .C2(n3244), .A(n3243), .B(n3242), .ZN(U3224)
         );
  INV_X1 U4079 ( .A(n3246), .ZN(n3247) );
  AOI21_X1 U4080 ( .B1(n3829), .B2(n3245), .A(n3247), .ZN(n4814) );
  OAI21_X1 U4081 ( .B1(n3829), .B2(n3249), .A(n3248), .ZN(n3254) );
  AOI22_X1 U4082 ( .A1(n4239), .A2(n4545), .B1(n3257), .B2(n4576), .ZN(n3250)
         );
  OAI21_X1 U4083 ( .B1(n3251), .B2(n4541), .A(n3250), .ZN(n3253) );
  NOR2_X1 U4084 ( .A1(n4814), .A2(n4479), .ZN(n3252) );
  AOI211_X1 U4085 ( .C1(n4531), .C2(n3254), .A(n3253), .B(n3252), .ZN(n4821)
         );
  OAI21_X1 U4086 ( .B1(n4814), .B2(n3255), .A(n4821), .ZN(n3265) );
  INV_X1 U4087 ( .A(n3256), .ZN(n3260) );
  NAND2_X1 U4088 ( .A1(n3258), .A2(n3257), .ZN(n3259) );
  NAND2_X1 U4089 ( .A1(n3260), .A2(n3259), .ZN(n4815) );
  OAI22_X1 U4090 ( .A1(n4629), .A2(n4815), .B1(n4910), .B2(n3261), .ZN(n3262)
         );
  AOI21_X1 U4091 ( .B1(n3265), .B2(n4910), .A(n3262), .ZN(n3263) );
  INV_X1 U4092 ( .A(n3263), .ZN(U3520) );
  INV_X1 U4093 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4122) );
  OAI22_X1 U4094 ( .A1(n4682), .A2(n4815), .B1(n4902), .B2(n4122), .ZN(n3264)
         );
  AOI21_X1 U4095 ( .B1(n3265), .B2(n4902), .A(n3264), .ZN(n3266) );
  INV_X1 U4096 ( .A(n3266), .ZN(U3471) );
  NAND2_X1 U4097 ( .A1(n3886), .A2(n3882), .ZN(n3851) );
  XNOR2_X1 U4098 ( .A(n3267), .B(n3851), .ZN(n3270) );
  OAI22_X1 U4099 ( .A1(n3300), .A2(n4541), .B1(n4565), .B2(n2355), .ZN(n3268)
         );
  AOI21_X1 U4100 ( .B1(n4545), .B2(n4237), .A(n3268), .ZN(n3269) );
  OAI21_X1 U4101 ( .B1(n3270), .B2(n4547), .A(n3269), .ZN(n3287) );
  INV_X1 U4102 ( .A(n3287), .ZN(n3277) );
  INV_X1 U4103 ( .A(n3333), .ZN(n3271) );
  AOI21_X1 U4104 ( .B1(n3303), .B2(n3272), .A(n3271), .ZN(n3292) );
  OAI22_X1 U4105 ( .A1(n4557), .A2(n2271), .B1(n3306), .B2(n4519), .ZN(n3273)
         );
  AOI21_X1 U4106 ( .B1(n3292), .B2(n4817), .A(n3273), .ZN(n3276) );
  XOR2_X1 U4107 ( .A(n3274), .B(n3851), .Z(n3288) );
  NAND2_X1 U4108 ( .A1(n3288), .A2(n4331), .ZN(n3275) );
  OAI211_X1 U4109 ( .C1(n3277), .C2(n4813), .A(n3276), .B(n3275), .ZN(U3284)
         );
  AOI22_X1 U4110 ( .A1(n3703), .A2(n4237), .B1(n3725), .B2(n4238), .ZN(n3278)
         );
  NAND2_X1 U4111 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n4274) );
  OAI211_X1 U4112 ( .C1(n3769), .C2(n3615), .A(n3278), .B(n4274), .ZN(n3285)
         );
  INV_X1 U4113 ( .A(n3280), .ZN(n3283) );
  INV_X1 U4114 ( .A(n3281), .ZN(n3282) );
  AOI211_X1 U4115 ( .C1(n3279), .C2(n3283), .A(n3790), .B(n3282), .ZN(n3284)
         );
  AOI211_X1 U4116 ( .C1(n3630), .C2(n3787), .A(n3285), .B(n3284), .ZN(n3286)
         );
  INV_X1 U4117 ( .A(n3286), .ZN(U3227) );
  AOI21_X1 U4118 ( .B1(n3288), .B2(n4891), .A(n3287), .ZN(n3294) );
  INV_X1 U4119 ( .A(n4682), .ZN(n4640) );
  INV_X1 U4120 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3289) );
  NOR2_X1 U4121 ( .A1(n4902), .A2(n3289), .ZN(n3290) );
  AOI21_X1 U4122 ( .B1(n3292), .B2(n4640), .A(n3290), .ZN(n3291) );
  OAI21_X1 U4123 ( .B1(n3294), .B2(n4900), .A(n3291), .ZN(U3479) );
  INV_X1 U4124 ( .A(n4629), .ZN(n4562) );
  AOI22_X1 U4125 ( .A1(n3292), .A2(n4562), .B1(n4908), .B2(REG1_REG_6__SCAN_IN), .ZN(n3293) );
  OAI21_X1 U4126 ( .B1(n3294), .B2(n4908), .A(n3293), .ZN(U3524) );
  XNOR2_X1 U4127 ( .A(n3297), .B(n3296), .ZN(n3298) );
  XNOR2_X1 U4128 ( .A(n3295), .B(n3298), .ZN(n3299) );
  NAND2_X1 U4129 ( .A1(n3299), .A2(n3757), .ZN(n3305) );
  OAI22_X1 U4130 ( .A1(n3624), .A2(n3781), .B1(n3780), .B2(n3300), .ZN(n3301)
         );
  AOI211_X1 U4131 ( .C1(n3303), .C2(n3784), .A(n3302), .B(n3301), .ZN(n3304)
         );
  OAI211_X1 U4132 ( .C1(n3762), .C2(n3306), .A(n3305), .B(n3304), .ZN(U3236)
         );
  XNOR2_X1 U4133 ( .A(n3308), .B(n3307), .ZN(n3314) );
  AOI22_X1 U4134 ( .A1(n3703), .A2(n3309), .B1(n3725), .B2(n3331), .ZN(n3311)
         );
  OAI211_X1 U4135 ( .C1(n3769), .C2(n3326), .A(n3311), .B(n3310), .ZN(n3312)
         );
  AOI21_X1 U4136 ( .B1(n3336), .B2(n3787), .A(n3312), .ZN(n3313) );
  OAI21_X1 U4137 ( .B1(n3314), .B2(n3790), .A(n3313), .ZN(U3210) );
  XNOR2_X1 U4138 ( .A(n3390), .B(n3351), .ZN(n3860) );
  XNOR2_X1 U4139 ( .A(n3315), .B(n3860), .ZN(n3319) );
  OAI22_X1 U4140 ( .A1(n3316), .A2(n4541), .B1(n4565), .B2(n3351), .ZN(n3317)
         );
  AOI21_X1 U4141 ( .B1(n4545), .B2(n4236), .A(n3317), .ZN(n3318) );
  OAI21_X1 U4142 ( .B1(n3319), .B2(n4547), .A(n3318), .ZN(n3356) );
  INV_X1 U4143 ( .A(n3356), .ZN(n3325) );
  XNOR2_X1 U4144 ( .A(n3320), .B(n3860), .ZN(n3357) );
  INV_X1 U4145 ( .A(n3334), .ZN(n3321) );
  OAI21_X1 U4146 ( .B1(n3321), .B2(n3351), .A(n2229), .ZN(n3361) );
  AOI22_X1 U4147 ( .A1(n4813), .A2(REG2_REG_8__SCAN_IN), .B1(n3353), .B2(n4826), .ZN(n3322) );
  OAI21_X1 U4148 ( .B1(n3361), .B2(n4555), .A(n3322), .ZN(n3323) );
  AOI21_X1 U4149 ( .B1(n3357), .B2(n4331), .A(n3323), .ZN(n3324) );
  OAI21_X1 U4150 ( .B1(n3325), .B2(n4813), .A(n3324), .ZN(U3282) );
  OAI22_X1 U4151 ( .A1(n3390), .A2(n4541), .B1(n3326), .B2(n4565), .ZN(n3330)
         );
  XOR2_X1 U4152 ( .A(n3827), .B(n3327), .Z(n3328) );
  NOR2_X1 U4153 ( .A1(n3328), .A2(n4547), .ZN(n3329) );
  AOI211_X1 U4154 ( .C1(n4545), .C2(n3331), .A(n3330), .B(n3329), .ZN(n4886)
         );
  AOI21_X1 U4155 ( .B1(n3333), .B2(n3332), .A(n4894), .ZN(n3335) );
  NAND2_X1 U4156 ( .A1(n3335), .A2(n3334), .ZN(n4885) );
  INV_X1 U4157 ( .A(n4885), .ZN(n3339) );
  INV_X1 U4158 ( .A(n3336), .ZN(n3337) );
  OAI22_X1 U4159 ( .A1(n4557), .A2(n3955), .B1(n3337), .B2(n4519), .ZN(n3338)
         );
  AOI21_X1 U4160 ( .B1(n3339), .B2(n4535), .A(n3338), .ZN(n3343) );
  NAND2_X1 U4161 ( .A1(n3341), .A2(n3827), .ZN(n4883) );
  NAND3_X1 U4162 ( .A1(n3340), .A2(n4883), .A3(n4331), .ZN(n3342) );
  OAI211_X1 U4163 ( .C1(n4886), .C2(n4813), .A(n3343), .B(n3342), .ZN(U3283)
         );
  INV_X1 U4164 ( .A(n3345), .ZN(n3347) );
  NOR2_X1 U4165 ( .A1(n3347), .A2(n3346), .ZN(n3348) );
  XNOR2_X1 U4166 ( .A(n3344), .B(n3348), .ZN(n3355) );
  AOI22_X1 U4167 ( .A1(n3725), .A2(n4236), .B1(n3703), .B2(n3481), .ZN(n3350)
         );
  OAI211_X1 U4168 ( .C1(n3769), .C2(n3351), .A(n3350), .B(n3349), .ZN(n3352)
         );
  AOI21_X1 U4169 ( .B1(n3353), .B2(n3787), .A(n3352), .ZN(n3354) );
  OAI21_X1 U4170 ( .B1(n3355), .B2(n3790), .A(n3354), .ZN(U3218) );
  INV_X1 U4171 ( .A(REG0_REG_8__SCAN_IN), .ZN(n4077) );
  AOI21_X1 U4172 ( .B1(n3357), .B2(n4891), .A(n3356), .ZN(n3359) );
  MUX2_X1 U4173 ( .A(n4077), .B(n3359), .S(n4902), .Z(n3358) );
  OAI21_X1 U4174 ( .B1(n3361), .B2(n4682), .A(n3358), .ZN(U3483) );
  MUX2_X1 U4175 ( .A(n2583), .B(n3359), .S(n4910), .Z(n3360) );
  OAI21_X1 U4176 ( .B1(n3361), .B2(n4629), .A(n3360), .ZN(U3526) );
  INV_X1 U4177 ( .A(n3362), .ZN(n3895) );
  NAND2_X1 U4178 ( .A1(n3895), .A2(n3892), .ZN(n3853) );
  XNOR2_X1 U4179 ( .A(n3363), .B(n3853), .ZN(n3367) );
  AOI22_X1 U4180 ( .A1(n3364), .A2(n4525), .B1(n4576), .B2(n3392), .ZN(n3365)
         );
  OAI21_X1 U4181 ( .B1(n3390), .B2(n4528), .A(n3365), .ZN(n3366) );
  AOI21_X1 U4182 ( .B1(n3367), .B2(n4531), .A(n3366), .ZN(n4888) );
  XOR2_X1 U4183 ( .A(n3853), .B(n3368), .Z(n4892) );
  NOR2_X1 U4184 ( .A1(n3370), .A2(n3369), .ZN(n3371) );
  OR2_X1 U4185 ( .A1(n3383), .A2(n3371), .ZN(n4889) );
  AOI22_X1 U4186 ( .A1(n4813), .A2(REG2_REG_9__SCAN_IN), .B1(n3393), .B2(n4826), .ZN(n3372) );
  OAI21_X1 U4187 ( .B1(n4889), .B2(n4555), .A(n3372), .ZN(n3373) );
  AOI21_X1 U4188 ( .B1(n4892), .B2(n4331), .A(n3373), .ZN(n3374) );
  OAI21_X1 U4189 ( .B1(n4813), .B2(n4888), .A(n3374), .ZN(U3281) );
  NAND2_X1 U4190 ( .A1(n3900), .A2(n3897), .ZN(n3852) );
  INV_X1 U4191 ( .A(n3852), .ZN(n3375) );
  XNOR2_X1 U4192 ( .A(n3376), .B(n3375), .ZN(n3381) );
  NAND2_X1 U4193 ( .A1(n3377), .A2(n4576), .ZN(n3379) );
  NAND2_X1 U4194 ( .A1(n3481), .A2(n4545), .ZN(n3378) );
  OAI211_X1 U4195 ( .C1(n3409), .C2(n4541), .A(n3379), .B(n3378), .ZN(n3380)
         );
  AOI21_X1 U4196 ( .B1(n3381), .B2(n4531), .A(n3380), .ZN(n3398) );
  XNOR2_X1 U4197 ( .A(n3382), .B(n3852), .ZN(n3397) );
  OR2_X1 U4198 ( .A1(n3383), .A2(n3483), .ZN(n3384) );
  NAND2_X1 U4199 ( .A1(n3441), .A2(n3384), .ZN(n3404) );
  AOI22_X1 U4200 ( .A1(n4813), .A2(REG2_REG_10__SCAN_IN), .B1(n3490), .B2(
        n4826), .ZN(n3385) );
  OAI21_X1 U4201 ( .B1(n3404), .B2(n4555), .A(n3385), .ZN(n3386) );
  AOI21_X1 U4202 ( .B1(n3397), .B2(n4331), .A(n3386), .ZN(n3387) );
  OAI21_X1 U4203 ( .B1(n3398), .B2(n4813), .A(n3387), .ZN(U3280) );
  XOR2_X1 U4204 ( .A(n3388), .B(n3389), .Z(n3396) );
  AND2_X1 U4205 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4712) );
  OAI22_X1 U4206 ( .A1(n3390), .A2(n3781), .B1(n3780), .B2(n3437), .ZN(n3391)
         );
  AOI211_X1 U4207 ( .C1(n3392), .C2(n3784), .A(n4712), .B(n3391), .ZN(n3395)
         );
  NAND2_X1 U4208 ( .A1(n3787), .A2(n3393), .ZN(n3394) );
  OAI211_X1 U4209 ( .C1(n3396), .C2(n3790), .A(n3395), .B(n3394), .ZN(U3228)
         );
  NAND2_X1 U4210 ( .A1(n3397), .A2(n4891), .ZN(n3399) );
  AND2_X1 U4211 ( .A1(n3399), .A2(n3398), .ZN(n3402) );
  INV_X1 U4212 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3400) );
  MUX2_X1 U4213 ( .A(n3402), .B(n3400), .S(n4900), .Z(n3401) );
  OAI21_X1 U4214 ( .B1(n3404), .B2(n4682), .A(n3401), .ZN(U3487) );
  MUX2_X1 U4215 ( .A(n3402), .B(n2619), .S(n4908), .Z(n3403) );
  OAI21_X1 U4216 ( .B1(n3404), .B2(n4629), .A(n3403), .ZN(U3528) );
  INV_X1 U4217 ( .A(n3405), .ZN(n3406) );
  AOI21_X1 U4218 ( .B1(n3431), .B2(n3407), .A(n3406), .ZN(n3521) );
  NAND2_X1 U4219 ( .A1(n3520), .A2(n3518), .ZN(n3854) );
  XNOR2_X1 U4220 ( .A(n3521), .B(n3854), .ZN(n3413) );
  OAI22_X1 U4221 ( .A1(n3408), .A2(n4541), .B1(n4565), .B2(n3499), .ZN(n3411)
         );
  NOR2_X1 U4222 ( .A1(n3409), .A2(n4528), .ZN(n3410) );
  OR2_X1 U4223 ( .A1(n3411), .A2(n3410), .ZN(n3412) );
  AOI21_X1 U4224 ( .B1(n3413), .B2(n4531), .A(n3412), .ZN(n3505) );
  NAND2_X1 U4225 ( .A1(n3442), .A2(n3414), .ZN(n3415) );
  NAND2_X1 U4226 ( .A1(n3528), .A2(n3415), .ZN(n3512) );
  INV_X1 U4227 ( .A(n3512), .ZN(n3419) );
  INV_X1 U4228 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3417) );
  INV_X1 U4229 ( .A(n3501), .ZN(n3416) );
  OAI22_X1 U4230 ( .A1(n4557), .A2(n3417), .B1(n3416), .B2(n4519), .ZN(n3418)
         );
  AOI21_X1 U4231 ( .B1(n3419), .B2(n4817), .A(n3418), .ZN(n3422) );
  XNOR2_X1 U4232 ( .A(n3420), .B(n3854), .ZN(n3504) );
  NAND2_X1 U4233 ( .A1(n3504), .A2(n4331), .ZN(n3421) );
  OAI211_X1 U4234 ( .C1(n3505), .C2(n4813), .A(n3422), .B(n3421), .ZN(U3278)
         );
  XOR2_X1 U4235 ( .A(n3425), .B(n3424), .Z(n3426) );
  XNOR2_X1 U4236 ( .A(n3423), .B(n3426), .ZN(n3430) );
  NOR2_X1 U4237 ( .A1(STATE_REG_SCAN_IN), .A2(n2636), .ZN(n4730) );
  OAI22_X1 U4238 ( .A1(n3539), .A2(n3780), .B1(n3781), .B2(n3437), .ZN(n3427)
         );
  AOI211_X1 U4239 ( .C1(n3435), .C2(n3784), .A(n4730), .B(n3427), .ZN(n3429)
         );
  NAND2_X1 U4240 ( .A1(n3787), .A2(n3445), .ZN(n3428) );
  OAI211_X1 U4241 ( .C1(n3430), .C2(n3790), .A(n3429), .B(n3428), .ZN(U3233)
         );
  XOR2_X1 U4242 ( .A(n3823), .B(n3431), .Z(n3440) );
  NAND2_X1 U4243 ( .A1(n3433), .A2(n3823), .ZN(n3434) );
  NAND2_X1 U4244 ( .A1(n3432), .A2(n3434), .ZN(n4898) );
  AOI22_X1 U4245 ( .A1(n4235), .A2(n4525), .B1(n3435), .B2(n4576), .ZN(n3436)
         );
  OAI21_X1 U4246 ( .B1(n3437), .B2(n4528), .A(n3436), .ZN(n3438) );
  AOI21_X1 U4247 ( .B1(n4898), .B2(n3626), .A(n3438), .ZN(n3439) );
  OAI21_X1 U4248 ( .B1(n4547), .B2(n3440), .A(n3439), .ZN(n4896) );
  INV_X1 U4249 ( .A(n4896), .ZN(n3450) );
  INV_X1 U4250 ( .A(n3441), .ZN(n3444) );
  OAI21_X1 U4251 ( .B1(n3444), .B2(n3443), .A(n3442), .ZN(n4895) );
  NOR2_X1 U4252 ( .A1(n4895), .A2(n4555), .ZN(n3448) );
  INV_X1 U4253 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3451) );
  INV_X1 U4254 ( .A(n3445), .ZN(n3446) );
  OAI22_X1 U4255 ( .A1(n3190), .A2(n3451), .B1(n3446), .B2(n4519), .ZN(n3447)
         );
  AOI211_X1 U4256 ( .C1(n4898), .C2(n4828), .A(n3448), .B(n3447), .ZN(n3449)
         );
  OAI21_X1 U4257 ( .B1(n3450), .B2(n4813), .A(n3449), .ZN(U3279) );
  NAND2_X1 U4258 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4855), .ZN(n3458) );
  INV_X1 U4259 ( .A(n4855), .ZN(n4737) );
  AOI22_X1 U4260 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4855), .B1(n4737), .B2(
        n3451), .ZN(n4734) );
  INV_X1 U4261 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3455) );
  AOI22_X1 U4262 ( .A1(n3467), .A2(REG2_REG_9__SCAN_IN), .B1(n3455), .B2(n4860), .ZN(n4716) );
  INV_X1 U4263 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3453) );
  OAI22_X1 U4264 ( .A1(n3454), .A2(n3453), .B1(n3452), .B2(n4692), .ZN(n4715)
         );
  NAND2_X1 U4265 ( .A1(n4716), .A2(n4715), .ZN(n4714) );
  OAI21_X1 U4266 ( .B1(n3455), .B2(n4860), .A(n4714), .ZN(n3456) );
  NAND2_X1 U4267 ( .A1(n4857), .A2(n3456), .ZN(n3457) );
  XNOR2_X1 U4268 ( .A(n3468), .B(n3456), .ZN(n4725) );
  NAND2_X1 U4269 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4725), .ZN(n4724) );
  NAND2_X1 U4270 ( .A1(n3459), .A2(n3460), .ZN(n3461) );
  NAND2_X1 U4271 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4745), .ZN(n4744) );
  INV_X1 U4272 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4108) );
  NOR2_X1 U4273 ( .A1(n3480), .A2(n4108), .ZN(n4293) );
  AOI21_X1 U4274 ( .B1(n4108), .B2(n3480), .A(n4293), .ZN(n3463) );
  AOI21_X1 U4275 ( .B1(n3463), .B2(n4294), .A(n4751), .ZN(n3462) );
  OAI21_X1 U4276 ( .B1(n4294), .B2(n3463), .A(n3462), .ZN(n3479) );
  AND2_X1 U4277 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n3541) );
  OAI21_X1 U4278 ( .B1(n3465), .B2(n4692), .A(n3464), .ZN(n3466) );
  INV_X1 U4279 ( .A(n3466), .ZN(n4711) );
  AOI22_X1 U4280 ( .A1(n3467), .A2(n2599), .B1(REG1_REG_9__SCAN_IN), .B2(n4860), .ZN(n4710) );
  NOR2_X1 U4281 ( .A1(n3469), .A2(n3468), .ZN(n3470) );
  AOI22_X1 U4282 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4737), .B1(n4855), .B2(
        n2639), .ZN(n4729) );
  NOR2_X1 U4283 ( .A1(n3471), .A2(n4854), .ZN(n3472) );
  XNOR2_X1 U4284 ( .A(n3471), .B(n4854), .ZN(n4739) );
  NAND2_X1 U4285 ( .A1(n4292), .A2(REG1_REG_13__SCAN_IN), .ZN(n4282) );
  NAND2_X1 U4286 ( .A1(n3480), .A2(n3577), .ZN(n3473) );
  NAND2_X1 U4287 ( .A1(n4282), .A2(n3473), .ZN(n3475) );
  INV_X1 U4288 ( .A(n4283), .ZN(n3474) );
  AOI211_X1 U4289 ( .C1(n3476), .C2(n3475), .A(n3474), .B(n4797), .ZN(n3477)
         );
  AOI211_X1 U4290 ( .C1(n4775), .C2(ADDR_REG_13__SCAN_IN), .A(n3541), .B(n3477), .ZN(n3478) );
  OAI211_X1 U4291 ( .C1(n4812), .C2(n3480), .A(n3479), .B(n3478), .ZN(U3253)
         );
  AOI22_X1 U4292 ( .A1(n3725), .A2(n3481), .B1(n3703), .B2(n3497), .ZN(n3482)
         );
  NAND2_X1 U4293 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4721) );
  OAI211_X1 U4294 ( .C1(n3769), .C2(n3483), .A(n3482), .B(n4721), .ZN(n3489)
         );
  INV_X1 U4295 ( .A(n3485), .ZN(n3486) );
  AOI211_X1 U4296 ( .C1(n3487), .C2(n3484), .A(n3790), .B(n3486), .ZN(n3488)
         );
  AOI211_X1 U4297 ( .C1(n3490), .C2(n3787), .A(n3489), .B(n3488), .ZN(n3491)
         );
  INV_X1 U4298 ( .A(n3491), .ZN(U3214) );
  INV_X1 U4299 ( .A(n3492), .ZN(n3494) );
  NOR2_X1 U4300 ( .A1(n3494), .A2(n3493), .ZN(n3495) );
  XNOR2_X1 U4301 ( .A(n3496), .B(n3495), .ZN(n3503) );
  AOI22_X1 U4302 ( .A1(n3725), .A2(n3497), .B1(n3703), .B2(n3583), .ZN(n3498)
         );
  NAND2_X1 U4303 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4741) );
  OAI211_X1 U4304 ( .C1(n3769), .C2(n3499), .A(n3498), .B(n4741), .ZN(n3500)
         );
  AOI21_X1 U4305 ( .B1(n3501), .B2(n3787), .A(n3500), .ZN(n3502) );
  OAI21_X1 U4306 ( .B1(n3503), .B2(n3790), .A(n3502), .ZN(U3221) );
  NAND2_X1 U4307 ( .A1(n3504), .A2(n4891), .ZN(n3506) );
  NAND2_X1 U4308 ( .A1(n3506), .A2(n3505), .ZN(n3509) );
  MUX2_X1 U4309 ( .A(n3509), .B(REG1_REG_12__SCAN_IN), .S(n4908), .Z(n3507) );
  INV_X1 U4310 ( .A(n3507), .ZN(n3508) );
  OAI21_X1 U4311 ( .B1(n4629), .B2(n3512), .A(n3508), .ZN(U3530) );
  MUX2_X1 U4312 ( .A(n3509), .B(REG0_REG_12__SCAN_IN), .S(n4900), .Z(n3510) );
  INV_X1 U4313 ( .A(n3510), .ZN(n3511) );
  OAI21_X1 U4314 ( .B1(n3512), .B2(n4682), .A(n3511), .ZN(U3491) );
  INV_X1 U4315 ( .A(n3513), .ZN(n3515) );
  OR2_X1 U4316 ( .A1(n3515), .A2(n3514), .ZN(n3850) );
  XOR2_X1 U4317 ( .A(n3850), .B(n3517), .Z(n3527) );
  INV_X1 U4318 ( .A(n3518), .ZN(n3519) );
  AOI21_X1 U4319 ( .B1(n3521), .B2(n3520), .A(n3519), .ZN(n3522) );
  XOR2_X1 U4320 ( .A(n3850), .B(n3522), .Z(n3525) );
  AOI22_X1 U4321 ( .A1(n3942), .A2(n4525), .B1(n4576), .B2(n3542), .ZN(n3523)
         );
  OAI21_X1 U4322 ( .B1(n3539), .B2(n4528), .A(n3523), .ZN(n3524) );
  AOI21_X1 U4323 ( .B1(n3525), .B2(n4531), .A(n3524), .ZN(n3526) );
  OAI21_X1 U4324 ( .B1(n3527), .B2(n4479), .A(n3526), .ZN(n3572) );
  INV_X1 U4325 ( .A(n3572), .ZN(n3534) );
  INV_X1 U4326 ( .A(n3527), .ZN(n3573) );
  INV_X1 U4327 ( .A(n3553), .ZN(n3530) );
  NAND2_X1 U4328 ( .A1(n3528), .A2(n3542), .ZN(n3529) );
  NAND2_X1 U4329 ( .A1(n3530), .A2(n3529), .ZN(n3579) );
  AOI22_X1 U4330 ( .A1(n4813), .A2(REG2_REG_13__SCAN_IN), .B1(n3543), .B2(
        n4826), .ZN(n3531) );
  OAI21_X1 U4331 ( .B1(n3579), .B2(n4555), .A(n3531), .ZN(n3532) );
  AOI21_X1 U4332 ( .B1(n3573), .B2(n4828), .A(n3532), .ZN(n3533) );
  OAI21_X1 U4333 ( .B1(n3534), .B2(n4813), .A(n3533), .ZN(U3277) );
  XOR2_X1 U4334 ( .A(n3536), .B(n3535), .Z(n3537) );
  XNOR2_X1 U4335 ( .A(n3538), .B(n3537), .ZN(n3546) );
  OAI22_X1 U4336 ( .A1(n3539), .A2(n3781), .B1(n3780), .B2(n3782), .ZN(n3540)
         );
  AOI211_X1 U4337 ( .C1(n3542), .C2(n3784), .A(n3541), .B(n3540), .ZN(n3545)
         );
  NAND2_X1 U4338 ( .A1(n3787), .A2(n3543), .ZN(n3544) );
  OAI211_X1 U4339 ( .C1(n3546), .C2(n3790), .A(n3545), .B(n3544), .ZN(U3231)
         );
  OAI21_X1 U4340 ( .B1(n3548), .B2(n3549), .A(n3547), .ZN(n3607) );
  INV_X1 U4341 ( .A(n3607), .ZN(n3558) );
  XNOR2_X1 U4342 ( .A(n3801), .B(n3549), .ZN(n3552) );
  OAI22_X1 U4343 ( .A1(n3603), .A2(n4541), .B1(n3585), .B2(n4565), .ZN(n3550)
         );
  AOI21_X1 U4344 ( .B1(n4545), .B2(n3583), .A(n3550), .ZN(n3551) );
  OAI21_X1 U4345 ( .B1(n3552), .B2(n4547), .A(n3551), .ZN(n3606) );
  OR2_X1 U4346 ( .A1(n3553), .A2(n3585), .ZN(n3554) );
  NAND2_X1 U4347 ( .A1(n3567), .A2(n3554), .ZN(n3612) );
  AOI22_X1 U4348 ( .A1(n4813), .A2(REG2_REG_14__SCAN_IN), .B1(n3587), .B2(
        n4826), .ZN(n3555) );
  OAI21_X1 U4349 ( .B1(n3612), .B2(n4555), .A(n3555), .ZN(n3556) );
  AOI21_X1 U4350 ( .B1(n3606), .B2(n4557), .A(n3556), .ZN(n3557) );
  OAI21_X1 U4351 ( .B1(n3558), .B2(n4559), .A(n3557), .ZN(U3276) );
  INV_X1 U4352 ( .A(n3559), .ZN(n3830) );
  XNOR2_X1 U4353 ( .A(n3560), .B(n3830), .ZN(n4639) );
  INV_X1 U4354 ( .A(n3561), .ZN(n3563) );
  OAI211_X1 U4355 ( .C1(n3563), .C2(n3830), .A(n4531), .B(n3562), .ZN(n3565)
         );
  AOI22_X1 U4356 ( .A1(n4544), .A2(n4525), .B1(n4576), .B2(n3785), .ZN(n3564)
         );
  OAI211_X1 U4357 ( .C1(n3782), .C2(n4528), .A(n3565), .B(n3564), .ZN(n4634)
         );
  XNOR2_X1 U4358 ( .A(n3567), .B(n3566), .ZN(n4635) );
  INV_X1 U4359 ( .A(n4635), .ZN(n3569) );
  AOI22_X1 U4360 ( .A1(n4813), .A2(REG2_REG_15__SCAN_IN), .B1(n3786), .B2(
        n4826), .ZN(n3568) );
  OAI21_X1 U4361 ( .B1(n3569), .B2(n4555), .A(n3568), .ZN(n3570) );
  AOI21_X1 U4362 ( .B1(n4634), .B2(n4557), .A(n3570), .ZN(n3571) );
  OAI21_X1 U4363 ( .B1(n4639), .B2(n4559), .A(n3571), .ZN(U3275) );
  INV_X1 U4364 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3574) );
  AOI21_X1 U4365 ( .B1(n4899), .B2(n3573), .A(n3572), .ZN(n3576) );
  MUX2_X1 U4366 ( .A(n3574), .B(n3576), .S(n4902), .Z(n3575) );
  OAI21_X1 U4367 ( .B1(n3579), .B2(n4682), .A(n3575), .ZN(U3493) );
  MUX2_X1 U4368 ( .A(n3577), .B(n3576), .S(n4910), .Z(n3578) );
  OAI21_X1 U4369 ( .B1(n4629), .B2(n3579), .A(n3578), .ZN(U3531) );
  NOR2_X1 U4370 ( .A1(n2394), .A2(n3581), .ZN(n3582) );
  XNOR2_X1 U4371 ( .A(n3580), .B(n3582), .ZN(n3589) );
  AOI22_X1 U4372 ( .A1(n3703), .A2(n3941), .B1(n3725), .B2(n3583), .ZN(n3584)
         );
  NAND2_X1 U4373 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4759) );
  OAI211_X1 U4374 ( .C1(n3769), .C2(n3585), .A(n3584), .B(n4759), .ZN(n3586)
         );
  AOI21_X1 U4375 ( .B1(n3587), .B2(n3787), .A(n3586), .ZN(n3588) );
  OAI21_X1 U4376 ( .B1(n3589), .B2(n3790), .A(n3588), .ZN(U3212) );
  OAI21_X1 U4377 ( .B1(n3592), .B2(n3591), .A(n3590), .ZN(n4633) );
  AOI21_X1 U4378 ( .B1(n3594), .B2(n3593), .A(n4550), .ZN(n4631) );
  INV_X1 U4379 ( .A(REG2_REG_16__SCAN_IN), .ZN(n3596) );
  INV_X1 U4380 ( .A(n3707), .ZN(n3595) );
  OAI22_X1 U4381 ( .A1(n3190), .A2(n3596), .B1(n3595), .B2(n4519), .ZN(n3597)
         );
  AOI21_X1 U4382 ( .B1(n4631), .B2(n4817), .A(n3597), .ZN(n3605) );
  OAI211_X1 U4383 ( .C1(n3599), .C2(n3842), .A(n3598), .B(n4531), .ZN(n3602)
         );
  OAI22_X1 U4384 ( .A1(n4529), .A2(n4541), .B1(n3705), .B2(n4565), .ZN(n3600)
         );
  INV_X1 U4385 ( .A(n3600), .ZN(n3601) );
  OAI211_X1 U4386 ( .C1(n3603), .C2(n4528), .A(n3602), .B(n3601), .ZN(n4630)
         );
  NAND2_X1 U4387 ( .A1(n4630), .A2(n4557), .ZN(n3604) );
  OAI211_X1 U4388 ( .C1(n4633), .C2(n4559), .A(n3605), .B(n3604), .ZN(U3274)
         );
  INV_X1 U4389 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3608) );
  AOI21_X1 U4390 ( .B1(n3607), .B2(n4891), .A(n3606), .ZN(n3610) );
  MUX2_X1 U4391 ( .A(n3608), .B(n3610), .S(n4902), .Z(n3609) );
  OAI21_X1 U4392 ( .B1(n3612), .B2(n4682), .A(n3609), .ZN(U3495) );
  MUX2_X1 U4393 ( .A(n4750), .B(n3610), .S(n4910), .Z(n3611) );
  OAI21_X1 U4394 ( .B1(n4629), .B2(n3612), .A(n3611), .ZN(U3532) );
  INV_X1 U4395 ( .A(n3613), .ZN(n3616) );
  OAI211_X1 U4396 ( .C1(n3616), .C2(n3615), .A(n4636), .B(n3614), .ZN(n4873)
         );
  NOR2_X1 U4397 ( .A1(n4873), .A2(n4691), .ZN(n3629) );
  XOR2_X1 U4398 ( .A(n3828), .B(n3618), .Z(n3628) );
  NAND2_X1 U4399 ( .A1(n3620), .A2(n3828), .ZN(n3621) );
  AND2_X1 U4400 ( .A1(n3619), .A2(n3621), .ZN(n4876) );
  AOI22_X1 U4401 ( .A1(n4238), .A2(n4545), .B1(n3622), .B2(n4576), .ZN(n3623)
         );
  OAI21_X1 U4402 ( .B1(n3624), .B2(n4541), .A(n3623), .ZN(n3625) );
  AOI21_X1 U4403 ( .B1(n4876), .B2(n3626), .A(n3625), .ZN(n3627) );
  OAI21_X1 U4404 ( .B1(n4547), .B2(n3628), .A(n3627), .ZN(n4874) );
  AOI211_X1 U4405 ( .C1(n4826), .C2(n3630), .A(n3629), .B(n4874), .ZN(n3632)
         );
  AOI22_X1 U4406 ( .A1(n4876), .A2(n4828), .B1(REG2_REG_4__SCAN_IN), .B2(n4813), .ZN(n3631) );
  OAI21_X1 U4407 ( .B1(n3632), .B2(n4813), .A(n3631), .ZN(U3286) );
  INV_X1 U4408 ( .A(n3633), .ZN(n3638) );
  AOI22_X1 U4409 ( .A1(n4813), .A2(REG2_REG_28__SCAN_IN), .B1(n3634), .B2(
        n4826), .ZN(n3635) );
  OAI21_X1 U4410 ( .B1(n3636), .B2(n4555), .A(n3635), .ZN(n3637) );
  AOI21_X1 U4411 ( .B1(n3638), .B2(n4557), .A(n3637), .ZN(n3639) );
  OAI21_X1 U4412 ( .B1(n3640), .B2(n4559), .A(n3639), .ZN(U3262) );
  OR2_X1 U4413 ( .A1(n3642), .A2(n3641), .ZN(n3643) );
  AND2_X1 U4414 ( .A1(n3644), .A2(n3643), .ZN(n4258) );
  AOI22_X1 U4415 ( .A1(n4258), .A2(n3757), .B1(n3645), .B2(n3784), .ZN(n3647)
         );
  NAND2_X1 U4416 ( .A1(n3673), .A2(REG3_REG_0__SCAN_IN), .ZN(n3646) );
  OAI211_X1 U4417 ( .C1(n2905), .C2(n3780), .A(n3647), .B(n3646), .ZN(U3229)
         );
  OAI21_X1 U4418 ( .B1(n3742), .B2(n3650), .A(n3649), .ZN(n3651) );
  NAND3_X1 U4419 ( .A1(n2338), .A2(n3757), .A3(n3651), .ZN(n3656) );
  NAND2_X1 U4420 ( .A1(n3703), .A2(n4420), .ZN(n3653) );
  AOI22_X1 U4421 ( .A1(n3784), .A2(n4419), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3652) );
  OAI211_X1 U4422 ( .C1(n4423), .C2(n3781), .A(n3653), .B(n3652), .ZN(n3654)
         );
  INV_X1 U4423 ( .A(n3654), .ZN(n3655) );
  OAI211_X1 U4424 ( .C1(n3762), .C2(n4427), .A(n3656), .B(n3655), .ZN(U3213)
         );
  INV_X1 U4425 ( .A(n3756), .ZN(n3659) );
  INV_X1 U4426 ( .A(n3753), .ZN(n3658) );
  OAI21_X1 U4427 ( .B1(n3756), .B2(n3753), .A(n3754), .ZN(n3657) );
  OAI21_X1 U4428 ( .B1(n3659), .B2(n3658), .A(n3657), .ZN(n3663) );
  NOR2_X1 U4429 ( .A1(n3661), .A2(n3660), .ZN(n3662) );
  XNOR2_X1 U4430 ( .A(n3663), .B(n3662), .ZN(n3668) );
  INV_X1 U4431 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4038) );
  NOR2_X1 U4432 ( .A1(n4038), .A2(STATE_REG_SCAN_IN), .ZN(n4305) );
  OAI22_X1 U4433 ( .A1(n4542), .A2(n3781), .B1(n3780), .B2(n4498), .ZN(n3664)
         );
  AOI211_X1 U4434 ( .C1(n3665), .C2(n3784), .A(n4305), .B(n3664), .ZN(n3667)
         );
  NAND2_X1 U4435 ( .A1(n3787), .A2(n4508), .ZN(n3666) );
  OAI211_X1 U4436 ( .C1(n3668), .C2(n3790), .A(n3667), .B(n3666), .ZN(U3216)
         );
  OAI211_X1 U4437 ( .C1(n3669), .C2(n3670), .A(n3671), .B(n3757), .ZN(n3676)
         );
  AOI22_X1 U4438 ( .A1(n3725), .A2(n2944), .B1(n2904), .B2(n3784), .ZN(n3675)
         );
  AOI22_X1 U4439 ( .A1(REG3_REG_1__SCAN_IN), .A2(n3673), .B1(n3703), .B2(n3672), .ZN(n3674) );
  NAND3_X1 U4440 ( .A1(n3676), .A2(n3675), .A3(n3674), .ZN(U3219) );
  INV_X1 U4441 ( .A(n3678), .ZN(n3680) );
  NAND2_X1 U4442 ( .A1(n3680), .A2(n3679), .ZN(n3684) );
  INV_X1 U4443 ( .A(n3735), .ZN(n3682) );
  OAI211_X1 U4444 ( .C1(n3681), .C2(n3682), .A(n3733), .B(n3684), .ZN(n3683)
         );
  OAI211_X1 U4445 ( .C1(n3677), .C2(n3684), .A(n3757), .B(n3683), .ZN(n3688)
         );
  OAI22_X1 U4446 ( .A1(n3769), .A2(n4459), .B1(STATE_REG_SCAN_IN), .B2(n4039), 
        .ZN(n3686) );
  OAI22_X1 U4447 ( .A1(n4498), .A2(n3781), .B1(n3780), .B2(n4423), .ZN(n3685)
         );
  AOI211_X1 U4448 ( .C1(n4462), .C2(n3787), .A(n3686), .B(n3685), .ZN(n3687)
         );
  NAND2_X1 U4449 ( .A1(n3688), .A2(n3687), .ZN(U3220) );
  INV_X1 U4450 ( .A(n3689), .ZN(n3691) );
  NAND2_X1 U4451 ( .A1(n3691), .A2(n3690), .ZN(n3692) );
  XNOR2_X1 U4452 ( .A(n3693), .B(n3692), .ZN(n3694) );
  NAND2_X1 U4453 ( .A1(n3694), .A2(n3757), .ZN(n3699) );
  NAND2_X1 U4454 ( .A1(n3725), .A2(n4420), .ZN(n3696) );
  AOI22_X1 U4455 ( .A1(n3784), .A2(n4377), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n3695) );
  OAI211_X1 U4456 ( .C1(n4345), .C2(n3780), .A(n3696), .B(n3695), .ZN(n3697)
         );
  INV_X1 U4457 ( .A(n3697), .ZN(n3698) );
  OAI211_X1 U4458 ( .C1(n3762), .C2(n4385), .A(n3699), .B(n3698), .ZN(U3222)
         );
  AOI21_X1 U4459 ( .B1(n3700), .B2(n3774), .A(n3776), .ZN(n3702) );
  XNOR2_X1 U4460 ( .A(n3702), .B(n3701), .ZN(n3709) );
  AOI22_X1 U4461 ( .A1(n3703), .A2(n3940), .B1(n3725), .B2(n3941), .ZN(n3704)
         );
  NAND2_X1 U4462 ( .A1(REG3_REG_16__SCAN_IN), .A2(U3149), .ZN(n4773) );
  OAI211_X1 U4463 ( .C1(n3769), .C2(n3705), .A(n3704), .B(n4773), .ZN(n3706)
         );
  AOI21_X1 U4464 ( .B1(n3707), .B2(n3787), .A(n3706), .ZN(n3708) );
  OAI21_X1 U4465 ( .B1(n3709), .B2(n3790), .A(n3708), .ZN(U3223) );
  NAND2_X1 U4466 ( .A1(n2192), .A2(n3711), .ZN(n3712) );
  XNOR2_X1 U4467 ( .A(n3710), .B(n3712), .ZN(n3717) );
  INV_X1 U4468 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4095) );
  NOR2_X1 U4469 ( .A1(STATE_REG_SCAN_IN), .A2(n4095), .ZN(n4785) );
  OAI22_X1 U4470 ( .A1(n3779), .A2(n3781), .B1(n3780), .B2(n4542), .ZN(n3713)
         );
  AOI211_X1 U4471 ( .C1(n3714), .C2(n3784), .A(n4785), .B(n3713), .ZN(n3716)
         );
  NAND2_X1 U4472 ( .A1(n3787), .A2(n4553), .ZN(n3715) );
  OAI211_X1 U4473 ( .C1(n3717), .C2(n3790), .A(n3716), .B(n3715), .ZN(U3225)
         );
  INV_X1 U4474 ( .A(n3718), .ZN(n3719) );
  NOR2_X1 U4475 ( .A1(n3720), .A2(n3719), .ZN(n3722) );
  XNOR2_X1 U4476 ( .A(n3722), .B(n3721), .ZN(n3723) );
  NAND2_X1 U4477 ( .A1(n3723), .A2(n3757), .ZN(n3731) );
  NAND2_X1 U4478 ( .A1(n3725), .A2(n3724), .ZN(n3728) );
  AOI22_X1 U4479 ( .A1(n3784), .A2(n3726), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3727) );
  OAI211_X1 U4480 ( .C1(n4359), .C2(n3780), .A(n3728), .B(n3727), .ZN(n3729)
         );
  INV_X1 U4481 ( .A(n3729), .ZN(n3730) );
  OAI211_X1 U4482 ( .C1(n3762), .C2(n4405), .A(n3731), .B(n3730), .ZN(U3226)
         );
  INV_X1 U4483 ( .A(n3732), .ZN(n3736) );
  AOI21_X1 U4484 ( .B1(n3733), .B2(n3735), .A(n3681), .ZN(n3734) );
  AOI21_X1 U4485 ( .B1(n3736), .B2(n3735), .A(n3734), .ZN(n3741) );
  INV_X1 U4486 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3737) );
  OAI22_X1 U4487 ( .A1(n3769), .A2(n4481), .B1(STATE_REG_SCAN_IN), .B2(n3737), 
        .ZN(n3739) );
  OAI22_X1 U4488 ( .A1(n4475), .A2(n3781), .B1(n3780), .B2(n3747), .ZN(n3738)
         );
  AOI211_X1 U4489 ( .C1(n4484), .C2(n3787), .A(n3739), .B(n3738), .ZN(n3740)
         );
  OAI21_X1 U4490 ( .B1(n3741), .B2(n3790), .A(n3740), .ZN(U3230) );
  AOI21_X1 U4491 ( .B1(n3744), .B2(n3743), .A(n3742), .ZN(n3752) );
  OAI22_X1 U4492 ( .A1(n3769), .A2(n3746), .B1(STATE_REG_SCAN_IN), .B2(n3745), 
        .ZN(n3749) );
  OAI22_X1 U4493 ( .A1(n4440), .A2(n3780), .B1(n3781), .B2(n3747), .ZN(n3748)
         );
  AOI211_X1 U4494 ( .C1(n3750), .C2(n3787), .A(n3749), .B(n3748), .ZN(n3751)
         );
  OAI21_X1 U4495 ( .B1(n3752), .B2(n3790), .A(n3751), .ZN(U3232) );
  XNOR2_X1 U4496 ( .A(n3754), .B(n3753), .ZN(n3755) );
  XNOR2_X1 U4497 ( .A(n3756), .B(n3755), .ZN(n3758) );
  NAND2_X1 U4498 ( .A1(n3758), .A2(n3757), .ZN(n3761) );
  AND2_X1 U4499 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4800) );
  OAI22_X1 U4500 ( .A1(n4475), .A2(n3780), .B1(n3781), .B2(n4529), .ZN(n3759)
         );
  AOI211_X1 U4501 ( .C1(n4524), .C2(n3784), .A(n4800), .B(n3759), .ZN(n3760)
         );
  OAI211_X1 U4502 ( .C1(n3762), .C2(n4520), .A(n3761), .B(n3760), .ZN(U3235)
         );
  INV_X1 U4503 ( .A(n3763), .ZN(n3765) );
  NAND2_X1 U4504 ( .A1(n3765), .A2(n3764), .ZN(n3766) );
  XNOR2_X1 U4505 ( .A(n3767), .B(n3766), .ZN(n3773) );
  OAI22_X1 U4506 ( .A1(n3769), .A2(n4365), .B1(STATE_REG_SCAN_IN), .B2(n3768), 
        .ZN(n3771) );
  OAI22_X1 U4507 ( .A1(n3865), .A2(n3780), .B1(n3781), .B2(n4359), .ZN(n3770)
         );
  AOI211_X1 U4508 ( .C1(n4367), .C2(n3787), .A(n3771), .B(n3770), .ZN(n3772)
         );
  OAI21_X1 U4509 ( .B1(n3773), .B2(n3790), .A(n3772), .ZN(U3237) );
  INV_X1 U4510 ( .A(n3774), .ZN(n3775) );
  NOR2_X1 U4511 ( .A1(n3776), .A2(n3775), .ZN(n3778) );
  XNOR2_X1 U4512 ( .A(n3778), .B(n3777), .ZN(n3791) );
  INV_X1 U4513 ( .A(REG3_REG_15__SCAN_IN), .ZN(n4020) );
  NOR2_X1 U4514 ( .A1(STATE_REG_SCAN_IN), .A2(n4020), .ZN(n4766) );
  OAI22_X1 U4515 ( .A1(n3782), .A2(n3781), .B1(n3780), .B2(n3779), .ZN(n3783)
         );
  AOI211_X1 U4516 ( .C1(n3785), .C2(n3784), .A(n4766), .B(n3783), .ZN(n3789)
         );
  NAND2_X1 U4517 ( .A1(n3787), .A2(n3786), .ZN(n3788) );
  OAI211_X1 U4518 ( .C1(n3791), .C2(n3790), .A(n3789), .B(n3788), .ZN(U3238)
         );
  AND2_X1 U4519 ( .A1(n3794), .A2(DATAI_29_), .ZN(n4333) );
  INV_X1 U4520 ( .A(n4333), .ZN(n4332) );
  AND2_X1 U4521 ( .A1(n3859), .A2(n4332), .ZN(n3792) );
  OR2_X1 U4522 ( .A1(n4312), .A2(n3792), .ZN(n3919) );
  INV_X1 U4523 ( .A(n3919), .ZN(n3797) );
  OR2_X1 U4524 ( .A1(n4313), .A2(n3799), .ZN(n3796) );
  AND2_X1 U4525 ( .A1(n3794), .A2(DATAI_30_), .ZN(n4577) );
  AOI222_X1 U4526 ( .A1(n2700), .A2(REG2_REG_31__SCAN_IN), .B1(n3793), .B2(
        REG1_REG_31__SCAN_IN), .C1(n2533), .C2(REG0_REG_31__SCAN_IN), .ZN(
        n4564) );
  NAND2_X1 U4527 ( .A1(n3794), .A2(DATAI_31_), .ZN(n4566) );
  INV_X1 U4528 ( .A(n4566), .ZN(n3795) );
  NOR2_X1 U4529 ( .A1(n4564), .A2(n3795), .ZN(n3925) );
  AOI21_X1 U4530 ( .B1(n4577), .B2(n4320), .A(n3925), .ZN(n3841) );
  OAI21_X1 U4531 ( .B1(n3859), .B2(n4332), .A(n3841), .ZN(n3798) );
  AOI21_X1 U4532 ( .B1(n3797), .B2(n3796), .A(n3798), .ZN(n3923) );
  NAND3_X1 U4533 ( .A1(n4340), .A2(n3797), .A3(n3838), .ZN(n3819) );
  NOR4_X1 U4534 ( .A1(n4313), .A2(n3799), .A3(n3915), .A4(n3798), .ZN(n3818)
         );
  INV_X1 U4535 ( .A(n3906), .ZN(n3805) );
  NAND2_X1 U4536 ( .A1(n3800), .A2(n3804), .ZN(n3904) );
  NOR3_X1 U4537 ( .A1(n3801), .A2(n3805), .A3(n3904), .ZN(n3803) );
  INV_X1 U4538 ( .A(n3802), .ZN(n3908) );
  OAI21_X1 U4539 ( .B1(n3803), .B2(n3908), .A(n3907), .ZN(n3813) );
  INV_X1 U4540 ( .A(n3804), .ZN(n3806) );
  AOI211_X1 U4541 ( .C1(n3808), .C2(n3807), .A(n3806), .B(n3805), .ZN(n3810)
         );
  OAI21_X1 U4542 ( .B1(n3810), .B2(n3809), .A(n3907), .ZN(n3812) );
  AND2_X1 U4543 ( .A1(n3812), .A2(n3811), .ZN(n3911) );
  NAND2_X1 U4544 ( .A1(n3813), .A2(n3911), .ZN(n3815) );
  AOI21_X1 U4545 ( .B1(n3914), .B2(n3815), .A(n3814), .ZN(n3816) );
  OAI21_X1 U4546 ( .B1(n3816), .B2(n3916), .A(n4354), .ZN(n3817) );
  AOI22_X1 U4547 ( .A1(n3923), .A2(n3819), .B1(n3818), .B2(n3817), .ZN(n3822)
         );
  INV_X1 U4548 ( .A(n4564), .ZN(n3938) );
  INV_X1 U4549 ( .A(n4577), .ZN(n4561) );
  NOR2_X1 U4550 ( .A1(n3938), .A2(n4561), .ZN(n3821) );
  NOR2_X1 U4551 ( .A1(n4320), .A2(n4577), .ZN(n3836) );
  NOR2_X1 U4552 ( .A1(n3836), .A2(n4564), .ZN(n3820) );
  OAI22_X1 U4553 ( .A1(n3822), .A2(n3821), .B1(n3820), .B2(n4566), .ZN(n3864)
         );
  INV_X1 U4554 ( .A(n4327), .ZN(n3835) );
  INV_X1 U4555 ( .A(n4515), .ZN(n4522) );
  NAND4_X1 U4556 ( .A1(n3825), .A2(n4522), .A3(n3824), .A4(n3823), .ZN(n3834)
         );
  INV_X1 U4557 ( .A(n2943), .ZN(n3826) );
  NAND4_X1 U4558 ( .A1(n3829), .A2(n3828), .A3(n3827), .A4(n3826), .ZN(n3833)
         );
  AND2_X1 U4559 ( .A1(n4491), .A2(n4490), .ZN(n4539) );
  NOR2_X1 U4560 ( .A1(n4412), .A2(n4414), .ZN(n4451) );
  NAND4_X1 U4561 ( .A1(n3831), .A2(n4539), .A3(n3830), .A4(n4451), .ZN(n3832)
         );
  NOR4_X1 U4562 ( .A1(n3835), .A2(n3834), .A3(n3833), .A4(n3832), .ZN(n3858)
         );
  INV_X1 U4563 ( .A(n3836), .ZN(n3837) );
  OAI21_X1 U4564 ( .B1(n3938), .B2(n4566), .A(n3837), .ZN(n3924) );
  NAND4_X1 U4565 ( .A1(n4340), .A2(n4358), .A3(n4375), .A4(n3841), .ZN(n3844)
         );
  NAND2_X1 U4566 ( .A1(n3842), .A2(n4434), .ZN(n3843) );
  NOR4_X1 U4567 ( .A1(n3924), .A2(n3844), .A3(n3843), .A4(n4827), .ZN(n3857)
         );
  NAND2_X1 U4568 ( .A1(n3845), .A2(n4392), .ZN(n4416) );
  NAND2_X1 U4569 ( .A1(n3846), .A2(n4374), .ZN(n4396) );
  INV_X1 U4570 ( .A(n3847), .ZN(n3849) );
  OR2_X1 U4571 ( .A1(n3849), .A2(n3848), .ZN(n4496) );
  NOR4_X1 U4572 ( .A1(n4416), .A2(n4396), .A3(n4496), .A4(n3850), .ZN(n3856)
         );
  NOR4_X1 U4573 ( .A1(n3854), .A2(n3853), .A3(n3852), .A4(n3851), .ZN(n3855)
         );
  AND4_X1 U4574 ( .A1(n3858), .A2(n3857), .A3(n3856), .A4(n3855), .ZN(n3861)
         );
  XNOR2_X1 U4575 ( .A(n3859), .B(n4333), .ZN(n4329) );
  XNOR2_X1 U4576 ( .A(n4498), .B(n4481), .ZN(n4470) );
  NAND4_X1 U4577 ( .A1(n3861), .A2(n4329), .A3(n4470), .A4(n3860), .ZN(n3863)
         );
  MUX2_X1 U4578 ( .A(n3864), .B(n3863), .S(n3862), .Z(n3931) );
  NOR2_X1 U4579 ( .A1(n3865), .A2(n4347), .ZN(n3922) );
  INV_X1 U4580 ( .A(n3866), .ZN(n3869) );
  OAI211_X1 U4581 ( .C1(n3869), .C2(n4689), .A(n3868), .B(n3867), .ZN(n3872)
         );
  NAND3_X1 U4582 ( .A1(n3872), .A2(n3871), .A3(n3870), .ZN(n3875) );
  NAND3_X1 U4583 ( .A1(n3875), .A2(n3874), .A3(n3873), .ZN(n3878) );
  NAND3_X1 U4584 ( .A1(n3878), .A2(n3877), .A3(n3876), .ZN(n3881) );
  NAND3_X1 U4585 ( .A1(n3881), .A2(n3880), .A3(n3879), .ZN(n3885) );
  INV_X1 U4586 ( .A(n3882), .ZN(n3883) );
  AOI21_X1 U4587 ( .B1(n3885), .B2(n3884), .A(n3883), .ZN(n3891) );
  NAND2_X1 U4588 ( .A1(n3887), .A2(n3886), .ZN(n3890) );
  OAI211_X1 U4589 ( .C1(n3891), .C2(n3890), .A(n3889), .B(n3888), .ZN(n3894)
         );
  NAND3_X1 U4590 ( .A1(n3894), .A2(n3893), .A3(n3892), .ZN(n3896) );
  NAND2_X1 U4591 ( .A1(n3896), .A2(n3895), .ZN(n3901) );
  INV_X1 U4592 ( .A(n3898), .ZN(n3899) );
  AOI211_X1 U4593 ( .C1(n3901), .C2(n3900), .A(n2228), .B(n3899), .ZN(n3905)
         );
  INV_X1 U4594 ( .A(n3902), .ZN(n3903) );
  NOR3_X1 U4595 ( .A1(n3905), .A2(n3904), .A3(n3903), .ZN(n3909) );
  OAI211_X1 U4596 ( .C1(n3909), .C2(n3908), .A(n3907), .B(n3906), .ZN(n3912)
         );
  INV_X1 U4597 ( .A(n4414), .ZN(n3910) );
  NAND3_X1 U4598 ( .A1(n3912), .A2(n3911), .A3(n3910), .ZN(n3913) );
  NAND2_X1 U4599 ( .A1(n3914), .A2(n3913), .ZN(n3917) );
  AOI211_X1 U4600 ( .C1(n3918), .C2(n3917), .A(n3916), .B(n3915), .ZN(n3921)
         );
  NOR4_X1 U4601 ( .A1(n3922), .A2(n3921), .A3(n3920), .A4(n3919), .ZN(n3928)
         );
  INV_X1 U4602 ( .A(n3923), .ZN(n3927) );
  INV_X1 U4603 ( .A(n3924), .ZN(n3926) );
  OAI22_X1 U4604 ( .A1(n3928), .A2(n3927), .B1(n3926), .B2(n3925), .ZN(n3930)
         );
  MUX2_X1 U4605 ( .A(n3931), .B(n3930), .S(n3929), .Z(n3932) );
  XNOR2_X1 U4606 ( .A(n3932), .B(n4307), .ZN(n3937) );
  NOR2_X1 U4607 ( .A1(n3933), .A2(n4251), .ZN(n3935) );
  OAI21_X1 U4608 ( .B1(n3936), .B2(n4688), .A(B_REG_SCAN_IN), .ZN(n3934) );
  OAI22_X1 U4609 ( .A1(n3937), .A2(n3936), .B1(n3935), .B2(n3934), .ZN(U3239)
         );
  MUX2_X1 U4610 ( .A(DATAO_REG_31__SCAN_IN), .B(n3938), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4611 ( .A(n4361), .B(DATAO_REG_27__SCAN_IN), .S(n4240), .Z(U3577)
         );
  MUX2_X1 U4612 ( .A(n4420), .B(DATAO_REG_24__SCAN_IN), .S(n4240), .Z(U3574)
         );
  MUX2_X1 U4613 ( .A(n4454), .B(DATAO_REG_22__SCAN_IN), .S(n4240), .Z(U3572)
         );
  MUX2_X1 U4614 ( .A(n4473), .B(DATAO_REG_21__SCAN_IN), .S(n4240), .Z(U3571)
         );
  MUX2_X1 U4615 ( .A(n4455), .B(DATAO_REG_20__SCAN_IN), .S(n4240), .Z(U3570)
         );
  MUX2_X1 U4616 ( .A(n4526), .B(DATAO_REG_19__SCAN_IN), .S(n4240), .Z(U3569)
         );
  MUX2_X1 U4617 ( .A(n3939), .B(DATAO_REG_18__SCAN_IN), .S(n4240), .Z(U3568)
         );
  MUX2_X1 U4618 ( .A(n3940), .B(DATAO_REG_17__SCAN_IN), .S(n4240), .Z(U3567)
         );
  MUX2_X1 U4619 ( .A(n4544), .B(DATAO_REG_16__SCAN_IN), .S(n4240), .Z(U3566)
         );
  MUX2_X1 U4620 ( .A(n3941), .B(DATAO_REG_15__SCAN_IN), .S(n4240), .Z(U3565)
         );
  MUX2_X1 U4621 ( .A(DATAO_REG_14__SCAN_IN), .B(n3942), .S(U4043), .Z(n4234)
         );
  INV_X1 U4622 ( .A(D_REG_13__SCAN_IN), .ZN(n4834) );
  AOI22_X1 U4623 ( .A1(n4834), .A2(keyinput88), .B1(keyinput45), .B2(n2593), 
        .ZN(n3943) );
  OAI221_X1 U4624 ( .B1(n4834), .B2(keyinput88), .C1(n2593), .C2(keyinput45), 
        .A(n3943), .ZN(n3953) );
  INV_X1 U4625 ( .A(D_REG_11__SCAN_IN), .ZN(n4835) );
  INV_X1 U4626 ( .A(keyinput33), .ZN(n3945) );
  AOI22_X1 U4627 ( .A1(n4835), .A2(keyinput41), .B1(DATAO_REG_28__SCAN_IN), 
        .B2(n3945), .ZN(n3944) );
  OAI221_X1 U4628 ( .B1(n4835), .B2(keyinput41), .C1(n3945), .C2(
        DATAO_REG_28__SCAN_IN), .A(n3944), .ZN(n3952) );
  INV_X1 U4629 ( .A(DATAI_19_), .ZN(n3947) );
  INV_X1 U4630 ( .A(D_REG_8__SCAN_IN), .ZN(n4838) );
  AOI22_X1 U4631 ( .A1(n3947), .A2(keyinput37), .B1(n4838), .B2(keyinput57), 
        .ZN(n3946) );
  OAI221_X1 U4632 ( .B1(n3947), .B2(keyinput37), .C1(n4838), .C2(keyinput57), 
        .A(n3946), .ZN(n3951) );
  INV_X1 U4633 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4599) );
  INV_X1 U4634 ( .A(REG2_REG_17__SCAN_IN), .ZN(n3949) );
  AOI22_X1 U4635 ( .A1(n4599), .A2(keyinput61), .B1(n3949), .B2(keyinput49), 
        .ZN(n3948) );
  OAI221_X1 U4636 ( .B1(n4599), .B2(keyinput61), .C1(n3949), .C2(keyinput49), 
        .A(n3948), .ZN(n3950) );
  NOR4_X1 U4637 ( .A1(n3953), .A2(n3952), .A3(n3951), .A4(n3950), .ZN(n3991)
         );
  INV_X1 U4638 ( .A(D_REG_9__SCAN_IN), .ZN(n4837) );
  AOI22_X1 U4639 ( .A1(n4837), .A2(keyinput9), .B1(keyinput25), .B2(n3955), 
        .ZN(n3954) );
  OAI221_X1 U4640 ( .B1(n4837), .B2(keyinput9), .C1(n3955), .C2(keyinput25), 
        .A(n3954), .ZN(n3965) );
  INV_X1 U4641 ( .A(keyinput17), .ZN(n3957) );
  AOI22_X1 U4642 ( .A1(n4750), .A2(keyinput29), .B1(DATAO_REG_6__SCAN_IN), 
        .B2(n3957), .ZN(n3956) );
  OAI221_X1 U4643 ( .B1(n4750), .B2(keyinput29), .C1(n3957), .C2(
        DATAO_REG_6__SCAN_IN), .A(n3956), .ZN(n3964) );
  XOR2_X1 U4644 ( .A(n3958), .B(keyinput13), .Z(n3962) );
  XNOR2_X1 U4645 ( .A(DATAI_4_), .B(keyinput5), .ZN(n3961) );
  XNOR2_X1 U4646 ( .A(IR_REG_17__SCAN_IN), .B(keyinput53), .ZN(n3960) );
  XNOR2_X1 U4647 ( .A(DATAI_3_), .B(keyinput1), .ZN(n3959) );
  NAND4_X1 U4648 ( .A1(n3962), .A2(n3961), .A3(n3960), .A4(n3959), .ZN(n3963)
         );
  NOR3_X1 U4649 ( .A1(n3965), .A2(n3964), .A3(n3963), .ZN(n3990) );
  INV_X1 U4650 ( .A(REG3_REG_12__SCAN_IN), .ZN(n3967) );
  INV_X1 U4651 ( .A(DATAI_23_), .ZN(n4844) );
  AOI22_X1 U4652 ( .A1(n3967), .A2(keyinput121), .B1(keyinput117), .B2(n4844), 
        .ZN(n3966) );
  OAI221_X1 U4653 ( .B1(n3967), .B2(keyinput121), .C1(n4844), .C2(keyinput117), 
        .A(n3966), .ZN(n3976) );
  INV_X1 U4654 ( .A(keyinput109), .ZN(n3969) );
  AOI22_X1 U4655 ( .A1(n2231), .A2(keyinput21), .B1(DATAO_REG_2__SCAN_IN), 
        .B2(n3969), .ZN(n3968) );
  OAI221_X1 U4656 ( .B1(n2231), .B2(keyinput21), .C1(n3969), .C2(
        DATAO_REG_2__SCAN_IN), .A(n3968), .ZN(n3975) );
  XOR2_X1 U4657 ( .A(n2419), .B(keyinput125), .Z(n3973) );
  XNOR2_X1 U4658 ( .A(REG3_REG_28__SCAN_IN), .B(keyinput105), .ZN(n3972) );
  XNOR2_X1 U4659 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput97), .ZN(n3971) );
  XNOR2_X1 U4660 ( .A(IR_REG_23__SCAN_IN), .B(keyinput101), .ZN(n3970) );
  NAND4_X1 U4661 ( .A1(n3973), .A2(n3972), .A3(n3971), .A4(n3970), .ZN(n3974)
         );
  NOR3_X1 U4662 ( .A1(n3976), .A2(n3975), .A3(n3974), .ZN(n3989) );
  INV_X1 U4663 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4754) );
  INV_X1 U4664 ( .A(DATAI_6_), .ZN(n3978) );
  AOI22_X1 U4665 ( .A1(n4754), .A2(keyinput113), .B1(keyinput77), .B2(n3978), 
        .ZN(n3977) );
  OAI221_X1 U4666 ( .B1(n4754), .B2(keyinput113), .C1(n3978), .C2(keyinput77), 
        .A(n3977), .ZN(n3987) );
  INV_X1 U4667 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4705) );
  INV_X1 U4668 ( .A(keyinput73), .ZN(n3980) );
  AOI22_X1 U4669 ( .A1(n4705), .A2(keyinput65), .B1(DATAO_REG_23__SCAN_IN), 
        .B2(n3980), .ZN(n3979) );
  OAI221_X1 U4670 ( .B1(n4705), .B2(keyinput65), .C1(n3980), .C2(
        DATAO_REG_23__SCAN_IN), .A(n3979), .ZN(n3986) );
  INV_X1 U4671 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4865) );
  INV_X1 U4672 ( .A(REG2_REG_20__SCAN_IN), .ZN(n3982) );
  AOI22_X1 U4673 ( .A1(n4865), .A2(keyinput69), .B1(n3982), .B2(keyinput89), 
        .ZN(n3981) );
  OAI221_X1 U4674 ( .B1(n4865), .B2(keyinput69), .C1(n3982), .C2(keyinput89), 
        .A(n3981), .ZN(n3985) );
  INV_X1 U4675 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4643) );
  INV_X1 U4676 ( .A(DATAI_28_), .ZN(n4700) );
  AOI22_X1 U4677 ( .A1(n4643), .A2(keyinput93), .B1(n4700), .B2(keyinput85), 
        .ZN(n3983) );
  OAI221_X1 U4678 ( .B1(n4643), .B2(keyinput93), .C1(n4700), .C2(keyinput85), 
        .A(n3983), .ZN(n3984) );
  NOR4_X1 U4679 ( .A1(n3987), .A2(n3986), .A3(n3985), .A4(n3984), .ZN(n3988)
         );
  NAND4_X1 U4680 ( .A1(n3991), .A2(n3990), .A3(n3989), .A4(n3988), .ZN(n4232)
         );
  INV_X1 U4681 ( .A(keyinput62), .ZN(n3994) );
  INV_X1 U4682 ( .A(keyinput50), .ZN(n3993) );
  AOI22_X1 U4683 ( .A1(n3994), .A2(DATAO_REG_11__SCAN_IN), .B1(
        DATAO_REG_13__SCAN_IN), .B2(n3993), .ZN(n3992) );
  OAI221_X1 U4684 ( .B1(n3994), .B2(DATAO_REG_11__SCAN_IN), .C1(n3993), .C2(
        DATAO_REG_13__SCAN_IN), .A(n3992), .ZN(n4004) );
  INV_X1 U4685 ( .A(keyinput22), .ZN(n4210) );
  INV_X1 U4686 ( .A(keyinput55), .ZN(n3996) );
  AOI22_X1 U4687 ( .A1(n4210), .A2(DATAO_REG_10__SCAN_IN), .B1(
        DATAO_REG_8__SCAN_IN), .B2(n3996), .ZN(n3995) );
  OAI221_X1 U4688 ( .B1(n4210), .B2(DATAO_REG_10__SCAN_IN), .C1(n3996), .C2(
        DATAO_REG_8__SCAN_IN), .A(n3995), .ZN(n4003) );
  INV_X1 U4689 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4303) );
  AOI22_X1 U4690 ( .A1(n4303), .A2(keyinput35), .B1(U3149), .B2(keyinput14), 
        .ZN(n3997) );
  OAI221_X1 U4691 ( .B1(n4303), .B2(keyinput35), .C1(U3149), .C2(keyinput14), 
        .A(n3997), .ZN(n4002) );
  INV_X1 U4692 ( .A(REG2_REG_25__SCAN_IN), .ZN(n3998) );
  XOR2_X1 U4693 ( .A(n3998), .B(keyinput30), .Z(n4000) );
  XNOR2_X1 U4694 ( .A(IR_REG_27__SCAN_IN), .B(keyinput81), .ZN(n3999) );
  NAND2_X1 U4695 ( .A1(n4000), .A2(n3999), .ZN(n4001) );
  NOR4_X1 U4696 ( .A1(n4004), .A2(n4003), .A3(n4002), .A4(n4001), .ZN(n4047)
         );
  INV_X1 U4697 ( .A(keyinput38), .ZN(n4006) );
  AOI22_X1 U4698 ( .A1(n4627), .A2(keyinput7), .B1(ADDR_REG_13__SCAN_IN), .B2(
        n4006), .ZN(n4005) );
  OAI221_X1 U4699 ( .B1(n4627), .B2(keyinput7), .C1(n4006), .C2(
        ADDR_REG_13__SCAN_IN), .A(n4005), .ZN(n4016) );
  AOI22_X1 U4700 ( .A1(n3065), .A2(keyinput18), .B1(n2271), .B2(keyinput19), 
        .ZN(n4007) );
  OAI221_X1 U4701 ( .B1(n3065), .B2(keyinput18), .C1(n2271), .C2(keyinput19), 
        .A(n4007), .ZN(n4015) );
  INV_X1 U4702 ( .A(DATAI_24_), .ZN(n4010) );
  INV_X1 U4703 ( .A(DATAI_22_), .ZN(n4009) );
  AOI22_X1 U4704 ( .A1(n4010), .A2(keyinput58), .B1(n4009), .B2(keyinput3), 
        .ZN(n4008) );
  OAI221_X1 U4705 ( .B1(n4010), .B2(keyinput58), .C1(n4009), .C2(keyinput3), 
        .A(n4008), .ZN(n4014) );
  XNOR2_X1 U4706 ( .A(REG1_REG_1__SCAN_IN), .B(keyinput6), .ZN(n4012) );
  XNOR2_X1 U4707 ( .A(REG1_REG_0__SCAN_IN), .B(keyinput15), .ZN(n4011) );
  NAND2_X1 U4708 ( .A1(n4012), .A2(n4011), .ZN(n4013) );
  NOR4_X1 U4709 ( .A1(n4016), .A2(n4015), .A3(n4014), .A4(n4013), .ZN(n4046)
         );
  INV_X1 U4710 ( .A(D_REG_25__SCAN_IN), .ZN(n4831) );
  INV_X1 U4711 ( .A(D_REG_3__SCAN_IN), .ZN(n4840) );
  AOI22_X1 U4712 ( .A1(n4831), .A2(keyinput23), .B1(keyinput54), .B2(n4840), 
        .ZN(n4017) );
  OAI221_X1 U4713 ( .B1(n4831), .B2(keyinput23), .C1(n4840), .C2(keyinput54), 
        .A(n4017), .ZN(n4027) );
  INV_X1 U4714 ( .A(keyinput10), .ZN(n4019) );
  AOI22_X1 U4715 ( .A1(n4020), .A2(keyinput39), .B1(ADDR_REG_18__SCAN_IN), 
        .B2(n4019), .ZN(n4018) );
  OAI221_X1 U4716 ( .B1(n4020), .B2(keyinput39), .C1(n4019), .C2(
        ADDR_REG_18__SCAN_IN), .A(n4018), .ZN(n4026) );
  INV_X1 U4717 ( .A(D_REG_16__SCAN_IN), .ZN(n4833) );
  INV_X1 U4718 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4671) );
  AOI22_X1 U4719 ( .A1(n4833), .A2(keyinput59), .B1(keyinput63), .B2(n4671), 
        .ZN(n4021) );
  OAI221_X1 U4720 ( .B1(n4833), .B2(keyinput59), .C1(n4671), .C2(keyinput63), 
        .A(n4021), .ZN(n4025) );
  INV_X1 U4721 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4877) );
  XOR2_X1 U4722 ( .A(n4877), .B(keyinput31), .Z(n4023) );
  XNOR2_X1 U4723 ( .A(IR_REG_20__SCAN_IN), .B(keyinput27), .ZN(n4022) );
  NAND2_X1 U4724 ( .A1(n4023), .A2(n4022), .ZN(n4024) );
  NOR4_X1 U4725 ( .A1(n4027), .A2(n4026), .A3(n4025), .A4(n4024), .ZN(n4045)
         );
  INV_X1 U4726 ( .A(keyinput11), .ZN(n4029) );
  AOI22_X1 U4727 ( .A1(n4030), .A2(keyinput43), .B1(DATAO_REG_26__SCAN_IN), 
        .B2(n4029), .ZN(n4028) );
  OAI221_X1 U4728 ( .B1(n4030), .B2(keyinput43), .C1(n4029), .C2(
        DATAO_REG_26__SCAN_IN), .A(n4028), .ZN(n4043) );
  AOI22_X1 U4729 ( .A1(n4033), .A2(keyinput2), .B1(keyinput34), .B2(n4032), 
        .ZN(n4031) );
  OAI221_X1 U4730 ( .B1(n4033), .B2(keyinput2), .C1(n4032), .C2(keyinput34), 
        .A(n4031), .ZN(n4042) );
  AOI22_X1 U4731 ( .A1(n4036), .A2(keyinput26), .B1(n4035), .B2(keyinput51), 
        .ZN(n4034) );
  OAI221_X1 U4732 ( .B1(n4036), .B2(keyinput26), .C1(n4035), .C2(keyinput51), 
        .A(n4034), .ZN(n4041) );
  AOI22_X1 U4733 ( .A1(n4039), .A2(keyinput47), .B1(keyinput42), .B2(n4038), 
        .ZN(n4037) );
  OAI221_X1 U4734 ( .B1(n4039), .B2(keyinput47), .C1(n4038), .C2(keyinput42), 
        .A(n4037), .ZN(n4040) );
  NOR4_X1 U4735 ( .A1(n4043), .A2(n4042), .A3(n4041), .A4(n4040), .ZN(n4044)
         );
  NAND4_X1 U4736 ( .A1(n4047), .A2(n4046), .A3(n4045), .A4(n4044), .ZN(n4231)
         );
  INV_X1 U4737 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4049) );
  AOI22_X1 U4738 ( .A1(n4050), .A2(keyinput70), .B1(keyinput67), .B2(n4049), 
        .ZN(n4048) );
  OAI221_X1 U4739 ( .B1(n4050), .B2(keyinput70), .C1(n4049), .C2(keyinput67), 
        .A(n4048), .ZN(n4061) );
  INV_X1 U4740 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4578) );
  INV_X1 U4741 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4052) );
  AOI22_X1 U4742 ( .A1(n4578), .A2(keyinput75), .B1(n4052), .B2(keyinput71), 
        .ZN(n4051) );
  OAI221_X1 U4743 ( .B1(n4578), .B2(keyinput75), .C1(n4052), .C2(keyinput71), 
        .A(n4051), .ZN(n4060) );
  INV_X1 U4744 ( .A(keyinput79), .ZN(n4053) );
  XNOR2_X1 U4745 ( .A(n4053), .B(DATAO_REG_4__SCAN_IN), .ZN(n4059) );
  INV_X1 U4746 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4054) );
  XOR2_X1 U4747 ( .A(n4054), .B(keyinput74), .Z(n4057) );
  XNOR2_X1 U4748 ( .A(IR_REG_28__SCAN_IN), .B(keyinput78), .ZN(n4056) );
  XNOR2_X1 U4749 ( .A(IR_REG_7__SCAN_IN), .B(keyinput82), .ZN(n4055) );
  NAND3_X1 U4750 ( .A1(n4057), .A2(n4056), .A3(n4055), .ZN(n4058) );
  NOR4_X1 U4751 ( .A1(n4061), .A2(n4060), .A3(n4059), .A4(n4058), .ZN(n4229)
         );
  INV_X1 U4752 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4650) );
  AOI22_X1 U4753 ( .A1(n4650), .A2(keyinput90), .B1(keyinput87), .B2(n2548), 
        .ZN(n4062) );
  OAI221_X1 U4754 ( .B1(n4650), .B2(keyinput90), .C1(n2548), .C2(keyinput87), 
        .A(n4062), .ZN(n4075) );
  INV_X1 U4755 ( .A(keyinput99), .ZN(n4064) );
  AOI22_X1 U4756 ( .A1(n4065), .A2(keyinput94), .B1(DATAO_REG_29__SCAN_IN), 
        .B2(n4064), .ZN(n4063) );
  OAI221_X1 U4757 ( .B1(n4065), .B2(keyinput94), .C1(n4064), .C2(
        DATAO_REG_29__SCAN_IN), .A(n4063), .ZN(n4074) );
  INV_X1 U4758 ( .A(REG0_REG_18__SCAN_IN), .ZN(n4068) );
  INV_X1 U4759 ( .A(REG2_REG_10__SCAN_IN), .ZN(n4067) );
  AOI22_X1 U4760 ( .A1(n4068), .A2(keyinput95), .B1(n4067), .B2(keyinput91), 
        .ZN(n4066) );
  OAI221_X1 U4761 ( .B1(n4068), .B2(keyinput95), .C1(n4067), .C2(keyinput91), 
        .A(n4066), .ZN(n4073) );
  XOR2_X1 U4762 ( .A(n4069), .B(keyinput83), .Z(n4071) );
  XNOR2_X1 U4763 ( .A(IR_REG_5__SCAN_IN), .B(keyinput86), .ZN(n4070) );
  NAND2_X1 U4764 ( .A1(n4071), .A2(n4070), .ZN(n4072) );
  NOR4_X1 U4765 ( .A1(n4075), .A2(n4074), .A3(n4073), .A4(n4072), .ZN(n4228)
         );
  INV_X1 U4766 ( .A(keyinput126), .ZN(n4079) );
  INV_X1 U4767 ( .A(D_REG_20__SCAN_IN), .ZN(n4832) );
  AOI22_X1 U4768 ( .A1(n4832), .A2(keyinput127), .B1(keyinput122), .B2(n4077), 
        .ZN(n4076) );
  OAI221_X1 U4769 ( .B1(n4832), .B2(keyinput127), .C1(n4077), .C2(keyinput122), 
        .A(n4076), .ZN(n4078) );
  AOI221_X1 U4770 ( .B1(REG1_REG_9__SCAN_IN), .B2(n4079), .C1(n2599), .C2(
        keyinput126), .A(n4078), .ZN(n4093) );
  INV_X1 U4771 ( .A(keyinput110), .ZN(n4081) );
  AOI22_X1 U4772 ( .A1(n2573), .A2(keyinput107), .B1(ADDR_REG_12__SCAN_IN), 
        .B2(n4081), .ZN(n4080) );
  OAI221_X1 U4773 ( .B1(n2573), .B2(keyinput107), .C1(n4081), .C2(
        ADDR_REG_12__SCAN_IN), .A(n4080), .ZN(n4091) );
  INV_X1 U4774 ( .A(REG3_REG_1__SCAN_IN), .ZN(n4083) );
  AOI22_X1 U4775 ( .A1(n4084), .A2(keyinput114), .B1(keyinput111), .B2(n4083), 
        .ZN(n4082) );
  OAI221_X1 U4776 ( .B1(n4084), .B2(keyinput114), .C1(n4083), .C2(keyinput111), 
        .A(n4082), .ZN(n4090) );
  INV_X1 U4777 ( .A(DATAI_14_), .ZN(n4853) );
  AOI22_X1 U4778 ( .A1(n4853), .A2(keyinput103), .B1(keyinput98), .B2(n3417), 
        .ZN(n4085) );
  OAI221_X1 U4779 ( .B1(n4853), .B2(keyinput103), .C1(n3417), .C2(keyinput98), 
        .A(n4085), .ZN(n4089) );
  INV_X1 U4780 ( .A(DATAI_1_), .ZN(n4087) );
  AOI22_X1 U4781 ( .A1(n2619), .A2(keyinput106), .B1(keyinput102), .B2(n4087), 
        .ZN(n4086) );
  OAI221_X1 U4782 ( .B1(n2619), .B2(keyinput106), .C1(n4087), .C2(keyinput102), 
        .A(n4086), .ZN(n4088) );
  NOR4_X1 U4783 ( .A1(n4091), .A2(n4090), .A3(n4089), .A4(n4088), .ZN(n4092)
         );
  OAI211_X1 U4784 ( .C1(keyinput46), .C2(n2498), .A(n4093), .B(n4092), .ZN(
        n4118) );
  AOI22_X1 U4785 ( .A1(n4095), .A2(keyinput0), .B1(keyinput112), .B2(n2542), 
        .ZN(n4094) );
  OAI221_X1 U4786 ( .B1(n4095), .B2(keyinput0), .C1(n2542), .C2(keyinput112), 
        .A(n4094), .ZN(n4100) );
  INV_X1 U4787 ( .A(keyinput119), .ZN(n4097) );
  AOI22_X1 U4788 ( .A1(n4098), .A2(keyinput115), .B1(DATAO_REG_27__SCAN_IN), 
        .B2(n4097), .ZN(n4096) );
  OAI221_X1 U4789 ( .B1(n4098), .B2(keyinput115), .C1(n4097), .C2(
        DATAO_REG_27__SCAN_IN), .A(n4096), .ZN(n4099) );
  NOR2_X1 U4790 ( .A1(n4100), .A2(n4099), .ZN(n4116) );
  INV_X1 U4791 ( .A(keyinput120), .ZN(n4101) );
  XNOR2_X1 U4792 ( .A(n4101), .B(ADDR_REG_1__SCAN_IN), .ZN(n4105) );
  XNOR2_X1 U4793 ( .A(IR_REG_24__SCAN_IN), .B(keyinput24), .ZN(n4103) );
  XNOR2_X1 U4794 ( .A(keyinput104), .B(REG2_REG_9__SCAN_IN), .ZN(n4102) );
  NAND2_X1 U4795 ( .A1(n4103), .A2(n4102), .ZN(n4104) );
  NOR2_X1 U4796 ( .A1(n4105), .A2(n4104), .ZN(n4115) );
  INV_X1 U4797 ( .A(keyinput116), .ZN(n4107) );
  AOI22_X1 U4798 ( .A1(n4108), .A2(keyinput124), .B1(DATAO_REG_9__SCAN_IN), 
        .B2(n4107), .ZN(n4106) );
  OAI221_X1 U4799 ( .B1(n4108), .B2(keyinput124), .C1(n4107), .C2(
        DATAO_REG_9__SCAN_IN), .A(n4106), .ZN(n4113) );
  XNOR2_X1 U4800 ( .A(IR_REG_31__SCAN_IN), .B(keyinput64), .ZN(n4111) );
  XNOR2_X1 U4801 ( .A(REG1_REG_28__SCAN_IN), .B(keyinput123), .ZN(n4110) );
  XNOR2_X1 U4802 ( .A(IR_REG_10__SCAN_IN), .B(keyinput118), .ZN(n4109) );
  NAND3_X1 U4803 ( .A1(n4111), .A2(n4110), .A3(n4109), .ZN(n4112) );
  NOR2_X1 U4804 ( .A1(n4113), .A2(n4112), .ZN(n4114) );
  NAND3_X1 U4805 ( .A1(n4116), .A2(n4115), .A3(n4114), .ZN(n4117) );
  NOR2_X1 U4806 ( .A1(n4118), .A2(n4117), .ZN(n4160) );
  INV_X1 U4807 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4680) );
  INV_X1 U4808 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n4120) );
  AOI22_X1 U4809 ( .A1(n4680), .A2(keyinput84), .B1(keyinput72), .B2(n4120), 
        .ZN(n4119) );
  OAI221_X1 U4810 ( .B1(n4680), .B2(keyinput84), .C1(n4120), .C2(keyinput72), 
        .A(n4119), .ZN(n4132) );
  INV_X1 U4811 ( .A(D_REG_10__SCAN_IN), .ZN(n4836) );
  AOI22_X1 U4812 ( .A1(n4836), .A2(keyinput96), .B1(keyinput92), .B2(n4122), 
        .ZN(n4121) );
  OAI221_X1 U4813 ( .B1(n4836), .B2(keyinput96), .C1(n4122), .C2(keyinput92), 
        .A(n4121), .ZN(n4131) );
  INV_X1 U4814 ( .A(DATAI_2_), .ZN(n4125) );
  INV_X1 U4815 ( .A(ADDR_REG_11__SCAN_IN), .ZN(n4124) );
  AOI22_X1 U4816 ( .A1(n4125), .A2(keyinput108), .B1(keyinput80), .B2(n4124), 
        .ZN(n4123) );
  OAI221_X1 U4817 ( .B1(n4125), .B2(keyinput108), .C1(n4124), .C2(keyinput80), 
        .A(n4123), .ZN(n4130) );
  INV_X1 U4818 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4128) );
  INV_X1 U4819 ( .A(ADDR_REG_15__SCAN_IN), .ZN(n4127) );
  AOI22_X1 U4820 ( .A1(n4128), .A2(keyinput76), .B1(keyinput100), .B2(n4127), 
        .ZN(n4126) );
  OAI221_X1 U4821 ( .B1(n4128), .B2(keyinput76), .C1(n4127), .C2(keyinput100), 
        .A(n4126), .ZN(n4129) );
  NOR4_X1 U4822 ( .A1(n4132), .A2(n4131), .A3(n4130), .A4(n4129), .ZN(n4159)
         );
  INV_X1 U4823 ( .A(D_REG_5__SCAN_IN), .ZN(n4839) );
  AOI22_X1 U4824 ( .A1(n2670), .A2(keyinput20), .B1(keyinput4), .B2(n4839), 
        .ZN(n4133) );
  OAI221_X1 U4825 ( .B1(n2670), .B2(keyinput20), .C1(n4839), .C2(keyinput4), 
        .A(n4133), .ZN(n4143) );
  INV_X1 U4826 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4893) );
  AOI22_X1 U4827 ( .A1(n4135), .A2(keyinput56), .B1(keyinput8), .B2(n4893), 
        .ZN(n4134) );
  OAI221_X1 U4828 ( .B1(n4135), .B2(keyinput56), .C1(n4893), .C2(keyinput8), 
        .A(n4134), .ZN(n4142) );
  INV_X1 U4829 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4658) );
  AOI22_X1 U4830 ( .A1(n2678), .A2(keyinput36), .B1(keyinput28), .B2(n4658), 
        .ZN(n4136) );
  OAI221_X1 U4831 ( .B1(n2678), .B2(keyinput36), .C1(n4658), .C2(keyinput28), 
        .A(n4136), .ZN(n4141) );
  INV_X1 U4832 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4138) );
  AOI22_X1 U4833 ( .A1(n4139), .A2(keyinput12), .B1(keyinput16), .B2(n4138), 
        .ZN(n4137) );
  OAI221_X1 U4834 ( .B1(n4139), .B2(keyinput12), .C1(n4138), .C2(keyinput16), 
        .A(n4137), .ZN(n4140) );
  NOR4_X1 U4835 ( .A1(n4143), .A2(n4142), .A3(n4141), .A4(n4140), .ZN(n4158)
         );
  AOI22_X1 U4836 ( .A1(n4145), .A2(keyinput52), .B1(n2636), .B2(keyinput40), 
        .ZN(n4144) );
  OAI221_X1 U4837 ( .B1(n4145), .B2(keyinput52), .C1(n2636), .C2(keyinput40), 
        .A(n4144), .ZN(n4156) );
  INV_X1 U4838 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4147) );
  INV_X1 U4839 ( .A(DATAI_15_), .ZN(n4851) );
  AOI22_X1 U4840 ( .A1(n4147), .A2(keyinput66), .B1(keyinput60), .B2(n4851), 
        .ZN(n4146) );
  OAI221_X1 U4841 ( .B1(n4147), .B2(keyinput66), .C1(n4851), .C2(keyinput60), 
        .A(n4146), .ZN(n4155) );
  INV_X1 U4842 ( .A(DATAI_26_), .ZN(n4150) );
  INV_X1 U4843 ( .A(keyinput48), .ZN(n4149) );
  AOI22_X1 U4844 ( .A1(n4150), .A2(keyinput68), .B1(DATAO_REG_25__SCAN_IN), 
        .B2(n4149), .ZN(n4148) );
  OAI221_X1 U4845 ( .B1(n4150), .B2(keyinput68), .C1(n4149), .C2(
        DATAO_REG_25__SCAN_IN), .A(n4148), .ZN(n4154) );
  INV_X1 U4846 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4887) );
  INV_X1 U4847 ( .A(keyinput32), .ZN(n4152) );
  AOI22_X1 U4848 ( .A1(n4887), .A2(keyinput44), .B1(ADDR_REG_3__SCAN_IN), .B2(
        n4152), .ZN(n4151) );
  OAI221_X1 U4849 ( .B1(n4887), .B2(keyinput44), .C1(n4152), .C2(
        ADDR_REG_3__SCAN_IN), .A(n4151), .ZN(n4153) );
  NOR4_X1 U4850 ( .A1(n4156), .A2(n4155), .A3(n4154), .A4(n4153), .ZN(n4157)
         );
  AND4_X1 U4851 ( .A1(n4160), .A2(n4159), .A3(n4158), .A4(n4157), .ZN(n4227)
         );
  INV_X1 U4852 ( .A(keyinput127), .ZN(n4161) );
  NAND4_X1 U4853 ( .A1(keyinput126), .A2(keyinput118), .A3(keyinput119), .A4(
        n4161), .ZN(n4162) );
  NOR4_X1 U4854 ( .A1(keyinput47), .A2(keyinput122), .A3(keyinput123), .A4(
        n4162), .ZN(n4174) );
  INV_X1 U4855 ( .A(keyinput102), .ZN(n4163) );
  NOR4_X1 U4856 ( .A1(keyinput107), .A2(keyinput106), .A3(keyinput103), .A4(
        n4163), .ZN(n4173) );
  NAND2_X1 U4857 ( .A1(keyinput111), .A2(keyinput115), .ZN(n4164) );
  NOR3_X1 U4858 ( .A1(keyinput114), .A2(keyinput110), .A3(n4164), .ZN(n4172)
         );
  NOR2_X1 U4859 ( .A1(keyinput94), .A2(keyinput87), .ZN(n4165) );
  NAND3_X1 U4860 ( .A1(keyinput95), .A2(keyinput86), .A3(n4165), .ZN(n4170) );
  NAND4_X1 U4861 ( .A1(keyinput98), .A2(keyinput99), .A3(keyinput91), .A4(
        keyinput90), .ZN(n4169) );
  NAND4_X1 U4862 ( .A1(keyinput79), .A2(keyinput78), .A3(keyinput71), .A4(
        keyinput70), .ZN(n4168) );
  NOR2_X1 U4863 ( .A1(keyinput83), .A2(keyinput74), .ZN(n4166) );
  NAND3_X1 U4864 ( .A1(keyinput82), .A2(keyinput75), .A3(n4166), .ZN(n4167) );
  NOR4_X1 U4865 ( .A1(n4170), .A2(n4169), .A3(n4168), .A4(n4167), .ZN(n4171)
         );
  NAND4_X1 U4866 ( .A1(n4174), .A2(n4173), .A3(n4172), .A4(n4171), .ZN(n4224)
         );
  NOR4_X1 U4867 ( .A1(keyinput109), .A2(keyinput105), .A3(keyinput97), .A4(
        keyinput101), .ZN(n4181) );
  NAND3_X1 U4868 ( .A1(keyinput121), .A2(keyinput125), .A3(keyinput21), .ZN(
        n4175) );
  NOR2_X1 U4869 ( .A1(keyinput17), .A2(n4175), .ZN(n4180) );
  INV_X1 U4870 ( .A(keyinput69), .ZN(n4176) );
  NOR4_X1 U4871 ( .A1(keyinput65), .A2(keyinput89), .A3(keyinput93), .A4(n4176), .ZN(n4179) );
  NAND3_X1 U4872 ( .A1(keyinput73), .A2(keyinput77), .A3(keyinput113), .ZN(
        n4177) );
  NOR2_X1 U4873 ( .A1(keyinput117), .A2(n4177), .ZN(n4178) );
  NAND4_X1 U4874 ( .A1(n4181), .A2(n4180), .A3(n4179), .A4(n4178), .ZN(n4223)
         );
  NAND2_X1 U4875 ( .A1(keyinput57), .A2(keyinput33), .ZN(n4182) );
  NOR3_X1 U4876 ( .A1(keyinput37), .A2(keyinput61), .A3(n4182), .ZN(n4188) );
  INV_X1 U4877 ( .A(keyinput45), .ZN(n4183) );
  NOR4_X1 U4878 ( .A1(keyinput80), .A2(keyinput88), .A3(keyinput41), .A4(n4183), .ZN(n4187) );
  NOR4_X1 U4879 ( .A1(keyinput5), .A2(keyinput1), .A3(keyinput13), .A4(
        keyinput9), .ZN(n4186) );
  NAND3_X1 U4880 ( .A1(keyinput29), .A2(keyinput25), .A3(keyinput49), .ZN(
        n4184) );
  NOR2_X1 U4881 ( .A1(keyinput53), .A2(n4184), .ZN(n4185) );
  NAND4_X1 U4882 ( .A1(n4188), .A2(n4187), .A3(n4186), .A4(n4185), .ZN(n4222)
         );
  NOR3_X1 U4883 ( .A1(keyinput64), .A2(keyinput0), .A3(keyinput104), .ZN(n4189) );
  NAND2_X1 U4884 ( .A1(keyinput116), .A2(n4189), .ZN(n4196) );
  NOR2_X1 U4885 ( .A1(keyinput28), .A2(keyinput120), .ZN(n4190) );
  NAND3_X1 U4886 ( .A1(keyinput24), .A2(keyinput124), .A3(n4190), .ZN(n4195)
         );
  NOR2_X1 U4887 ( .A1(keyinput100), .A2(keyinput76), .ZN(n4191) );
  NAND3_X1 U4888 ( .A1(keyinput72), .A2(keyinput108), .A3(n4191), .ZN(n4194)
         );
  NOR2_X1 U4889 ( .A1(keyinput112), .A2(keyinput84), .ZN(n4192) );
  NAND3_X1 U4890 ( .A1(keyinput96), .A2(keyinput92), .A3(n4192), .ZN(n4193) );
  NOR4_X1 U4891 ( .A1(n4196), .A2(n4195), .A3(n4194), .A4(n4193), .ZN(n4220)
         );
  NOR2_X1 U4892 ( .A1(keyinput44), .A2(keyinput68), .ZN(n4197) );
  NAND3_X1 U4893 ( .A1(keyinput40), .A2(keyinput32), .A3(n4197), .ZN(n4202) );
  INV_X1 U4894 ( .A(keyinput60), .ZN(n4198) );
  NAND4_X1 U4895 ( .A1(keyinput66), .A2(keyinput67), .A3(keyinput52), .A4(
        n4198), .ZN(n4201) );
  NAND4_X1 U4896 ( .A1(keyinput4), .A2(keyinput12), .A3(keyinput16), .A4(
        keyinput36), .ZN(n4200) );
  NAND4_X1 U4897 ( .A1(keyinput48), .A2(keyinput56), .A3(keyinput8), .A4(
        keyinput20), .ZN(n4199) );
  NOR4_X1 U4898 ( .A1(n4202), .A2(n4201), .A3(n4200), .A4(n4199), .ZN(n4219)
         );
  NOR2_X1 U4899 ( .A1(keyinput27), .A2(keyinput59), .ZN(n4203) );
  NAND3_X1 U4900 ( .A1(keyinput23), .A2(keyinput54), .A3(n4203), .ZN(n4209) );
  NAND4_X1 U4901 ( .A1(keyinput6), .A2(keyinput10), .A3(keyinput39), .A4(
        keyinput31), .ZN(n4208) );
  NOR2_X1 U4902 ( .A1(keyinput34), .A2(keyinput51), .ZN(n4204) );
  NAND3_X1 U4903 ( .A1(keyinput26), .A2(keyinput42), .A3(n4204), .ZN(n4207) );
  NOR2_X1 U4904 ( .A1(keyinput11), .A2(keyinput2), .ZN(n4205) );
  NAND3_X1 U4905 ( .A1(keyinput63), .A2(keyinput43), .A3(n4205), .ZN(n4206) );
  NOR4_X1 U4906 ( .A1(n4209), .A2(n4208), .A3(n4207), .A4(n4206), .ZN(n4218)
         );
  NAND4_X1 U4907 ( .A1(keyinput14), .A2(keyinput55), .A3(keyinput62), .A4(
        n4210), .ZN(n4216) );
  NOR2_X1 U4908 ( .A1(keyinput85), .A2(keyinput30), .ZN(n4211) );
  NAND3_X1 U4909 ( .A1(keyinput81), .A2(keyinput35), .A3(n4211), .ZN(n4215) );
  INV_X1 U4910 ( .A(keyinput7), .ZN(n4212) );
  NAND4_X1 U4911 ( .A1(keyinput38), .A2(keyinput19), .A3(keyinput15), .A4(
        n4212), .ZN(n4214) );
  NAND4_X1 U4912 ( .A1(keyinput50), .A2(keyinput58), .A3(keyinput3), .A4(
        keyinput18), .ZN(n4213) );
  NOR4_X1 U4913 ( .A1(n4216), .A2(n4215), .A3(n4214), .A4(n4213), .ZN(n4217)
         );
  NAND4_X1 U4914 ( .A1(n4220), .A2(n4219), .A3(n4218), .A4(n4217), .ZN(n4221)
         );
  NOR4_X1 U4915 ( .A1(n4224), .A2(n4223), .A3(n4222), .A4(n4221), .ZN(n4225)
         );
  OAI21_X1 U4916 ( .B1(keyinput46), .B2(n4225), .A(n2498), .ZN(n4226) );
  NAND4_X1 U4917 ( .A1(n4229), .A2(n4228), .A3(n4227), .A4(n4226), .ZN(n4230)
         );
  NOR3_X1 U4918 ( .A1(n4232), .A2(n4231), .A3(n4230), .ZN(n4233) );
  XOR2_X1 U4919 ( .A(n4234), .B(n4233), .Z(U3564) );
  MUX2_X1 U4920 ( .A(n4235), .B(DATAO_REG_12__SCAN_IN), .S(n4240), .Z(U3562)
         );
  MUX2_X1 U4921 ( .A(n4236), .B(DATAO_REG_7__SCAN_IN), .S(n4240), .Z(U3557) );
  MUX2_X1 U4922 ( .A(n4237), .B(DATAO_REG_5__SCAN_IN), .S(n4240), .Z(U3555) );
  MUX2_X1 U4923 ( .A(n4238), .B(DATAO_REG_3__SCAN_IN), .S(n4240), .Z(U3553) );
  MUX2_X1 U4924 ( .A(n4239), .B(DATAO_REG_1__SCAN_IN), .S(n4240), .Z(U3551) );
  MUX2_X1 U4925 ( .A(n2944), .B(DATAO_REG_0__SCAN_IN), .S(n4240), .Z(U3550) );
  NOR2_X1 U4926 ( .A1(n2419), .A2(n3071), .ZN(n4252) );
  MUX2_X1 U4927 ( .A(REG2_REG_1__SCAN_IN), .B(n3070), .S(n4699), .Z(n4242) );
  INV_X1 U4928 ( .A(n4241), .ZN(n4263) );
  OAI211_X1 U4929 ( .C1(n4252), .C2(n4242), .A(n4809), .B(n4263), .ZN(n4249)
         );
  AOI22_X1 U4930 ( .A1(n4775), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4248) );
  NAND2_X1 U4931 ( .A1(n4758), .A2(n4699), .ZN(n4247) );
  OAI211_X1 U4932 ( .C1(n4245), .C2(n4244), .A(n4794), .B(n4243), .ZN(n4246)
         );
  NAND4_X1 U4933 ( .A1(n4249), .A2(n4248), .A3(n4247), .A4(n4246), .ZN(U3241)
         );
  NAND2_X1 U4934 ( .A1(n4250), .A2(n4318), .ZN(n4257) );
  INV_X1 U4935 ( .A(n4251), .ZN(n4253) );
  AOI22_X1 U4936 ( .A1(n4254), .A2(n2419), .B1(n4253), .B2(n4252), .ZN(n4255)
         );
  OAI211_X1 U4937 ( .C1(n4258), .C2(n4257), .A(U4043), .B(n4255), .ZN(n4279)
         );
  AOI22_X1 U4938 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4775), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n4270) );
  XNOR2_X1 U4939 ( .A(n4260), .B(n4259), .ZN(n4261) );
  AOI22_X1 U4940 ( .A1(n4698), .A2(n4758), .B1(n4794), .B2(n4261), .ZN(n4269)
         );
  MUX2_X1 U4941 ( .A(n3075), .B(REG2_REG_2__SCAN_IN), .S(n4698), .Z(n4265) );
  INV_X1 U4942 ( .A(n4262), .ZN(n4264) );
  NAND3_X1 U4943 ( .A1(n4265), .A2(n4264), .A3(n4263), .ZN(n4266) );
  NAND3_X1 U4944 ( .A1(n4809), .A2(n4267), .A3(n4266), .ZN(n4268) );
  NAND4_X1 U4945 ( .A1(n4279), .A2(n4270), .A3(n4269), .A4(n4268), .ZN(U3242)
         );
  XNOR2_X1 U4946 ( .A(n4271), .B(REG1_REG_4__SCAN_IN), .ZN(n4277) );
  XNOR2_X1 U4947 ( .A(n4272), .B(REG2_REG_4__SCAN_IN), .ZN(n4275) );
  NAND2_X1 U4948 ( .A1(n4758), .A2(n4696), .ZN(n4273) );
  OAI211_X1 U4949 ( .C1(n4751), .C2(n4275), .A(n4274), .B(n4273), .ZN(n4276)
         );
  AOI21_X1 U4950 ( .B1(n4794), .B2(n4277), .A(n4276), .ZN(n4280) );
  NAND2_X1 U4951 ( .A1(n4775), .A2(ADDR_REG_4__SCAN_IN), .ZN(n4278) );
  NAND3_X1 U4952 ( .A1(n4280), .A2(n4279), .A3(n4278), .ZN(U3244) );
  INV_X1 U4953 ( .A(n4302), .ZN(n4846) );
  AOI22_X1 U4954 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4846), .B1(n4302), .B2(
        n4281), .ZN(n4798) );
  AOI22_X1 U4955 ( .A1(n4301), .A2(REG1_REG_17__SCAN_IN), .B1(n4627), .B2(
        n4848), .ZN(n4788) );
  NOR2_X1 U4956 ( .A1(n4284), .A2(n2282), .ZN(n4285) );
  NOR2_X1 U4957 ( .A1(n4750), .A2(n4749), .ZN(n4748) );
  INV_X1 U4958 ( .A(n4298), .ZN(n4852) );
  AOI22_X1 U4959 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4852), .B1(n4298), .B2(
        n4286), .ZN(n4763) );
  NAND2_X1 U4960 ( .A1(n4287), .A2(n4850), .ZN(n4288) );
  NAND2_X1 U4961 ( .A1(n4288), .A2(n4776), .ZN(n4787) );
  NAND2_X1 U4962 ( .A1(n4788), .A2(n4787), .ZN(n4786) );
  OAI21_X1 U4963 ( .B1(n4301), .B2(REG1_REG_17__SCAN_IN), .A(n4786), .ZN(n4799) );
  XNOR2_X1 U4964 ( .A(n4691), .B(REG1_REG_19__SCAN_IN), .ZN(n4289) );
  NAND2_X1 U4965 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4302), .ZN(n4290) );
  OAI21_X1 U4966 ( .B1(REG2_REG_18__SCAN_IN), .B2(n4302), .A(n4290), .ZN(n4807) );
  NOR2_X1 U4967 ( .A1(n4301), .A2(REG2_REG_17__SCAN_IN), .ZN(n4291) );
  AOI21_X1 U4968 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4301), .A(n4291), .ZN(n4791) );
  NOR2_X1 U4969 ( .A1(n2282), .A2(n4295), .ZN(n4296) );
  NOR2_X1 U4970 ( .A1(n4296), .A2(n4752), .ZN(n4768) );
  INV_X1 U4971 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4297) );
  AOI22_X1 U4972 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4852), .B1(n4298), .B2(
        n4297), .ZN(n4769) );
  NOR2_X1 U4973 ( .A1(n4768), .A2(n4769), .ZN(n4767) );
  NAND2_X1 U4974 ( .A1(n4299), .A2(n4850), .ZN(n4300) );
  NAND2_X1 U4975 ( .A1(n4791), .A2(n4790), .ZN(n4789) );
  MUX2_X1 U4976 ( .A(REG2_REG_19__SCAN_IN), .B(n4303), .S(n4691), .Z(n4304) );
  AOI21_X1 U4977 ( .B1(n4775), .B2(ADDR_REG_19__SCAN_IN), .A(n4305), .ZN(n4306) );
  OAI21_X1 U4978 ( .B1(n4812), .B2(n4307), .A(n4306), .ZN(n4308) );
  AOI21_X1 U4979 ( .B1(n4309), .B2(n4809), .A(n4308), .ZN(n4310) );
  INV_X1 U4980 ( .A(n4311), .ZN(n4324) );
  INV_X1 U4981 ( .A(n4329), .ZN(n4317) );
  INV_X1 U4982 ( .A(n4312), .ZN(n4314) );
  AOI21_X1 U4983 ( .B1(n4315), .B2(n4314), .A(n4313), .ZN(n4316) );
  XOR2_X1 U4984 ( .A(n4317), .B(n4316), .Z(n4323) );
  INV_X1 U4985 ( .A(B_REG_SCAN_IN), .ZN(n4319) );
  OAI21_X1 U4986 ( .B1(n4319), .B2(n4318), .A(n4525), .ZN(n4563) );
  OAI22_X1 U4987 ( .A1(n4320), .A2(n4563), .B1(n4332), .B2(n4565), .ZN(n4321)
         );
  AOI21_X1 U4988 ( .B1(n4342), .B2(n4545), .A(n4321), .ZN(n4322) );
  OAI21_X1 U4989 ( .B1(n4323), .B2(n4547), .A(n4322), .ZN(n4581) );
  AOI21_X1 U4990 ( .B1(n4324), .B2(n4826), .A(n4581), .ZN(n4336) );
  XNOR2_X1 U4991 ( .A(n4330), .B(n4329), .ZN(n4580) );
  NAND2_X1 U4992 ( .A1(n4580), .A2(n4331), .ZN(n4335) );
  AOI21_X1 U4993 ( .B1(n4333), .B2(n2180), .A(n4570), .ZN(n4582) );
  AOI22_X1 U4994 ( .A1(n4582), .A2(n4817), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4813), .ZN(n4334) );
  OAI211_X1 U4995 ( .C1(n4813), .C2(n4336), .A(n4335), .B(n4334), .ZN(U3354)
         );
  XOR2_X1 U4996 ( .A(n4340), .B(n4337), .Z(n4588) );
  OAI21_X1 U4997 ( .B1(n4340), .B2(n4339), .A(n4338), .ZN(n4341) );
  NAND2_X1 U4998 ( .A1(n4341), .A2(n4531), .ZN(n4344) );
  AOI22_X1 U4999 ( .A1(n4342), .A2(n4525), .B1(n4576), .B2(n4347), .ZN(n4343)
         );
  OAI211_X1 U5000 ( .C1(n4345), .C2(n4528), .A(n4344), .B(n4343), .ZN(n4585)
         );
  AOI21_X1 U5001 ( .B1(n4347), .B2(n4364), .A(n4346), .ZN(n4586) );
  INV_X1 U5002 ( .A(n4586), .ZN(n4350) );
  AOI22_X1 U5003 ( .A1(n4813), .A2(REG2_REG_27__SCAN_IN), .B1(n4348), .B2(
        n4826), .ZN(n4349) );
  OAI21_X1 U5004 ( .B1(n4350), .B2(n4555), .A(n4349), .ZN(n4351) );
  AOI21_X1 U5005 ( .B1(n4585), .B2(n4557), .A(n4351), .ZN(n4352) );
  OAI21_X1 U5006 ( .B1(n4588), .B2(n4559), .A(n4352), .ZN(U3263) );
  XOR2_X1 U5007 ( .A(n4358), .B(n4353), .Z(n4590) );
  INV_X1 U5008 ( .A(n4590), .ZN(n4371) );
  INV_X1 U5009 ( .A(n4354), .ZN(n4356) );
  OAI21_X1 U5010 ( .B1(n4373), .B2(n4356), .A(n4355), .ZN(n4357) );
  XOR2_X1 U5011 ( .A(n4358), .B(n4357), .Z(n4363) );
  OAI22_X1 U5012 ( .A1(n4359), .A2(n4528), .B1(n4365), .B2(n4565), .ZN(n4360)
         );
  AOI21_X1 U5013 ( .B1(n4525), .B2(n4361), .A(n4360), .ZN(n4362) );
  OAI21_X1 U5014 ( .B1(n4363), .B2(n4547), .A(n4362), .ZN(n4589) );
  INV_X1 U5015 ( .A(n4384), .ZN(n4366) );
  OAI21_X1 U5016 ( .B1(n4366), .B2(n4365), .A(n4364), .ZN(n4652) );
  AOI22_X1 U5017 ( .A1(n4813), .A2(REG2_REG_26__SCAN_IN), .B1(n4367), .B2(
        n4826), .ZN(n4368) );
  OAI21_X1 U5018 ( .B1(n4652), .B2(n4555), .A(n4368), .ZN(n4369) );
  AOI21_X1 U5019 ( .B1(n4589), .B2(n4557), .A(n4369), .ZN(n4370) );
  OAI21_X1 U5020 ( .B1(n4371), .B2(n4559), .A(n4370), .ZN(U3264) );
  XNOR2_X1 U5021 ( .A(n4372), .B(n4375), .ZN(n4594) );
  INV_X1 U5022 ( .A(n4594), .ZN(n4390) );
  NAND2_X1 U5023 ( .A1(n2204), .A2(n4374), .ZN(n4376) );
  XNOR2_X1 U5024 ( .A(n4376), .B(n4375), .ZN(n4381) );
  AOI22_X1 U5025 ( .A1(n4420), .A2(n4545), .B1(n4377), .B2(n4576), .ZN(n4380)
         );
  NAND2_X1 U5026 ( .A1(n4378), .A2(n4525), .ZN(n4379) );
  OAI211_X1 U5027 ( .C1(n4381), .C2(n4547), .A(n4380), .B(n4379), .ZN(n4593)
         );
  OR2_X1 U5028 ( .A1(n4401), .A2(n4382), .ZN(n4383) );
  NAND2_X1 U5029 ( .A1(n4384), .A2(n4383), .ZN(n4656) );
  INV_X1 U5030 ( .A(n4385), .ZN(n4386) );
  AOI22_X1 U5031 ( .A1(n4813), .A2(REG2_REG_25__SCAN_IN), .B1(n4386), .B2(
        n4826), .ZN(n4387) );
  OAI21_X1 U5032 ( .B1(n4656), .B2(n4555), .A(n4387), .ZN(n4388) );
  AOI21_X1 U5033 ( .B1(n4593), .B2(n4557), .A(n4388), .ZN(n4389) );
  OAI21_X1 U5034 ( .B1(n4390), .B2(n4559), .A(n4389), .ZN(U3265) );
  XNOR2_X1 U5035 ( .A(n4391), .B(n4396), .ZN(n4598) );
  INV_X1 U5036 ( .A(n4598), .ZN(n4410) );
  INV_X1 U5037 ( .A(n4392), .ZN(n4393) );
  NOR2_X1 U5038 ( .A1(n4394), .A2(n4393), .ZN(n4395) );
  XOR2_X1 U5039 ( .A(n4396), .B(n4395), .Z(n4400) );
  OAI22_X1 U5040 ( .A1(n4440), .A2(n4528), .B1(n4403), .B2(n4565), .ZN(n4397)
         );
  AOI21_X1 U5041 ( .B1(n4525), .B2(n4398), .A(n4397), .ZN(n4399) );
  OAI21_X1 U5042 ( .B1(n4400), .B2(n4547), .A(n4399), .ZN(n4597) );
  INV_X1 U5043 ( .A(n4424), .ZN(n4404) );
  INV_X1 U5044 ( .A(n4401), .ZN(n4402) );
  OAI21_X1 U5045 ( .B1(n4404), .B2(n4403), .A(n4402), .ZN(n4660) );
  NOR2_X1 U5046 ( .A1(n4660), .A2(n4555), .ZN(n4408) );
  INV_X1 U5047 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4406) );
  OAI22_X1 U5048 ( .A1(n4557), .A2(n4406), .B1(n4405), .B2(n4519), .ZN(n4407)
         );
  AOI211_X1 U5049 ( .C1(n4597), .C2(n4557), .A(n4408), .B(n4407), .ZN(n4409)
         );
  OAI21_X1 U5050 ( .B1(n4410), .B2(n4559), .A(n4409), .ZN(U3266) );
  XOR2_X1 U5051 ( .A(n4416), .B(n4411), .Z(n4602) );
  INV_X1 U5052 ( .A(n4602), .ZN(n4431) );
  INV_X1 U5053 ( .A(n4412), .ZN(n4413) );
  OAI21_X1 U5054 ( .B1(n4452), .B2(n4414), .A(n4413), .ZN(n4435) );
  AND2_X1 U5055 ( .A1(n4435), .A2(n4434), .ZN(n4437) );
  NOR2_X1 U5056 ( .A1(n4437), .A2(n4415), .ZN(n4417) );
  XNOR2_X1 U5057 ( .A(n4417), .B(n4416), .ZN(n4418) );
  NAND2_X1 U5058 ( .A1(n4418), .A2(n4531), .ZN(n4422) );
  AOI22_X1 U5059 ( .A1(n4420), .A2(n4525), .B1(n4576), .B2(n4419), .ZN(n4421)
         );
  OAI211_X1 U5060 ( .C1(n4423), .C2(n4528), .A(n4422), .B(n4421), .ZN(n4601)
         );
  INV_X1 U5061 ( .A(n4606), .ZN(n4426) );
  OAI21_X1 U5062 ( .B1(n4426), .B2(n4425), .A(n4424), .ZN(n4664) );
  NOR2_X1 U5063 ( .A1(n4664), .A2(n4555), .ZN(n4429) );
  OAI22_X1 U5064 ( .A1(n4557), .A2(n4138), .B1(n4427), .B2(n4519), .ZN(n4428)
         );
  AOI211_X1 U5065 ( .C1(n4601), .C2(n4557), .A(n4429), .B(n4428), .ZN(n4430)
         );
  OAI21_X1 U5066 ( .B1(n4431), .B2(n4559), .A(n4430), .ZN(U3267) );
  OAI21_X1 U5067 ( .B1(n4433), .B2(n2934), .A(n4432), .ZN(n4609) );
  NOR2_X1 U5068 ( .A1(n4435), .A2(n4434), .ZN(n4436) );
  OR2_X1 U5069 ( .A1(n4437), .A2(n4436), .ZN(n4442) );
  NAND2_X1 U5070 ( .A1(n4445), .A2(n4576), .ZN(n4439) );
  NAND2_X1 U5071 ( .A1(n4473), .A2(n4545), .ZN(n4438) );
  OAI211_X1 U5072 ( .C1(n4440), .C2(n4541), .A(n4439), .B(n4438), .ZN(n4441)
         );
  AOI21_X1 U5073 ( .B1(n4442), .B2(n4531), .A(n4441), .ZN(n4608) );
  OAI22_X1 U5074 ( .A1(n4557), .A2(n4049), .B1(n4443), .B2(n4519), .ZN(n4444)
         );
  INV_X1 U5075 ( .A(n4444), .ZN(n4447) );
  NAND2_X1 U5076 ( .A1(n4461), .A2(n4445), .ZN(n4605) );
  NAND3_X1 U5077 ( .A1(n4606), .A2(n4817), .A3(n4605), .ZN(n4446) );
  OAI211_X1 U5078 ( .C1(n4608), .C2(n4813), .A(n4447), .B(n4446), .ZN(n4448)
         );
  INV_X1 U5079 ( .A(n4448), .ZN(n4449) );
  OAI21_X1 U5080 ( .B1(n4609), .B2(n4559), .A(n4449), .ZN(U3268) );
  XOR2_X1 U5081 ( .A(n4451), .B(n4450), .Z(n4611) );
  INV_X1 U5082 ( .A(n4611), .ZN(n4466) );
  XNOR2_X1 U5083 ( .A(n4452), .B(n4451), .ZN(n4458) );
  NOR2_X1 U5084 ( .A1(n4459), .A2(n4565), .ZN(n4453) );
  AOI21_X1 U5085 ( .B1(n4454), .B2(n4525), .A(n4453), .ZN(n4457) );
  NAND2_X1 U5086 ( .A1(n4455), .A2(n4545), .ZN(n4456) );
  OAI211_X1 U5087 ( .C1(n4458), .C2(n4547), .A(n4457), .B(n4456), .ZN(n4610)
         );
  OR2_X1 U5088 ( .A1(n4483), .A2(n4459), .ZN(n4460) );
  NAND2_X1 U5089 ( .A1(n4461), .A2(n4460), .ZN(n4669) );
  AOI22_X1 U5090 ( .A1(n4813), .A2(REG2_REG_21__SCAN_IN), .B1(n4462), .B2(
        n4826), .ZN(n4463) );
  OAI21_X1 U5091 ( .B1(n4669), .B2(n4555), .A(n4463), .ZN(n4464) );
  AOI21_X1 U5092 ( .B1(n4610), .B2(n4557), .A(n4464), .ZN(n4465) );
  OAI21_X1 U5093 ( .B1(n4466), .B2(n4559), .A(n4465), .ZN(U3269) );
  XOR2_X1 U5094 ( .A(n4470), .B(n4467), .Z(n4480) );
  NAND2_X1 U5095 ( .A1(n4469), .A2(n4468), .ZN(n4471) );
  XNOR2_X1 U5096 ( .A(n4471), .B(n4470), .ZN(n4477) );
  AOI22_X1 U5097 ( .A1(n4473), .A2(n4525), .B1(n4576), .B2(n4472), .ZN(n4474)
         );
  OAI21_X1 U5098 ( .B1(n4475), .B2(n4528), .A(n4474), .ZN(n4476) );
  AOI21_X1 U5099 ( .B1(n4477), .B2(n4531), .A(n4476), .ZN(n4478) );
  OAI21_X1 U5100 ( .B1(n4480), .B2(n4479), .A(n4478), .ZN(n4614) );
  INV_X1 U5101 ( .A(n4614), .ZN(n4488) );
  INV_X1 U5102 ( .A(n4480), .ZN(n4615) );
  NOR2_X1 U5103 ( .A1(n4504), .A2(n4481), .ZN(n4482) );
  OR2_X1 U5104 ( .A1(n4483), .A2(n4482), .ZN(n4673) );
  AOI22_X1 U5105 ( .A1(n4813), .A2(REG2_REG_20__SCAN_IN), .B1(n4484), .B2(
        n4826), .ZN(n4485) );
  OAI21_X1 U5106 ( .B1(n4673), .B2(n4555), .A(n4485), .ZN(n4486) );
  AOI21_X1 U5107 ( .B1(n4615), .B2(n4828), .A(n4486), .ZN(n4487) );
  OAI21_X1 U5108 ( .B1(n4488), .B2(n4813), .A(n4487), .ZN(U3270) );
  XNOR2_X1 U5109 ( .A(n4489), .B(n4496), .ZN(n4619) );
  INV_X1 U5110 ( .A(n4619), .ZN(n4512) );
  INV_X1 U5111 ( .A(n4490), .ZN(n4492) );
  OAI21_X1 U5112 ( .B1(n4540), .B2(n4492), .A(n4491), .ZN(n4523) );
  INV_X1 U5113 ( .A(n4493), .ZN(n4495) );
  OAI21_X1 U5114 ( .B1(n4523), .B2(n4495), .A(n4494), .ZN(n4497) );
  XNOR2_X1 U5115 ( .A(n4497), .B(n4496), .ZN(n4501) );
  NOR2_X1 U5116 ( .A1(n4542), .A2(n4528), .ZN(n4500) );
  OAI22_X1 U5117 ( .A1(n4498), .A2(n4541), .B1(n4565), .B2(n4506), .ZN(n4499)
         );
  AOI211_X1 U5118 ( .C1(n4501), .C2(n4531), .A(n4500), .B(n4499), .ZN(n4502)
         );
  INV_X1 U5119 ( .A(n4502), .ZN(n4618) );
  INV_X1 U5120 ( .A(n4503), .ZN(n4507) );
  INV_X1 U5121 ( .A(n4504), .ZN(n4505) );
  OAI21_X1 U5122 ( .B1(n4507), .B2(n4506), .A(n4505), .ZN(n4677) );
  AOI22_X1 U5123 ( .A1(n4813), .A2(REG2_REG_19__SCAN_IN), .B1(n4508), .B2(
        n4826), .ZN(n4509) );
  OAI21_X1 U5124 ( .B1(n4677), .B2(n4555), .A(n4509), .ZN(n4510) );
  AOI21_X1 U5125 ( .B1(n4618), .B2(n4557), .A(n4510), .ZN(n4511) );
  OAI21_X1 U5126 ( .B1(n4512), .B2(n4559), .A(n4511), .ZN(U3271) );
  OAI21_X1 U5127 ( .B1(n4513), .B2(n4515), .A(n4514), .ZN(n4516) );
  INV_X1 U5128 ( .A(n4516), .ZN(n4624) );
  XNOR2_X1 U5129 ( .A(n4552), .B(n4517), .ZN(n4518) );
  NAND2_X1 U5130 ( .A1(n4518), .A2(n4636), .ZN(n4622) );
  INV_X1 U5131 ( .A(n4622), .ZN(n4536) );
  INV_X1 U5132 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4521) );
  OAI22_X1 U5133 ( .A1(n4557), .A2(n4521), .B1(n4520), .B2(n4519), .ZN(n4534)
         );
  XNOR2_X1 U5134 ( .A(n4523), .B(n4522), .ZN(n4532) );
  AOI22_X1 U5135 ( .A1(n4526), .A2(n4525), .B1(n4524), .B2(n4576), .ZN(n4527)
         );
  OAI21_X1 U5136 ( .B1(n4529), .B2(n4528), .A(n4527), .ZN(n4530) );
  AOI21_X1 U5137 ( .B1(n4532), .B2(n4531), .A(n4530), .ZN(n4623) );
  NOR2_X1 U5138 ( .A1(n4623), .A2(n4813), .ZN(n4533) );
  AOI211_X1 U5139 ( .C1(n4536), .C2(n4535), .A(n4534), .B(n4533), .ZN(n4537)
         );
  OAI21_X1 U5140 ( .B1(n4624), .B2(n4559), .A(n4537), .ZN(U3272) );
  XNOR2_X1 U5141 ( .A(n4538), .B(n4539), .ZN(n4626) );
  INV_X1 U5142 ( .A(n4626), .ZN(n4560) );
  XNOR2_X1 U5143 ( .A(n4540), .B(n4539), .ZN(n4548) );
  OAI22_X1 U5144 ( .A1(n4542), .A2(n4541), .B1(n4565), .B2(n4549), .ZN(n4543)
         );
  AOI21_X1 U5145 ( .B1(n4545), .B2(n4544), .A(n4543), .ZN(n4546) );
  OAI21_X1 U5146 ( .B1(n4548), .B2(n4547), .A(n4546), .ZN(n4625) );
  OR2_X1 U5147 ( .A1(n4550), .A2(n4549), .ZN(n4551) );
  NAND2_X1 U5148 ( .A1(n4552), .A2(n4551), .ZN(n4683) );
  AOI22_X1 U5149 ( .A1(n4813), .A2(REG2_REG_17__SCAN_IN), .B1(n4553), .B2(
        n4826), .ZN(n4554) );
  OAI21_X1 U5150 ( .B1(n4683), .B2(n4555), .A(n4554), .ZN(n4556) );
  AOI21_X1 U5151 ( .B1(n4625), .B2(n4557), .A(n4556), .ZN(n4558) );
  OAI21_X1 U5152 ( .B1(n4560), .B2(n4559), .A(n4558), .ZN(U3273) );
  INV_X1 U5153 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4569) );
  NAND2_X1 U5154 ( .A1(n4570), .A2(n4561), .ZN(n4571) );
  XNOR2_X1 U5155 ( .A(n4571), .B(n4566), .ZN(n4703) );
  NAND2_X1 U5156 ( .A1(n4703), .A2(n4562), .ZN(n4568) );
  OR2_X1 U5157 ( .A1(n4564), .A2(n4563), .ZN(n4574) );
  OAI21_X1 U5158 ( .B1(n4566), .B2(n4565), .A(n4574), .ZN(n4702) );
  NAND2_X1 U5159 ( .A1(n4702), .A2(n4910), .ZN(n4567) );
  OAI211_X1 U5160 ( .C1(n4910), .C2(n4569), .A(n4568), .B(n4567), .ZN(U3549)
         );
  INV_X1 U5161 ( .A(n4570), .ZN(n4573) );
  INV_X1 U5162 ( .A(n4571), .ZN(n4572) );
  AOI21_X1 U5163 ( .B1(n4577), .B2(n4573), .A(n4572), .ZN(n4706) );
  INV_X1 U5164 ( .A(n4706), .ZN(n4646) );
  INV_X1 U5165 ( .A(n4574), .ZN(n4575) );
  AOI21_X1 U5166 ( .B1(n4577), .B2(n4576), .A(n4575), .ZN(n4708) );
  MUX2_X1 U5167 ( .A(n4578), .B(n4708), .S(n4910), .Z(n4579) );
  OAI21_X1 U5168 ( .B1(n4646), .B2(n4629), .A(n4579), .ZN(U3548) );
  NAND2_X1 U5169 ( .A1(n4580), .A2(n4891), .ZN(n4584) );
  NAND2_X1 U5170 ( .A1(n4584), .A2(n4583), .ZN(n4647) );
  MUX2_X1 U5171 ( .A(REG1_REG_29__SCAN_IN), .B(n4647), .S(n4910), .Z(U3547) );
  AOI21_X1 U5172 ( .B1(n4636), .B2(n4586), .A(n4585), .ZN(n4587) );
  OAI21_X1 U5173 ( .B1(n4588), .B2(n4638), .A(n4587), .ZN(n4648) );
  MUX2_X1 U5174 ( .A(REG1_REG_27__SCAN_IN), .B(n4648), .S(n4910), .Z(U3545) );
  AOI21_X1 U5175 ( .B1(n4590), .B2(n4891), .A(n4589), .ZN(n4649) );
  MUX2_X1 U5176 ( .A(n4591), .B(n4649), .S(n4910), .Z(n4592) );
  OAI21_X1 U5177 ( .B1(n4629), .B2(n4652), .A(n4592), .ZN(U3544) );
  INV_X1 U5178 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4595) );
  AOI21_X1 U5179 ( .B1(n4594), .B2(n4891), .A(n4593), .ZN(n4653) );
  MUX2_X1 U5180 ( .A(n4595), .B(n4653), .S(n4910), .Z(n4596) );
  OAI21_X1 U5181 ( .B1(n4629), .B2(n4656), .A(n4596), .ZN(U3543) );
  AOI21_X1 U5182 ( .B1(n4598), .B2(n4891), .A(n4597), .ZN(n4657) );
  MUX2_X1 U5183 ( .A(n4599), .B(n4657), .S(n4910), .Z(n4600) );
  OAI21_X1 U5184 ( .B1(n4629), .B2(n4660), .A(n4600), .ZN(U3542) );
  INV_X1 U5185 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4603) );
  AOI21_X1 U5186 ( .B1(n4602), .B2(n4891), .A(n4601), .ZN(n4661) );
  MUX2_X1 U5187 ( .A(n4603), .B(n4661), .S(n4910), .Z(n4604) );
  OAI21_X1 U5188 ( .B1(n4629), .B2(n4664), .A(n4604), .ZN(U3541) );
  NAND3_X1 U5189 ( .A1(n4606), .A2(n4636), .A3(n4605), .ZN(n4607) );
  OAI211_X1 U5190 ( .C1(n4609), .C2(n4638), .A(n4608), .B(n4607), .ZN(n4665)
         );
  MUX2_X1 U5191 ( .A(REG1_REG_22__SCAN_IN), .B(n4665), .S(n4910), .Z(U3540) );
  AOI21_X1 U5192 ( .B1(n4611), .B2(n4891), .A(n4610), .ZN(n4666) );
  MUX2_X1 U5193 ( .A(n4612), .B(n4666), .S(n4910), .Z(n4613) );
  OAI21_X1 U5194 ( .B1(n4629), .B2(n4669), .A(n4613), .ZN(U3539) );
  AOI21_X1 U5195 ( .B1(n4899), .B2(n4615), .A(n4614), .ZN(n4670) );
  MUX2_X1 U5196 ( .A(n4616), .B(n4670), .S(n4910), .Z(n4617) );
  OAI21_X1 U5197 ( .B1(n4629), .B2(n4673), .A(n4617), .ZN(U3538) );
  AOI21_X1 U5198 ( .B1(n4619), .B2(n4891), .A(n4618), .ZN(n4674) );
  MUX2_X1 U5199 ( .A(n4620), .B(n4674), .S(n4910), .Z(n4621) );
  OAI21_X1 U5200 ( .B1(n4629), .B2(n4677), .A(n4621), .ZN(U3537) );
  OAI211_X1 U5201 ( .C1(n4624), .C2(n4638), .A(n4623), .B(n4622), .ZN(n4678)
         );
  MUX2_X1 U5202 ( .A(REG1_REG_18__SCAN_IN), .B(n4678), .S(n4910), .Z(U3536) );
  AOI21_X1 U5203 ( .B1(n4626), .B2(n4891), .A(n4625), .ZN(n4679) );
  MUX2_X1 U5204 ( .A(n4627), .B(n4679), .S(n4910), .Z(n4628) );
  OAI21_X1 U5205 ( .B1(n4629), .B2(n4683), .A(n4628), .ZN(U3535) );
  AOI21_X1 U5206 ( .B1(n4636), .B2(n4631), .A(n4630), .ZN(n4632) );
  OAI21_X1 U5207 ( .B1(n4633), .B2(n4638), .A(n4632), .ZN(n4684) );
  MUX2_X1 U5208 ( .A(REG1_REG_16__SCAN_IN), .B(n4684), .S(n4910), .Z(U3534) );
  AOI21_X1 U5209 ( .B1(n4636), .B2(n4635), .A(n4634), .ZN(n4637) );
  OAI21_X1 U5210 ( .B1(n4639), .B2(n4638), .A(n4637), .ZN(n4685) );
  MUX2_X1 U5211 ( .A(REG1_REG_15__SCAN_IN), .B(n4685), .S(n4910), .Z(U3533) );
  NAND2_X1 U5212 ( .A1(n4703), .A2(n4640), .ZN(n4642) );
  NAND2_X1 U5213 ( .A1(n4702), .A2(n4902), .ZN(n4641) );
  OAI211_X1 U5214 ( .C1(n4902), .C2(n4643), .A(n4642), .B(n4641), .ZN(U3517)
         );
  INV_X1 U5215 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4644) );
  MUX2_X1 U5216 ( .A(n4644), .B(n4708), .S(n4902), .Z(n4645) );
  OAI21_X1 U5217 ( .B1(n4646), .B2(n4682), .A(n4645), .ZN(U3516) );
  MUX2_X1 U5218 ( .A(REG0_REG_29__SCAN_IN), .B(n4647), .S(n4902), .Z(U3515) );
  MUX2_X1 U5219 ( .A(REG0_REG_27__SCAN_IN), .B(n4648), .S(n4902), .Z(U3513) );
  MUX2_X1 U5220 ( .A(n4650), .B(n4649), .S(n4902), .Z(n4651) );
  OAI21_X1 U5221 ( .B1(n4652), .B2(n4682), .A(n4651), .ZN(U3512) );
  INV_X1 U5222 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4654) );
  MUX2_X1 U5223 ( .A(n4654), .B(n4653), .S(n4902), .Z(n4655) );
  OAI21_X1 U5224 ( .B1(n4656), .B2(n4682), .A(n4655), .ZN(U3511) );
  MUX2_X1 U5225 ( .A(n4658), .B(n4657), .S(n4902), .Z(n4659) );
  OAI21_X1 U5226 ( .B1(n4660), .B2(n4682), .A(n4659), .ZN(U3510) );
  INV_X1 U5227 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4662) );
  MUX2_X1 U5228 ( .A(n4662), .B(n4661), .S(n4902), .Z(n4663) );
  OAI21_X1 U5229 ( .B1(n4664), .B2(n4682), .A(n4663), .ZN(U3509) );
  MUX2_X1 U5230 ( .A(REG0_REG_22__SCAN_IN), .B(n4665), .S(n4902), .Z(U3508) );
  INV_X1 U5231 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4667) );
  MUX2_X1 U5232 ( .A(n4667), .B(n4666), .S(n4902), .Z(n4668) );
  OAI21_X1 U5233 ( .B1(n4669), .B2(n4682), .A(n4668), .ZN(U3507) );
  MUX2_X1 U5234 ( .A(n4671), .B(n4670), .S(n4902), .Z(n4672) );
  OAI21_X1 U5235 ( .B1(n4673), .B2(n4682), .A(n4672), .ZN(U3506) );
  INV_X1 U5236 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4675) );
  MUX2_X1 U5237 ( .A(n4675), .B(n4674), .S(n4902), .Z(n4676) );
  OAI21_X1 U5238 ( .B1(n4677), .B2(n4682), .A(n4676), .ZN(U3505) );
  MUX2_X1 U5239 ( .A(REG0_REG_18__SCAN_IN), .B(n4678), .S(n4902), .Z(U3503) );
  MUX2_X1 U5240 ( .A(n4680), .B(n4679), .S(n4902), .Z(n4681) );
  OAI21_X1 U5241 ( .B1(n4683), .B2(n4682), .A(n4681), .ZN(U3501) );
  MUX2_X1 U5242 ( .A(REG0_REG_16__SCAN_IN), .B(n4684), .S(n4902), .Z(U3499) );
  MUX2_X1 U5243 ( .A(REG0_REG_15__SCAN_IN), .B(n4685), .S(n4902), .Z(U3497) );
  MUX2_X1 U5244 ( .A(n4686), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U5245 ( .A(n4687), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5246 ( .A(DATAI_24_), .B(n2852), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U5247 ( .A(n4688), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U5248 ( .A(n4689), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U5249 ( .A(DATAI_20_), .B(n4690), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5250 ( .A(n4691), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U5251 ( .A(DATAI_8_), .B(n2252), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U5252 ( .A(n4693), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U5253 ( .A(n4694), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5254 ( .A(n4695), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5255 ( .A(DATAI_4_), .B(n4696), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5256 ( .A(n4697), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5257 ( .A(n4698), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5258 ( .A(n4699), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  AOI22_X1 U5259 ( .A1(STATE_REG_SCAN_IN), .A2(n4701), .B1(n4700), .B2(U3149), 
        .ZN(U3324) );
  AOI22_X1 U5260 ( .A1(n4703), .A2(n4817), .B1(n3190), .B2(n4702), .ZN(n4704)
         );
  OAI21_X1 U5261 ( .B1(n3190), .B2(n4705), .A(n4704), .ZN(U3260) );
  AOI22_X1 U5262 ( .A1(n4706), .A2(n4817), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4813), .ZN(n4707) );
  OAI21_X1 U5263 ( .B1(n4813), .B2(n4708), .A(n4707), .ZN(U3261) );
  AOI211_X1 U5264 ( .C1(n4711), .C2(n4710), .A(n4709), .B(n4797), .ZN(n4713)
         );
  AOI211_X1 U5265 ( .C1(n4775), .C2(ADDR_REG_9__SCAN_IN), .A(n4713), .B(n4712), 
        .ZN(n4718) );
  OAI211_X1 U5266 ( .C1(n4716), .C2(n4715), .A(n4809), .B(n4714), .ZN(n4717)
         );
  OAI211_X1 U5267 ( .C1(n4812), .C2(n4860), .A(n4718), .B(n4717), .ZN(U3249)
         );
  AOI211_X1 U5268 ( .C1(n2619), .C2(n4720), .A(n4719), .B(n4797), .ZN(n4723)
         );
  INV_X1 U5269 ( .A(n4721), .ZN(n4722) );
  AOI211_X1 U5270 ( .C1(n4775), .C2(ADDR_REG_10__SCAN_IN), .A(n4723), .B(n4722), .ZN(n4727) );
  OAI211_X1 U5271 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4725), .A(n4809), .B(n4724), .ZN(n4726) );
  OAI211_X1 U5272 ( .C1(n4812), .C2(n3468), .A(n4727), .B(n4726), .ZN(U3250)
         );
  AOI211_X1 U5273 ( .C1(n2193), .C2(n4729), .A(n4728), .B(n4797), .ZN(n4731)
         );
  AOI211_X1 U5274 ( .C1(n4775), .C2(ADDR_REG_11__SCAN_IN), .A(n4731), .B(n4730), .ZN(n4736) );
  OAI211_X1 U5275 ( .C1(n4734), .C2(n4733), .A(n4809), .B(n4732), .ZN(n4735)
         );
  OAI211_X1 U5276 ( .C1(n4812), .C2(n4737), .A(n4736), .B(n4735), .ZN(U3251)
         );
  AOI211_X1 U5277 ( .C1(n4740), .C2(n4739), .A(n4738), .B(n4797), .ZN(n4743)
         );
  INV_X1 U5278 ( .A(n4741), .ZN(n4742) );
  AOI211_X1 U5279 ( .C1(n4775), .C2(ADDR_REG_12__SCAN_IN), .A(n4743), .B(n4742), .ZN(n4747) );
  OAI211_X1 U5280 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4745), .A(n4809), .B(n4744), .ZN(n4746) );
  OAI211_X1 U5281 ( .C1(n4812), .C2(n4854), .A(n4747), .B(n4746), .ZN(U3252)
         );
  NAND2_X1 U5282 ( .A1(ADDR_REG_14__SCAN_IN), .A2(n4775), .ZN(n4761) );
  AOI211_X1 U5283 ( .C1(n4750), .C2(n4749), .A(n4748), .B(n4797), .ZN(n4756)
         );
  AOI211_X1 U5284 ( .C1(n4754), .C2(n4753), .A(n4752), .B(n4751), .ZN(n4755)
         );
  AOI211_X1 U5285 ( .C1(n4758), .C2(n4757), .A(n4756), .B(n4755), .ZN(n4760)
         );
  NAND3_X1 U5286 ( .A1(n4761), .A2(n4760), .A3(n4759), .ZN(U3254) );
  AOI211_X1 U5287 ( .C1(n4764), .C2(n4763), .A(n4762), .B(n4797), .ZN(n4765)
         );
  AOI211_X1 U5288 ( .C1(n4775), .C2(ADDR_REG_15__SCAN_IN), .A(n4766), .B(n4765), .ZN(n4772) );
  AOI21_X1 U5289 ( .B1(n4769), .B2(n4768), .A(n4767), .ZN(n4770) );
  NAND2_X1 U5290 ( .A1(n4809), .A2(n4770), .ZN(n4771) );
  OAI211_X1 U5291 ( .C1(n4812), .C2(n4852), .A(n4772), .B(n4771), .ZN(U3255)
         );
  INV_X1 U5292 ( .A(n4773), .ZN(n4774) );
  AOI21_X1 U5293 ( .B1(n4775), .B2(ADDR_REG_16__SCAN_IN), .A(n4774), .ZN(n4784) );
  OAI21_X1 U5294 ( .B1(n4778), .B2(n4777), .A(n4776), .ZN(n4782) );
  OAI21_X1 U5295 ( .B1(n4780), .B2(n3596), .A(n4779), .ZN(n4781) );
  AOI22_X1 U5296 ( .A1(n4794), .A2(n4782), .B1(n4809), .B2(n4781), .ZN(n4783)
         );
  OAI211_X1 U5297 ( .C1(n4850), .C2(n4812), .A(n4784), .B(n4783), .ZN(U3256)
         );
  AOI21_X1 U5298 ( .B1(n4775), .B2(ADDR_REG_17__SCAN_IN), .A(n4785), .ZN(n4796) );
  OAI21_X1 U5299 ( .B1(n4788), .B2(n4787), .A(n4786), .ZN(n4793) );
  OAI21_X1 U5300 ( .B1(n4791), .B2(n4790), .A(n4789), .ZN(n4792) );
  AOI22_X1 U5301 ( .A1(n4794), .A2(n4793), .B1(n4809), .B2(n4792), .ZN(n4795)
         );
  OAI211_X1 U5302 ( .C1(n4848), .C2(n4812), .A(n4796), .B(n4795), .ZN(U3257)
         );
  AOI21_X1 U5303 ( .B1(n4799), .B2(n4798), .A(n4797), .ZN(n4804) );
  NAND2_X1 U5304 ( .A1(n4775), .A2(ADDR_REG_18__SCAN_IN), .ZN(n4802) );
  INV_X1 U5305 ( .A(n4800), .ZN(n4801) );
  AOI21_X1 U5306 ( .B1(n4807), .B2(n4806), .A(n4805), .ZN(n4808) );
  NAND2_X1 U5307 ( .A1(n4809), .A2(n4808), .ZN(n4810) );
  OAI211_X1 U5308 ( .C1(n4812), .C2(n4846), .A(n4811), .B(n4810), .ZN(U3258)
         );
  AOI22_X1 U5309 ( .A1(REG2_REG_2__SCAN_IN), .A2(n4813), .B1(
        REG3_REG_2__SCAN_IN), .B2(n4826), .ZN(n4820) );
  INV_X1 U5310 ( .A(n4814), .ZN(n4818) );
  INV_X1 U5311 ( .A(n4815), .ZN(n4816) );
  AOI22_X1 U5312 ( .A1(n4818), .A2(n4828), .B1(n4817), .B2(n4816), .ZN(n4819)
         );
  OAI211_X1 U5313 ( .C1(n4813), .C2(n4821), .A(n4820), .B(n4819), .ZN(U3288)
         );
  INV_X1 U5314 ( .A(n4822), .ZN(n4824) );
  AOI21_X1 U5315 ( .B1(n4825), .B2(n4824), .A(n4823), .ZN(n4830) );
  AOI22_X1 U5316 ( .A1(n4828), .A2(n4827), .B1(REG3_REG_0__SCAN_IN), .B2(n4826), .ZN(n4829) );
  OAI221_X1 U5317 ( .B1(n4813), .B2(n4830), .C1(n3190), .C2(n3071), .A(n4829), 
        .ZN(U3290) );
  AND2_X1 U5318 ( .A1(D_REG_31__SCAN_IN), .A2(n4842), .ZN(U3291) );
  AND2_X1 U5319 ( .A1(D_REG_30__SCAN_IN), .A2(n4842), .ZN(U3292) );
  AND2_X1 U5320 ( .A1(D_REG_29__SCAN_IN), .A2(n4842), .ZN(U3293) );
  AND2_X1 U5321 ( .A1(D_REG_28__SCAN_IN), .A2(n4842), .ZN(U3294) );
  AND2_X1 U5322 ( .A1(D_REG_27__SCAN_IN), .A2(n4842), .ZN(U3295) );
  AND2_X1 U5323 ( .A1(D_REG_26__SCAN_IN), .A2(n4842), .ZN(U3296) );
  NOR2_X1 U5324 ( .A1(n4841), .A2(n4831), .ZN(U3297) );
  AND2_X1 U5325 ( .A1(D_REG_24__SCAN_IN), .A2(n4842), .ZN(U3298) );
  AND2_X1 U5326 ( .A1(D_REG_23__SCAN_IN), .A2(n4842), .ZN(U3299) );
  AND2_X1 U5327 ( .A1(D_REG_22__SCAN_IN), .A2(n4842), .ZN(U3300) );
  AND2_X1 U5328 ( .A1(D_REG_21__SCAN_IN), .A2(n4842), .ZN(U3301) );
  NOR2_X1 U5329 ( .A1(n4841), .A2(n4832), .ZN(U3302) );
  AND2_X1 U5330 ( .A1(D_REG_19__SCAN_IN), .A2(n4842), .ZN(U3303) );
  AND2_X1 U5331 ( .A1(D_REG_18__SCAN_IN), .A2(n4842), .ZN(U3304) );
  AND2_X1 U5332 ( .A1(D_REG_17__SCAN_IN), .A2(n4842), .ZN(U3305) );
  NOR2_X1 U5333 ( .A1(n4841), .A2(n4833), .ZN(U3306) );
  AND2_X1 U5334 ( .A1(D_REG_15__SCAN_IN), .A2(n4842), .ZN(U3307) );
  AND2_X1 U5335 ( .A1(D_REG_14__SCAN_IN), .A2(n4842), .ZN(U3308) );
  NOR2_X1 U5336 ( .A1(n4841), .A2(n4834), .ZN(U3309) );
  AND2_X1 U5337 ( .A1(D_REG_12__SCAN_IN), .A2(n4842), .ZN(U3310) );
  NOR2_X1 U5338 ( .A1(n4841), .A2(n4835), .ZN(U3311) );
  NOR2_X1 U5339 ( .A1(n4841), .A2(n4836), .ZN(U3312) );
  NOR2_X1 U5340 ( .A1(n4841), .A2(n4837), .ZN(U3313) );
  NOR2_X1 U5341 ( .A1(n4841), .A2(n4838), .ZN(U3314) );
  AND2_X1 U5342 ( .A1(D_REG_7__SCAN_IN), .A2(n4842), .ZN(U3315) );
  AND2_X1 U5343 ( .A1(D_REG_6__SCAN_IN), .A2(n4842), .ZN(U3316) );
  NOR2_X1 U5344 ( .A1(n4841), .A2(n4839), .ZN(U3317) );
  AND2_X1 U5345 ( .A1(D_REG_4__SCAN_IN), .A2(n4842), .ZN(U3318) );
  NOR2_X1 U5346 ( .A1(n4841), .A2(n4840), .ZN(U3319) );
  AND2_X1 U5347 ( .A1(D_REG_2__SCAN_IN), .A2(n4842), .ZN(U3320) );
  AOI21_X1 U5348 ( .B1(U3149), .B2(n4844), .A(n4843), .ZN(U3329) );
  INV_X1 U5349 ( .A(DATAI_18_), .ZN(n4845) );
  AOI22_X1 U5350 ( .A1(STATE_REG_SCAN_IN), .A2(n4846), .B1(n4845), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U5351 ( .A1(STATE_REG_SCAN_IN), .A2(n4848), .B1(n4847), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U5352 ( .A(DATAI_16_), .ZN(n4849) );
  AOI22_X1 U5353 ( .A1(STATE_REG_SCAN_IN), .A2(n4850), .B1(n4849), .B2(U3149), 
        .ZN(U3336) );
  AOI22_X1 U5354 ( .A1(STATE_REG_SCAN_IN), .A2(n4852), .B1(n4851), .B2(U3149), 
        .ZN(U3337) );
  AOI22_X1 U5355 ( .A1(STATE_REG_SCAN_IN), .A2(n2282), .B1(n4853), .B2(U3149), 
        .ZN(U3338) );
  AOI22_X1 U5356 ( .A1(STATE_REG_SCAN_IN), .A2(n4854), .B1(n2655), .B2(U3149), 
        .ZN(U3340) );
  OAI22_X1 U5357 ( .A1(U3149), .A2(n4855), .B1(DATAI_11_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4856) );
  INV_X1 U5358 ( .A(n4856), .ZN(U3341) );
  OAI22_X1 U5359 ( .A1(U3149), .A2(n4857), .B1(DATAI_10_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4858) );
  INV_X1 U5360 ( .A(n4858), .ZN(U3342) );
  INV_X1 U5361 ( .A(DATAI_9_), .ZN(n4859) );
  AOI22_X1 U5362 ( .A1(STATE_REG_SCAN_IN), .A2(n4860), .B1(n4859), .B2(U3149), 
        .ZN(U3343) );
  INV_X1 U5363 ( .A(DATAI_0_), .ZN(n4862) );
  AOI22_X1 U5364 ( .A1(STATE_REG_SCAN_IN), .A2(n2419), .B1(n4862), .B2(U3149), 
        .ZN(U3352) );
  INV_X1 U5365 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4863) );
  AOI22_X1 U5366 ( .A1(n4902), .A2(n4864), .B1(n4863), .B2(n4900), .ZN(U3467)
         );
  AOI22_X1 U5367 ( .A1(n4902), .A2(n4866), .B1(n4865), .B2(n4900), .ZN(U3469)
         );
  NOR2_X1 U5368 ( .A1(n4867), .A2(n4894), .ZN(n4868) );
  AOI21_X1 U5369 ( .B1(n4869), .B2(n4899), .A(n4868), .ZN(n4870) );
  AND2_X1 U5370 ( .A1(n4871), .A2(n4870), .ZN(n4903) );
  INV_X1 U5371 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4872) );
  AOI22_X1 U5372 ( .A1(n4902), .A2(n4903), .B1(n4872), .B2(n4900), .ZN(U3473)
         );
  INV_X1 U5373 ( .A(n4873), .ZN(n4875) );
  AOI211_X1 U5374 ( .C1(n4876), .C2(n4899), .A(n4875), .B(n4874), .ZN(n4904)
         );
  AOI22_X1 U5375 ( .A1(n4902), .A2(n4904), .B1(n4877), .B2(n4900), .ZN(U3475)
         );
  OAI21_X1 U5376 ( .B1(n4894), .B2(n4879), .A(n4878), .ZN(n4880) );
  AOI21_X1 U5377 ( .B1(n4881), .B2(n4891), .A(n4880), .ZN(n4905) );
  INV_X1 U5378 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4882) );
  AOI22_X1 U5379 ( .A1(n4902), .A2(n4905), .B1(n4882), .B2(n4900), .ZN(U3477)
         );
  NAND3_X1 U5380 ( .A1(n3340), .A2(n4883), .A3(n4891), .ZN(n4884) );
  AND3_X1 U5381 ( .A1(n4886), .A2(n4885), .A3(n4884), .ZN(n4906) );
  AOI22_X1 U5382 ( .A1(n4902), .A2(n4906), .B1(n4887), .B2(n4900), .ZN(U3481)
         );
  OAI21_X1 U5383 ( .B1(n4894), .B2(n4889), .A(n4888), .ZN(n4890) );
  AOI21_X1 U5384 ( .B1(n4892), .B2(n4891), .A(n4890), .ZN(n4907) );
  AOI22_X1 U5385 ( .A1(n4902), .A2(n4907), .B1(n4893), .B2(n4900), .ZN(U3485)
         );
  NOR2_X1 U5386 ( .A1(n4895), .A2(n4894), .ZN(n4897) );
  AOI211_X1 U5387 ( .C1(n4899), .C2(n4898), .A(n4897), .B(n4896), .ZN(n4909)
         );
  INV_X1 U5388 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4901) );
  AOI22_X1 U5389 ( .A1(n4902), .A2(n4909), .B1(n4901), .B2(n4900), .ZN(U3489)
         );
  AOI22_X1 U5390 ( .A1(n4910), .A2(n4903), .B1(n2498), .B2(n4908), .ZN(U3521)
         );
  AOI22_X1 U5391 ( .A1(n4910), .A2(n4904), .B1(n3065), .B2(n4908), .ZN(U3522)
         );
  AOI22_X1 U5392 ( .A1(n4910), .A2(n4905), .B1(n3068), .B2(n4908), .ZN(U3523)
         );
  AOI22_X1 U5393 ( .A1(n4910), .A2(n4906), .B1(n2573), .B2(n4908), .ZN(U3525)
         );
  AOI22_X1 U5394 ( .A1(n4910), .A2(n4907), .B1(n2599), .B2(n4908), .ZN(U3527)
         );
  AOI22_X1 U5395 ( .A1(n4910), .A2(n4909), .B1(n2639), .B2(n4908), .ZN(U3529)
         );
  CLKBUF_X1 U2405 ( .A(n2484), .Z(n2975) );
endmodule

