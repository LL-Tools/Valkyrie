

module b20_C_AntiSAT_k_256_2 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, ADD_1068_U4, ADD_1068_U55, 
        ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, 
        ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, 
        ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, 
        ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, 
        P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, 
        P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, 
        P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, 
        P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, 
        P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, 
        P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, 
        P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, 
        P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, 
        P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, 
        P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, 
        P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, 
        P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, 
        P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, 
        P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, 
        P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, 
        P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, 
        P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, 
        P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, 
        P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, 
        P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, 
        P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, 
        P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4491, n4492, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438;

  AND2_X1 U4997 ( .A1(n7844), .A2(n7843), .ZN(n8596) );
  INV_X2 U4999 ( .A(n7841), .ZN(n4814) );
  CLKBUF_X2 U5000 ( .A(n5599), .Z(n9477) );
  INV_X1 U5002 ( .A(n9621), .ZN(n5281) );
  INV_X1 U5003 ( .A(n7595), .ZN(n4617) );
  INV_X1 U5004 ( .A(n7893), .ZN(n7892) );
  OR2_X1 U5005 ( .A1(n7357), .A2(n7932), .ZN(n7471) );
  INV_X1 U5006 ( .A(n5716), .ZN(n8208) );
  INV_X1 U5007 ( .A(n7903), .ZN(n7865) );
  CLKBUF_X2 U5008 ( .A(n8097), .Z(n4495) );
  INV_X1 U5009 ( .A(n5702), .ZN(n8182) );
  AND2_X1 U5010 ( .A1(n7625), .A2(n7595), .ZN(n5707) );
  NAND2_X1 U5011 ( .A1(n5175), .A2(n5176), .ZN(n5589) );
  INV_X1 U5012 ( .A(n5911), .ZN(n6700) );
  INV_X1 U5013 ( .A(n5741), .ZN(n6339) );
  INV_X1 U5014 ( .A(n9325), .ZN(n5736) );
  AOI21_X1 U5015 ( .B1(n7398), .B2(n7397), .A(n4958), .ZN(n7401) );
  INV_X1 U5016 ( .A(n7977), .ZN(n6547) );
  NAND4_X2 U5017 ( .A1(n5300), .A2(n5298), .A3(n5299), .A4(n4616), .ZN(n5593)
         );
  OAI21_X2 U5018 ( .B1(n5133), .B2(n7250), .A(n5134), .ZN(n5761) );
  OAI21_X2 U5019 ( .B1(n6371), .B2(n6370), .A(n6369), .ZN(n6554) );
  NOR2_X2 U5020 ( .A1(n6265), .A2(n6266), .ZN(n6371) );
  XNOR2_X2 U5021 ( .A(n5777), .B(P2_IR_REG_20__SCAN_IN), .ZN(n7977) );
  OAI21_X1 U5022 ( .B1(n9987), .B2(n4561), .A(n4915), .ZN(n4611) );
  AND2_X1 U5023 ( .A1(n9319), .A2(n5706), .ZN(n5719) );
  BUF_X2 U5024 ( .A(n5708), .Z(n9476) );
  CLKBUF_X1 U5025 ( .A(n5786), .Z(n7973) );
  CLKBUF_X3 U5026 ( .A(n5895), .Z(n9473) );
  CLKBUF_X2 U5027 ( .A(n5707), .Z(n4491) );
  CLKBUF_X2 U5028 ( .A(n5707), .Z(n4492) );
  XNOR2_X1 U5029 ( .A(n5261), .B(n5260), .ZN(n9577) );
  AND2_X1 U5030 ( .A1(n9827), .A2(n9826), .ZN(n10048) );
  OAI21_X1 U5031 ( .B1(n4591), .B2(n9341), .A(n9340), .ZN(n9343) );
  NAND2_X1 U5032 ( .A1(n4602), .A2(n9838), .ZN(n9792) );
  NAND2_X1 U5033 ( .A1(n7891), .A2(n7890), .ZN(n4813) );
  NOR2_X1 U5034 ( .A1(n10040), .A2(n4839), .ZN(n10043) );
  MUX2_X1 U5035 ( .A(n7887), .B(n7886), .S(n7892), .Z(n7891) );
  NOR2_X1 U5036 ( .A1(n8163), .A2(n8161), .ZN(n4998) );
  INV_X1 U5037 ( .A(n4614), .ZN(n9920) );
  AOI21_X1 U5038 ( .B1(n8386), .B2(n8558), .A(n5003), .ZN(n8281) );
  NAND2_X1 U5039 ( .A1(n8606), .A2(n7964), .ZN(n8585) );
  OAI21_X1 U5040 ( .B1(n10000), .B2(n9977), .A(n9781), .ZN(n9952) );
  NAND2_X1 U5041 ( .A1(n9868), .A2(n9873), .ZN(n9867) );
  XNOR2_X1 U5042 ( .A(n4965), .B(n4509), .ZN(n8301) );
  INV_X1 U5043 ( .A(n4611), .ZN(n9974) );
  NAND2_X1 U5044 ( .A1(n9895), .A2(n4529), .ZN(n9828) );
  OR2_X1 U5045 ( .A1(n8642), .A2(n8415), .ZN(n8614) );
  NAND2_X1 U5046 ( .A1(n6790), .A2(n4517), .ZN(n6968) );
  AND2_X1 U5047 ( .A1(n7018), .A2(n4866), .ZN(n4865) );
  NOR2_X1 U5048 ( .A1(n4526), .A2(n4868), .ZN(n4867) );
  NAND2_X1 U5049 ( .A1(n7467), .A2(n7466), .ZN(n8331) );
  NAND2_X1 U5050 ( .A1(n4590), .A2(n4589), .ZN(n4586) );
  NOR2_X1 U5051 ( .A1(n7836), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n7859) );
  OR2_X1 U5052 ( .A1(n7826), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n7836) );
  NAND2_X1 U5053 ( .A1(n5634), .A2(n5633), .ZN(n4953) );
  INV_X2 U5054 ( .A(n10028), .ZN(n9986) );
  INV_X2 U5055 ( .A(n8139), .ZN(n8258) );
  NOR2_X1 U5056 ( .A1(n6470), .A2(n5911), .ZN(n6431) );
  AND2_X1 U5057 ( .A1(n7651), .A2(n7649), .ZN(n7916) );
  NAND2_X1 U5058 ( .A1(n4817), .A2(n5149), .ZN(n5194) );
  NOR2_X1 U5059 ( .A1(n5743), .A2(n6705), .ZN(n6802) );
  AND3_X1 U5060 ( .A1(n5711), .A2(n5710), .A3(n5709), .ZN(n6804) );
  NAND3_X1 U5061 ( .A1(n5297), .A2(n5296), .A3(n5295), .ZN(n5594) );
  AND2_X2 U5062 ( .A1(n6985), .A2(n5033), .ZN(P1_U3973) );
  INV_X1 U5063 ( .A(n5597), .ZN(n5743) );
  NAND2_X2 U5064 ( .A1(n7973), .A2(n7986), .ZN(n7893) );
  NAND4_X1 U5065 ( .A1(n5800), .A2(n5799), .A3(n5798), .A4(n5797), .ZN(n8430)
         );
  INV_X2 U5066 ( .A(n6564), .ZN(n7873) );
  OR2_X1 U5067 ( .A1(n5281), .A2(n5280), .ZN(n5520) );
  NAND4_X2 U5068 ( .A1(n5794), .A2(n5793), .A3(n5792), .A4(n5791), .ZN(n8429)
         );
  OAI211_X1 U5069 ( .C1(n5894), .C2(n7994), .A(n5700), .B(n5699), .ZN(n9325)
         );
  INV_X2 U5070 ( .A(n5894), .ZN(n9467) );
  OAI211_X1 U5071 ( .C1(n5894), .C2(n5715), .A(n5714), .B(n5713), .ZN(n5741)
         );
  NAND2_X1 U5072 ( .A1(n9531), .A2(n9577), .ZN(n6278) );
  XNOR2_X1 U5073 ( .A(n5047), .B(P2_IR_REG_25__SCAN_IN), .ZN(n7250) );
  OAI21_X1 U5074 ( .B1(n5589), .B2(n5279), .A(n5278), .ZN(n6705) );
  NOR2_X1 U5075 ( .A1(n7318), .A2(n7315), .ZN(n5032) );
  NAND2_X1 U5076 ( .A1(n5810), .A2(n5085), .ZN(n6564) );
  NAND2_X2 U5077 ( .A1(n5810), .A2(n7901), .ZN(n7874) );
  NAND2_X1 U5078 ( .A1(n5056), .A2(n5055), .ZN(n7395) );
  NAND2_X1 U5079 ( .A1(n5027), .A2(n5030), .ZN(n7318) );
  NAND2_X1 U5080 ( .A1(n5030), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5031) );
  AND2_X2 U5081 ( .A1(n5293), .A2(n7595), .ZN(n5599) );
  NAND2_X2 U5082 ( .A1(n5320), .A2(n5321), .ZN(n7288) );
  OR2_X1 U5083 ( .A1(n5054), .A2(n5053), .ZN(n5056) );
  AND2_X2 U5084 ( .A1(n7593), .A2(n5320), .ZN(n7903) );
  INV_X1 U5085 ( .A(n5320), .ZN(n9218) );
  MUX2_X1 U5086 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5290), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5292) );
  MUX2_X1 U5087 ( .A(n5077), .B(P2_IR_REG_31__SCAN_IN), .S(n5073), .Z(n5079)
         );
  XNOR2_X1 U5088 ( .A(n5288), .B(n5287), .ZN(n7625) );
  XNOR2_X1 U5089 ( .A(n5029), .B(n5022), .ZN(n7315) );
  MUX2_X1 U5090 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5170), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5171) );
  NAND2_X1 U5091 ( .A1(n5991), .A2(n5253), .ZN(n6062) );
  OR2_X1 U5092 ( .A1(n6119), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n5778) );
  NAND2_X1 U5093 ( .A1(n5252), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5991) );
  AND2_X1 U5094 ( .A1(n4609), .A2(n4631), .ZN(n5286) );
  NAND2_X2 U5095 ( .A1(n7901), .A2(P1_U3086), .ZN(n10173) );
  AND2_X1 U5096 ( .A1(n4504), .A2(n5167), .ZN(n4607) );
  AND3_X1 U5097 ( .A1(n5021), .A2(n4516), .A3(n5256), .ZN(n5168) );
  AND2_X1 U5098 ( .A1(n5166), .A2(n5165), .ZN(n5167) );
  AND2_X1 U5099 ( .A1(n4966), .A2(n5374), .ZN(n4969) );
  AND2_X1 U5100 ( .A1(n5006), .A2(n5150), .ZN(n5007) );
  NAND3_X1 U5101 ( .A1(n4711), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4955) );
  AND2_X1 U5102 ( .A1(n5008), .A2(n5236), .ZN(n4993) );
  AND2_X1 U5103 ( .A1(n5375), .A2(n4967), .ZN(n4966) );
  AND2_X1 U5104 ( .A1(n5016), .A2(n5005), .ZN(n5006) );
  AND3_X1 U5105 ( .A1(n4910), .A2(n4909), .A3(n4908), .ZN(n5021) );
  INV_X1 U5106 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n9084) );
  INV_X1 U5107 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n6421) );
  NOR2_X1 U5108 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n4909) );
  NOR2_X1 U5109 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n4910) );
  INV_X1 U5110 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5156) );
  INV_X1 U5111 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n4967) );
  INV_X1 U5112 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5236) );
  NOR2_X1 U5113 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5100) );
  NOR2_X1 U5114 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4569) );
  INV_X1 U5115 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4712) );
  INV_X1 U5116 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5004) );
  NOR2_X1 U5117 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n4912) );
  NOR2_X1 U5118 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n4911) );
  INV_X4 U5119 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  XNOR2_X2 U5120 ( .A(n5107), .B(SI_3_), .ZN(n5105) );
  XNOR2_X1 U5121 ( .A(n8254), .B(n8252), .ZN(n8386) );
  NOR2_X2 U5122 ( .A1(n5626), .A2(n5627), .ZN(n9322) );
  NOR2_X2 U5123 ( .A1(n6577), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6579) );
  XNOR2_X2 U5124 ( .A(n5164), .B(n5166), .ZN(n5175) );
  OAI21_X2 U5125 ( .B1(n7230), .B2(n7229), .A(n7228), .ZN(n7413) );
  NAND2_X2 U5126 ( .A1(n4570), .A2(n7019), .ZN(n7230) );
  AND2_X4 U5127 ( .A1(n5293), .A2(n4617), .ZN(n5720) );
  NAND2_X4 U5128 ( .A1(n9218), .A2(n5321), .ZN(n6581) );
  NOR2_X2 U5129 ( .A1(n7286), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7359) );
  OR2_X2 U5130 ( .A1(n7266), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7286) );
  OAI22_X4 U5131 ( .A1(n8575), .A2(n8576), .B1(n8566), .B2(n8582), .ZN(n8537)
         );
  AOI21_X2 U5132 ( .B1(n8585), .B2(n7966), .A(n7965), .ZN(n8575) );
  NOR2_X4 U5133 ( .A1(n4851), .A2(n5122), .ZN(n5538) );
  NAND2_X2 U5134 ( .A1(n4852), .A2(n5004), .ZN(n5122) );
  XOR2_X2 U5135 ( .A(n8562), .B(n8537), .Z(n8733) );
  XNOR2_X2 U5136 ( .A(n5031), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5247) );
  INV_X1 U5137 ( .A(n5589), .ZN(n4494) );
  AND2_X4 U5138 ( .A1(n5515), .A2(n5519), .ZN(n5521) );
  NAND2_X2 U5139 ( .A1(n5032), .A2(n5247), .ZN(n5519) );
  NAND3_X1 U5140 ( .A1(n5520), .A2(n5519), .A3(n6278), .ZN(n8097) );
  INV_X1 U5141 ( .A(n7735), .ZN(n4779) );
  AND2_X1 U5142 ( .A1(n7184), .A2(n7177), .ZN(n7248) );
  OAI21_X2 U5143 ( .B1(n5480), .B2(n4744), .A(n4742), .ZN(n5634) );
  INV_X1 U5144 ( .A(n4745), .ZN(n4744) );
  AOI21_X1 U5145 ( .B1(n4743), .B2(n4745), .A(n4535), .ZN(n4742) );
  NOR2_X1 U5146 ( .A1(n5546), .A2(n4746), .ZN(n4745) );
  OAI22_X1 U5147 ( .A1(n8316), .A2(n8317), .B1(n8251), .B2(n8639), .ZN(n8254)
         );
  NAND2_X1 U5148 ( .A1(n5074), .A2(n5073), .ZN(n5078) );
  NAND2_X1 U5149 ( .A1(n5520), .A2(n5517), .ZN(n5518) );
  NAND2_X1 U5150 ( .A1(n4593), .A2(n4592), .ZN(n9778) );
  AOI21_X1 U5151 ( .B1(n4595), .B2(n4597), .A(n4531), .ZN(n4592) );
  NAND2_X1 U5152 ( .A1(n6837), .A2(n4595), .ZN(n4593) );
  NAND2_X1 U5153 ( .A1(n7702), .A2(n7893), .ZN(n4794) );
  NOR2_X1 U5154 ( .A1(n4778), .A2(n4511), .ZN(n4777) );
  NAND2_X1 U5155 ( .A1(n4770), .A2(n7734), .ZN(n4769) );
  NAND2_X1 U5156 ( .A1(n4779), .A2(n4771), .ZN(n4770) );
  OAI21_X1 U5157 ( .B1(n9551), .B2(n9395), .A(n4643), .ZN(n4640) );
  NAND2_X1 U5158 ( .A1(n4638), .A2(n9471), .ZN(n4637) );
  NAND2_X1 U5159 ( .A1(n4542), .A2(n9404), .ZN(n4638) );
  NAND2_X1 U5160 ( .A1(n4732), .A2(n6606), .ZN(n6604) );
  NAND2_X1 U5161 ( .A1(n4733), .A2(n6905), .ZN(n4732) );
  INV_X1 U5162 ( .A(n7921), .ZN(n4733) );
  AND2_X1 U5163 ( .A1(n7311), .A2(n7248), .ZN(n7186) );
  NOR2_X1 U5164 ( .A1(n5216), .A2(n4754), .ZN(n4753) );
  INV_X1 U5165 ( .A(n5196), .ZN(n4754) );
  INV_X1 U5166 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5613) );
  INV_X1 U5167 ( .A(n7593), .ZN(n5321) );
  OR2_X1 U5168 ( .A1(n8427), .A2(n10306), .ZN(n7674) );
  NOR2_X1 U5169 ( .A1(n4522), .A2(n4731), .ZN(n4729) );
  OR2_X1 U5170 ( .A1(n8393), .A2(n8329), .ZN(n7724) );
  OAI21_X2 U5171 ( .B1(n5778), .B2(P2_IR_REG_19__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5777) );
  OR2_X1 U5172 ( .A1(n5974), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5988) );
  NAND2_X1 U5173 ( .A1(n5374), .A2(n5375), .ZN(n5129) );
  OR2_X1 U5174 ( .A1(n8008), .A2(n8007), .ZN(n4882) );
  NOR2_X1 U5175 ( .A1(n9281), .A2(n4906), .ZN(n4905) );
  INV_X1 U5176 ( .A(n8021), .ZN(n4906) );
  AND2_X1 U5177 ( .A1(n4663), .A2(n4532), .ZN(n4662) );
  AND2_X1 U5178 ( .A1(n9622), .A2(n9597), .ZN(n4663) );
  NAND2_X1 U5179 ( .A1(n9867), .A2(n4524), .ZN(n9837) );
  AOI21_X1 U5180 ( .B1(n4923), .B2(n4925), .A(n4534), .ZN(n4922) );
  NAND2_X1 U5181 ( .A1(n10071), .A2(n9891), .ZN(n4933) );
  OR2_X1 U5182 ( .A1(n10071), .A2(n9924), .ZN(n9486) );
  NOR2_X1 U5183 ( .A1(n9944), .A2(n9784), .ZN(n4615) );
  INV_X1 U5184 ( .A(n4596), .ZN(n4595) );
  OAI21_X1 U5185 ( .B1(n4598), .B2(n4597), .A(n7209), .ZN(n4596) );
  OR2_X1 U5186 ( .A1(n9418), .A2(n9629), .ZN(n7209) );
  AND2_X1 U5187 ( .A1(n7196), .A2(n7194), .ZN(n7206) );
  INV_X1 U5188 ( .A(n5233), .ZN(n5012) );
  INV_X1 U5189 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5010) );
  INV_X1 U5190 ( .A(n4947), .ZN(n4946) );
  OAI21_X1 U5191 ( .B1(n4950), .B2(n4948), .A(n6292), .ZN(n4947) );
  NAND2_X1 U5192 ( .A1(n5231), .A2(n4515), .ZN(n5480) );
  NAND2_X1 U5193 ( .A1(n6099), .A2(n4978), .ZN(n6232) );
  NOR2_X1 U5194 ( .A1(n6102), .A2(n4979), .ZN(n4978) );
  INV_X1 U5195 ( .A(n6098), .ZN(n4979) );
  NAND2_X1 U5196 ( .A1(n7602), .A2(n4974), .ZN(n4972) );
  OR2_X1 U5197 ( .A1(n7601), .A2(n8421), .ZN(n4974) );
  OR2_X1 U5198 ( .A1(n7865), .A2(n5823), .ZN(n5827) );
  XNOR2_X1 U5199 ( .A(n8473), .B(n8477), .ZN(n8454) );
  AND2_X1 U5200 ( .A1(n7707), .A2(n7708), .ZN(n7928) );
  OR2_X1 U5201 ( .A1(n8772), .A2(n8341), .ZN(n8697) );
  OR2_X1 U5202 ( .A1(n7973), .A2(n7986), .ZN(n10352) );
  NAND2_X1 U5203 ( .A1(n7250), .A2(n5057), .ZN(n5834) );
  NOR2_X1 U5204 ( .A1(n7208), .A2(n7395), .ZN(n5057) );
  NAND2_X1 U5205 ( .A1(n9214), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5313) );
  INV_X1 U5206 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4980) );
  INV_X1 U5207 ( .A(n5074), .ZN(n5076) );
  AOI21_X1 U5208 ( .B1(n8166), .B2(n8162), .A(n4890), .ZN(n4889) );
  INV_X1 U5209 ( .A(n9263), .ZN(n4890) );
  AOI22_X1 U5210 ( .A1(n4648), .A2(n4645), .B1(n9458), .B2(n4643), .ZN(n9466)
         );
  AOI21_X1 U5211 ( .B1(n4662), .B2(n9596), .A(n4656), .ZN(n4655) );
  OR2_X1 U5212 ( .A1(n4657), .A2(n9574), .ZN(n4656) );
  AND2_X1 U5213 ( .A1(n4659), .A2(n4661), .ZN(n4657) );
  INV_X1 U5214 ( .A(n4491), .ZN(n8175) );
  AND2_X1 U5215 ( .A1(n7625), .A2(n4617), .ZN(n5708) );
  AND2_X1 U5216 ( .A1(n9720), .A2(n9719), .ZN(n9717) );
  AND2_X1 U5217 ( .A1(n10111), .A2(n9775), .ZN(n9776) );
  OR2_X1 U5218 ( .A1(n7031), .A2(n9633), .ZN(n6680) );
  OR2_X1 U5219 ( .A1(n7002), .A2(n9635), .ZN(n6447) );
  INV_X1 U5220 ( .A(n4605), .ZN(n4604) );
  INV_X1 U5221 ( .A(n6192), .ZN(n4606) );
  NAND2_X1 U5222 ( .A1(n9602), .A2(n9652), .ZN(n10011) );
  NAND2_X1 U5223 ( .A1(n9475), .A2(n9474), .ZN(n9766) );
  XNOR2_X1 U5224 ( .A(n7249), .B(n7248), .ZN(n8167) );
  AND2_X2 U5225 ( .A1(n4956), .A2(n4955), .ZN(n5085) );
  AND2_X1 U5226 ( .A1(n8248), .A2(n8415), .ZN(n8249) );
  OR2_X2 U5227 ( .A1(n6040), .A2(n6039), .ZN(n6099) );
  NAND2_X1 U5228 ( .A1(n9312), .A2(n8098), .ZN(n4580) );
  OAI21_X1 U5229 ( .B1(n9312), .B2(n8098), .A(n9309), .ZN(n8099) );
  AOI21_X1 U5230 ( .B1(n7669), .B2(n7668), .A(n7917), .ZN(n7675) );
  AOI21_X1 U5231 ( .B1(n7709), .B2(n7708), .A(n7893), .ZN(n4792) );
  NAND2_X1 U5232 ( .A1(n4680), .A2(n4688), .ZN(n4675) );
  NAND2_X1 U5233 ( .A1(n9378), .A2(n4682), .ZN(n4681) );
  OAI21_X1 U5234 ( .B1(n9376), .B2(n4678), .A(n4676), .ZN(n4690) );
  INV_X1 U5235 ( .A(n4679), .ZN(n4678) );
  AOI21_X1 U5236 ( .B1(n4686), .B2(n4679), .A(n4677), .ZN(n4676) );
  AND2_X1 U5237 ( .A1(n4683), .A2(n9381), .ZN(n4679) );
  NAND2_X1 U5238 ( .A1(n7281), .A2(n4797), .ZN(n4796) );
  INV_X1 U5239 ( .A(n7713), .ZN(n4797) );
  AND2_X1 U5240 ( .A1(n4792), .A2(n4793), .ZN(n4790) );
  INV_X1 U5241 ( .A(n7708), .ZN(n4793) );
  AOI21_X1 U5242 ( .B1(n7704), .B2(n4785), .A(n4513), .ZN(n4791) );
  AND2_X1 U5243 ( .A1(n4795), .A2(n4794), .ZN(n4785) );
  NAND2_X1 U5244 ( .A1(n7703), .A2(n7893), .ZN(n4795) );
  OAI21_X1 U5245 ( .B1(n7705), .B2(n4787), .A(n4781), .ZN(n4786) );
  OAI21_X1 U5246 ( .B1(n4769), .B2(n4773), .A(n7747), .ZN(n4766) );
  AND2_X1 U5247 ( .A1(n4779), .A2(n4774), .ZN(n4773) );
  INV_X1 U5248 ( .A(n4769), .ZN(n4768) );
  OAI22_X1 U5249 ( .A1(n4637), .A2(n4639), .B1(n4640), .B2(n4641), .ZN(n4636)
         );
  AND2_X1 U5250 ( .A1(n9404), .A2(n4644), .ZN(n4639) );
  NOR2_X1 U5251 ( .A1(n9395), .A2(n4642), .ZN(n4641) );
  NAND2_X1 U5252 ( .A1(n4668), .A2(n9520), .ZN(n4667) );
  NAND2_X1 U5253 ( .A1(n4670), .A2(n4669), .ZN(n4668) );
  NAND2_X1 U5254 ( .A1(n9521), .A2(n9471), .ZN(n4669) );
  NAND2_X1 U5255 ( .A1(n4673), .A2(n4671), .ZN(n4670) );
  INV_X1 U5256 ( .A(n4666), .ZN(n4665) );
  OAI21_X1 U5257 ( .B1(n9471), .B2(n9588), .A(n4823), .ZN(n4666) );
  OAI21_X1 U5258 ( .B1(n7822), .B2(n8621), .A(n7821), .ZN(n4800) );
  NAND2_X1 U5259 ( .A1(n8778), .A2(n7969), .ZN(n4763) );
  AND2_X1 U5260 ( .A1(n6602), .A2(n6604), .ZN(n6603) );
  NAND2_X1 U5261 ( .A1(n4735), .A2(n4734), .ZN(n7357) );
  AND2_X1 U5262 ( .A1(n7351), .A2(n7352), .ZN(n4734) );
  NAND2_X1 U5263 ( .A1(n7349), .A2(n7348), .ZN(n4735) );
  INV_X1 U5264 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5041) );
  AOI21_X1 U5265 ( .B1(n9449), .B2(n9448), .A(n9447), .ZN(n9454) );
  AND2_X1 U5266 ( .A1(n10155), .A2(n4859), .ZN(n4858) );
  OR2_X1 U5267 ( .A1(n7179), .A2(n7244), .ZN(n7185) );
  INV_X1 U5268 ( .A(n5977), .ZN(n5011) );
  INV_X1 U5269 ( .A(SI_12_), .ZN(n9082) );
  AND2_X1 U5270 ( .A1(n8367), .A2(n4963), .ZN(n4962) );
  NAND2_X1 U5271 ( .A1(n8244), .A2(n8243), .ZN(n4963) );
  AND2_X1 U5272 ( .A1(n7120), .A2(n6967), .ZN(n4987) );
  INV_X1 U5273 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5067) );
  INV_X1 U5274 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5040) );
  INV_X1 U5275 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5038) );
  NAND2_X1 U5276 ( .A1(n5389), .A2(n5500), .ZN(n5570) );
  NAND2_X1 U5277 ( .A1(n6137), .A2(n4708), .ZN(n6138) );
  OR2_X1 U5278 ( .A1(n6570), .A2(n6013), .ZN(n4708) );
  NAND2_X1 U5279 ( .A1(n6393), .A2(n4709), .ZN(n6527) );
  NAND2_X1 U5280 ( .A1(n6145), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4709) );
  NAND2_X1 U5281 ( .A1(n6865), .A2(n4706), .ZN(n6943) );
  NAND2_X1 U5282 ( .A1(n6534), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4706) );
  NAND2_X1 U5283 ( .A1(n8456), .A2(n4566), .ZN(n8494) );
  AOI21_X1 U5284 ( .B1(n7934), .B2(n4727), .A(n4726), .ZN(n4725) );
  INV_X1 U5285 ( .A(n7469), .ZN(n4727) );
  INV_X1 U5286 ( .A(n7551), .ZN(n4726) );
  OR2_X1 U5287 ( .A1(n7977), .A2(n8523), .ZN(n5866) );
  INV_X1 U5288 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n4804) );
  OR2_X1 U5289 ( .A1(n5687), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n5688) );
  INV_X1 U5290 ( .A(n6991), .ZN(n4869) );
  AND2_X1 U5291 ( .A1(n8039), .A2(n9280), .ZN(n4904) );
  NAND2_X1 U5292 ( .A1(n8060), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n8075) );
  NOR2_X1 U5293 ( .A1(n9977), .A2(n10099), .ZN(n4859) );
  INV_X1 U5294 ( .A(n9582), .ZN(n4835) );
  INV_X1 U5295 ( .A(n4834), .ZN(n4833) );
  OAI21_X1 U5296 ( .B1(n9580), .B2(n4835), .A(n9583), .ZN(n4834) );
  NOR2_X1 U5297 ( .A1(n9488), .A2(n4848), .ZN(n4847) );
  OR2_X1 U5298 ( .A1(n6661), .A2(n6660), .ZN(n6669) );
  OR2_X1 U5299 ( .A1(n6214), .A2(n6213), .ZN(n6300) );
  OR2_X1 U5300 ( .A1(n7002), .A2(n7113), .ZN(n6642) );
  INV_X1 U5301 ( .A(n9814), .ZN(n10042) );
  NAND2_X1 U5302 ( .A1(n4862), .A2(n4861), .ZN(n6855) );
  NAND2_X1 U5303 ( .A1(n5247), .A2(n5249), .ZN(n5273) );
  XNOR2_X1 U5304 ( .A(n7615), .B(n7616), .ZN(n7613) );
  NAND2_X1 U5305 ( .A1(n7197), .A2(n7196), .ZN(n7382) );
  AND2_X1 U5306 ( .A1(n7204), .A2(n7206), .ZN(n7195) );
  NAND2_X1 U5307 ( .A1(n6542), .A2(n6541), .ZN(n6716) );
  OR2_X1 U5308 ( .A1(n6540), .A2(n6539), .ZN(n6542) );
  AND2_X1 U5309 ( .A1(n4951), .A2(n6058), .ZN(n4950) );
  NAND2_X1 U5310 ( .A1(n5982), .A2(n5981), .ZN(n4951) );
  NAND2_X1 U5311 ( .A1(n5966), .A2(n5965), .ZN(n5983) );
  INV_X1 U5312 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5017) );
  NAND2_X1 U5313 ( .A1(n4749), .A2(n4748), .ZN(n5231) );
  INV_X1 U5314 ( .A(n4753), .ZN(n4752) );
  AOI21_X1 U5315 ( .B1(n5192), .B2(n4753), .A(n4751), .ZN(n4750) );
  INV_X1 U5316 ( .A(n5215), .ZN(n4751) );
  NAND2_X1 U5317 ( .A1(n5141), .A2(n5140), .ZN(n5147) );
  OAI21_X1 U5318 ( .B1(n5085), .B2(n5083), .A(n5082), .ZN(n5092) );
  INV_X1 U5319 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5083) );
  INV_X2 U5320 ( .A(n5085), .ZN(n5110) );
  OR2_X1 U5321 ( .A1(n8138), .A2(n4985), .ZN(n4982) );
  NOR2_X1 U5322 ( .A1(n8132), .A2(n4986), .ZN(n4985) );
  AND2_X1 U5323 ( .A1(n5882), .A2(n5886), .ZN(n5838) );
  AND2_X1 U5324 ( .A1(n7868), .A2(n7867), .ZN(n8566) );
  NAND2_X1 U5325 ( .A1(n4696), .A2(n4695), .ZN(n5502) );
  NAND2_X1 U5326 ( .A1(n7993), .A2(n4697), .ZN(n4695) );
  OR2_X1 U5327 ( .A1(n7993), .A2(n4697), .ZN(n4696) );
  NAND2_X1 U5328 ( .A1(n6007), .A2(n6008), .ZN(n6137) );
  NAND2_X1 U5329 ( .A1(n6146), .A2(n4692), .ZN(n6147) );
  OR2_X1 U5330 ( .A1(n6570), .A2(n6012), .ZN(n4692) );
  NAND2_X1 U5331 ( .A1(n6140), .A2(n6141), .ZN(n6393) );
  XNOR2_X1 U5332 ( .A(n6527), .B(n6730), .ZN(n6394) );
  NAND2_X1 U5333 ( .A1(n6531), .A2(n6532), .ZN(n6865) );
  XNOR2_X1 U5334 ( .A(n6943), .B(n7253), .ZN(n6866) );
  NAND2_X1 U5335 ( .A1(n8453), .A2(n4565), .ZN(n8473) );
  NAND2_X1 U5336 ( .A1(n8454), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8474) );
  NAND2_X1 U5337 ( .A1(n7882), .A2(n7881), .ZN(n8562) );
  AND4_X1 U5338 ( .A1(n6585), .A2(n6584), .A3(n6583), .A4(n6582), .ZN(n6969)
         );
  OR2_X1 U5339 ( .A1(n7841), .A2(n6576), .ZN(n6584) );
  AND2_X1 U5340 ( .A1(n5881), .A2(n5880), .ZN(n6172) );
  NAND2_X1 U5341 ( .A1(n9163), .A2(n8560), .ZN(n4937) );
  AND2_X1 U5342 ( .A1(n8630), .A2(n8555), .ZN(n8619) );
  AOI21_X1 U5343 ( .B1(n8668), .B2(n4703), .A(n7785), .ZN(n4702) );
  INV_X1 U5344 ( .A(n7953), .ZN(n4703) );
  OR2_X1 U5345 ( .A1(n7954), .A2(n8648), .ZN(n4701) );
  AND2_X1 U5346 ( .A1(n4540), .A2(n7956), .ZN(n8652) );
  AND2_X1 U5347 ( .A1(n7953), .A2(n7912), .ZN(n8678) );
  OR2_X1 U5348 ( .A1(n8718), .A2(n7947), .ZN(n8716) );
  NAND2_X1 U5349 ( .A1(n7548), .A2(n7547), .ZN(n7946) );
  AND4_X1 U5350 ( .A1(n7479), .A2(n7478), .A3(n7477), .A4(n7476), .ZN(n8721)
         );
  OR2_X1 U5351 ( .A1(n5872), .A2(n7893), .ZN(n10192) );
  INV_X1 U5352 ( .A(n8703), .ZN(n10194) );
  INV_X1 U5353 ( .A(n4724), .ZN(n7552) );
  AOI21_X1 U5354 ( .B1(n7471), .B2(n7469), .A(n7470), .ZN(n4724) );
  NAND2_X1 U5355 ( .A1(n4700), .A2(n4698), .ZN(n7464) );
  AOI21_X1 U5356 ( .B1(n7370), .B2(n4499), .A(n4699), .ZN(n4698) );
  NAND2_X1 U5357 ( .A1(n5870), .A2(n5869), .ZN(n8706) );
  INV_X1 U5358 ( .A(n10192), .ZN(n8701) );
  OR2_X1 U5359 ( .A1(n7272), .A2(n4499), .ZN(n7371) );
  INV_X1 U5360 ( .A(n8706), .ZN(n10296) );
  INV_X1 U5361 ( .A(n7208), .ZN(n5134) );
  INV_X1 U5362 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5316) );
  AND2_X1 U5363 ( .A1(n5073), .A2(n5312), .ZN(n4816) );
  XNOR2_X1 U5364 ( .A(n5075), .B(n5312), .ZN(n5820) );
  NAND2_X1 U5365 ( .A1(n5078), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5075) );
  NOR3_X1 U5366 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n5048) );
  AND2_X1 U5367 ( .A1(n5058), .A2(n5046), .ZN(n5054) );
  OR2_X1 U5368 ( .A1(n5314), .A2(n5059), .ZN(n5046) );
  INV_X1 U5369 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5053) );
  NAND2_X1 U5370 ( .A1(n5054), .A2(n5053), .ZN(n5055) );
  AND2_X1 U5371 ( .A1(n5130), .A2(n5184), .ZN(n6035) );
  INV_X1 U5372 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4693) );
  INV_X1 U5373 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5375) );
  INV_X1 U5374 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5019) );
  AOI21_X1 U5375 ( .B1(n4878), .B2(n4876), .A(n4558), .ZN(n4875) );
  INV_X1 U5376 ( .A(n4880), .ZN(n4876) );
  NAND2_X1 U5377 ( .A1(n4880), .A2(n4884), .ZN(n4874) );
  NAND2_X1 U5378 ( .A1(n8230), .A2(n8215), .ZN(n4897) );
  INV_X1 U5379 ( .A(n6261), .ZN(n4900) );
  NAND2_X1 U5380 ( .A1(n6264), .A2(n6263), .ZN(n6363) );
  NAND2_X1 U5381 ( .A1(n4586), .A2(n4588), .ZN(n6264) );
  INV_X1 U5382 ( .A(n4583), .ZN(n4582) );
  OAI21_X1 U5383 ( .B1(n4584), .B2(n4905), .A(n8040), .ZN(n4583) );
  NAND2_X1 U5384 ( .A1(n4885), .A2(n4889), .ZN(n9339) );
  OR2_X1 U5385 ( .A1(n4662), .A2(n4659), .ZN(n4658) );
  NOR2_X1 U5386 ( .A1(n4658), .A2(n9615), .ZN(n4653) );
  NOR2_X1 U5387 ( .A1(n9614), .A2(n4643), .ZN(n4652) );
  NAND2_X1 U5388 ( .A1(n4655), .A2(n5280), .ZN(n4654) );
  NOR2_X1 U5389 ( .A1(n4629), .A2(n7595), .ZN(n4991) );
  NAND2_X1 U5390 ( .A1(n7625), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4629) );
  NOR2_X1 U5391 ( .A1(n9717), .A2(n4564), .ZN(n7501) );
  INV_X1 U5392 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5081) );
  AND4_X1 U5393 ( .A1(n8207), .A2(n8206), .A3(n8205), .A4(n8204), .ZN(n9859)
         );
  NAND2_X1 U5394 ( .A1(n4924), .A2(n4496), .ZN(n4923) );
  INV_X1 U5395 ( .A(n4927), .ZN(n4924) );
  AOI21_X1 U5396 ( .B1(n4930), .B2(n4928), .A(n4502), .ZN(n4927) );
  AND2_X1 U5397 ( .A1(n10145), .A2(n9904), .ZN(n9895) );
  NOR2_X2 U5398 ( .A1(n10071), .A2(n9925), .ZN(n9904) );
  NOR2_X1 U5399 ( .A1(n10079), .A2(n9914), .ZN(n4934) );
  AND2_X1 U5400 ( .A1(n8002), .A2(n8001), .ZN(n9924) );
  NAND2_X1 U5401 ( .A1(n9588), .A2(n4827), .ZN(n4826) );
  INV_X1 U5402 ( .A(n9587), .ZN(n4827) );
  AND2_X1 U5403 ( .A1(n9962), .A2(n9972), .ZN(n9782) );
  NOR2_X1 U5404 ( .A1(n7213), .A2(n8833), .ZN(n8046) );
  NAND2_X1 U5405 ( .A1(n10099), .A2(n9971), .ZN(n4915) );
  AND4_X1 U5406 ( .A1(n7095), .A2(n7094), .A3(n7093), .A4(n7092), .ZN(n10012)
         );
  NOR2_X1 U5407 ( .A1(n4917), .A2(n4599), .ZN(n4598) );
  INV_X1 U5408 ( .A(n6836), .ZN(n4599) );
  NAND2_X1 U5409 ( .A1(n4921), .A2(n7073), .ZN(n4917) );
  INV_X1 U5410 ( .A(n4919), .ZN(n4918) );
  OAI21_X1 U5411 ( .B1(n9502), .B2(n4920), .A(n7078), .ZN(n4919) );
  NAND2_X1 U5412 ( .A1(n7074), .A2(n7073), .ZN(n7333) );
  NAND2_X1 U5413 ( .A1(n6843), .A2(n6844), .ZN(n7087) );
  OR2_X1 U5414 ( .A1(n7012), .A2(n9634), .ZN(n6679) );
  OR2_X1 U5415 ( .A1(n6550), .A2(n9636), .ZN(n6313) );
  AND4_X1 U5416 ( .A1(n5905), .A2(n5904), .A3(n5903), .A4(n5902), .ZN(n8270)
         );
  NAND2_X1 U5417 ( .A1(n5910), .A2(n6220), .ZN(n6193) );
  NAND2_X1 U5418 ( .A1(n9535), .A2(n5746), .ZN(n9490) );
  INV_X1 U5419 ( .A(n9999), .ZN(n10013) );
  INV_X1 U5420 ( .A(n10041), .ZN(n4841) );
  NAND2_X1 U5421 ( .A1(n10042), .A2(n10117), .ZN(n4840) );
  NAND2_X1 U5422 ( .A1(n6317), .A2(n10120), .ZN(n10276) );
  OAI22_X1 U5423 ( .A1(n5273), .A2(P1_D_REG_0__SCAN_IN), .B1(n5247), .B2(n5272), .ZN(n6273) );
  NOR2_X1 U5424 ( .A1(n5162), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n5165) );
  INV_X1 U5425 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5166) );
  XNOR2_X1 U5426 ( .A(n7382), .B(n7381), .ZN(n8200) );
  XNOR2_X1 U5427 ( .A(n7207), .B(n7206), .ZN(n8183) );
  XNOR2_X1 U5428 ( .A(n7314), .B(n7313), .ZN(n8149) );
  OAI21_X1 U5429 ( .B1(n7183), .B2(n4941), .A(n4938), .ZN(n7314) );
  AOI21_X1 U5430 ( .B1(n7308), .B2(n4940), .A(n4939), .ZN(n4938) );
  NAND2_X1 U5431 ( .A1(n7183), .A2(n7180), .ZN(n7309) );
  OAI21_X1 U5432 ( .B1(n5157), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5155) );
  NAND2_X1 U5433 ( .A1(n5155), .A2(n5156), .ZN(n5154) );
  NAND2_X1 U5434 ( .A1(n4953), .A2(n5636), .ZN(n5755) );
  XNOR2_X1 U5435 ( .A(n5634), .B(n5632), .ZN(n7252) );
  CLKBUF_X1 U5436 ( .A(n5122), .Z(n5124) );
  AND3_X1 U5437 ( .A1(n7560), .A2(n7559), .A3(n7558), .ZN(n8341) );
  NAND2_X1 U5438 ( .A1(n7453), .A2(n7452), .ZN(n7602) );
  AND4_X1 U5439 ( .A1(n7293), .A2(n7292), .A3(n7291), .A4(n7290), .ZN(n8329)
         );
  AND4_X1 U5440 ( .A1(n6620), .A2(n6619), .A3(n6618), .A4(n6617), .ZN(n7404)
         );
  AND3_X1 U5441 ( .A1(n7744), .A2(n7743), .A3(n7742), .ZN(n8720) );
  INV_X1 U5442 ( .A(n8253), .ZN(n8252) );
  NAND2_X1 U5443 ( .A1(n5076), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5077) );
  NAND2_X1 U5444 ( .A1(n7980), .A2(n7979), .ZN(n7982) );
  XNOR2_X1 U5445 ( .A(n5071), .B(P2_IR_REG_22__SCAN_IN), .ZN(n7986) );
  NAND2_X1 U5446 ( .A1(n5065), .A2(n4990), .ZN(n5070) );
  NAND2_X1 U5447 ( .A1(n7759), .A2(n7758), .ZN(n8704) );
  NAND4_X1 U5448 ( .A1(n5828), .A2(n5827), .A3(n5826), .A4(n5825), .ZN(n8427)
         );
  OR2_X1 U5449 ( .A1(P2_U3150), .A2(n5362), .ZN(n5939) );
  NAND2_X1 U5450 ( .A1(n6940), .A2(n6941), .ZN(n7157) );
  AND2_X1 U5451 ( .A1(n7859), .A2(n7858), .ZN(n8572) );
  NAND2_X1 U5452 ( .A1(n7871), .A2(n7870), .ZN(n8582) );
  NAND2_X1 U5453 ( .A1(n7728), .A2(n7727), .ZN(n8772) );
  AND3_X1 U5454 ( .A1(n6096), .A2(n6095), .A3(n6094), .ZN(n10309) );
  NAND2_X1 U5455 ( .A1(n7739), .A2(n7738), .ZN(n9205) );
  AND2_X1 U5456 ( .A1(n7208), .A2(n7395), .ZN(n5762) );
  INV_X1 U5457 ( .A(n9907), .ZN(n10071) );
  INV_X1 U5458 ( .A(n10159), .ZN(n9977) );
  NOR2_X1 U5459 ( .A1(n4894), .A2(n9365), .ZN(n4892) );
  NOR2_X1 U5460 ( .A1(n4895), .A2(n4898), .ZN(n4894) );
  NOR2_X1 U5461 ( .A1(n8230), .A2(n8215), .ZN(n4898) );
  INV_X1 U5462 ( .A(n4897), .ZN(n4895) );
  NAND2_X1 U5463 ( .A1(n4897), .A2(n4899), .ZN(n4896) );
  INV_X1 U5464 ( .A(n8230), .ZN(n4899) );
  AND4_X1 U5465 ( .A1(n6674), .A2(n6673), .A3(n6672), .A4(n6671), .ZN(n7414)
         );
  NAND2_X1 U5466 ( .A1(n8169), .A2(n8168), .ZN(n9877) );
  AND3_X1 U5467 ( .A1(n8079), .A2(n8078), .A3(n8077), .ZN(n9957) );
  AOI21_X1 U5468 ( .B1(n4889), .B2(n4887), .A(n4528), .ZN(n4886) );
  INV_X1 U5469 ( .A(n4889), .ZN(n4888) );
  NAND2_X1 U5470 ( .A1(n9980), .A2(n5533), .ZN(n9363) );
  NAND2_X1 U5471 ( .A1(n8178), .A2(n8177), .ZN(n9890) );
  OR2_X1 U5472 ( .A1(n9879), .A2(n8172), .ZN(n8178) );
  NAND2_X1 U5473 ( .A1(n5708), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4616) );
  NOR2_X1 U5474 ( .A1(n5457), .A2(n5456), .ZN(n5485) );
  NAND2_X1 U5475 ( .A1(n9759), .A2(n9758), .ZN(n4622) );
  OAI22_X1 U5476 ( .A1(n9754), .A2(n9752), .B1(n9757), .B2(n9751), .ZN(n4619)
         );
  OR2_X1 U5477 ( .A1(n9761), .A2(n5081), .ZN(n4620) );
  OAI21_X1 U5478 ( .B1(n4602), .B2(n4601), .A(n4600), .ZN(n4603) );
  INV_X1 U5479 ( .A(n4913), .ZN(n4601) );
  AOI21_X1 U5480 ( .B1(n4913), .B2(n9836), .A(n4562), .ZN(n4600) );
  NAND2_X1 U5481 ( .A1(n4842), .A2(n9809), .ZN(n10040) );
  NAND2_X1 U5482 ( .A1(n4843), .A2(n10009), .ZN(n4842) );
  OR2_X1 U5483 ( .A1(n5532), .A2(n10239), .ZN(n9980) );
  INV_X1 U5484 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5279) );
  NAND2_X1 U5485 ( .A1(n5589), .A2(n10175), .ZN(n5278) );
  INV_X1 U5486 ( .A(n9766), .ZN(n10125) );
  AOI21_X1 U5487 ( .B1(n4855), .B2(n10072), .A(n4854), .ZN(n10123) );
  INV_X1 U5488 ( .A(n10035), .ZN(n4854) );
  INV_X1 U5489 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10169) );
  NAND2_X1 U5490 ( .A1(n4994), .A2(n4999), .ZN(n4573) );
  NAND2_X1 U5491 ( .A1(n5991), .A2(n4572), .ZN(n4574) );
  MUX2_X1 U5492 ( .A(n7648), .B(n7647), .S(n7973), .Z(n7658) );
  NAND2_X1 U5493 ( .A1(n9374), .A2(n9471), .ZN(n4682) );
  AOI22_X1 U5494 ( .A1(n4685), .A2(n9374), .B1(n9379), .B2(n4684), .ZN(n4683)
         );
  NOR2_X1 U5495 ( .A1(n9380), .A2(n4643), .ZN(n4685) );
  NAND2_X1 U5496 ( .A1(n9375), .A2(n9379), .ZN(n4686) );
  OAI21_X1 U5497 ( .B1(n4808), .B2(n7682), .A(n7892), .ZN(n4807) );
  AOI21_X1 U5498 ( .B1(n7678), .B2(n4500), .A(n4539), .ZN(n4808) );
  OAI21_X1 U5499 ( .B1(n4806), .B2(n7673), .A(n7893), .ZN(n4805) );
  AOI21_X1 U5500 ( .B1(n7672), .B2(n4501), .A(n4538), .ZN(n4806) );
  AND2_X1 U5501 ( .A1(n4556), .A2(n4780), .ZN(n4775) );
  AND2_X1 U5502 ( .A1(n4774), .A2(n4772), .ZN(n4771) );
  INV_X1 U5503 ( .A(n4775), .ZN(n4772) );
  INV_X1 U5504 ( .A(n4674), .ZN(n4687) );
  AOI21_X1 U5505 ( .B1(n9376), .B2(n4520), .A(n4675), .ZN(n4674) );
  INV_X1 U5506 ( .A(n4782), .ZN(n4781) );
  OAI21_X1 U5507 ( .B1(n4784), .B2(n4791), .A(n4783), .ZN(n4782) );
  NAND2_X1 U5508 ( .A1(n4796), .A2(n7711), .ZN(n4783) );
  NAND2_X1 U5509 ( .A1(n4537), .A2(n4796), .ZN(n4784) );
  NAND2_X1 U5510 ( .A1(n4789), .A2(n4523), .ZN(n4787) );
  NAND2_X1 U5511 ( .A1(n4791), .A2(n4530), .ZN(n4789) );
  INV_X1 U5512 ( .A(n4790), .ZN(n4788) );
  NAND2_X1 U5513 ( .A1(n4775), .A2(n4776), .ZN(n4774) );
  INV_X1 U5514 ( .A(n4766), .ZN(n4765) );
  NOR2_X1 U5515 ( .A1(n4525), .A2(n4636), .ZN(n4635) );
  NAND2_X1 U5516 ( .A1(n7789), .A2(n7788), .ZN(n7805) );
  NAND2_X1 U5517 ( .A1(n7780), .A2(n7893), .ZN(n7789) );
  NAND2_X1 U5518 ( .A1(n9430), .A2(n9471), .ZN(n4673) );
  NOR2_X1 U5519 ( .A1(n9435), .A2(n4672), .ZN(n4671) );
  AND2_X1 U5520 ( .A1(n9429), .A2(n4643), .ZN(n4672) );
  NAND2_X1 U5521 ( .A1(n4667), .A2(n4665), .ZN(n9439) );
  AND2_X1 U5522 ( .A1(n6639), .A2(n6638), .ZN(n9384) );
  NAND2_X1 U5523 ( .A1(n9396), .A2(n6642), .ZN(n9388) );
  NAND2_X1 U5524 ( .A1(n7592), .A2(n7591), .ZN(n7615) );
  NAND2_X1 U5525 ( .A1(n6289), .A2(n6060), .ZN(n4948) );
  NOR2_X1 U5526 ( .A1(n4948), .A2(n4944), .ZN(n4943) );
  INV_X1 U5527 ( .A(n5981), .ZN(n4944) );
  INV_X1 U5528 ( .A(n5481), .ZN(n4746) );
  INV_X1 U5529 ( .A(n5479), .ZN(n4743) );
  INV_X1 U5530 ( .A(n8119), .ZN(n4986) );
  NOR2_X1 U5531 ( .A1(n8138), .A2(n4984), .ZN(n4981) );
  OAI21_X1 U5532 ( .B1(n8537), .B2(n7967), .A(n4533), .ZN(n4761) );
  AND2_X1 U5533 ( .A1(n4764), .A2(n4763), .ZN(n4762) );
  INV_X1 U5534 ( .A(n7968), .ZN(n4764) );
  NAND2_X1 U5535 ( .A1(n4813), .A2(n7883), .ZN(n4810) );
  NAND2_X1 U5536 ( .A1(n7167), .A2(n4707), .ZN(n7520) );
  NAND2_X1 U5537 ( .A1(n6959), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4707) );
  OR2_X1 U5538 ( .A1(n6608), .A2(n6607), .ZN(n6609) );
  AND2_X1 U5539 ( .A1(n6900), .A2(n7689), .ZN(n7922) );
  OAI21_X1 U5540 ( .B1(n5774), .B2(n5773), .A(n5772), .ZN(n5886) );
  NAND2_X1 U5541 ( .A1(n5810), .A2(P2_B_REG_SCAN_IN), .ZN(n8531) );
  OR2_X1 U5542 ( .A1(n7961), .A2(n7960), .ZN(n8601) );
  AND2_X1 U5543 ( .A1(n4548), .A2(n7956), .ZN(n4756) );
  NAND2_X1 U5544 ( .A1(n4545), .A2(n4957), .ZN(n8630) );
  INV_X1 U5545 ( .A(n8632), .ZN(n4957) );
  INV_X1 U5546 ( .A(n8542), .ZN(n4741) );
  NOR2_X1 U5547 ( .A1(n10189), .A2(n7256), .ZN(n7259) );
  INV_X1 U5548 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5059) );
  XNOR2_X1 U5549 ( .A(n5069), .B(P2_IR_REG_21__SCAN_IN), .ZN(n5786) );
  NAND2_X1 U5550 ( .A1(n5068), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5069) );
  OR2_X1 U5551 ( .A1(n4988), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n5064) );
  INV_X1 U5552 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5689) );
  AND2_X1 U5553 ( .A1(n5065), .A2(n5406), .ZN(n5614) );
  AND4_X1 U5554 ( .A1(n5223), .A2(n5036), .A3(n5035), .A4(n5034), .ZN(n4992)
         );
  INV_X1 U5555 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5034) );
  NOR2_X1 U5556 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5035) );
  NAND2_X1 U5557 ( .A1(n4992), .A2(n4968), .ZN(n5240) );
  INV_X1 U5558 ( .A(n5129), .ZN(n4968) );
  OR2_X1 U5559 ( .A1(n5205), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5225) );
  NOR2_X1 U5560 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5223) );
  NOR2_X1 U5561 ( .A1(n8009), .A2(n4881), .ZN(n4880) );
  INV_X1 U5562 ( .A(n7412), .ZN(n4881) );
  AND2_X1 U5563 ( .A1(n4878), .A2(n4872), .ZN(n4871) );
  NAND2_X1 U5564 ( .A1(n4880), .A2(n4873), .ZN(n4872) );
  NOR2_X1 U5565 ( .A1(n6556), .A2(n4869), .ZN(n4868) );
  NAND2_X1 U5566 ( .A1(n9456), .A2(n9457), .ZN(n4648) );
  AOI21_X1 U5567 ( .B1(n4647), .B2(n4646), .A(n9455), .ZN(n4645) );
  NOR2_X1 U5568 ( .A1(n9519), .A2(n9471), .ZN(n4646) );
  NAND2_X1 U5569 ( .A1(n9454), .A2(n9453), .ZN(n4647) );
  NAND2_X1 U5570 ( .A1(n9954), .A2(n9588), .ZN(n9795) );
  AND2_X1 U5571 ( .A1(n4664), .A2(n4660), .ZN(n4659) );
  OR2_X1 U5572 ( .A1(n9596), .A2(n4643), .ZN(n4660) );
  OR2_X1 U5573 ( .A1(n9367), .A2(n9845), .ZN(n9804) );
  OR2_X1 U5574 ( .A1(n9846), .A2(n9859), .ZN(n9803) );
  OR2_X1 U5575 ( .A1(n8075), .A2(n9256), .ZN(n8088) );
  OR2_X1 U5576 ( .A1(n7090), .A2(n9085), .ZN(n7213) );
  INV_X1 U5577 ( .A(n4497), .ZN(n4597) );
  INV_X1 U5578 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6846) );
  INV_X1 U5579 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6668) );
  OR2_X1 U5580 ( .A1(n7238), .A2(n9632), .ZN(n6836) );
  INV_X1 U5581 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6660) );
  AND2_X1 U5582 ( .A1(n6451), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6651) );
  INV_X1 U5583 ( .A(n4838), .ZN(n6643) );
  OAI21_X1 U5584 ( .B1(n9388), .B2(n9384), .A(n9398), .ZN(n4838) );
  NOR2_X1 U5585 ( .A1(n6300), .A2(n6299), .ZN(n6451) );
  NAND2_X1 U5586 ( .A1(n4837), .A2(n4836), .ZN(n9396) );
  INV_X1 U5587 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6213) );
  AND2_X1 U5588 ( .A1(n5736), .A2(n6339), .ZN(n4853) );
  NAND2_X1 U5589 ( .A1(n5745), .A2(n4521), .ZN(n9537) );
  NAND2_X1 U5590 ( .A1(n9895), .A2(n4498), .ZN(n9860) );
  NAND2_X1 U5591 ( .A1(n10018), .A2(n4527), .ZN(n9942) );
  NAND2_X1 U5592 ( .A1(n5745), .A2(n5744), .ZN(n4633) );
  INV_X1 U5593 ( .A(n9490), .ZN(n4632) );
  INV_X1 U5594 ( .A(n7315), .ZN(n5272) );
  NOR2_X1 U5595 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n4908) );
  AND2_X1 U5596 ( .A1(n7383), .A2(n7201), .ZN(n7381) );
  OR2_X1 U5597 ( .A1(n7188), .A2(n7187), .ZN(n7189) );
  AND2_X1 U5598 ( .A1(n7181), .A2(n7184), .ZN(n7182) );
  INV_X1 U5599 ( .A(n7180), .ZN(n4940) );
  INV_X1 U5600 ( .A(n7310), .ZN(n4939) );
  INV_X1 U5601 ( .A(n7308), .ZN(n4941) );
  OR2_X1 U5602 ( .A1(n6979), .A2(n6978), .ZN(n7183) );
  NAND2_X1 U5603 ( .A1(n5255), .A2(n6063), .ZN(n5020) );
  INV_X1 U5604 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5255) );
  INV_X1 U5605 ( .A(n5756), .ZN(n5757) );
  OAI21_X1 U5606 ( .B1(n5085), .B2(P2_DATAO_REG_2__SCAN_IN), .A(n4849), .ZN(
        n5095) );
  NAND2_X1 U5607 ( .A1(n5085), .A2(n4850), .ZN(n4849) );
  NAND3_X1 U5608 ( .A1(n6421), .A2(n5081), .A3(n4712), .ZN(n4956) );
  INV_X1 U5609 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4711) );
  AOI21_X1 U5610 ( .B1(n4962), .B2(n4960), .A(n4543), .ZN(n4959) );
  INV_X1 U5611 ( .A(n4962), .ZN(n4961) );
  INV_X1 U5612 ( .A(n8243), .ZN(n4960) );
  NOR2_X1 U5613 ( .A1(n7605), .A2(n4971), .ZN(n4970) );
  INV_X1 U5614 ( .A(n4973), .ZN(n4971) );
  NAND2_X1 U5615 ( .A1(n7601), .A2(n8421), .ZN(n4973) );
  NAND2_X1 U5616 ( .A1(n8241), .A2(n8242), .ZN(n8243) );
  NAND2_X1 U5617 ( .A1(n5821), .A2(n5810), .ZN(n5872) );
  OR3_X1 U5618 ( .A1(n7973), .A2(n6547), .A3(n5869), .ZN(n6085) );
  NAND2_X1 U5619 ( .A1(n8296), .A2(n8119), .ZN(n8396) );
  NAND2_X1 U5620 ( .A1(n4758), .A2(n4757), .ZN(n7976) );
  NAND2_X1 U5621 ( .A1(n4761), .A2(n4759), .ZN(n4758) );
  NAND2_X1 U5622 ( .A1(n7974), .A2(n4760), .ZN(n4757) );
  AOI21_X1 U5623 ( .B1(n7971), .B2(n7970), .A(n4760), .ZN(n4759) );
  NAND2_X1 U5624 ( .A1(n4811), .A2(n4809), .ZN(n7909) );
  AOI21_X1 U5625 ( .B1(n4813), .B2(n4812), .A(n7907), .ZN(n4811) );
  NAND2_X1 U5626 ( .A1(n4810), .A2(n7893), .ZN(n4809) );
  NOR2_X1 U5627 ( .A1(n7943), .A2(n7893), .ZN(n4812) );
  AND4_X1 U5628 ( .A1(n5044), .A2(n5043), .A3(n5063), .A4(n5042), .ZN(n4990)
         );
  AND4_X1 U5629 ( .A1(n5067), .A2(n5040), .A3(n5039), .A4(n5613), .ZN(n5043)
         );
  AND2_X1 U5630 ( .A1(n7800), .A2(n7799), .ZN(n8415) );
  NAND2_X1 U5631 ( .A1(n5501), .A2(n5502), .ZN(n5500) );
  XNOR2_X1 U5632 ( .A(n5954), .B(n5953), .ZN(n6005) );
  OAI22_X1 U5633 ( .A1(n6005), .A2(n6929), .B1(n6573), .B2(n6006), .ZN(n6007)
         );
  NAND2_X1 U5634 ( .A1(n6155), .A2(n6139), .ZN(n6140) );
  NAND2_X1 U5635 ( .A1(n6167), .A2(n6148), .ZN(n6149) );
  NAND2_X1 U5636 ( .A1(n6149), .A2(n6150), .ZN(n6380) );
  NAND2_X1 U5637 ( .A1(n6380), .A2(n4694), .ZN(n6511) );
  NAND2_X1 U5638 ( .A1(n6145), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4694) );
  NAND2_X1 U5639 ( .A1(n6529), .A2(n6530), .ZN(n6531) );
  NAND2_X1 U5640 ( .A1(n6945), .A2(n6946), .ZN(n6947) );
  NAND2_X1 U5641 ( .A1(n6947), .A2(n6948), .ZN(n7167) );
  XNOR2_X1 U5642 ( .A(n7514), .B(n7527), .ZN(n7158) );
  XNOR2_X1 U5643 ( .A(n7520), .B(n7527), .ZN(n7168) );
  NAND2_X1 U5644 ( .A1(n7157), .A2(n4691), .ZN(n7514) );
  NAND2_X1 U5645 ( .A1(n6959), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4691) );
  XNOR2_X1 U5646 ( .A(n8494), .B(n8477), .ZN(n8459) );
  NAND2_X1 U5647 ( .A1(n8459), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8498) );
  NOR2_X1 U5648 ( .A1(n7793), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n7814) );
  OR2_X1 U5649 ( .A1(n7642), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n7767) );
  NAND2_X1 U5650 ( .A1(n7954), .A2(n7953), .ZN(n8669) );
  INV_X1 U5651 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n7640) );
  NAND2_X1 U5652 ( .A1(n7754), .A2(n7640), .ZN(n7642) );
  INV_X1 U5653 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7751) );
  AND2_X1 U5654 ( .A1(n7752), .A2(n7751), .ZN(n7754) );
  OR2_X1 U5655 ( .A1(n7554), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n7740) );
  NOR2_X1 U5656 ( .A1(n7740), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n7752) );
  INV_X1 U5657 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7536) );
  AND2_X1 U5658 ( .A1(n7359), .A2(n7536), .ZN(n7474) );
  AND4_X1 U5659 ( .A1(n7271), .A2(n7270), .A3(n7269), .A4(n7268), .ZN(n10193)
         );
  AND4_X1 U5660 ( .A1(n6742), .A2(n6741), .A3(n6740), .A4(n6739), .ZN(n10191)
         );
  NAND2_X1 U5661 ( .A1(n6747), .A2(n6746), .ZN(n4704) );
  OR2_X1 U5662 ( .A1(n6614), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6616) );
  AND2_X1 U5663 ( .A1(n7706), .A2(n7701), .ZN(n7927) );
  INV_X1 U5664 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5348) );
  OR2_X1 U5665 ( .A1(n6934), .A2(n6969), .ZN(n6900) );
  AND2_X1 U5666 ( .A1(n7683), .A2(n7690), .ZN(n7921) );
  NAND2_X1 U5667 ( .A1(n6605), .A2(n7922), .ZN(n6905) );
  INV_X1 U5668 ( .A(n7922), .ZN(n7687) );
  OR2_X1 U5669 ( .A1(n6240), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6577) );
  AND2_X1 U5670 ( .A1(n6567), .A2(n6566), .ZN(n6771) );
  NAND2_X1 U5671 ( .A1(n6483), .A2(n6482), .ZN(n6497) );
  OR2_X1 U5672 ( .A1(n6480), .A2(n6479), .ZN(n6483) );
  AND2_X1 U5673 ( .A1(n7674), .A2(n7670), .ZN(n7915) );
  NAND2_X1 U5674 ( .A1(n6176), .A2(n6175), .ZN(n6180) );
  NAND2_X1 U5675 ( .A1(n7916), .A2(n6351), .ZN(n6350) );
  OR2_X1 U5676 ( .A1(n8430), .A2(n5995), .ZN(n7648) );
  INV_X1 U5677 ( .A(n8562), .ZN(n4716) );
  OR2_X1 U5678 ( .A1(n8532), .A2(n8564), .ZN(n8776) );
  AND2_X1 U5679 ( .A1(n7963), .A2(n8605), .ZN(n7964) );
  NAND2_X1 U5680 ( .A1(n8548), .A2(n8675), .ZN(n8680) );
  INV_X1 U5681 ( .A(n8678), .ZN(n8675) );
  AND2_X1 U5682 ( .A1(n7750), .A2(n7749), .ZN(n8547) );
  AOI21_X1 U5683 ( .B1(n7947), .B2(n4512), .A(n4740), .ZN(n4739) );
  NOR2_X1 U5684 ( .A1(n8543), .A2(n8720), .ZN(n4740) );
  NAND2_X1 U5685 ( .A1(n4738), .A2(n4736), .ZN(n8688) );
  NOR2_X1 U5686 ( .A1(n4737), .A2(n8545), .ZN(n4736) );
  INV_X1 U5687 ( .A(n4739), .ZN(n4737) );
  AOI21_X1 U5688 ( .B1(n7471), .B2(n4725), .A(n4722), .ZN(n4721) );
  NAND2_X1 U5689 ( .A1(n4723), .A2(n7550), .ZN(n4722) );
  NAND2_X1 U5690 ( .A1(n4725), .A2(n7470), .ZN(n4723) );
  NAND2_X1 U5691 ( .A1(n6735), .A2(n6734), .ZN(n7349) );
  OR2_X1 U5692 ( .A1(n7259), .A2(n7930), .ZN(n7273) );
  NAND2_X1 U5693 ( .A1(n5865), .A2(n6177), .ZN(n10336) );
  AND3_X1 U5694 ( .A1(n6237), .A2(n6236), .A3(n6235), .ZN(n10314) );
  AND2_X1 U5695 ( .A1(n5785), .A2(n4976), .ZN(n4975) );
  INV_X1 U5696 ( .A(n5819), .ZN(n5885) );
  AND2_X1 U5697 ( .A1(n5988), .A2(n5975), .ZN(n8458) );
  INV_X1 U5698 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5406) );
  NAND2_X1 U5699 ( .A1(n6555), .A2(n6556), .ZN(n6992) );
  AND2_X1 U5700 ( .A1(n8089), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8101) );
  AND2_X1 U5701 ( .A1(n8165), .A2(n8160), .ZN(n9290) );
  NAND2_X1 U5702 ( .A1(n4867), .A2(n4869), .ZN(n4866) );
  NAND2_X1 U5703 ( .A1(n4903), .A2(n4901), .ZN(n9331) );
  AND2_X1 U5704 ( .A1(n4902), .A2(n4904), .ZN(n4901) );
  NAND2_X1 U5705 ( .A1(n4905), .A2(n8022), .ZN(n4902) );
  INV_X1 U5706 ( .A(n8166), .ZN(n4887) );
  NAND2_X1 U5707 ( .A1(n4579), .A2(n9236), .ZN(n4578) );
  INV_X1 U5708 ( .A(n5301), .ZN(n9602) );
  AND4_X1 U5709 ( .A1(n6457), .A2(n6456), .A3(n6455), .A4(n6454), .ZN(n7013)
         );
  NAND2_X1 U5710 ( .A1(n9477), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5711) );
  NOR2_X1 U5711 ( .A1(n4989), .A2(n4996), .ZN(n5710) );
  AND2_X1 U5712 ( .A1(n9715), .A2(n9716), .ZN(n9713) );
  INV_X1 U5713 ( .A(n5176), .ZN(n9652) );
  NOR2_X1 U5714 ( .A1(n7503), .A2(n7502), .ZN(n7581) );
  NOR2_X1 U5715 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5018) );
  INV_X1 U5716 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5005) );
  OR2_X1 U5717 ( .A1(n9731), .A2(n9732), .ZN(n9749) );
  XNOR2_X1 U5718 ( .A(n4844), .B(n9805), .ZN(n4843) );
  NAND2_X1 U5719 ( .A1(n9818), .A2(n9804), .ZN(n4844) );
  AND2_X1 U5720 ( .A1(n8232), .A2(n8221), .ZN(n9829) );
  NOR2_X1 U5721 ( .A1(n9824), .A2(n4914), .ZN(n4913) );
  INV_X1 U5722 ( .A(n9791), .ZN(n4914) );
  AND4_X1 U5723 ( .A1(n8191), .A2(n8190), .A3(n8189), .A4(n8188), .ZN(n9842)
         );
  INV_X1 U5724 ( .A(n8203), .ZN(n8219) );
  OAI21_X1 U5725 ( .B1(n4614), .B2(n4613), .A(n4922), .ZN(n9788) );
  INV_X1 U5726 ( .A(n4923), .ZN(n4613) );
  NAND2_X1 U5727 ( .A1(n4928), .A2(n4496), .ZN(n4925) );
  NAND2_X1 U5728 ( .A1(n9895), .A2(n10141), .ZN(n9874) );
  NAND2_X1 U5729 ( .A1(n4820), .A2(n4818), .ZN(n9908) );
  INV_X1 U5730 ( .A(n4819), .ZN(n4818) );
  OAI21_X1 U5731 ( .B1(n4822), .B2(n9588), .A(n9796), .ZN(n4819) );
  NAND2_X1 U5732 ( .A1(n9969), .A2(n9587), .ZN(n9954) );
  AND2_X1 U5733 ( .A1(n9487), .A2(n9587), .ZN(n9975) );
  NAND2_X1 U5734 ( .A1(n10018), .A2(n4859), .ZN(n9979) );
  AOI21_X1 U5735 ( .B1(n4833), .B2(n4835), .A(n4831), .ZN(n4830) );
  INV_X1 U5736 ( .A(n9584), .ZN(n4831) );
  NAND2_X1 U5737 ( .A1(n10018), .A2(n9993), .ZN(n9988) );
  NAND2_X1 U5738 ( .A1(n4612), .A2(n4916), .ZN(n9987) );
  NAND2_X1 U5739 ( .A1(n10165), .A2(n9779), .ZN(n4916) );
  AND2_X1 U5740 ( .A1(n9585), .A2(n9586), .ZN(n9996) );
  NAND2_X1 U5741 ( .A1(n4832), .A2(n9582), .ZN(n10008) );
  NAND2_X1 U5742 ( .A1(n9581), .A2(n9580), .ZN(n4832) );
  OAI21_X1 U5743 ( .B1(n4847), .B2(n4846), .A(n4845), .ZN(n7088) );
  INV_X1 U5744 ( .A(n9412), .ZN(n4846) );
  NAND2_X1 U5745 ( .A1(n6837), .A2(n6836), .ZN(n6840) );
  NAND2_X1 U5746 ( .A1(n6840), .A2(n9502), .ZN(n7074) );
  OR2_X1 U5747 ( .A1(n6996), .A2(n4836), .ZN(n6677) );
  NAND2_X1 U5748 ( .A1(n6449), .A2(n6450), .ZN(n6678) );
  NAND2_X1 U5749 ( .A1(n6430), .A2(n6199), .ZN(n6210) );
  AND4_X1 U5750 ( .A1(n6205), .A2(n6204), .A3(n6203), .A4(n6202), .ZN(n6549)
         );
  AND2_X1 U5751 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5901) );
  INV_X1 U5752 ( .A(n5742), .ZN(n6254) );
  NAND2_X1 U5753 ( .A1(n6802), .A2(n5736), .ZN(n6801) );
  AND2_X1 U5754 ( .A1(n5529), .A2(n5526), .ZN(n6276) );
  NAND2_X1 U5755 ( .A1(n8151), .A2(n8150), .ZN(n9786) );
  INV_X1 U5756 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4608) );
  INV_X1 U5757 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5158) );
  INV_X1 U5758 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5260) );
  NOR2_X1 U5759 ( .A1(n5020), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n5013) );
  INV_X1 U5760 ( .A(n5252), .ZN(n4870) );
  AND2_X1 U5761 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5257) );
  INV_X1 U5762 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U5763 ( .A1(n4945), .A2(n6060), .ZN(n6293) );
  NAND2_X1 U5764 ( .A1(n4952), .A2(n4950), .ZN(n4945) );
  NAND2_X1 U5765 ( .A1(n5983), .A2(n5981), .ZN(n4952) );
  NAND2_X1 U5766 ( .A1(n4949), .A2(n5981), .ZN(n6059) );
  NAND2_X1 U5767 ( .A1(n4747), .A2(n5481), .ZN(n5547) );
  XNOR2_X1 U5768 ( .A(n5229), .B(n5228), .ZN(n6587) );
  INV_X1 U5769 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5016) );
  XNOR2_X1 U5770 ( .A(n5194), .B(n5192), .ZN(n6206) );
  NAND2_X1 U5771 ( .A1(n5094), .A2(n5093), .ZN(n5698) );
  OR2_X1 U5772 ( .A1(n5100), .A2(n10169), .ZN(n5410) );
  BUF_X8 U5773 ( .A(n5110), .Z(n7901) );
  AND2_X1 U5774 ( .A1(n6790), .A2(n6773), .ZN(n6775) );
  NAND2_X1 U5775 ( .A1(n8116), .A2(n8293), .ZN(n8296) );
  AND2_X1 U5776 ( .A1(n7802), .A2(n7801), .ZN(n8550) );
  AND4_X1 U5777 ( .A1(n7364), .A2(n7363), .A3(n7362), .A4(n7361), .ZN(n8345)
         );
  NAND2_X1 U5778 ( .A1(n7792), .A2(n7791), .ZN(n8642) );
  NAND2_X1 U5779 ( .A1(n4972), .A2(n4973), .ZN(n7604) );
  OAI21_X1 U5780 ( .B1(n8245), .B2(n8244), .A(n8243), .ZN(n8366) );
  NOR2_X1 U5781 ( .A1(n7399), .A2(n8422), .ZN(n4958) );
  NAND2_X1 U5782 ( .A1(n7825), .A2(n7824), .ZN(n8557) );
  NAND2_X1 U5783 ( .A1(n5841), .A2(n5840), .ZN(n8406) );
  INV_X1 U5784 ( .A(n8566), .ZN(n8588) );
  INV_X1 U5785 ( .A(n8596), .ZN(n8560) );
  INV_X1 U5786 ( .A(n8415), .ZN(n8653) );
  NAND2_X1 U5787 ( .A1(n7773), .A2(n7772), .ZN(n8662) );
  INV_X1 U5788 ( .A(n8416), .ZN(n8681) );
  INV_X1 U5789 ( .A(n8329), .ZN(n8418) );
  INV_X1 U5790 ( .A(n10191), .ZN(n8421) );
  AND4_X1 U5791 ( .A1(n5333), .A2(n5332), .A3(n5331), .A4(n5330), .ZN(n7066)
         );
  AND4_X1 U5792 ( .A1(n5354), .A2(n5353), .A3(n5352), .A4(n5351), .ZN(n7443)
         );
  AND4_X1 U5793 ( .A1(n5326), .A2(n5325), .A3(n5324), .A4(n5323), .ZN(n7439)
         );
  NAND4_X1 U5794 ( .A1(n5817), .A2(n5816), .A3(n5815), .A4(n5814), .ZN(n8428)
         );
  OR2_X1 U5795 ( .A1(n7288), .A2(n5931), .ZN(n5792) );
  OR2_X1 U5796 ( .A1(n5834), .A2(n5060), .ZN(n8485) );
  INV_X1 U5797 ( .A(n5939), .ZN(n8519) );
  XNOR2_X1 U5798 ( .A(n5185), .B(P2_IR_REG_4__SCAN_IN), .ZN(n8447) );
  XNOR2_X1 U5799 ( .A(n6147), .B(n6588), .ZN(n6168) );
  XNOR2_X1 U5800 ( .A(n6511), .B(n6730), .ZN(n6381) );
  NAND2_X1 U5801 ( .A1(n6938), .A2(n6939), .ZN(n6940) );
  NAND2_X1 U5802 ( .A1(n8474), .A2(n8475), .ZN(n8504) );
  AOI21_X1 U5803 ( .B1(n8498), .B2(n8496), .A(n8497), .ZN(n8507) );
  AOI21_X1 U5804 ( .B1(n9459), .B2(n7873), .A(n7848), .ZN(n8735) );
  AND2_X1 U5805 ( .A1(n4714), .A2(n4715), .ZN(n8737) );
  INV_X1 U5806 ( .A(n8569), .ZN(n4715) );
  OR2_X1 U5807 ( .A1(n8572), .A2(n7860), .ZN(n8581) );
  NAND2_X1 U5808 ( .A1(n8669), .A2(n8668), .ZN(n8757) );
  NAND2_X1 U5809 ( .A1(n6572), .A2(n6571), .ZN(n10333) );
  NAND2_X1 U5810 ( .A1(n6575), .A2(n6574), .ZN(n6934) );
  NAND2_X1 U5811 ( .A1(n6206), .A2(n7873), .ZN(n6575) );
  AOI22_X1 U5812 ( .A1(n7737), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7736), .B2(
        n6573), .ZN(n6574) );
  AND3_X1 U5813 ( .A1(n6038), .A2(n6037), .A3(n6036), .ZN(n10306) );
  NAND2_X1 U5814 ( .A1(n8724), .A2(n10196), .ZN(n8729) );
  NOR2_X2 U5815 ( .A1(n5883), .A2(n5819), .ZN(n8709) );
  INV_X1 U5816 ( .A(n8729), .ZN(n8670) );
  INV_X1 U5817 ( .A(n8610), .ZN(n8726) );
  INV_X1 U5818 ( .A(n8752), .ZN(n8768) );
  AND3_X2 U5819 ( .A1(n6172), .A2(n5889), .A3(n6174), .ZN(n10381) );
  INV_X1 U5820 ( .A(n8582), .ZN(n9157) );
  AND2_X1 U5821 ( .A1(n4730), .A2(n4936), .ZN(n8577) );
  NAND2_X1 U5822 ( .A1(n7835), .A2(n7834), .ZN(n9163) );
  INV_X1 U5823 ( .A(n8557), .ZN(n9170) );
  NAND2_X1 U5824 ( .A1(n7813), .A2(n7812), .ZN(n9173) );
  INV_X1 U5825 ( .A(n8550), .ZN(n9185) );
  NAND2_X1 U5826 ( .A1(n4701), .A2(n4702), .ZN(n8647) );
  NAND2_X1 U5827 ( .A1(n7639), .A2(n7638), .ZN(n9192) );
  INV_X1 U5828 ( .A(n8547), .ZN(n9198) );
  NAND2_X1 U5829 ( .A1(n8716), .A2(n8542), .ZN(n8700) );
  NAND2_X1 U5830 ( .A1(n7946), .A2(n7945), .ZN(n8713) );
  AND2_X1 U5831 ( .A1(n7482), .A2(n7481), .ZN(n7488) );
  NAND2_X1 U5832 ( .A1(n7355), .A2(n7354), .ZN(n8393) );
  NAND2_X1 U5833 ( .A1(n7371), .A2(n7370), .ZN(n7372) );
  NAND2_X1 U5834 ( .A1(n7264), .A2(n7263), .ZN(n8299) );
  INV_X1 U5835 ( .A(n9178), .ZN(n9204) );
  NAND2_X1 U5836 ( .A1(n10364), .A2(n10358), .ZN(n9212) );
  NAND2_X1 U5837 ( .A1(n10364), .A2(n10363), .ZN(n9178) );
  AND2_X1 U5838 ( .A1(n6089), .A2(n6088), .ZN(n10366) );
  OR2_X1 U5839 ( .A1(n6084), .A2(n6083), .ZN(n6089) );
  OR2_X1 U5840 ( .A1(n6087), .A2(n6086), .ZN(n6088) );
  AND2_X1 U5841 ( .A1(n5833), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5214) );
  AND2_X1 U5842 ( .A1(n4816), .A2(n5316), .ZN(n4815) );
  XNOR2_X1 U5843 ( .A(n5317), .B(n5316), .ZN(n7593) );
  OR2_X1 U5844 ( .A1(n5315), .A2(n5314), .ZN(n5317) );
  NAND2_X1 U5845 ( .A1(n5076), .A2(n5052), .ZN(n7208) );
  INV_X1 U5846 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7811) );
  NAND2_X1 U5847 ( .A1(n5055), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5047) );
  INV_X1 U5848 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7790) );
  INV_X1 U5849 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8788) );
  INV_X1 U5850 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8840) );
  INV_X1 U5851 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7637) );
  INV_X1 U5852 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7748) );
  INV_X1 U5853 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6298) );
  INV_X1 U5854 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6122) );
  INV_X1 U5855 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n5990) );
  INV_X1 U5856 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5976) );
  INV_X1 U5857 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n9068) );
  INV_X1 U5858 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n8874) );
  XNOR2_X1 U5859 ( .A(n5376), .B(n5375), .ZN(n7993) );
  NAND2_X1 U5860 ( .A1(n5154), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5014) );
  AND3_X1 U5861 ( .A1(n8064), .A2(n8063), .A3(n8062), .ZN(n9941) );
  NAND2_X1 U5862 ( .A1(n6363), .A2(n4587), .ZN(n6265) );
  INV_X1 U5863 ( .A(n6263), .ZN(n4585) );
  AND3_X1 U5864 ( .A1(n8037), .A2(n8036), .A3(n8035), .ZN(n10014) );
  NAND2_X1 U5865 ( .A1(n4907), .A2(n8021), .ZN(n9283) );
  NOR2_X1 U5866 ( .A1(n5719), .A2(n5718), .ZN(n8268) );
  AND4_X1 U5867 ( .A1(n6219), .A2(n6218), .A3(n6217), .A4(n6216), .ZN(n7113)
         );
  NAND2_X1 U5868 ( .A1(n5726), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9314) );
  AOI21_X1 U5869 ( .B1(n9248), .B2(n9249), .A(n8056), .ZN(n9302) );
  AOI21_X1 U5870 ( .B1(n7413), .B2(n7412), .A(n4877), .ZN(n8010) );
  INV_X1 U5871 ( .A(n4883), .ZN(n4877) );
  NAND2_X1 U5872 ( .A1(n9254), .A2(n9255), .ZN(n4581) );
  AND4_X1 U5873 ( .A1(n6666), .A2(n6665), .A3(n6664), .A4(n6663), .ZN(n7420)
         );
  NAND2_X1 U5874 ( .A1(n6650), .A2(n6649), .ZN(n7031) );
  INV_X1 U5875 ( .A(n9360), .ZN(n9334) );
  INV_X1 U5876 ( .A(n9339), .ZN(n4591) );
  NAND2_X1 U5877 ( .A1(n7080), .A2(n7079), .ZN(n9418) );
  NAND2_X1 U5878 ( .A1(n4650), .A2(n4655), .ZN(n9616) );
  NAND2_X1 U5879 ( .A1(n9481), .A2(n4658), .ZN(n4650) );
  INV_X1 U5880 ( .A(n9577), .ZN(n9604) );
  AOI21_X1 U5881 ( .B1(n4653), .B2(n4655), .A(n4652), .ZN(n4651) );
  NAND2_X1 U5882 ( .A1(n8107), .A2(n8106), .ZN(n9913) );
  OR2_X1 U5883 ( .A1(n9897), .A2(n8172), .ZN(n8107) );
  INV_X1 U5884 ( .A(n9924), .ZN(n9891) );
  INV_X1 U5885 ( .A(n10014), .ZN(n9971) );
  INV_X1 U5886 ( .A(n10012), .ZN(n9775) );
  INV_X1 U5887 ( .A(n6549), .ZN(n9636) );
  INV_X1 U5888 ( .A(n8270), .ZN(n9638) );
  AND2_X1 U5889 ( .A1(n5601), .A2(n5600), .ZN(n5603) );
  NAND2_X1 U5890 ( .A1(n9687), .A2(n9688), .ZN(n9686) );
  NOR2_X1 U5891 ( .A1(n5443), .A2(n5442), .ZN(n5441) );
  AND2_X1 U5892 ( .A1(n9686), .A2(n4628), .ZN(n5443) );
  NAND2_X1 U5893 ( .A1(n9685), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4628) );
  NOR2_X1 U5894 ( .A1(n5466), .A2(n4557), .ZN(n5457) );
  NOR2_X1 U5895 ( .A1(n5485), .A2(n4623), .ZN(n5486) );
  NOR2_X1 U5896 ( .A1(n4625), .A2(n4624), .ZN(n4623) );
  INV_X1 U5897 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n4624) );
  INV_X1 U5898 ( .A(n6309), .ZN(n4625) );
  NAND2_X1 U5899 ( .A1(n5486), .A2(n5487), .ZN(n5679) );
  NOR2_X1 U5900 ( .A1(n5857), .A2(n5858), .ZN(n6075) );
  NOR2_X1 U5901 ( .A1(n5855), .A2(n4627), .ZN(n5858) );
  AND2_X1 U5902 ( .A1(n6644), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4627) );
  NOR2_X1 U5903 ( .A1(n6075), .A2(n4626), .ZN(n6078) );
  AND2_X1 U5904 ( .A1(n6648), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4626) );
  NAND2_X1 U5905 ( .A1(n6078), .A2(n6077), .ZN(n7140) );
  XNOR2_X1 U5906 ( .A(n7501), .B(n7500), .ZN(n7145) );
  NOR2_X1 U5907 ( .A1(n7145), .A2(n7144), .ZN(n7502) );
  AND2_X1 U5908 ( .A1(n9753), .A2(n5176), .ZN(n9755) );
  AND2_X1 U5909 ( .A1(n9461), .A2(n9460), .ZN(n9814) );
  NAND2_X1 U5910 ( .A1(n9867), .A2(n9800), .ZN(n9855) );
  NAND2_X1 U5911 ( .A1(n4926), .A2(n4928), .ZN(n9885) );
  NAND2_X1 U5912 ( .A1(n9920), .A2(n4929), .ZN(n4926) );
  AOI21_X1 U5913 ( .B1(n7995), .B2(n9467), .A(n4997), .ZN(n9907) );
  INV_X1 U5914 ( .A(n4934), .ZN(n4931) );
  NAND2_X1 U5915 ( .A1(n9920), .A2(n9785), .ZN(n4932) );
  NAND2_X1 U5916 ( .A1(n4824), .A2(n4507), .ZN(n9922) );
  NAND2_X1 U5917 ( .A1(n4825), .A2(n9588), .ZN(n4824) );
  NAND2_X1 U5918 ( .A1(n7212), .A2(n7211), .ZN(n10111) );
  NAND2_X1 U5919 ( .A1(n4594), .A2(n4497), .ZN(n7210) );
  NAND2_X1 U5920 ( .A1(n6837), .A2(n4598), .ZN(n4594) );
  NAND2_X1 U5921 ( .A1(n7087), .A2(n9553), .ZN(n7334) );
  NAND2_X1 U5922 ( .A1(n6193), .A2(n6192), .ZN(n6428) );
  INV_X1 U5923 ( .A(n10030), .ZN(n9976) );
  INV_X2 U5924 ( .A(n10290), .ZN(n10293) );
  NAND2_X1 U5925 ( .A1(n4841), .A2(n4840), .ZN(n4839) );
  INV_X1 U5926 ( .A(n9877), .ZN(n10141) );
  INV_X1 U5927 ( .A(n9786), .ZN(n10145) );
  AND2_X1 U5928 ( .A1(n8045), .A2(n8044), .ZN(n10159) );
  INV_X1 U5929 ( .A(n9418), .ZN(n7432) );
  NAND2_X1 U5930 ( .A1(n6839), .A2(n6838), .ZN(n7422) );
  INV_X1 U5931 ( .A(n6550), .ZN(n6633) );
  NAND2_X1 U5932 ( .A1(n5712), .A2(n5783), .ZN(n5592) );
  NAND2_X1 U5933 ( .A1(n6985), .A2(n5246), .ZN(n10239) );
  AND2_X1 U5934 ( .A1(n5519), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5246) );
  INV_X1 U5935 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5287) );
  NAND2_X1 U5936 ( .A1(n5291), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5288) );
  NAND2_X1 U5937 ( .A1(n5163), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5164) );
  INV_X1 U5938 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9079) );
  INV_X1 U5939 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7316) );
  INV_X1 U5940 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n9073) );
  XNOR2_X1 U5941 ( .A(n7309), .B(n7308), .ZN(n7995) );
  INV_X1 U5942 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7991) );
  INV_X1 U5943 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6811) );
  INV_X1 U5944 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8277) );
  INV_X1 U5945 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5992) );
  INV_X1 U5946 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n5850) );
  OR2_X1 U5947 ( .A1(n5542), .A2(n5541), .ZN(n7150) );
  INV_X1 U5948 ( .A(n6206), .ZN(n5209) );
  INV_X1 U5949 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5015) );
  AND2_X1 U5950 ( .A1(n5126), .A2(n5125), .ZN(n5906) );
  XNOR2_X1 U5951 ( .A(n5410), .B(P1_IR_REG_2__SCAN_IN), .ZN(n9658) );
  NAND2_X1 U5952 ( .A1(n5368), .A2(n5810), .ZN(n5080) );
  NAND2_X1 U5953 ( .A1(n6099), .A2(n6098), .ZN(n6101) );
  XNOR2_X1 U5954 ( .A(n7982), .B(n8523), .ZN(n7989) );
  NAND2_X1 U5955 ( .A1(n4896), .A2(n9342), .ZN(n4893) );
  NAND2_X1 U5956 ( .A1(n4619), .A2(n9621), .ZN(n4618) );
  NAND2_X1 U5957 ( .A1(n4622), .A2(n5281), .ZN(n4621) );
  OAI21_X1 U5958 ( .B1(n10123), .B2(n10278), .A(n4856), .ZN(P1_U3521) );
  INV_X1 U5959 ( .A(n4857), .ZN(n4856) );
  OAI22_X1 U5960 ( .A1(n10125), .A2(n10164), .B1(n10280), .B2(n10124), .ZN(
        n4857) );
  OR2_X1 U5962 ( .A1(n9786), .A2(n9913), .ZN(n4496) );
  NAND2_X1 U5963 ( .A1(n7957), .A2(n7956), .ZN(n8599) );
  INV_X1 U5964 ( .A(n9921), .ZN(n4823) );
  OR2_X1 U5965 ( .A1(n4918), .A2(n7077), .ZN(n4497) );
  NAND2_X1 U5966 ( .A1(n8087), .A2(n8086), .ZN(n10079) );
  AND2_X1 U5967 ( .A1(n10141), .A2(n4864), .ZN(n4498) );
  OR2_X1 U5968 ( .A1(n7273), .A2(n7714), .ZN(n4499) );
  AND2_X1 U5969 ( .A1(n7677), .A2(n7676), .ZN(n4500) );
  AND4_X1 U5970 ( .A1(n5919), .A2(n5918), .A3(n5917), .A4(n5916), .ZN(n6365)
         );
  NAND2_X1 U5971 ( .A1(n5100), .A2(n4569), .ZN(n5112) );
  AND2_X1 U5972 ( .A1(n7671), .A2(n7679), .ZN(n4501) );
  AND2_X1 U5973 ( .A1(n9786), .A2(n9913), .ZN(n4502) );
  INV_X1 U5974 ( .A(n10165), .ZN(n10020) );
  AND2_X1 U5975 ( .A1(n8025), .A2(n8024), .ZN(n10165) );
  AND2_X1 U5976 ( .A1(n4498), .A2(n4863), .ZN(n4503) );
  AND2_X1 U5977 ( .A1(n4630), .A2(n4608), .ZN(n4504) );
  INV_X1 U5978 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4630) );
  AND2_X1 U5979 ( .A1(n8074), .A2(n8073), .ZN(n10151) );
  INV_X1 U5980 ( .A(n10151), .ZN(n9944) );
  AND4_X1 U5981 ( .A1(n6305), .A2(n6304), .A3(n6303), .A4(n6302), .ZN(n7041)
         );
  INV_X1 U5982 ( .A(n7041), .ZN(n4836) );
  NAND2_X1 U5983 ( .A1(n9621), .A2(n9577), .ZN(n5516) );
  INV_X1 U5984 ( .A(n7238), .ZN(n4861) );
  AND2_X1 U5985 ( .A1(n5690), .A2(n5759), .ZN(n7262) );
  INV_X1 U5986 ( .A(n10300), .ZN(n5868) );
  AND2_X1 U5987 ( .A1(n5280), .A2(n5281), .ZN(n9471) );
  AND2_X1 U5988 ( .A1(n5589), .A2(n5085), .ZN(n5895) );
  NAND2_X1 U5989 ( .A1(n4983), .A2(n4982), .ZN(n8309) );
  XNOR2_X1 U5990 ( .A(n5313), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5320) );
  INV_X1 U5991 ( .A(n5589), .ZN(n8043) );
  NAND2_X1 U5992 ( .A1(n7630), .A2(n7629), .ZN(n8246) );
  AND2_X1 U5993 ( .A1(n9895), .A2(n4503), .ZN(n4505) );
  AND3_X1 U5994 ( .A1(n5724), .A2(n5723), .A3(n5722), .ZN(n4506) );
  AND2_X1 U5995 ( .A1(n7726), .A2(n7729), .ZN(n7470) );
  AND2_X1 U5996 ( .A1(n4826), .A2(n9794), .ZN(n4507) );
  AND2_X1 U5997 ( .A1(n9381), .A2(n9543), .ZN(n4508) );
  XOR2_X1 U5998 ( .A(n8550), .B(n8258), .Z(n4509) );
  INV_X1 U5999 ( .A(n6804), .ZN(n5739) );
  AND2_X1 U6000 ( .A1(n4969), .A2(n4992), .ZN(n5065) );
  OAI21_X1 U6001 ( .B1(n9927), .B2(n8172), .A(n8095), .ZN(n9914) );
  NOR2_X1 U6002 ( .A1(n4801), .A2(n4802), .ZN(n5049) );
  AND2_X1 U6003 ( .A1(n5589), .A2(n7901), .ZN(n5712) );
  NAND4_X1 U6004 ( .A1(n4610), .A2(n4607), .A3(n4631), .A4(n5168), .ZN(n5291)
         );
  INV_X1 U6005 ( .A(n7276), .ZN(n7714) );
  AND2_X1 U6006 ( .A1(n7718), .A2(n7717), .ZN(n7276) );
  OR2_X1 U6007 ( .A1(n8550), .A2(n8549), .ZN(n4510) );
  AND3_X1 U6008 ( .A1(n8393), .A2(n8329), .A3(n7892), .ZN(n4511) );
  INV_X1 U6009 ( .A(n9553), .ZN(n4848) );
  INV_X1 U6010 ( .A(n9588), .ZN(n4828) );
  NOR2_X1 U6011 ( .A1(n4741), .A2(n8544), .ZN(n4512) );
  NAND2_X1 U6012 ( .A1(n5725), .A2(n4506), .ZN(n5742) );
  AND3_X1 U6013 ( .A1(n10362), .A2(n10191), .A3(n7893), .ZN(n4513) );
  OR2_X1 U6014 ( .A1(n5810), .A2(n5784), .ZN(n4514) );
  NAND2_X1 U6015 ( .A1(n8099), .A2(n4580), .ZN(n8163) );
  AND2_X1 U6016 ( .A1(n5336), .A2(n5230), .ZN(n4515) );
  AND4_X1 U6017 ( .A1(n5156), .A2(n5158), .A3(n5260), .A4(n5019), .ZN(n4516)
         );
  AND2_X1 U6018 ( .A1(n6774), .A2(n6773), .ZN(n4517) );
  AND2_X1 U6019 ( .A1(n9907), .A2(n9924), .ZN(n4518) );
  OR2_X1 U6020 ( .A1(n8331), .A2(n8345), .ZN(n7726) );
  INV_X1 U6021 ( .A(n7726), .ZN(n4776) );
  NOR2_X1 U6022 ( .A1(n7901), .A2(n5783), .ZN(n4519) );
  AND2_X1 U6023 ( .A1(n9375), .A2(n4508), .ZN(n4520) );
  INV_X1 U6024 ( .A(n9574), .ZN(n9614) );
  AND2_X1 U6025 ( .A1(n5744), .A2(n5746), .ZN(n4521) );
  NOR2_X1 U6026 ( .A1(n8582), .A2(n8588), .ZN(n4522) );
  INV_X1 U6027 ( .A(n10116), .ZN(n9247) );
  NAND2_X1 U6028 ( .A1(n7076), .A2(n7075), .ZN(n10116) );
  AND2_X1 U6029 ( .A1(n4796), .A2(n4788), .ZN(n4523) );
  XNOR2_X1 U6030 ( .A(n4603), .B(n9793), .ZN(n10039) );
  AND2_X1 U6031 ( .A1(n9801), .A2(n9800), .ZN(n4524) );
  AND2_X1 U6032 ( .A1(n8031), .A2(n8030), .ZN(n9993) );
  INV_X1 U6033 ( .A(n9993), .ZN(n10099) );
  AND2_X1 U6034 ( .A1(n9406), .A2(n9405), .ZN(n4525) );
  INV_X1 U6035 ( .A(n9367), .ZN(n10133) );
  NAND2_X1 U6036 ( .A1(n8218), .A2(n8217), .ZN(n9367) );
  OR2_X1 U6037 ( .A1(n7006), .A2(n7003), .ZN(n4526) );
  AND2_X1 U6038 ( .A1(n4858), .A2(n10151), .ZN(n4527) );
  OR2_X1 U6039 ( .A1(n9340), .A2(n9341), .ZN(n4528) );
  AND2_X1 U6040 ( .A1(n4503), .A2(n10133), .ZN(n4529) );
  AND2_X1 U6041 ( .A1(n9804), .A2(n9483), .ZN(n9824) );
  NAND2_X1 U6042 ( .A1(n7704), .A2(n4794), .ZN(n4530) );
  NOR2_X1 U6043 ( .A1(n10116), .A2(n9630), .ZN(n7077) );
  INV_X1 U6044 ( .A(n7073), .ZN(n4920) );
  OR2_X1 U6045 ( .A1(n7422), .A2(n9631), .ZN(n7073) );
  INV_X1 U6046 ( .A(n6198), .ZN(n10254) );
  NOR2_X1 U6047 ( .A1(n7432), .A2(n9241), .ZN(n4531) );
  OR2_X1 U6048 ( .A1(n8246), .A2(n8416), .ZN(n7955) );
  OR2_X1 U6049 ( .A1(n4661), .A2(n9471), .ZN(n4532) );
  INV_X1 U6050 ( .A(n7229), .ZN(n4884) );
  INV_X1 U6051 ( .A(n4879), .ZN(n4878) );
  OAI21_X1 U6052 ( .B1(n8009), .B2(n4883), .A(n4882), .ZN(n4879) );
  AND2_X1 U6053 ( .A1(n7972), .A2(n4762), .ZN(n4533) );
  NOR2_X1 U6054 ( .A1(n9877), .A2(n9890), .ZN(n4534) );
  INV_X1 U6055 ( .A(n4710), .ZN(n5374) );
  NAND2_X1 U6056 ( .A1(n4693), .A2(n5805), .ZN(n4710) );
  AND2_X1 U6057 ( .A1(n5545), .A2(SI_12_), .ZN(n4535) );
  NAND2_X1 U6058 ( .A1(n9293), .A2(n9292), .ZN(n4536) );
  INV_X1 U6059 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5253) );
  NOR2_X1 U6060 ( .A1(n4790), .A2(n4792), .ZN(n4537) );
  NAND2_X1 U6061 ( .A1(n4507), .A2(n4823), .ZN(n4822) );
  NAND2_X1 U6062 ( .A1(n7681), .A2(n7676), .ZN(n4538) );
  NAND2_X1 U6063 ( .A1(n7680), .A2(n7679), .ZN(n4539) );
  NAND2_X1 U6064 ( .A1(n8550), .A2(n8662), .ZN(n4540) );
  OR2_X1 U6065 ( .A1(n4934), .A2(n4518), .ZN(n4541) );
  INV_X1 U6066 ( .A(n4930), .ZN(n4929) );
  NAND2_X1 U6067 ( .A1(n4933), .A2(n9785), .ZN(n4930) );
  NAND2_X1 U6068 ( .A1(n9554), .A2(n9403), .ZN(n4542) );
  AND2_X1 U6069 ( .A1(n7955), .A2(n7766), .ZN(n8668) );
  AND2_X1 U6070 ( .A1(n8247), .A2(n8416), .ZN(n4543) );
  NAND2_X1 U6071 ( .A1(n4541), .A2(n4933), .ZN(n4928) );
  OR2_X1 U6072 ( .A1(n5810), .A2(n7993), .ZN(n4544) );
  NAND2_X1 U6073 ( .A1(n5286), .A2(n5285), .ZN(n5289) );
  OR2_X1 U6074 ( .A1(n8266), .A2(n8267), .ZN(n6258) );
  NAND2_X1 U6075 ( .A1(n4508), .A2(n4681), .ZN(n4680) );
  NAND2_X1 U6076 ( .A1(n9470), .A2(n9469), .ZN(n9596) );
  INV_X1 U6077 ( .A(n9596), .ZN(n4661) );
  NAND2_X1 U6078 ( .A1(n5292), .A2(n5291), .ZN(n7595) );
  AND2_X1 U6079 ( .A1(n8553), .A2(n8633), .ZN(n4545) );
  AND2_X1 U6080 ( .A1(n5048), .A2(n4980), .ZN(n4546) );
  AND2_X1 U6081 ( .A1(n4932), .A2(n4931), .ZN(n4547) );
  NOR2_X1 U6082 ( .A1(n8600), .A2(n7962), .ZN(n4548) );
  AND2_X1 U6083 ( .A1(n7724), .A2(n7356), .ZN(n7932) );
  INV_X1 U6084 ( .A(n7932), .ZN(n4699) );
  INV_X1 U6085 ( .A(n10155), .ZN(n9962) );
  AND2_X1 U6086 ( .A1(n8059), .A2(n8058), .ZN(n10155) );
  AND2_X1 U6087 ( .A1(n6844), .A2(n9412), .ZN(n4549) );
  AND2_X1 U6088 ( .A1(n7947), .A2(n7945), .ZN(n4550) );
  AND2_X1 U6089 ( .A1(n5013), .A2(n5260), .ZN(n4551) );
  AND2_X1 U6090 ( .A1(n4540), .A2(n4702), .ZN(n4552) );
  OR2_X1 U6091 ( .A1(n9157), .A2(n8566), .ZN(n4553) );
  AND2_X1 U6092 ( .A1(n7901), .A2(n4977), .ZN(n4554) );
  AND2_X1 U6093 ( .A1(n5757), .A2(n5636), .ZN(n4555) );
  OR2_X1 U6094 ( .A1(n4777), .A2(n4776), .ZN(n4556) );
  INV_X1 U6095 ( .A(n4936), .ZN(n4731) );
  NAND2_X1 U6096 ( .A1(n8561), .A2(n8596), .ZN(n4936) );
  INV_X1 U6097 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n4697) );
  AND2_X1 U6098 ( .A1(n6968), .A2(n6967), .ZN(n7121) );
  NAND2_X1 U6099 ( .A1(n6992), .A2(n6991), .ZN(n7034) );
  NAND2_X1 U6100 ( .A1(n4972), .A2(n4970), .ZN(n8115) );
  NAND2_X1 U6101 ( .A1(n6568), .A2(n7680), .ZN(n6747) );
  NAND2_X1 U6102 ( .A1(n8185), .A2(n8184), .ZN(n10058) );
  INV_X1 U6103 ( .A(n10058), .ZN(n4864) );
  AND2_X1 U6104 ( .A1(n9803), .A2(n9484), .ZN(n9836) );
  AND2_X1 U6105 ( .A1(n6207), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4557) );
  INV_X1 U6106 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4850) );
  XNOR2_X1 U6107 ( .A(n7399), .B(n7404), .ZN(n7398) );
  XOR2_X1 U6108 ( .A(n8011), .B(n4495), .Z(n4558) );
  INV_X1 U6109 ( .A(n9382), .ZN(n4677) );
  INV_X1 U6110 ( .A(n9543), .ZN(n4684) );
  NAND2_X1 U6111 ( .A1(n8202), .A2(n8201), .ZN(n9846) );
  INV_X1 U6112 ( .A(n9846), .ZN(n4863) );
  INV_X1 U6113 ( .A(n9550), .ZN(n4642) );
  INV_X1 U6114 ( .A(n9779), .ZN(n9998) );
  AND4_X1 U6115 ( .A1(n7218), .A2(n7217), .A3(n7216), .A4(n7215), .ZN(n9779)
         );
  AND2_X1 U6116 ( .A1(n4738), .A2(n4739), .ZN(n4559) );
  NAND2_X1 U6117 ( .A1(n10018), .A2(n4858), .ZN(n4860) );
  AND2_X1 U6118 ( .A1(n7087), .A2(n4847), .ZN(n4560) );
  AND2_X1 U6119 ( .A1(n9993), .A2(n10014), .ZN(n4561) );
  NOR2_X1 U6120 ( .A1(n10133), .A2(n9845), .ZN(n4562) );
  NAND2_X1 U6121 ( .A1(n9330), .A2(n8041), .ZN(n9248) );
  AND2_X1 U6122 ( .A1(n6891), .A2(n6717), .ZN(n4563) );
  INV_X1 U6123 ( .A(n8293), .ZN(n4984) );
  NOR2_X1 U6124 ( .A1(n6821), .A2(n7031), .ZN(n4862) );
  NAND2_X1 U6125 ( .A1(n5171), .A2(n5289), .ZN(n5176) );
  INV_X2 U6126 ( .A(n10278), .ZN(n10280) );
  INV_X1 U6127 ( .A(n7228), .ZN(n4873) );
  AND2_X1 U6128 ( .A1(n9712), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4564) );
  NAND2_X1 U6129 ( .A1(n5045), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5058) );
  OR2_X1 U6130 ( .A1(n6706), .A2(n9604), .ZN(n10266) );
  INV_X1 U6131 ( .A(n10266), .ZN(n10072) );
  NAND2_X1 U6132 ( .A1(n5284), .A2(n9617), .ZN(n10009) );
  INV_X1 U6133 ( .A(n8477), .ZN(n8493) );
  AND3_X1 U6134 ( .A1(n5527), .A2(n6275), .A3(n5534), .ZN(n9342) );
  OR2_X1 U6135 ( .A1(n8458), .A2(n9090), .ZN(n4565) );
  OR2_X1 U6136 ( .A1(n8458), .A2(n8457), .ZN(n4566) );
  NOR2_X1 U6137 ( .A1(n8268), .A2(n6258), .ZN(n4567) );
  AND2_X1 U6138 ( .A1(n4620), .A2(n9760), .ZN(n4568) );
  NAND3_X1 U6139 ( .A1(n5604), .A2(n5603), .A3(n5602), .ZN(n5735) );
  XNOR2_X1 U6140 ( .A(n5779), .B(P2_IR_REG_19__SCAN_IN), .ZN(n7981) );
  NAND3_X1 U6141 ( .A1(n5258), .A2(n4574), .A3(n4573), .ZN(n9621) );
  INV_X1 U6142 ( .A(n7973), .ZN(n4760) );
  NAND2_X1 U6143 ( .A1(n4571), .A2(n4865), .ZN(n4570) );
  NAND2_X1 U6144 ( .A1(n6555), .A2(n4867), .ZN(n4571) );
  NAND2_X1 U6145 ( .A1(n6554), .A2(n6553), .ZN(n6555) );
  NOR2_X1 U6146 ( .A1(n5020), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n4572) );
  INV_X1 U6147 ( .A(n4578), .ZN(n9351) );
  NAND2_X1 U6148 ( .A1(n8015), .A2(n4575), .ZN(n9270) );
  NAND2_X1 U6149 ( .A1(n4576), .A2(n9352), .ZN(n4575) );
  NAND2_X1 U6150 ( .A1(n4578), .A2(n4577), .ZN(n4576) );
  INV_X1 U6151 ( .A(n9353), .ZN(n4577) );
  NAND2_X1 U6152 ( .A1(n9235), .A2(n9237), .ZN(n4579) );
  NAND2_X2 U6153 ( .A1(n4581), .A2(n8084), .ZN(n9312) );
  OAI21_X2 U6154 ( .B1(n4907), .B2(n4584), .A(n4582), .ZN(n9330) );
  INV_X1 U6155 ( .A(n9280), .ZN(n4584) );
  NAND3_X1 U6156 ( .A1(n4586), .A2(n4588), .A3(n4585), .ZN(n4587) );
  NAND2_X1 U6157 ( .A1(n6258), .A2(n4900), .ZN(n4588) );
  NOR2_X1 U6158 ( .A1(n5718), .A2(n6261), .ZN(n4589) );
  INV_X1 U6159 ( .A(n5719), .ZN(n4590) );
  NAND3_X1 U6160 ( .A1(n4852), .A2(n5004), .A3(n5007), .ZN(n5233) );
  NAND2_X1 U6161 ( .A1(n9792), .A2(n4913), .ZN(n9827) );
  INV_X1 U6162 ( .A(n9835), .ZN(n4602) );
  OAI21_X1 U6163 ( .B1(n6220), .B2(n4606), .A(n6427), .ZN(n4605) );
  OAI21_X2 U6164 ( .B1(n5910), .B2(n4606), .A(n4604), .ZN(n6430) );
  AND2_X1 U6165 ( .A1(n5168), .A2(n5167), .ZN(n5285) );
  NOR2_X1 U6166 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(n5122), .ZN(n4609) );
  INV_X1 U6167 ( .A(n5122), .ZN(n4610) );
  NAND2_X1 U6168 ( .A1(n10005), .A2(n9780), .ZN(n4612) );
  AOI21_X2 U6169 ( .B1(n9934), .B2(n5000), .A(n4615), .ZN(n4614) );
  NAND3_X1 U6170 ( .A1(n4621), .A2(n4568), .A3(n4618), .ZN(P1_U3262) );
  INV_X1 U6171 ( .A(n5112), .ZN(n4852) );
  INV_X1 U6172 ( .A(n4851), .ZN(n4631) );
  NAND2_X1 U6173 ( .A1(n5289), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5290) );
  XNOR2_X1 U6174 ( .A(n4633), .B(n4632), .ZN(n6806) );
  OR2_X1 U6175 ( .A1(n9402), .A2(n4637), .ZN(n4634) );
  OAI211_X1 U6176 ( .C1(n9394), .C2(n4640), .A(n4634), .B(n4635), .ZN(n9424)
         );
  INV_X1 U6177 ( .A(n9471), .ZN(n4643) );
  AND2_X1 U6178 ( .A1(n9401), .A2(n9548), .ZN(n4644) );
  OR2_X1 U6179 ( .A1(n9481), .A2(n4654), .ZN(n4649) );
  NAND2_X1 U6180 ( .A1(n4649), .A2(n4651), .ZN(n9620) );
  AND2_X1 U6181 ( .A1(n9766), .A2(n9627), .ZN(n4664) );
  NAND2_X1 U6182 ( .A1(n4689), .A2(n4687), .ZN(n9387) );
  NOR2_X1 U6183 ( .A1(n4677), .A2(n9471), .ZN(n4688) );
  NAND2_X1 U6184 ( .A1(n4690), .A2(n9471), .ZN(n4689) );
  NAND2_X1 U6185 ( .A1(n6003), .A2(n6004), .ZN(n6146) );
  OAI22_X1 U6186 ( .A1(n6001), .A2(n6580), .B1(n6002), .B2(n6573), .ZN(n6003)
         );
  NAND2_X1 U6187 ( .A1(n7272), .A2(n7370), .ZN(n4700) );
  NAND2_X1 U6188 ( .A1(n4701), .A2(n4552), .ZN(n7957) );
  INV_X2 U6189 ( .A(n5810), .ZN(n7736) );
  MUX2_X1 U6190 ( .A(n5805), .B(n9223), .S(n5810), .Z(n5995) );
  NAND3_X1 U6191 ( .A1(n5811), .A2(n5812), .A3(n4544), .ZN(n6355) );
  NAND2_X1 U6192 ( .A1(n7902), .A2(n5810), .ZN(n8778) );
  NAND3_X1 U6193 ( .A1(n4704), .A2(n7701), .A3(n6750), .ZN(n7068) );
  NOR2_X2 U6194 ( .A1(n4802), .A2(n4803), .ZN(n5074) );
  OR2_X2 U6195 ( .A1(n8569), .A2(n4705), .ZN(n8782) );
  NAND3_X1 U6196 ( .A1(n8736), .A2(n5001), .A3(n4714), .ZN(n4705) );
  NAND2_X1 U6197 ( .A1(n4710), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5376) );
  NAND2_X1 U6198 ( .A1(n4713), .A2(n8706), .ZN(n4714) );
  XNOR2_X1 U6199 ( .A(n8563), .B(n4716), .ZN(n4713) );
  NAND2_X1 U6200 ( .A1(n8782), .A2(n10364), .ZN(n8785) );
  NAND2_X1 U6201 ( .A1(n4717), .A2(n5109), .ZN(n4718) );
  INV_X1 U6202 ( .A(n5105), .ZN(n4717) );
  NAND3_X1 U6203 ( .A1(n4719), .A2(n4718), .A3(n5115), .ZN(n5120) );
  NAND3_X1 U6204 ( .A1(n5109), .A2(n5097), .A3(n5098), .ZN(n4719) );
  NAND2_X1 U6205 ( .A1(n5098), .A2(n5097), .ZN(n5106) );
  NAND2_X1 U6206 ( .A1(n4720), .A2(n5109), .ZN(n5116) );
  NAND2_X1 U6207 ( .A1(n5106), .A2(n5105), .ZN(n4720) );
  INV_X1 U6208 ( .A(n4721), .ZN(n8541) );
  INV_X1 U6209 ( .A(n8587), .ZN(n4728) );
  NAND2_X1 U6210 ( .A1(n4728), .A2(n4937), .ZN(n4730) );
  NAND2_X1 U6211 ( .A1(n4730), .A2(n4729), .ZN(n4935) );
  NAND2_X1 U6212 ( .A1(n8718), .A2(n4512), .ZN(n4738) );
  XNOR2_X2 U6213 ( .A(n8428), .B(n6355), .ZN(n7914) );
  XNOR2_X1 U6214 ( .A(n5092), .B(SI_1_), .ZN(n5089) );
  NAND2_X1 U6215 ( .A1(n4755), .A2(n5196), .ZN(n5217) );
  NAND2_X1 U6216 ( .A1(n8620), .A2(n8556), .ZN(n8594) );
  NAND2_X1 U6217 ( .A1(n4935), .A2(n4553), .ZN(n8563) );
  NAND2_X1 U6218 ( .A1(n5480), .A2(n5479), .ZN(n4747) );
  NAND2_X1 U6219 ( .A1(n5194), .A2(n4750), .ZN(n4749) );
  NAND2_X1 U6220 ( .A1(n5194), .A2(n5193), .ZN(n4755) );
  OAI21_X1 U6221 ( .B1(n5194), .B2(n4752), .A(n4750), .ZN(n5229) );
  AOI21_X1 U6222 ( .B1(n4750), .B2(n4752), .A(n5222), .ZN(n4748) );
  NAND2_X1 U6223 ( .A1(n7946), .A2(n4550), .ZN(n8715) );
  NAND2_X1 U6224 ( .A1(n7957), .A2(n4756), .ZN(n8606) );
  NAND2_X1 U6225 ( .A1(n4767), .A2(n4765), .ZN(n7782) );
  NAND2_X1 U6226 ( .A1(n7723), .A2(n4768), .ZN(n4767) );
  INV_X1 U6227 ( .A(n7729), .ZN(n4778) );
  INV_X1 U6228 ( .A(n7725), .ZN(n4780) );
  INV_X1 U6229 ( .A(n4786), .ZN(n7716) );
  NAND2_X1 U6230 ( .A1(n4798), .A2(n7857), .ZN(n7889) );
  NAND2_X1 U6231 ( .A1(n4799), .A2(n5002), .ZN(n4798) );
  NAND2_X1 U6232 ( .A1(n4800), .A2(n8603), .ZN(n4799) );
  INV_X1 U6233 ( .A(n4990), .ZN(n4801) );
  NAND3_X1 U6234 ( .A1(n4969), .A2(n4804), .A3(n4992), .ZN(n4802) );
  NAND2_X1 U6235 ( .A1(n4990), .A2(n4546), .ZN(n4803) );
  NAND3_X1 U6236 ( .A1(n4807), .A2(n4805), .A3(n7688), .ZN(n7700) );
  NAND2_X2 U6237 ( .A1(n9218), .A2(n7593), .ZN(n7841) );
  NAND2_X1 U6238 ( .A1(n4814), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5797) );
  AND2_X1 U6239 ( .A1(n5074), .A2(n4816), .ZN(n5315) );
  NAND2_X1 U6240 ( .A1(n5074), .A2(n4815), .ZN(n9214) );
  NAND2_X1 U6241 ( .A1(n5147), .A2(n5146), .ZN(n4817) );
  INV_X1 U6242 ( .A(n9969), .ZN(n4825) );
  NAND2_X1 U6243 ( .A1(n4821), .A2(n9969), .ZN(n4820) );
  INV_X1 U6244 ( .A(n4822), .ZN(n4821) );
  NAND2_X1 U6245 ( .A1(n9581), .A2(n4833), .ZN(n4829) );
  NAND2_X1 U6246 ( .A1(n4829), .A2(n4830), .ZN(n9995) );
  INV_X1 U6247 ( .A(n6996), .ZN(n4837) );
  NAND2_X1 U6248 ( .A1(n7002), .A2(n7113), .ZN(n6639) );
  NAND2_X1 U6249 ( .A1(n6843), .A2(n4549), .ZN(n4845) );
  NAND4_X1 U6250 ( .A1(n4993), .A2(n4912), .A3(n5017), .A4(n4911), .ZN(n4851)
         );
  NAND2_X1 U6251 ( .A1(n6802), .A2(n4853), .ZN(n5912) );
  INV_X1 U6252 ( .A(n10032), .ZN(n4855) );
  INV_X1 U6253 ( .A(n4860), .ZN(n9961) );
  AND2_X2 U6254 ( .A1(n7338), .A2(n9247), .ZN(n7339) );
  NOR2_X2 U6255 ( .A1(n6855), .A2(n7422), .ZN(n7338) );
  NAND2_X1 U6256 ( .A1(n4870), .A2(n5013), .ZN(n5259) );
  NAND2_X1 U6257 ( .A1(n4870), .A2(n4551), .ZN(n5157) );
  OAI21_X1 U6258 ( .B1(n7230), .B2(n4874), .A(n4871), .ZN(n8012) );
  OAI21_X2 U6259 ( .B1(n7413), .B2(n4879), .A(n4875), .ZN(n9235) );
  NAND2_X1 U6260 ( .A1(n7411), .A2(n7410), .ZN(n4883) );
  NAND2_X1 U6261 ( .A1(n8163), .A2(n8166), .ZN(n4885) );
  OAI21_X1 U6262 ( .B1(n8163), .B2(n4888), .A(n4886), .ZN(n9226) );
  NAND2_X1 U6263 ( .A1(n9293), .A2(n8166), .ZN(n9262) );
  OR2_X1 U6264 ( .A1(n8163), .A2(n8162), .ZN(n9293) );
  NAND2_X1 U6265 ( .A1(n9225), .A2(n4892), .ZN(n4891) );
  OAI211_X1 U6266 ( .C1(n9225), .C2(n4893), .A(n4891), .B(n8240), .ZN(P1_U3220) );
  NAND2_X1 U6267 ( .A1(n9270), .A2(n4905), .ZN(n4903) );
  OR2_X1 U6268 ( .A1(n9270), .A2(n8022), .ZN(n4907) );
  NAND2_X1 U6269 ( .A1(n9792), .A2(n9791), .ZN(n9825) );
  INV_X1 U6270 ( .A(n7077), .ZN(n4921) );
  OAI21_X1 U6271 ( .B1(n9920), .B2(n4925), .A(n4923), .ZN(n9872) );
  NAND2_X1 U6272 ( .A1(n5983), .A2(n4943), .ZN(n4942) );
  NAND2_X1 U6273 ( .A1(n4942), .A2(n4946), .ZN(n6540) );
  OR2_X1 U6274 ( .A1(n5983), .A2(n5982), .ZN(n4949) );
  NAND2_X1 U6275 ( .A1(n4953), .A2(n4555), .ZN(n5962) );
  NAND2_X1 U6276 ( .A1(n5231), .A2(n5230), .ZN(n5335) );
  NAND2_X1 U6277 ( .A1(n6716), .A2(n6715), .ZN(n4954) );
  NAND2_X1 U6278 ( .A1(n4954), .A2(n6717), .ZN(n6890) );
  NAND2_X1 U6279 ( .A1(n4954), .A2(n4563), .ZN(n6895) );
  NAND3_X1 U6280 ( .A1(n4956), .A2(P1_DATAO_REG_1__SCAN_IN), .A3(n4955), .ZN(
        n5082) );
  NAND3_X1 U6281 ( .A1(n8631), .A2(n8621), .A3(n8619), .ZN(n8620) );
  OAI21_X2 U6282 ( .B1(n8301), .B2(n8662), .A(n4964), .ZN(n8349) );
  OAI21_X2 U6283 ( .B1(n8245), .B2(n4961), .A(n4959), .ZN(n4965) );
  NAND2_X1 U6284 ( .A1(n4965), .A2(n4509), .ZN(n4964) );
  NAND2_X1 U6285 ( .A1(n4514), .A2(n4975), .ZN(n10300) );
  NAND2_X1 U6286 ( .A1(n5810), .A2(n4554), .ZN(n4976) );
  INV_X1 U6287 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4977) );
  NAND2_X1 U6288 ( .A1(n6232), .A2(n6231), .ZN(n6767) );
  NAND2_X1 U6289 ( .A1(n5049), .A2(n5048), .ZN(n5050) );
  NAND2_X1 U6290 ( .A1(n8116), .A2(n4981), .ZN(n4983) );
  NAND2_X1 U6291 ( .A1(n6968), .A2(n4987), .ZN(n7128) );
  INV_X1 U6292 ( .A(n6733), .ZN(n6735) );
  NAND2_X1 U6293 ( .A1(n6469), .A2(n6468), .ZN(n6467) );
  NAND2_X1 U6294 ( .A1(n5736), .A2(n5735), .ZN(n9535) );
  INV_X1 U6295 ( .A(n5735), .ZN(n5737) );
  OAI21_X1 U6296 ( .B1(n8733), .B2(n10336), .A(n8568), .ZN(n8569) );
  OR2_X1 U6297 ( .A1(n8396), .A2(n8395), .ZN(n8397) );
  NOR2_X2 U6298 ( .A1(n9783), .A2(n9782), .ZN(n9934) );
  XNOR2_X1 U6299 ( .A(n5868), .B(n6033), .ZN(n5807) );
  NAND2_X1 U6300 ( .A1(n8281), .A2(n8280), .ZN(n8279) );
  NAND2_X2 U6301 ( .A1(n5820), .A2(n8512), .ZN(n5810) );
  OAI21_X1 U6302 ( .B1(n10159), .B2(n9956), .A(n9974), .ZN(n9781) );
  INV_X1 U6303 ( .A(n7625), .ZN(n5293) );
  NAND2_X1 U6304 ( .A1(n5063), .A2(n5062), .ZN(n4988) );
  AND2_X1 U6305 ( .A1(n4491), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n4989) );
  OR2_X1 U6306 ( .A1(n5255), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4994) );
  AND2_X1 U6307 ( .A1(n5011), .A2(n5010), .ZN(n4995) );
  AND2_X1 U6308 ( .A1(n5708), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4996) );
  INV_X1 U6309 ( .A(n9630), .ZN(n9361) );
  AND2_X1 U6310 ( .A1(n9473), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n4997) );
  NAND2_X1 U6311 ( .A1(n10181), .A2(n5818), .ZN(n8390) );
  NAND2_X2 U6312 ( .A1(n6180), .A2(n10181), .ZN(n8724) );
  NAND2_X1 U6313 ( .A1(n5254), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4999) );
  OR2_X1 U6314 ( .A1(n10151), .A2(n9957), .ZN(n5000) );
  INV_X1 U6315 ( .A(n8712), .ZN(n7947) );
  OR2_X1 U6316 ( .A1(n8735), .A2(n10352), .ZN(n5001) );
  AND2_X1 U6317 ( .A1(n8586), .A2(n7846), .ZN(n5002) );
  AND2_X1 U6318 ( .A1(n8254), .A2(n8253), .ZN(n5003) );
  NAND2_X2 U6319 ( .A1(n6277), .A2(n9980), .ZN(n10028) );
  AND2_X1 U6320 ( .A1(n8668), .A2(n7953), .ZN(n7779) );
  NAND2_X1 U6321 ( .A1(n7787), .A2(n7892), .ZN(n7788) );
  NOR2_X1 U6322 ( .A1(n8562), .A2(n7856), .ZN(n7857) );
  INV_X1 U6323 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5037) );
  INV_X1 U6324 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5039) );
  INV_X1 U6325 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5008) );
  NAND2_X1 U6326 ( .A1(n5161), .A2(n5160), .ZN(n5162) );
  INV_X1 U6327 ( .A(n7975), .ZN(n7907) );
  NAND2_X1 U6328 ( .A1(n6988), .A2(n6990), .ZN(n6991) );
  OR2_X1 U6329 ( .A1(n7322), .A2(n7321), .ZN(n7016) );
  INV_X1 U6330 ( .A(n9856), .ZN(n9801) );
  INV_X1 U6331 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9085) );
  INV_X1 U6332 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8996) );
  INV_X1 U6333 ( .A(n5761), .ZN(n5772) );
  NAND2_X1 U6334 ( .A1(n6547), .A2(n8523), .ZN(n5831) );
  NOR2_X1 U6335 ( .A1(n5064), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5066) );
  AND2_X1 U6336 ( .A1(n6260), .A2(n6259), .ZN(n6261) );
  AND2_X1 U6337 ( .A1(n7017), .A2(n7016), .ZN(n7018) );
  INV_X1 U6338 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8833) );
  OR2_X1 U6339 ( .A1(n6669), .A2(n6668), .ZN(n6847) );
  INV_X1 U6340 ( .A(SI_26_), .ZN(n7191) );
  INV_X1 U6341 ( .A(SI_24_), .ZN(n9065) );
  INV_X1 U6342 ( .A(SI_20_), .ZN(n6543) );
  INV_X1 U6343 ( .A(SI_17_), .ZN(n5984) );
  INV_X1 U6344 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5318) );
  NOR2_X1 U6345 ( .A1(n7944), .A2(n7977), .ZN(n7908) );
  INV_X1 U6346 ( .A(n6581), .ZN(n7862) );
  INV_X1 U6347 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7869) );
  INV_X1 U6348 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7473) );
  INV_X1 U6349 ( .A(n8567), .ZN(n8568) );
  OR2_X1 U6350 ( .A1(n7893), .A2(n5831), .ZN(n6177) );
  AND2_X1 U6351 ( .A1(n9227), .A2(n9228), .ZN(n8214) );
  NAND2_X1 U6352 ( .A1(n7322), .A2(n7321), .ZN(n7019) );
  NOR2_X1 U6353 ( .A1(n9265), .A2(n8170), .ZN(n8186) );
  NAND2_X1 U6354 ( .A1(n8101), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8170) );
  NOR2_X1 U6355 ( .A1(n6847), .A2(n6846), .ZN(n7081) );
  AND2_X1 U6356 ( .A1(n5707), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5294) );
  OAI22_X1 U6357 ( .A1(n9845), .A2(n10011), .B1(n9807), .B2(n9806), .ZN(n9808)
         );
  NAND2_X1 U6358 ( .A1(n10020), .A2(n9998), .ZN(n9780) );
  INV_X1 U6359 ( .A(n9980), .ZN(n10022) );
  NAND2_X1 U6360 ( .A1(n5739), .A2(n6339), .ZN(n9534) );
  OR2_X1 U6361 ( .A1(n7190), .A2(n7189), .ZN(n7204) );
  AND2_X1 U6362 ( .A1(n6579), .A2(n5318), .ZN(n5349) );
  INV_X1 U6363 ( .A(n8623), .ZN(n8558) );
  INV_X1 U6364 ( .A(n8704), .ZN(n8546) );
  INV_X1 U6365 ( .A(n8662), .ZN(n8549) );
  INV_X1 U6366 ( .A(n8639), .ZN(n8595) );
  INV_X2 U6367 ( .A(n7288), .ZN(n7861) );
  INV_X1 U6368 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5312) );
  AND2_X1 U6369 ( .A1(n5368), .A2(n7385), .ZN(n5373) );
  NAND2_X1 U6370 ( .A1(n7474), .A2(n7473), .ZN(n7554) );
  INV_X1 U6371 ( .A(n7928), .ZN(n6734) );
  INV_X1 U6372 ( .A(n5872), .ZN(n5873) );
  INV_X1 U6373 ( .A(n8709), .ZN(n10181) );
  OR2_X1 U6374 ( .A1(n7893), .A2(n5832), .ZN(n5888) );
  OR2_X1 U6375 ( .A1(n10352), .A2(n5866), .ZN(n5883) );
  INV_X1 U6376 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8783) );
  OR2_X1 U6377 ( .A1(n5704), .A2(n5703), .ZN(n5706) );
  INV_X1 U6378 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9256) );
  INV_X1 U6379 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6299) );
  INV_X1 U6380 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9313) );
  AND2_X1 U6381 ( .A1(n5706), .A2(n5705), .ZN(n9320) );
  OR2_X1 U6382 ( .A1(n5628), .A2(n10013), .ZN(n9345) );
  OR2_X1 U6383 ( .A1(n5628), .A2(n10011), .ZN(n9360) );
  NOR2_X1 U6384 ( .A1(n8088), .A2(n9313), .ZN(n8089) );
  AND2_X1 U6385 ( .A1(n8046), .A2(n7996), .ZN(n8060) );
  INV_X1 U6386 ( .A(n9914), .ZN(n9940) );
  AND2_X1 U6387 ( .A1(n9561), .A2(n9557), .ZN(n9505) );
  NAND2_X1 U6388 ( .A1(n6756), .A2(n9500), .ZN(n6755) );
  OR2_X1 U6389 ( .A1(n5280), .A2(n5514), .ZN(n5301) );
  NAND2_X1 U6390 ( .A1(n6316), .A2(n6315), .ZN(n6448) );
  INV_X1 U6391 ( .A(n10009), .ZN(n9938) );
  NAND2_X1 U6392 ( .A1(n7384), .A2(n7383), .ZN(n7588) );
  AND2_X1 U6393 ( .A1(n7310), .A2(n6984), .ZN(n7308) );
  AND2_X1 U6394 ( .A1(n6717), .A2(n6546), .ZN(n6715) );
  AND2_X1 U6395 ( .A1(n6060), .A2(n5987), .ZN(n6058) );
  INV_X1 U6396 ( .A(n5222), .ZN(n5228) );
  INV_X1 U6397 ( .A(n8382), .ZN(n8402) );
  INV_X1 U6398 ( .A(n8394), .ZN(n8302) );
  AND2_X1 U6399 ( .A1(n7636), .A2(n7635), .ZN(n8416) );
  OR2_X1 U6400 ( .A1(n7841), .A2(n5822), .ZN(n5828) );
  NAND2_X1 U6401 ( .A1(n7903), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5800) );
  INV_X1 U6402 ( .A(n8522), .ZN(n8448) );
  INV_X1 U6403 ( .A(n8529), .ZN(n8442) );
  INV_X1 U6404 ( .A(n8517), .ZN(n8464) );
  AND2_X1 U6405 ( .A1(n5373), .A2(n5383), .ZN(n8526) );
  OR2_X1 U6406 ( .A1(n10352), .A2(n6185), .ZN(n10183) );
  NOR2_X2 U6407 ( .A1(n7893), .A2(n5873), .ZN(n8703) );
  INV_X1 U6408 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9090) );
  AND2_X1 U6409 ( .A1(n5888), .A2(n5887), .ZN(n6174) );
  AND2_X1 U6410 ( .A1(n7563), .A2(n7562), .ZN(n7570) );
  NAND2_X1 U6411 ( .A1(n10336), .A2(n10344), .ZN(n10358) );
  INV_X1 U6412 ( .A(n10352), .ZN(n10363) );
  XNOR2_X1 U6413 ( .A(n5058), .B(n5059), .ZN(n5833) );
  AND2_X1 U6414 ( .A1(n5210), .A2(n5208), .ZN(n6573) );
  INV_X1 U6415 ( .A(n9345), .ZN(n9355) );
  INV_X1 U6416 ( .A(n9314), .ZN(n9357) );
  AND4_X1 U6417 ( .A1(n8225), .A2(n8224), .A3(n8223), .A4(n8222), .ZN(n9845)
         );
  INV_X1 U6418 ( .A(n5720), .ZN(n8172) );
  AND4_X1 U6419 ( .A1(n6656), .A2(n6655), .A3(n6654), .A4(n6653), .ZN(n7327)
         );
  INV_X1 U6420 ( .A(n9751), .ZN(n9756) );
  OR2_X1 U6421 ( .A1(n5429), .A2(n5428), .ZN(n9752) );
  INV_X1 U6422 ( .A(n9752), .ZN(n9740) );
  AND3_X1 U6423 ( .A1(n9979), .A2(n10072), .A3(n9978), .ZN(n10094) );
  INV_X1 U6424 ( .A(n6317), .ZN(n7337) );
  INV_X1 U6425 ( .A(n10011), .ZN(n9997) );
  INV_X1 U6426 ( .A(n6705), .ZN(n9530) );
  INV_X1 U6427 ( .A(n10276), .ZN(n10113) );
  AND2_X1 U6428 ( .A1(n5525), .A2(n5516), .ZN(n10117) );
  AND2_X1 U6429 ( .A1(n9471), .A2(n9577), .ZN(n6916) );
  INV_X1 U6430 ( .A(n5273), .ZN(n10205) );
  AND2_X1 U6431 ( .A1(n5645), .A2(n5846), .ZN(n9712) );
  AND2_X1 U6432 ( .A1(n5238), .A2(n5345), .ZN(n6440) );
  AND2_X2 U6433 ( .A1(n5782), .A2(n5781), .ZN(n8394) );
  INV_X1 U6434 ( .A(n8390), .ZN(n8410) );
  NAND2_X1 U6435 ( .A1(n7832), .A2(n7831), .ZN(n8623) );
  INV_X1 U6436 ( .A(n8720), .ZN(n8690) );
  OR2_X1 U6437 ( .A1(n8485), .A2(n7983), .ZN(n8517) );
  OR2_X1 U6438 ( .A1(n5384), .A2(n5383), .ZN(n8529) );
  OR2_X1 U6439 ( .A1(n6180), .A2(n10183), .ZN(n8610) );
  INV_X1 U6440 ( .A(n8724), .ZN(n10198) );
  NAND2_X1 U6441 ( .A1(n10381), .A2(n10358), .ZN(n8775) );
  INV_X1 U6442 ( .A(n10381), .ZN(n10378) );
  INV_X1 U6443 ( .A(n7969), .ZN(n8781) );
  AND2_X1 U6444 ( .A1(n7549), .A2(n7946), .ZN(n7574) );
  INV_X2 U6445 ( .A(n10366), .ZN(n10364) );
  INV_X1 U6446 ( .A(n5305), .ZN(n5311) );
  NAND2_X1 U6447 ( .A1(n5834), .A2(n5214), .ZN(n5819) );
  INV_X1 U6448 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7823) );
  INV_X1 U6449 ( .A(n7981), .ZN(n8523) );
  INV_X1 U6450 ( .A(n6573), .ZN(n5953) );
  INV_X1 U6451 ( .A(n7048), .ZN(n7594) );
  XNOR2_X1 U6452 ( .A(n5014), .B(n5019), .ZN(n6985) );
  INV_X1 U6453 ( .A(n9342), .ZN(n9365) );
  INV_X1 U6454 ( .A(n9842), .ZN(n9869) );
  INV_X1 U6455 ( .A(n9941), .ZN(n9972) );
  INV_X1 U6456 ( .A(n7420), .ZN(n9632) );
  OR2_X1 U6457 ( .A1(n5429), .A2(n9762), .ZN(n9751) );
  OAI21_X2 U6458 ( .B1(n7337), .B2(n6318), .A(n10028), .ZN(n10030) );
  NAND2_X1 U6459 ( .A1(n10293), .A2(n10117), .ZN(n10108) );
  OR2_X1 U6460 ( .A1(n5692), .A2(n6273), .ZN(n10290) );
  NAND2_X1 U6461 ( .A1(n10280), .A2(n10117), .ZN(n10164) );
  OR2_X1 U6462 ( .A1(n5692), .A2(n10168), .ZN(n10278) );
  INV_X1 U6463 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8114) );
  INV_X1 U6464 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n6797) );
  INV_X1 U6465 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n8877) );
  INV_X1 U6466 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5355) );
  INV_X1 U6467 ( .A(n8485), .ZN(P2_U3893) );
  INV_X2 U6468 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U6469 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5150) );
  NOR2_X1 U6470 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5009) );
  NAND4_X1 U6471 ( .A1(n5018), .A2(n4993), .A3(n5009), .A4(n9084), .ZN(n5977)
         );
  NAND2_X1 U6472 ( .A1(n5012), .A2(n4995), .ZN(n5252) );
  INV_X1 U6473 ( .A(n5020), .ZN(n5256) );
  NAND2_X1 U6474 ( .A1(n5538), .A2(n5168), .ZN(n5028) );
  INV_X1 U6475 ( .A(n5028), .ZN(n5023) );
  INV_X1 U6476 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5022) );
  NAND2_X1 U6477 ( .A1(n5023), .A2(n5022), .ZN(n5025) );
  NAND2_X1 U6478 ( .A1(n5025), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5024) );
  MUX2_X1 U6479 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5024), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n5027) );
  INV_X1 U6480 ( .A(n5025), .ZN(n5026) );
  NAND2_X1 U6481 ( .A1(n5026), .A2(n5160), .ZN(n5030) );
  NAND2_X1 U6482 ( .A1(n5028), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5029) );
  NOR2_X1 U6483 ( .A1(n5519), .A2(P1_U3086), .ZN(n5033) );
  NOR2_X1 U6484 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5036) );
  NAND2_X1 U6485 ( .A1(n5038), .A2(n5037), .ZN(n5061) );
  NOR2_X1 U6486 ( .A1(n5061), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5044) );
  NAND2_X1 U6487 ( .A1(n5689), .A2(n5041), .ZN(n5971) );
  INV_X1 U6488 ( .A(n5971), .ZN(n5063) );
  NOR2_X1 U6489 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5042) );
  INV_X1 U6490 ( .A(n5049), .ZN(n5045) );
  NAND2_X1 U6491 ( .A1(n5050), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5051) );
  MUX2_X1 U6492 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5051), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5052) );
  INV_X1 U6493 ( .A(n5214), .ZN(n5060) );
  INV_X1 U6494 ( .A(n5061), .ZN(n5062) );
  NAND2_X1 U6495 ( .A1(n5066), .A2(n5614), .ZN(n6119) );
  NAND2_X1 U6496 ( .A1(n5777), .A2(n5067), .ZN(n5068) );
  NAND2_X1 U6497 ( .A1(n5070), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5071) );
  NAND2_X1 U6498 ( .A1(n7893), .A2(n5834), .ZN(n5072) );
  NAND2_X1 U6499 ( .A1(n5072), .A2(n5833), .ZN(n5368) );
  INV_X1 U6500 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5073) );
  NAND2_X4 U6501 ( .A1(n5079), .A2(n5078), .ZN(n8512) );
  NAND2_X1 U6502 ( .A1(n5080), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  AND2_X1 U6503 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5084) );
  NAND2_X1 U6504 ( .A1(n5110), .A2(n5084), .ZN(n5276) );
  AND2_X1 U6505 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5086) );
  NAND2_X1 U6506 ( .A1(n5085), .A2(n5086), .ZN(n5803) );
  NAND2_X1 U6507 ( .A1(n5276), .A2(n5803), .ZN(n5090) );
  XNOR2_X1 U6508 ( .A(n5089), .B(n5090), .ZN(n5783) );
  INV_X1 U6509 ( .A(n5783), .ZN(n5132) );
  NAND2_X1 U6510 ( .A1(n5085), .A2(P1_U3086), .ZN(n8278) );
  INV_X1 U6511 ( .A(n8278), .ZN(n10171) );
  NAND2_X1 U6512 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5087) );
  XNOR2_X1 U6513 ( .A(n5087), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9645) );
  AOI22_X1 U6514 ( .A1(n10171), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(n9645), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n5088) );
  OAI21_X1 U6515 ( .B1(n5132), .B2(n10173), .A(n5088), .ZN(P1_U3354) );
  INV_X1 U6516 ( .A(n5089), .ZN(n5091) );
  NAND2_X1 U6517 ( .A1(n5091), .A2(n5090), .ZN(n5094) );
  NAND2_X1 U6518 ( .A1(n5092), .A2(SI_1_), .ZN(n5093) );
  XNOR2_X1 U6519 ( .A(n5095), .B(SI_2_), .ZN(n5697) );
  NAND2_X1 U6520 ( .A1(n5698), .A2(n5697), .ZN(n5098) );
  INV_X1 U6521 ( .A(n5095), .ZN(n5096) );
  NAND2_X1 U6522 ( .A1(n5096), .A2(SI_2_), .ZN(n5097) );
  INV_X1 U6523 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6034) );
  INV_X1 U6524 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n5099) );
  MUX2_X1 U6525 ( .A(n6034), .B(n5099), .S(n5110), .Z(n5107) );
  XNOR2_X1 U6526 ( .A(n5106), .B(n5105), .ZN(n5715) );
  INV_X1 U6527 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5101) );
  NAND2_X1 U6528 ( .A1(n5410), .A2(n5101), .ZN(n5102) );
  NAND2_X1 U6529 ( .A1(n5102), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5103) );
  XNOR2_X1 U6530 ( .A(n5103), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9671) );
  AOI22_X1 U6531 ( .A1(n9671), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n10171), .ZN(n5104) );
  OAI21_X1 U6532 ( .B1(n5715), .B2(n10173), .A(n5104), .ZN(P1_U3352) );
  INV_X1 U6533 ( .A(n5107), .ZN(n5108) );
  NAND2_X1 U6534 ( .A1(n5108), .A2(SI_3_), .ZN(n5109) );
  INV_X1 U6535 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6093) );
  INV_X1 U6536 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n5111) );
  MUX2_X1 U6537 ( .A(n6093), .B(n5111), .S(n5110), .Z(n5117) );
  XNOR2_X1 U6538 ( .A(n5117), .B(SI_4_), .ZN(n5115) );
  XNOR2_X1 U6539 ( .A(n5116), .B(n5115), .ZN(n5898) );
  NAND2_X1 U6540 ( .A1(n5112), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5113) );
  XNOR2_X1 U6541 ( .A(n5113), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9685) );
  AOI22_X1 U6542 ( .A1(n9685), .A2(P1_STATE_REG_SCAN_IN), .B1(n10171), .B2(
        P2_DATAO_REG_4__SCAN_IN), .ZN(n5114) );
  OAI21_X1 U6543 ( .B1(n5898), .B2(n10173), .A(n5114), .ZN(P1_U3351) );
  INV_X1 U6544 ( .A(n5117), .ZN(n5118) );
  NAND2_X1 U6545 ( .A1(n5118), .A2(SI_4_), .ZN(n5119) );
  NAND2_X1 U6546 ( .A1(n5120), .A2(n5119), .ZN(n5137) );
  INV_X1 U6547 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6234) );
  INV_X1 U6548 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n5121) );
  MUX2_X1 U6549 ( .A(n6234), .B(n5121), .S(n7901), .Z(n5138) );
  XNOR2_X1 U6550 ( .A(n5138), .B(SI_5_), .ZN(n5136) );
  XNOR2_X1 U6551 ( .A(n5137), .B(n5136), .ZN(n5909) );
  NAND2_X1 U6552 ( .A1(n5124), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5123) );
  MUX2_X1 U6553 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5123), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5126) );
  NOR2_X1 U6554 ( .A1(n5124), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5142) );
  INV_X1 U6555 ( .A(n5142), .ZN(n5125) );
  AOI22_X1 U6556 ( .A1(n5906), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n10171), .ZN(n5127) );
  OAI21_X1 U6557 ( .B1(n5909), .B2(n10173), .A(n5127), .ZN(P1_U3350) );
  NOR2_X1 U6558 ( .A1(n5085), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9216) );
  INV_X2 U6559 ( .A(n9216), .ZN(n9222) );
  NAND2_X1 U6560 ( .A1(n5085), .A2(P2_U3151), .ZN(n9220) );
  NAND2_X1 U6561 ( .A1(n5129), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5128) );
  MUX2_X1 U6562 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5128), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5130) );
  OR2_X1 U6563 ( .A1(n5129), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n5184) );
  INV_X1 U6564 ( .A(n6035), .ZN(n5576) );
  OAI222_X1 U6565 ( .A1(n9222), .A2(n6034), .B1(n9220), .B2(n5715), .C1(
        P2_U3151), .C2(n5576), .ZN(P2_U3292) );
  NAND2_X1 U6566 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5131) );
  XNOR2_X1 U6567 ( .A(n5131), .B(P2_IR_REG_1__SCAN_IN), .ZN(n5784) );
  INV_X1 U6568 ( .A(n5784), .ZN(n5394) );
  OAI222_X1 U6569 ( .A1(n9222), .A2(n4977), .B1(n9220), .B2(n5132), .C1(
        P2_U3151), .C2(n5394), .ZN(P2_U3294) );
  INV_X1 U6570 ( .A(P2_B_REG_SCAN_IN), .ZN(n8863) );
  XNOR2_X1 U6571 ( .A(n7395), .B(n8863), .ZN(n5133) );
  OAI22_X1 U6572 ( .A1(n5761), .A2(P2_D_REG_1__SCAN_IN), .B1(n7250), .B2(n5134), .ZN(n5877) );
  NAND2_X1 U6573 ( .A1(n5819), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5135) );
  OAI21_X1 U6574 ( .B1(n5877), .B2(n5819), .A(n5135), .ZN(P2_U3377) );
  INV_X1 U6575 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n5144) );
  NAND2_X1 U6576 ( .A1(n5137), .A2(n5136), .ZN(n5141) );
  INV_X1 U6577 ( .A(n5138), .ZN(n5139) );
  NAND2_X1 U6578 ( .A1(n5139), .A2(SI_5_), .ZN(n5140) );
  MUX2_X1 U6579 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7901), .Z(n5148) );
  XNOR2_X1 U6580 ( .A(n5148), .B(SI_6_), .ZN(n5145) );
  XNOR2_X1 U6581 ( .A(n5147), .B(n5145), .ZN(n6194) );
  INV_X1 U6582 ( .A(n6194), .ZN(n5190) );
  OR2_X1 U6583 ( .A1(n5142), .A2(n10169), .ZN(n5143) );
  XNOR2_X1 U6584 ( .A(n5143), .B(n5015), .ZN(n6197) );
  OAI222_X1 U6585 ( .A1(n8278), .A2(n5144), .B1(n10173), .B2(n5190), .C1(
        P1_U3086), .C2(n6197), .ZN(P1_U3349) );
  INV_X1 U6586 ( .A(n5145), .ZN(n5146) );
  NAND2_X1 U6587 ( .A1(n5148), .A2(SI_6_), .ZN(n5149) );
  MUX2_X1 U6588 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7901), .Z(n5195) );
  XNOR2_X1 U6589 ( .A(n5195), .B(SI_7_), .ZN(n5192) );
  AND2_X1 U6590 ( .A1(n4610), .A2(n5150), .ZN(n5201) );
  OR2_X1 U6591 ( .A1(n5201), .A2(n10169), .ZN(n5151) );
  XNOR2_X1 U6592 ( .A(n5151), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6207) );
  AOI22_X1 U6593 ( .A1(n6207), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n10171), .ZN(n5152) );
  OAI21_X1 U6594 ( .B1(n5209), .B2(n10173), .A(n5152), .ZN(P1_U3348) );
  INV_X1 U6595 ( .A(n5519), .ZN(n5522) );
  AOI21_X1 U6596 ( .B1(n6985), .B2(n5522), .A(P1_U3086), .ZN(n5173) );
  NAND2_X1 U6597 ( .A1(n5157), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5159) );
  XNOR2_X1 U6598 ( .A(n5159), .B(n5158), .ZN(n5514) );
  INV_X1 U6599 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5161) );
  INV_X1 U6600 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5160) );
  NAND3_X1 U6601 ( .A1(n5538), .A2(n5168), .A3(n5165), .ZN(n5163) );
  NAND2_X1 U6602 ( .A1(n5538), .A2(n5285), .ZN(n5169) );
  NAND2_X1 U6603 ( .A1(n5169), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5170) );
  AOI21_X1 U6604 ( .B1(n9602), .B2(n6985), .A(n8043), .ZN(n5174) );
  INV_X1 U6605 ( .A(n5174), .ZN(n5172) );
  NAND2_X1 U6606 ( .A1(n5173), .A2(n5172), .ZN(n9761) );
  INV_X1 U6607 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n5180) );
  NAND2_X1 U6608 ( .A1(n5174), .A2(n5173), .ZN(n5429) );
  INV_X1 U6609 ( .A(n5429), .ZN(n9753) );
  INV_X1 U6610 ( .A(n5175), .ZN(n9762) );
  INV_X1 U6611 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6714) );
  AOI21_X1 U6612 ( .B1(n9762), .B2(n6714), .A(n5176), .ZN(n9655) );
  OAI21_X1 U6613 ( .B1(n9762), .B2(P1_REG1_REG_0__SCAN_IN), .A(n9655), .ZN(
        n5177) );
  XNOR2_X1 U6614 ( .A(n5177), .B(P1_IR_REG_0__SCAN_IN), .ZN(n5178) );
  AOI22_X1 U6615 ( .A1(n9753), .A2(n5178), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n5179) );
  OAI21_X1 U6616 ( .B1(n9761), .B2(n5180), .A(n5179), .ZN(P1_U3243) );
  INV_X1 U6617 ( .A(n9220), .ZN(n7048) );
  INV_X1 U6618 ( .A(n5184), .ZN(n5182) );
  INV_X1 U6619 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5181) );
  NAND2_X1 U6620 ( .A1(n5182), .A2(n5181), .ZN(n5186) );
  NAND2_X1 U6621 ( .A1(n5186), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5183) );
  XNOR2_X1 U6622 ( .A(n5183), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6233) );
  INV_X1 U6623 ( .A(n6233), .ZN(n5664) );
  OAI222_X1 U6624 ( .A1(n9222), .A2(n6234), .B1(n7594), .B2(n5909), .C1(
        P2_U3151), .C2(n5664), .ZN(P2_U3290) );
  NAND2_X1 U6625 ( .A1(n5184), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5185) );
  INV_X1 U6626 ( .A(n8447), .ZN(n5565) );
  OAI222_X1 U6627 ( .A1(n9222), .A2(n6093), .B1(n7594), .B2(n5898), .C1(
        P2_U3151), .C2(n5565), .ZN(P2_U3291) );
  INV_X1 U6628 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n5191) );
  INV_X1 U6629 ( .A(n5186), .ZN(n5188) );
  INV_X1 U6630 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5187) );
  NAND2_X1 U6631 ( .A1(n5188), .A2(n5187), .ZN(n5205) );
  NAND2_X1 U6632 ( .A1(n5205), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5189) );
  XNOR2_X1 U6633 ( .A(n5189), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6565) );
  INV_X1 U6634 ( .A(n6565), .ZN(n5952) );
  OAI222_X1 U6635 ( .A1(n9222), .A2(n5191), .B1(n7594), .B2(n5190), .C1(
        P2_U3151), .C2(n5952), .ZN(P2_U3289) );
  INV_X1 U6636 ( .A(n5192), .ZN(n5193) );
  NAND2_X1 U6637 ( .A1(n5195), .A2(SI_7_), .ZN(n5196) );
  INV_X1 U6638 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n5213) );
  INV_X1 U6639 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5327) );
  MUX2_X1 U6640 ( .A(n5213), .B(n5327), .S(n7901), .Z(n5198) );
  INV_X1 U6641 ( .A(SI_8_), .ZN(n5197) );
  NAND2_X1 U6642 ( .A1(n5198), .A2(n5197), .ZN(n5215) );
  INV_X1 U6643 ( .A(n5198), .ZN(n5199) );
  NAND2_X1 U6644 ( .A1(n5199), .A2(SI_8_), .ZN(n5200) );
  NAND2_X1 U6645 ( .A1(n5215), .A2(n5200), .ZN(n5216) );
  XNOR2_X1 U6646 ( .A(n5217), .B(n5216), .ZN(n6569) );
  INV_X1 U6647 ( .A(n6569), .ZN(n5212) );
  NAND2_X1 U6648 ( .A1(n5201), .A2(n5016), .ZN(n5202) );
  NAND2_X1 U6649 ( .A1(n5202), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5203) );
  XNOR2_X1 U6650 ( .A(n5203), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6309) );
  AOI22_X1 U6651 ( .A1(n6309), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n10171), .ZN(n5204) );
  OAI21_X1 U6652 ( .B1(n5212), .B2(n10173), .A(n5204), .ZN(P1_U3347) );
  INV_X1 U6653 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n8994) );
  NAND2_X1 U6654 ( .A1(n5225), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5207) );
  INV_X1 U6655 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5206) );
  NAND2_X1 U6656 ( .A1(n5207), .A2(n5206), .ZN(n5210) );
  OR2_X1 U6657 ( .A1(n5207), .A2(n5206), .ZN(n5208) );
  OAI222_X1 U6658 ( .A1(n9222), .A2(n8994), .B1(n7594), .B2(n5209), .C1(
        P2_U3151), .C2(n5953), .ZN(P2_U3288) );
  INV_X1 U6659 ( .A(n9761), .ZN(n9644) );
  NOR2_X1 U6660 ( .A1(n9644), .A2(P1_U3973), .ZN(P1_U3085) );
  NAND2_X1 U6661 ( .A1(n5210), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5211) );
  XNOR2_X1 U6662 ( .A(n5211), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6570) );
  INV_X1 U6663 ( .A(n6570), .ZN(n6015) );
  OAI222_X1 U6664 ( .A1(n9222), .A2(n5213), .B1(n7594), .B2(n5212), .C1(
        P2_U3151), .C2(n6015), .ZN(P2_U3287) );
  NAND2_X1 U6665 ( .A1(n5885), .A2(n5761), .ZN(n5305) );
  INV_X1 U6666 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5763) );
  AOI22_X1 U6667 ( .A1(n5305), .A2(n5763), .B1(n5214), .B2(n5762), .ZN(
        P2_U3376) );
  INV_X1 U6668 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5227) );
  MUX2_X1 U6669 ( .A(n5227), .B(n5355), .S(n7901), .Z(n5219) );
  INV_X1 U6670 ( .A(SI_9_), .ZN(n5218) );
  NAND2_X1 U6671 ( .A1(n5219), .A2(n5218), .ZN(n5230) );
  INV_X1 U6672 ( .A(n5219), .ZN(n5220) );
  NAND2_X1 U6673 ( .A1(n5220), .A2(SI_9_), .ZN(n5221) );
  NAND2_X1 U6674 ( .A1(n5230), .A2(n5221), .ZN(n5222) );
  INV_X1 U6675 ( .A(n6587), .ZN(n5239) );
  INV_X1 U6676 ( .A(n5223), .ZN(n5224) );
  OAI21_X1 U6677 ( .B1(n5225), .B2(n5224), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5226) );
  XNOR2_X1 U6678 ( .A(n5226), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6588) );
  INV_X1 U6679 ( .A(n6588), .ZN(n6158) );
  OAI222_X1 U6680 ( .A1(n9220), .A2(n5239), .B1(n6158), .B2(P2_U3151), .C1(
        n5227), .C2(n9222), .ZN(P2_U3286) );
  INV_X1 U6681 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5244) );
  INV_X1 U6682 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5232) );
  MUX2_X1 U6683 ( .A(n5244), .B(n5232), .S(n7901), .Z(n5337) );
  XNOR2_X1 U6684 ( .A(n5337), .B(SI_10_), .ZN(n5336) );
  XNOR2_X1 U6685 ( .A(n5335), .B(n5336), .ZN(n6722) );
  INV_X1 U6686 ( .A(n6722), .ZN(n5245) );
  OR2_X1 U6687 ( .A1(n5233), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5345) );
  NAND2_X1 U6688 ( .A1(n5345), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5234) );
  XNOR2_X1 U6689 ( .A(n5234), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6644) );
  AOI22_X1 U6690 ( .A1(n6644), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10171), .ZN(n5235) );
  OAI21_X1 U6691 ( .B1(n5245), .B2(n10173), .A(n5235), .ZN(P1_U3345) );
  NAND2_X1 U6692 ( .A1(n5233), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5237) );
  MUX2_X1 U6693 ( .A(n5237), .B(P1_IR_REG_31__SCAN_IN), .S(n5236), .Z(n5238)
         );
  INV_X1 U6694 ( .A(n6440), .ZN(n5494) );
  OAI222_X1 U6695 ( .A1(n8278), .A2(n5355), .B1(n10173), .B2(n5239), .C1(n5494), .C2(P1_U3086), .ZN(P1_U3346) );
  NAND2_X1 U6696 ( .A1(n5240), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5241) );
  MUX2_X1 U6697 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5241), .S(
        P2_IR_REG_10__SCAN_IN), .Z(n5242) );
  INV_X1 U6698 ( .A(n5242), .ZN(n5243) );
  NOR2_X1 U6699 ( .A1(n5243), .A2(n5065), .ZN(n6723) );
  INV_X1 U6700 ( .A(n6723), .ZN(n6145) );
  OAI222_X1 U6701 ( .A1(n7594), .A2(n5245), .B1(n6145), .B2(P2_U3151), .C1(
        n5244), .C2(n9222), .ZN(P2_U3285) );
  AND2_X1 U6702 ( .A1(n5305), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U6703 ( .A1(n5305), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U6704 ( .A1(n5305), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U6705 ( .A1(n5305), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U6706 ( .A1(n5305), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U6707 ( .A1(n5305), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U6708 ( .A1(n5305), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U6709 ( .A1(n5305), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U6710 ( .A1(n5305), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U6711 ( .A1(n5305), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U6712 ( .A1(n5305), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U6713 ( .A1(n5305), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U6714 ( .A1(n5305), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U6715 ( .A1(n5305), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U6716 ( .A1(n5305), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U6717 ( .A1(n5305), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U6718 ( .A1(n5305), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U6719 ( .A1(n5305), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U6720 ( .A1(n5305), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U6721 ( .A1(n5305), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U6722 ( .A1(n5305), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  NAND2_X1 U6723 ( .A1(n7318), .A2(P1_B_REG_SCAN_IN), .ZN(n5248) );
  MUX2_X1 U6724 ( .A(n5248), .B(P1_B_REG_SCAN_IN), .S(n5272), .Z(n5249) );
  INV_X1 U6725 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10238) );
  INV_X1 U6726 ( .A(n7318), .ZN(n5250) );
  NOR2_X1 U6727 ( .A1(n5247), .A2(n5250), .ZN(n5251) );
  AOI21_X1 U6728 ( .B1(n10205), .B2(n10238), .A(n5251), .ZN(n6274) );
  NOR2_X1 U6729 ( .A1(n10239), .A2(n6274), .ZN(n10237) );
  NAND2_X1 U6730 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n5254) );
  NAND2_X1 U6731 ( .A1(n6062), .A2(n5257), .ZN(n5258) );
  NAND2_X1 U6732 ( .A1(n5259), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5261) );
  NAND2_X1 U6733 ( .A1(n9602), .A2(n5516), .ZN(n5529) );
  NOR2_X1 U6734 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n5265) );
  NOR4_X1 U6735 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5264) );
  NOR4_X1 U6736 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n5263) );
  NOR4_X1 U6737 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n5262) );
  NAND4_X1 U6738 ( .A1(n5265), .A2(n5264), .A3(n5263), .A4(n5262), .ZN(n5271)
         );
  NOR4_X1 U6739 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5269) );
  NOR4_X1 U6740 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5268) );
  NOR4_X1 U6741 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5267) );
  NOR4_X1 U6742 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n5266) );
  NAND4_X1 U6743 ( .A1(n5269), .A2(n5268), .A3(n5267), .A4(n5266), .ZN(n5270)
         );
  OAI21_X1 U6744 ( .B1(n5271), .B2(n5270), .A(n10205), .ZN(n5526) );
  NAND2_X1 U6745 ( .A1(n6916), .A2(n5514), .ZN(n5532) );
  NAND3_X1 U6746 ( .A1(n10237), .A2(n6276), .A3(n5532), .ZN(n5692) );
  INV_X1 U6747 ( .A(n6273), .ZN(n10168) );
  INV_X1 U6748 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5304) );
  NAND2_X1 U6749 ( .A1(n5280), .A2(n5514), .ZN(n6706) );
  INV_X1 U6750 ( .A(SI_0_), .ZN(n5275) );
  INV_X1 U6751 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5274) );
  OAI21_X1 U6752 ( .B1(n5085), .B2(n5275), .A(n5274), .ZN(n5277) );
  AND2_X1 U6753 ( .A1(n5277), .A2(n5276), .ZN(n10175) );
  NAND2_X1 U6754 ( .A1(n5520), .A2(n5516), .ZN(n5282) );
  AND2_X1 U6755 ( .A1(n5282), .A2(n6706), .ZN(n5283) );
  INV_X1 U6756 ( .A(n5516), .ZN(n5535) );
  NAND2_X1 U6757 ( .A1(n9602), .A2(n5535), .ZN(n6707) );
  NAND2_X1 U6758 ( .A1(n5283), .A2(n6707), .ZN(n6317) );
  INV_X1 U6759 ( .A(n6916), .ZN(n10120) );
  OR2_X1 U6760 ( .A1(n5280), .A2(n9621), .ZN(n5284) );
  INV_X1 U6761 ( .A(n5514), .ZN(n9531) );
  NAND2_X1 U6762 ( .A1(n9531), .A2(n9604), .ZN(n9617) );
  NAND2_X1 U6763 ( .A1(n5599), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5297) );
  NAND2_X1 U6764 ( .A1(n5720), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5296) );
  NOR2_X1 U6765 ( .A1(n4991), .A2(n5294), .ZN(n5295) );
  XNOR2_X1 U6766 ( .A(n5594), .B(n9530), .ZN(n9489) );
  OAI21_X1 U6767 ( .B1(n10276), .B2(n10009), .A(n9489), .ZN(n5302) );
  NAND2_X1 U6768 ( .A1(n5707), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5300) );
  NAND2_X1 U6769 ( .A1(n5720), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5299) );
  NAND2_X1 U6770 ( .A1(n5599), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5298) );
  NOR2_X2 U6771 ( .A1(n5301), .A2(n9652), .ZN(n9999) );
  NAND2_X1 U6772 ( .A1(n5593), .A2(n9999), .ZN(n6708) );
  OAI211_X1 U6773 ( .C1(n6706), .C2(n9530), .A(n5302), .B(n6708), .ZN(n10122)
         );
  NAND2_X1 U6774 ( .A1(n10122), .A2(n10280), .ZN(n5303) );
  OAI21_X1 U6775 ( .B1(n10280), .B2(n5304), .A(n5303), .ZN(P1_U3453) );
  INV_X1 U6776 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n8988) );
  NOR2_X1 U6777 ( .A1(n5311), .A2(n8988), .ZN(P2_U3255) );
  INV_X1 U6778 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n9071) );
  NOR2_X1 U6779 ( .A1(n5311), .A2(n9071), .ZN(P2_U3258) );
  INV_X1 U6780 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n8965) );
  NOR2_X1 U6781 ( .A1(n5311), .A2(n8965), .ZN(P2_U3259) );
  INV_X1 U6782 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n5306) );
  NOR2_X1 U6783 ( .A1(n5311), .A2(n5306), .ZN(P2_U3262) );
  INV_X1 U6784 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n8855) );
  NOR2_X1 U6785 ( .A1(n5311), .A2(n8855), .ZN(P2_U3251) );
  INV_X1 U6786 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n5307) );
  NOR2_X1 U6787 ( .A1(n5311), .A2(n5307), .ZN(P2_U3254) );
  INV_X1 U6788 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n5308) );
  NOR2_X1 U6789 ( .A1(n5311), .A2(n5308), .ZN(P2_U3241) );
  INV_X1 U6790 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n5309) );
  NOR2_X1 U6791 ( .A1(n5311), .A2(n5309), .ZN(P2_U3250) );
  INV_X1 U6792 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n5310) );
  NOR2_X1 U6793 ( .A1(n5311), .A2(n5310), .ZN(P2_U3240) );
  INV_X1 U6794 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5314) );
  NOR2_X1 U6795 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6105) );
  INV_X1 U6796 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U6797 ( .A1(n6105), .A2(n6104), .ZN(n6240) );
  NOR2_X1 U6798 ( .A1(n6579), .A2(n5318), .ZN(n5319) );
  OR2_X1 U6799 ( .A1(n5349), .A2(n5319), .ZN(n6974) );
  NAND2_X1 U6800 ( .A1(n7861), .A2(n6974), .ZN(n5326) );
  INV_X1 U6801 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6013) );
  OR2_X1 U6802 ( .A1(n7865), .A2(n6013), .ZN(n5325) );
  INV_X1 U6803 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6012) );
  OR2_X1 U6804 ( .A1(n6581), .A2(n6012), .ZN(n5324) );
  INV_X1 U6805 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5322) );
  OR2_X1 U6806 ( .A1(n7841), .A2(n5322), .ZN(n5323) );
  MUX2_X1 U6807 ( .A(n5327), .B(n7439), .S(P2_U3893), .Z(n5328) );
  INV_X1 U6808 ( .A(n5328), .ZN(P2_U3499) );
  INV_X1 U6809 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6810 ( .A1(n4814), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5333) );
  INV_X1 U6811 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6383) );
  OR2_X1 U6812 ( .A1(n7865), .A2(n6383), .ZN(n5332) );
  NAND2_X1 U6813 ( .A1(n5349), .A2(n5348), .ZN(n6614) );
  OR2_X2 U6814 ( .A1(n6616), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6737) );
  NAND2_X1 U6815 ( .A1(n6616), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5329) );
  AND2_X1 U6816 ( .A1(n6737), .A2(n5329), .ZN(n6751) );
  OR2_X1 U6817 ( .A1(n7288), .A2(n6751), .ZN(n5331) );
  INV_X1 U6818 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6382) );
  OR2_X1 U6819 ( .A1(n6581), .A2(n6382), .ZN(n5330) );
  MUX2_X1 U6820 ( .A(n5339), .B(n7066), .S(P2_U3893), .Z(n5334) );
  INV_X1 U6821 ( .A(n5334), .ZN(P2_U3502) );
  INV_X1 U6822 ( .A(n5337), .ZN(n5338) );
  NAND2_X1 U6823 ( .A1(n5338), .A2(SI_10_), .ZN(n5477) );
  NAND2_X1 U6824 ( .A1(n5480), .A2(n5477), .ZN(n5344) );
  INV_X1 U6825 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5409) );
  MUX2_X1 U6826 ( .A(n5409), .B(n5339), .S(n7901), .Z(n5341) );
  INV_X1 U6827 ( .A(SI_11_), .ZN(n5340) );
  NAND2_X1 U6828 ( .A1(n5341), .A2(n5340), .ZN(n5481) );
  INV_X1 U6829 ( .A(n5341), .ZN(n5342) );
  NAND2_X1 U6830 ( .A1(n5342), .A2(SI_11_), .ZN(n5343) );
  NAND2_X1 U6831 ( .A1(n5481), .A2(n5343), .ZN(n5476) );
  XNOR2_X1 U6832 ( .A(n5344), .B(n5476), .ZN(n6729) );
  INV_X1 U6833 ( .A(n6729), .ZN(n5408) );
  OAI21_X1 U6834 ( .B1(n5345), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5346) );
  XNOR2_X1 U6835 ( .A(n5346), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6648) );
  AOI22_X1 U6836 ( .A1(n6648), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n10171), .ZN(n5347) );
  OAI21_X1 U6837 ( .B1(n5408), .B2(n10173), .A(n5347), .ZN(P1_U3344) );
  NAND2_X1 U6838 ( .A1(n4814), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5354) );
  INV_X1 U6839 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6624) );
  OR2_X1 U6840 ( .A1(n7865), .A2(n6624), .ZN(n5353) );
  OR2_X1 U6841 ( .A1(n5349), .A2(n5348), .ZN(n5350) );
  AND2_X1 U6842 ( .A1(n6614), .A2(n5350), .ZN(n7435) );
  OR2_X1 U6843 ( .A1(n7288), .A2(n7435), .ZN(n5352) );
  INV_X1 U6844 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6123) );
  OR2_X1 U6845 ( .A1(n6581), .A2(n6123), .ZN(n5351) );
  MUX2_X1 U6846 ( .A(n5355), .B(n7443), .S(P2_U3893), .Z(n5356) );
  INV_X1 U6847 ( .A(n5356), .ZN(P2_U3500) );
  INV_X1 U6848 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6849 ( .A1(n9476), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5359) );
  NAND2_X1 U6850 ( .A1(n9477), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5358) );
  NAND2_X1 U6851 ( .A1(n4491), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5357) );
  AND3_X1 U6852 ( .A1(n5359), .A2(n5358), .A3(n5357), .ZN(n9482) );
  INV_X1 U6853 ( .A(n9482), .ZN(n9765) );
  NAND2_X1 U6854 ( .A1(n9765), .A2(P1_U3973), .ZN(n5360) );
  OAI21_X1 U6855 ( .B1(P1_U3973), .B2(n5361), .A(n5360), .ZN(P1_U3585) );
  INV_X1 U6856 ( .A(n5833), .ZN(n7049) );
  NOR2_X1 U6857 ( .A1(n5834), .A2(n7049), .ZN(n5362) );
  INV_X1 U6858 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n5372) );
  NOR2_X1 U6859 ( .A1(n5820), .A2(P2_U3151), .ZN(n7385) );
  INV_X1 U6860 ( .A(n5373), .ZN(n5384) );
  INV_X1 U6861 ( .A(n5820), .ZN(n7983) );
  INV_X1 U6862 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5363) );
  INV_X1 U6863 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5795) );
  MUX2_X1 U6864 ( .A(n5363), .B(n5795), .S(n8512), .Z(n5364) );
  NAND2_X1 U6865 ( .A1(n5364), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n5550) );
  MUX2_X1 U6866 ( .A(P2_REG2_REG_0__SCAN_IN), .B(P2_REG1_REG_0__SCAN_IN), .S(
        n8512), .Z(n5365) );
  INV_X1 U6867 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n5805) );
  NAND2_X1 U6868 ( .A1(n5365), .A2(n5805), .ZN(n5366) );
  AOI22_X1 U6869 ( .A1(n5384), .A2(n8517), .B1(n5550), .B2(n5366), .ZN(n5367)
         );
  AOI21_X1 U6870 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .A(n5367), .ZN(
        n5371) );
  NOR2_X1 U6871 ( .A1(n8512), .A2(P2_U3151), .ZN(n7202) );
  NAND2_X1 U6872 ( .A1(n5368), .A2(n7202), .ZN(n5369) );
  MUX2_X1 U6873 ( .A(n8485), .B(n5369), .S(n5820), .Z(n8522) );
  NAND2_X1 U6874 ( .A1(n8448), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n5370) );
  OAI211_X1 U6875 ( .C1(n5939), .C2(n5372), .A(n5371), .B(n5370), .ZN(P2_U3182) );
  INV_X1 U6876 ( .A(n8512), .ZN(n5383) );
  INV_X1 U6877 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6189) );
  XNOR2_X1 U6878 ( .A(n7993), .B(n6189), .ZN(n5505) );
  AND2_X1 U6879 ( .A1(n5374), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5378) );
  NAND2_X1 U6880 ( .A1(n5805), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5377) );
  OAI22_X1 U6881 ( .A1(n5378), .A2(n5784), .B1(n5374), .B2(n5377), .ZN(n5552)
         );
  NAND2_X1 U6882 ( .A1(n5552), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5379) );
  OAI21_X1 U6883 ( .B1(n5363), .B2(n4710), .A(n5379), .ZN(n5506) );
  NAND2_X1 U6884 ( .A1(n5505), .A2(n5506), .ZN(n5381) );
  NAND2_X1 U6885 ( .A1(n7993), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5380) );
  NAND2_X1 U6886 ( .A1(n5381), .A2(n5380), .ZN(n5577) );
  XNOR2_X1 U6887 ( .A(n5577), .B(n6035), .ZN(n5575) );
  XNOR2_X1 U6888 ( .A(n5575), .B(P2_REG2_REG_3__SCAN_IN), .ZN(n5393) );
  INV_X1 U6889 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5382) );
  NOR2_X1 U6890 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5382), .ZN(n6050) );
  INV_X1 U6891 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n5391) );
  AND2_X1 U6892 ( .A1(n5374), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5386) );
  NAND2_X1 U6893 ( .A1(n5805), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5385) );
  OAI22_X1 U6894 ( .A1(n5386), .A2(n5784), .B1(n5374), .B2(n5385), .ZN(n5553)
         );
  NAND2_X1 U6895 ( .A1(n5553), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5388) );
  INV_X1 U6896 ( .A(n5386), .ZN(n5387) );
  NAND2_X1 U6897 ( .A1(n5388), .A2(n5387), .ZN(n5501) );
  NAND2_X1 U6898 ( .A1(n7993), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5389) );
  XNOR2_X1 U6899 ( .A(n5570), .B(n6035), .ZN(n5569) );
  INV_X1 U6900 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5824) );
  XNOR2_X1 U6901 ( .A(n5569), .B(n5824), .ZN(n5390) );
  OAI22_X1 U6902 ( .A1(n5939), .A2(n5391), .B1(n8529), .B2(n5390), .ZN(n5392)
         );
  AOI211_X1 U6903 ( .C1(n8526), .C2(n5393), .A(n6050), .B(n5392), .ZN(n5405)
         );
  MUX2_X1 U6904 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8512), .Z(n5395) );
  XNOR2_X1 U6905 ( .A(n5395), .B(n5784), .ZN(n5551) );
  NAND2_X1 U6906 ( .A1(n5551), .A2(n5550), .ZN(n5397) );
  NAND2_X1 U6907 ( .A1(n5395), .A2(n5394), .ZN(n5396) );
  NAND2_X1 U6908 ( .A1(n5397), .A2(n5396), .ZN(n5499) );
  MUX2_X1 U6909 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8512), .Z(n5398) );
  INV_X1 U6910 ( .A(n7993), .ZN(n5511) );
  XNOR2_X1 U6911 ( .A(n5398), .B(n5511), .ZN(n5498) );
  INV_X1 U6912 ( .A(n5398), .ZN(n5399) );
  NOR2_X1 U6913 ( .A1(n5399), .A2(n5511), .ZN(n5400) );
  AOI21_X1 U6914 ( .B1(n5499), .B2(n5498), .A(n5400), .ZN(n5402) );
  MUX2_X1 U6915 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8512), .Z(n5562) );
  XNOR2_X1 U6916 ( .A(n5562), .B(n6035), .ZN(n5401) );
  NAND2_X1 U6917 ( .A1(n5402), .A2(n5401), .ZN(n8431) );
  OAI21_X1 U6918 ( .B1(n5402), .B2(n5401), .A(n8431), .ZN(n5403) );
  NAND2_X1 U6919 ( .A1(n5403), .A2(n8464), .ZN(n5404) );
  OAI211_X1 U6920 ( .C1(n8522), .C2(n5576), .A(n5405), .B(n5404), .ZN(P2_U3185) );
  OR2_X1 U6921 ( .A1(n5065), .A2(n5314), .ZN(n5407) );
  XNOR2_X1 U6922 ( .A(n5407), .B(n5406), .ZN(n6528) );
  OAI222_X1 U6923 ( .A1(n9222), .A2(n5409), .B1(n7594), .B2(n5408), .C1(
        P2_U3151), .C2(n6528), .ZN(P2_U3284) );
  INV_X1 U6924 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10281) );
  MUX2_X1 U6925 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10281), .S(n9658), .Z(n9661)
         );
  INV_X1 U6926 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n5411) );
  XNOR2_X1 U6927 ( .A(n9645), .B(n5411), .ZN(n9643) );
  AND2_X1 U6928 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9642) );
  NAND2_X1 U6929 ( .A1(n9643), .A2(n9642), .ZN(n9641) );
  NAND2_X1 U6930 ( .A1(n9645), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5412) );
  NAND2_X1 U6931 ( .A1(n9641), .A2(n5412), .ZN(n9660) );
  NAND2_X1 U6932 ( .A1(n9661), .A2(n9660), .ZN(n9659) );
  NAND2_X1 U6933 ( .A1(n9658), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5413) );
  NAND2_X1 U6934 ( .A1(n9659), .A2(n5413), .ZN(n9673) );
  INV_X1 U6935 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n5414) );
  XNOR2_X1 U6936 ( .A(n9671), .B(n5414), .ZN(n9674) );
  NAND2_X1 U6937 ( .A1(n9673), .A2(n9674), .ZN(n9672) );
  NAND2_X1 U6938 ( .A1(n9671), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5415) );
  NAND2_X1 U6939 ( .A1(n9672), .A2(n5415), .ZN(n9690) );
  INV_X1 U6940 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5416) );
  XNOR2_X1 U6941 ( .A(n9685), .B(n5416), .ZN(n9691) );
  NAND2_X1 U6942 ( .A1(n9690), .A2(n9691), .ZN(n9689) );
  INV_X1 U6943 ( .A(n9689), .ZN(n5417) );
  AOI21_X1 U6944 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n9685), .A(n5417), .ZN(
        n5437) );
  XNOR2_X1 U6945 ( .A(n5906), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n5436) );
  NOR2_X1 U6946 ( .A1(n5437), .A2(n5436), .ZN(n5435) );
  AOI21_X1 U6947 ( .B1(n5906), .B2(P1_REG1_REG_5__SCAN_IN), .A(n5435), .ZN(
        n5419) );
  XOR2_X1 U6948 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6197), .Z(n5418) );
  NOR2_X1 U6949 ( .A1(n5419), .A2(n5418), .ZN(n5447) );
  AOI211_X1 U6950 ( .C1(n5419), .C2(n5418), .A(n5447), .B(n9751), .ZN(n5434)
         );
  INV_X1 U6951 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n5421) );
  INV_X1 U6952 ( .A(n6197), .ZN(n5453) );
  NAND2_X1 U6953 ( .A1(n9755), .A2(n5453), .ZN(n5420) );
  NAND2_X1 U6954 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6374) );
  OAI211_X1 U6955 ( .C1(n5421), .C2(n9761), .A(n5420), .B(n6374), .ZN(n5433)
         );
  INV_X1 U6956 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5422) );
  MUX2_X1 U6957 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n5422), .S(n9658), .Z(n9664)
         );
  INV_X1 U6958 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6281) );
  XNOR2_X1 U6959 ( .A(n9645), .B(n6281), .ZN(n9640) );
  AND2_X1 U6960 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9651) );
  NAND2_X1 U6961 ( .A1(n9640), .A2(n9651), .ZN(n9639) );
  NAND2_X1 U6962 ( .A1(n9645), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5423) );
  NAND2_X1 U6963 ( .A1(n9639), .A2(n5423), .ZN(n9663) );
  NAND2_X1 U6964 ( .A1(n9664), .A2(n9663), .ZN(n9662) );
  NAND2_X1 U6965 ( .A1(n9658), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5424) );
  NAND2_X1 U6966 ( .A1(n9662), .A2(n5424), .ZN(n9676) );
  INV_X1 U6967 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5425) );
  XNOR2_X1 U6968 ( .A(n9671), .B(n5425), .ZN(n9677) );
  NAND2_X1 U6969 ( .A1(n9676), .A2(n9677), .ZN(n9675) );
  NAND2_X1 U6970 ( .A1(n9671), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5426) );
  NAND2_X1 U6971 ( .A1(n9675), .A2(n5426), .ZN(n9687) );
  INV_X1 U6972 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5427) );
  XNOR2_X1 U6973 ( .A(n9685), .B(n5427), .ZN(n9688) );
  XNOR2_X1 U6974 ( .A(n5906), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n5442) );
  AOI21_X1 U6975 ( .B1(n5906), .B2(P1_REG2_REG_5__SCAN_IN), .A(n5441), .ZN(
        n5431) );
  XOR2_X1 U6976 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6197), .Z(n5430) );
  NOR2_X1 U6977 ( .A1(n5431), .A2(n5430), .ZN(n5452) );
  NAND2_X1 U6978 ( .A1(n9652), .A2(n9762), .ZN(n5428) );
  AOI211_X1 U6979 ( .C1(n5431), .C2(n5430), .A(n5452), .B(n9752), .ZN(n5432)
         );
  OR3_X1 U6980 ( .A1(n5434), .A2(n5433), .A3(n5432), .ZN(P1_U3249) );
  AOI211_X1 U6981 ( .C1(n5437), .C2(n5436), .A(n5435), .B(n9751), .ZN(n5446)
         );
  INV_X1 U6982 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n5440) );
  NAND2_X1 U6983 ( .A1(n9755), .A2(n5906), .ZN(n5439) );
  INV_X1 U6984 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n8970) );
  NOR2_X1 U6985 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8970), .ZN(n6269) );
  INV_X1 U6986 ( .A(n6269), .ZN(n5438) );
  OAI211_X1 U6987 ( .C1(n5440), .C2(n9761), .A(n5439), .B(n5438), .ZN(n5445)
         );
  AOI211_X1 U6988 ( .C1(n5443), .C2(n5442), .A(n5441), .B(n9752), .ZN(n5444)
         );
  OR3_X1 U6989 ( .A1(n5446), .A2(n5445), .A3(n5444), .ZN(P1_U3248) );
  AOI21_X1 U6990 ( .B1(n5453), .B2(P1_REG1_REG_6__SCAN_IN), .A(n5447), .ZN(
        n5465) );
  INV_X1 U6991 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5448) );
  MUX2_X1 U6992 ( .A(n5448), .B(P1_REG1_REG_7__SCAN_IN), .S(n6207), .Z(n5464)
         );
  NOR2_X1 U6993 ( .A1(n5465), .A2(n5464), .ZN(n5463) );
  AOI21_X1 U6994 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n6207), .A(n5463), .ZN(
        n5451) );
  INV_X1 U6995 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n5449) );
  MUX2_X1 U6996 ( .A(n5449), .B(P1_REG1_REG_8__SCAN_IN), .S(n6309), .Z(n5450)
         );
  NOR2_X1 U6997 ( .A1(n5451), .A2(n5450), .ZN(n5488) );
  AOI211_X1 U6998 ( .C1(n5451), .C2(n5450), .A(n5488), .B(n9751), .ZN(n5462)
         );
  AOI21_X1 U6999 ( .B1(n5453), .B2(P1_REG2_REG_6__SCAN_IN), .A(n5452), .ZN(
        n5468) );
  NAND2_X1 U7000 ( .A1(n6207), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5454) );
  OAI21_X1 U7001 ( .B1(n6207), .B2(P1_REG2_REG_7__SCAN_IN), .A(n5454), .ZN(
        n5467) );
  NOR2_X1 U7002 ( .A1(n5468), .A2(n5467), .ZN(n5466) );
  NAND2_X1 U7003 ( .A1(n6309), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5455) );
  OAI21_X1 U7004 ( .B1(n6309), .B2(P1_REG2_REG_8__SCAN_IN), .A(n5455), .ZN(
        n5456) );
  AOI211_X1 U7005 ( .C1(n5457), .C2(n5456), .A(n5485), .B(n9752), .ZN(n5461)
         );
  INV_X1 U7006 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U7007 ( .A1(n9755), .A2(n6309), .ZN(n5458) );
  NAND2_X1 U7008 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7039) );
  OAI211_X1 U7009 ( .C1(n5459), .C2(n9761), .A(n5458), .B(n7039), .ZN(n5460)
         );
  OR3_X1 U7010 ( .A1(n5462), .A2(n5461), .A3(n5460), .ZN(P1_U3251) );
  AOI211_X1 U7011 ( .C1(n5465), .C2(n5464), .A(n9751), .B(n5463), .ZN(n5475)
         );
  AOI211_X1 U7012 ( .C1(n5468), .C2(n5467), .A(n9752), .B(n5466), .ZN(n5474)
         );
  INV_X1 U7013 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U7014 ( .A1(n9755), .A2(n6207), .ZN(n5471) );
  INV_X1 U7015 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5469) );
  NOR2_X1 U7016 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5469), .ZN(n6560) );
  INV_X1 U7017 ( .A(n6560), .ZN(n5470) );
  OAI211_X1 U7018 ( .C1(n5472), .C2(n9761), .A(n5471), .B(n5470), .ZN(n5473)
         );
  OR3_X1 U7019 ( .A1(n5475), .A2(n5474), .A3(n5473), .ZN(P1_U3250) );
  INV_X1 U7020 ( .A(n5476), .ZN(n5478) );
  AND2_X1 U7021 ( .A1(n5478), .A2(n5477), .ZN(n5479) );
  MUX2_X1 U7022 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n7901), .Z(n5545) );
  XNOR2_X1 U7023 ( .A(n5545), .B(n9082), .ZN(n5544) );
  XNOR2_X1 U7024 ( .A(n5547), .B(n5544), .ZN(n7060) );
  INV_X1 U7025 ( .A(n7060), .ZN(n5543) );
  OR2_X1 U7026 ( .A1(n5614), .A2(n5314), .ZN(n5482) );
  XNOR2_X1 U7027 ( .A(n5482), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7061) );
  INV_X1 U7028 ( .A(n7061), .ZN(n6534) );
  INV_X1 U7029 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5483) );
  OAI222_X1 U7030 ( .A1(n7594), .A2(n5543), .B1(n6534), .B2(P2_U3151), .C1(
        n5483), .C2(n9222), .ZN(P2_U3283) );
  NOR2_X1 U7031 ( .A1(n6440), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5484) );
  AOI21_X1 U7032 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n6440), .A(n5484), .ZN(
        n5487) );
  OAI21_X1 U7033 ( .B1(n5487), .B2(n5486), .A(n5679), .ZN(n5496) );
  INV_X1 U7034 ( .A(n9755), .ZN(n7509) );
  INV_X1 U7035 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10286) );
  AOI22_X1 U7036 ( .A1(n6440), .A2(P1_REG1_REG_9__SCAN_IN), .B1(n10286), .B2(
        n5494), .ZN(n5490) );
  AOI21_X1 U7037 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n6309), .A(n5488), .ZN(
        n5489) );
  NAND2_X1 U7038 ( .A1(n5490), .A2(n5489), .ZN(n5675) );
  OAI21_X1 U7039 ( .B1(n5490), .B2(n5489), .A(n5675), .ZN(n5491) );
  NAND2_X1 U7040 ( .A1(n5491), .A2(n9756), .ZN(n5493) );
  NOR2_X1 U7041 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6299), .ZN(n7116) );
  AOI21_X1 U7042 ( .B1(n9644), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n7116), .ZN(
        n5492) );
  OAI211_X1 U7043 ( .C1(n7509), .C2(n5494), .A(n5493), .B(n5492), .ZN(n5495)
         );
  AOI21_X1 U7044 ( .B1(n9740), .B2(n5496), .A(n5495), .ZN(n5497) );
  INV_X1 U7045 ( .A(n5497), .ZN(P1_U3252) );
  XNOR2_X1 U7046 ( .A(n5499), .B(n5498), .ZN(n5513) );
  INV_X1 U7047 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9093) );
  OAI21_X1 U7048 ( .B1(n5502), .B2(n5501), .A(n5500), .ZN(n5503) );
  NAND2_X1 U7049 ( .A1(n8442), .A2(n5503), .ZN(n5504) );
  OAI21_X1 U7050 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n9093), .A(n5504), .ZN(n5510) );
  INV_X1 U7051 ( .A(n8526), .ZN(n5558) );
  XOR2_X1 U7052 ( .A(n5506), .B(n5505), .Z(n5508) );
  INV_X1 U7053 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n5507) );
  OAI22_X1 U7054 ( .A1(n5558), .A2(n5508), .B1(n5507), .B2(n5939), .ZN(n5509)
         );
  AOI211_X1 U7055 ( .C1(n5511), .C2(n8448), .A(n5510), .B(n5509), .ZN(n5512)
         );
  OAI21_X1 U7056 ( .B1(n8517), .B2(n5513), .A(n5512), .ZN(P2_U3184) );
  INV_X1 U7057 ( .A(n5594), .ZN(n5605) );
  INV_X1 U7058 ( .A(n6278), .ZN(n5515) );
  INV_X4 U7059 ( .A(n5521), .ZN(n8226) );
  NAND2_X1 U7060 ( .A1(n6278), .A2(n5516), .ZN(n5517) );
  NAND2_X4 U7061 ( .A1(n5518), .A2(n5519), .ZN(n5702) );
  AND2_X2 U7062 ( .A1(n5702), .A2(n8097), .ZN(n5716) );
  OAI22_X1 U7063 ( .A1(n5605), .A2(n8226), .B1(n5716), .B2(n9530), .ZN(n5618)
         );
  AOI21_X1 U7064 ( .B1(P1_REG1_REG_0__SCAN_IN), .B2(n5522), .A(n5618), .ZN(
        n5620) );
  NAND2_X1 U7065 ( .A1(n5594), .A2(n8182), .ZN(n5524) );
  AOI22_X1 U7066 ( .A1(n6705), .A2(n5521), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n5522), .ZN(n5523) );
  AND2_X1 U7067 ( .A1(n5524), .A2(n5523), .ZN(n5619) );
  XNOR2_X1 U7068 ( .A(n5620), .B(n5619), .ZN(n9650) );
  INV_X1 U7069 ( .A(n6706), .ZN(n5525) );
  NOR2_X1 U7070 ( .A1(n10117), .A2(n9602), .ZN(n5527) );
  INV_X1 U7071 ( .A(n10239), .ZN(n6275) );
  AND3_X1 U7072 ( .A1(n10168), .A2(n6274), .A3(n5526), .ZN(n5534) );
  INV_X1 U7073 ( .A(n10117), .ZN(n10274) );
  NOR2_X1 U7074 ( .A1(n6706), .A2(n9577), .ZN(n6282) );
  INV_X1 U7075 ( .A(n5534), .ZN(n5528) );
  OAI21_X1 U7076 ( .B1(n10274), .B2(n6282), .A(n5528), .ZN(n5531) );
  AND3_X1 U7077 ( .A1(n5529), .A2(n6985), .A3(n5519), .ZN(n5530) );
  NAND2_X1 U7078 ( .A1(n5531), .A2(n5530), .ZN(n5726) );
  OR2_X1 U7079 ( .A1(n5726), .A2(P1_U3086), .ZN(n9326) );
  NAND3_X1 U7080 ( .A1(n6275), .A2(n5534), .A3(n6282), .ZN(n5533) );
  INV_X1 U7081 ( .A(n9363), .ZN(n9350) );
  NAND3_X1 U7082 ( .A1(n6275), .A2(n5535), .A3(n5534), .ZN(n5628) );
  INV_X1 U7083 ( .A(n5593), .ZN(n5732) );
  OAI22_X1 U7084 ( .A1(n9350), .A2(n9530), .B1(n9345), .B2(n5732), .ZN(n5536)
         );
  AOI21_X1 U7085 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n9326), .A(n5536), .ZN(
        n5537) );
  OAI21_X1 U7086 ( .B1(n9650), .B2(n9365), .A(n5537), .ZN(P1_U3232) );
  INV_X1 U7087 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n8998) );
  NOR2_X1 U7088 ( .A1(n5538), .A2(n10169), .ZN(n5539) );
  MUX2_X1 U7089 ( .A(n10169), .B(n5539), .S(P1_IR_REG_12__SCAN_IN), .Z(n5542)
         );
  INV_X1 U7090 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5540) );
  NAND2_X1 U7091 ( .A1(n5538), .A2(n5540), .ZN(n5642) );
  INV_X1 U7092 ( .A(n5642), .ZN(n5541) );
  OAI222_X1 U7093 ( .A1(n8278), .A2(n8998), .B1(n10173), .B2(n5543), .C1(n7150), .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U7094 ( .A(n5544), .ZN(n5546) );
  MUX2_X1 U7095 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n7901), .Z(n5635) );
  XNOR2_X1 U7096 ( .A(n5635), .B(SI_13_), .ZN(n5632) );
  INV_X1 U7097 ( .A(n7252), .ZN(n5616) );
  NAND2_X1 U7098 ( .A1(n5642), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5548) );
  XNOR2_X1 U7099 ( .A(n5548), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9699) );
  AOI22_X1 U7100 ( .A1(n9699), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n10171), .ZN(n5549) );
  OAI21_X1 U7101 ( .B1(n5616), .B2(n10173), .A(n5549), .ZN(P1_U3342) );
  XNOR2_X1 U7102 ( .A(n5551), .B(n5550), .ZN(n5561) );
  INV_X1 U7103 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6348) );
  XNOR2_X1 U7104 ( .A(n5552), .B(n6348), .ZN(n5557) );
  XNOR2_X1 U7105 ( .A(n5553), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n5554) );
  AOI22_X1 U7106 ( .A1(n8519), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(n8442), .B2(
        n5554), .ZN(n5556) );
  NAND2_X1 U7107 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(P2_U3151), .ZN(n5555) );
  OAI211_X1 U7108 ( .C1(n5558), .C2(n5557), .A(n5556), .B(n5555), .ZN(n5559)
         );
  AOI21_X1 U7109 ( .B1(n5784), .B2(n8448), .A(n5559), .ZN(n5560) );
  OAI21_X1 U7110 ( .B1(n8517), .B2(n5561), .A(n5560), .ZN(P2_U3183) );
  MUX2_X1 U7111 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8512), .Z(n5652) );
  XNOR2_X1 U7112 ( .A(n5652), .B(n6233), .ZN(n5650) );
  INV_X1 U7113 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6042) );
  INV_X1 U7114 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6043) );
  MUX2_X1 U7115 ( .A(n6042), .B(n6043), .S(n8512), .Z(n5564) );
  XNOR2_X1 U7116 ( .A(n5564), .B(n8447), .ZN(n8432) );
  NOR2_X1 U7117 ( .A1(n5562), .A2(n5576), .ZN(n8433) );
  NOR2_X1 U7118 ( .A1(n8432), .A2(n8433), .ZN(n5563) );
  NAND2_X1 U7119 ( .A1(n8431), .A2(n5563), .ZN(n8435) );
  INV_X1 U7120 ( .A(n5564), .ZN(n5566) );
  NAND2_X1 U7121 ( .A1(n5566), .A2(n5565), .ZN(n5567) );
  NAND2_X1 U7122 ( .A1(n8435), .A2(n5567), .ZN(n5651) );
  XOR2_X1 U7123 ( .A(n5650), .B(n5651), .Z(n5587) );
  NAND2_X1 U7124 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3151), .ZN(n6247) );
  INV_X1 U7125 ( .A(n6247), .ZN(n5568) );
  AOI21_X1 U7126 ( .B1(n8519), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n5568), .ZN(
        n5585) );
  NAND2_X1 U7127 ( .A1(n5569), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5572) );
  NAND2_X1 U7128 ( .A1(n5570), .A2(n5576), .ZN(n5571) );
  NAND2_X1 U7129 ( .A1(n5572), .A2(n5571), .ZN(n8438) );
  MUX2_X1 U7130 ( .A(n6043), .B(P2_REG1_REG_4__SCAN_IN), .S(n8447), .Z(n8439)
         );
  NAND2_X1 U7131 ( .A1(n8438), .A2(n8439), .ZN(n8437) );
  OR2_X1 U7132 ( .A1(n8447), .A2(n6043), .ZN(n5573) );
  NAND2_X1 U7133 ( .A1(n8437), .A2(n5573), .ZN(n5663) );
  XNOR2_X1 U7134 ( .A(n5663), .B(n6233), .ZN(n5665) );
  INV_X1 U7135 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6107) );
  XNOR2_X1 U7136 ( .A(n5665), .B(n6107), .ZN(n5574) );
  OR2_X1 U7137 ( .A1(n8529), .A2(n5574), .ZN(n5584) );
  NAND2_X1 U7138 ( .A1(n5575), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5579) );
  NAND2_X1 U7139 ( .A1(n5577), .A2(n5576), .ZN(n5578) );
  NAND2_X1 U7140 ( .A1(n5579), .A2(n5578), .ZN(n8444) );
  MUX2_X1 U7141 ( .A(n6042), .B(P2_REG2_REG_4__SCAN_IN), .S(n8447), .Z(n8445)
         );
  NAND2_X1 U7142 ( .A1(n8444), .A2(n8445), .ZN(n8443) );
  OR2_X1 U7143 ( .A1(n8447), .A2(n6042), .ZN(n5580) );
  NAND2_X1 U7144 ( .A1(n8443), .A2(n5580), .ZN(n5658) );
  XNOR2_X1 U7145 ( .A(n5658), .B(n6233), .ZN(n5659) );
  XNOR2_X1 U7146 ( .A(n5659), .B(P2_REG2_REG_5__SCAN_IN), .ZN(n5581) );
  NAND2_X1 U7147 ( .A1(n8526), .A2(n5581), .ZN(n5583) );
  OR2_X1 U7148 ( .A1(n8522), .A2(n5664), .ZN(n5582) );
  NAND4_X1 U7149 ( .A1(n5585), .A2(n5584), .A3(n5583), .A4(n5582), .ZN(n5586)
         );
  AOI21_X1 U7150 ( .B1(n5587), .B2(n8464), .A(n5586), .ZN(n5588) );
  INV_X1 U7151 ( .A(n5588), .ZN(P2_U3187) );
  NAND2_X1 U7152 ( .A1(n5895), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5591) );
  NAND2_X1 U7153 ( .A1(n8043), .A2(n9645), .ZN(n5590) );
  AND3_X2 U7154 ( .A1(n5592), .A2(n5591), .A3(n5590), .ZN(n5597) );
  XNOR2_X1 U7155 ( .A(n5593), .B(n5597), .ZN(n5595) );
  NAND2_X1 U7156 ( .A1(n5594), .A2(n6705), .ZN(n5596) );
  NAND2_X1 U7157 ( .A1(n5596), .A2(n5595), .ZN(n5734) );
  OAI21_X1 U7158 ( .B1(n5595), .B2(n5596), .A(n5734), .ZN(n5609) );
  AOI211_X1 U7159 ( .C1(n6705), .C2(n5743), .A(n10266), .B(n6802), .ZN(n6285)
         );
  INV_X1 U7160 ( .A(n5609), .ZN(n6288) );
  INV_X1 U7161 ( .A(n5595), .ZN(n9492) );
  NOR2_X1 U7162 ( .A1(n5594), .A2(n9530), .ZN(n5598) );
  NAND2_X1 U7163 ( .A1(n9492), .A2(n5598), .ZN(n5745) );
  OAI21_X1 U7164 ( .B1(n9492), .B2(n5598), .A(n5745), .ZN(n5607) );
  NAND2_X1 U7165 ( .A1(n5720), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5604) );
  NAND2_X1 U7166 ( .A1(n5708), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5601) );
  NAND2_X1 U7167 ( .A1(n5599), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5600) );
  NAND2_X1 U7168 ( .A1(n4492), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5602) );
  OAI22_X1 U7169 ( .A1(n5605), .A2(n10011), .B1(n5737), .B2(n10013), .ZN(n5606) );
  AOI21_X1 U7170 ( .B1(n5607), .B2(n10009), .A(n5606), .ZN(n5608) );
  OAI21_X1 U7171 ( .B1(n6288), .B2(n6317), .A(n5608), .ZN(n6279) );
  AOI211_X1 U7172 ( .C1(n6916), .C2(n5609), .A(n6285), .B(n6279), .ZN(n5695)
         );
  INV_X1 U7173 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5610) );
  OAI22_X1 U7174 ( .A1(n10164), .A2(n5597), .B1(n10280), .B2(n5610), .ZN(n5611) );
  INV_X1 U7175 ( .A(n5611), .ZN(n5612) );
  OAI21_X1 U7176 ( .B1(n5695), .B2(n10278), .A(n5612), .ZN(P1_U3456) );
  INV_X1 U7177 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U7178 ( .A1(n5614), .A2(n5613), .ZN(n5687) );
  NAND2_X1 U7179 ( .A1(n5687), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5615) );
  XNOR2_X1 U7180 ( .A(n5615), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7253) );
  INV_X1 U7181 ( .A(n7253), .ZN(n6944) );
  OAI222_X1 U7182 ( .A1(n9222), .A2(n5617), .B1(n9220), .B2(n5616), .C1(
        P2_U3151), .C2(n6944), .ZN(P2_U3282) );
  OAI22_X1 U7183 ( .A1(n5620), .A2(n5619), .B1(n4495), .B2(n5618), .ZN(n5627)
         );
  NAND2_X1 U7184 ( .A1(n5593), .A2(n5521), .ZN(n5621) );
  OAI21_X1 U7185 ( .B1(n5716), .B2(n5597), .A(n5621), .ZN(n5622) );
  XNOR2_X1 U7186 ( .A(n5622), .B(n8194), .ZN(n5624) );
  AOI22_X1 U7187 ( .A1(n5593), .A2(n8182), .B1(n5743), .B2(n5521), .ZN(n5623)
         );
  NAND2_X1 U7188 ( .A1(n5624), .A2(n5623), .ZN(n5696) );
  OR2_X1 U7189 ( .A1(n5624), .A2(n5623), .ZN(n5625) );
  NAND2_X1 U7190 ( .A1(n5696), .A2(n5625), .ZN(n5626) );
  AOI21_X1 U7191 ( .B1(n5627), .B2(n5626), .A(n9322), .ZN(n5631) );
  AOI22_X1 U7192 ( .A1(n9334), .A2(n5594), .B1(n5743), .B2(n9363), .ZN(n5630)
         );
  AOI22_X1 U7193 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(n9326), .B1(n9355), .B2(
        n5735), .ZN(n5629) );
  OAI211_X1 U7194 ( .C1(n5631), .C2(n9365), .A(n5630), .B(n5629), .ZN(P1_U3222) );
  INV_X1 U7195 ( .A(n5632), .ZN(n5633) );
  NAND2_X1 U7196 ( .A1(n5635), .A2(SI_13_), .ZN(n5636) );
  INV_X1 U7197 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n5637) );
  MUX2_X1 U7198 ( .A(n8874), .B(n5637), .S(n7901), .Z(n5639) );
  INV_X1 U7199 ( .A(SI_14_), .ZN(n5638) );
  NAND2_X1 U7200 ( .A1(n5639), .A2(n5638), .ZN(n5959) );
  INV_X1 U7201 ( .A(n5639), .ZN(n5640) );
  NAND2_X1 U7202 ( .A1(n5640), .A2(SI_14_), .ZN(n5641) );
  NAND2_X1 U7203 ( .A1(n5959), .A2(n5641), .ZN(n5756) );
  XNOR2_X1 U7204 ( .A(n5755), .B(n5756), .ZN(n7261) );
  INV_X1 U7205 ( .A(n7261), .ZN(n5691) );
  OR2_X1 U7206 ( .A1(n5642), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5643) );
  NAND2_X1 U7207 ( .A1(n5643), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5644) );
  OR2_X1 U7208 ( .A1(n5644), .A2(n9084), .ZN(n5645) );
  NAND2_X1 U7209 ( .A1(n5644), .A2(n9084), .ZN(n5846) );
  AOI22_X1 U7210 ( .A1(n9712), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n10171), .ZN(n5646) );
  OAI21_X1 U7211 ( .B1(n5691), .B2(n10173), .A(n5646), .ZN(P1_U3341) );
  INV_X1 U7212 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6239) );
  INV_X1 U7213 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6242) );
  MUX2_X1 U7214 ( .A(n6239), .B(n6242), .S(n8512), .Z(n5647) );
  NAND2_X1 U7215 ( .A1(n5647), .A2(n6565), .ZN(n5946) );
  INV_X1 U7216 ( .A(n5647), .ZN(n5648) );
  NAND2_X1 U7217 ( .A1(n5648), .A2(n5952), .ZN(n5649) );
  NAND2_X1 U7218 ( .A1(n5946), .A2(n5649), .ZN(n5657) );
  NAND2_X1 U7219 ( .A1(n5651), .A2(n5650), .ZN(n5654) );
  NAND2_X1 U7220 ( .A1(n5652), .A2(n5664), .ZN(n5653) );
  NAND2_X1 U7221 ( .A1(n5654), .A2(n5653), .ZN(n5656) );
  OR2_X1 U7222 ( .A1(n5656), .A2(n5657), .ZN(n5947) );
  INV_X1 U7223 ( .A(n5947), .ZN(n5655) );
  AOI21_X1 U7224 ( .B1(n5657), .B2(n5656), .A(n5655), .ZN(n5674) );
  MUX2_X1 U7225 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6239), .S(n6565), .Z(n5661)
         );
  AOI22_X1 U7226 ( .A1(n5659), .A2(P2_REG2_REG_5__SCAN_IN), .B1(n5664), .B2(
        n5658), .ZN(n5660) );
  NOR2_X1 U7227 ( .A1(n5660), .A2(n5661), .ZN(n5951) );
  AOI21_X1 U7228 ( .B1(n5661), .B2(n5660), .A(n5951), .ZN(n5662) );
  INV_X1 U7229 ( .A(n5662), .ZN(n5672) );
  MUX2_X1 U7230 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6242), .S(n6565), .Z(n5667)
         );
  AOI22_X1 U7231 ( .A1(n5665), .A2(P2_REG1_REG_5__SCAN_IN), .B1(n5664), .B2(
        n5663), .ZN(n5666) );
  NOR2_X1 U7232 ( .A1(n5666), .A2(n5667), .ZN(n5936) );
  AOI21_X1 U7233 ( .B1(n5667), .B2(n5666), .A(n5936), .ZN(n5668) );
  NOR2_X1 U7234 ( .A1(n5668), .A2(n8529), .ZN(n5671) );
  AND2_X1 U7235 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6784) );
  AOI21_X1 U7236 ( .B1(n8519), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n6784), .ZN(
        n5669) );
  OAI21_X1 U7237 ( .B1(n5952), .B2(n8522), .A(n5669), .ZN(n5670) );
  AOI211_X1 U7238 ( .C1(n8526), .C2(n5672), .A(n5671), .B(n5670), .ZN(n5673)
         );
  OAI21_X1 U7239 ( .B1(n5674), .B2(n8517), .A(n5673), .ZN(P2_U3188) );
  MUX2_X1 U7240 ( .A(n10288), .B(P1_REG1_REG_10__SCAN_IN), .S(n6644), .Z(n5677) );
  OAI21_X1 U7241 ( .B1(n6440), .B2(P1_REG1_REG_9__SCAN_IN), .A(n5675), .ZN(
        n5676) );
  NOR2_X1 U7242 ( .A1(n5676), .A2(n5677), .ZN(n5851) );
  AOI211_X1 U7243 ( .C1(n5677), .C2(n5676), .A(n9751), .B(n5851), .ZN(n5686)
         );
  INV_X1 U7244 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n5678) );
  MUX2_X1 U7245 ( .A(n5678), .B(P1_REG2_REG_10__SCAN_IN), .S(n6644), .Z(n5681)
         );
  OAI21_X1 U7246 ( .B1(n6440), .B2(P1_REG2_REG_9__SCAN_IN), .A(n5679), .ZN(
        n5680) );
  NOR2_X1 U7247 ( .A1(n5680), .A2(n5681), .ZN(n5855) );
  AOI211_X1 U7248 ( .C1(n5681), .C2(n5680), .A(n9752), .B(n5855), .ZN(n5685)
         );
  INV_X1 U7249 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U7250 ( .A1(n9755), .A2(n6644), .ZN(n5682) );
  NAND2_X1 U7251 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7326) );
  OAI211_X1 U7252 ( .C1(n5683), .C2(n9761), .A(n5682), .B(n7326), .ZN(n5684)
         );
  OR3_X1 U7253 ( .A1(n5686), .A2(n5685), .A3(n5684), .ZN(P1_U3253) );
  NAND2_X1 U7254 ( .A1(n5688), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5973) );
  OR2_X1 U7255 ( .A1(n5973), .A2(n5689), .ZN(n5690) );
  NAND2_X1 U7256 ( .A1(n5973), .A2(n5689), .ZN(n5759) );
  INV_X1 U7257 ( .A(n7262), .ZN(n6959) );
  OAI222_X1 U7258 ( .A1(n9222), .A2(n8874), .B1(n9220), .B2(n5691), .C1(
        P2_U3151), .C2(n6959), .ZN(P2_U3281) );
  OAI22_X1 U7259 ( .A1(n10108), .A2(n5597), .B1(n10293), .B2(n5411), .ZN(n5693) );
  INV_X1 U7260 ( .A(n5693), .ZN(n5694) );
  OAI21_X1 U7261 ( .B1(n5695), .B2(n10290), .A(n5694), .ZN(P1_U3523) );
  INV_X1 U7262 ( .A(n5696), .ZN(n9321) );
  XNOR2_X1 U7263 ( .A(n5698), .B(n5697), .ZN(n7994) );
  NAND2_X1 U7264 ( .A1(n5895), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U7265 ( .A1(n4494), .A2(n9658), .ZN(n5699) );
  OAI22_X1 U7266 ( .A1(n5737), .A2(n8226), .B1(n5736), .B2(n5716), .ZN(n5701)
         );
  XNOR2_X1 U7267 ( .A(n5701), .B(n4495), .ZN(n5704) );
  OAI22_X1 U7268 ( .A1(n5737), .A2(n5702), .B1(n5736), .B2(n8226), .ZN(n5703)
         );
  NAND2_X1 U7269 ( .A1(n5704), .A2(n5703), .ZN(n5705) );
  OAI21_X1 U7270 ( .B1(n9322), .B2(n9321), .A(n9320), .ZN(n9319) );
  INV_X1 U7271 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6336) );
  NAND2_X1 U7272 ( .A1(n5720), .A2(n6336), .ZN(n5709) );
  INV_X1 U7273 ( .A(n5712), .ZN(n5894) );
  NAND2_X1 U7274 ( .A1(n4494), .A2(n9671), .ZN(n5714) );
  NAND2_X1 U7275 ( .A1(n5895), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5713) );
  AOI22_X1 U7276 ( .A1(n5739), .A2(n8182), .B1(n5521), .B2(n5741), .ZN(n6255)
         );
  OAI22_X1 U7277 ( .A1(n6804), .A2(n8226), .B1(n6339), .B2(n5716), .ZN(n5717)
         );
  XNOR2_X1 U7278 ( .A(n5717), .B(n4495), .ZN(n6257) );
  XOR2_X1 U7279 ( .A(n6255), .B(n6257), .Z(n5718) );
  AOI21_X1 U7280 ( .B1(n5719), .B2(n5718), .A(n8268), .ZN(n5731) );
  NAND2_X1 U7281 ( .A1(n4492), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5725) );
  NOR2_X1 U7282 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5721) );
  NOR2_X1 U7283 ( .A1(n5901), .A2(n5721), .ZN(n8272) );
  NAND2_X1 U7284 ( .A1(n5720), .A2(n8272), .ZN(n5724) );
  NAND2_X1 U7285 ( .A1(n5599), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5723) );
  NAND2_X1 U7286 ( .A1(n5708), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5722) );
  AOI22_X1 U7287 ( .A1(n9334), .A2(n5735), .B1(n9355), .B2(n5742), .ZN(n5730)
         );
  NAND2_X1 U7288 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9668) );
  INV_X1 U7289 ( .A(n9668), .ZN(n5728) );
  NOR2_X1 U7290 ( .A1(n9350), .A2(n6339), .ZN(n5727) );
  AOI211_X1 U7291 ( .C1(n9357), .C2(n6336), .A(n5728), .B(n5727), .ZN(n5729)
         );
  OAI211_X1 U7292 ( .C1(n5731), .C2(n9365), .A(n5730), .B(n5729), .ZN(P1_U3218) );
  NAND2_X1 U7293 ( .A1(n5732), .A2(n5597), .ZN(n5733) );
  NAND2_X1 U7294 ( .A1(n5734), .A2(n5733), .ZN(n6800) );
  NAND2_X1 U7295 ( .A1(n5737), .A2(n9325), .ZN(n5746) );
  NAND2_X1 U7296 ( .A1(n6800), .A2(n9490), .ZN(n6799) );
  NAND2_X1 U7297 ( .A1(n5737), .A2(n5736), .ZN(n5738) );
  NAND2_X1 U7298 ( .A1(n6799), .A2(n5738), .ZN(n5740) );
  NAND2_X1 U7299 ( .A1(n6804), .A2(n5741), .ZN(n9538) );
  NAND2_X1 U7300 ( .A1(n9534), .A2(n9538), .ZN(n9491) );
  NAND2_X1 U7301 ( .A1(n5740), .A2(n9491), .ZN(n5893) );
  OAI21_X1 U7302 ( .B1(n5740), .B2(n9491), .A(n5893), .ZN(n6341) );
  INV_X1 U7303 ( .A(n5912), .ZN(n6471) );
  AOI211_X1 U7304 ( .C1(n5741), .C2(n6801), .A(n10266), .B(n6471), .ZN(n6335)
         );
  NAND2_X1 U7305 ( .A1(n5732), .A2(n5743), .ZN(n5744) );
  NAND2_X1 U7306 ( .A1(n9537), .A2(n9535), .ZN(n9370) );
  OR2_X1 U7307 ( .A1(n9370), .A2(n9491), .ZN(n9371) );
  INV_X1 U7308 ( .A(n9371), .ZN(n5747) );
  AOI21_X1 U7309 ( .B1(n9370), .B2(n9491), .A(n5747), .ZN(n5748) );
  OAI222_X1 U7310 ( .A1(n10013), .A2(n6254), .B1(n10011), .B2(n5737), .C1(
        n9938), .C2(n5748), .ZN(n6334) );
  AOI211_X1 U7311 ( .C1(n10276), .C2(n6341), .A(n6335), .B(n6334), .ZN(n5754)
         );
  INV_X1 U7312 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5749) );
  OAI22_X1 U7313 ( .A1(n10164), .A2(n6339), .B1(n10280), .B2(n5749), .ZN(n5750) );
  INV_X1 U7314 ( .A(n5750), .ZN(n5751) );
  OAI21_X1 U7315 ( .B1(n5754), .B2(n10278), .A(n5751), .ZN(P1_U3462) );
  OAI22_X1 U7316 ( .A1(n10108), .A2(n6339), .B1(n10293), .B2(n5414), .ZN(n5752) );
  INV_X1 U7317 ( .A(n5752), .ZN(n5753) );
  OAI21_X1 U7318 ( .B1(n5754), .B2(n10290), .A(n5753), .ZN(P1_U3525) );
  NAND2_X1 U7319 ( .A1(n5962), .A2(n5959), .ZN(n5758) );
  MUX2_X1 U7320 ( .A(n9068), .B(n5850), .S(n7901), .Z(n5963) );
  XNOR2_X1 U7321 ( .A(n5963), .B(SI_15_), .ZN(n5960) );
  XNOR2_X1 U7322 ( .A(n5758), .B(n5960), .ZN(n7353) );
  INV_X1 U7323 ( .A(n7353), .ZN(n5849) );
  NAND2_X1 U7324 ( .A1(n5759), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5760) );
  XNOR2_X1 U7325 ( .A(n5760), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7527) );
  INV_X1 U7326 ( .A(n7527), .ZN(n7521) );
  OAI222_X1 U7327 ( .A1(n7594), .A2(n5849), .B1(n7521), .B2(P2_U3151), .C1(
        n9068), .C2(n9222), .ZN(P2_U3280) );
  AOI21_X2 U7328 ( .B1(n5772), .B2(n5763), .A(n5762), .ZN(n5878) );
  INV_X1 U7329 ( .A(n5878), .ZN(n5780) );
  OR2_X1 U7330 ( .A1(n5877), .A2(n5780), .ZN(n6173) );
  INV_X1 U7331 ( .A(n6173), .ZN(n5775) );
  NOR2_X1 U7332 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .ZN(
        n5767) );
  NOR4_X1 U7333 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n5766) );
  NOR4_X1 U7334 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n5765) );
  NOR4_X1 U7335 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n5764) );
  NAND4_X1 U7336 ( .A1(n5767), .A2(n5766), .A3(n5765), .A4(n5764), .ZN(n5774)
         );
  NOR4_X1 U7337 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5771) );
  NOR4_X1 U7338 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n5770) );
  NOR4_X1 U7339 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n5769) );
  NOR4_X1 U7340 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n5768) );
  NAND4_X1 U7341 ( .A1(n5771), .A2(n5770), .A3(n5769), .A4(n5768), .ZN(n5773)
         );
  NAND2_X1 U7342 ( .A1(n5775), .A2(n5886), .ZN(n5830) );
  INV_X1 U7343 ( .A(n5830), .ZN(n5776) );
  NAND2_X1 U7344 ( .A1(n5776), .A2(n5885), .ZN(n6087) );
  NAND2_X1 U7345 ( .A1(n5778), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5779) );
  NAND2_X1 U7346 ( .A1(n7981), .A2(n7986), .ZN(n5869) );
  NAND3_X1 U7347 ( .A1(n10352), .A2(n6085), .A3(n7893), .ZN(n5829) );
  OR2_X1 U7348 ( .A1(n6087), .A2(n5829), .ZN(n5782) );
  AND2_X1 U7349 ( .A1(n5877), .A2(n5780), .ZN(n5882) );
  NAND2_X1 U7350 ( .A1(n5838), .A2(n5885), .ZN(n6083) );
  OR2_X1 U7351 ( .A1(n6083), .A2(n6085), .ZN(n5781) );
  NAND2_X1 U7352 ( .A1(n5810), .A2(n4519), .ZN(n5785) );
  XNOR2_X1 U7353 ( .A(n5786), .B(n6547), .ZN(n5787) );
  NAND2_X1 U7354 ( .A1(n5787), .A2(n5878), .ZN(n5788) );
  NAND2_X2 U7355 ( .A1(n5788), .A2(n5831), .ZN(n6033) );
  INV_X1 U7356 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n5789) );
  OR2_X1 U7357 ( .A1(n6581), .A2(n5789), .ZN(n5794) );
  NAND2_X1 U7358 ( .A1(n7903), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5793) );
  INV_X1 U7359 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n5931) );
  INV_X1 U7360 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5790) );
  OR2_X1 U7361 ( .A1(n7841), .A2(n5790), .ZN(n5791) );
  XNOR2_X1 U7362 ( .A(n5807), .B(n8429), .ZN(n5928) );
  OR2_X1 U7363 ( .A1(n6581), .A2(n5795), .ZN(n5799) );
  INV_X1 U7364 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n5999) );
  OR2_X1 U7365 ( .A1(n7288), .A2(n5999), .ZN(n5798) );
  INV_X1 U7366 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5796) );
  NAND2_X1 U7367 ( .A1(n5085), .A2(SI_0_), .ZN(n5802) );
  INV_X1 U7368 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5801) );
  NAND2_X1 U7369 ( .A1(n5802), .A2(n5801), .ZN(n5804) );
  NAND2_X1 U7370 ( .A1(n5804), .A2(n5803), .ZN(n9223) );
  INV_X1 U7371 ( .A(n5995), .ZN(n10299) );
  OR2_X1 U7372 ( .A1(n6033), .A2(n10299), .ZN(n5806) );
  NAND2_X1 U7373 ( .A1(n7648), .A2(n5806), .ZN(n5929) );
  NAND2_X1 U7374 ( .A1(n5928), .A2(n5929), .ZN(n5809) );
  INV_X1 U7375 ( .A(n8429), .ZN(n5994) );
  NAND2_X1 U7376 ( .A1(n5807), .A2(n5994), .ZN(n5808) );
  NAND2_X1 U7377 ( .A1(n5809), .A2(n5808), .ZN(n6029) );
  OR2_X1 U7378 ( .A1(n6564), .A2(n7994), .ZN(n5812) );
  OR2_X1 U7379 ( .A1(n7874), .A2(n4850), .ZN(n5811) );
  XNOR2_X1 U7380 ( .A(n6033), .B(n6355), .ZN(n6030) );
  NAND2_X1 U7381 ( .A1(n7903), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5817) );
  INV_X1 U7382 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5813) );
  OR2_X1 U7383 ( .A1(n7841), .A2(n5813), .ZN(n5816) );
  OR2_X1 U7384 ( .A1(n7288), .A2(n9093), .ZN(n5815) );
  OR2_X1 U7385 ( .A1(n6581), .A2(n4697), .ZN(n5814) );
  XNOR2_X1 U7386 ( .A(n6030), .B(n8428), .ZN(n6028) );
  XOR2_X1 U7387 ( .A(n6029), .B(n6028), .Z(n5845) );
  OR2_X1 U7388 ( .A1(n6087), .A2(n10352), .ZN(n5818) );
  NOR2_X1 U7389 ( .A1(n6177), .A2(n5819), .ZN(n7984) );
  OR2_X1 U7390 ( .A1(n8512), .A2(n5820), .ZN(n5821) );
  NAND3_X1 U7391 ( .A1(n7984), .A2(n5838), .A3(n5873), .ZN(n8404) );
  NAND3_X1 U7392 ( .A1(n7984), .A2(n5838), .A3(n5872), .ZN(n8382) );
  INV_X1 U7393 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5822) );
  INV_X1 U7394 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5823) );
  OR2_X1 U7395 ( .A1(n7288), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5826) );
  OR2_X1 U7396 ( .A1(n6581), .A2(n5824), .ZN(n5825) );
  INV_X1 U7397 ( .A(n8427), .ZN(n6114) );
  OAI22_X1 U7398 ( .A1(n5994), .A2(n8404), .B1(n8382), .B2(n6114), .ZN(n5843)
         );
  INV_X1 U7399 ( .A(n5866), .ZN(n6185) );
  NAND2_X1 U7400 ( .A1(n5829), .A2(n10183), .ZN(n6082) );
  NAND2_X1 U7401 ( .A1(n6082), .A2(n5830), .ZN(n5836) );
  INV_X1 U7402 ( .A(n5831), .ZN(n5832) );
  AND3_X1 U7403 ( .A1(n5888), .A2(n5834), .A3(n5833), .ZN(n5835) );
  OAI211_X1 U7404 ( .C1(n5838), .C2(n6085), .A(n5836), .B(n5835), .ZN(n5837)
         );
  NAND2_X1 U7405 ( .A1(n5837), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5841) );
  INV_X1 U7406 ( .A(n5838), .ZN(n5839) );
  NAND2_X1 U7407 ( .A1(n7984), .A2(n5839), .ZN(n5840) );
  NOR2_X1 U7408 ( .A1(n8406), .A2(P2_U3151), .ZN(n6000) );
  NOR2_X1 U7409 ( .A1(n6000), .A2(n9093), .ZN(n5842) );
  AOI211_X1 U7410 ( .C1(n6355), .C2(n8390), .A(n5843), .B(n5842), .ZN(n5844)
         );
  OAI21_X1 U7411 ( .B1(n8394), .B2(n5845), .A(n5844), .ZN(P2_U3177) );
  NAND2_X1 U7412 ( .A1(n5846), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5848) );
  INV_X1 U7413 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5847) );
  XNOR2_X1 U7414 ( .A(n5848), .B(n5847), .ZN(n7500) );
  OAI222_X1 U7415 ( .A1(n8278), .A2(n5850), .B1(n10173), .B2(n5849), .C1(n7500), .C2(P1_U3086), .ZN(P1_U3340) );
  AOI21_X1 U7416 ( .B1(n6644), .B2(P1_REG1_REG_10__SCAN_IN), .A(n5851), .ZN(
        n5854) );
  INV_X1 U7417 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n5852) );
  MUX2_X1 U7418 ( .A(n5852), .B(P1_REG1_REG_11__SCAN_IN), .S(n6648), .Z(n5853)
         );
  NOR2_X1 U7419 ( .A1(n5854), .A2(n5853), .ZN(n6068) );
  AOI211_X1 U7420 ( .C1(n5854), .C2(n5853), .A(n9751), .B(n6068), .ZN(n5863)
         );
  NAND2_X1 U7421 ( .A1(n6648), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5856) );
  OAI21_X1 U7422 ( .B1(n6648), .B2(P1_REG2_REG_11__SCAN_IN), .A(n5856), .ZN(
        n5857) );
  AOI211_X1 U7423 ( .C1(n5858), .C2(n5857), .A(n9752), .B(n6075), .ZN(n5862)
         );
  INV_X1 U7424 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n5860) );
  NAND2_X1 U7425 ( .A1(n9755), .A2(n6648), .ZN(n5859) );
  NAND2_X1 U7426 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n7028) );
  OAI211_X1 U7427 ( .C1(n5860), .C2(n9761), .A(n5859), .B(n7028), .ZN(n5861)
         );
  OR3_X1 U7428 ( .A1(n5863), .A2(n5862), .A3(n5861), .ZN(P1_U3254) );
  INV_X1 U7429 ( .A(n7986), .ZN(n7646) );
  AOI21_X1 U7430 ( .B1(n7977), .B2(n7646), .A(n7981), .ZN(n5864) );
  AND2_X1 U7431 ( .A1(n10352), .A2(n5864), .ZN(n5865) );
  NOR2_X1 U7432 ( .A1(n5866), .A2(n7986), .ZN(n10318) );
  INV_X1 U7433 ( .A(n10318), .ZN(n10344) );
  OR2_X1 U7434 ( .A1(n8429), .A2(n10300), .ZN(n7651) );
  NAND2_X1 U7435 ( .A1(n8429), .A2(n10300), .ZN(n7649) );
  NOR2_X1 U7436 ( .A1(n8430), .A2(n5995), .ZN(n6351) );
  NAND2_X1 U7437 ( .A1(n6350), .A2(n7651), .ZN(n5867) );
  NAND2_X1 U7438 ( .A1(n5867), .A2(n7914), .ZN(n6359) );
  OAI21_X1 U7439 ( .B1(n5867), .B2(n7914), .A(n6359), .ZN(n6184) );
  INV_X1 U7440 ( .A(n7914), .ZN(n7656) );
  AND2_X1 U7441 ( .A1(n8430), .A2(n10299), .ZN(n6344) );
  OAI22_X1 U7442 ( .A1(n7916), .A2(n6344), .B1(n5868), .B2(n8429), .ZN(n6354)
         );
  XNOR2_X1 U7443 ( .A(n7656), .B(n6354), .ZN(n5871) );
  NAND2_X1 U7444 ( .A1(n7973), .A2(n7977), .ZN(n5870) );
  NAND2_X1 U7445 ( .A1(n5871), .A2(n8706), .ZN(n5875) );
  AOI22_X1 U7446 ( .A1(n8701), .A2(n8429), .B1(n8427), .B2(n8703), .ZN(n5874)
         );
  NAND2_X1 U7447 ( .A1(n5875), .A2(n5874), .ZN(n6187) );
  AOI21_X1 U7448 ( .B1(n10358), .B2(n6184), .A(n6187), .ZN(n6092) );
  NAND3_X1 U7449 ( .A1(n7977), .A2(n7986), .A3(n8523), .ZN(n5876) );
  NAND2_X1 U7450 ( .A1(n7893), .A2(n5876), .ZN(n5879) );
  OR2_X1 U7451 ( .A1(n5879), .A2(n5877), .ZN(n5881) );
  NAND2_X1 U7452 ( .A1(n5879), .A2(n5878), .ZN(n5880) );
  INV_X1 U7453 ( .A(n5882), .ZN(n5884) );
  AND2_X1 U7454 ( .A1(n5884), .A2(n5883), .ZN(n5889) );
  AND2_X1 U7455 ( .A1(n5886), .A2(n5885), .ZN(n5887) );
  NAND2_X1 U7456 ( .A1(n10381), .A2(n10363), .ZN(n8752) );
  INV_X1 U7457 ( .A(n6355), .ZN(n7661) );
  OAI22_X1 U7458 ( .A1(n8752), .A2(n7661), .B1(n10381), .B2(n4697), .ZN(n5890)
         );
  INV_X1 U7459 ( .A(n5890), .ZN(n5891) );
  OAI21_X1 U7460 ( .B1(n6092), .B2(n10378), .A(n5891), .ZN(P2_U3461) );
  NAND2_X1 U7461 ( .A1(n6804), .A2(n6339), .ZN(n5892) );
  NAND2_X1 U7462 ( .A1(n5893), .A2(n5892), .ZN(n6469) );
  NAND2_X1 U7463 ( .A1(n5895), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5897) );
  NAND2_X1 U7464 ( .A1(n8043), .A2(n9685), .ZN(n5896) );
  OAI211_X1 U7465 ( .C1(n5894), .C2(n5898), .A(n5897), .B(n5896), .ZN(n5899)
         );
  NAND2_X1 U7466 ( .A1(n6254), .A2(n5899), .ZN(n9377) );
  INV_X1 U7467 ( .A(n5899), .ZN(n10247) );
  NAND2_X1 U7468 ( .A1(n5742), .A2(n10247), .ZN(n9541) );
  NAND2_X1 U7469 ( .A1(n9377), .A2(n9541), .ZN(n6468) );
  NAND2_X1 U7470 ( .A1(n6254), .A2(n10247), .ZN(n5900) );
  NAND2_X1 U7471 ( .A1(n6467), .A2(n5900), .ZN(n5910) );
  NAND2_X1 U7472 ( .A1(n5901), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5914) );
  OAI21_X1 U7473 ( .B1(n5901), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5914), .ZN(
        n6267) );
  INV_X1 U7474 ( .A(n6267), .ZN(n6697) );
  NAND2_X1 U7475 ( .A1(n5720), .A2(n6697), .ZN(n5905) );
  NAND2_X1 U7476 ( .A1(n9476), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5904) );
  NAND2_X1 U7477 ( .A1(n5599), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5903) );
  NAND2_X1 U7478 ( .A1(n4491), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5902) );
  NAND2_X1 U7479 ( .A1(n9473), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5908) );
  NAND2_X1 U7480 ( .A1(n4494), .A2(n5906), .ZN(n5907) );
  OAI211_X1 U7481 ( .C1(n5894), .C2(n5909), .A(n5908), .B(n5907), .ZN(n5911)
         );
  NAND2_X1 U7482 ( .A1(n8270), .A2(n5911), .ZN(n9379) );
  NAND2_X1 U7483 ( .A1(n9638), .A2(n6700), .ZN(n9543) );
  NAND2_X1 U7484 ( .A1(n9379), .A2(n9543), .ZN(n6220) );
  OAI21_X1 U7485 ( .B1(n5910), .B2(n6220), .A(n6193), .ZN(n6702) );
  OR2_X1 U7486 ( .A1(n5912), .A2(n5899), .ZN(n6470) );
  AOI211_X1 U7487 ( .C1(n5911), .C2(n6470), .A(n10266), .B(n6431), .ZN(n6696)
         );
  NAND2_X1 U7488 ( .A1(n9476), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5919) );
  INV_X1 U7489 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5913) );
  NOR2_X1 U7490 ( .A1(n5914), .A2(n5913), .ZN(n6200) );
  AND2_X1 U7491 ( .A1(n5914), .A2(n5913), .ZN(n5915) );
  NOR2_X1 U7492 ( .A1(n6200), .A2(n5915), .ZN(n6434) );
  NAND2_X1 U7493 ( .A1(n5720), .A2(n6434), .ZN(n5918) );
  NAND2_X1 U7494 ( .A1(n5599), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5917) );
  NAND2_X1 U7495 ( .A1(n4491), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5916) );
  NAND2_X1 U7496 ( .A1(n9371), .A2(n9538), .ZN(n6465) );
  INV_X1 U7497 ( .A(n6468), .ZN(n9494) );
  NAND2_X1 U7498 ( .A1(n6465), .A2(n9494), .ZN(n6464) );
  NAND2_X1 U7499 ( .A1(n6464), .A2(n9377), .ZN(n6221) );
  XNOR2_X1 U7500 ( .A(n6221), .B(n6220), .ZN(n5920) );
  OAI222_X1 U7501 ( .A1(n10013), .A2(n6365), .B1(n10011), .B2(n6254), .C1(
        n5920), .C2(n9938), .ZN(n6695) );
  AOI211_X1 U7502 ( .C1(n10276), .C2(n6702), .A(n6696), .B(n6695), .ZN(n5927)
         );
  INV_X1 U7503 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5921) );
  OAI22_X1 U7504 ( .A1(n10164), .A2(n6700), .B1(n10280), .B2(n5921), .ZN(n5922) );
  INV_X1 U7505 ( .A(n5922), .ZN(n5923) );
  OAI21_X1 U7506 ( .B1(n5927), .B2(n10278), .A(n5923), .ZN(P1_U3468) );
  INV_X1 U7507 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5924) );
  OAI22_X1 U7508 ( .A1(n10108), .A2(n6700), .B1(n10293), .B2(n5924), .ZN(n5925) );
  INV_X1 U7509 ( .A(n5925), .ZN(n5926) );
  OAI21_X1 U7510 ( .B1(n5927), .B2(n10290), .A(n5926), .ZN(P1_U3527) );
  XOR2_X1 U7511 ( .A(n5929), .B(n5928), .Z(n5935) );
  INV_X1 U7512 ( .A(n8428), .ZN(n6053) );
  INV_X1 U7513 ( .A(n8430), .ZN(n5930) );
  OAI22_X1 U7514 ( .A1(n6053), .A2(n8382), .B1(n8404), .B2(n5930), .ZN(n5933)
         );
  NOR2_X1 U7515 ( .A1(n6000), .A2(n5931), .ZN(n5932) );
  AOI211_X1 U7516 ( .C1(n5868), .C2(n8390), .A(n5933), .B(n5932), .ZN(n5934)
         );
  OAI21_X1 U7517 ( .B1(n8394), .B2(n5935), .A(n5934), .ZN(P2_U3162) );
  AOI21_X1 U7518 ( .B1(n5952), .B2(P2_REG1_REG_6__SCAN_IN), .A(n5936), .ZN(
        n6002) );
  INV_X1 U7519 ( .A(n6002), .ZN(n5937) );
  XNOR2_X1 U7520 ( .A(n5937), .B(n5953), .ZN(n6001) );
  XNOR2_X1 U7521 ( .A(n6001), .B(P2_REG1_REG_7__SCAN_IN), .ZN(n5958) );
  INV_X1 U7522 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n5938) );
  INV_X1 U7523 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8866) );
  OR2_X1 U7524 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8866), .ZN(n6779) );
  OAI21_X1 U7525 ( .B1(n5939), .B2(n5938), .A(n6779), .ZN(n5950) );
  NAND2_X1 U7526 ( .A1(n5947), .A2(n5946), .ZN(n5944) );
  INV_X1 U7527 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6929) );
  INV_X1 U7528 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6580) );
  MUX2_X1 U7529 ( .A(n6929), .B(n6580), .S(n8512), .Z(n5940) );
  NAND2_X1 U7530 ( .A1(n5940), .A2(n6573), .ZN(n6021) );
  INV_X1 U7531 ( .A(n5940), .ZN(n5941) );
  NAND2_X1 U7532 ( .A1(n5941), .A2(n5953), .ZN(n5942) );
  NAND2_X1 U7533 ( .A1(n6021), .A2(n5942), .ZN(n5945) );
  INV_X1 U7534 ( .A(n5945), .ZN(n5943) );
  NAND2_X1 U7535 ( .A1(n5944), .A2(n5943), .ZN(n6022) );
  NAND3_X1 U7536 ( .A1(n5947), .A2(n5946), .A3(n5945), .ZN(n5948) );
  AOI21_X1 U7537 ( .B1(n6022), .B2(n5948), .A(n8517), .ZN(n5949) );
  AOI211_X1 U7538 ( .C1(n8448), .C2(n6573), .A(n5950), .B(n5949), .ZN(n5957)
         );
  AOI21_X1 U7539 ( .B1(n5952), .B2(P2_REG2_REG_6__SCAN_IN), .A(n5951), .ZN(
        n6006) );
  INV_X1 U7540 ( .A(n6006), .ZN(n5954) );
  XNOR2_X1 U7541 ( .A(n6005), .B(n6929), .ZN(n5955) );
  NAND2_X1 U7542 ( .A1(n5955), .A2(n8526), .ZN(n5956) );
  OAI211_X1 U7543 ( .C1(n5958), .C2(n8529), .A(n5957), .B(n5956), .ZN(P2_U3189) );
  AND2_X1 U7544 ( .A1(n5960), .A2(n5959), .ZN(n5961) );
  NAND2_X1 U7545 ( .A1(n5962), .A2(n5961), .ZN(n5966) );
  INV_X1 U7546 ( .A(n5963), .ZN(n5964) );
  NAND2_X1 U7547 ( .A1(n5964), .A2(SI_15_), .ZN(n5965) );
  MUX2_X1 U7548 ( .A(n5976), .B(n8877), .S(n7901), .Z(n5968) );
  INV_X1 U7549 ( .A(SI_16_), .ZN(n5967) );
  NAND2_X1 U7550 ( .A1(n5968), .A2(n5967), .ZN(n5981) );
  INV_X1 U7551 ( .A(n5968), .ZN(n5969) );
  NAND2_X1 U7552 ( .A1(n5969), .A2(SI_16_), .ZN(n5970) );
  NAND2_X1 U7553 ( .A1(n5981), .A2(n5970), .ZN(n5982) );
  XNOR2_X1 U7554 ( .A(n5983), .B(n5982), .ZN(n7465) );
  INV_X1 U7555 ( .A(n7465), .ZN(n5980) );
  NAND2_X1 U7556 ( .A1(n5971), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5972) );
  NAND2_X1 U7557 ( .A1(n5973), .A2(n5972), .ZN(n5974) );
  NAND2_X1 U7558 ( .A1(n5974), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5975) );
  INV_X1 U7559 ( .A(n8458), .ZN(n7538) );
  OAI222_X1 U7560 ( .A1(n9222), .A2(n5976), .B1(n9220), .B2(n5980), .C1(
        P2_U3151), .C2(n7538), .ZN(P2_U3279) );
  OR2_X1 U7561 ( .A1(n5233), .A2(n5977), .ZN(n5978) );
  NAND2_X1 U7562 ( .A1(n5978), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5979) );
  XNOR2_X1 U7563 ( .A(n5979), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7584) );
  INV_X1 U7564 ( .A(n7584), .ZN(n7496) );
  OAI222_X1 U7565 ( .A1(n8278), .A2(n8877), .B1(n10173), .B2(n5980), .C1(
        P1_U3086), .C2(n7496), .ZN(P1_U3339) );
  MUX2_X1 U7566 ( .A(n5990), .B(n5992), .S(n7901), .Z(n5985) );
  NAND2_X1 U7567 ( .A1(n5985), .A2(n5984), .ZN(n6060) );
  INV_X1 U7568 ( .A(n5985), .ZN(n5986) );
  NAND2_X1 U7569 ( .A1(n5986), .A2(SI_17_), .ZN(n5987) );
  XNOR2_X1 U7570 ( .A(n6059), .B(n6058), .ZN(n8023) );
  INV_X1 U7571 ( .A(n8023), .ZN(n5993) );
  NAND2_X1 U7572 ( .A1(n5988), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5989) );
  XNOR2_X1 U7573 ( .A(n5989), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8477) );
  OAI222_X1 U7574 ( .A1(n7594), .A2(n5993), .B1(n8493), .B2(P2_U3151), .C1(
        n5990), .C2(n9222), .ZN(P2_U3278) );
  XNOR2_X1 U7575 ( .A(n5991), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9735) );
  INV_X1 U7576 ( .A(n9735), .ZN(n7508) );
  OAI222_X1 U7577 ( .A1(P1_U3086), .A2(n7508), .B1(n10173), .B2(n5993), .C1(
        n5992), .C2(n8278), .ZN(P1_U3338) );
  NAND2_X1 U7578 ( .A1(n8430), .A2(n5995), .ZN(n7653) );
  AND2_X1 U7579 ( .A1(n7648), .A2(n7653), .ZN(n10295) );
  INV_X1 U7580 ( .A(n10295), .ZN(n5997) );
  OAI22_X1 U7581 ( .A1(n8410), .A2(n5995), .B1(n5994), .B2(n8382), .ZN(n5996)
         );
  AOI21_X1 U7582 ( .B1(n5997), .B2(n8302), .A(n5996), .ZN(n5998) );
  OAI21_X1 U7583 ( .B1(n6000), .B2(n5999), .A(n5998), .ZN(P2_U3172) );
  MUX2_X1 U7584 ( .A(n6012), .B(P2_REG1_REG_8__SCAN_IN), .S(n6570), .Z(n6004)
         );
  OAI21_X1 U7585 ( .B1(n6004), .B2(n6003), .A(n6146), .ZN(n6026) );
  MUX2_X1 U7586 ( .A(n6013), .B(P2_REG2_REG_8__SCAN_IN), .S(n6570), .Z(n6008)
         );
  OAI21_X1 U7587 ( .B1(n6008), .B2(n6007), .A(n6137), .ZN(n6009) );
  NAND2_X1 U7588 ( .A1(n6009), .A2(n8526), .ZN(n6011) );
  AND2_X1 U7589 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6970) );
  AOI21_X1 U7590 ( .B1(n8519), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6970), .ZN(
        n6010) );
  OAI211_X1 U7591 ( .C1(n8522), .C2(n6015), .A(n6011), .B(n6010), .ZN(n6025)
         );
  NAND2_X1 U7592 ( .A1(n6022), .A2(n6021), .ZN(n6019) );
  MUX2_X1 U7593 ( .A(n6013), .B(n6012), .S(n8512), .Z(n6014) );
  NAND2_X1 U7594 ( .A1(n6014), .A2(n6570), .ZN(n6160) );
  INV_X1 U7595 ( .A(n6014), .ZN(n6016) );
  NAND2_X1 U7596 ( .A1(n6016), .A2(n6015), .ZN(n6017) );
  NAND2_X1 U7597 ( .A1(n6160), .A2(n6017), .ZN(n6020) );
  INV_X1 U7598 ( .A(n6020), .ZN(n6018) );
  NAND2_X1 U7599 ( .A1(n6019), .A2(n6018), .ZN(n6161) );
  NAND3_X1 U7600 ( .A1(n6022), .A2(n6021), .A3(n6020), .ZN(n6023) );
  AOI21_X1 U7601 ( .B1(n6161), .B2(n6023), .A(n8517), .ZN(n6024) );
  AOI211_X1 U7602 ( .C1(n8442), .C2(n6026), .A(n6025), .B(n6024), .ZN(n6027)
         );
  INV_X1 U7603 ( .A(n6027), .ZN(P2_U3190) );
  INV_X1 U7604 ( .A(n8406), .ZN(n8291) );
  NAND2_X1 U7605 ( .A1(n6029), .A2(n6028), .ZN(n6032) );
  NAND2_X1 U7606 ( .A1(n6030), .A2(n6053), .ZN(n6031) );
  NAND2_X1 U7607 ( .A1(n6032), .A2(n6031), .ZN(n6040) );
  INV_X2 U7608 ( .A(n6033), .ZN(n8139) );
  INV_X1 U7609 ( .A(n8139), .ZN(n6238) );
  OR2_X1 U7610 ( .A1(n6564), .A2(n5715), .ZN(n6038) );
  OR2_X1 U7611 ( .A1(n7874), .A2(n6034), .ZN(n6037) );
  NAND2_X1 U7612 ( .A1(n7736), .A2(n6035), .ZN(n6036) );
  XNOR2_X1 U7613 ( .A(n6238), .B(n10306), .ZN(n6097) );
  XNOR2_X1 U7614 ( .A(n6097), .B(n8427), .ZN(n6039) );
  AOI21_X1 U7615 ( .B1(n6040), .B2(n6039), .A(n8394), .ZN(n6041) );
  NAND2_X1 U7616 ( .A1(n6041), .A2(n6099), .ZN(n6057) );
  INV_X1 U7617 ( .A(n10306), .ZN(n6481) );
  AND2_X1 U7618 ( .A1(n8390), .A2(n6481), .ZN(n6055) );
  NAND2_X1 U7619 ( .A1(n4814), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6048) );
  OR2_X1 U7620 ( .A1(n7865), .A2(n6042), .ZN(n6047) );
  OR2_X1 U7621 ( .A1(n6581), .A2(n6043), .ZN(n6046) );
  AND2_X1 U7622 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6044) );
  NOR2_X1 U7623 ( .A1(n6105), .A2(n6044), .ZN(n6478) );
  OR2_X1 U7624 ( .A1(n7288), .A2(n6478), .ZN(n6045) );
  NAND4_X1 U7625 ( .A1(n6048), .A2(n6047), .A3(n6046), .A4(n6045), .ZN(n8426)
         );
  INV_X1 U7626 ( .A(n8426), .ZN(n6049) );
  OR2_X1 U7627 ( .A1(n8382), .A2(n6049), .ZN(n6052) );
  INV_X1 U7628 ( .A(n6050), .ZN(n6051) );
  OAI211_X1 U7629 ( .C1(n8404), .C2(n6053), .A(n6052), .B(n6051), .ZN(n6054)
         );
  NOR2_X1 U7630 ( .A1(n6055), .A2(n6054), .ZN(n6056) );
  OAI211_X1 U7631 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8291), .A(n6057), .B(
        n6056), .ZN(P2_U3158) );
  INV_X1 U7632 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6061) );
  MUX2_X1 U7633 ( .A(n6122), .B(n6061), .S(n7901), .Z(n6290) );
  XNOR2_X1 U7634 ( .A(n6290), .B(SI_18_), .ZN(n6289) );
  XNOR2_X1 U7635 ( .A(n6293), .B(n6289), .ZN(n8029) );
  INV_X1 U7636 ( .A(n8029), .ZN(n6121) );
  NAND2_X1 U7637 ( .A1(n6062), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6064) );
  OR2_X1 U7638 ( .A1(n6064), .A2(n6063), .ZN(n6066) );
  NAND2_X1 U7639 ( .A1(n6064), .A2(n6063), .ZN(n6065) );
  AND2_X1 U7640 ( .A1(n6066), .A2(n6065), .ZN(n9738) );
  AOI22_X1 U7641 ( .A1(n9738), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10171), .ZN(n6067) );
  OAI21_X1 U7642 ( .B1(n6121), .B2(n10173), .A(n6067), .ZN(P1_U3337) );
  AOI21_X1 U7643 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n6648), .A(n6068), .ZN(
        n6070) );
  MUX2_X1 U7644 ( .A(n10291), .B(P1_REG1_REG_12__SCAN_IN), .S(n7150), .Z(n6069) );
  NAND2_X1 U7645 ( .A1(n6070), .A2(n6069), .ZN(n7148) );
  OAI21_X1 U7646 ( .B1(n6070), .B2(n6069), .A(n7148), .ZN(n6074) );
  INV_X1 U7647 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n6072) );
  INV_X1 U7648 ( .A(n7150), .ZN(n6657) );
  NAND2_X1 U7649 ( .A1(n9755), .A2(n6657), .ZN(n6071) );
  NAND2_X1 U7650 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n7235) );
  OAI211_X1 U7651 ( .C1(n6072), .C2(n9761), .A(n6071), .B(n7235), .ZN(n6073)
         );
  AOI21_X1 U7652 ( .B1(n6074), .B2(n9756), .A(n6073), .ZN(n6081) );
  NOR2_X1 U7653 ( .A1(n6657), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6076) );
  AOI21_X1 U7654 ( .B1(n6657), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6076), .ZN(
        n6077) );
  OAI21_X1 U7655 ( .B1(n6078), .B2(n6077), .A(n7140), .ZN(n6079) );
  NAND2_X1 U7656 ( .A1(n6079), .A2(n9740), .ZN(n6080) );
  NAND2_X1 U7657 ( .A1(n6081), .A2(n6080), .ZN(P1_U3255) );
  INV_X1 U7658 ( .A(n6082), .ZN(n6084) );
  AND2_X1 U7659 ( .A1(n6177), .A2(n6085), .ZN(n6086) );
  OAI22_X1 U7660 ( .A1(n9178), .A2(n7661), .B1(n5813), .B2(n10364), .ZN(n6090)
         );
  INV_X1 U7661 ( .A(n6090), .ZN(n6091) );
  OAI21_X1 U7662 ( .B1(n6092), .B2(n10366), .A(n6091), .ZN(P2_U3396) );
  OR2_X1 U7663 ( .A1(n6564), .A2(n5898), .ZN(n6096) );
  OR2_X1 U7664 ( .A1(n7874), .A2(n6093), .ZN(n6095) );
  NAND2_X1 U7665 ( .A1(n7736), .A2(n8447), .ZN(n6094) );
  XNOR2_X1 U7666 ( .A(n6238), .B(n10309), .ZN(n6230) );
  XNOR2_X1 U7667 ( .A(n6230), .B(n8426), .ZN(n6102) );
  NAND2_X1 U7668 ( .A1(n6097), .A2(n8427), .ZN(n6098) );
  INV_X1 U7669 ( .A(n6232), .ZN(n6100) );
  AOI21_X1 U7670 ( .B1(n6102), .B2(n6101), .A(n6100), .ZN(n6118) );
  INV_X1 U7671 ( .A(n10309), .ZN(n6498) );
  NAND2_X1 U7672 ( .A1(n7903), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6111) );
  INV_X1 U7673 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6103) );
  OR2_X1 U7674 ( .A1(n7841), .A2(n6103), .ZN(n6110) );
  OR2_X1 U7675 ( .A1(n6105), .A2(n6104), .ZN(n6106) );
  AND2_X1 U7676 ( .A1(n6240), .A2(n6106), .ZN(n6505) );
  OR2_X1 U7677 ( .A1(n7288), .A2(n6505), .ZN(n6109) );
  OR2_X1 U7678 ( .A1(n6581), .A2(n6107), .ZN(n6108) );
  NAND4_X1 U7679 ( .A1(n6111), .A2(n6110), .A3(n6109), .A4(n6108), .ZN(n8425)
         );
  INV_X1 U7680 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6112) );
  NOR2_X1 U7681 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6112), .ZN(n8440) );
  AOI21_X1 U7682 ( .B1(n8402), .B2(n8425), .A(n8440), .ZN(n6113) );
  OAI21_X1 U7683 ( .B1(n6114), .B2(n8404), .A(n6113), .ZN(n6116) );
  NOR2_X1 U7684 ( .A1(n8291), .A2(n6478), .ZN(n6115) );
  AOI211_X1 U7685 ( .C1(n6498), .C2(n8390), .A(n6116), .B(n6115), .ZN(n6117)
         );
  OAI21_X1 U7686 ( .B1(n6118), .B2(n8394), .A(n6117), .ZN(P2_U3170) );
  NAND2_X1 U7687 ( .A1(n6119), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6120) );
  XNOR2_X1 U7688 ( .A(n6120), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8495) );
  INV_X1 U7689 ( .A(n8495), .ZN(n8508) );
  OAI222_X1 U7690 ( .A1(n9222), .A2(n6122), .B1(n8508), .B2(P2_U3151), .C1(
        n7594), .C2(n6121), .ZN(P2_U3277) );
  NAND2_X1 U7691 ( .A1(n6161), .A2(n6160), .ZN(n6128) );
  MUX2_X1 U7692 ( .A(n6624), .B(n6123), .S(n8512), .Z(n6124) );
  NAND2_X1 U7693 ( .A1(n6124), .A2(n6588), .ZN(n6135) );
  INV_X1 U7694 ( .A(n6124), .ZN(n6125) );
  NAND2_X1 U7695 ( .A1(n6125), .A2(n6158), .ZN(n6126) );
  NAND2_X1 U7696 ( .A1(n6135), .A2(n6126), .ZN(n6159) );
  INV_X1 U7697 ( .A(n6159), .ZN(n6127) );
  NAND2_X1 U7698 ( .A1(n6128), .A2(n6127), .ZN(n6163) );
  NAND2_X1 U7699 ( .A1(n6163), .A2(n6135), .ZN(n6133) );
  INV_X1 U7700 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6612) );
  INV_X1 U7701 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6613) );
  MUX2_X1 U7702 ( .A(n6612), .B(n6613), .S(n8512), .Z(n6129) );
  NAND2_X1 U7703 ( .A1(n6129), .A2(n6723), .ZN(n6390) );
  INV_X1 U7704 ( .A(n6129), .ZN(n6130) );
  NAND2_X1 U7705 ( .A1(n6130), .A2(n6145), .ZN(n6131) );
  NAND2_X1 U7706 ( .A1(n6390), .A2(n6131), .ZN(n6134) );
  INV_X1 U7707 ( .A(n6134), .ZN(n6132) );
  NAND2_X1 U7708 ( .A1(n6133), .A2(n6132), .ZN(n6391) );
  NAND3_X1 U7709 ( .A1(n6163), .A2(n6135), .A3(n6134), .ZN(n6136) );
  AND2_X1 U7710 ( .A1(n6391), .A2(n6136), .ZN(n6154) );
  AOI22_X1 U7711 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n6145), .B1(n6723), .B2(
        n6612), .ZN(n6141) );
  NAND2_X1 U7712 ( .A1(n6138), .A2(n6158), .ZN(n6139) );
  XNOR2_X1 U7713 ( .A(n6138), .B(n6588), .ZN(n6156) );
  NAND2_X1 U7714 ( .A1(P2_REG2_REG_9__SCAN_IN), .A2(n6156), .ZN(n6155) );
  OAI21_X1 U7715 ( .B1(n6141), .B2(n6140), .A(n6393), .ZN(n6144) );
  NAND2_X1 U7716 ( .A1(n8519), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n6142) );
  NAND2_X1 U7717 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7129) );
  OAI211_X1 U7718 ( .C1(n8522), .C2(n6145), .A(n6142), .B(n7129), .ZN(n6143)
         );
  AOI21_X1 U7719 ( .B1(n6144), .B2(n8526), .A(n6143), .ZN(n6153) );
  AOI22_X1 U7720 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n6145), .B1(n6723), .B2(
        n6613), .ZN(n6150) );
  NAND2_X1 U7721 ( .A1(n6147), .A2(n6158), .ZN(n6148) );
  NAND2_X1 U7722 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(n6168), .ZN(n6167) );
  OAI21_X1 U7723 ( .B1(n6150), .B2(n6149), .A(n6380), .ZN(n6151) );
  NAND2_X1 U7724 ( .A1(n6151), .A2(n8442), .ZN(n6152) );
  OAI211_X1 U7725 ( .C1(n6154), .C2(n8517), .A(n6153), .B(n6152), .ZN(P2_U3192) );
  OAI21_X1 U7726 ( .B1(n6156), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6155), .ZN(
        n6166) );
  NAND2_X1 U7727 ( .A1(n8519), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n6157) );
  NAND2_X1 U7728 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7433) );
  OAI211_X1 U7729 ( .C1(n8522), .C2(n6158), .A(n6157), .B(n7433), .ZN(n6165)
         );
  NAND3_X1 U7730 ( .A1(n6161), .A2(n6160), .A3(n6159), .ZN(n6162) );
  AOI21_X1 U7731 ( .B1(n6163), .B2(n6162), .A(n8517), .ZN(n6164) );
  AOI211_X1 U7732 ( .C1(n8526), .C2(n6166), .A(n6165), .B(n6164), .ZN(n6171)
         );
  OAI21_X1 U7733 ( .B1(n6168), .B2(P2_REG1_REG_9__SCAN_IN), .A(n6167), .ZN(
        n6169) );
  NAND2_X1 U7734 ( .A1(n6169), .A2(n8442), .ZN(n6170) );
  NAND2_X1 U7735 ( .A1(n6171), .A2(n6170), .ZN(P2_U3191) );
  INV_X1 U7736 ( .A(n6172), .ZN(n6176) );
  AND2_X1 U7737 ( .A1(n6174), .A2(n6173), .ZN(n6175) );
  NAND2_X1 U7738 ( .A1(n6177), .A2(n10352), .ZN(n6179) );
  NAND2_X1 U7739 ( .A1(n8429), .A2(n8703), .ZN(n10294) );
  NAND2_X1 U7740 ( .A1(n8709), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6178) );
  OAI211_X1 U7741 ( .C1(n10295), .C2(n6179), .A(n10294), .B(n6178), .ZN(n6181)
         );
  MUX2_X1 U7742 ( .A(n6181), .B(P2_REG2_REG_0__SCAN_IN), .S(n10198), .Z(n6182)
         );
  AOI21_X1 U7743 ( .B1(n8726), .B2(n10299), .A(n6182), .ZN(n6183) );
  INV_X1 U7744 ( .A(n6183), .ZN(P2_U3233) );
  INV_X1 U7745 ( .A(n6184), .ZN(n6191) );
  NAND2_X1 U7746 ( .A1(n6185), .A2(n7973), .ZN(n8570) );
  NAND2_X1 U7747 ( .A1(n10336), .A2(n8570), .ZN(n10196) );
  OAI22_X1 U7748 ( .A1(n10181), .A2(n9093), .B1(n7661), .B2(n10183), .ZN(n6186) );
  NOR2_X1 U7749 ( .A1(n6187), .A2(n6186), .ZN(n6188) );
  MUX2_X1 U7750 ( .A(n6189), .B(n6188), .S(n8724), .Z(n6190) );
  OAI21_X1 U7751 ( .B1(n6191), .B2(n8729), .A(n6190), .ZN(P2_U3231) );
  NAND2_X1 U7752 ( .A1(n8270), .A2(n6700), .ZN(n6192) );
  NAND2_X1 U7753 ( .A1(n6194), .A2(n9467), .ZN(n6196) );
  NAND2_X1 U7754 ( .A1(n9473), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n6195) );
  OAI211_X1 U7755 ( .C1(n5589), .C2(n6197), .A(n6196), .B(n6195), .ZN(n6198)
         );
  NAND2_X1 U7756 ( .A1(n6365), .A2(n6198), .ZN(n9382) );
  INV_X1 U7757 ( .A(n6365), .ZN(n9637) );
  NAND2_X1 U7758 ( .A1(n9637), .A2(n10254), .ZN(n9381) );
  NAND2_X1 U7759 ( .A1(n9382), .A2(n9381), .ZN(n6427) );
  NAND2_X1 U7760 ( .A1(n10254), .A2(n6365), .ZN(n6199) );
  NAND2_X1 U7761 ( .A1(n6200), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6214) );
  OR2_X1 U7762 ( .A1(n6200), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6201) );
  AND2_X1 U7763 ( .A1(n6214), .A2(n6201), .ZN(n6630) );
  NAND2_X1 U7764 ( .A1(n5720), .A2(n6630), .ZN(n6205) );
  NAND2_X1 U7765 ( .A1(n9476), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6204) );
  NAND2_X1 U7766 ( .A1(n4491), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6203) );
  NAND2_X1 U7767 ( .A1(n5599), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6202) );
  NAND2_X1 U7768 ( .A1(n6206), .A2(n9467), .ZN(n6209) );
  AOI22_X1 U7769 ( .A1(n9473), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n4494), .B2(
        n6207), .ZN(n6208) );
  NAND2_X1 U7770 ( .A1(n6209), .A2(n6208), .ZN(n6550) );
  NAND2_X1 U7771 ( .A1(n6549), .A2(n6550), .ZN(n6638) );
  NAND2_X1 U7772 ( .A1(n6633), .A2(n9636), .ZN(n6641) );
  NAND2_X1 U7773 ( .A1(n6638), .A2(n6641), .ZN(n9386) );
  NAND2_X1 U7774 ( .A1(n6210), .A2(n9386), .ZN(n6314) );
  OAI21_X1 U7775 ( .B1(n6210), .B2(n9386), .A(n6314), .ZN(n6635) );
  AND2_X1 U7776 ( .A1(n6431), .A2(n10254), .ZN(n6432) );
  INV_X1 U7777 ( .A(n6432), .ZN(n6212) );
  NAND2_X1 U7778 ( .A1(n6432), .A2(n6633), .ZN(n6320) );
  INV_X1 U7779 ( .A(n6320), .ZN(n6211) );
  AOI211_X1 U7780 ( .C1(n6550), .C2(n6212), .A(n10266), .B(n6211), .ZN(n6629)
         );
  NAND2_X1 U7781 ( .A1(n6214), .A2(n6213), .ZN(n6215) );
  AND2_X1 U7782 ( .A1(n6300), .A2(n6215), .ZN(n7040) );
  NAND2_X1 U7783 ( .A1(n5720), .A2(n7040), .ZN(n6219) );
  NAND2_X1 U7784 ( .A1(n9476), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6218) );
  NAND2_X1 U7785 ( .A1(n4492), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U7786 ( .A1(n5599), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6216) );
  INV_X1 U7787 ( .A(n6220), .ZN(n9493) );
  NAND2_X1 U7788 ( .A1(n6221), .A2(n9493), .ZN(n6222) );
  NAND2_X1 U7789 ( .A1(n6222), .A2(n9379), .ZN(n6640) );
  INV_X1 U7790 ( .A(n6427), .ZN(n6424) );
  NAND2_X1 U7791 ( .A1(n6640), .A2(n6424), .ZN(n6223) );
  NAND2_X1 U7792 ( .A1(n6223), .A2(n9382), .ZN(n6307) );
  XNOR2_X1 U7793 ( .A(n6307), .B(n9386), .ZN(n6224) );
  OAI222_X1 U7794 ( .A1(n10013), .A2(n7113), .B1(n10011), .B2(n6365), .C1(
        n6224), .C2(n9938), .ZN(n6628) );
  AOI211_X1 U7795 ( .C1(n10276), .C2(n6635), .A(n6629), .B(n6628), .ZN(n6229)
         );
  INV_X1 U7796 ( .A(n10108), .ZN(n6885) );
  AOI22_X1 U7797 ( .A1(n6885), .A2(n6550), .B1(n10290), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n6225) );
  OAI21_X1 U7798 ( .B1(n6229), .B2(n10290), .A(n6225), .ZN(P1_U3529) );
  INV_X1 U7799 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n6226) );
  OAI22_X1 U7800 ( .A1(n10164), .A2(n6633), .B1(n10280), .B2(n6226), .ZN(n6227) );
  INV_X1 U7801 ( .A(n6227), .ZN(n6228) );
  OAI21_X1 U7802 ( .B1(n6229), .B2(n10278), .A(n6228), .ZN(P1_U3474) );
  OR2_X1 U7803 ( .A1(n6230), .A2(n8426), .ZN(n6231) );
  OR2_X1 U7804 ( .A1(n5909), .A2(n6564), .ZN(n6237) );
  NAND2_X1 U7805 ( .A1(n7736), .A2(n6233), .ZN(n6236) );
  OR2_X1 U7806 ( .A1(n7874), .A2(n6234), .ZN(n6235) );
  XNOR2_X1 U7807 ( .A(n6238), .B(n10314), .ZN(n6768) );
  INV_X1 U7808 ( .A(n8425), .ZN(n6789) );
  XNOR2_X1 U7809 ( .A(n6768), .B(n6789), .ZN(n6766) );
  XOR2_X1 U7810 ( .A(n6767), .B(n6766), .Z(n6252) );
  INV_X1 U7811 ( .A(n10314), .ZN(n6508) );
  INV_X1 U7812 ( .A(n8404), .ZN(n8379) );
  NAND2_X1 U7813 ( .A1(n4814), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6246) );
  OR2_X1 U7814 ( .A1(n7865), .A2(n6239), .ZN(n6245) );
  NAND2_X1 U7815 ( .A1(n6240), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6241) );
  AND2_X1 U7816 ( .A1(n6577), .A2(n6241), .ZN(n6785) );
  OR2_X1 U7817 ( .A1(n7288), .A2(n6785), .ZN(n6244) );
  OR2_X1 U7818 ( .A1(n6581), .A2(n6242), .ZN(n6243) );
  NAND4_X1 U7819 ( .A1(n6246), .A2(n6245), .A3(n6244), .A4(n6243), .ZN(n8424)
         );
  INV_X1 U7820 ( .A(n8424), .ZN(n6778) );
  OAI21_X1 U7821 ( .B1(n8382), .B2(n6778), .A(n6247), .ZN(n6248) );
  AOI21_X1 U7822 ( .B1(n8379), .B2(n8426), .A(n6248), .ZN(n6249) );
  OAI21_X1 U7823 ( .B1(n6505), .B2(n8291), .A(n6249), .ZN(n6250) );
  AOI21_X1 U7824 ( .B1(n6508), .B2(n8390), .A(n6250), .ZN(n6251) );
  OAI21_X1 U7825 ( .B1(n6252), .B2(n8394), .A(n6251), .ZN(P2_U3167) );
  OAI22_X1 U7826 ( .A1(n8270), .A2(n5702), .B1(n6700), .B2(n8226), .ZN(n6266)
         );
  OAI22_X1 U7827 ( .A1(n6254), .A2(n8226), .B1(n10247), .B2(n5716), .ZN(n6253)
         );
  XNOR2_X1 U7828 ( .A(n6253), .B(n4495), .ZN(n6260) );
  OAI22_X1 U7829 ( .A1(n6254), .A2(n5702), .B1(n10247), .B2(n8226), .ZN(n6259)
         );
  XNOR2_X1 U7830 ( .A(n6260), .B(n6259), .ZN(n8266) );
  INV_X1 U7831 ( .A(n6255), .ZN(n6256) );
  NOR2_X1 U7832 ( .A1(n6257), .A2(n6256), .ZN(n8267) );
  AOI22_X1 U7833 ( .A1(n9638), .A2(n5521), .B1(n5911), .B2(n8208), .ZN(n6262)
         );
  XNOR2_X1 U7834 ( .A(n6262), .B(n4495), .ZN(n6263) );
  AOI21_X1 U7835 ( .B1(n6266), .B2(n6265), .A(n6371), .ZN(n6272) );
  OAI22_X1 U7836 ( .A1(n9314), .A2(n6267), .B1(n6365), .B2(n9345), .ZN(n6268)
         );
  AOI211_X1 U7837 ( .C1(n9334), .C2(n5742), .A(n6269), .B(n6268), .ZN(n6271)
         );
  NAND2_X1 U7838 ( .A1(n9363), .A2(n5911), .ZN(n6270) );
  OAI211_X1 U7839 ( .C1(n6272), .C2(n9365), .A(n6271), .B(n6270), .ZN(P1_U3227) );
  NAND4_X1 U7840 ( .A1(n6276), .A2(n6275), .A3(n6274), .A4(n6273), .ZN(n6277)
         );
  NOR2_X1 U7841 ( .A1(n6278), .A2(n9621), .ZN(n6318) );
  NAND2_X1 U7842 ( .A1(n10028), .A2(n6318), .ZN(n7343) );
  NAND2_X1 U7843 ( .A1(n6279), .A2(n10028), .ZN(n6287) );
  AND2_X2 U7844 ( .A1(n10028), .A2(n9621), .ZN(n10021) );
  INV_X1 U7845 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6280) );
  OAI22_X1 U7846 ( .A1(n10028), .A2(n6281), .B1(n6280), .B2(n9980), .ZN(n6284)
         );
  NAND2_X2 U7847 ( .A1(n10028), .A2(n6282), .ZN(n10026) );
  NOR2_X1 U7848 ( .A1(n10026), .A2(n5597), .ZN(n6283) );
  AOI211_X1 U7849 ( .C1(n6285), .C2(n10021), .A(n6284), .B(n6283), .ZN(n6286)
         );
  OAI211_X1 U7850 ( .C1(n6288), .C2(n7343), .A(n6287), .B(n6286), .ZN(P1_U3292) );
  INV_X1 U7851 ( .A(n6290), .ZN(n6291) );
  NAND2_X1 U7852 ( .A1(n6291), .A2(SI_18_), .ZN(n6292) );
  MUX2_X1 U7853 ( .A(n6298), .B(n8277), .S(n7901), .Z(n6295) );
  INV_X1 U7854 ( .A(SI_19_), .ZN(n6294) );
  NAND2_X1 U7855 ( .A1(n6295), .A2(n6294), .ZN(n6541) );
  INV_X1 U7856 ( .A(n6295), .ZN(n6296) );
  NAND2_X1 U7857 ( .A1(n6296), .A2(SI_19_), .ZN(n6297) );
  NAND2_X1 U7858 ( .A1(n6541), .A2(n6297), .ZN(n6539) );
  XNOR2_X1 U7859 ( .A(n6540), .B(n6539), .ZN(n8042) );
  INV_X1 U7860 ( .A(n8042), .ZN(n8276) );
  OAI222_X1 U7861 ( .A1(n9222), .A2(n6298), .B1(n9220), .B2(n8276), .C1(
        P2_U3151), .C2(n8523), .ZN(P2_U3276) );
  NAND2_X1 U7862 ( .A1(n9476), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6305) );
  AND2_X1 U7863 ( .A1(n6300), .A2(n6299), .ZN(n6301) );
  NOR2_X1 U7864 ( .A1(n6451), .A2(n6301), .ZN(n7112) );
  NAND2_X1 U7865 ( .A1(n5720), .A2(n7112), .ZN(n6304) );
  NAND2_X1 U7866 ( .A1(n9477), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6303) );
  NAND2_X1 U7867 ( .A1(n4491), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6302) );
  INV_X1 U7868 ( .A(n9386), .ZN(n6306) );
  NAND2_X1 U7869 ( .A1(n6307), .A2(n6306), .ZN(n6308) );
  NAND2_X1 U7870 ( .A1(n6308), .A2(n6638), .ZN(n6439) );
  NAND2_X1 U7871 ( .A1(n6569), .A2(n9467), .ZN(n6311) );
  AOI22_X1 U7872 ( .A1(n9473), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n4494), .B2(
        n6309), .ZN(n6310) );
  NAND2_X1 U7873 ( .A1(n6311), .A2(n6310), .ZN(n7002) );
  NAND2_X1 U7874 ( .A1(n6642), .A2(n6639), .ZN(n6315) );
  XNOR2_X1 U7875 ( .A(n6439), .B(n6315), .ZN(n6312) );
  OAI222_X1 U7876 ( .A1(n10013), .A2(n7041), .B1(n10011), .B2(n6549), .C1(
        n6312), .C2(n9938), .ZN(n6326) );
  INV_X1 U7877 ( .A(n6326), .ZN(n6325) );
  NAND2_X1 U7878 ( .A1(n6314), .A2(n6313), .ZN(n6316) );
  OAI21_X1 U7879 ( .B1(n6316), .B2(n6315), .A(n6448), .ZN(n6328) );
  INV_X1 U7880 ( .A(n7002), .ZN(n7047) );
  OR2_X1 U7881 ( .A1(n6320), .A2(n7002), .ZN(n6682) );
  INV_X1 U7882 ( .A(n6682), .ZN(n6319) );
  AOI211_X1 U7883 ( .C1(n7002), .C2(n6320), .A(n10266), .B(n6319), .ZN(n6327)
         );
  NAND2_X1 U7884 ( .A1(n6327), .A2(n10021), .ZN(n6322) );
  AOI22_X1 U7885 ( .A1(n9986), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7040), .B2(
        n10022), .ZN(n6321) );
  OAI211_X1 U7886 ( .C1(n7047), .C2(n10026), .A(n6322), .B(n6321), .ZN(n6323)
         );
  AOI21_X1 U7887 ( .B1(n6328), .B2(n9976), .A(n6323), .ZN(n6324) );
  OAI21_X1 U7888 ( .B1(n6325), .B2(n9986), .A(n6324), .ZN(P1_U3285) );
  AOI211_X1 U7889 ( .C1(n10276), .C2(n6328), .A(n6327), .B(n6326), .ZN(n6333)
         );
  INV_X1 U7890 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n6329) );
  OAI22_X1 U7891 ( .A1(n10164), .A2(n7047), .B1(n10280), .B2(n6329), .ZN(n6330) );
  INV_X1 U7892 ( .A(n6330), .ZN(n6331) );
  OAI21_X1 U7893 ( .B1(n6333), .B2(n10278), .A(n6331), .ZN(P1_U3477) );
  AOI22_X1 U7894 ( .A1(n6885), .A2(n7002), .B1(n10290), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n6332) );
  OAI21_X1 U7895 ( .B1(n6333), .B2(n10290), .A(n6332), .ZN(P1_U3530) );
  INV_X1 U7896 ( .A(n6334), .ZN(n6343) );
  NAND2_X1 U7897 ( .A1(n6335), .A2(n10021), .ZN(n6338) );
  AOI22_X1 U7898 ( .A1(n9986), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10022), .B2(
        n6336), .ZN(n6337) );
  OAI211_X1 U7899 ( .C1(n6339), .C2(n10026), .A(n6338), .B(n6337), .ZN(n6340)
         );
  AOI21_X1 U7900 ( .B1(n9976), .B2(n6341), .A(n6340), .ZN(n6342) );
  OAI21_X1 U7901 ( .B1(n6343), .B2(n9986), .A(n6342), .ZN(P1_U3290) );
  XNOR2_X1 U7902 ( .A(n7916), .B(n6344), .ZN(n6345) );
  NAND2_X1 U7903 ( .A1(n6345), .A2(n8706), .ZN(n6347) );
  AOI22_X1 U7904 ( .A1(n8703), .A2(n8428), .B1(n8430), .B2(n8701), .ZN(n6346)
         );
  NAND2_X1 U7905 ( .A1(n6347), .A2(n6346), .ZN(n10303) );
  AOI21_X1 U7906 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n8709), .A(n10303), .ZN(
        n6349) );
  MUX2_X1 U7907 ( .A(n6349), .B(n6348), .S(n10198), .Z(n6353) );
  OAI21_X1 U7908 ( .B1(n7916), .B2(n6351), .A(n6350), .ZN(n10304) );
  AOI22_X1 U7909 ( .A1(n8670), .A2(n10304), .B1(n5868), .B2(n8726), .ZN(n6352)
         );
  NAND2_X1 U7910 ( .A1(n6353), .A2(n6352), .ZN(P2_U3232) );
  NAND2_X1 U7911 ( .A1(n8427), .A2(n10306), .ZN(n7670) );
  NAND2_X1 U7912 ( .A1(n6354), .A2(n7656), .ZN(n6357) );
  OR2_X1 U7913 ( .A1(n8428), .A2(n6355), .ZN(n6356) );
  NAND2_X1 U7914 ( .A1(n6357), .A2(n6356), .ZN(n6480) );
  XOR2_X1 U7915 ( .A(n7915), .B(n6480), .Z(n6358) );
  AOI222_X1 U7916 ( .A1(n8706), .A2(n6358), .B1(n8428), .B2(n8701), .C1(n8426), 
        .C2(n8703), .ZN(n10305) );
  OR2_X1 U7917 ( .A1(n8428), .A2(n7661), .ZN(n7662) );
  NAND2_X1 U7918 ( .A1(n6359), .A2(n7662), .ZN(n6476) );
  XNOR2_X1 U7919 ( .A(n6476), .B(n7915), .ZN(n10308) );
  NOR2_X1 U7920 ( .A1(n8724), .A2(n5823), .ZN(n6361) );
  OAI22_X1 U7921 ( .A1(n8610), .A2(n10306), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n10181), .ZN(n6360) );
  AOI211_X1 U7922 ( .C1(n10308), .C2(n8670), .A(n6361), .B(n6360), .ZN(n6362)
         );
  OAI21_X1 U7923 ( .B1(n10305), .B2(n10198), .A(n6362), .ZN(P2_U3230) );
  INV_X1 U7924 ( .A(n6363), .ZN(n6370) );
  OAI22_X1 U7925 ( .A1(n6365), .A2(n8226), .B1(n10254), .B2(n5716), .ZN(n6364)
         );
  XNOR2_X1 U7926 ( .A(n6364), .B(n4495), .ZN(n6367) );
  OAI22_X1 U7927 ( .A1(n6365), .A2(n5702), .B1(n10254), .B2(n8226), .ZN(n6366)
         );
  OR2_X1 U7928 ( .A1(n6367), .A2(n6366), .ZN(n6553) );
  NAND2_X1 U7929 ( .A1(n6367), .A2(n6366), .ZN(n6368) );
  AND2_X1 U7930 ( .A1(n6553), .A2(n6368), .ZN(n6369) );
  INV_X1 U7931 ( .A(n6554), .ZN(n6373) );
  NOR3_X1 U7932 ( .A1(n6371), .A2(n6370), .A3(n6369), .ZN(n6372) );
  OAI21_X1 U7933 ( .B1(n6373), .B2(n6372), .A(n9342), .ZN(n6379) );
  INV_X1 U7934 ( .A(n6374), .ZN(n6377) );
  INV_X1 U7935 ( .A(n6434), .ZN(n6375) );
  OAI22_X1 U7936 ( .A1(n9314), .A2(n6375), .B1(n6549), .B2(n9345), .ZN(n6376)
         );
  AOI211_X1 U7937 ( .C1(n9334), .C2(n9638), .A(n6377), .B(n6376), .ZN(n6378)
         );
  OAI211_X1 U7938 ( .C1(n10254), .C2(n9350), .A(n6379), .B(n6378), .ZN(
        P1_U3239) );
  NAND2_X1 U7939 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n6381), .ZN(n6512) );
  OAI21_X1 U7940 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n6381), .A(n6512), .ZN(
        n6401) );
  NAND2_X1 U7941 ( .A1(n6391), .A2(n6390), .ZN(n6388) );
  MUX2_X1 U7942 ( .A(n6383), .B(n6382), .S(n8512), .Z(n6384) );
  INV_X1 U7943 ( .A(n6528), .ZN(n6730) );
  NAND2_X1 U7944 ( .A1(n6384), .A2(n6730), .ZN(n6522) );
  INV_X1 U7945 ( .A(n6384), .ZN(n6385) );
  NAND2_X1 U7946 ( .A1(n6385), .A2(n6528), .ZN(n6386) );
  NAND2_X1 U7947 ( .A1(n6522), .A2(n6386), .ZN(n6389) );
  INV_X1 U7948 ( .A(n6389), .ZN(n6387) );
  NAND2_X1 U7949 ( .A1(n6388), .A2(n6387), .ZN(n6523) );
  NAND3_X1 U7950 ( .A1(n6391), .A2(n6390), .A3(n6389), .ZN(n6392) );
  AOI21_X1 U7951 ( .B1(n6523), .B2(n6392), .A(n8517), .ZN(n6400) );
  NAND2_X1 U7952 ( .A1(P2_REG2_REG_11__SCAN_IN), .A2(n6394), .ZN(n6529) );
  OAI21_X1 U7953 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n6394), .A(n6529), .ZN(
        n6395) );
  NAND2_X1 U7954 ( .A1(n6395), .A2(n8526), .ZN(n6398) );
  INV_X1 U7955 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n6396) );
  NOR2_X1 U7956 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6396), .ZN(n7402) );
  AOI21_X1 U7957 ( .B1(n8519), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7402), .ZN(
        n6397) );
  OAI211_X1 U7958 ( .C1(n8522), .C2(n6528), .A(n6398), .B(n6397), .ZN(n6399)
         );
  AOI211_X1 U7959 ( .C1(n8442), .C2(n6401), .A(n6400), .B(n6399), .ZN(n6402)
         );
  INV_X1 U7960 ( .A(n6402), .ZN(P2_U3193) );
  INV_X1 U7961 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10388) );
  NOR2_X1 U7962 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n6403) );
  AOI21_X1 U7963 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n6403), .ZN(n10393) );
  NOR2_X1 U7964 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n6404) );
  AOI21_X1 U7965 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n6404), .ZN(n10396) );
  NOR2_X1 U7966 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(P2_ADDR_REG_15__SCAN_IN), 
        .ZN(n6405) );
  AOI21_X1 U7967 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n6405), .ZN(n10399) );
  NOR2_X1 U7968 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n6406) );
  AOI21_X1 U7969 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n6406), .ZN(n10402) );
  NOR2_X1 U7970 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n6407) );
  AOI21_X1 U7971 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n6407), .ZN(n10405) );
  NOR2_X1 U7972 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n6408) );
  AOI21_X1 U7973 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n6408), .ZN(n10408) );
  NOR2_X1 U7974 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n6409) );
  AOI21_X1 U7975 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n6409), .ZN(n10411) );
  NOR2_X1 U7976 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n6410) );
  AOI21_X1 U7977 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n6410), .ZN(n10414) );
  NOR2_X1 U7978 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n6411) );
  AOI21_X1 U7979 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n6411), .ZN(n10423) );
  NOR2_X1 U7980 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n6412) );
  AOI21_X1 U7981 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n6412), .ZN(n10429) );
  NOR2_X1 U7982 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n6413) );
  AOI21_X1 U7983 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n6413), .ZN(n10426) );
  NOR2_X1 U7984 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n6414) );
  AOI21_X1 U7985 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n6414), .ZN(n10417) );
  NOR2_X1 U7986 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n6415) );
  AOI21_X1 U7987 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n6415), .ZN(n10420) );
  AND2_X1 U7988 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n6416) );
  NOR2_X1 U7989 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n6416), .ZN(n10383) );
  INV_X1 U7990 ( .A(n10383), .ZN(n10384) );
  INV_X1 U7991 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10386) );
  NAND3_X1 U7992 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10385) );
  NAND2_X1 U7993 ( .A1(n10386), .A2(n10385), .ZN(n10382) );
  NAND2_X1 U7994 ( .A1(n10384), .A2(n10382), .ZN(n10432) );
  NAND2_X1 U7995 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n6417) );
  OAI21_X1 U7996 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n6417), .ZN(n10431) );
  NOR2_X1 U7997 ( .A1(n10432), .A2(n10431), .ZN(n10430) );
  AOI21_X1 U7998 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10430), .ZN(n10435) );
  NAND2_X1 U7999 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n6418) );
  OAI21_X1 U8000 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n6418), .ZN(n10434) );
  NOR2_X1 U8001 ( .A1(n10435), .A2(n10434), .ZN(n10433) );
  AOI21_X1 U8002 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10433), .ZN(n10438) );
  NOR2_X1 U8003 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n6419) );
  AOI21_X1 U8004 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n6419), .ZN(n10437) );
  NAND2_X1 U8005 ( .A1(n10438), .A2(n10437), .ZN(n10436) );
  OAI21_X1 U8006 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10436), .ZN(n10419) );
  NAND2_X1 U8007 ( .A1(n10420), .A2(n10419), .ZN(n10418) );
  OAI21_X1 U8008 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10418), .ZN(n10416) );
  NAND2_X1 U8009 ( .A1(n10417), .A2(n10416), .ZN(n10415) );
  OAI21_X1 U8010 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10415), .ZN(n10425) );
  NAND2_X1 U8011 ( .A1(n10426), .A2(n10425), .ZN(n10424) );
  OAI21_X1 U8012 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10424), .ZN(n10428) );
  NAND2_X1 U8013 ( .A1(n10429), .A2(n10428), .ZN(n10427) );
  OAI21_X1 U8014 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10427), .ZN(n10422) );
  NAND2_X1 U8015 ( .A1(n10423), .A2(n10422), .ZN(n10421) );
  OAI21_X1 U8016 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10421), .ZN(n10413) );
  NAND2_X1 U8017 ( .A1(n10414), .A2(n10413), .ZN(n10412) );
  OAI21_X1 U8018 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10412), .ZN(n10410) );
  NAND2_X1 U8019 ( .A1(n10411), .A2(n10410), .ZN(n10409) );
  OAI21_X1 U8020 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10409), .ZN(n10407) );
  NAND2_X1 U8021 ( .A1(n10408), .A2(n10407), .ZN(n10406) );
  OAI21_X1 U8022 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10406), .ZN(n10404) );
  NAND2_X1 U8023 ( .A1(n10405), .A2(n10404), .ZN(n10403) );
  OAI21_X1 U8024 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10403), .ZN(n10401) );
  NAND2_X1 U8025 ( .A1(n10402), .A2(n10401), .ZN(n10400) );
  OAI21_X1 U8026 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10400), .ZN(n10398) );
  NAND2_X1 U8027 ( .A1(n10399), .A2(n10398), .ZN(n10397) );
  OAI21_X1 U8028 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10397), .ZN(n10395) );
  NAND2_X1 U8029 ( .A1(n10396), .A2(n10395), .ZN(n10394) );
  OAI21_X1 U8030 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10394), .ZN(n10392) );
  NAND2_X1 U8031 ( .A1(n10393), .A2(n10392), .ZN(n10391) );
  OAI21_X1 U8032 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10391), .ZN(n10389) );
  NOR2_X1 U8033 ( .A1(n10388), .A2(n10389), .ZN(n6420) );
  NAND2_X1 U8034 ( .A1(n10388), .A2(n10389), .ZN(n10387) );
  OAI21_X1 U8035 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n6420), .A(n10387), .ZN(
        n6423) );
  XNOR2_X1 U8036 ( .A(n6421), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n6422) );
  XNOR2_X1 U8037 ( .A(n6423), .B(n6422), .ZN(ADD_1068_U4) );
  XNOR2_X1 U8038 ( .A(n6640), .B(n6424), .ZN(n6426) );
  OAI22_X1 U8039 ( .A1(n8270), .A2(n10011), .B1(n6549), .B2(n10013), .ZN(n6425) );
  AOI21_X1 U8040 ( .B1(n6426), .B2(n10009), .A(n6425), .ZN(n10258) );
  OR2_X1 U8041 ( .A1(n6428), .A2(n6427), .ZN(n6429) );
  NAND2_X1 U8042 ( .A1(n6430), .A2(n6429), .ZN(n10256) );
  OAI21_X1 U8043 ( .B1(n6431), .B2(n10254), .A(n10072), .ZN(n6433) );
  OR2_X1 U8044 ( .A1(n6433), .A2(n6432), .ZN(n10253) );
  INV_X1 U8045 ( .A(n10021), .ZN(n9774) );
  AOI22_X1 U8046 ( .A1(n9986), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n6434), .B2(
        n10022), .ZN(n6436) );
  INV_X1 U8047 ( .A(n10026), .ZN(n6824) );
  NAND2_X1 U8048 ( .A1(n6824), .A2(n6198), .ZN(n6435) );
  OAI211_X1 U8049 ( .C1(n10253), .C2(n9774), .A(n6436), .B(n6435), .ZN(n6437)
         );
  AOI21_X1 U8050 ( .B1(n10256), .B2(n9976), .A(n6437), .ZN(n6438) );
  OAI21_X1 U8051 ( .B1(n10258), .B2(n9986), .A(n6438), .ZN(P1_U3287) );
  INV_X1 U8052 ( .A(n6639), .ZN(n9389) );
  OAI21_X1 U8053 ( .B1(n6439), .B2(n9389), .A(n6642), .ZN(n6443) );
  NAND2_X1 U8054 ( .A1(n6587), .A2(n9467), .ZN(n6442) );
  AOI22_X1 U8055 ( .A1(n9473), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8043), .B2(
        n6440), .ZN(n6441) );
  NAND2_X1 U8056 ( .A1(n6442), .A2(n6441), .ZN(n6996) );
  NAND2_X1 U8057 ( .A1(n6996), .A2(n7041), .ZN(n9398) );
  NAND2_X1 U8058 ( .A1(n9396), .A2(n9398), .ZN(n6450) );
  XNOR2_X1 U8059 ( .A(n6443), .B(n6450), .ZN(n6444) );
  NAND2_X1 U8060 ( .A1(n6444), .A2(n10009), .ZN(n6446) );
  OR2_X1 U8061 ( .A1(n7113), .A2(n10011), .ZN(n6445) );
  NAND2_X1 U8062 ( .A1(n6446), .A2(n6445), .ZN(n10261) );
  INV_X1 U8063 ( .A(n10261), .ZN(n6463) );
  INV_X1 U8064 ( .A(n7113), .ZN(n9635) );
  NAND2_X1 U8065 ( .A1(n6448), .A2(n6447), .ZN(n6449) );
  OAI21_X1 U8066 ( .B1(n6449), .B2(n6450), .A(n6678), .ZN(n10263) );
  XNOR2_X1 U8067 ( .A(n6682), .B(n4837), .ZN(n6458) );
  NAND2_X1 U8068 ( .A1(n9476), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6457) );
  NOR2_X1 U8069 ( .A1(n6451), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6452) );
  OR2_X1 U8070 ( .A1(n6651), .A2(n6452), .ZN(n7328) );
  INV_X1 U8071 ( .A(n7328), .ZN(n6453) );
  NAND2_X1 U8072 ( .A1(n5720), .A2(n6453), .ZN(n6456) );
  NAND2_X1 U8073 ( .A1(n9477), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6455) );
  NAND2_X1 U8074 ( .A1(n4492), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6454) );
  INV_X1 U8075 ( .A(n7013), .ZN(n9634) );
  AOI22_X1 U8076 ( .A1(n6458), .A2(n10072), .B1(n9999), .B2(n9634), .ZN(n10260) );
  AOI22_X1 U8077 ( .A1(n9986), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7112), .B2(
        n10022), .ZN(n6460) );
  NAND2_X1 U8078 ( .A1(n6824), .A2(n6996), .ZN(n6459) );
  OAI211_X1 U8079 ( .C1(n10260), .C2(n9774), .A(n6460), .B(n6459), .ZN(n6461)
         );
  AOI21_X1 U8080 ( .B1(n10263), .B2(n9976), .A(n6461), .ZN(n6462) );
  OAI21_X1 U8081 ( .B1(n6463), .B2(n9986), .A(n6462), .ZN(P1_U3284) );
  OAI21_X1 U8082 ( .B1(n9494), .B2(n6465), .A(n6464), .ZN(n6466) );
  AOI222_X1 U8083 ( .A1(n10009), .A2(n6466), .B1(n9638), .B2(n9999), .C1(n5739), .C2(n9997), .ZN(n10248) );
  OAI21_X1 U8084 ( .B1(n6469), .B2(n6468), .A(n6467), .ZN(n10251) );
  OAI211_X1 U8085 ( .C1(n6471), .C2(n10247), .A(n10072), .B(n6470), .ZN(n10246) );
  AOI22_X1 U8086 ( .A1(n9986), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n8272), .B2(
        n10022), .ZN(n6473) );
  NAND2_X1 U8087 ( .A1(n6824), .A2(n5899), .ZN(n6472) );
  OAI211_X1 U8088 ( .C1(n10246), .C2(n9774), .A(n6473), .B(n6472), .ZN(n6474)
         );
  AOI21_X1 U8089 ( .B1(n10251), .B2(n9976), .A(n6474), .ZN(n6475) );
  OAI21_X1 U8090 ( .B1(n10248), .B2(n9986), .A(n6475), .ZN(P1_U3289) );
  NAND2_X1 U8091 ( .A1(n6476), .A2(n7915), .ZN(n6477) );
  NAND2_X1 U8092 ( .A1(n6477), .A2(n7674), .ZN(n6491) );
  OR2_X1 U8093 ( .A1(n8426), .A2(n10309), .ZN(n7671) );
  NAND2_X1 U8094 ( .A1(n8426), .A2(n10309), .ZN(n7677) );
  NAND2_X1 U8095 ( .A1(n7671), .A2(n7677), .ZN(n7917) );
  XOR2_X1 U8096 ( .A(n6491), .B(n7917), .Z(n10312) );
  OAI22_X1 U8097 ( .A1(n8610), .A2(n10309), .B1(n6478), .B2(n10181), .ZN(n6489) );
  NOR2_X1 U8098 ( .A1(n8427), .A2(n6481), .ZN(n6479) );
  NAND2_X1 U8099 ( .A1(n8427), .A2(n6481), .ZN(n6482) );
  INV_X1 U8100 ( .A(n7917), .ZN(n6484) );
  XNOR2_X1 U8101 ( .A(n6497), .B(n6484), .ZN(n6485) );
  NAND2_X1 U8102 ( .A1(n6485), .A2(n8706), .ZN(n6487) );
  AOI22_X1 U8103 ( .A1(n8703), .A2(n8425), .B1(n8427), .B2(n8701), .ZN(n6486)
         );
  NAND2_X1 U8104 ( .A1(n6487), .A2(n6486), .ZN(n10310) );
  MUX2_X1 U8105 ( .A(n10310), .B(P2_REG2_REG_4__SCAN_IN), .S(n10198), .Z(n6488) );
  AOI211_X1 U8106 ( .C1(n8670), .C2(n10312), .A(n6489), .B(n6488), .ZN(n6490)
         );
  INV_X1 U8107 ( .A(n6490), .ZN(P2_U3229) );
  INV_X1 U8108 ( .A(n8570), .ZN(n6504) );
  NAND2_X1 U8109 ( .A1(n6491), .A2(n7677), .ZN(n6492) );
  NAND2_X1 U8110 ( .A1(n6492), .A2(n7671), .ZN(n6494) );
  NAND2_X1 U8111 ( .A1(n8425), .A2(n10314), .ZN(n7676) );
  NAND2_X1 U8112 ( .A1(n6494), .A2(n7676), .ZN(n6563) );
  OR2_X1 U8113 ( .A1(n8425), .A2(n10314), .ZN(n7679) );
  INV_X1 U8114 ( .A(n7679), .ZN(n6495) );
  OR2_X1 U8115 ( .A1(n8425), .A2(n6508), .ZN(n6599) );
  NAND2_X1 U8116 ( .A1(n8425), .A2(n6508), .ZN(n6689) );
  AND2_X1 U8117 ( .A1(n6599), .A2(n6689), .ZN(n7918) );
  INV_X1 U8118 ( .A(n7918), .ZN(n6493) );
  OAI22_X1 U8119 ( .A1(n6563), .A2(n6495), .B1(n6494), .B2(n6493), .ZN(n10317)
         );
  OR2_X1 U8120 ( .A1(n8426), .A2(n6498), .ZN(n6496) );
  NAND2_X1 U8121 ( .A1(n6497), .A2(n6496), .ZN(n6500) );
  NAND2_X1 U8122 ( .A1(n8426), .A2(n6498), .ZN(n6499) );
  NAND2_X1 U8123 ( .A1(n6500), .A2(n6499), .ZN(n6600) );
  XNOR2_X1 U8124 ( .A(n6600), .B(n7918), .ZN(n6503) );
  INV_X1 U8125 ( .A(n10336), .ZN(n10349) );
  NAND2_X1 U8126 ( .A1(n10317), .A2(n10349), .ZN(n6502) );
  AOI22_X1 U8127 ( .A1(n8701), .A2(n8426), .B1(n8424), .B2(n8703), .ZN(n6501)
         );
  OAI211_X1 U8128 ( .C1(n10296), .C2(n6503), .A(n6502), .B(n6501), .ZN(n10315)
         );
  AOI21_X1 U8129 ( .B1(n6504), .B2(n10317), .A(n10315), .ZN(n6510) );
  INV_X1 U8130 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6506) );
  OAI22_X1 U8131 ( .A1(n8724), .A2(n6506), .B1(n6505), .B2(n10181), .ZN(n6507)
         );
  AOI21_X1 U8132 ( .B1(n8726), .B2(n6508), .A(n6507), .ZN(n6509) );
  OAI21_X1 U8133 ( .B1(n6510), .B2(n10198), .A(n6509), .ZN(P2_U3228) );
  INV_X1 U8134 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10379) );
  AOI22_X1 U8135 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n6534), .B1(n7061), .B2(
        n10379), .ZN(n6515) );
  NAND2_X1 U8136 ( .A1(n6528), .A2(n6511), .ZN(n6513) );
  NAND2_X1 U8137 ( .A1(n6513), .A2(n6512), .ZN(n6514) );
  NAND2_X1 U8138 ( .A1(n6515), .A2(n6514), .ZN(n6862) );
  OAI21_X1 U8139 ( .B1(n6515), .B2(n6514), .A(n6862), .ZN(n6526) );
  NAND2_X1 U8140 ( .A1(n6523), .A2(n6522), .ZN(n6520) );
  INV_X1 U8141 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6736) );
  MUX2_X1 U8142 ( .A(n6736), .B(n10379), .S(n8512), .Z(n6516) );
  NAND2_X1 U8143 ( .A1(n6516), .A2(n7061), .ZN(n6873) );
  INV_X1 U8144 ( .A(n6516), .ZN(n6517) );
  NAND2_X1 U8145 ( .A1(n6517), .A2(n6534), .ZN(n6518) );
  NAND2_X1 U8146 ( .A1(n6873), .A2(n6518), .ZN(n6521) );
  INV_X1 U8147 ( .A(n6521), .ZN(n6519) );
  NAND2_X1 U8148 ( .A1(n6520), .A2(n6519), .ZN(n6874) );
  NAND3_X1 U8149 ( .A1(n6523), .A2(n6522), .A3(n6521), .ZN(n6524) );
  AOI21_X1 U8150 ( .B1(n6874), .B2(n6524), .A(n8517), .ZN(n6525) );
  AOI21_X1 U8151 ( .B1(n6526), .B2(n8442), .A(n6525), .ZN(n6538) );
  AOI22_X1 U8152 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n6534), .B1(n7061), .B2(
        n6736), .ZN(n6532) );
  NAND2_X1 U8153 ( .A1(n6528), .A2(n6527), .ZN(n6530) );
  OAI21_X1 U8154 ( .B1(n6532), .B2(n6531), .A(n6865), .ZN(n6536) );
  NAND2_X1 U8155 ( .A1(n8519), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n6533) );
  NAND2_X1 U8156 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7455) );
  OAI211_X1 U8157 ( .C1(n8522), .C2(n6534), .A(n6533), .B(n7455), .ZN(n6535)
         );
  AOI21_X1 U8158 ( .B1(n6536), .B2(n8526), .A(n6535), .ZN(n6537) );
  NAND2_X1 U8159 ( .A1(n6538), .A2(n6537), .ZN(P2_U3194) );
  MUX2_X1 U8160 ( .A(n7748), .B(n6811), .S(n7901), .Z(n6544) );
  NAND2_X1 U8161 ( .A1(n6544), .A2(n6543), .ZN(n6717) );
  INV_X1 U8162 ( .A(n6544), .ZN(n6545) );
  NAND2_X1 U8163 ( .A1(n6545), .A2(SI_20_), .ZN(n6546) );
  XNOR2_X1 U8164 ( .A(n6716), .B(n6715), .ZN(n8057) );
  INV_X1 U8165 ( .A(n8057), .ZN(n6812) );
  OAI222_X1 U8166 ( .A1(n9220), .A2(n6812), .B1(n6547), .B2(P2_U3151), .C1(
        n7748), .C2(n9222), .ZN(P2_U3275) );
  AOI22_X1 U8167 ( .A1(n9636), .A2(n5521), .B1(n6550), .B2(n8208), .ZN(n6548)
         );
  XNOR2_X1 U8168 ( .A(n6548), .B(n4495), .ZN(n6988) );
  OR2_X1 U8169 ( .A1(n6549), .A2(n5702), .ZN(n6552) );
  NAND2_X1 U8170 ( .A1(n6550), .A2(n5521), .ZN(n6551) );
  NAND2_X1 U8171 ( .A1(n6552), .A2(n6551), .ZN(n6989) );
  XNOR2_X1 U8172 ( .A(n6988), .B(n6989), .ZN(n6556) );
  OAI21_X1 U8173 ( .B1(n6556), .B2(n6555), .A(n6992), .ZN(n6557) );
  NAND2_X1 U8174 ( .A1(n6557), .A2(n9342), .ZN(n6562) );
  INV_X1 U8175 ( .A(n6630), .ZN(n6558) );
  OAI22_X1 U8176 ( .A1(n9314), .A2(n6558), .B1(n7113), .B2(n9345), .ZN(n6559)
         );
  AOI211_X1 U8177 ( .C1(n9334), .C2(n9637), .A(n6560), .B(n6559), .ZN(n6561)
         );
  OAI211_X1 U8178 ( .C1(n6633), .C2(n9350), .A(n6562), .B(n6561), .ZN(P1_U3213) );
  NAND2_X1 U8179 ( .A1(n6563), .A2(n7679), .ZN(n6688) );
  INV_X1 U8180 ( .A(n6688), .ZN(n6568) );
  NAND2_X1 U8181 ( .A1(n6194), .A2(n7873), .ZN(n6567) );
  INV_X2 U8182 ( .A(n7874), .ZN(n7737) );
  AOI22_X1 U8183 ( .A1(n7737), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7736), .B2(
        n6565), .ZN(n6566) );
  OR2_X1 U8184 ( .A1(n8424), .A2(n6771), .ZN(n7680) );
  INV_X1 U8185 ( .A(n7680), .ZN(n7673) );
  NAND2_X1 U8186 ( .A1(n8424), .A2(n6771), .ZN(n7681) );
  NAND2_X1 U8187 ( .A1(n6569), .A2(n7873), .ZN(n6572) );
  AOI22_X1 U8188 ( .A1(n7737), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7736), .B2(
        n6570), .ZN(n6571) );
  NAND2_X1 U8189 ( .A1(n10333), .A2(n7439), .ZN(n7690) );
  INV_X1 U8190 ( .A(n7690), .ZN(n6586) );
  OR2_X1 U8191 ( .A1(n10333), .A2(n7439), .ZN(n7683) );
  NAND2_X1 U8192 ( .A1(n7903), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6585) );
  INV_X1 U8193 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6576) );
  AND2_X1 U8194 ( .A1(n6577), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6578) );
  NOR2_X1 U8195 ( .A1(n6579), .A2(n6578), .ZN(n6777) );
  OR2_X1 U8196 ( .A1(n7288), .A2(n6777), .ZN(n6583) );
  OR2_X1 U8197 ( .A1(n6581), .A2(n6580), .ZN(n6582) );
  AND2_X1 U8198 ( .A1(n7683), .A2(n6900), .ZN(n7694) );
  OR2_X1 U8199 ( .A1(n6586), .A2(n7694), .ZN(n6591) );
  AND2_X1 U8200 ( .A1(n7681), .A2(n6591), .ZN(n6745) );
  NAND2_X1 U8201 ( .A1(n6747), .A2(n6745), .ZN(n6596) );
  NAND2_X1 U8202 ( .A1(n6587), .A2(n7873), .ZN(n6590) );
  AOI22_X1 U8203 ( .A1(n7737), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7736), .B2(
        n6588), .ZN(n6589) );
  NAND2_X1 U8204 ( .A1(n6590), .A2(n6589), .ZN(n10334) );
  OR2_X1 U8205 ( .A1(n10334), .A2(n7443), .ZN(n7684) );
  NAND2_X1 U8206 ( .A1(n10334), .A2(n7443), .ZN(n7691) );
  NAND2_X1 U8207 ( .A1(n7684), .A2(n7691), .ZN(n7924) );
  INV_X1 U8208 ( .A(n7924), .ZN(n6594) );
  INV_X1 U8209 ( .A(n6591), .ZN(n6593) );
  NAND2_X1 U8210 ( .A1(n6934), .A2(n6969), .ZN(n7689) );
  AND2_X1 U8211 ( .A1(n7922), .A2(n7690), .ZN(n6592) );
  OR2_X1 U8212 ( .A1(n6593), .A2(n6592), .ZN(n6595) );
  AND2_X1 U8213 ( .A1(n6594), .A2(n6595), .ZN(n6748) );
  NAND2_X1 U8214 ( .A1(n6596), .A2(n6748), .ZN(n6829) );
  NAND2_X1 U8215 ( .A1(n6596), .A2(n6595), .ZN(n6597) );
  NAND2_X1 U8216 ( .A1(n6597), .A2(n7924), .ZN(n6598) );
  NAND2_X1 U8217 ( .A1(n6829), .A2(n6598), .ZN(n10337) );
  NAND2_X1 U8218 ( .A1(n6600), .A2(n6599), .ZN(n6690) );
  INV_X1 U8219 ( .A(n6771), .ZN(n10322) );
  AND2_X1 U8220 ( .A1(n10322), .A2(n8424), .ZN(n6902) );
  INV_X1 U8221 ( .A(n6902), .ZN(n6601) );
  AND2_X1 U8222 ( .A1(n6601), .A2(n6689), .ZN(n6602) );
  INV_X1 U8223 ( .A(n7439), .ZN(n7441) );
  OR2_X1 U8224 ( .A1(n10333), .A2(n7441), .ZN(n6606) );
  INV_X1 U8225 ( .A(n6934), .ZN(n10324) );
  NAND2_X1 U8226 ( .A1(n10324), .A2(n6969), .ZN(n6605) );
  NAND2_X1 U8227 ( .A1(n6690), .A2(n6603), .ZN(n6610) );
  INV_X1 U8228 ( .A(n6604), .ZN(n6608) );
  NAND2_X1 U8229 ( .A1(n6778), .A2(n6771), .ZN(n6921) );
  AND2_X1 U8230 ( .A1(n6921), .A2(n6605), .ZN(n6904) );
  AND2_X1 U8231 ( .A1(n6904), .A2(n6606), .ZN(n6607) );
  NAND2_X1 U8232 ( .A1(n6610), .A2(n6609), .ZN(n6719) );
  XNOR2_X1 U8233 ( .A(n6719), .B(n7924), .ZN(n6611) );
  NAND2_X1 U8234 ( .A1(n6611), .A2(n8706), .ZN(n6623) );
  NAND2_X1 U8235 ( .A1(n4814), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6620) );
  OR2_X1 U8236 ( .A1(n7865), .A2(n6612), .ZN(n6619) );
  OR2_X1 U8237 ( .A1(n6581), .A2(n6613), .ZN(n6618) );
  NAND2_X1 U8238 ( .A1(n6614), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6615) );
  AND2_X1 U8239 ( .A1(n6616), .A2(n6615), .ZN(n7133) );
  OR2_X1 U8240 ( .A1(n7288), .A2(n7133), .ZN(n6617) );
  OAI22_X1 U8241 ( .A1(n7439), .A2(n10192), .B1(n7404), .B2(n10194), .ZN(n6621) );
  INV_X1 U8242 ( .A(n6621), .ZN(n6622) );
  NAND2_X1 U8243 ( .A1(n6623), .A2(n6622), .ZN(n10340) );
  NAND2_X1 U8244 ( .A1(n10340), .A2(n8724), .ZN(n6627) );
  OAI22_X1 U8245 ( .A1(n8724), .A2(n6624), .B1(n7435), .B2(n10181), .ZN(n6625)
         );
  AOI21_X1 U8246 ( .B1(n8726), .B2(n10334), .A(n6625), .ZN(n6626) );
  OAI211_X1 U8247 ( .C1(n8729), .C2(n10337), .A(n6627), .B(n6626), .ZN(
        P2_U3224) );
  INV_X1 U8248 ( .A(n6628), .ZN(n6637) );
  NAND2_X1 U8249 ( .A1(n6629), .A2(n10021), .ZN(n6632) );
  AOI22_X1 U8250 ( .A1(n9986), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n6630), .B2(
        n10022), .ZN(n6631) );
  OAI211_X1 U8251 ( .C1(n6633), .C2(n10026), .A(n6632), .B(n6631), .ZN(n6634)
         );
  AOI21_X1 U8252 ( .B1(n6635), .B2(n9976), .A(n6634), .ZN(n6636) );
  OAI21_X1 U8253 ( .B1(n6637), .B2(n9986), .A(n6636), .ZN(P1_U3286) );
  NAND2_X1 U8254 ( .A1(n6643), .A2(n9382), .ZN(n9544) );
  OR2_X1 U8255 ( .A1(n6640), .A2(n9544), .ZN(n6817) );
  AND2_X1 U8256 ( .A1(n6642), .A2(n6641), .ZN(n9383) );
  NAND3_X1 U8257 ( .A1(n9396), .A2(n9383), .A3(n9381), .ZN(n9497) );
  NAND2_X1 U8258 ( .A1(n6643), .A2(n9497), .ZN(n9547) );
  NAND2_X1 U8259 ( .A1(n6722), .A2(n9467), .ZN(n6646) );
  AOI22_X1 U8260 ( .A1(n9473), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n8043), .B2(
        n6644), .ZN(n6645) );
  NAND2_X1 U8261 ( .A1(n6646), .A2(n6645), .ZN(n7012) );
  OR2_X1 U8262 ( .A1(n7012), .A2(n7013), .ZN(n9548) );
  NAND2_X1 U8263 ( .A1(n7012), .A2(n7013), .ZN(n9399) );
  NAND2_X1 U8264 ( .A1(n9548), .A2(n9399), .ZN(n9498) );
  INV_X1 U8265 ( .A(n9498), .ZN(n6816) );
  AND2_X1 U8266 ( .A1(n9547), .A2(n6816), .ZN(n6647) );
  NAND2_X1 U8267 ( .A1(n6817), .A2(n6647), .ZN(n6815) );
  NAND2_X1 U8268 ( .A1(n6729), .A2(n9467), .ZN(n6650) );
  AOI22_X1 U8269 ( .A1(n9473), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n4494), .B2(
        n6648), .ZN(n6649) );
  NAND2_X1 U8270 ( .A1(n6651), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6661) );
  OR2_X1 U8271 ( .A1(n6651), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6652) );
  AND2_X1 U8272 ( .A1(n6661), .A2(n6652), .ZN(n7027) );
  NAND2_X1 U8273 ( .A1(n5720), .A2(n7027), .ZN(n6656) );
  NAND2_X1 U8274 ( .A1(n9476), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6655) );
  NAND2_X1 U8275 ( .A1(n9477), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6654) );
  NAND2_X1 U8276 ( .A1(n4491), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6653) );
  NAND2_X1 U8277 ( .A1(n7031), .A2(n7327), .ZN(n9403) );
  AND2_X1 U8278 ( .A1(n9403), .A2(n9399), .ZN(n9550) );
  NAND2_X1 U8279 ( .A1(n6815), .A2(n9550), .ZN(n6841) );
  OR2_X1 U8280 ( .A1(n7031), .A2(n7327), .ZN(n9401) );
  NAND2_X1 U8281 ( .A1(n6841), .A2(n9401), .ZN(n6667) );
  NAND2_X1 U8282 ( .A1(n7060), .A2(n9467), .ZN(n6659) );
  AOI22_X1 U8283 ( .A1(n9473), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n8043), .B2(
        n6657), .ZN(n6658) );
  NAND2_X1 U8284 ( .A1(n6659), .A2(n6658), .ZN(n7238) );
  NAND2_X1 U8285 ( .A1(n6661), .A2(n6660), .ZN(n6662) );
  AND2_X1 U8286 ( .A1(n6669), .A2(n6662), .ZN(n7234) );
  NAND2_X1 U8287 ( .A1(n5720), .A2(n7234), .ZN(n6666) );
  NAND2_X1 U8288 ( .A1(n9476), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6665) );
  NAND2_X1 U8289 ( .A1(n4492), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6664) );
  NAND2_X1 U8290 ( .A1(n9477), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6663) );
  OR2_X1 U8291 ( .A1(n7238), .A2(n7420), .ZN(n9404) );
  NAND2_X1 U8292 ( .A1(n7238), .A2(n7420), .ZN(n9554) );
  NAND2_X1 U8293 ( .A1(n9404), .A2(n9554), .ZN(n9501) );
  XNOR2_X1 U8294 ( .A(n6667), .B(n9501), .ZN(n6676) );
  NAND2_X1 U8295 ( .A1(n9476), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6674) );
  NAND2_X1 U8296 ( .A1(n6669), .A2(n6668), .ZN(n6670) );
  AND2_X1 U8297 ( .A1(n6847), .A2(n6670), .ZN(n7418) );
  NAND2_X1 U8298 ( .A1(n5720), .A2(n7418), .ZN(n6673) );
  NAND2_X1 U8299 ( .A1(n9477), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6672) );
  NAND2_X1 U8300 ( .A1(n4491), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6671) );
  OAI22_X1 U8301 ( .A1(n7414), .A2(n10013), .B1(n7327), .B2(n10011), .ZN(n6675) );
  AOI21_X1 U8302 ( .B1(n6676), .B2(n10009), .A(n6675), .ZN(n10273) );
  NAND2_X1 U8303 ( .A1(n6678), .A2(n6677), .ZN(n6814) );
  NAND2_X1 U8304 ( .A1(n6814), .A2(n9498), .ZN(n6813) );
  NAND2_X1 U8305 ( .A1(n6813), .A2(n6679), .ZN(n6756) );
  NAND2_X1 U8306 ( .A1(n9401), .A2(n9403), .ZN(n9500) );
  INV_X1 U8307 ( .A(n7327), .ZN(n9633) );
  NAND2_X1 U8308 ( .A1(n6755), .A2(n6680), .ZN(n6681) );
  NAND2_X2 U8309 ( .A1(n6681), .A2(n9501), .ZN(n6837) );
  OAI21_X1 U8310 ( .B1(n6681), .B2(n9501), .A(n6837), .ZN(n10277) );
  NAND2_X1 U8311 ( .A1(n10277), .A2(n9976), .ZN(n6687) );
  NOR2_X2 U8312 ( .A1(n6682), .A2(n6996), .ZN(n6822) );
  INV_X1 U8313 ( .A(n7012), .ZN(n10265) );
  NAND2_X1 U8314 ( .A1(n6822), .A2(n10265), .ZN(n6821) );
  OAI211_X1 U8315 ( .C1(n4862), .C2(n4861), .A(n10072), .B(n6855), .ZN(n10272)
         );
  INV_X1 U8316 ( .A(n10272), .ZN(n6685) );
  AOI22_X1 U8317 ( .A1(n9986), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7234), .B2(
        n10022), .ZN(n6683) );
  OAI21_X1 U8318 ( .B1(n4861), .B2(n10026), .A(n6683), .ZN(n6684) );
  AOI21_X1 U8319 ( .B1(n6685), .B2(n10021), .A(n6684), .ZN(n6686) );
  OAI211_X1 U8320 ( .C1(n9986), .C2(n10273), .A(n6687), .B(n6686), .ZN(
        P1_U3281) );
  AND2_X1 U8321 ( .A1(n7680), .A2(n7681), .ZN(n7920) );
  XOR2_X1 U8322 ( .A(n7920), .B(n6688), .Z(n10319) );
  NAND2_X1 U8323 ( .A1(n6690), .A2(n6689), .ZN(n6903) );
  XOR2_X1 U8324 ( .A(n7920), .B(n6903), .Z(n6691) );
  OAI222_X1 U8325 ( .A1(n10194), .A2(n6969), .B1(n10192), .B2(n6789), .C1(
        n6691), .C2(n10296), .ZN(n10320) );
  NAND2_X1 U8326 ( .A1(n10320), .A2(n8724), .ZN(n6694) );
  OAI22_X1 U8327 ( .A1(n8724), .A2(n6239), .B1(n6785), .B2(n10181), .ZN(n6692)
         );
  AOI21_X1 U8328 ( .B1(n8726), .B2(n10322), .A(n6692), .ZN(n6693) );
  OAI211_X1 U8329 ( .C1(n8729), .C2(n10319), .A(n6694), .B(n6693), .ZN(
        P2_U3227) );
  INV_X1 U8330 ( .A(n6695), .ZN(n6704) );
  NAND2_X1 U8331 ( .A1(n6696), .A2(n10021), .ZN(n6699) );
  AOI22_X1 U8332 ( .A1(n9986), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n6697), .B2(
        n10022), .ZN(n6698) );
  OAI211_X1 U8333 ( .C1(n6700), .C2(n10026), .A(n6699), .B(n6698), .ZN(n6701)
         );
  AOI21_X1 U8334 ( .B1(n9976), .B2(n6702), .A(n6701), .ZN(n6703) );
  OAI21_X1 U8335 ( .B1(n6704), .B2(n9986), .A(n6703), .ZN(P1_U3288) );
  NAND2_X1 U8336 ( .A1(n10021), .A2(n10072), .ZN(n9769) );
  INV_X1 U8337 ( .A(n9769), .ZN(n9918) );
  OAI21_X1 U8338 ( .B1(n9918), .B2(n6824), .A(n6705), .ZN(n6713) );
  INV_X1 U8339 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6710) );
  NAND3_X1 U8340 ( .A1(n9489), .A2(n6707), .A3(n6706), .ZN(n6709) );
  OAI211_X1 U8341 ( .C1(n9980), .C2(n6710), .A(n6709), .B(n6708), .ZN(n6711)
         );
  NAND2_X1 U8342 ( .A1(n6711), .A2(n10028), .ZN(n6712) );
  OAI211_X1 U8343 ( .C1(n6714), .C2(n10028), .A(n6713), .B(n6712), .ZN(
        P1_U3293) );
  MUX2_X1 U8344 ( .A(n7637), .B(n6797), .S(n7901), .Z(n6892) );
  XNOR2_X1 U8345 ( .A(n6892), .B(SI_21_), .ZN(n6891) );
  XNOR2_X1 U8346 ( .A(n6890), .B(n6891), .ZN(n8072) );
  INV_X1 U8347 ( .A(n8072), .ZN(n6798) );
  OAI222_X1 U8348 ( .A1(n9220), .A2(n6798), .B1(n4760), .B2(P2_U3151), .C1(
        n7637), .C2(n9222), .ZN(P2_U3274) );
  INV_X1 U8349 ( .A(n7443), .ZN(n7123) );
  NAND2_X1 U8350 ( .A1(n10334), .A2(n7123), .ZN(n6718) );
  NAND2_X1 U8351 ( .A1(n6719), .A2(n6718), .ZN(n6721) );
  OR2_X1 U8352 ( .A1(n10334), .A2(n7123), .ZN(n6720) );
  NAND2_X1 U8353 ( .A1(n6721), .A2(n6720), .ZN(n6831) );
  NAND2_X1 U8354 ( .A1(n6722), .A2(n7873), .ZN(n6725) );
  AOI22_X1 U8355 ( .A1(n7737), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7736), .B2(
        n6723), .ZN(n6724) );
  NAND2_X1 U8356 ( .A1(n6725), .A2(n6724), .ZN(n10342) );
  INV_X1 U8357 ( .A(n7404), .ZN(n8422) );
  NAND2_X1 U8358 ( .A1(n10342), .A2(n8422), .ZN(n6726) );
  NAND2_X1 U8359 ( .A1(n6831), .A2(n6726), .ZN(n6728) );
  OR2_X1 U8360 ( .A1(n10342), .A2(n8422), .ZN(n6727) );
  NAND2_X1 U8361 ( .A1(n6728), .A2(n6727), .ZN(n6733) );
  NAND2_X1 U8362 ( .A1(n6729), .A2(n7873), .ZN(n6732) );
  AOI22_X1 U8363 ( .A1(n7737), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n7736), .B2(
        n6730), .ZN(n6731) );
  NAND2_X1 U8364 ( .A1(n6732), .A2(n6731), .ZN(n7059) );
  OR2_X1 U8365 ( .A1(n7059), .A2(n7066), .ZN(n7707) );
  NAND2_X1 U8366 ( .A1(n7059), .A2(n7066), .ZN(n7708) );
  AOI21_X1 U8367 ( .B1(n6733), .B2(n7928), .A(n10296), .ZN(n6744) );
  NAND2_X1 U8368 ( .A1(n4814), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6742) );
  OR2_X1 U8369 ( .A1(n7865), .A2(n6736), .ZN(n6741) );
  NOR2_X2 U8370 ( .A1(n6737), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7052) );
  AND2_X1 U8371 ( .A1(n6737), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6738) );
  NOR2_X1 U8372 ( .A1(n7052), .A2(n6738), .ZN(n7460) );
  OR2_X1 U8373 ( .A1(n7288), .A2(n7460), .ZN(n6740) );
  OR2_X1 U8374 ( .A1(n6581), .A2(n10379), .ZN(n6739) );
  OAI22_X1 U8375 ( .A1(n7404), .A2(n10192), .B1(n10191), .B2(n10194), .ZN(
        n6743) );
  AOI21_X1 U8376 ( .B1(n6744), .B2(n7349), .A(n6743), .ZN(n10351) );
  OR2_X1 U8377 ( .A1(n10342), .A2(n7404), .ZN(n7706) );
  AND2_X1 U8378 ( .A1(n7706), .A2(n7684), .ZN(n7693) );
  AND2_X1 U8379 ( .A1(n6745), .A2(n7693), .ZN(n6746) );
  INV_X1 U8380 ( .A(n7693), .ZN(n6749) );
  OR2_X1 U8381 ( .A1(n6749), .A2(n6748), .ZN(n6750) );
  NAND2_X1 U8382 ( .A1(n10342), .A2(n7404), .ZN(n7701) );
  XNOR2_X1 U8383 ( .A(n7068), .B(n7928), .ZN(n10355) );
  INV_X1 U8384 ( .A(n7059), .ZN(n10353) );
  INV_X1 U8385 ( .A(n6751), .ZN(n7406) );
  AOI22_X1 U8386 ( .A1(n10198), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n8709), .B2(
        n7406), .ZN(n6752) );
  OAI21_X1 U8387 ( .B1(n10353), .B2(n8610), .A(n6752), .ZN(n6753) );
  AOI21_X1 U8388 ( .B1(n10355), .B2(n8670), .A(n6753), .ZN(n6754) );
  OAI21_X1 U8389 ( .B1(n10351), .B2(n10198), .A(n6754), .ZN(P2_U3222) );
  OAI21_X1 U8390 ( .B1(n6756), .B2(n9500), .A(n6755), .ZN(n6915) );
  INV_X1 U8391 ( .A(n6915), .ZN(n6765) );
  NAND2_X1 U8392 ( .A1(n6815), .A2(n9399), .ZN(n6757) );
  XNOR2_X1 U8393 ( .A(n6757), .B(n9500), .ZN(n6760) );
  NAND2_X1 U8394 ( .A1(n6915), .A2(n7337), .ZN(n6759) );
  AOI22_X1 U8395 ( .A1(n9997), .A2(n9634), .B1(n9632), .B2(n9999), .ZN(n6758)
         );
  OAI211_X1 U8396 ( .C1(n9938), .C2(n6760), .A(n6759), .B(n6758), .ZN(n6913)
         );
  NAND2_X1 U8397 ( .A1(n6913), .A2(n10028), .ZN(n6764) );
  AOI211_X1 U8398 ( .C1(n7031), .C2(n6821), .A(n10266), .B(n4862), .ZN(n6914)
         );
  INV_X1 U8399 ( .A(n7031), .ZN(n6920) );
  AOI22_X1 U8400 ( .A1(n9986), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7027), .B2(
        n10022), .ZN(n6761) );
  OAI21_X1 U8401 ( .B1(n6920), .B2(n10026), .A(n6761), .ZN(n6762) );
  AOI21_X1 U8402 ( .B1(n6914), .B2(n10021), .A(n6762), .ZN(n6763) );
  OAI211_X1 U8403 ( .C1(n6765), .C2(n7343), .A(n6764), .B(n6763), .ZN(P1_U3282) );
  NAND2_X1 U8404 ( .A1(n6767), .A2(n6766), .ZN(n6770) );
  OR2_X1 U8405 ( .A1(n6768), .A2(n8425), .ZN(n6769) );
  NAND2_X1 U8406 ( .A1(n6770), .A2(n6769), .ZN(n6792) );
  XNOR2_X1 U8407 ( .A(n6771), .B(n8258), .ZN(n6772) );
  XNOR2_X1 U8408 ( .A(n6772), .B(n8424), .ZN(n6793) );
  OR2_X2 U8409 ( .A1(n6792), .A2(n6793), .ZN(n6790) );
  NAND2_X1 U8410 ( .A1(n6772), .A2(n8424), .ZN(n6773) );
  XNOR2_X1 U8411 ( .A(n6934), .B(n8139), .ZN(n6965) );
  XNOR2_X1 U8412 ( .A(n6965), .B(n6969), .ZN(n6774) );
  OAI21_X1 U8413 ( .B1(n6775), .B2(n6774), .A(n6968), .ZN(n6776) );
  NAND2_X1 U8414 ( .A1(n6776), .A2(n8302), .ZN(n6783) );
  INV_X1 U8415 ( .A(n6777), .ZN(n6927) );
  OR2_X1 U8416 ( .A1(n8404), .A2(n6778), .ZN(n6780) );
  OAI211_X1 U8417 ( .C1(n8382), .C2(n7439), .A(n6780), .B(n6779), .ZN(n6781)
         );
  AOI21_X1 U8418 ( .B1(n6927), .B2(n8406), .A(n6781), .ZN(n6782) );
  OAI211_X1 U8419 ( .C1(n10324), .C2(n8410), .A(n6783), .B(n6782), .ZN(
        P2_U3153) );
  INV_X1 U8420 ( .A(n6969), .ZN(n8423) );
  AOI21_X1 U8421 ( .B1(n8402), .B2(n8423), .A(n6784), .ZN(n6788) );
  INV_X1 U8422 ( .A(n6785), .ZN(n6786) );
  NAND2_X1 U8423 ( .A1(n8406), .A2(n6786), .ZN(n6787) );
  OAI211_X1 U8424 ( .C1(n6789), .C2(n8404), .A(n6788), .B(n6787), .ZN(n6795)
         );
  INV_X1 U8425 ( .A(n6790), .ZN(n6791) );
  AOI211_X1 U8426 ( .C1(n6793), .C2(n6792), .A(n8394), .B(n6791), .ZN(n6794)
         );
  AOI211_X1 U8427 ( .C1(n10322), .C2(n8390), .A(n6795), .B(n6794), .ZN(n6796)
         );
  INV_X1 U8428 ( .A(n6796), .ZN(P2_U3179) );
  OAI222_X1 U8429 ( .A1(P1_U3086), .A2(n5514), .B1(n10173), .B2(n6798), .C1(
        n6797), .C2(n8278), .ZN(P1_U3334) );
  OAI21_X1 U8430 ( .B1(n6800), .B2(n9490), .A(n6799), .ZN(n10244) );
  OAI21_X1 U8431 ( .B1(n5736), .B2(n6802), .A(n6801), .ZN(n10240) );
  OAI22_X1 U8432 ( .A1(n9769), .A2(n10240), .B1(n5736), .B2(n10026), .ZN(n6809) );
  INV_X1 U8433 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9656) );
  NAND2_X1 U8434 ( .A1(n5593), .A2(n9997), .ZN(n6803) );
  OAI21_X1 U8435 ( .B1(n6804), .B2(n10013), .A(n6803), .ZN(n6805) );
  AOI21_X1 U8436 ( .B1(n6806), .B2(n10009), .A(n6805), .ZN(n10241) );
  OAI21_X1 U8437 ( .B1(n9656), .B2(n9980), .A(n10241), .ZN(n6807) );
  MUX2_X1 U8438 ( .A(n6807), .B(P1_REG2_REG_2__SCAN_IN), .S(n9986), .Z(n6808)
         );
  AOI211_X1 U8439 ( .C1(n9976), .C2(n10244), .A(n6809), .B(n6808), .ZN(n6810)
         );
  INV_X1 U8440 ( .A(n6810), .ZN(P1_U3291) );
  OAI222_X1 U8441 ( .A1(P1_U3086), .A2(n9577), .B1(n10173), .B2(n6812), .C1(
        n6811), .C2(n8278), .ZN(P1_U3335) );
  OAI21_X1 U8442 ( .B1(n6814), .B2(n9498), .A(n6813), .ZN(n10270) );
  INV_X1 U8443 ( .A(n10270), .ZN(n6828) );
  INV_X1 U8444 ( .A(n6815), .ZN(n6819) );
  AOI21_X1 U8445 ( .B1(n6817), .B2(n9547), .A(n6816), .ZN(n6818) );
  NOR2_X1 U8446 ( .A1(n6819), .A2(n6818), .ZN(n6820) );
  OAI222_X1 U8447 ( .A1(n10013), .A2(n7327), .B1(n10011), .B2(n7041), .C1(
        n9938), .C2(n6820), .ZN(n10269) );
  OAI21_X1 U8448 ( .B1(n6822), .B2(n10265), .A(n6821), .ZN(n10267) );
  OAI22_X1 U8449 ( .A1(n10028), .A2(n5678), .B1(n7328), .B2(n9980), .ZN(n6823)
         );
  AOI21_X1 U8450 ( .B1(n7012), .B2(n6824), .A(n6823), .ZN(n6825) );
  OAI21_X1 U8451 ( .B1(n10267), .B2(n9769), .A(n6825), .ZN(n6826) );
  AOI21_X1 U8452 ( .B1(n10269), .B2(n10028), .A(n6826), .ZN(n6827) );
  OAI21_X1 U8453 ( .B1(n6828), .B2(n10030), .A(n6827), .ZN(P1_U3283) );
  NAND2_X1 U8454 ( .A1(n6829), .A2(n7684), .ZN(n6830) );
  XOR2_X1 U8455 ( .A(n7927), .B(n6830), .Z(n10348) );
  INV_X1 U8456 ( .A(n10348), .ZN(n10345) );
  XNOR2_X1 U8457 ( .A(n6831), .B(n7927), .ZN(n6832) );
  OAI222_X1 U8458 ( .A1(n10194), .A2(n7066), .B1(n10192), .B2(n7443), .C1(
        n10296), .C2(n6832), .ZN(n10346) );
  NAND2_X1 U8459 ( .A1(n10346), .A2(n8724), .ZN(n6835) );
  OAI22_X1 U8460 ( .A1(n8724), .A2(n6612), .B1(n7133), .B2(n10181), .ZN(n6833)
         );
  AOI21_X1 U8461 ( .B1(n10342), .B2(n8726), .A(n6833), .ZN(n6834) );
  OAI211_X1 U8462 ( .C1(n10345), .C2(n8729), .A(n6835), .B(n6834), .ZN(
        P2_U3223) );
  NAND2_X1 U8463 ( .A1(n7252), .A2(n9467), .ZN(n6839) );
  AOI22_X1 U8464 ( .A1(n9473), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n4494), .B2(
        n9699), .ZN(n6838) );
  OR2_X1 U8465 ( .A1(n7422), .A2(n7414), .ZN(n9411) );
  NAND2_X1 U8466 ( .A1(n7422), .A2(n7414), .ZN(n9553) );
  NAND2_X1 U8467 ( .A1(n9411), .A2(n9553), .ZN(n9502) );
  OAI21_X1 U8468 ( .B1(n6840), .B2(n9502), .A(n7074), .ZN(n6884) );
  INV_X1 U8469 ( .A(n6884), .ZN(n6861) );
  INV_X1 U8470 ( .A(n9502), .ZN(n6844) );
  AND2_X1 U8471 ( .A1(n9404), .A2(n9401), .ZN(n9551) );
  NAND2_X1 U8472 ( .A1(n6841), .A2(n9551), .ZN(n6842) );
  NAND2_X1 U8473 ( .A1(n6842), .A2(n9554), .ZN(n6843) );
  OAI21_X1 U8474 ( .B1(n6844), .B2(n6843), .A(n7087), .ZN(n6845) );
  NAND2_X1 U8475 ( .A1(n6845), .A2(n10009), .ZN(n6854) );
  NAND2_X1 U8476 ( .A1(n9476), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6852) );
  AND2_X1 U8477 ( .A1(n6847), .A2(n6846), .ZN(n6848) );
  NOR2_X1 U8478 ( .A1(n7081), .A2(n6848), .ZN(n9240) );
  NAND2_X1 U8479 ( .A1(n5720), .A2(n9240), .ZN(n6851) );
  NAND2_X1 U8480 ( .A1(n9477), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6850) );
  NAND2_X1 U8481 ( .A1(n4492), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6849) );
  NAND4_X1 U8482 ( .A1(n6852), .A2(n6851), .A3(n6850), .A4(n6849), .ZN(n9630)
         );
  AOI22_X1 U8483 ( .A1(n9632), .A2(n9997), .B1(n9999), .B2(n9630), .ZN(n6853)
         );
  NAND2_X1 U8484 ( .A1(n6854), .A2(n6853), .ZN(n6882) );
  INV_X1 U8485 ( .A(n7422), .ZN(n6858) );
  AOI211_X1 U8486 ( .C1(n7422), .C2(n6855), .A(n10266), .B(n7338), .ZN(n6883)
         );
  NAND2_X1 U8487 ( .A1(n6883), .A2(n10021), .ZN(n6857) );
  AOI22_X1 U8488 ( .A1(n9986), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7418), .B2(
        n10022), .ZN(n6856) );
  OAI211_X1 U8489 ( .C1(n6858), .C2(n10026), .A(n6857), .B(n6856), .ZN(n6859)
         );
  AOI21_X1 U8490 ( .B1(n10028), .B2(n6882), .A(n6859), .ZN(n6860) );
  OAI21_X1 U8491 ( .B1(n6861), .B2(n10030), .A(n6860), .ZN(P1_U3280) );
  OAI21_X1 U8492 ( .B1(n7061), .B2(n10379), .A(n6862), .ZN(n6937) );
  XNOR2_X1 U8493 ( .A(n7253), .B(n6937), .ZN(n6863) );
  NAND2_X1 U8494 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n6863), .ZN(n6938) );
  OAI21_X1 U8495 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n6863), .A(n6938), .ZN(
        n6864) );
  INV_X1 U8496 ( .A(n6864), .ZN(n6881) );
  NAND2_X1 U8497 ( .A1(P2_REG2_REG_13__SCAN_IN), .A2(n6866), .ZN(n6945) );
  OAI21_X1 U8498 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n6866), .A(n6945), .ZN(
        n6879) );
  NAND2_X1 U8499 ( .A1(n6874), .A2(n6873), .ZN(n6871) );
  INV_X1 U8500 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7051) );
  INV_X1 U8501 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7054) );
  MUX2_X1 U8502 ( .A(n7051), .B(n7054), .S(n8512), .Z(n6867) );
  NAND2_X1 U8503 ( .A1(n6867), .A2(n7253), .ZN(n6955) );
  INV_X1 U8504 ( .A(n6867), .ZN(n6868) );
  NAND2_X1 U8505 ( .A1(n6868), .A2(n6944), .ZN(n6869) );
  NAND2_X1 U8506 ( .A1(n6955), .A2(n6869), .ZN(n6872) );
  INV_X1 U8507 ( .A(n6872), .ZN(n6870) );
  NAND2_X1 U8508 ( .A1(n6871), .A2(n6870), .ZN(n6956) );
  NAND3_X1 U8509 ( .A1(n6874), .A2(n6873), .A3(n6872), .ZN(n6875) );
  AOI21_X1 U8510 ( .B1(n6956), .B2(n6875), .A(n8517), .ZN(n6878) );
  NAND2_X1 U8511 ( .A1(n8519), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n6876) );
  NAND2_X1 U8512 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7606) );
  OAI211_X1 U8513 ( .C1(n8522), .C2(n6944), .A(n6876), .B(n7606), .ZN(n6877)
         );
  AOI211_X1 U8514 ( .C1(n6879), .C2(n8526), .A(n6878), .B(n6877), .ZN(n6880)
         );
  OAI21_X1 U8515 ( .B1(n8529), .B2(n6881), .A(n6880), .ZN(P2_U3195) );
  AOI211_X1 U8516 ( .C1(n6884), .C2(n10276), .A(n6883), .B(n6882), .ZN(n6889)
         );
  AOI22_X1 U8517 ( .A1(n7422), .A2(n6885), .B1(P1_REG1_REG_13__SCAN_IN), .B2(
        n10290), .ZN(n6886) );
  OAI21_X1 U8518 ( .B1(n6889), .B2(n10290), .A(n6886), .ZN(P1_U3535) );
  INV_X1 U8519 ( .A(n10164), .ZN(n6887) );
  AOI22_X1 U8520 ( .A1(n7422), .A2(n6887), .B1(P1_REG0_REG_13__SCAN_IN), .B2(
        n10278), .ZN(n6888) );
  OAI21_X1 U8521 ( .B1(n6889), .B2(n10278), .A(n6888), .ZN(P1_U3492) );
  INV_X1 U8522 ( .A(n6892), .ZN(n6893) );
  NAND2_X1 U8523 ( .A1(n6893), .A2(SI_21_), .ZN(n6894) );
  NAND2_X1 U8524 ( .A1(n6895), .A2(n6894), .ZN(n6979) );
  MUX2_X1 U8525 ( .A(n8840), .B(n7991), .S(n7901), .Z(n6897) );
  INV_X1 U8526 ( .A(SI_22_), .ZN(n6896) );
  NAND2_X1 U8527 ( .A1(n6897), .A2(n6896), .ZN(n7180) );
  INV_X1 U8528 ( .A(n6897), .ZN(n6898) );
  NAND2_X1 U8529 ( .A1(n6898), .A2(SI_22_), .ZN(n6899) );
  NAND2_X1 U8530 ( .A1(n7180), .A2(n6899), .ZN(n6978) );
  XNOR2_X1 U8531 ( .A(n6979), .B(n6978), .ZN(n8085) );
  INV_X1 U8532 ( .A(n8085), .ZN(n7990) );
  OAI222_X1 U8533 ( .A1(n9222), .A2(n8840), .B1(n9220), .B2(n7990), .C1(
        P2_U3151), .C2(n7646), .ZN(P2_U3273) );
  NAND2_X1 U8534 ( .A1(n6747), .A2(n7681), .ZN(n6930) );
  NAND2_X1 U8535 ( .A1(n6930), .A2(n7922), .ZN(n6931) );
  NAND2_X1 U8536 ( .A1(n6931), .A2(n6900), .ZN(n6901) );
  XNOR2_X1 U8537 ( .A(n6901), .B(n7921), .ZN(n10330) );
  OR2_X1 U8538 ( .A1(n6903), .A2(n6902), .ZN(n6922) );
  NAND2_X1 U8539 ( .A1(n6922), .A2(n6904), .ZN(n6906) );
  AND2_X1 U8540 ( .A1(n6906), .A2(n6905), .ZN(n6907) );
  XNOR2_X1 U8541 ( .A(n6907), .B(n7921), .ZN(n6908) );
  OAI222_X1 U8542 ( .A1(n10194), .A2(n7443), .B1(n10192), .B2(n6969), .C1(
        n10296), .C2(n6908), .ZN(n10331) );
  NAND2_X1 U8543 ( .A1(n10331), .A2(n8724), .ZN(n6912) );
  INV_X1 U8544 ( .A(n6974), .ZN(n6909) );
  OAI22_X1 U8545 ( .A1(n8724), .A2(n6013), .B1(n6909), .B2(n10181), .ZN(n6910)
         );
  AOI21_X1 U8546 ( .B1(n8726), .B2(n10333), .A(n6910), .ZN(n6911) );
  OAI211_X1 U8547 ( .C1(n10330), .C2(n8729), .A(n6912), .B(n6911), .ZN(
        P2_U3225) );
  INV_X1 U8548 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n8846) );
  AOI211_X1 U8549 ( .C1(n6916), .C2(n6915), .A(n6914), .B(n6913), .ZN(n6918)
         );
  MUX2_X1 U8550 ( .A(n8846), .B(n6918), .S(n10280), .Z(n6917) );
  OAI21_X1 U8551 ( .B1(n6920), .B2(n10164), .A(n6917), .ZN(P1_U3486) );
  MUX2_X1 U8552 ( .A(n5852), .B(n6918), .S(n10293), .Z(n6919) );
  OAI21_X1 U8553 ( .B1(n6920), .B2(n10108), .A(n6919), .ZN(P1_U3533) );
  NAND2_X1 U8554 ( .A1(n6922), .A2(n6921), .ZN(n6923) );
  XNOR2_X1 U8555 ( .A(n6923), .B(n7687), .ZN(n6924) );
  NAND2_X1 U8556 ( .A1(n6924), .A2(n8706), .ZN(n6926) );
  AOI22_X1 U8557 ( .A1(n7441), .A2(n8703), .B1(n8701), .B2(n8424), .ZN(n6925)
         );
  NAND2_X1 U8558 ( .A1(n6926), .A2(n6925), .ZN(n10327) );
  AOI21_X1 U8559 ( .B1(n8709), .B2(n6927), .A(n10327), .ZN(n6928) );
  MUX2_X1 U8560 ( .A(n6929), .B(n6928), .S(n8724), .Z(n6936) );
  INV_X1 U8561 ( .A(n6930), .ZN(n6933) );
  INV_X1 U8562 ( .A(n6931), .ZN(n6932) );
  AOI21_X1 U8563 ( .B1(n6933), .B2(n7687), .A(n6932), .ZN(n10328) );
  AOI22_X1 U8564 ( .A1(n10328), .A2(n8670), .B1(n8726), .B2(n6934), .ZN(n6935)
         );
  NAND2_X1 U8565 ( .A1(n6936), .A2(n6935), .ZN(P2_U3226) );
  INV_X1 U8566 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7295) );
  AOI22_X1 U8567 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n6959), .B1(n7262), .B2(
        n7295), .ZN(n6941) );
  NAND2_X1 U8568 ( .A1(n6944), .A2(n6937), .ZN(n6939) );
  OAI21_X1 U8569 ( .B1(n6941), .B2(n6940), .A(n7157), .ZN(n6942) );
  INV_X1 U8570 ( .A(n6942), .ZN(n6964) );
  INV_X1 U8571 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7265) );
  AOI22_X1 U8572 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n6959), .B1(n7262), .B2(
        n7265), .ZN(n6948) );
  NAND2_X1 U8573 ( .A1(n6944), .A2(n6943), .ZN(n6946) );
  OAI21_X1 U8574 ( .B1(n6948), .B2(n6947), .A(n7167), .ZN(n6962) );
  NAND2_X1 U8575 ( .A1(n6956), .A2(n6955), .ZN(n6953) );
  MUX2_X1 U8576 ( .A(n7265), .B(n7295), .S(n8512), .Z(n6949) );
  NAND2_X1 U8577 ( .A1(n6949), .A2(n7262), .ZN(n7160) );
  INV_X1 U8578 ( .A(n6949), .ZN(n6950) );
  NAND2_X1 U8579 ( .A1(n6950), .A2(n6959), .ZN(n6951) );
  NAND2_X1 U8580 ( .A1(n7160), .A2(n6951), .ZN(n6954) );
  INV_X1 U8581 ( .A(n6954), .ZN(n6952) );
  NAND2_X1 U8582 ( .A1(n6953), .A2(n6952), .ZN(n7161) );
  NAND3_X1 U8583 ( .A1(n6956), .A2(n6955), .A3(n6954), .ZN(n6957) );
  AOI21_X1 U8584 ( .B1(n7161), .B2(n6957), .A(n8517), .ZN(n6961) );
  NAND2_X1 U8585 ( .A1(n8519), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n6958) );
  NAND2_X1 U8586 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8286) );
  OAI211_X1 U8587 ( .C1(n8522), .C2(n6959), .A(n6958), .B(n8286), .ZN(n6960)
         );
  AOI211_X1 U8588 ( .C1(n6962), .C2(n8526), .A(n6961), .B(n6960), .ZN(n6963)
         );
  OAI21_X1 U8589 ( .B1(n8529), .B2(n6964), .A(n6963), .ZN(P2_U3196) );
  INV_X1 U8590 ( .A(n6965), .ZN(n6966) );
  NAND2_X1 U8591 ( .A1(n6966), .A2(n6969), .ZN(n6967) );
  XNOR2_X1 U8592 ( .A(n10333), .B(n8258), .ZN(n7119) );
  INV_X1 U8593 ( .A(n7119), .ZN(n7440) );
  XNOR2_X1 U8594 ( .A(n7121), .B(n7440), .ZN(n7442) );
  XNOR2_X1 U8595 ( .A(n7442), .B(n7439), .ZN(n6977) );
  OR2_X1 U8596 ( .A1(n8404), .A2(n6969), .ZN(n6972) );
  INV_X1 U8597 ( .A(n6970), .ZN(n6971) );
  OAI211_X1 U8598 ( .C1(n8382), .C2(n7443), .A(n6972), .B(n6971), .ZN(n6973)
         );
  AOI21_X1 U8599 ( .B1(n6974), .B2(n8406), .A(n6973), .ZN(n6976) );
  NAND2_X1 U8600 ( .A1(n8390), .A2(n10333), .ZN(n6975) );
  OAI211_X1 U8601 ( .C1(n6977), .C2(n8394), .A(n6976), .B(n6975), .ZN(P2_U3161) );
  INV_X1 U8602 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n6980) );
  MUX2_X1 U8603 ( .A(n8788), .B(n6980), .S(n7901), .Z(n6982) );
  INV_X1 U8604 ( .A(SI_23_), .ZN(n6981) );
  NAND2_X1 U8605 ( .A1(n6982), .A2(n6981), .ZN(n7310) );
  INV_X1 U8606 ( .A(n6982), .ZN(n6983) );
  NAND2_X1 U8607 ( .A1(n6983), .A2(SI_23_), .ZN(n6984) );
  INV_X1 U8608 ( .A(n7995), .ZN(n6987) );
  OR2_X1 U8609 ( .A1(n6985), .A2(P1_U3086), .ZN(n9618) );
  INV_X1 U8610 ( .A(n9618), .ZN(n9610) );
  AOI21_X1 U8611 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n10171), .A(n9610), .ZN(
        n6986) );
  OAI21_X1 U8612 ( .B1(n6987), .B2(n10173), .A(n6986), .ZN(P1_U3332) );
  INV_X1 U8613 ( .A(n6989), .ZN(n6990) );
  NAND2_X1 U8614 ( .A1(n6996), .A2(n8208), .ZN(n6994) );
  OR2_X1 U8615 ( .A1(n7041), .A2(n8226), .ZN(n6993) );
  NAND2_X1 U8616 ( .A1(n6994), .A2(n6993), .ZN(n6995) );
  XNOR2_X1 U8617 ( .A(n6995), .B(n4495), .ZN(n7107) );
  NAND2_X1 U8618 ( .A1(n6996), .A2(n5521), .ZN(n6998) );
  OR2_X1 U8619 ( .A1(n7041), .A2(n5702), .ZN(n6997) );
  NAND2_X1 U8620 ( .A1(n6998), .A2(n6997), .ZN(n7004) );
  NAND2_X1 U8621 ( .A1(n7107), .A2(n7004), .ZN(n7319) );
  NAND2_X1 U8622 ( .A1(n7002), .A2(n8208), .ZN(n7000) );
  OR2_X1 U8623 ( .A1(n7113), .A2(n8226), .ZN(n6999) );
  NAND2_X1 U8624 ( .A1(n7000), .A2(n6999), .ZN(n7001) );
  XNOR2_X1 U8625 ( .A(n7001), .B(n8194), .ZN(n7105) );
  AOI22_X1 U8626 ( .A1(n9635), .A2(n8182), .B1(n7002), .B2(n5521), .ZN(n7037)
         );
  NOR2_X1 U8627 ( .A1(n7105), .A2(n7037), .ZN(n7003) );
  INV_X1 U8628 ( .A(n7107), .ZN(n7008) );
  INV_X1 U8629 ( .A(n7004), .ZN(n7106) );
  INV_X1 U8630 ( .A(n7319), .ZN(n7006) );
  INV_X1 U8631 ( .A(n7037), .ZN(n7005) );
  INV_X1 U8632 ( .A(n7105), .ZN(n7035) );
  NOR3_X1 U8633 ( .A1(n7006), .A2(n7005), .A3(n7035), .ZN(n7007) );
  AOI21_X1 U8634 ( .B1(n7008), .B2(n7106), .A(n7007), .ZN(n7017) );
  NAND2_X1 U8635 ( .A1(n7012), .A2(n8208), .ZN(n7010) );
  OR2_X1 U8636 ( .A1(n7013), .A2(n8226), .ZN(n7009) );
  NAND2_X1 U8637 ( .A1(n7010), .A2(n7009), .ZN(n7011) );
  XNOR2_X1 U8638 ( .A(n7011), .B(n4495), .ZN(n7322) );
  NAND2_X1 U8639 ( .A1(n7012), .A2(n5521), .ZN(n7015) );
  OR2_X1 U8640 ( .A1(n7013), .A2(n5702), .ZN(n7014) );
  NAND2_X1 U8641 ( .A1(n7015), .A2(n7014), .ZN(n7321) );
  NAND2_X1 U8642 ( .A1(n7031), .A2(n8208), .ZN(n7021) );
  OR2_X1 U8643 ( .A1(n7327), .A2(n8226), .ZN(n7020) );
  NAND2_X1 U8644 ( .A1(n7021), .A2(n7020), .ZN(n7022) );
  XNOR2_X1 U8645 ( .A(n7022), .B(n8194), .ZN(n7025) );
  NOR2_X1 U8646 ( .A1(n7327), .A2(n5702), .ZN(n7023) );
  AOI21_X1 U8647 ( .B1(n7031), .B2(n5521), .A(n7023), .ZN(n7024) );
  NOR2_X1 U8648 ( .A1(n7025), .A2(n7024), .ZN(n7229) );
  NAND2_X1 U8649 ( .A1(n7025), .A2(n7024), .ZN(n7228) );
  NOR2_X1 U8650 ( .A1(n7229), .A2(n4873), .ZN(n7026) );
  XNOR2_X1 U8651 ( .A(n7230), .B(n7026), .ZN(n7033) );
  AOI22_X1 U8652 ( .A1(n9357), .A2(n7027), .B1(n9334), .B2(n9634), .ZN(n7029)
         );
  OAI211_X1 U8653 ( .C1(n7420), .C2(n9345), .A(n7029), .B(n7028), .ZN(n7030)
         );
  AOI21_X1 U8654 ( .B1(n7031), .B2(n9363), .A(n7030), .ZN(n7032) );
  OAI21_X1 U8655 ( .B1(n7033), .B2(n9365), .A(n7032), .ZN(P1_U3236) );
  XNOR2_X1 U8656 ( .A(n7034), .B(n7035), .ZN(n7036) );
  NAND2_X1 U8657 ( .A1(n7036), .A2(n7037), .ZN(n7109) );
  OAI21_X1 U8658 ( .B1(n7037), .B2(n7036), .A(n7109), .ZN(n7038) );
  NAND2_X1 U8659 ( .A1(n7038), .A2(n9342), .ZN(n7046) );
  INV_X1 U8660 ( .A(n7039), .ZN(n7044) );
  INV_X1 U8661 ( .A(n7040), .ZN(n7042) );
  OAI22_X1 U8662 ( .A1(n9314), .A2(n7042), .B1(n7041), .B2(n9345), .ZN(n7043)
         );
  AOI211_X1 U8663 ( .C1(n9334), .C2(n9636), .A(n7044), .B(n7043), .ZN(n7045)
         );
  OAI211_X1 U8664 ( .C1(n7047), .C2(n9350), .A(n7046), .B(n7045), .ZN(P1_U3221) );
  NAND2_X1 U8665 ( .A1(n7995), .A2(n7048), .ZN(n7050) );
  NAND2_X1 U8666 ( .A1(n7049), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7988) );
  OAI211_X1 U8667 ( .C1(n8788), .C2(n9222), .A(n7050), .B(n7988), .ZN(P2_U3272) );
  NAND2_X1 U8668 ( .A1(n4814), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n7058) );
  OR2_X1 U8669 ( .A1(n7865), .A2(n7051), .ZN(n7057) );
  OR2_X1 U8670 ( .A1(n7052), .A2(n8996), .ZN(n7053) );
  NAND2_X1 U8671 ( .A1(n7052), .A2(n8996), .ZN(n7266) );
  AND2_X1 U8672 ( .A1(n7053), .A2(n7266), .ZN(n10182) );
  OR2_X1 U8673 ( .A1(n7288), .A2(n10182), .ZN(n7056) );
  OR2_X1 U8674 ( .A1(n6581), .A2(n7054), .ZN(n7055) );
  NAND4_X1 U8675 ( .A1(n7058), .A2(n7057), .A3(n7056), .A4(n7055), .ZN(n8420)
         );
  INV_X1 U8676 ( .A(n8420), .ZN(n8287) );
  INV_X1 U8677 ( .A(n7066), .ZN(n7458) );
  NAND2_X1 U8678 ( .A1(n7059), .A2(n7458), .ZN(n7279) );
  NAND2_X1 U8679 ( .A1(n7349), .A2(n7279), .ZN(n10185) );
  NAND2_X1 U8680 ( .A1(n7060), .A2(n7873), .ZN(n7063) );
  AOI22_X1 U8681 ( .A1(n7737), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7736), .B2(
        n7061), .ZN(n7062) );
  NAND2_X1 U8682 ( .A1(n7063), .A2(n7062), .ZN(n10362) );
  OR2_X1 U8683 ( .A1(n10362), .A2(n10191), .ZN(n10176) );
  NAND2_X1 U8684 ( .A1(n10362), .A2(n10191), .ZN(n7064) );
  NAND2_X1 U8685 ( .A1(n10176), .A2(n7064), .ZN(n7930) );
  XNOR2_X1 U8686 ( .A(n10185), .B(n7930), .ZN(n7065) );
  OAI222_X1 U8687 ( .A1(n10192), .A2(n7066), .B1(n10194), .B2(n8287), .C1(
        n7065), .C2(n10296), .ZN(n10360) );
  INV_X1 U8688 ( .A(n10360), .ZN(n7072) );
  OAI22_X1 U8689 ( .A1(n8724), .A2(n6736), .B1(n7460), .B2(n10181), .ZN(n7067)
         );
  AOI21_X1 U8690 ( .B1(n10362), .B2(n8726), .A(n7067), .ZN(n7071) );
  NAND2_X1 U8691 ( .A1(n7068), .A2(n7928), .ZN(n7069) );
  NAND2_X1 U8692 ( .A1(n7069), .A2(n7708), .ZN(n7272) );
  OR2_X1 U8693 ( .A1(n7272), .A2(n7930), .ZN(n10359) );
  NAND2_X1 U8694 ( .A1(n7272), .A2(n7930), .ZN(n10357) );
  NAND3_X1 U8695 ( .A1(n10359), .A2(n10357), .A3(n8670), .ZN(n7070) );
  OAI211_X1 U8696 ( .C1(n7072), .C2(n10198), .A(n7071), .B(n7070), .ZN(
        P2_U3221) );
  INV_X1 U8697 ( .A(n7414), .ZN(n9631) );
  NAND2_X1 U8698 ( .A1(n7261), .A2(n9467), .ZN(n7076) );
  AOI22_X1 U8699 ( .A1(n9473), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n8043), .B2(
        n9712), .ZN(n7075) );
  NAND2_X1 U8700 ( .A1(n10116), .A2(n9630), .ZN(n7078) );
  NAND2_X1 U8701 ( .A1(n7353), .A2(n9467), .ZN(n7080) );
  INV_X1 U8702 ( .A(n7500), .ZN(n7146) );
  AOI22_X1 U8703 ( .A1(n9473), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n4494), .B2(
        n7146), .ZN(n7079) );
  NAND2_X1 U8704 ( .A1(n9476), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n7086) );
  OR2_X1 U8705 ( .A1(n7081), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7082) );
  NAND2_X1 U8706 ( .A1(n7081), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7090) );
  AND2_X1 U8707 ( .A1(n7082), .A2(n7090), .ZN(n9356) );
  NAND2_X1 U8708 ( .A1(n5720), .A2(n9356), .ZN(n7085) );
  NAND2_X1 U8709 ( .A1(n9477), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n7084) );
  NAND2_X1 U8710 ( .A1(n4492), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n7083) );
  NAND4_X1 U8711 ( .A1(n7086), .A2(n7085), .A3(n7084), .A4(n7083), .ZN(n9629)
         );
  INV_X1 U8712 ( .A(n9629), .ZN(n9241) );
  OR2_X1 U8713 ( .A1(n9418), .A2(n9241), .ZN(n9561) );
  NAND2_X1 U8714 ( .A1(n9418), .A2(n9241), .ZN(n9557) );
  XNOR2_X1 U8715 ( .A(n7210), .B(n9505), .ZN(n7427) );
  INV_X1 U8716 ( .A(n7427), .ZN(n7104) );
  OR2_X1 U8717 ( .A1(n10116), .A2(n9361), .ZN(n9412) );
  NAND2_X1 U8718 ( .A1(n10116), .A2(n9361), .ZN(n9556) );
  NAND2_X1 U8719 ( .A1(n9412), .A2(n9556), .ZN(n9488) );
  NAND2_X1 U8720 ( .A1(n7088), .A2(n9505), .ZN(n7219) );
  OAI21_X1 U8721 ( .B1(n9505), .B2(n7088), .A(n7219), .ZN(n7089) );
  NAND2_X1 U8722 ( .A1(n7089), .A2(n10009), .ZN(n7097) );
  NAND2_X1 U8723 ( .A1(n7090), .A2(n9085), .ZN(n7091) );
  AND2_X1 U8724 ( .A1(n7213), .A2(n7091), .ZN(n9274) );
  NAND2_X1 U8725 ( .A1(n5720), .A2(n9274), .ZN(n7095) );
  NAND2_X1 U8726 ( .A1(n9476), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n7094) );
  NAND2_X1 U8727 ( .A1(n5599), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7093) );
  NAND2_X1 U8728 ( .A1(n4491), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n7092) );
  AOI22_X1 U8729 ( .A1(n9775), .A2(n9999), .B1(n9997), .B2(n9630), .ZN(n7096)
         );
  NAND2_X1 U8730 ( .A1(n7097), .A2(n7096), .ZN(n7425) );
  INV_X1 U8731 ( .A(n7339), .ZN(n7099) );
  NAND2_X1 U8732 ( .A1(n7339), .A2(n7432), .ZN(n7222) );
  INV_X1 U8733 ( .A(n7222), .ZN(n7098) );
  AOI211_X1 U8734 ( .C1(n9418), .C2(n7099), .A(n10266), .B(n7098), .ZN(n7426)
         );
  NAND2_X1 U8735 ( .A1(n7426), .A2(n10021), .ZN(n7101) );
  AOI22_X1 U8736 ( .A1(n9986), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9356), .B2(
        n10022), .ZN(n7100) );
  OAI211_X1 U8737 ( .C1(n7432), .C2(n10026), .A(n7101), .B(n7100), .ZN(n7102)
         );
  AOI21_X1 U8738 ( .B1(n10028), .B2(n7425), .A(n7102), .ZN(n7103) );
  OAI21_X1 U8739 ( .B1(n7104), .B2(n10030), .A(n7103), .ZN(P1_U3278) );
  NAND2_X1 U8740 ( .A1(n7034), .A2(n7105), .ZN(n7108) );
  AND2_X1 U8741 ( .A1(n7109), .A2(n7108), .ZN(n7111) );
  XNOR2_X1 U8742 ( .A(n7107), .B(n7106), .ZN(n7110) );
  NAND3_X1 U8743 ( .A1(n7109), .A2(n7110), .A3(n7108), .ZN(n7320) );
  OAI211_X1 U8744 ( .C1(n7111), .C2(n7110), .A(n9342), .B(n7320), .ZN(n7118)
         );
  INV_X1 U8745 ( .A(n7112), .ZN(n7114) );
  OAI22_X1 U8746 ( .A1(n9314), .A2(n7114), .B1(n7113), .B2(n9360), .ZN(n7115)
         );
  AOI211_X1 U8747 ( .C1(n9355), .C2(n9634), .A(n7116), .B(n7115), .ZN(n7117)
         );
  OAI211_X1 U8748 ( .C1(n4837), .C2(n9350), .A(n7118), .B(n7117), .ZN(P1_U3231) );
  XNOR2_X1 U8749 ( .A(n10334), .B(n8258), .ZN(n7444) );
  AOI22_X1 U8750 ( .A1(n7444), .A2(n7443), .B1(n7439), .B2(n7119), .ZN(n7120)
         );
  INV_X1 U8751 ( .A(n7444), .ZN(n7126) );
  NAND2_X1 U8752 ( .A1(n7440), .A2(n7441), .ZN(n7122) );
  NAND2_X1 U8753 ( .A1(n7122), .A2(n7443), .ZN(n7125) );
  INV_X1 U8754 ( .A(n7122), .ZN(n7124) );
  AOI22_X1 U8755 ( .A1(n7126), .A2(n7125), .B1(n7124), .B2(n7123), .ZN(n7127)
         );
  NAND2_X1 U8756 ( .A1(n7128), .A2(n7127), .ZN(n7399) );
  XNOR2_X1 U8757 ( .A(n10342), .B(n8258), .ZN(n7397) );
  XOR2_X1 U8758 ( .A(n7398), .B(n7397), .Z(n7136) );
  INV_X1 U8759 ( .A(n7129), .ZN(n7131) );
  NOR2_X1 U8760 ( .A1(n8404), .A2(n7443), .ZN(n7130) );
  AOI211_X1 U8761 ( .C1(n8402), .C2(n7458), .A(n7131), .B(n7130), .ZN(n7132)
         );
  OAI21_X1 U8762 ( .B1(n7133), .B2(n8291), .A(n7132), .ZN(n7134) );
  AOI21_X1 U8763 ( .B1(n10342), .B2(n8390), .A(n7134), .ZN(n7135) );
  OAI21_X1 U8764 ( .B1(n7136), .B2(n8394), .A(n7135), .ZN(P2_U3157) );
  NAND2_X1 U8765 ( .A1(n9712), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7137) );
  OAI21_X1 U8766 ( .B1(n9712), .B2(P1_REG2_REG_14__SCAN_IN), .A(n7137), .ZN(
        n7138) );
  INV_X1 U8767 ( .A(n7138), .ZN(n9720) );
  INV_X1 U8768 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7139) );
  XNOR2_X1 U8769 ( .A(n9699), .B(n7139), .ZN(n9702) );
  INV_X1 U8770 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7142) );
  INV_X1 U8771 ( .A(n7140), .ZN(n7141) );
  AOI21_X1 U8772 ( .B1(n7150), .B2(n7142), .A(n7141), .ZN(n9701) );
  NAND2_X1 U8773 ( .A1(n9702), .A2(n9701), .ZN(n9700) );
  NAND2_X1 U8774 ( .A1(n9699), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7143) );
  NAND2_X1 U8775 ( .A1(n9700), .A2(n7143), .ZN(n9719) );
  INV_X1 U8776 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7144) );
  AOI211_X1 U8777 ( .C1(n7145), .C2(n7144), .A(n7502), .B(n9752), .ZN(n7156)
         );
  INV_X1 U8778 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n8854) );
  NAND2_X1 U8779 ( .A1(n9755), .A2(n7146), .ZN(n7147) );
  NAND2_X1 U8780 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9358) );
  OAI211_X1 U8781 ( .C1(n8854), .C2(n9761), .A(n7147), .B(n9358), .ZN(n7155)
         );
  INV_X1 U8782 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n8879) );
  XNOR2_X1 U8783 ( .A(n9699), .B(n8879), .ZN(n9705) );
  INV_X1 U8784 ( .A(n7148), .ZN(n7149) );
  AOI21_X1 U8785 ( .B1(n7150), .B2(n10291), .A(n7149), .ZN(n9704) );
  NAND2_X1 U8786 ( .A1(n9705), .A2(n9704), .ZN(n9703) );
  NAND2_X1 U8787 ( .A1(n9699), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7151) );
  NAND2_X1 U8788 ( .A1(n9703), .A2(n7151), .ZN(n9715) );
  INV_X1 U8789 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7152) );
  XNOR2_X1 U8790 ( .A(n9712), .B(n7152), .ZN(n9716) );
  AOI21_X1 U8791 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9712), .A(n9713), .ZN(
        n7492) );
  XNOR2_X1 U8792 ( .A(n7500), .B(n7492), .ZN(n7153) );
  INV_X1 U8793 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n8835) );
  NOR2_X1 U8794 ( .A1(n8835), .A2(n7153), .ZN(n7493) );
  AOI211_X1 U8795 ( .C1(n7153), .C2(n8835), .A(n7493), .B(n9751), .ZN(n7154)
         );
  OR3_X1 U8796 ( .A1(n7156), .A2(n7155), .A3(n7154), .ZN(P1_U3258) );
  NAND2_X1 U8797 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n7158), .ZN(n7515) );
  OAI21_X1 U8798 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n7158), .A(n7515), .ZN(
        n7159) );
  INV_X1 U8799 ( .A(n7159), .ZN(n7172) );
  NAND2_X1 U8800 ( .A1(n7161), .A2(n7160), .ZN(n7163) );
  MUX2_X1 U8801 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8512), .Z(n7526) );
  XNOR2_X1 U8802 ( .A(n7526), .B(n7527), .ZN(n7162) );
  NAND2_X1 U8803 ( .A1(n7163), .A2(n7162), .ZN(n7530) );
  OAI21_X1 U8804 ( .B1(n7163), .B2(n7162), .A(n7530), .ZN(n7166) );
  NAND2_X1 U8805 ( .A1(n8519), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n7164) );
  NAND2_X1 U8806 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8400) );
  OAI211_X1 U8807 ( .C1(n8522), .C2(n7521), .A(n7164), .B(n8400), .ZN(n7165)
         );
  AOI21_X1 U8808 ( .B1(n7166), .B2(n8464), .A(n7165), .ZN(n7171) );
  NAND2_X1 U8809 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n7168), .ZN(n7522) );
  OAI21_X1 U8810 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n7168), .A(n7522), .ZN(
        n7169) );
  NAND2_X1 U8811 ( .A1(n7169), .A2(n8526), .ZN(n7170) );
  OAI211_X1 U8812 ( .C1(n7172), .C2(n8529), .A(n7171), .B(n7170), .ZN(P2_U3197) );
  MUX2_X1 U8813 ( .A(n7790), .B(n9073), .S(n7901), .Z(n7178) );
  INV_X1 U8814 ( .A(n7178), .ZN(n7173) );
  NAND2_X1 U8815 ( .A1(n7173), .A2(SI_24_), .ZN(n7311) );
  MUX2_X1 U8816 ( .A(n7811), .B(n7316), .S(n7901), .Z(n7175) );
  INV_X1 U8817 ( .A(SI_25_), .ZN(n7174) );
  NAND2_X1 U8818 ( .A1(n7175), .A2(n7174), .ZN(n7184) );
  INV_X1 U8819 ( .A(n7175), .ZN(n7176) );
  NAND2_X1 U8820 ( .A1(n7176), .A2(SI_25_), .ZN(n7177) );
  INV_X1 U8821 ( .A(n7186), .ZN(n7179) );
  NAND2_X1 U8822 ( .A1(n7178), .A2(n9065), .ZN(n7312) );
  AND2_X1 U8823 ( .A1(n7310), .A2(n7312), .ZN(n7244) );
  AND2_X1 U8824 ( .A1(n7180), .A2(n7185), .ZN(n7181) );
  NAND2_X1 U8825 ( .A1(n7183), .A2(n7182), .ZN(n7205) );
  INV_X1 U8826 ( .A(n7184), .ZN(n7190) );
  INV_X1 U8827 ( .A(n7185), .ZN(n7188) );
  AND2_X1 U8828 ( .A1(n7308), .A2(n7186), .ZN(n7187) );
  MUX2_X1 U8829 ( .A(n7823), .B(n9079), .S(n7901), .Z(n7192) );
  NAND2_X1 U8830 ( .A1(n7192), .A2(n7191), .ZN(n7196) );
  INV_X1 U8831 ( .A(n7192), .ZN(n7193) );
  NAND2_X1 U8832 ( .A1(n7193), .A2(SI_26_), .ZN(n7194) );
  NAND2_X1 U8833 ( .A1(n7205), .A2(n7195), .ZN(n7197) );
  INV_X1 U8834 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7833) );
  MUX2_X1 U8835 ( .A(n7833), .B(n8114), .S(n7901), .Z(n7199) );
  INV_X1 U8836 ( .A(SI_27_), .ZN(n7198) );
  NAND2_X1 U8837 ( .A1(n7199), .A2(n7198), .ZN(n7383) );
  INV_X1 U8838 ( .A(n7199), .ZN(n7200) );
  NAND2_X1 U8839 ( .A1(n7200), .A2(SI_27_), .ZN(n7201) );
  INV_X1 U8840 ( .A(n8200), .ZN(n8113) );
  AOI21_X1 U8841 ( .B1(n9216), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n7202), .ZN(
        n7203) );
  OAI21_X1 U8842 ( .B1(n8113), .B2(n9220), .A(n7203), .ZN(P2_U3268) );
  AND2_X1 U8843 ( .A1(n7205), .A2(n7204), .ZN(n7207) );
  INV_X1 U8844 ( .A(n8183), .ZN(n7241) );
  OAI222_X1 U8845 ( .A1(n7594), .A2(n7241), .B1(P2_U3151), .B2(n7208), .C1(
        n7823), .C2(n9222), .ZN(P2_U3269) );
  NAND2_X1 U8846 ( .A1(n7465), .A2(n9467), .ZN(n7212) );
  AOI22_X1 U8847 ( .A1(n9473), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n4494), .B2(
        n7584), .ZN(n7211) );
  OR2_X1 U8848 ( .A1(n10111), .A2(n10012), .ZN(n9562) );
  NAND2_X1 U8849 ( .A1(n10111), .A2(n10012), .ZN(n9582) );
  NAND2_X1 U8850 ( .A1(n9562), .A2(n9582), .ZN(n9777) );
  XNOR2_X1 U8851 ( .A(n9778), .B(n9777), .ZN(n10114) );
  AND2_X1 U8852 ( .A1(n7213), .A2(n8833), .ZN(n7214) );
  NOR2_X1 U8853 ( .A1(n8046), .A2(n7214), .ZN(n10023) );
  NAND2_X1 U8854 ( .A1(n10023), .A2(n5720), .ZN(n7218) );
  NAND2_X1 U8855 ( .A1(n4492), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n7217) );
  NAND2_X1 U8856 ( .A1(n9477), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7216) );
  NAND2_X1 U8857 ( .A1(n9476), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7215) );
  NAND2_X1 U8858 ( .A1(n7219), .A2(n9557), .ZN(n9581) );
  XNOR2_X1 U8859 ( .A(n9581), .B(n9777), .ZN(n7220) );
  OAI222_X1 U8860 ( .A1(n10013), .A2(n9779), .B1(n10011), .B2(n9241), .C1(
        n7220), .C2(n9938), .ZN(n10109) );
  INV_X1 U8861 ( .A(n10111), .ZN(n7225) );
  OR2_X1 U8862 ( .A1(n7222), .A2(n10111), .ZN(n10019) );
  INV_X1 U8863 ( .A(n10019), .ZN(n7221) );
  AOI211_X1 U8864 ( .C1(n10111), .C2(n7222), .A(n10266), .B(n7221), .ZN(n10110) );
  NAND2_X1 U8865 ( .A1(n10110), .A2(n10021), .ZN(n7224) );
  AOI22_X1 U8866 ( .A1(n9986), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9274), .B2(
        n10022), .ZN(n7223) );
  OAI211_X1 U8867 ( .C1(n7225), .C2(n10026), .A(n7224), .B(n7223), .ZN(n7226)
         );
  AOI21_X1 U8868 ( .B1(n10109), .B2(n10028), .A(n7226), .ZN(n7227) );
  OAI21_X1 U8869 ( .B1(n10114), .B2(n10030), .A(n7227), .ZN(P1_U3277) );
  NAND2_X1 U8870 ( .A1(n7238), .A2(n8208), .ZN(n7232) );
  OR2_X1 U8871 ( .A1(n7420), .A2(n8226), .ZN(n7231) );
  NAND2_X1 U8872 ( .A1(n7232), .A2(n7231), .ZN(n7233) );
  XNOR2_X1 U8873 ( .A(n7233), .B(n4495), .ZN(n7409) );
  AOI22_X1 U8874 ( .A1(n7238), .A2(n5521), .B1(n8182), .B2(n9632), .ZN(n7410)
         );
  XNOR2_X1 U8875 ( .A(n7409), .B(n7410), .ZN(n7412) );
  XOR2_X1 U8876 ( .A(n7413), .B(n7412), .Z(n7240) );
  AOI22_X1 U8877 ( .A1(n9357), .A2(n7234), .B1(n9334), .B2(n9633), .ZN(n7236)
         );
  OAI211_X1 U8878 ( .C1(n7414), .C2(n9345), .A(n7236), .B(n7235), .ZN(n7237)
         );
  AOI21_X1 U8879 ( .B1(n7238), .B2(n9363), .A(n7237), .ZN(n7239) );
  OAI21_X1 U8880 ( .B1(n7240), .B2(n9365), .A(n7239), .ZN(P1_U3224) );
  INV_X1 U8881 ( .A(n5247), .ZN(n7242) );
  OAI222_X1 U8882 ( .A1(n7242), .A2(P1_U3086), .B1(n10173), .B2(n7241), .C1(
        n9079), .C2(n8278), .ZN(P1_U3329) );
  AND2_X1 U8883 ( .A1(n7308), .A2(n7311), .ZN(n7243) );
  NAND2_X1 U8884 ( .A1(n7309), .A2(n7243), .ZN(n7247) );
  INV_X1 U8885 ( .A(n7311), .ZN(n7245) );
  OR2_X1 U8886 ( .A1(n7245), .A2(n7244), .ZN(n7246) );
  NAND2_X1 U8887 ( .A1(n7247), .A2(n7246), .ZN(n7249) );
  INV_X1 U8888 ( .A(n8167), .ZN(n7317) );
  INV_X1 U8889 ( .A(n7250), .ZN(n7251) );
  OAI222_X1 U8890 ( .A1(n7594), .A2(n7317), .B1(P2_U3151), .B2(n7251), .C1(
        n7811), .C2(n9222), .ZN(P2_U3270) );
  NAND2_X1 U8891 ( .A1(n7252), .A2(n7873), .ZN(n7255) );
  AOI22_X1 U8892 ( .A1(n7737), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7736), .B2(
        n7253), .ZN(n7254) );
  NAND2_X1 U8893 ( .A1(n7255), .A2(n7254), .ZN(n10180) );
  OR2_X1 U8894 ( .A1(n10180), .A2(n8287), .ZN(n7257) );
  INV_X1 U8895 ( .A(n7257), .ZN(n7256) );
  OR2_X1 U8896 ( .A1(n10180), .A2(n8420), .ZN(n7281) );
  NAND2_X1 U8897 ( .A1(n10180), .A2(n8420), .ZN(n7712) );
  NAND2_X1 U8898 ( .A1(n7281), .A2(n7712), .ZN(n10189) );
  OR2_X1 U8899 ( .A1(n7272), .A2(n7273), .ZN(n7260) );
  AND2_X1 U8900 ( .A1(n10176), .A2(n7257), .ZN(n7258) );
  OR2_X1 U8901 ( .A1(n7259), .A2(n7258), .ZN(n7274) );
  NAND2_X1 U8902 ( .A1(n7260), .A2(n7274), .ZN(n7277) );
  NAND2_X1 U8903 ( .A1(n7261), .A2(n7873), .ZN(n7264) );
  AOI22_X1 U8904 ( .A1(n7737), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7736), .B2(
        n7262), .ZN(n7263) );
  NAND2_X1 U8905 ( .A1(n4814), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n7271) );
  OR2_X1 U8906 ( .A1(n7865), .A2(n7265), .ZN(n7270) );
  NAND2_X1 U8907 ( .A1(n7266), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7267) );
  AND2_X1 U8908 ( .A1(n7286), .A2(n7267), .ZN(n8292) );
  OR2_X1 U8909 ( .A1(n7288), .A2(n8292), .ZN(n7269) );
  OR2_X1 U8910 ( .A1(n6581), .A2(n7295), .ZN(n7268) );
  OR2_X1 U8911 ( .A1(n8299), .A2(n10193), .ZN(n7718) );
  NAND2_X1 U8912 ( .A1(n8299), .A2(n10193), .ZN(n7717) );
  OR2_X1 U8913 ( .A1(n7714), .A2(n7274), .ZN(n7369) );
  AND2_X1 U8914 ( .A1(n7371), .A2(n7369), .ZN(n7275) );
  OAI21_X1 U8915 ( .B1(n7277), .B2(n7276), .A(n7275), .ZN(n7307) );
  INV_X1 U8916 ( .A(n7281), .ZN(n7710) );
  NAND2_X1 U8917 ( .A1(n10362), .A2(n8421), .ZN(n10186) );
  AND2_X1 U8918 ( .A1(n7712), .A2(n10186), .ZN(n7278) );
  OR2_X1 U8919 ( .A1(n7710), .A2(n7278), .ZN(n7280) );
  AND2_X1 U8920 ( .A1(n7279), .A2(n7280), .ZN(n7347) );
  NAND2_X1 U8921 ( .A1(n7349), .A2(n7347), .ZN(n7284) );
  INV_X1 U8922 ( .A(n7280), .ZN(n7283) );
  OR2_X1 U8923 ( .A1(n10362), .A2(n8421), .ZN(n10184) );
  AND2_X1 U8924 ( .A1(n10184), .A2(n7281), .ZN(n7282) );
  OR2_X1 U8925 ( .A1(n7283), .A2(n7282), .ZN(n7350) );
  NAND2_X1 U8926 ( .A1(n7284), .A2(n7350), .ZN(n7285) );
  XNOR2_X1 U8927 ( .A(n7285), .B(n7714), .ZN(n7294) );
  NAND2_X1 U8928 ( .A1(n4814), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n7293) );
  INV_X1 U8929 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7388) );
  OR2_X1 U8930 ( .A1(n7865), .A2(n7388), .ZN(n7292) );
  AND2_X1 U8931 ( .A1(n7286), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7287) );
  NOR2_X1 U8932 ( .A1(n7359), .A2(n7287), .ZN(n8399) );
  OR2_X1 U8933 ( .A1(n7288), .A2(n8399), .ZN(n7291) );
  INV_X1 U8934 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7289) );
  OR2_X1 U8935 ( .A1(n6581), .A2(n7289), .ZN(n7290) );
  AOI222_X1 U8936 ( .A1(n8706), .A2(n7294), .B1(n8418), .B2(n8703), .C1(n8420), 
        .C2(n8701), .ZN(n7301) );
  MUX2_X1 U8937 ( .A(n7295), .B(n7301), .S(n10381), .Z(n7297) );
  NAND2_X1 U8938 ( .A1(n8299), .A2(n8768), .ZN(n7296) );
  OAI211_X1 U8939 ( .C1(n8775), .C2(n7307), .A(n7297), .B(n7296), .ZN(P2_U3473) );
  INV_X1 U8940 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7298) );
  MUX2_X1 U8941 ( .A(n7298), .B(n7301), .S(n10364), .Z(n7300) );
  NAND2_X1 U8942 ( .A1(n8299), .A2(n9204), .ZN(n7299) );
  OAI211_X1 U8943 ( .C1(n7307), .C2(n9212), .A(n7300), .B(n7299), .ZN(P2_U3432) );
  INV_X1 U8944 ( .A(n7301), .ZN(n7304) );
  INV_X1 U8945 ( .A(n8299), .ZN(n7302) );
  OAI22_X1 U8946 ( .A1(n7302), .A2(n10183), .B1(n8292), .B2(n10181), .ZN(n7303) );
  OAI21_X1 U8947 ( .B1(n7304), .B2(n7303), .A(n8724), .ZN(n7306) );
  NAND2_X1 U8948 ( .A1(n10198), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7305) );
  OAI211_X1 U8949 ( .C1(n7307), .C2(n8729), .A(n7306), .B(n7305), .ZN(P2_U3219) );
  AND2_X1 U8950 ( .A1(n7312), .A2(n7311), .ZN(n7313) );
  INV_X1 U8951 ( .A(n8149), .ZN(n7396) );
  OAI222_X1 U8952 ( .A1(n7315), .A2(P1_U3086), .B1(n10173), .B2(n7396), .C1(
        n9073), .C2(n8278), .ZN(P1_U3331) );
  OAI222_X1 U8953 ( .A1(n7318), .A2(P1_U3086), .B1(n10173), .B2(n7317), .C1(
        n7316), .C2(n8278), .ZN(P1_U3330) );
  NAND2_X1 U8954 ( .A1(n7320), .A2(n7319), .ZN(n7324) );
  XNOR2_X1 U8955 ( .A(n7322), .B(n7321), .ZN(n7323) );
  XNOR2_X1 U8956 ( .A(n7324), .B(n7323), .ZN(n7325) );
  NAND2_X1 U8957 ( .A1(n7325), .A2(n9342), .ZN(n7332) );
  INV_X1 U8958 ( .A(n7326), .ZN(n7330) );
  OAI22_X1 U8959 ( .A1(n9314), .A2(n7328), .B1(n7327), .B2(n9345), .ZN(n7329)
         );
  AOI211_X1 U8960 ( .C1(n9334), .C2(n4836), .A(n7330), .B(n7329), .ZN(n7331)
         );
  OAI211_X1 U8961 ( .C1(n10265), .C2(n9350), .A(n7332), .B(n7331), .ZN(
        P1_U3217) );
  XNOR2_X1 U8962 ( .A(n7333), .B(n9488), .ZN(n7342) );
  AOI211_X1 U8963 ( .C1(n9488), .C2(n7334), .A(n9938), .B(n4560), .ZN(n7336)
         );
  OAI22_X1 U8964 ( .A1(n9241), .A2(n10013), .B1(n7414), .B2(n10011), .ZN(n7335) );
  AOI211_X1 U8965 ( .C1(n7342), .C2(n7337), .A(n7336), .B(n7335), .ZN(n10119)
         );
  INV_X1 U8966 ( .A(n7338), .ZN(n7340) );
  AOI211_X1 U8967 ( .C1(n10116), .C2(n7340), .A(n10266), .B(n7339), .ZN(n10115) );
  AOI22_X1 U8968 ( .A1(n9986), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9240), .B2(
        n10022), .ZN(n7341) );
  OAI21_X1 U8969 ( .B1(n9247), .B2(n10026), .A(n7341), .ZN(n7345) );
  INV_X1 U8970 ( .A(n7342), .ZN(n10121) );
  NOR2_X1 U8971 ( .A1(n10121), .A2(n7343), .ZN(n7344) );
  AOI211_X1 U8972 ( .C1(n10115), .C2(n10021), .A(n7345), .B(n7344), .ZN(n7346)
         );
  OAI21_X1 U8973 ( .B1(n9986), .B2(n10119), .A(n7346), .ZN(P1_U3279) );
  AND2_X1 U8974 ( .A1(n7347), .A2(n7714), .ZN(n7348) );
  OR2_X1 U8975 ( .A1(n7276), .A2(n7350), .ZN(n7351) );
  INV_X1 U8976 ( .A(n10193), .ZN(n8419) );
  OR2_X1 U8977 ( .A1(n8299), .A2(n8419), .ZN(n7352) );
  NAND2_X1 U8978 ( .A1(n7353), .A2(n7873), .ZN(n7355) );
  AOI22_X1 U8979 ( .A1(n7737), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n7736), .B2(
        n7527), .ZN(n7354) );
  NAND2_X1 U8980 ( .A1(n8393), .A2(n8329), .ZN(n7356) );
  NAND2_X1 U8981 ( .A1(n7357), .A2(n7932), .ZN(n7358) );
  NAND3_X1 U8982 ( .A1(n7471), .A2(n8706), .A3(n7358), .ZN(n7367) );
  NOR2_X1 U8983 ( .A1(n7359), .A2(n7536), .ZN(n7360) );
  OR2_X1 U8984 ( .A1(n7474), .A2(n7360), .ZN(n8326) );
  NAND2_X1 U8985 ( .A1(n7861), .A2(n8326), .ZN(n7364) );
  INV_X1 U8986 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n7483) );
  OR2_X1 U8987 ( .A1(n7841), .A2(n7483), .ZN(n7363) );
  INV_X1 U8988 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8457) );
  OR2_X1 U8989 ( .A1(n7865), .A2(n8457), .ZN(n7362) );
  OR2_X1 U8990 ( .A1(n6581), .A2(n9090), .ZN(n7361) );
  OAI22_X1 U8991 ( .A1(n10193), .A2(n10192), .B1(n8345), .B2(n10194), .ZN(
        n7365) );
  INV_X1 U8992 ( .A(n7365), .ZN(n7366) );
  NAND2_X1 U8993 ( .A1(n7367), .A2(n7366), .ZN(n7387) );
  MUX2_X1 U8994 ( .A(n7387), .B(P2_REG1_REG_15__SCAN_IN), .S(n10378), .Z(n7368) );
  INV_X1 U8995 ( .A(n7368), .ZN(n7376) );
  AND2_X1 U8996 ( .A1(n7369), .A2(n7718), .ZN(n7370) );
  OR2_X1 U8997 ( .A1(n7372), .A2(n7932), .ZN(n7373) );
  AND2_X1 U8998 ( .A1(n7464), .A2(n7373), .ZN(n7392) );
  INV_X1 U8999 ( .A(n8775), .ZN(n7374) );
  AOI22_X1 U9000 ( .A1(n7392), .A2(n7374), .B1(n8768), .B2(n8393), .ZN(n7375)
         );
  NAND2_X1 U9001 ( .A1(n7376), .A2(n7375), .ZN(P2_U3474) );
  MUX2_X1 U9002 ( .A(n7387), .B(P2_REG0_REG_15__SCAN_IN), .S(n10366), .Z(n7377) );
  INV_X1 U9003 ( .A(n7377), .ZN(n7380) );
  INV_X1 U9004 ( .A(n9212), .ZN(n7378) );
  AOI22_X1 U9005 ( .A1(n7392), .A2(n7378), .B1(n9204), .B2(n8393), .ZN(n7379)
         );
  NAND2_X1 U9006 ( .A1(n7380), .A2(n7379), .ZN(P2_U3435) );
  NAND2_X1 U9007 ( .A1(n7382), .A2(n7381), .ZN(n7384) );
  INV_X1 U9008 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7628) );
  MUX2_X1 U9009 ( .A(n7869), .B(n7628), .S(n7901), .Z(n7590) );
  XNOR2_X1 U9010 ( .A(n7590), .B(SI_28_), .ZN(n7587) );
  XNOR2_X1 U9011 ( .A(n7588), .B(n7587), .ZN(n8216) );
  INV_X1 U9012 ( .A(n8216), .ZN(n7627) );
  AOI21_X1 U9013 ( .B1(n9216), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n7385), .ZN(
        n7386) );
  OAI21_X1 U9014 ( .B1(n7627), .B2(n9220), .A(n7386), .ZN(P2_U3267) );
  INV_X1 U9015 ( .A(n7387), .ZN(n7389) );
  MUX2_X1 U9016 ( .A(n7389), .B(n7388), .S(n10198), .Z(n7394) );
  NAND2_X1 U9017 ( .A1(n8393), .A2(n8726), .ZN(n7390) );
  OAI21_X1 U9018 ( .B1(n8399), .B2(n10181), .A(n7390), .ZN(n7391) );
  AOI21_X1 U9019 ( .B1(n7392), .B2(n8670), .A(n7391), .ZN(n7393) );
  NAND2_X1 U9020 ( .A1(n7394), .A2(n7393), .ZN(P2_U3218) );
  OAI222_X1 U9021 ( .A1(n7594), .A2(n7396), .B1(P2_U3151), .B2(n7395), .C1(
        n7790), .C2(n9222), .ZN(P2_U3271) );
  XNOR2_X1 U9022 ( .A(n7928), .B(n8139), .ZN(n7451) );
  INV_X1 U9023 ( .A(n7451), .ZN(n7400) );
  NAND2_X1 U9024 ( .A1(n7401), .A2(n7400), .ZN(n7453) );
  OAI211_X1 U9025 ( .C1(n7401), .C2(n7400), .A(n8302), .B(n7453), .ZN(n7408)
         );
  AOI21_X1 U9026 ( .B1(n8402), .B2(n8421), .A(n7402), .ZN(n7403) );
  OAI21_X1 U9027 ( .B1(n7404), .B2(n8404), .A(n7403), .ZN(n7405) );
  AOI21_X1 U9028 ( .B1(n7406), .B2(n8406), .A(n7405), .ZN(n7407) );
  OAI211_X1 U9029 ( .C1(n10353), .C2(n8410), .A(n7408), .B(n7407), .ZN(
        P2_U3176) );
  INV_X1 U9030 ( .A(n7409), .ZN(n7411) );
  AOI22_X1 U9031 ( .A1(n7422), .A2(n5521), .B1(n8182), .B2(n9631), .ZN(n8006)
         );
  NAND2_X1 U9032 ( .A1(n7422), .A2(n8208), .ZN(n7416) );
  OR2_X1 U9033 ( .A1(n7414), .A2(n8226), .ZN(n7415) );
  NAND2_X1 U9034 ( .A1(n7416), .A2(n7415), .ZN(n7417) );
  XNOR2_X1 U9035 ( .A(n7417), .B(n4495), .ZN(n8008) );
  XOR2_X1 U9036 ( .A(n8006), .B(n8008), .Z(n8009) );
  XOR2_X1 U9037 ( .A(n8010), .B(n8009), .Z(n7424) );
  AOI22_X1 U9038 ( .A1(n9357), .A2(n7418), .B1(n9355), .B2(n9630), .ZN(n7419)
         );
  NAND2_X1 U9039 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n9696) );
  OAI211_X1 U9040 ( .C1(n7420), .C2(n9360), .A(n7419), .B(n9696), .ZN(n7421)
         );
  AOI21_X1 U9041 ( .B1(n7422), .B2(n9363), .A(n7421), .ZN(n7423) );
  OAI21_X1 U9042 ( .B1(n7424), .B2(n9365), .A(n7423), .ZN(P1_U3234) );
  AOI211_X1 U9043 ( .C1(n7427), .C2(n10276), .A(n7426), .B(n7425), .ZN(n7429)
         );
  MUX2_X1 U9044 ( .A(n8835), .B(n7429), .S(n10293), .Z(n7428) );
  OAI21_X1 U9045 ( .B1(n7432), .B2(n10108), .A(n7428), .ZN(P1_U3537) );
  INV_X1 U9046 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n7430) );
  MUX2_X1 U9047 ( .A(n7430), .B(n7429), .S(n10280), .Z(n7431) );
  OAI21_X1 U9048 ( .B1(n7432), .B2(n10164), .A(n7431), .ZN(P1_U3498) );
  INV_X1 U9049 ( .A(n7433), .ZN(n7434) );
  AOI21_X1 U9050 ( .B1(n8402), .B2(n8422), .A(n7434), .ZN(n7438) );
  INV_X1 U9051 ( .A(n7435), .ZN(n7436) );
  NAND2_X1 U9052 ( .A1(n8406), .A2(n7436), .ZN(n7437) );
  OAI211_X1 U9053 ( .C1(n7439), .C2(n8404), .A(n7438), .B(n7437), .ZN(n7449)
         );
  OAI22_X1 U9054 ( .A1(n7442), .A2(n7441), .B1(n7121), .B2(n7440), .ZN(n7446)
         );
  XNOR2_X1 U9055 ( .A(n7444), .B(n7443), .ZN(n7445) );
  XNOR2_X1 U9056 ( .A(n7446), .B(n7445), .ZN(n7447) );
  NOR2_X1 U9057 ( .A1(n7447), .A2(n8394), .ZN(n7448) );
  AOI211_X1 U9058 ( .C1(n10334), .C2(n8390), .A(n7449), .B(n7448), .ZN(n7450)
         );
  INV_X1 U9059 ( .A(n7450), .ZN(P2_U3171) );
  NAND2_X1 U9060 ( .A1(n7451), .A2(n7458), .ZN(n7452) );
  XNOR2_X1 U9061 ( .A(n10362), .B(n8139), .ZN(n7601) );
  XNOR2_X1 U9062 ( .A(n7601), .B(n10191), .ZN(n7454) );
  XNOR2_X1 U9063 ( .A(n7602), .B(n7454), .ZN(n7463) );
  INV_X1 U9064 ( .A(n7455), .ZN(n7457) );
  NOR2_X1 U9065 ( .A1(n8382), .A2(n8287), .ZN(n7456) );
  AOI211_X1 U9066 ( .C1(n8379), .C2(n7458), .A(n7457), .B(n7456), .ZN(n7459)
         );
  OAI21_X1 U9067 ( .B1(n7460), .B2(n8291), .A(n7459), .ZN(n7461) );
  AOI21_X1 U9068 ( .B1(n10362), .B2(n8390), .A(n7461), .ZN(n7462) );
  OAI21_X1 U9069 ( .B1(n7463), .B2(n8394), .A(n7462), .ZN(P2_U3164) );
  NAND2_X1 U9070 ( .A1(n7464), .A2(n7724), .ZN(n7468) );
  NAND2_X1 U9071 ( .A1(n7465), .A2(n7873), .ZN(n7467) );
  AOI22_X1 U9072 ( .A1(n7737), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7736), .B2(
        n8458), .ZN(n7466) );
  NAND2_X1 U9073 ( .A1(n8331), .A2(n8345), .ZN(n7729) );
  NAND2_X1 U9074 ( .A1(n7468), .A2(n7470), .ZN(n7548) );
  OAI21_X1 U9075 ( .B1(n7468), .B2(n7470), .A(n7548), .ZN(n7491) );
  NAND2_X1 U9076 ( .A1(n8393), .A2(n8418), .ZN(n7469) );
  INV_X1 U9077 ( .A(n7470), .ZN(n7934) );
  NAND3_X1 U9078 ( .A1(n7471), .A2(n7470), .A3(n7469), .ZN(n7472) );
  NAND3_X1 U9079 ( .A1(n7552), .A2(n8706), .A3(n7472), .ZN(n7482) );
  OR2_X1 U9080 ( .A1(n7474), .A2(n7473), .ZN(n7475) );
  NAND2_X1 U9081 ( .A1(n7554), .A2(n7475), .ZN(n8342) );
  NAND2_X1 U9082 ( .A1(n8342), .A2(n7861), .ZN(n7479) );
  INV_X1 U9083 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n7567) );
  OR2_X1 U9084 ( .A1(n7865), .A2(n7567), .ZN(n7478) );
  INV_X1 U9085 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n7571) );
  OR2_X1 U9086 ( .A1(n6581), .A2(n7571), .ZN(n7477) );
  NAND2_X1 U9087 ( .A1(n4814), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n7476) );
  OAI22_X1 U9088 ( .A1(n8721), .A2(n10194), .B1(n8329), .B2(n10192), .ZN(n7480) );
  INV_X1 U9089 ( .A(n7480), .ZN(n7481) );
  MUX2_X1 U9090 ( .A(n7488), .B(n7483), .S(n10366), .Z(n7485) );
  NAND2_X1 U9091 ( .A1(n8331), .A2(n9204), .ZN(n7484) );
  OAI211_X1 U9092 ( .C1(n7491), .C2(n9212), .A(n7485), .B(n7484), .ZN(P2_U3438) );
  MUX2_X1 U9093 ( .A(n7488), .B(n8457), .S(n10198), .Z(n7487) );
  AOI22_X1 U9094 ( .A1(n8331), .A2(n8726), .B1(n8709), .B2(n8326), .ZN(n7486)
         );
  OAI211_X1 U9095 ( .C1(n7491), .C2(n8729), .A(n7487), .B(n7486), .ZN(P2_U3217) );
  MUX2_X1 U9096 ( .A(n9090), .B(n7488), .S(n10381), .Z(n7490) );
  NAND2_X1 U9097 ( .A1(n8331), .A2(n8768), .ZN(n7489) );
  OAI211_X1 U9098 ( .C1(n8775), .C2(n7491), .A(n7490), .B(n7489), .ZN(P2_U3475) );
  INV_X1 U9099 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10106) );
  XNOR2_X1 U9100 ( .A(n9735), .B(n10106), .ZN(n9726) );
  NOR2_X1 U9101 ( .A1(n7492), .A2(n7500), .ZN(n7494) );
  NOR2_X1 U9102 ( .A1(n7494), .A2(n7493), .ZN(n7575) );
  INV_X1 U9103 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7495) );
  XNOR2_X1 U9104 ( .A(n7584), .B(n7495), .ZN(n7576) );
  NAND2_X1 U9105 ( .A1(n7575), .A2(n7576), .ZN(n7498) );
  NAND2_X1 U9106 ( .A1(n7496), .A2(n7495), .ZN(n7497) );
  NAND2_X1 U9107 ( .A1(n7498), .A2(n7497), .ZN(n9727) );
  XOR2_X1 U9108 ( .A(n9726), .B(n9727), .Z(n7513) );
  INV_X1 U9109 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n7499) );
  XNOR2_X1 U9110 ( .A(n9735), .B(n7499), .ZN(n7506) );
  NOR2_X1 U9111 ( .A1(n7501), .A2(n7500), .ZN(n7503) );
  XNOR2_X1 U9112 ( .A(n7584), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n7580) );
  OR2_X1 U9113 ( .A1(n7581), .A2(n7580), .ZN(n7578) );
  NAND2_X1 U9114 ( .A1(n7584), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7504) );
  AND2_X1 U9115 ( .A1(n7578), .A2(n7504), .ZN(n7505) );
  NAND2_X1 U9116 ( .A1(n7505), .A2(n7506), .ZN(n9737) );
  OAI21_X1 U9117 ( .B1(n7506), .B2(n7505), .A(n9737), .ZN(n7511) );
  NAND2_X1 U9118 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9284) );
  NAND2_X1 U9119 ( .A1(n9644), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n7507) );
  OAI211_X1 U9120 ( .C1(n7509), .C2(n7508), .A(n9284), .B(n7507), .ZN(n7510)
         );
  AOI21_X1 U9121 ( .B1(n7511), .B2(n9740), .A(n7510), .ZN(n7512) );
  OAI21_X1 U9122 ( .B1(n9751), .B2(n7513), .A(n7512), .ZN(P1_U3260) );
  AOI22_X1 U9123 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n7538), .B1(n8458), .B2(
        n9090), .ZN(n7518) );
  NAND2_X1 U9124 ( .A1(n7521), .A2(n7514), .ZN(n7516) );
  NAND2_X1 U9125 ( .A1(n7516), .A2(n7515), .ZN(n7517) );
  NAND2_X1 U9126 ( .A1(n7518), .A2(n7517), .ZN(n8453) );
  OAI21_X1 U9127 ( .B1(n7518), .B2(n7517), .A(n8453), .ZN(n7519) );
  INV_X1 U9128 ( .A(n7519), .ZN(n7543) );
  AOI22_X1 U9129 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n7538), .B1(n8458), .B2(
        n8457), .ZN(n7525) );
  NAND2_X1 U9130 ( .A1(n7521), .A2(n7520), .ZN(n7523) );
  NAND2_X1 U9131 ( .A1(n7523), .A2(n7522), .ZN(n7524) );
  NAND2_X1 U9132 ( .A1(n7525), .A2(n7524), .ZN(n8456) );
  OAI21_X1 U9133 ( .B1(n7525), .B2(n7524), .A(n8456), .ZN(n7541) );
  INV_X1 U9134 ( .A(n7526), .ZN(n7528) );
  NAND2_X1 U9135 ( .A1(n7528), .A2(n7527), .ZN(n7529) );
  NAND2_X1 U9136 ( .A1(n7530), .A2(n7529), .ZN(n7532) );
  MUX2_X1 U9137 ( .A(n8457), .B(n9090), .S(n8512), .Z(n7531) );
  NAND2_X1 U9138 ( .A1(n7532), .A2(n7531), .ZN(n8460) );
  OR2_X1 U9139 ( .A1(n7532), .A2(n7531), .ZN(n7533) );
  NAND2_X1 U9140 ( .A1(n8460), .A2(n7533), .ZN(n7534) );
  OR2_X1 U9141 ( .A1(n7534), .A2(n7538), .ZN(n8461) );
  NAND2_X1 U9142 ( .A1(n7534), .A2(n7538), .ZN(n7535) );
  AOI21_X1 U9143 ( .B1(n8461), .B2(n7535), .A(n8517), .ZN(n7540) );
  NOR2_X1 U9144 ( .A1(n7536), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8325) );
  AOI21_X1 U9145 ( .B1(n8519), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8325), .ZN(
        n7537) );
  OAI21_X1 U9146 ( .B1(n7538), .B2(n8522), .A(n7537), .ZN(n7539) );
  AOI211_X1 U9147 ( .C1(n7541), .C2(n8526), .A(n7540), .B(n7539), .ZN(n7542)
         );
  OAI21_X1 U9148 ( .B1(n8529), .B2(n7543), .A(n7542), .ZN(P2_U3198) );
  NAND2_X1 U9149 ( .A1(n7548), .A2(n7726), .ZN(n7546) );
  NAND2_X1 U9150 ( .A1(n8023), .A2(n7873), .ZN(n7545) );
  AOI22_X1 U9151 ( .A1(n7737), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7736), .B2(
        n8477), .ZN(n7544) );
  NAND2_X2 U9152 ( .A1(n7545), .A2(n7544), .ZN(n8539) );
  OR2_X1 U9153 ( .A1(n8539), .A2(n8721), .ZN(n7730) );
  NAND2_X1 U9154 ( .A1(n8539), .A2(n8721), .ZN(n7945) );
  NAND2_X1 U9155 ( .A1(n7730), .A2(n7945), .ZN(n7550) );
  NAND2_X1 U9156 ( .A1(n7546), .A2(n7550), .ZN(n7549) );
  NOR2_X1 U9157 ( .A1(n7550), .A2(n4776), .ZN(n7547) );
  INV_X1 U9158 ( .A(n8345), .ZN(n8417) );
  NAND2_X1 U9159 ( .A1(n8331), .A2(n8417), .ZN(n7551) );
  INV_X1 U9160 ( .A(n7550), .ZN(n7936) );
  NAND3_X1 U9161 ( .A1(n7552), .A2(n7936), .A3(n7551), .ZN(n7553) );
  NAND3_X1 U9162 ( .A1(n8541), .A2(n8706), .A3(n7553), .ZN(n7563) );
  NAND2_X1 U9163 ( .A1(n7554), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n7555) );
  NAND2_X1 U9164 ( .A1(n7740), .A2(n7555), .ZN(n8722) );
  NAND2_X1 U9165 ( .A1(n8722), .A2(n7861), .ZN(n7560) );
  INV_X1 U9166 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9210) );
  OR2_X1 U9167 ( .A1(n7841), .A2(n9210), .ZN(n7557) );
  INV_X1 U9168 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8876) );
  OR2_X1 U9169 ( .A1(n7865), .A2(n8876), .ZN(n7556) );
  AND2_X1 U9170 ( .A1(n7557), .A2(n7556), .ZN(n7559) );
  NAND2_X1 U9171 ( .A1(n7862), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n7558) );
  OAI22_X1 U9172 ( .A1(n8341), .A2(n10194), .B1(n8345), .B2(n10192), .ZN(n7561) );
  INV_X1 U9173 ( .A(n7561), .ZN(n7562) );
  INV_X1 U9174 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n7564) );
  MUX2_X1 U9175 ( .A(n7570), .B(n7564), .S(n10366), .Z(n7566) );
  NAND2_X1 U9176 ( .A1(n8539), .A2(n9204), .ZN(n7565) );
  OAI211_X1 U9177 ( .C1(n7574), .C2(n9212), .A(n7566), .B(n7565), .ZN(P2_U3441) );
  MUX2_X1 U9178 ( .A(n7570), .B(n7567), .S(n10198), .Z(n7569) );
  AOI22_X1 U9179 ( .A1(n8539), .A2(n8726), .B1(n8709), .B2(n8342), .ZN(n7568)
         );
  OAI211_X1 U9180 ( .C1(n7574), .C2(n8729), .A(n7569), .B(n7568), .ZN(P2_U3216) );
  MUX2_X1 U9181 ( .A(n7571), .B(n7570), .S(n10381), .Z(n7573) );
  NAND2_X1 U9182 ( .A1(n8539), .A2(n8768), .ZN(n7572) );
  OAI211_X1 U9183 ( .C1(n7574), .C2(n8775), .A(n7573), .B(n7572), .ZN(P2_U3476) );
  XOR2_X1 U9184 ( .A(n7576), .B(n7575), .Z(n7586) );
  INV_X1 U9185 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7577) );
  NAND2_X1 U9186 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9275) );
  OAI21_X1 U9187 ( .B1(n9761), .B2(n7577), .A(n9275), .ZN(n7583) );
  INV_X1 U9188 ( .A(n7578), .ZN(n7579) );
  AOI211_X1 U9189 ( .C1(n7581), .C2(n7580), .A(n9752), .B(n7579), .ZN(n7582)
         );
  AOI211_X1 U9190 ( .C1(n9755), .C2(n7584), .A(n7583), .B(n7582), .ZN(n7585)
         );
  OAI21_X1 U9191 ( .B1(n7586), .B2(n9751), .A(n7585), .ZN(P1_U3259) );
  NAND2_X1 U9192 ( .A1(n7588), .A2(n7587), .ZN(n7592) );
  INV_X1 U9193 ( .A(SI_28_), .ZN(n7589) );
  NAND2_X1 U9194 ( .A1(n7590), .A2(n7589), .ZN(n7591) );
  INV_X1 U9195 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7847) );
  INV_X1 U9196 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7597) );
  MUX2_X1 U9197 ( .A(n7847), .B(n7597), .S(n7901), .Z(n7616) );
  XNOR2_X1 U9198 ( .A(n7613), .B(SI_29_), .ZN(n9459) );
  INV_X1 U9199 ( .A(n9459), .ZN(n7596) );
  OAI222_X1 U9200 ( .A1(n7594), .A2(n7596), .B1(n7593), .B2(P2_U3151), .C1(
        n7847), .C2(n9222), .ZN(P2_U3266) );
  OAI222_X1 U9201 ( .A1(n8278), .A2(n7597), .B1(n10173), .B2(n7596), .C1(n7595), .C2(P1_U3086), .ZN(P1_U3326) );
  XNOR2_X1 U9202 ( .A(n10180), .B(n8258), .ZN(n7598) );
  NAND2_X1 U9203 ( .A1(n7598), .A2(n8287), .ZN(n8294) );
  INV_X1 U9204 ( .A(n7598), .ZN(n7599) );
  NAND2_X1 U9205 ( .A1(n7599), .A2(n8420), .ZN(n7600) );
  NAND2_X1 U9206 ( .A1(n8294), .A2(n7600), .ZN(n7605) );
  INV_X1 U9207 ( .A(n8115), .ZN(n7603) );
  AOI21_X1 U9208 ( .B1(n7605), .B2(n7604), .A(n7603), .ZN(n7612) );
  INV_X1 U9209 ( .A(n7606), .ZN(n7608) );
  NOR2_X1 U9210 ( .A1(n8404), .A2(n10191), .ZN(n7607) );
  AOI211_X1 U9211 ( .C1(n8402), .C2(n8419), .A(n7608), .B(n7607), .ZN(n7609)
         );
  OAI21_X1 U9212 ( .B1(n10182), .B2(n8291), .A(n7609), .ZN(n7610) );
  AOI21_X1 U9213 ( .B1(n10180), .B2(n8390), .A(n7610), .ZN(n7611) );
  OAI21_X1 U9214 ( .B1(n7612), .B2(n8394), .A(n7611), .ZN(P2_U3174) );
  INV_X1 U9215 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7626) );
  INV_X1 U9216 ( .A(n7613), .ZN(n7614) );
  NAND2_X1 U9217 ( .A1(n7614), .A2(SI_29_), .ZN(n7620) );
  INV_X1 U9218 ( .A(n7615), .ZN(n7618) );
  INV_X1 U9219 ( .A(n7616), .ZN(n7617) );
  NAND2_X1 U9220 ( .A1(n7618), .A2(n7617), .ZN(n7619) );
  NAND2_X1 U9221 ( .A1(n7620), .A2(n7619), .ZN(n7896) );
  INV_X1 U9222 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9221) );
  MUX2_X1 U9223 ( .A(n9221), .B(n7626), .S(n7901), .Z(n7622) );
  INV_X1 U9224 ( .A(SI_30_), .ZN(n7621) );
  NAND2_X1 U9225 ( .A1(n7622), .A2(n7621), .ZN(n7894) );
  INV_X1 U9226 ( .A(n7622), .ZN(n7623) );
  NAND2_X1 U9227 ( .A1(n7623), .A2(SI_30_), .ZN(n7624) );
  NAND2_X1 U9228 ( .A1(n7894), .A2(n7624), .ZN(n7895) );
  XNOR2_X1 U9229 ( .A(n7896), .B(n7895), .ZN(n9468) );
  INV_X1 U9230 ( .A(n9468), .ZN(n9219) );
  OAI222_X1 U9231 ( .A1(n8278), .A2(n7626), .B1(n10173), .B2(n9219), .C1(
        P1_U3086), .C2(n7625), .ZN(P1_U3325) );
  OAI222_X1 U9232 ( .A1(n8278), .A2(n7628), .B1(n10173), .B2(n7627), .C1(n5176), .C2(P1_U3086), .ZN(P1_U3327) );
  NAND2_X1 U9233 ( .A1(n8085), .A2(n7873), .ZN(n7630) );
  OR2_X1 U9234 ( .A1(n7874), .A2(n8840), .ZN(n7629) );
  NAND2_X1 U9235 ( .A1(n7642), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n7631) );
  NAND2_X1 U9236 ( .A1(n7767), .A2(n7631), .ZN(n8664) );
  NAND2_X1 U9237 ( .A1(n8664), .A2(n7861), .ZN(n7636) );
  INV_X1 U9238 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8832) );
  NAND2_X1 U9239 ( .A1(n7903), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n7633) );
  NAND2_X1 U9240 ( .A1(n7862), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n7632) );
  OAI211_X1 U9241 ( .C1(n7841), .C2(n8832), .A(n7633), .B(n7632), .ZN(n7634)
         );
  INV_X1 U9242 ( .A(n7634), .ZN(n7635) );
  NAND2_X1 U9243 ( .A1(n8246), .A2(n8416), .ZN(n7766) );
  NAND2_X1 U9244 ( .A1(n8072), .A2(n7873), .ZN(n7639) );
  OR2_X1 U9245 ( .A1(n7874), .A2(n7637), .ZN(n7638) );
  OR2_X1 U9246 ( .A1(n7754), .A2(n7640), .ZN(n7641) );
  NAND2_X1 U9247 ( .A1(n7642), .A2(n7641), .ZN(n8684) );
  INV_X1 U9248 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8762) );
  NAND2_X1 U9249 ( .A1(n7903), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n7644) );
  NAND2_X1 U9250 ( .A1(n4814), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n7643) );
  OAI211_X1 U9251 ( .C1(n8762), .C2(n6581), .A(n7644), .B(n7643), .ZN(n7645)
         );
  AOI21_X1 U9252 ( .B1(n8684), .B2(n7861), .A(n7645), .ZN(n8242) );
  OR2_X1 U9253 ( .A1(n9192), .A2(n8242), .ZN(n7953) );
  NAND2_X1 U9254 ( .A1(n7653), .A2(n7646), .ZN(n7647) );
  INV_X1 U9255 ( .A(n7649), .ZN(n7650) );
  OAI21_X1 U9256 ( .B1(n7658), .B2(n7650), .A(n7651), .ZN(n7652) );
  MUX2_X1 U9257 ( .A(n7652), .B(n7651), .S(n7892), .Z(n7660) );
  INV_X1 U9258 ( .A(n7916), .ZN(n7655) );
  INV_X1 U9259 ( .A(n7653), .ZN(n7654) );
  NOR2_X1 U9260 ( .A1(n7655), .A2(n7654), .ZN(n7657) );
  AOI21_X1 U9261 ( .B1(n7658), .B2(n7657), .A(n7656), .ZN(n7659) );
  NAND2_X1 U9262 ( .A1(n7660), .A2(n7659), .ZN(n7669) );
  NAND2_X1 U9263 ( .A1(n7674), .A2(n7893), .ZN(n7664) );
  NAND3_X1 U9264 ( .A1(n7664), .A2(n7661), .A3(n8428), .ZN(n7667) );
  INV_X1 U9265 ( .A(n7662), .ZN(n7665) );
  INV_X1 U9266 ( .A(n7670), .ZN(n7663) );
  OAI22_X1 U9267 ( .A1(n7665), .A2(n7664), .B1(n7663), .B2(n7893), .ZN(n7666)
         );
  AND2_X1 U9268 ( .A1(n7667), .A2(n7666), .ZN(n7668) );
  NAND2_X1 U9269 ( .A1(n7675), .A2(n7670), .ZN(n7672) );
  NAND2_X1 U9270 ( .A1(n7675), .A2(n7674), .ZN(n7678) );
  INV_X1 U9271 ( .A(n7681), .ZN(n7682) );
  NAND2_X1 U9272 ( .A1(n7691), .A2(n7690), .ZN(n7686) );
  NAND2_X1 U9273 ( .A1(n7684), .A2(n7683), .ZN(n7685) );
  MUX2_X1 U9274 ( .A(n7686), .B(n7685), .S(n7892), .Z(n7695) );
  NOR2_X1 U9275 ( .A1(n7695), .A2(n7687), .ZN(n7688) );
  AND2_X1 U9276 ( .A1(n7690), .A2(n7689), .ZN(n7692) );
  OAI211_X1 U9277 ( .C1(n7695), .C2(n7692), .A(n7691), .B(n7701), .ZN(n7697)
         );
  OAI21_X1 U9278 ( .B1(n7695), .B2(n7694), .A(n7693), .ZN(n7696) );
  MUX2_X1 U9279 ( .A(n7697), .B(n7696), .S(n7893), .Z(n7698) );
  INV_X1 U9280 ( .A(n7698), .ZN(n7699) );
  NAND2_X1 U9281 ( .A1(n7700), .A2(n7699), .ZN(n7705) );
  AND2_X1 U9282 ( .A1(n7708), .A2(n7701), .ZN(n7703) );
  INV_X1 U9283 ( .A(n7707), .ZN(n7702) );
  INV_X1 U9284 ( .A(n7930), .ZN(n7704) );
  NAND2_X1 U9285 ( .A1(n7707), .A2(n7706), .ZN(n7709) );
  NOR2_X1 U9286 ( .A1(n10176), .A2(n7893), .ZN(n7711) );
  MUX2_X1 U9287 ( .A(n8420), .B(n10180), .S(n7893), .Z(n7713) );
  NAND2_X1 U9288 ( .A1(n7713), .A2(n7712), .ZN(n7715) );
  AOI21_X1 U9289 ( .B1(n7716), .B2(n7715), .A(n7714), .ZN(n7722) );
  INV_X1 U9290 ( .A(n7717), .ZN(n7720) );
  INV_X1 U9291 ( .A(n7718), .ZN(n7719) );
  MUX2_X1 U9292 ( .A(n7720), .B(n7719), .S(n7892), .Z(n7721) );
  OR3_X1 U9293 ( .A1(n7722), .A2(n7721), .A3(n4699), .ZN(n7723) );
  AOI21_X1 U9294 ( .B1(n7726), .B2(n7724), .A(n7892), .ZN(n7725) );
  NAND2_X1 U9295 ( .A1(n8029), .A2(n7873), .ZN(n7728) );
  AOI22_X1 U9296 ( .A1(n7737), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7736), .B2(
        n8495), .ZN(n7727) );
  NAND2_X1 U9297 ( .A1(n8772), .A2(n8341), .ZN(n7913) );
  OAI211_X1 U9298 ( .C1(n7892), .C2(n7729), .A(n7936), .B(n7913), .ZN(n7735)
         );
  AND2_X1 U9299 ( .A1(n7913), .A2(n7893), .ZN(n7733) );
  NAND2_X1 U9300 ( .A1(n8697), .A2(n7730), .ZN(n7732) );
  NAND2_X1 U9301 ( .A1(n7913), .A2(n7945), .ZN(n7731) );
  AOI22_X1 U9302 ( .A1(n7733), .A2(n7732), .B1(n7731), .B2(n7892), .ZN(n7734)
         );
  NAND2_X1 U9303 ( .A1(n8042), .A2(n7873), .ZN(n7739) );
  AOI22_X1 U9304 ( .A1(n7737), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7981), .B2(
        n7736), .ZN(n7738) );
  AND2_X1 U9305 ( .A1(n7740), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n7741) );
  OR2_X1 U9306 ( .A1(n7741), .A2(n7752), .ZN(n8708) );
  NAND2_X1 U9307 ( .A1(n8708), .A2(n7861), .ZN(n7744) );
  AOI22_X1 U9308 ( .A1(n4814), .A2(P2_REG0_REG_19__SCAN_IN), .B1(n7903), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n7743) );
  INV_X1 U9309 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9081) );
  OR2_X1 U9310 ( .A1(n6581), .A2(n9081), .ZN(n7742) );
  OR2_X1 U9311 ( .A1(n9205), .A2(n8720), .ZN(n7760) );
  AND2_X1 U9312 ( .A1(n7760), .A2(n8697), .ZN(n7948) );
  INV_X1 U9313 ( .A(n7948), .ZN(n7746) );
  NAND2_X1 U9314 ( .A1(n9205), .A2(n8720), .ZN(n7949) );
  INV_X1 U9315 ( .A(n7949), .ZN(n7745) );
  AOI21_X1 U9316 ( .B1(n7746), .B2(n7892), .A(n7745), .ZN(n7747) );
  NAND2_X1 U9317 ( .A1(n8057), .A2(n7873), .ZN(n7750) );
  OR2_X1 U9318 ( .A1(n7874), .A2(n7748), .ZN(n7749) );
  NOR2_X1 U9319 ( .A1(n7752), .A2(n7751), .ZN(n7753) );
  OR2_X1 U9320 ( .A1(n7754), .A2(n7753), .ZN(n8694) );
  NAND2_X1 U9321 ( .A1(n8694), .A2(n7861), .ZN(n7759) );
  INV_X1 U9322 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9197) );
  NAND2_X1 U9323 ( .A1(n7862), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n7756) );
  NAND2_X1 U9324 ( .A1(n7903), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n7755) );
  OAI211_X1 U9325 ( .C1(n7841), .C2(n9197), .A(n7756), .B(n7755), .ZN(n7757)
         );
  INV_X1 U9326 ( .A(n7757), .ZN(n7758) );
  NAND2_X1 U9327 ( .A1(n8547), .A2(n8704), .ZN(n7951) );
  NAND2_X1 U9328 ( .A1(n9198), .A2(n8546), .ZN(n8673) );
  NAND2_X1 U9329 ( .A1(n7951), .A2(n8673), .ZN(n8689) );
  INV_X1 U9330 ( .A(n8689), .ZN(n8545) );
  NAND3_X1 U9331 ( .A1(n7782), .A2(n7760), .A3(n8545), .ZN(n7764) );
  NAND2_X1 U9332 ( .A1(n7953), .A2(n7951), .ZN(n7762) );
  NAND2_X1 U9333 ( .A1(n9192), .A2(n8242), .ZN(n7912) );
  AND2_X1 U9334 ( .A1(n7912), .A2(n8673), .ZN(n7952) );
  INV_X1 U9335 ( .A(n7952), .ZN(n7761) );
  MUX2_X1 U9336 ( .A(n7762), .B(n7761), .S(n7893), .Z(n7781) );
  INV_X1 U9337 ( .A(n7781), .ZN(n7763) );
  NAND2_X1 U9338 ( .A1(n7764), .A2(n7763), .ZN(n7778) );
  NAND2_X1 U9339 ( .A1(n7995), .A2(n7873), .ZN(n7802) );
  OR2_X1 U9340 ( .A1(n7874), .A2(n8788), .ZN(n7801) );
  AND2_X1 U9341 ( .A1(n7801), .A2(n7766), .ZN(n7765) );
  NAND2_X1 U9342 ( .A1(n7802), .A2(n7765), .ZN(n7776) );
  INV_X1 U9343 ( .A(n7766), .ZN(n7774) );
  OR2_X2 U9344 ( .A1(n7767), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n7793) );
  NAND2_X1 U9345 ( .A1(n7767), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n7768) );
  NAND2_X1 U9346 ( .A1(n7793), .A2(n7768), .ZN(n8656) );
  NAND2_X1 U9347 ( .A1(n8656), .A2(n7861), .ZN(n7773) );
  INV_X1 U9348 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8971) );
  NAND2_X1 U9349 ( .A1(n7903), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n7770) );
  INV_X1 U9350 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9184) );
  OR2_X1 U9351 ( .A1(n7841), .A2(n9184), .ZN(n7769) );
  OAI211_X1 U9352 ( .C1(n8971), .C2(n6581), .A(n7770), .B(n7769), .ZN(n7771)
         );
  INV_X1 U9353 ( .A(n7771), .ZN(n7772) );
  OR2_X1 U9354 ( .A1(n7774), .A2(n8549), .ZN(n7775) );
  AND2_X1 U9355 ( .A1(n7776), .A2(n7775), .ZN(n7777) );
  AOI21_X1 U9356 ( .B1(n7779), .B2(n7778), .A(n7777), .ZN(n7780) );
  NAND2_X1 U9357 ( .A1(n7781), .A2(n7912), .ZN(n7784) );
  NAND3_X1 U9358 ( .A1(n7782), .A2(n7952), .A3(n7949), .ZN(n7783) );
  NAND2_X1 U9359 ( .A1(n7784), .A2(n7783), .ZN(n7786) );
  INV_X1 U9360 ( .A(n7955), .ZN(n7785) );
  AOI21_X1 U9361 ( .B1(n7786), .B2(n8668), .A(n7785), .ZN(n7787) );
  INV_X1 U9362 ( .A(n7805), .ZN(n7804) );
  NAND2_X1 U9363 ( .A1(n8149), .A2(n7873), .ZN(n7792) );
  OR2_X1 U9364 ( .A1(n7874), .A2(n7790), .ZN(n7791) );
  INV_X1 U9365 ( .A(n7814), .ZN(n7795) );
  NAND2_X1 U9366 ( .A1(n7793), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n7794) );
  NAND2_X1 U9367 ( .A1(n7795), .A2(n7794), .ZN(n8644) );
  NAND2_X1 U9368 ( .A1(n8644), .A2(n7861), .ZN(n7800) );
  INV_X1 U9369 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8813) );
  NAND2_X1 U9370 ( .A1(n7903), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n7797) );
  NAND2_X1 U9371 ( .A1(n4814), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n7796) );
  OAI211_X1 U9372 ( .C1(n8813), .C2(n6581), .A(n7797), .B(n7796), .ZN(n7798)
         );
  INV_X1 U9373 ( .A(n7798), .ZN(n7799) );
  AND2_X1 U9374 ( .A1(n8614), .A2(n4540), .ZN(n7803) );
  AND2_X1 U9375 ( .A1(n8642), .A2(n8415), .ZN(n8613) );
  AOI21_X1 U9376 ( .B1(n7804), .B2(n7803), .A(n8613), .ZN(n7810) );
  NAND2_X1 U9377 ( .A1(n7805), .A2(n4540), .ZN(n7808) );
  NAND2_X1 U9378 ( .A1(n9185), .A2(n8549), .ZN(n7956) );
  AND2_X1 U9379 ( .A1(n7911), .A2(n7956), .ZN(n7807) );
  INV_X1 U9380 ( .A(n8614), .ZN(n7806) );
  AOI21_X1 U9381 ( .B1(n7808), .B2(n7807), .A(n7806), .ZN(n7809) );
  MUX2_X1 U9382 ( .A(n7810), .B(n7809), .S(n7892), .Z(n7822) );
  NAND2_X1 U9383 ( .A1(n8167), .A2(n7873), .ZN(n7813) );
  OR2_X1 U9384 ( .A1(n7874), .A2(n7811), .ZN(n7812) );
  INV_X1 U9385 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8318) );
  NAND2_X1 U9386 ( .A1(n7814), .A2(n8318), .ZN(n7826) );
  OR2_X1 U9387 ( .A1(n7814), .A2(n8318), .ZN(n7815) );
  NAND2_X1 U9388 ( .A1(n7826), .A2(n7815), .ZN(n8627) );
  NAND2_X1 U9389 ( .A1(n8627), .A2(n7861), .ZN(n7820) );
  INV_X1 U9390 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8749) );
  NAND2_X1 U9391 ( .A1(n7903), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n7817) );
  NAND2_X1 U9392 ( .A1(n4814), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n7816) );
  OAI211_X1 U9393 ( .C1(n8749), .C2(n6581), .A(n7817), .B(n7816), .ZN(n7818)
         );
  INV_X1 U9394 ( .A(n7818), .ZN(n7819) );
  NAND2_X1 U9395 ( .A1(n7820), .A2(n7819), .ZN(n8639) );
  XNOR2_X1 U9396 ( .A(n9173), .B(n8639), .ZN(n8617) );
  INV_X1 U9397 ( .A(n8617), .ZN(n8621) );
  OR2_X1 U9398 ( .A1(n9173), .A2(n8595), .ZN(n7959) );
  NAND2_X1 U9399 ( .A1(n9173), .A2(n8595), .ZN(n7958) );
  MUX2_X1 U9400 ( .A(n7959), .B(n7958), .S(n7893), .Z(n7821) );
  NAND2_X1 U9401 ( .A1(n8183), .A2(n7873), .ZN(n7825) );
  OR2_X1 U9402 ( .A1(n7874), .A2(n7823), .ZN(n7824) );
  NAND2_X1 U9403 ( .A1(n7826), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n7827) );
  NAND2_X1 U9404 ( .A1(n7836), .A2(n7827), .ZN(n8607) );
  NAND2_X1 U9405 ( .A1(n8607), .A2(n7861), .ZN(n7832) );
  INV_X1 U9406 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9168) );
  NAND2_X1 U9407 ( .A1(n7903), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n7829) );
  NAND2_X1 U9408 ( .A1(n7862), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n7828) );
  OAI211_X1 U9409 ( .C1(n9168), .C2(n7841), .A(n7829), .B(n7828), .ZN(n7830)
         );
  INV_X1 U9410 ( .A(n7830), .ZN(n7831) );
  XNOR2_X1 U9411 ( .A(n8557), .B(n8623), .ZN(n8603) );
  NAND2_X1 U9412 ( .A1(n8200), .A2(n7873), .ZN(n7835) );
  OR2_X1 U9413 ( .A1(n7874), .A2(n7833), .ZN(n7834) );
  INV_X1 U9414 ( .A(n7859), .ZN(n7838) );
  NAND2_X1 U9415 ( .A1(n7836), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n7837) );
  NAND2_X1 U9416 ( .A1(n7838), .A2(n7837), .ZN(n8591) );
  NAND2_X1 U9417 ( .A1(n8591), .A2(n7861), .ZN(n7844) );
  INV_X1 U9418 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9162) );
  NAND2_X1 U9419 ( .A1(n7903), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n7840) );
  NAND2_X1 U9420 ( .A1(n7862), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n7839) );
  OAI211_X1 U9421 ( .C1(n9162), .C2(n7841), .A(n7840), .B(n7839), .ZN(n7842)
         );
  INV_X1 U9422 ( .A(n7842), .ZN(n7843) );
  XNOR2_X1 U9423 ( .A(n9163), .B(n8560), .ZN(n8586) );
  NAND2_X1 U9424 ( .A1(n8557), .A2(n8558), .ZN(n7845) );
  OR2_X1 U9425 ( .A1(n8557), .A2(n8558), .ZN(n7963) );
  MUX2_X1 U9426 ( .A(n7845), .B(n7963), .S(n7892), .Z(n7846) );
  NOR2_X1 U9427 ( .A1(n7874), .A2(n7847), .ZN(n7848) );
  INV_X1 U9428 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7858) );
  NAND2_X1 U9429 ( .A1(n8572), .A2(n7861), .ZN(n7905) );
  INV_X1 U9430 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n7851) );
  NAND2_X1 U9431 ( .A1(n7903), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n7850) );
  NAND2_X1 U9432 ( .A1(n4814), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n7849) );
  OAI211_X1 U9433 ( .C1(n6581), .C2(n7851), .A(n7850), .B(n7849), .ZN(n7852)
         );
  INV_X1 U9434 ( .A(n7852), .ZN(n7853) );
  NAND2_X1 U9435 ( .A1(n7905), .A2(n7853), .ZN(n8414) );
  AND2_X1 U9436 ( .A1(n8735), .A2(n8414), .ZN(n7967) );
  INV_X1 U9437 ( .A(n7967), .ZN(n7882) );
  INV_X1 U9438 ( .A(n8735), .ZN(n7854) );
  INV_X1 U9439 ( .A(n8414), .ZN(n8579) );
  NAND2_X1 U9440 ( .A1(n7854), .A2(n8579), .ZN(n7881) );
  NAND2_X1 U9441 ( .A1(n9163), .A2(n8596), .ZN(n7966) );
  INV_X1 U9442 ( .A(n7966), .ZN(n7855) );
  NOR2_X1 U9443 ( .A1(n9163), .A2(n8596), .ZN(n7965) );
  MUX2_X1 U9444 ( .A(n7855), .B(n7965), .S(n7893), .Z(n7856) );
  NOR2_X1 U9445 ( .A1(n7859), .A2(n7858), .ZN(n7860) );
  NAND2_X1 U9446 ( .A1(n8581), .A2(n7861), .ZN(n7868) );
  INV_X1 U9447 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8962) );
  NAND2_X1 U9448 ( .A1(n7862), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n7864) );
  NAND2_X1 U9449 ( .A1(n4814), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7863) );
  OAI211_X1 U9450 ( .C1(n7865), .C2(n8962), .A(n7864), .B(n7863), .ZN(n7866)
         );
  INV_X1 U9451 ( .A(n7866), .ZN(n7867) );
  NAND2_X1 U9452 ( .A1(n8216), .A2(n7873), .ZN(n7871) );
  OR2_X1 U9453 ( .A1(n7874), .A2(n7869), .ZN(n7870) );
  MUX2_X1 U9454 ( .A(n8566), .B(n9157), .S(n7893), .Z(n7888) );
  OR2_X1 U9455 ( .A1(n8562), .A2(n7888), .ZN(n7872) );
  NAND2_X1 U9456 ( .A1(n7889), .A2(n7872), .ZN(n7885) );
  NAND2_X1 U9457 ( .A1(n9468), .A2(n7873), .ZN(n7876) );
  OR2_X1 U9458 ( .A1(n7874), .A2(n9221), .ZN(n7875) );
  NAND2_X1 U9459 ( .A1(n7876), .A2(n7875), .ZN(n7969) );
  INV_X1 U9460 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8868) );
  NAND2_X1 U9461 ( .A1(n4814), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n7878) );
  NAND2_X1 U9462 ( .A1(n7903), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n7877) );
  OAI211_X1 U9463 ( .C1(n8868), .C2(n6581), .A(n7878), .B(n7877), .ZN(n7879)
         );
  INV_X1 U9464 ( .A(n7879), .ZN(n7880) );
  AND2_X1 U9465 ( .A1(n7905), .A2(n7880), .ZN(n8565) );
  NAND2_X1 U9466 ( .A1(n7969), .A2(n8565), .ZN(n7910) );
  NAND2_X1 U9467 ( .A1(n7910), .A2(n7881), .ZN(n7968) );
  AOI21_X1 U9468 ( .B1(n7885), .B2(n8566), .A(n7968), .ZN(n7887) );
  INV_X1 U9469 ( .A(n8565), .ZN(n8413) );
  AND2_X1 U9470 ( .A1(n8781), .A2(n8413), .ZN(n7970) );
  INV_X1 U9471 ( .A(n7970), .ZN(n7883) );
  NAND2_X1 U9472 ( .A1(n7883), .A2(n7882), .ZN(n7884) );
  AOI21_X1 U9473 ( .B1(n7885), .B2(n9157), .A(n7884), .ZN(n7886) );
  OR2_X1 U9474 ( .A1(n7889), .A2(n7888), .ZN(n7890) );
  OAI21_X1 U9475 ( .B1(n7896), .B2(n7895), .A(n7894), .ZN(n7900) );
  INV_X1 U9476 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n7897) );
  MUX2_X1 U9477 ( .A(n5361), .B(n7897), .S(n7901), .Z(n7898) );
  XNOR2_X1 U9478 ( .A(n7898), .B(SI_31_), .ZN(n7899) );
  XNOR2_X1 U9479 ( .A(n7900), .B(n7899), .ZN(n9472) );
  MUX2_X1 U9480 ( .A(n9472), .B(P1_DATAO_REG_31__SCAN_IN), .S(n7901), .Z(n7902) );
  INV_X1 U9481 ( .A(n8778), .ZN(n7971) );
  INV_X1 U9482 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7906) );
  AOI22_X1 U9483 ( .A1(n4814), .A2(P2_REG0_REG_31__SCAN_IN), .B1(n7903), .B2(
        P2_REG2_REG_31__SCAN_IN), .ZN(n7904) );
  OAI211_X1 U9484 ( .C1(n6581), .C2(n7906), .A(n7905), .B(n7904), .ZN(n8412)
         );
  INV_X1 U9485 ( .A(n8412), .ZN(n8532) );
  NAND2_X1 U9486 ( .A1(n7971), .A2(n8532), .ZN(n7975) );
  NAND2_X1 U9487 ( .A1(n8778), .A2(n8412), .ZN(n7972) );
  INV_X1 U9488 ( .A(n7972), .ZN(n7944) );
  NAND2_X1 U9489 ( .A1(n7909), .A2(n7908), .ZN(n7980) );
  INV_X1 U9490 ( .A(n7910), .ZN(n7943) );
  XNOR2_X1 U9491 ( .A(n8582), .B(n8566), .ZN(n8576) );
  NAND2_X1 U9492 ( .A1(n8642), .A2(n8415), .ZN(n7911) );
  NAND2_X1 U9493 ( .A1(n8614), .A2(n7911), .ZN(n8553) );
  INV_X1 U9494 ( .A(n8553), .ZN(n8635) );
  XNOR2_X1 U9495 ( .A(n9205), .B(n8720), .ZN(n8699) );
  NAND2_X1 U9496 ( .A1(n8697), .A2(n7913), .ZN(n8712) );
  NAND4_X1 U9497 ( .A1(n7916), .A2(n7915), .A3(n10295), .A4(n7914), .ZN(n7919)
         );
  NOR3_X1 U9498 ( .A1(n7919), .A2(n7918), .A3(n7917), .ZN(n7923) );
  NAND4_X1 U9499 ( .A1(n7923), .A2(n7922), .A3(n7921), .A4(n7920), .ZN(n7925)
         );
  NOR2_X1 U9500 ( .A1(n7925), .A2(n7924), .ZN(n7926) );
  NAND3_X1 U9501 ( .A1(n7928), .A2(n7927), .A3(n7926), .ZN(n7929) );
  NOR2_X1 U9502 ( .A1(n7930), .A2(n7929), .ZN(n7931) );
  NAND4_X1 U9503 ( .A1(n7932), .A2(n7276), .A3(n7931), .A4(n10189), .ZN(n7933)
         );
  NOR2_X1 U9504 ( .A1(n7934), .A2(n7933), .ZN(n7935) );
  NAND2_X1 U9505 ( .A1(n7936), .A2(n7935), .ZN(n7937) );
  NOR4_X1 U9506 ( .A1(n8689), .A2(n8699), .A3(n8712), .A4(n7937), .ZN(n7938)
         );
  NAND4_X1 U9507 ( .A1(n8652), .A2(n8668), .A3(n8678), .A4(n7938), .ZN(n7939)
         );
  NOR2_X1 U9508 ( .A1(n8553), .A2(n7939), .ZN(n7940) );
  NAND4_X1 U9509 ( .A1(n8586), .A2(n7940), .A3(n8603), .A4(n8617), .ZN(n7941)
         );
  OR3_X1 U9510 ( .A1(n8562), .A2(n8576), .A3(n7941), .ZN(n7942) );
  NOR4_X1 U9511 ( .A1(n7944), .A2(n7970), .A3(n7943), .A4(n7942), .ZN(n7974)
         );
  NAND2_X1 U9512 ( .A1(n8715), .A2(n7948), .ZN(n7950) );
  NAND2_X1 U9513 ( .A1(n7950), .A2(n7949), .ZN(n8687) );
  NAND2_X1 U9514 ( .A1(n8687), .A2(n7951), .ZN(n8674) );
  NAND2_X1 U9515 ( .A1(n8674), .A2(n7952), .ZN(n7954) );
  INV_X1 U9516 ( .A(n7958), .ZN(n7961) );
  OR2_X1 U9517 ( .A1(n7961), .A2(n8613), .ZN(n8600) );
  INV_X1 U9518 ( .A(n8603), .ZN(n7962) );
  AND2_X1 U9519 ( .A1(n8614), .A2(n7959), .ZN(n7960) );
  OR2_X1 U9520 ( .A1(n7962), .A2(n8601), .ZN(n8605) );
  NAND2_X1 U9521 ( .A1(n7976), .A2(n7975), .ZN(n7978) );
  NAND2_X1 U9522 ( .A1(n7978), .A2(n7977), .ZN(n7979) );
  NAND3_X1 U9523 ( .A1(n7984), .A2(n7983), .A3(n8512), .ZN(n7985) );
  OAI211_X1 U9524 ( .C1(n7986), .C2(n7988), .A(n7985), .B(P2_B_REG_SCAN_IN), 
        .ZN(n7987) );
  OAI21_X1 U9525 ( .B1(n7989), .B2(n7988), .A(n7987), .ZN(P2_U3296) );
  OAI222_X1 U9526 ( .A1(n8278), .A2(n7991), .B1(n10173), .B2(n7990), .C1(
        P1_U3086), .C2(n5280), .ZN(P1_U3333) );
  AOI22_X1 U9527 ( .A1(n10171), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n9658), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n7992) );
  OAI21_X1 U9528 ( .B1(n7994), .B2(n10173), .A(n7992), .ZN(P1_U3353) );
  OAI222_X1 U9529 ( .A1(n9222), .A2(n4850), .B1(n9220), .B2(n7994), .C1(
        P2_U3151), .C2(n7993), .ZN(P2_U3293) );
  AND2_X1 U9530 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n7996) );
  NOR2_X1 U9531 ( .A1(n8089), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n7997) );
  OR2_X1 U9532 ( .A1(n8101), .A2(n7997), .ZN(n8108) );
  INV_X1 U9533 ( .A(n8108), .ZN(n9905) );
  NAND2_X1 U9534 ( .A1(n9905), .A2(n5720), .ZN(n8002) );
  INV_X1 U9535 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n8842) );
  NAND2_X1 U9536 ( .A1(n9476), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n7999) );
  NAND2_X1 U9537 ( .A1(n9477), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n7998) );
  OAI211_X1 U9538 ( .C1(n8842), .C2(n8175), .A(n7999), .B(n7998), .ZN(n8000)
         );
  INV_X1 U9539 ( .A(n8000), .ZN(n8001) );
  AOI22_X1 U9540 ( .A1(n10071), .A2(n8208), .B1(n5521), .B2(n9891), .ZN(n8003)
         );
  XNOR2_X1 U9541 ( .A(n8003), .B(n4495), .ZN(n8005) );
  AOI22_X1 U9542 ( .A1(n10071), .A2(n5521), .B1(n8182), .B2(n9891), .ZN(n8004)
         );
  NAND2_X1 U9543 ( .A1(n8005), .A2(n8004), .ZN(n9289) );
  OAI21_X1 U9544 ( .B1(n8005), .B2(n8004), .A(n9289), .ZN(n8161) );
  INV_X1 U9545 ( .A(n8006), .ZN(n8007) );
  AOI22_X1 U9546 ( .A1(n10116), .A2(n8208), .B1(n5521), .B2(n9630), .ZN(n8011)
         );
  OAI22_X1 U9547 ( .A1(n9247), .A2(n8226), .B1(n9361), .B2(n5702), .ZN(n9237)
         );
  INV_X1 U9548 ( .A(n8012), .ZN(n8013) );
  NAND2_X1 U9549 ( .A1(n8013), .A2(n4558), .ZN(n9236) );
  AOI22_X1 U9550 ( .A1(n9418), .A2(n8208), .B1(n5521), .B2(n9629), .ZN(n8014)
         );
  XNOR2_X1 U9551 ( .A(n8014), .B(n4495), .ZN(n9353) );
  AOI22_X1 U9552 ( .A1(n9418), .A2(n5521), .B1(n8182), .B2(n9629), .ZN(n9352)
         );
  NAND2_X1 U9553 ( .A1(n9351), .A2(n9353), .ZN(n8015) );
  NAND2_X1 U9554 ( .A1(n10111), .A2(n8208), .ZN(n8017) );
  OR2_X1 U9555 ( .A1(n10012), .A2(n8226), .ZN(n8016) );
  NAND2_X1 U9556 ( .A1(n8017), .A2(n8016), .ZN(n8018) );
  XNOR2_X1 U9557 ( .A(n8018), .B(n4495), .ZN(n9272) );
  NAND2_X1 U9558 ( .A1(n10111), .A2(n5521), .ZN(n8020) );
  OR2_X1 U9559 ( .A1(n10012), .A2(n5702), .ZN(n8019) );
  NAND2_X1 U9560 ( .A1(n8020), .A2(n8019), .ZN(n9271) );
  NOR2_X1 U9561 ( .A1(n9272), .A2(n9271), .ZN(n8022) );
  NAND2_X1 U9562 ( .A1(n9272), .A2(n9271), .ZN(n8021) );
  NAND2_X1 U9563 ( .A1(n8023), .A2(n9467), .ZN(n8025) );
  AOI22_X1 U9564 ( .A1(n9473), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n8043), .B2(
        n9735), .ZN(n8024) );
  OAI22_X1 U9565 ( .A1(n10165), .A2(n5716), .B1(n9779), .B2(n8226), .ZN(n8026)
         );
  XNOR2_X1 U9566 ( .A(n8026), .B(n4495), .ZN(n8028) );
  OAI22_X1 U9567 ( .A1(n10165), .A2(n8226), .B1(n9779), .B2(n5702), .ZN(n8027)
         );
  AND2_X1 U9568 ( .A1(n8028), .A2(n8027), .ZN(n9281) );
  OR2_X1 U9569 ( .A1(n8028), .A2(n8027), .ZN(n9280) );
  NAND2_X1 U9570 ( .A1(n8029), .A2(n9467), .ZN(n8031) );
  AOI22_X1 U9571 ( .A1(n9473), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n4494), .B2(
        n9738), .ZN(n8030) );
  NAND2_X1 U9572 ( .A1(n9477), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8033) );
  NAND2_X1 U9573 ( .A1(n4491), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n8032) );
  AND2_X1 U9574 ( .A1(n8033), .A2(n8032), .ZN(n8037) );
  INV_X1 U9575 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8034) );
  XNOR2_X1 U9576 ( .A(n8046), .B(n8034), .ZN(n9991) );
  NAND2_X1 U9577 ( .A1(n9991), .A2(n5720), .ZN(n8036) );
  NAND2_X1 U9578 ( .A1(n9476), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8035) );
  AOI22_X1 U9579 ( .A1(n10099), .A2(n8208), .B1(n5521), .B2(n9971), .ZN(n8038)
         );
  XNOR2_X1 U9580 ( .A(n8038), .B(n4495), .ZN(n8040) );
  INV_X1 U9581 ( .A(n8040), .ZN(n8039) );
  AOI22_X1 U9582 ( .A1(n10099), .A2(n5521), .B1(n8182), .B2(n9971), .ZN(n9332)
         );
  NAND2_X1 U9583 ( .A1(n9331), .A2(n9332), .ZN(n8041) );
  NAND2_X1 U9584 ( .A1(n8042), .A2(n9467), .ZN(n8045) );
  AOI22_X1 U9585 ( .A1(n9473), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n8043), .B2(
        n5281), .ZN(n8044) );
  AOI21_X1 U9586 ( .B1(n8046), .B2(P1_REG3_REG_18__SCAN_IN), .A(
        P1_REG3_REG_19__SCAN_IN), .ZN(n8047) );
  OR2_X1 U9587 ( .A1(n8060), .A2(n8047), .ZN(n9981) );
  NAND2_X1 U9588 ( .A1(n4491), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8049) );
  NAND2_X1 U9589 ( .A1(n9477), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n8048) );
  AND2_X1 U9590 ( .A1(n8049), .A2(n8048), .ZN(n8051) );
  NAND2_X1 U9591 ( .A1(n9476), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n8050) );
  OAI211_X1 U9592 ( .C1(n9981), .C2(n8172), .A(n8051), .B(n8050), .ZN(n10000)
         );
  INV_X1 U9593 ( .A(n10000), .ZN(n9956) );
  OAI22_X1 U9594 ( .A1(n10159), .A2(n5716), .B1(n9956), .B2(n8226), .ZN(n8052)
         );
  XNOR2_X1 U9595 ( .A(n8052), .B(n4495), .ZN(n8055) );
  AOI22_X1 U9596 ( .A1(n9977), .A2(n5521), .B1(n8182), .B2(n10000), .ZN(n8053)
         );
  XNOR2_X1 U9597 ( .A(n8055), .B(n8053), .ZN(n9249) );
  INV_X1 U9598 ( .A(n8053), .ZN(n8054) );
  NOR2_X1 U9599 ( .A1(n8055), .A2(n8054), .ZN(n8056) );
  NAND2_X1 U9600 ( .A1(n8057), .A2(n9467), .ZN(n8059) );
  NAND2_X1 U9601 ( .A1(n9473), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8058) );
  OR2_X1 U9602 ( .A1(n8060), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n8061) );
  AND2_X1 U9603 ( .A1(n8075), .A2(n8061), .ZN(n9963) );
  NAND2_X1 U9604 ( .A1(n9963), .A2(n5720), .ZN(n8064) );
  AOI22_X1 U9605 ( .A1(n4492), .A2(P1_REG0_REG_20__SCAN_IN), .B1(n5599), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n8063) );
  NAND2_X1 U9606 ( .A1(n9476), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n8062) );
  OAI22_X1 U9607 ( .A1(n10155), .A2(n5716), .B1(n9941), .B2(n8226), .ZN(n8065)
         );
  XNOR2_X1 U9608 ( .A(n8065), .B(n8194), .ZN(n9300) );
  NOR2_X1 U9609 ( .A1(n9941), .A2(n5702), .ZN(n8066) );
  AOI21_X1 U9610 ( .B1(n9962), .B2(n5521), .A(n8066), .ZN(n8068) );
  NAND2_X1 U9611 ( .A1(n9300), .A2(n8068), .ZN(n8067) );
  NAND2_X1 U9612 ( .A1(n9302), .A2(n8067), .ZN(n8071) );
  INV_X1 U9613 ( .A(n9300), .ZN(n8069) );
  INV_X1 U9614 ( .A(n8068), .ZN(n9299) );
  NAND2_X1 U9615 ( .A1(n8069), .A2(n9299), .ZN(n8070) );
  NAND2_X1 U9616 ( .A1(n8071), .A2(n8070), .ZN(n9254) );
  NAND2_X1 U9617 ( .A1(n8072), .A2(n9467), .ZN(n8074) );
  NAND2_X1 U9618 ( .A1(n9473), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8073) );
  NAND2_X1 U9619 ( .A1(n8075), .A2(n9256), .ZN(n8076) );
  AND2_X1 U9620 ( .A1(n8088), .A2(n8076), .ZN(n9945) );
  NAND2_X1 U9621 ( .A1(n9945), .A2(n5720), .ZN(n8079) );
  AOI22_X1 U9622 ( .A1(n9476), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n9477), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n8078) );
  NAND2_X1 U9623 ( .A1(n4492), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8077) );
  OAI22_X1 U9624 ( .A1(n10151), .A2(n5716), .B1(n9957), .B2(n8226), .ZN(n8080)
         );
  XNOR2_X1 U9625 ( .A(n8080), .B(n4495), .ZN(n8083) );
  INV_X1 U9626 ( .A(n9957), .ZN(n9784) );
  AOI22_X1 U9627 ( .A1(n9944), .A2(n5521), .B1(n8182), .B2(n9784), .ZN(n8081)
         );
  XNOR2_X1 U9628 ( .A(n8083), .B(n8081), .ZN(n9255) );
  INV_X1 U9629 ( .A(n8081), .ZN(n8082) );
  NAND2_X1 U9630 ( .A1(n8083), .A2(n8082), .ZN(n8084) );
  NAND2_X1 U9631 ( .A1(n8085), .A2(n9467), .ZN(n8087) );
  NAND2_X1 U9632 ( .A1(n9473), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8086) );
  AND2_X1 U9633 ( .A1(n8088), .A2(n9313), .ZN(n8090) );
  OR2_X1 U9634 ( .A1(n8090), .A2(n8089), .ZN(n9927) );
  INV_X1 U9635 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n8093) );
  NAND2_X1 U9636 ( .A1(n9476), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8092) );
  NAND2_X1 U9637 ( .A1(n9477), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8091) );
  OAI211_X1 U9638 ( .C1(n8175), .C2(n8093), .A(n8092), .B(n8091), .ZN(n8094)
         );
  INV_X1 U9639 ( .A(n8094), .ZN(n8095) );
  AOI22_X1 U9640 ( .A1(n10079), .A2(n8208), .B1(n5521), .B2(n9914), .ZN(n8096)
         );
  XOR2_X1 U9641 ( .A(n4495), .B(n8096), .Z(n8098) );
  INV_X1 U9642 ( .A(n8098), .ZN(n9310) );
  INV_X1 U9643 ( .A(n10079), .ZN(n9931) );
  OAI22_X1 U9644 ( .A1(n9931), .A2(n8226), .B1(n9940), .B2(n5702), .ZN(n9309)
         );
  AOI21_X1 U9645 ( .B1(n8161), .B2(n8163), .A(n4998), .ZN(n8112) );
  INV_X1 U9646 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8100) );
  OAI22_X1 U9647 ( .A1(n9940), .A2(n9360), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8100), .ZN(n8110) );
  OR2_X1 U9648 ( .A1(n8101), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8102) );
  NAND2_X1 U9649 ( .A1(n8170), .A2(n8102), .ZN(n9897) );
  INV_X1 U9650 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n10143) );
  NAND2_X1 U9651 ( .A1(n9476), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8104) );
  NAND2_X1 U9652 ( .A1(n5599), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8103) );
  OAI211_X1 U9653 ( .C1(n8175), .C2(n10143), .A(n8104), .B(n8103), .ZN(n8105)
         );
  INV_X1 U9654 ( .A(n8105), .ZN(n8106) );
  INV_X1 U9655 ( .A(n9913), .ZN(n9443) );
  OAI22_X1 U9656 ( .A1(n9443), .A2(n9345), .B1(n8108), .B2(n9314), .ZN(n8109)
         );
  AOI211_X1 U9657 ( .C1(n10071), .C2(n9363), .A(n8110), .B(n8109), .ZN(n8111)
         );
  OAI21_X1 U9658 ( .B1(n8112), .B2(n9365), .A(n8111), .ZN(P1_U3216) );
  OAI222_X1 U9659 ( .A1(n8278), .A2(n8114), .B1(n10173), .B2(n8113), .C1(n5175), .C2(P1_U3086), .ZN(P1_U3328) );
  NAND2_X1 U9660 ( .A1(n8115), .A2(n8294), .ZN(n8116) );
  XNOR2_X1 U9661 ( .A(n8299), .B(n8139), .ZN(n8117) );
  XNOR2_X1 U9662 ( .A(n8117), .B(n10193), .ZN(n8293) );
  INV_X1 U9663 ( .A(n8117), .ZN(n8118) );
  NAND2_X1 U9664 ( .A1(n8118), .A2(n10193), .ZN(n8119) );
  XNOR2_X1 U9665 ( .A(n8393), .B(n8258), .ZN(n8133) );
  XNOR2_X1 U9666 ( .A(n8133), .B(n8329), .ZN(n8395) );
  XNOR2_X1 U9667 ( .A(n8772), .B(n8258), .ZN(n8120) );
  NAND2_X1 U9668 ( .A1(n8120), .A2(n8341), .ZN(n8129) );
  INV_X1 U9669 ( .A(n8129), .ZN(n8127) );
  XNOR2_X1 U9670 ( .A(n8120), .B(n8341), .ZN(n8378) );
  INV_X1 U9671 ( .A(n8378), .ZN(n8125) );
  XNOR2_X1 U9672 ( .A(n8539), .B(n8258), .ZN(n8121) );
  NAND2_X1 U9673 ( .A1(n8121), .A2(n8721), .ZN(n8334) );
  INV_X1 U9674 ( .A(n8334), .ZN(n8124) );
  XNOR2_X1 U9675 ( .A(n8331), .B(n8139), .ZN(n8128) );
  NAND2_X1 U9676 ( .A1(n8128), .A2(n8417), .ZN(n8337) );
  INV_X1 U9677 ( .A(n8121), .ZN(n8122) );
  INV_X1 U9678 ( .A(n8721), .ZN(n8538) );
  NAND2_X1 U9679 ( .A1(n8122), .A2(n8538), .ZN(n8335) );
  AND2_X1 U9680 ( .A1(n8337), .A2(n8335), .ZN(n8123) );
  OR2_X1 U9681 ( .A1(n8124), .A2(n8123), .ZN(n8375) );
  AND2_X1 U9682 ( .A1(n8125), .A2(n8375), .ZN(n8126) );
  OR2_X1 U9683 ( .A1(n8127), .A2(n8126), .ZN(n8135) );
  INV_X1 U9684 ( .A(n8135), .ZN(n8131) );
  XNOR2_X1 U9685 ( .A(n8128), .B(n8345), .ZN(n8336) );
  AND2_X1 U9686 ( .A1(n8336), .A2(n8334), .ZN(n8373) );
  AND2_X1 U9687 ( .A1(n8373), .A2(n8129), .ZN(n8130) );
  NOR2_X1 U9688 ( .A1(n8131), .A2(n8130), .ZN(n8137) );
  OR2_X1 U9689 ( .A1(n8395), .A2(n8137), .ZN(n8132) );
  INV_X1 U9690 ( .A(n8133), .ZN(n8134) );
  NAND2_X1 U9691 ( .A1(n8134), .A2(n8418), .ZN(n8324) );
  AND2_X1 U9692 ( .A1(n8324), .A2(n8135), .ZN(n8136) );
  NOR2_X1 U9693 ( .A1(n8137), .A2(n8136), .ZN(n8138) );
  XNOR2_X1 U9694 ( .A(n8547), .B(n8258), .ZN(n8358) );
  XNOR2_X1 U9695 ( .A(n9205), .B(n8139), .ZN(n8310) );
  AOI22_X1 U9696 ( .A1(n8358), .A2(n8704), .B1(n8310), .B2(n8690), .ZN(n8143)
         );
  INV_X1 U9697 ( .A(n8310), .ZN(n8356) );
  AOI21_X1 U9698 ( .B1(n8356), .B2(n8720), .A(n8546), .ZN(n8141) );
  NAND3_X1 U9699 ( .A1(n8356), .A2(n8720), .A3(n8546), .ZN(n8140) );
  OAI21_X1 U9700 ( .B1(n8358), .B2(n8141), .A(n8140), .ZN(n8142) );
  AOI21_X2 U9701 ( .B1(n8309), .B2(n8143), .A(n8142), .ZN(n8245) );
  XNOR2_X1 U9702 ( .A(n9192), .B(n8258), .ZN(n8241) );
  XNOR2_X1 U9703 ( .A(n8241), .B(n8242), .ZN(n8244) );
  XOR2_X1 U9704 ( .A(n8245), .B(n8244), .Z(n8148) );
  AOI22_X1 U9705 ( .A1(n8704), .A2(n8379), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8145) );
  NAND2_X1 U9706 ( .A1(n8684), .A2(n8406), .ZN(n8144) );
  OAI211_X1 U9707 ( .C1(n8416), .C2(n8382), .A(n8145), .B(n8144), .ZN(n8146)
         );
  AOI21_X1 U9708 ( .B1(n9192), .B2(n8390), .A(n8146), .ZN(n8147) );
  OAI21_X1 U9709 ( .B1(n8148), .B2(n8394), .A(n8147), .ZN(P2_U3163) );
  NAND2_X1 U9710 ( .A1(n8149), .A2(n9467), .ZN(n8151) );
  NAND2_X1 U9711 ( .A1(n9473), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8150) );
  NAND2_X1 U9712 ( .A1(n9786), .A2(n8208), .ZN(n8153) );
  NAND2_X1 U9713 ( .A1(n9913), .A2(n5521), .ZN(n8152) );
  NAND2_X1 U9714 ( .A1(n8153), .A2(n8152), .ZN(n8154) );
  XNOR2_X1 U9715 ( .A(n8154), .B(n8194), .ZN(n8156) );
  AND2_X1 U9716 ( .A1(n9913), .A2(n8182), .ZN(n8155) );
  AOI21_X1 U9717 ( .B1(n9786), .B2(n5521), .A(n8155), .ZN(n8157) );
  NAND2_X1 U9718 ( .A1(n8156), .A2(n8157), .ZN(n8165) );
  INV_X1 U9719 ( .A(n8156), .ZN(n8159) );
  INV_X1 U9720 ( .A(n8157), .ZN(n8158) );
  NAND2_X1 U9721 ( .A1(n8159), .A2(n8158), .ZN(n8160) );
  INV_X1 U9722 ( .A(n9290), .ZN(n8164) );
  OR2_X1 U9723 ( .A1(n8161), .A2(n8164), .ZN(n8162) );
  OR2_X1 U9724 ( .A1(n8164), .A2(n9289), .ZN(n9292) );
  AND2_X1 U9725 ( .A1(n8165), .A2(n9292), .ZN(n8166) );
  NAND2_X1 U9726 ( .A1(n8167), .A2(n9467), .ZN(n8169) );
  NAND2_X1 U9727 ( .A1(n9473), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8168) );
  NAND2_X1 U9728 ( .A1(n9877), .A2(n8208), .ZN(n8180) );
  INV_X1 U9729 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9265) );
  NAND2_X1 U9730 ( .A1(n8170), .A2(n9265), .ZN(n8171) );
  INV_X1 U9731 ( .A(n8186), .ZN(n8187) );
  NAND2_X1 U9732 ( .A1(n8171), .A2(n8187), .ZN(n9879) );
  INV_X1 U9733 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10139) );
  NAND2_X1 U9734 ( .A1(n9476), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8174) );
  NAND2_X1 U9735 ( .A1(n9477), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8173) );
  OAI211_X1 U9736 ( .C1(n10139), .C2(n8175), .A(n8174), .B(n8173), .ZN(n8176)
         );
  INV_X1 U9737 ( .A(n8176), .ZN(n8177) );
  NAND2_X1 U9738 ( .A1(n9890), .A2(n5521), .ZN(n8179) );
  NAND2_X1 U9739 ( .A1(n8180), .A2(n8179), .ZN(n8181) );
  XNOR2_X1 U9740 ( .A(n8181), .B(n4495), .ZN(n8199) );
  AOI22_X1 U9741 ( .A1(n9877), .A2(n5521), .B1(n8182), .B2(n9890), .ZN(n8197)
         );
  XNOR2_X1 U9742 ( .A(n8199), .B(n8197), .ZN(n9263) );
  NAND2_X1 U9743 ( .A1(n8183), .A2(n9467), .ZN(n8185) );
  NAND2_X1 U9744 ( .A1(n9473), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8184) );
  NAND2_X1 U9745 ( .A1(n10058), .A2(n8208), .ZN(n8193) );
  INV_X1 U9746 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9344) );
  NAND2_X1 U9747 ( .A1(n8186), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8203) );
  AOI21_X1 U9748 ( .B1(n9344), .B2(n8187), .A(n8219), .ZN(n9862) );
  NAND2_X1 U9749 ( .A1(n5720), .A2(n9862), .ZN(n8191) );
  NAND2_X1 U9750 ( .A1(n9476), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8190) );
  NAND2_X1 U9751 ( .A1(n9477), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8189) );
  NAND2_X1 U9752 ( .A1(n4492), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8188) );
  OR2_X1 U9753 ( .A1(n9842), .A2(n8226), .ZN(n8192) );
  NAND2_X1 U9754 ( .A1(n8193), .A2(n8192), .ZN(n8195) );
  XNOR2_X1 U9755 ( .A(n8195), .B(n8194), .ZN(n8213) );
  NOR2_X1 U9756 ( .A1(n9842), .A2(n5702), .ZN(n8196) );
  AOI21_X1 U9757 ( .B1(n10058), .B2(n5521), .A(n8196), .ZN(n8212) );
  XNOR2_X1 U9758 ( .A(n8213), .B(n8212), .ZN(n9340) );
  INV_X1 U9759 ( .A(n8197), .ZN(n8198) );
  NOR2_X1 U9760 ( .A1(n8199), .A2(n8198), .ZN(n9341) );
  NAND2_X1 U9761 ( .A1(n8200), .A2(n9467), .ZN(n8202) );
  NAND2_X1 U9762 ( .A1(n9473), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8201) );
  XNOR2_X1 U9763 ( .A(P1_REG3_REG_27__SCAN_IN), .B(n8203), .ZN(n9847) );
  NAND2_X1 U9764 ( .A1(n5720), .A2(n9847), .ZN(n8207) );
  NAND2_X1 U9765 ( .A1(n9476), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8206) );
  NAND2_X1 U9766 ( .A1(n4491), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8205) );
  NAND2_X1 U9767 ( .A1(n5599), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8204) );
  INV_X1 U9768 ( .A(n9859), .ZN(n9821) );
  AOI22_X1 U9769 ( .A1(n9846), .A2(n8208), .B1(n5521), .B2(n9821), .ZN(n8209)
         );
  XOR2_X1 U9770 ( .A(n4495), .B(n8209), .Z(n8211) );
  OAI22_X1 U9771 ( .A1(n4863), .A2(n8226), .B1(n9859), .B2(n5702), .ZN(n8210)
         );
  NOR2_X1 U9772 ( .A1(n8211), .A2(n8210), .ZN(n8215) );
  AOI21_X1 U9773 ( .B1(n8211), .B2(n8210), .A(n8215), .ZN(n9227) );
  OR2_X1 U9774 ( .A1(n8213), .A2(n8212), .ZN(n9228) );
  NAND2_X1 U9775 ( .A1(n9226), .A2(n8214), .ZN(n9225) );
  NAND2_X1 U9776 ( .A1(n8216), .A2(n9467), .ZN(n8218) );
  NAND2_X1 U9777 ( .A1(n9473), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8217) );
  NAND3_X1 U9778 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_REG3_REG_27__SCAN_IN), 
        .A3(n8219), .ZN(n8232) );
  INV_X1 U9779 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8231) );
  NAND2_X1 U9780 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n8219), .ZN(n8220) );
  NAND2_X1 U9781 ( .A1(n8231), .A2(n8220), .ZN(n8221) );
  NAND2_X1 U9782 ( .A1(n5720), .A2(n9829), .ZN(n8225) );
  NAND2_X1 U9783 ( .A1(n9476), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8224) );
  NAND2_X1 U9784 ( .A1(n9477), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8223) );
  NAND2_X1 U9785 ( .A1(n4491), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8222) );
  OAI22_X1 U9786 ( .A1(n10133), .A2(n8226), .B1(n9845), .B2(n5702), .ZN(n8229)
         );
  OAI22_X1 U9787 ( .A1(n10133), .A2(n5716), .B1(n9845), .B2(n8226), .ZN(n8227)
         );
  XNOR2_X1 U9788 ( .A(n8227), .B(n4495), .ZN(n8228) );
  XOR2_X1 U9789 ( .A(n8229), .B(n8228), .Z(n8230) );
  OAI22_X1 U9790 ( .A1(n9360), .A2(n9859), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8231), .ZN(n8239) );
  INV_X1 U9791 ( .A(n9829), .ZN(n8237) );
  INV_X1 U9792 ( .A(n8232), .ZN(n9811) );
  NAND2_X1 U9793 ( .A1(n5720), .A2(n9811), .ZN(n8236) );
  NAND2_X1 U9794 ( .A1(n9476), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8235) );
  NAND2_X1 U9795 ( .A1(n4492), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8234) );
  NAND2_X1 U9796 ( .A1(n5599), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8233) );
  NAND4_X1 U9797 ( .A1(n8236), .A2(n8235), .A3(n8234), .A4(n8233), .ZN(n9820)
         );
  INV_X1 U9798 ( .A(n9820), .ZN(n9462) );
  OAI22_X1 U9799 ( .A1(n9314), .A2(n8237), .B1(n9462), .B2(n9345), .ZN(n8238)
         );
  AOI211_X1 U9800 ( .C1(n9367), .C2(n9363), .A(n8239), .B(n8238), .ZN(n8240)
         );
  INV_X1 U9801 ( .A(n8242), .ZN(n8691) );
  XNOR2_X1 U9802 ( .A(n8246), .B(n8258), .ZN(n8247) );
  XOR2_X1 U9803 ( .A(n8416), .B(n8247), .Z(n8367) );
  XNOR2_X1 U9804 ( .A(n8642), .B(n8258), .ZN(n8248) );
  XOR2_X1 U9805 ( .A(n8415), .B(n8248), .Z(n8350) );
  AOI21_X2 U9806 ( .B1(n8349), .B2(n8350), .A(n8249), .ZN(n8316) );
  XNOR2_X1 U9807 ( .A(n9173), .B(n8258), .ZN(n8250) );
  XNOR2_X1 U9808 ( .A(n8250), .B(n8595), .ZN(n8317) );
  INV_X1 U9809 ( .A(n8250), .ZN(n8251) );
  XNOR2_X1 U9810 ( .A(n8557), .B(n8258), .ZN(n8253) );
  XNOR2_X1 U9811 ( .A(n9163), .B(n8258), .ZN(n8255) );
  NOR2_X1 U9812 ( .A1(n8255), .A2(n8596), .ZN(n8256) );
  AOI21_X1 U9813 ( .B1(n8596), .B2(n8255), .A(n8256), .ZN(n8280) );
  INV_X1 U9814 ( .A(n8256), .ZN(n8257) );
  NAND2_X1 U9815 ( .A1(n8279), .A2(n8257), .ZN(n8260) );
  XOR2_X1 U9816 ( .A(n8258), .B(n8576), .Z(n8259) );
  XNOR2_X1 U9817 ( .A(n8260), .B(n8259), .ZN(n8265) );
  NOR2_X1 U9818 ( .A1(n8579), .A2(n8382), .ZN(n8263) );
  AOI22_X1 U9819 ( .A1(n8581), .A2(n8406), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8261) );
  OAI21_X1 U9820 ( .B1(n8596), .B2(n8404), .A(n8261), .ZN(n8262) );
  AOI211_X1 U9821 ( .C1(n8582), .C2(n8390), .A(n8263), .B(n8262), .ZN(n8264)
         );
  OAI21_X1 U9822 ( .B1(n8265), .B2(n8394), .A(n8264), .ZN(P2_U3160) );
  OAI21_X1 U9823 ( .B1(n8268), .B2(n8267), .A(n8266), .ZN(n8269) );
  NAND2_X1 U9824 ( .A1(n8269), .A2(n9342), .ZN(n8275) );
  AOI22_X1 U9825 ( .A1(n9334), .A2(n5739), .B1(n5899), .B2(n9363), .ZN(n8274)
         );
  AND2_X1 U9826 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9681) );
  NOR2_X1 U9827 ( .A1(n9345), .A2(n8270), .ZN(n8271) );
  AOI211_X1 U9828 ( .C1(n9357), .C2(n8272), .A(n9681), .B(n8271), .ZN(n8273)
         );
  OAI211_X1 U9829 ( .C1(n4567), .C2(n8275), .A(n8274), .B(n8273), .ZN(P1_U3230) );
  OAI222_X1 U9830 ( .A1(n8278), .A2(n8277), .B1(n10173), .B2(n8276), .C1(
        P1_U3086), .C2(n9621), .ZN(P1_U3336) );
  INV_X1 U9831 ( .A(n9163), .ZN(n8561) );
  OAI211_X1 U9832 ( .C1(n8281), .C2(n8280), .A(n8279), .B(n8302), .ZN(n8285)
         );
  AOI22_X1 U9833 ( .A1(n8591), .A2(n8406), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8282) );
  OAI21_X1 U9834 ( .B1(n8558), .B2(n8404), .A(n8282), .ZN(n8283) );
  AOI21_X1 U9835 ( .B1(n8588), .B2(n8402), .A(n8283), .ZN(n8284) );
  OAI211_X1 U9836 ( .C1(n8561), .C2(n8410), .A(n8285), .B(n8284), .ZN(P2_U3154) );
  INV_X1 U9837 ( .A(n8286), .ZN(n8289) );
  NOR2_X1 U9838 ( .A1(n8404), .A2(n8287), .ZN(n8288) );
  AOI211_X1 U9839 ( .C1(n8402), .C2(n8418), .A(n8289), .B(n8288), .ZN(n8290)
         );
  OAI21_X1 U9840 ( .B1(n8292), .B2(n8291), .A(n8290), .ZN(n8298) );
  NAND3_X1 U9841 ( .A1(n8115), .A2(n4984), .A3(n8294), .ZN(n8295) );
  AOI21_X1 U9842 ( .B1(n8296), .B2(n8295), .A(n8394), .ZN(n8297) );
  AOI211_X1 U9843 ( .C1(n8299), .C2(n8390), .A(n8298), .B(n8297), .ZN(n8300)
         );
  INV_X1 U9844 ( .A(n8300), .ZN(P2_U3155) );
  XNOR2_X1 U9845 ( .A(n8301), .B(n8662), .ZN(n8303) );
  NAND2_X1 U9846 ( .A1(n8303), .A2(n8302), .ZN(n8308) );
  INV_X1 U9847 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8304) );
  OAI22_X1 U9848 ( .A1(n8416), .A2(n8404), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8304), .ZN(n8306) );
  NOR2_X1 U9849 ( .A1(n8415), .A2(n8382), .ZN(n8305) );
  AOI211_X1 U9850 ( .C1(n8656), .C2(n8406), .A(n8306), .B(n8305), .ZN(n8307)
         );
  OAI211_X1 U9851 ( .C1(n8550), .C2(n8410), .A(n8308), .B(n8307), .ZN(P2_U3156) );
  XNOR2_X1 U9852 ( .A(n8309), .B(n8310), .ZN(n8357) );
  XNOR2_X1 U9853 ( .A(n8357), .B(n8690), .ZN(n8315) );
  NAND2_X1 U9854 ( .A1(n8704), .A2(n8402), .ZN(n8311) );
  NAND2_X1 U9855 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8520) );
  OAI211_X1 U9856 ( .C1(n8341), .C2(n8404), .A(n8311), .B(n8520), .ZN(n8313)
         );
  INV_X1 U9857 ( .A(n9205), .ZN(n8543) );
  NOR2_X1 U9858 ( .A1(n8543), .A2(n8410), .ZN(n8312) );
  AOI211_X1 U9859 ( .C1(n8708), .C2(n8406), .A(n8313), .B(n8312), .ZN(n8314)
         );
  OAI21_X1 U9860 ( .B1(n8315), .B2(n8394), .A(n8314), .ZN(P2_U3159) );
  XOR2_X1 U9861 ( .A(n8317), .B(n8316), .Z(n8323) );
  OAI22_X1 U9862 ( .A1(n8415), .A2(n8404), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8318), .ZN(n8319) );
  AOI21_X1 U9863 ( .B1(n8627), .B2(n8406), .A(n8319), .ZN(n8320) );
  OAI21_X1 U9864 ( .B1(n8558), .B2(n8382), .A(n8320), .ZN(n8321) );
  AOI21_X1 U9865 ( .B1(n9173), .B2(n8390), .A(n8321), .ZN(n8322) );
  OAI21_X1 U9866 ( .B1(n8323), .B2(n8394), .A(n8322), .ZN(P2_U3165) );
  NAND2_X1 U9867 ( .A1(n8397), .A2(n8324), .ZN(n8374) );
  XNOR2_X1 U9868 ( .A(n8374), .B(n8336), .ZN(n8333) );
  AOI21_X1 U9869 ( .B1(n8402), .B2(n8538), .A(n8325), .ZN(n8328) );
  NAND2_X1 U9870 ( .A1(n8406), .A2(n8326), .ZN(n8327) );
  OAI211_X1 U9871 ( .C1(n8329), .C2(n8404), .A(n8328), .B(n8327), .ZN(n8330)
         );
  AOI21_X1 U9872 ( .B1(n8331), .B2(n8390), .A(n8330), .ZN(n8332) );
  OAI21_X1 U9873 ( .B1(n8333), .B2(n8394), .A(n8332), .ZN(P2_U3166) );
  NAND2_X1 U9874 ( .A1(n8335), .A2(n8334), .ZN(n8340) );
  NAND2_X1 U9875 ( .A1(n8374), .A2(n8336), .ZN(n8338) );
  NAND2_X1 U9876 ( .A1(n8338), .A2(n8337), .ZN(n8339) );
  XOR2_X1 U9877 ( .A(n8340), .B(n8339), .Z(n8348) );
  INV_X1 U9878 ( .A(n8341), .ZN(n8702) );
  AND2_X1 U9879 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8466) );
  AOI21_X1 U9880 ( .B1(n8702), .B2(n8402), .A(n8466), .ZN(n8344) );
  NAND2_X1 U9881 ( .A1(n8406), .A2(n8342), .ZN(n8343) );
  OAI211_X1 U9882 ( .C1(n8345), .C2(n8404), .A(n8344), .B(n8343), .ZN(n8346)
         );
  AOI21_X1 U9883 ( .B1(n8539), .B2(n8390), .A(n8346), .ZN(n8347) );
  OAI21_X1 U9884 ( .B1(n8348), .B2(n8394), .A(n8347), .ZN(P2_U3168) );
  XOR2_X1 U9885 ( .A(n8350), .B(n8349), .Z(n8355) );
  AOI22_X1 U9886 ( .A1(n8662), .A2(n8379), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8352) );
  NAND2_X1 U9887 ( .A1(n8644), .A2(n8406), .ZN(n8351) );
  OAI211_X1 U9888 ( .C1(n8595), .C2(n8382), .A(n8352), .B(n8351), .ZN(n8353)
         );
  AOI21_X1 U9889 ( .B1(n8642), .B2(n8390), .A(n8353), .ZN(n8354) );
  OAI21_X1 U9890 ( .B1(n8355), .B2(n8394), .A(n8354), .ZN(P2_U3169) );
  AOI22_X1 U9891 ( .A1(n8357), .A2(n8720), .B1(n8309), .B2(n8356), .ZN(n8360)
         );
  XNOR2_X1 U9892 ( .A(n8358), .B(n8546), .ZN(n8359) );
  XNOR2_X1 U9893 ( .A(n8360), .B(n8359), .ZN(n8365) );
  AOI22_X1 U9894 ( .A1(n8691), .A2(n8402), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8362) );
  NAND2_X1 U9895 ( .A1(n8406), .A2(n8694), .ZN(n8361) );
  OAI211_X1 U9896 ( .C1(n8720), .C2(n8404), .A(n8362), .B(n8361), .ZN(n8363)
         );
  AOI21_X1 U9897 ( .B1(n9198), .B2(n8390), .A(n8363), .ZN(n8364) );
  OAI21_X1 U9898 ( .B1(n8365), .B2(n8394), .A(n8364), .ZN(P2_U3173) );
  XOR2_X1 U9899 ( .A(n8367), .B(n8366), .Z(n8372) );
  AOI22_X1 U9900 ( .A1(n8691), .A2(n8379), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8369) );
  NAND2_X1 U9901 ( .A1(n8664), .A2(n8406), .ZN(n8368) );
  OAI211_X1 U9902 ( .C1(n8549), .C2(n8382), .A(n8369), .B(n8368), .ZN(n8370)
         );
  AOI21_X1 U9903 ( .B1(n8246), .B2(n8390), .A(n8370), .ZN(n8371) );
  OAI21_X1 U9904 ( .B1(n8372), .B2(n8394), .A(n8371), .ZN(P2_U3175) );
  NAND2_X1 U9905 ( .A1(n8374), .A2(n8373), .ZN(n8376) );
  NAND2_X1 U9906 ( .A1(n8376), .A2(n8375), .ZN(n8377) );
  XOR2_X1 U9907 ( .A(n8378), .B(n8377), .Z(n8385) );
  INV_X1 U9908 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9070) );
  NOR2_X1 U9909 ( .A1(n9070), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8488) );
  AOI21_X1 U9910 ( .B1(n8379), .B2(n8538), .A(n8488), .ZN(n8381) );
  NAND2_X1 U9911 ( .A1(n8406), .A2(n8722), .ZN(n8380) );
  OAI211_X1 U9912 ( .C1(n8720), .C2(n8382), .A(n8381), .B(n8380), .ZN(n8383)
         );
  AOI21_X1 U9913 ( .B1(n8772), .B2(n8390), .A(n8383), .ZN(n8384) );
  OAI21_X1 U9914 ( .B1(n8385), .B2(n8394), .A(n8384), .ZN(P2_U3178) );
  XNOR2_X1 U9915 ( .A(n8386), .B(n8623), .ZN(n8392) );
  NAND2_X1 U9916 ( .A1(n8560), .A2(n8402), .ZN(n8388) );
  AOI22_X1 U9917 ( .A1(n8607), .A2(n8406), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8387) );
  OAI211_X1 U9918 ( .C1(n8595), .C2(n8404), .A(n8388), .B(n8387), .ZN(n8389)
         );
  AOI21_X1 U9919 ( .B1(n8557), .B2(n8390), .A(n8389), .ZN(n8391) );
  OAI21_X1 U9920 ( .B1(n8392), .B2(n8394), .A(n8391), .ZN(P2_U3180) );
  INV_X1 U9921 ( .A(n8393), .ZN(n8411) );
  AOI21_X1 U9922 ( .B1(n8396), .B2(n8395), .A(n8394), .ZN(n8398) );
  NAND2_X1 U9923 ( .A1(n8398), .A2(n8397), .ZN(n8409) );
  INV_X1 U9924 ( .A(n8399), .ZN(n8407) );
  INV_X1 U9925 ( .A(n8400), .ZN(n8401) );
  AOI21_X1 U9926 ( .B1(n8402), .B2(n8417), .A(n8401), .ZN(n8403) );
  OAI21_X1 U9927 ( .B1(n10193), .B2(n8404), .A(n8403), .ZN(n8405) );
  AOI21_X1 U9928 ( .B1(n8407), .B2(n8406), .A(n8405), .ZN(n8408) );
  OAI211_X1 U9929 ( .C1(n8411), .C2(n8410), .A(n8409), .B(n8408), .ZN(P2_U3181) );
  MUX2_X1 U9930 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8412), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U9931 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8413), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9932 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8414), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U9933 ( .A(n8588), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8485), .Z(
        P2_U3519) );
  MUX2_X1 U9934 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8560), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9935 ( .A(n8623), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8485), .Z(
        P2_U3517) );
  MUX2_X1 U9936 ( .A(n8639), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8485), .Z(
        P2_U3516) );
  MUX2_X1 U9937 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8653), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9938 ( .A(n8662), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8485), .Z(
        P2_U3514) );
  MUX2_X1 U9939 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8681), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9940 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8691), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9941 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8704), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9942 ( .A(n8690), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8485), .Z(
        P2_U3510) );
  MUX2_X1 U9943 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8702), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U9944 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8538), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9945 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8417), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9946 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8418), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U9947 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8419), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U9948 ( .A(n8420), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8485), .Z(
        P2_U3504) );
  MUX2_X1 U9949 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8421), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U9950 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8422), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U9951 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8423), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U9952 ( .A(n8424), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8485), .Z(
        P2_U3497) );
  MUX2_X1 U9953 ( .A(n8425), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8485), .Z(
        P2_U3496) );
  MUX2_X1 U9954 ( .A(n8426), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8485), .Z(
        P2_U3495) );
  MUX2_X1 U9955 ( .A(n8427), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8485), .Z(
        P2_U3494) );
  MUX2_X1 U9956 ( .A(n8428), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8485), .Z(
        P2_U3493) );
  MUX2_X1 U9957 ( .A(n8429), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8485), .Z(
        P2_U3492) );
  MUX2_X1 U9958 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8430), .S(P2_U3893), .Z(
        P2_U3491) );
  INV_X1 U9959 ( .A(n8431), .ZN(n8434) );
  OAI21_X1 U9960 ( .B1(n8434), .B2(n8433), .A(n8432), .ZN(n8436) );
  NAND3_X1 U9961 ( .A1(n8436), .A2(n8464), .A3(n8435), .ZN(n8452) );
  OAI21_X1 U9962 ( .B1(n8439), .B2(n8438), .A(n8437), .ZN(n8441) );
  AOI21_X1 U9963 ( .B1(n8442), .B2(n8441), .A(n8440), .ZN(n8451) );
  OAI21_X1 U9964 ( .B1(n8445), .B2(n8444), .A(n8443), .ZN(n8446) );
  AOI22_X1 U9965 ( .A1(n8519), .A2(P2_ADDR_REG_4__SCAN_IN), .B1(n8526), .B2(
        n8446), .ZN(n8450) );
  NAND2_X1 U9966 ( .A1(n8448), .A2(n8447), .ZN(n8449) );
  NAND4_X1 U9967 ( .A1(n8452), .A2(n8451), .A3(n8450), .A4(n8449), .ZN(
        P2_U3186) );
  OAI21_X1 U9968 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8454), .A(n8474), .ZN(
        n8455) );
  INV_X1 U9969 ( .A(n8455), .ZN(n8472) );
  OAI21_X1 U9970 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n8459), .A(n8498), .ZN(
        n8470) );
  NAND2_X1 U9971 ( .A1(n8461), .A2(n8460), .ZN(n8463) );
  MUX2_X1 U9972 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n8512), .Z(n8476) );
  XNOR2_X1 U9973 ( .A(n8476), .B(n8477), .ZN(n8462) );
  NAND2_X1 U9974 ( .A1(n8463), .A2(n8462), .ZN(n8480) );
  OAI21_X1 U9975 ( .B1(n8463), .B2(n8462), .A(n8480), .ZN(n8465) );
  NAND2_X1 U9976 ( .A1(n8465), .A2(n8464), .ZN(n8468) );
  AOI21_X1 U9977 ( .B1(n8519), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8466), .ZN(
        n8467) );
  OAI211_X1 U9978 ( .C1(n8522), .C2(n8493), .A(n8468), .B(n8467), .ZN(n8469)
         );
  AOI21_X1 U9979 ( .B1(n8470), .B2(n8526), .A(n8469), .ZN(n8471) );
  OAI21_X1 U9980 ( .B1(n8472), .B2(n8529), .A(n8471), .ZN(P2_U3199) );
  XNOR2_X1 U9981 ( .A(n8495), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8503) );
  NAND2_X1 U9982 ( .A1(n8493), .A2(n8473), .ZN(n8475) );
  XOR2_X1 U9983 ( .A(n8503), .B(n8504), .Z(n8502) );
  INV_X1 U9984 ( .A(n8476), .ZN(n8478) );
  NAND2_X1 U9985 ( .A1(n8478), .A2(n8477), .ZN(n8479) );
  AND2_X1 U9986 ( .A1(n8480), .A2(n8479), .ZN(n8481) );
  MUX2_X1 U9987 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8512), .Z(n8482) );
  NAND2_X1 U9988 ( .A1(n8481), .A2(n8482), .ZN(n8487) );
  NAND2_X1 U9989 ( .A1(n8487), .A2(n8495), .ZN(n8511) );
  INV_X1 U9990 ( .A(n8481), .ZN(n8484) );
  INV_X1 U9991 ( .A(n8482), .ZN(n8483) );
  NAND2_X1 U9992 ( .A1(n8484), .A2(n8483), .ZN(n8510) );
  INV_X1 U9993 ( .A(n8510), .ZN(n8486) );
  NOR3_X1 U9994 ( .A1(n8511), .A2(n8486), .A3(n8485), .ZN(n8492) );
  AOI211_X1 U9995 ( .C1(n8487), .C2(n8510), .A(n8495), .B(n8517), .ZN(n8491)
         );
  AOI21_X1 U9996 ( .B1(n8519), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8488), .ZN(
        n8489) );
  OAI21_X1 U9997 ( .B1(n8508), .B2(n8522), .A(n8489), .ZN(n8490) );
  NOR3_X1 U9998 ( .A1(n8492), .A2(n8491), .A3(n8490), .ZN(n8501) );
  NAND2_X1 U9999 ( .A1(n8494), .A2(n8493), .ZN(n8496) );
  XNOR2_X1 U10000 ( .A(n8495), .B(n8876), .ZN(n8497) );
  AND3_X1 U10001 ( .A1(n8498), .A2(n8497), .A3(n8496), .ZN(n8499) );
  OAI21_X1 U10002 ( .B1(n8507), .B2(n8499), .A(n8526), .ZN(n8500) );
  OAI211_X1 U10003 ( .C1(n8502), .C2(n8529), .A(n8501), .B(n8500), .ZN(
        P2_U3200) );
  AOI22_X1 U10004 ( .A1(n8504), .A2(n8503), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n8508), .ZN(n8506) );
  XNOR2_X1 U10005 ( .A(n8523), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8513) );
  INV_X1 U10006 ( .A(n8513), .ZN(n8505) );
  XNOR2_X1 U10007 ( .A(n8506), .B(n8505), .ZN(n8530) );
  AOI21_X1 U10008 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n8508), .A(n8507), .ZN(
        n8509) );
  XNOR2_X1 U10009 ( .A(n8523), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8514) );
  XNOR2_X1 U10010 ( .A(n8509), .B(n8514), .ZN(n8527) );
  NAND2_X1 U10011 ( .A1(n8511), .A2(n8510), .ZN(n8516) );
  MUX2_X1 U10012 ( .A(n8514), .B(n8513), .S(n8512), .Z(n8515) );
  XNOR2_X1 U10013 ( .A(n8516), .B(n8515), .ZN(n8518) );
  NOR2_X1 U10014 ( .A1(n8518), .A2(n8517), .ZN(n8525) );
  NAND2_X1 U10015 ( .A1(n8519), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8521) );
  OAI211_X1 U10016 ( .C1(n8523), .C2(n8522), .A(n8521), .B(n8520), .ZN(n8524)
         );
  AOI211_X1 U10017 ( .C1(n8527), .C2(n8526), .A(n8525), .B(n8524), .ZN(n8528)
         );
  OAI21_X1 U10018 ( .B1(n8530), .B2(n8529), .A(n8528), .ZN(P2_U3201) );
  NAND2_X1 U10019 ( .A1(n8709), .A2(n8572), .ZN(n8533) );
  NAND2_X1 U10020 ( .A1(n8703), .A2(n8531), .ZN(n8564) );
  AOI21_X1 U10021 ( .B1(n8533), .B2(n8776), .A(n10198), .ZN(n8535) );
  AOI21_X1 U10022 ( .B1(n10198), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8535), .ZN(
        n8534) );
  OAI21_X1 U10023 ( .B1(n8778), .B2(n8610), .A(n8534), .ZN(P2_U3202) );
  AOI21_X1 U10024 ( .B1(n10198), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8535), .ZN(
        n8536) );
  OAI21_X1 U10025 ( .B1(n8781), .B2(n8610), .A(n8536), .ZN(P2_U3203) );
  NAND2_X1 U10026 ( .A1(n8539), .A2(n8538), .ZN(n8540) );
  NAND2_X1 U10027 ( .A1(n8541), .A2(n8540), .ZN(n8718) );
  OR2_X1 U10028 ( .A1(n8772), .A2(n8702), .ZN(n8542) );
  NOR2_X1 U10029 ( .A1(n9205), .A2(n8690), .ZN(n8544) );
  NAND2_X1 U10030 ( .A1(n8547), .A2(n8546), .ZN(n8677) );
  NAND2_X1 U10031 ( .A1(n8688), .A2(n8677), .ZN(n8548) );
  OR2_X1 U10032 ( .A1(n9192), .A2(n8691), .ZN(n8659) );
  OR2_X1 U10033 ( .A1(n8246), .A2(n8681), .ZN(n8650) );
  NAND2_X1 U10034 ( .A1(n8550), .A2(n8549), .ZN(n8551) );
  NAND2_X1 U10035 ( .A1(n8650), .A2(n8551), .ZN(n8552) );
  NAND2_X1 U10036 ( .A1(n4510), .A2(n8552), .ZN(n8633) );
  AND2_X1 U10037 ( .A1(n8659), .A2(n4545), .ZN(n8554) );
  NAND2_X1 U10038 ( .A1(n8680), .A2(n8554), .ZN(n8631) );
  NAND2_X1 U10039 ( .A1(n8642), .A2(n8653), .ZN(n8555) );
  INV_X1 U10040 ( .A(n8668), .ZN(n8648) );
  AND2_X1 U10041 ( .A1(n4510), .A2(n8648), .ZN(n8632) );
  OR2_X1 U10042 ( .A1(n9173), .A2(n8639), .ZN(n8556) );
  NOR2_X1 U10043 ( .A1(n8557), .A2(n8623), .ZN(n8559) );
  OAI22_X2 U10044 ( .A1(n8594), .A2(n8559), .B1(n8558), .B2(n9170), .ZN(n8587)
         );
  OAI22_X1 U10045 ( .A1(n8566), .A2(n10192), .B1(n8565), .B2(n8564), .ZN(n8567) );
  OAI21_X1 U10046 ( .B1(n8733), .B2(n8570), .A(n8737), .ZN(n8571) );
  NAND2_X1 U10047 ( .A1(n8571), .A2(n8724), .ZN(n8574) );
  AOI22_X1 U10048 ( .A1(n8572), .A2(n8709), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n10198), .ZN(n8573) );
  OAI211_X1 U10049 ( .C1(n8735), .C2(n8610), .A(n8574), .B(n8573), .ZN(
        P2_U3204) );
  XNOR2_X1 U10050 ( .A(n8575), .B(n8576), .ZN(n9158) );
  XNOR2_X1 U10051 ( .A(n8577), .B(n8576), .ZN(n8578) );
  OAI222_X1 U10052 ( .A1(n10192), .A2(n8596), .B1(n10194), .B2(n8579), .C1(
        n8578), .C2(n10296), .ZN(n9156) );
  INV_X1 U10053 ( .A(n9156), .ZN(n8580) );
  MUX2_X1 U10054 ( .A(n8962), .B(n8580), .S(n8724), .Z(n8584) );
  AOI22_X1 U10055 ( .A1(n8582), .A2(n8726), .B1(n8709), .B2(n8581), .ZN(n8583)
         );
  OAI211_X1 U10056 ( .C1(n9158), .C2(n8729), .A(n8584), .B(n8583), .ZN(
        P2_U3205) );
  XNOR2_X1 U10057 ( .A(n8585), .B(n8586), .ZN(n9166) );
  INV_X1 U10058 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8590) );
  XNOR2_X1 U10059 ( .A(n8587), .B(n8586), .ZN(n8589) );
  AOI222_X1 U10060 ( .A1(n8706), .A2(n8589), .B1(n8588), .B2(n8703), .C1(n8623), .C2(n8701), .ZN(n9161) );
  MUX2_X1 U10061 ( .A(n8590), .B(n9161), .S(n8724), .Z(n8593) );
  AOI22_X1 U10062 ( .A1(n9163), .A2(n8726), .B1(n8709), .B2(n8591), .ZN(n8592)
         );
  OAI211_X1 U10063 ( .C1(n9166), .C2(n8729), .A(n8593), .B(n8592), .ZN(
        P2_U3206) );
  XNOR2_X1 U10064 ( .A(n8594), .B(n7962), .ZN(n8598) );
  OAI22_X1 U10065 ( .A1(n8596), .A2(n10194), .B1(n8595), .B2(n10192), .ZN(
        n8597) );
  AOI21_X1 U10066 ( .B1(n8598), .B2(n8706), .A(n8597), .ZN(n8746) );
  NOR2_X1 U10067 ( .A1(n8746), .A2(n10198), .ZN(n8612) );
  OR2_X1 U10068 ( .A1(n8599), .A2(n8600), .ZN(n8602) );
  NAND2_X1 U10069 ( .A1(n8602), .A2(n8601), .ZN(n8604) );
  OR2_X1 U10070 ( .A1(n8604), .A2(n8603), .ZN(n8744) );
  AND2_X1 U10071 ( .A1(n8606), .A2(n8605), .ZN(n8743) );
  NAND3_X1 U10072 ( .A1(n8744), .A2(n8743), .A3(n8670), .ZN(n8609) );
  AOI22_X1 U10073 ( .A1(n8607), .A2(n8709), .B1(n10198), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8608) );
  OAI211_X1 U10074 ( .C1(n9170), .C2(n8610), .A(n8609), .B(n8608), .ZN(n8611)
         );
  OR2_X1 U10075 ( .A1(n8612), .A2(n8611), .ZN(P2_U3207) );
  OR2_X1 U10076 ( .A1(n8599), .A2(n8613), .ZN(n8615) );
  NAND2_X1 U10077 ( .A1(n8615), .A2(n8614), .ZN(n8618) );
  NAND2_X1 U10078 ( .A1(n8618), .A2(n8617), .ZN(n8616) );
  OAI21_X1 U10079 ( .B1(n8618), .B2(n8617), .A(n8616), .ZN(n9176) );
  INV_X1 U10080 ( .A(n9173), .ZN(n8625) );
  AND2_X1 U10081 ( .A1(n8631), .A2(n8619), .ZN(n8622) );
  OAI21_X1 U10082 ( .B1(n8622), .B2(n8621), .A(n8620), .ZN(n8624) );
  AOI222_X1 U10083 ( .A1(n8706), .A2(n8624), .B1(n8623), .B2(n8703), .C1(n8653), .C2(n8701), .ZN(n9171) );
  OAI21_X1 U10084 ( .B1(n8625), .B2(n10183), .A(n9171), .ZN(n8626) );
  NAND2_X1 U10085 ( .A1(n8626), .A2(n8724), .ZN(n8629) );
  AOI22_X1 U10086 ( .A1(n8627), .A2(n8709), .B1(n10198), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n8628) );
  OAI211_X1 U10087 ( .C1(n9176), .C2(n8729), .A(n8629), .B(n8628), .ZN(
        P2_U3208) );
  XNOR2_X1 U10088 ( .A(n8599), .B(n8553), .ZN(n9180) );
  AND2_X1 U10089 ( .A1(n8631), .A2(n8630), .ZN(n8638) );
  NAND2_X1 U10090 ( .A1(n8680), .A2(n8659), .ZN(n8649) );
  NAND2_X1 U10091 ( .A1(n8649), .A2(n8632), .ZN(n8634) );
  NAND2_X1 U10092 ( .A1(n8634), .A2(n8633), .ZN(n8636) );
  NAND2_X1 U10093 ( .A1(n8636), .A2(n8635), .ZN(n8637) );
  NAND3_X1 U10094 ( .A1(n8638), .A2(n8706), .A3(n8637), .ZN(n8641) );
  AOI22_X1 U10095 ( .A1(n8639), .A2(n8703), .B1(n8701), .B2(n8662), .ZN(n8640)
         );
  NAND2_X1 U10096 ( .A1(n8641), .A2(n8640), .ZN(n9177) );
  INV_X1 U10097 ( .A(n8642), .ZN(n9179) );
  NOR2_X1 U10098 ( .A1(n9179), .A2(n10183), .ZN(n8643) );
  OAI21_X1 U10099 ( .B1(n9177), .B2(n8643), .A(n8724), .ZN(n8646) );
  AOI22_X1 U10100 ( .A1(n8644), .A2(n8709), .B1(n10198), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n8645) );
  OAI211_X1 U10101 ( .C1(n9180), .C2(n8729), .A(n8646), .B(n8645), .ZN(
        P2_U3209) );
  XNOR2_X1 U10102 ( .A(n8647), .B(n8652), .ZN(n9188) );
  INV_X1 U10103 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8655) );
  NAND2_X1 U10104 ( .A1(n8649), .A2(n8648), .ZN(n8661) );
  NAND2_X1 U10105 ( .A1(n8661), .A2(n8650), .ZN(n8651) );
  XOR2_X1 U10106 ( .A(n8652), .B(n8651), .Z(n8654) );
  AOI222_X1 U10107 ( .A1(n8706), .A2(n8654), .B1(n8653), .B2(n8703), .C1(n8681), .C2(n8701), .ZN(n9183) );
  MUX2_X1 U10108 ( .A(n8655), .B(n9183), .S(n8724), .Z(n8658) );
  AOI22_X1 U10109 ( .A1(n9185), .A2(n8726), .B1(n8709), .B2(n8656), .ZN(n8657)
         );
  OAI211_X1 U10110 ( .C1(n9188), .C2(n8729), .A(n8658), .B(n8657), .ZN(
        P2_U3210) );
  NAND3_X1 U10111 ( .A1(n8680), .A2(n8668), .A3(n8659), .ZN(n8660) );
  NAND2_X1 U10112 ( .A1(n8661), .A2(n8660), .ZN(n8663) );
  AOI222_X1 U10113 ( .A1(n8706), .A2(n8663), .B1(n8691), .B2(n8701), .C1(n8662), .C2(n8703), .ZN(n8760) );
  INV_X1 U10114 ( .A(n8664), .ZN(n8666) );
  INV_X1 U10115 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8665) );
  OAI22_X1 U10116 ( .A1(n8666), .A2(n10181), .B1(n8724), .B2(n8665), .ZN(n8667) );
  AOI21_X1 U10117 ( .B1(n8246), .B2(n8726), .A(n8667), .ZN(n8672) );
  OR2_X1 U10118 ( .A1(n8669), .A2(n8668), .ZN(n8758) );
  NAND3_X1 U10119 ( .A1(n8758), .A2(n8757), .A3(n8670), .ZN(n8671) );
  OAI211_X1 U10120 ( .C1(n8760), .C2(n10198), .A(n8672), .B(n8671), .ZN(
        P2_U3211) );
  NAND2_X1 U10121 ( .A1(n8674), .A2(n8673), .ZN(n8676) );
  XNOR2_X1 U10122 ( .A(n8676), .B(n8675), .ZN(n9195) );
  INV_X1 U10123 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8683) );
  NAND3_X1 U10124 ( .A1(n8688), .A2(n8678), .A3(n8677), .ZN(n8679) );
  NAND2_X1 U10125 ( .A1(n8680), .A2(n8679), .ZN(n8682) );
  AOI222_X1 U10126 ( .A1(n8706), .A2(n8682), .B1(n8704), .B2(n8701), .C1(n8681), .C2(n8703), .ZN(n9190) );
  MUX2_X1 U10127 ( .A(n8683), .B(n9190), .S(n8724), .Z(n8686) );
  AOI22_X1 U10128 ( .A1(n9192), .A2(n8726), .B1(n8709), .B2(n8684), .ZN(n8685)
         );
  OAI211_X1 U10129 ( .C1(n9195), .C2(n8729), .A(n8686), .B(n8685), .ZN(
        P2_U3212) );
  XNOR2_X1 U10130 ( .A(n8687), .B(n8689), .ZN(n9201) );
  INV_X1 U10131 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8693) );
  OAI21_X1 U10132 ( .B1(n4559), .B2(n8689), .A(n8688), .ZN(n8692) );
  AOI222_X1 U10133 ( .A1(n8706), .A2(n8692), .B1(n8691), .B2(n8703), .C1(n8690), .C2(n8701), .ZN(n9196) );
  MUX2_X1 U10134 ( .A(n8693), .B(n9196), .S(n8724), .Z(n8696) );
  AOI22_X1 U10135 ( .A1(n9198), .A2(n8726), .B1(n8709), .B2(n8694), .ZN(n8695)
         );
  OAI211_X1 U10136 ( .C1(n9201), .C2(n8729), .A(n8696), .B(n8695), .ZN(
        P2_U3213) );
  NAND2_X1 U10137 ( .A1(n8715), .A2(n8697), .ZN(n8698) );
  XOR2_X1 U10138 ( .A(n8699), .B(n8698), .Z(n9208) );
  INV_X1 U10139 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8707) );
  XNOR2_X1 U10140 ( .A(n8700), .B(n8699), .ZN(n8705) );
  AOI222_X1 U10141 ( .A1(n8706), .A2(n8705), .B1(n8704), .B2(n8703), .C1(n8702), .C2(n8701), .ZN(n9202) );
  MUX2_X1 U10142 ( .A(n8707), .B(n9202), .S(n8724), .Z(n8711) );
  AOI22_X1 U10143 ( .A1(n9205), .A2(n8726), .B1(n8709), .B2(n8708), .ZN(n8710)
         );
  OAI211_X1 U10144 ( .C1(n9208), .C2(n8729), .A(n8711), .B(n8710), .ZN(
        P2_U3214) );
  NAND2_X1 U10145 ( .A1(n8713), .A2(n8712), .ZN(n8714) );
  NAND2_X1 U10146 ( .A1(n8715), .A2(n8714), .ZN(n9213) );
  INV_X1 U10147 ( .A(n8716), .ZN(n8717) );
  AOI21_X1 U10148 ( .B1(n7947), .B2(n8718), .A(n8717), .ZN(n8719) );
  OAI222_X1 U10149 ( .A1(n10192), .A2(n8721), .B1(n10194), .B2(n8720), .C1(
        n10296), .C2(n8719), .ZN(n8771) );
  NAND2_X1 U10150 ( .A1(n8771), .A2(n8724), .ZN(n8728) );
  INV_X1 U10151 ( .A(n8722), .ZN(n8723) );
  OAI22_X1 U10152 ( .A1(n8724), .A2(n8876), .B1(n8723), .B2(n10181), .ZN(n8725) );
  AOI21_X1 U10153 ( .B1(n8772), .B2(n8726), .A(n8725), .ZN(n8727) );
  OAI211_X1 U10154 ( .C1(n9213), .C2(n8729), .A(n8728), .B(n8727), .ZN(
        P2_U3215) );
  NOR2_X1 U10155 ( .A1(n8776), .A2(n10378), .ZN(n8731) );
  AOI21_X1 U10156 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n10378), .A(n8731), .ZN(
        n8730) );
  OAI21_X1 U10157 ( .B1(n8778), .B2(n8752), .A(n8730), .ZN(P2_U3490) );
  AOI21_X1 U10158 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n10378), .A(n8731), .ZN(
        n8732) );
  OAI21_X1 U10159 ( .B1(n8781), .B2(n8752), .A(n8732), .ZN(P2_U3489) );
  INV_X1 U10160 ( .A(n8733), .ZN(n8734) );
  NAND2_X1 U10161 ( .A1(n8734), .A2(n10318), .ZN(n8736) );
  MUX2_X1 U10162 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8782), .S(n10381), .Z(
        P2_U3488) );
  MUX2_X1 U10163 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9156), .S(n10381), .Z(
        n8739) );
  OAI22_X1 U10164 ( .A1(n9158), .A2(n8775), .B1(n9157), .B2(n8752), .ZN(n8738)
         );
  OR2_X1 U10165 ( .A1(n8739), .A2(n8738), .ZN(P2_U3487) );
  INV_X1 U10166 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8740) );
  MUX2_X1 U10167 ( .A(n8740), .B(n9161), .S(n10381), .Z(n8742) );
  NAND2_X1 U10168 ( .A1(n9163), .A2(n8768), .ZN(n8741) );
  OAI211_X1 U10169 ( .C1(n8775), .C2(n9166), .A(n8742), .B(n8741), .ZN(
        P2_U3486) );
  INV_X1 U10170 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8747) );
  NAND3_X1 U10171 ( .A1(n8744), .A2(n8743), .A3(n10358), .ZN(n8745) );
  AND2_X1 U10172 ( .A1(n8746), .A2(n8745), .ZN(n9167) );
  MUX2_X1 U10173 ( .A(n8747), .B(n9167), .S(n10381), .Z(n8748) );
  OAI21_X1 U10174 ( .B1(n9170), .B2(n8752), .A(n8748), .ZN(P2_U3485) );
  MUX2_X1 U10175 ( .A(n8749), .B(n9171), .S(n10381), .Z(n8751) );
  NAND2_X1 U10176 ( .A1(n9173), .A2(n8768), .ZN(n8750) );
  OAI211_X1 U10177 ( .C1(n8775), .C2(n9176), .A(n8751), .B(n8750), .ZN(
        P2_U3484) );
  MUX2_X1 U10178 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9177), .S(n10381), .Z(
        n8754) );
  OAI22_X1 U10179 ( .A1(n9180), .A2(n8775), .B1(n9179), .B2(n8752), .ZN(n8753)
         );
  OR2_X1 U10180 ( .A1(n8754), .A2(n8753), .ZN(P2_U3483) );
  MUX2_X1 U10181 ( .A(n8971), .B(n9183), .S(n10381), .Z(n8756) );
  NAND2_X1 U10182 ( .A1(n9185), .A2(n8768), .ZN(n8755) );
  OAI211_X1 U10183 ( .C1(n9188), .C2(n8775), .A(n8756), .B(n8755), .ZN(
        P2_U3482) );
  INV_X1 U10184 ( .A(n8246), .ZN(n8761) );
  NAND3_X1 U10185 ( .A1(n8758), .A2(n8757), .A3(n10358), .ZN(n8759) );
  OAI211_X1 U10186 ( .C1(n8761), .C2(n10352), .A(n8760), .B(n8759), .ZN(n9189)
         );
  MUX2_X1 U10187 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9189), .S(n10381), .Z(
        P2_U3481) );
  MUX2_X1 U10188 ( .A(n8762), .B(n9190), .S(n10381), .Z(n8764) );
  NAND2_X1 U10189 ( .A1(n9192), .A2(n8768), .ZN(n8763) );
  OAI211_X1 U10190 ( .C1(n8775), .C2(n9195), .A(n8764), .B(n8763), .ZN(
        P2_U3480) );
  INV_X1 U10191 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8765) );
  MUX2_X1 U10192 ( .A(n8765), .B(n9196), .S(n10381), .Z(n8767) );
  NAND2_X1 U10193 ( .A1(n9198), .A2(n8768), .ZN(n8766) );
  OAI211_X1 U10194 ( .C1(n8775), .C2(n9201), .A(n8767), .B(n8766), .ZN(
        P2_U3479) );
  MUX2_X1 U10195 ( .A(n9081), .B(n9202), .S(n10381), .Z(n8770) );
  NAND2_X1 U10196 ( .A1(n9205), .A2(n8768), .ZN(n8769) );
  OAI211_X1 U10197 ( .C1(n8775), .C2(n9208), .A(n8770), .B(n8769), .ZN(
        P2_U3478) );
  INV_X1 U10198 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8773) );
  AOI21_X1 U10199 ( .B1(n10363), .B2(n8772), .A(n8771), .ZN(n9209) );
  MUX2_X1 U10200 ( .A(n8773), .B(n9209), .S(n10381), .Z(n8774) );
  OAI21_X1 U10201 ( .B1(n8775), .B2(n9213), .A(n8774), .ZN(P2_U3477) );
  NOR2_X1 U10202 ( .A1(n8776), .A2(n10366), .ZN(n8779) );
  AOI21_X1 U10203 ( .B1(n10366), .B2(P2_REG0_REG_31__SCAN_IN), .A(n8779), .ZN(
        n8777) );
  OAI21_X1 U10204 ( .B1(n8778), .B2(n9178), .A(n8777), .ZN(P2_U3458) );
  AOI21_X1 U10205 ( .B1(n10366), .B2(P2_REG0_REG_30__SCAN_IN), .A(n8779), .ZN(
        n8780) );
  OAI21_X1 U10206 ( .B1(n8781), .B2(n9178), .A(n8780), .ZN(P2_U3457) );
  OR2_X1 U10207 ( .A1(n10364), .A2(n8783), .ZN(n8784) );
  NAND2_X1 U10208 ( .A1(n8785), .A2(n8784), .ZN(n9155) );
  AOI22_X1 U10209 ( .A1(n5322), .A2(keyinput68), .B1(n9079), .B2(keyinput79), 
        .ZN(n8786) );
  OAI221_X1 U10210 ( .B1(n5322), .B2(keyinput68), .C1(n9079), .C2(keyinput79), 
        .A(n8786), .ZN(n8799) );
  AOI22_X1 U10211 ( .A1(n9084), .A2(keyinput2), .B1(keyinput34), .B2(n8788), 
        .ZN(n8787) );
  OAI221_X1 U10212 ( .B1(n9084), .B2(keyinput2), .C1(n8788), .C2(keyinput34), 
        .A(n8787), .ZN(n8798) );
  XNOR2_X1 U10213 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput70), .ZN(n8792) );
  XNOR2_X1 U10214 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput37), .ZN(n8791) );
  XNOR2_X1 U10215 ( .A(P2_REG2_REG_28__SCAN_IN), .B(keyinput96), .ZN(n8790) );
  XNOR2_X1 U10216 ( .A(P1_REG0_REG_29__SCAN_IN), .B(keyinput118), .ZN(n8789)
         );
  AND4_X1 U10217 ( .A1(n8792), .A2(n8791), .A3(n8790), .A4(n8789), .ZN(n8796)
         );
  XNOR2_X1 U10218 ( .A(keyinput15), .B(P1_REG2_REG_23__SCAN_IN), .ZN(n8795) );
  XNOR2_X1 U10219 ( .A(P1_REG2_REG_1__SCAN_IN), .B(keyinput20), .ZN(n8794) );
  XNOR2_X1 U10220 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(keyinput101), .ZN(n8793)
         );
  NAND4_X1 U10221 ( .A1(n8796), .A2(n8795), .A3(n8794), .A4(n8793), .ZN(n8797)
         );
  NOR3_X1 U10222 ( .A1(n8799), .A2(n8798), .A3(n8797), .ZN(n8820) );
  INV_X1 U10223 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n8801) );
  OAI22_X1 U10224 ( .A1(n8801), .A2(keyinput78), .B1(n9197), .B2(keyinput105), 
        .ZN(n8800) );
  AOI221_X1 U10225 ( .B1(n8801), .B2(keyinput78), .C1(keyinput105), .C2(n9197), 
        .A(n8800), .ZN(n8819) );
  XNOR2_X1 U10226 ( .A(P2_REG2_REG_2__SCAN_IN), .B(keyinput62), .ZN(n8805) );
  XNOR2_X1 U10227 ( .A(P1_REG1_REG_0__SCAN_IN), .B(keyinput102), .ZN(n8804) );
  XNOR2_X1 U10228 ( .A(P1_REG0_REG_30__SCAN_IN), .B(keyinput11), .ZN(n8803) );
  XNOR2_X1 U10229 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput123), .ZN(n8802)
         );
  NAND4_X1 U10230 ( .A1(n8805), .A2(n8804), .A3(n8803), .A4(n8802), .ZN(n8811)
         );
  XNOR2_X1 U10231 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(keyinput22), .ZN(n8809) );
  XNOR2_X1 U10232 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(keyinput23), .ZN(n8808) );
  XNOR2_X1 U10233 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput114), .ZN(n8807) );
  XNOR2_X1 U10234 ( .A(P2_IR_REG_27__SCAN_IN), .B(keyinput71), .ZN(n8806) );
  NAND4_X1 U10235 ( .A1(n8809), .A2(n8808), .A3(n8807), .A4(n8806), .ZN(n8810)
         );
  NOR2_X1 U10236 ( .A1(n8811), .A2(n8810), .ZN(n8818) );
  INV_X1 U10237 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10222) );
  AOI22_X1 U10238 ( .A1(n10222), .A2(keyinput81), .B1(keyinput29), .B2(n8813), 
        .ZN(n8812) );
  OAI221_X1 U10239 ( .B1(n10222), .B2(keyinput81), .C1(n8813), .C2(keyinput29), 
        .A(n8812), .ZN(n8816) );
  INV_X1 U10240 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n10054) );
  AOI22_X1 U10241 ( .A1(n8034), .A2(keyinput24), .B1(keyinput44), .B2(n10054), 
        .ZN(n8814) );
  OAI221_X1 U10242 ( .B1(n8034), .B2(keyinput24), .C1(n10054), .C2(keyinput44), 
        .A(n8814), .ZN(n8815) );
  NOR2_X1 U10243 ( .A1(n8816), .A2(n8815), .ZN(n8817) );
  AND4_X1 U10244 ( .A1(n8820), .A2(n8819), .A3(n8818), .A4(n8817), .ZN(n8829)
         );
  OAI22_X1 U10245 ( .A1(n8994), .A2(keyinput4), .B1(n5824), .B2(keyinput41), 
        .ZN(n8821) );
  AOI221_X1 U10246 ( .B1(n8994), .B2(keyinput4), .C1(keyinput41), .C2(n5824), 
        .A(n8821), .ZN(n8828) );
  INV_X1 U10247 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10090) );
  INV_X1 U10248 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n8823) );
  OAI22_X1 U10249 ( .A1(n10090), .A2(keyinput103), .B1(n8823), .B2(keyinput91), 
        .ZN(n8822) );
  AOI221_X1 U10250 ( .B1(n10090), .B2(keyinput103), .C1(keyinput91), .C2(n8823), .A(n8822), .ZN(n8827) );
  INV_X1 U10251 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8825) );
  OAI22_X1 U10252 ( .A1(n8825), .A2(keyinput93), .B1(n8965), .B2(keyinput60), 
        .ZN(n8824) );
  AOI221_X1 U10253 ( .B1(n8825), .B2(keyinput93), .C1(keyinput60), .C2(n8965), 
        .A(n8824), .ZN(n8826) );
  AND4_X1 U10254 ( .A1(n8829), .A2(n8828), .A3(n8827), .A4(n8826), .ZN(n8887)
         );
  INV_X1 U10255 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10209) );
  AOI22_X1 U10256 ( .A1(n8988), .A2(keyinput30), .B1(n10209), .B2(keyinput33), 
        .ZN(n8830) );
  OAI221_X1 U10257 ( .B1(n8988), .B2(keyinput30), .C1(n10209), .C2(keyinput33), 
        .A(n8830), .ZN(n8838) );
  AOI22_X1 U10258 ( .A1(n8833), .A2(keyinput115), .B1(keyinput26), .B2(n8832), 
        .ZN(n8831) );
  OAI221_X1 U10259 ( .B1(n8833), .B2(keyinput115), .C1(n8832), .C2(keyinput26), 
        .A(n8831), .ZN(n8837) );
  AOI22_X1 U10260 ( .A1(n8835), .A2(keyinput127), .B1(n9085), .B2(keyinput86), 
        .ZN(n8834) );
  OAI221_X1 U10261 ( .B1(n8835), .B2(keyinput127), .C1(n9085), .C2(keyinput86), 
        .A(n8834), .ZN(n8836) );
  NOR3_X1 U10262 ( .A1(n8838), .A2(n8837), .A3(n8836), .ZN(n8861) );
  INV_X1 U10263 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10291) );
  AOI22_X1 U10264 ( .A1(n10291), .A2(keyinput94), .B1(n8840), .B2(keyinput90), 
        .ZN(n8839) );
  OAI221_X1 U10265 ( .B1(n10291), .B2(keyinput94), .C1(n8840), .C2(keyinput90), 
        .A(n8839), .ZN(n8844) );
  AOI22_X1 U10266 ( .A1(n7051), .A2(keyinput122), .B1(n8842), .B2(keyinput61), 
        .ZN(n8841) );
  OAI221_X1 U10267 ( .B1(n7051), .B2(keyinput122), .C1(n8842), .C2(keyinput61), 
        .A(n8841), .ZN(n8843) );
  NOR2_X1 U10268 ( .A1(n8844), .A2(n8843), .ZN(n8860) );
  AOI22_X1 U10269 ( .A1(n9221), .A2(keyinput77), .B1(n8846), .B2(keyinput5), 
        .ZN(n8845) );
  OAI221_X1 U10270 ( .B1(n9221), .B2(keyinput77), .C1(n8846), .C2(keyinput5), 
        .A(n8845), .ZN(n8852) );
  AOI22_X1 U10271 ( .A1(n9168), .A2(keyinput16), .B1(n9265), .B2(keyinput12), 
        .ZN(n8847) );
  OAI221_X1 U10272 ( .B1(n9168), .B2(keyinput16), .C1(n9265), .C2(keyinput12), 
        .A(n8847), .ZN(n8851) );
  XNOR2_X1 U10273 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput43), .ZN(n8849) );
  XNOR2_X1 U10274 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput108), .ZN(n8848) );
  NAND2_X1 U10275 ( .A1(n8849), .A2(n8848), .ZN(n8850) );
  NOR3_X1 U10276 ( .A1(n8852), .A2(n8851), .A3(n8850), .ZN(n8859) );
  INV_X1 U10277 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9101) );
  AOI22_X1 U10278 ( .A1(n9101), .A2(keyinput36), .B1(keyinput99), .B2(n8854), 
        .ZN(n8853) );
  OAI221_X1 U10279 ( .B1(n9101), .B2(keyinput36), .C1(n8854), .C2(keyinput99), 
        .A(n8853), .ZN(n8857) );
  XNOR2_X1 U10280 ( .A(n8855), .B(keyinput97), .ZN(n8856) );
  NOR2_X1 U10281 ( .A1(n8857), .A2(n8856), .ZN(n8858) );
  AND4_X1 U10282 ( .A1(n8861), .A2(n8860), .A3(n8859), .A4(n8858), .ZN(n8872)
         );
  INV_X1 U10283 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n8864) );
  OAI22_X1 U10284 ( .A1(n8864), .A2(keyinput40), .B1(n8863), .B2(keyinput19), 
        .ZN(n8862) );
  AOI221_X1 U10285 ( .B1(n8864), .B2(keyinput40), .C1(keyinput19), .C2(n8863), 
        .A(n8862), .ZN(n8871) );
  OAI22_X1 U10286 ( .A1(n10286), .A2(keyinput38), .B1(n8866), .B2(keyinput32), 
        .ZN(n8865) );
  AOI221_X1 U10287 ( .B1(n10286), .B2(keyinput38), .C1(keyinput32), .C2(n8866), 
        .A(n8865), .ZN(n8870) );
  OAI22_X1 U10288 ( .A1(n5678), .A2(keyinput49), .B1(n8868), .B2(keyinput75), 
        .ZN(n8867) );
  AOI221_X1 U10289 ( .B1(n5678), .B2(keyinput49), .C1(keyinput75), .C2(n8868), 
        .A(n8867), .ZN(n8869) );
  AND4_X1 U10290 ( .A1(n8872), .A2(n8871), .A3(n8870), .A4(n8869), .ZN(n8886)
         );
  AOI22_X1 U10291 ( .A1(n8874), .A2(keyinput113), .B1(keyinput55), .B2(n7388), 
        .ZN(n8873) );
  OAI221_X1 U10292 ( .B1(n8874), .B2(keyinput113), .C1(n7388), .C2(keyinput55), 
        .A(n8873), .ZN(n8884) );
  AOI22_X1 U10293 ( .A1(n8877), .A2(keyinput107), .B1(keyinput59), .B2(n8876), 
        .ZN(n8875) );
  OAI221_X1 U10294 ( .B1(n8877), .B2(keyinput107), .C1(n8876), .C2(keyinput59), 
        .A(n8875), .ZN(n8883) );
  INV_X1 U10295 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10224) );
  AOI22_X1 U10296 ( .A1(n8879), .A2(keyinput119), .B1(n10224), .B2(keyinput65), 
        .ZN(n8878) );
  OAI221_X1 U10297 ( .B1(n8879), .B2(keyinput119), .C1(n10224), .C2(keyinput65), .A(n8878), .ZN(n8882) );
  INV_X1 U10298 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n10228) );
  AOI22_X1 U10299 ( .A1(n10228), .A2(keyinput27), .B1(keyinput106), .B2(n9071), 
        .ZN(n8880) );
  OAI221_X1 U10300 ( .B1(n10228), .B2(keyinput27), .C1(n9071), .C2(keyinput106), .A(n8880), .ZN(n8881) );
  NOR4_X1 U10301 ( .A1(n8884), .A2(n8883), .A3(n8882), .A4(n8881), .ZN(n8885)
         );
  AND3_X1 U10302 ( .A1(n8887), .A2(n8886), .A3(n8885), .ZN(n9153) );
  OAI22_X1 U10303 ( .A1(P2_D_REG_3__SCAN_IN), .A2(keyinput53), .B1(keyinput100), .B2(P2_REG3_REG_12__SCAN_IN), .ZN(n8888) );
  AOI221_X1 U10304 ( .B1(P2_D_REG_3__SCAN_IN), .B2(keyinput53), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput100), .A(n8888), .ZN(n8895) );
  OAI22_X1 U10305 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(keyinput76), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(keyinput104), .ZN(n8889) );
  AOI221_X1 U10306 ( .B1(P1_DATAO_REG_21__SCAN_IN), .B2(keyinput76), .C1(
        keyinput104), .C2(P1_DATAO_REG_15__SCAN_IN), .A(n8889), .ZN(n8894) );
  OAI22_X1 U10307 ( .A1(P1_REG0_REG_9__SCAN_IN), .A2(keyinput54), .B1(
        P1_ADDR_REG_2__SCAN_IN), .B2(keyinput110), .ZN(n8890) );
  AOI221_X1 U10308 ( .B1(P1_REG0_REG_9__SCAN_IN), .B2(keyinput54), .C1(
        keyinput110), .C2(P1_ADDR_REG_2__SCAN_IN), .A(n8890), .ZN(n8893) );
  OAI22_X1 U10309 ( .A1(SI_24_), .A2(keyinput52), .B1(keyinput14), .B2(
        P2_REG0_REG_5__SCAN_IN), .ZN(n8891) );
  AOI221_X1 U10310 ( .B1(SI_24_), .B2(keyinput52), .C1(P2_REG0_REG_5__SCAN_IN), 
        .C2(keyinput14), .A(n8891), .ZN(n8892) );
  NAND4_X1 U10311 ( .A1(n8895), .A2(n8894), .A3(n8893), .A4(n8892), .ZN(n8923)
         );
  OAI22_X1 U10312 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(keyinput51), .B1(
        keyinput56), .B2(P1_RD_REG_SCAN_IN), .ZN(n8896) );
  AOI221_X1 U10313 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(keyinput51), .C1(
        P1_RD_REG_SCAN_IN), .C2(keyinput56), .A(n8896), .ZN(n8903) );
  OAI22_X1 U10314 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(keyinput82), .B1(
        P2_REG1_REG_13__SCAN_IN), .B2(keyinput46), .ZN(n8897) );
  AOI221_X1 U10315 ( .B1(P2_IR_REG_1__SCAN_IN), .B2(keyinput82), .C1(
        keyinput46), .C2(P2_REG1_REG_13__SCAN_IN), .A(n8897), .ZN(n8902) );
  OAI22_X1 U10316 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(keyinput48), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(keyinput88), .ZN(n8898) );
  AOI221_X1 U10317 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput48), .C1(
        keyinput88), .C2(P2_REG3_REG_1__SCAN_IN), .A(n8898), .ZN(n8901) );
  OAI22_X1 U10318 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(keyinput31), .B1(
        keyinput85), .B2(P1_REG3_REG_10__SCAN_IN), .ZN(n8899) );
  AOI221_X1 U10319 ( .B1(P1_IR_REG_26__SCAN_IN), .B2(keyinput31), .C1(
        P1_REG3_REG_10__SCAN_IN), .C2(keyinput85), .A(n8899), .ZN(n8900) );
  NAND4_X1 U10320 ( .A1(n8903), .A2(n8902), .A3(n8901), .A4(n8900), .ZN(n8922)
         );
  OAI22_X1 U10321 ( .A1(SI_20_), .A2(keyinput58), .B1(keyinput50), .B2(SI_0_), 
        .ZN(n8904) );
  AOI221_X1 U10322 ( .B1(SI_20_), .B2(keyinput58), .C1(SI_0_), .C2(keyinput50), 
        .A(n8904), .ZN(n8911) );
  OAI22_X1 U10323 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(keyinput84), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(keyinput109), .ZN(n8905) );
  AOI221_X1 U10324 ( .B1(P2_IR_REG_17__SCAN_IN), .B2(keyinput84), .C1(
        keyinput109), .C2(P2_REG3_REG_0__SCAN_IN), .A(n8905), .ZN(n8910) );
  OAI22_X1 U10325 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(keyinput69), .B1(
        keyinput80), .B2(P1_REG1_REG_18__SCAN_IN), .ZN(n8906) );
  AOI221_X1 U10326 ( .B1(P1_IR_REG_27__SCAN_IN), .B2(keyinput69), .C1(
        P1_REG1_REG_18__SCAN_IN), .C2(keyinput80), .A(n8906), .ZN(n8909) );
  OAI22_X1 U10327 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(keyinput95), .B1(
        keyinput124), .B2(P2_REG1_REG_16__SCAN_IN), .ZN(n8907) );
  AOI221_X1 U10328 ( .B1(P1_DATAO_REG_2__SCAN_IN), .B2(keyinput95), .C1(
        P2_REG1_REG_16__SCAN_IN), .C2(keyinput124), .A(n8907), .ZN(n8908) );
  NAND4_X1 U10329 ( .A1(n8911), .A2(n8910), .A3(n8909), .A4(n8908), .ZN(n8921)
         );
  OAI22_X1 U10330 ( .A1(P2_REG0_REG_2__SCAN_IN), .A2(keyinput66), .B1(
        P2_REG1_REG_23__SCAN_IN), .B2(keyinput42), .ZN(n8912) );
  AOI221_X1 U10331 ( .B1(P2_REG0_REG_2__SCAN_IN), .B2(keyinput66), .C1(
        keyinput42), .C2(P2_REG1_REG_23__SCAN_IN), .A(n8912), .ZN(n8919) );
  OAI22_X1 U10332 ( .A1(P1_REG2_REG_19__SCAN_IN), .A2(keyinput116), .B1(
        P2_D_REG_25__SCAN_IN), .B2(keyinput47), .ZN(n8913) );
  AOI221_X1 U10333 ( .B1(P1_REG2_REG_19__SCAN_IN), .B2(keyinput116), .C1(
        keyinput47), .C2(P2_D_REG_25__SCAN_IN), .A(n8913), .ZN(n8918) );
  OAI22_X1 U10334 ( .A1(P1_D_REG_12__SCAN_IN), .A2(keyinput10), .B1(
        P2_REG2_REG_31__SCAN_IN), .B2(keyinput64), .ZN(n8914) );
  AOI221_X1 U10335 ( .B1(P1_D_REG_12__SCAN_IN), .B2(keyinput10), .C1(
        keyinput64), .C2(P2_REG2_REG_31__SCAN_IN), .A(n8914), .ZN(n8917) );
  OAI22_X1 U10336 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(keyinput98), .B1(
        P2_D_REG_11__SCAN_IN), .B2(keyinput17), .ZN(n8915) );
  AOI221_X1 U10337 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(keyinput98), .C1(
        keyinput17), .C2(P2_D_REG_11__SCAN_IN), .A(n8915), .ZN(n8916) );
  NAND4_X1 U10338 ( .A1(n8919), .A2(n8918), .A3(n8917), .A4(n8916), .ZN(n8920)
         );
  NOR4_X1 U10339 ( .A1(n8923), .A2(n8922), .A3(n8921), .A4(n8920), .ZN(n9152)
         );
  OAI22_X1 U10340 ( .A1(P2_REG0_REG_27__SCAN_IN), .A2(keyinput126), .B1(
        keyinput112), .B2(P2_REG2_REG_17__SCAN_IN), .ZN(n8924) );
  AOI221_X1 U10341 ( .B1(P2_REG0_REG_27__SCAN_IN), .B2(keyinput126), .C1(
        P2_REG2_REG_17__SCAN_IN), .C2(keyinput112), .A(n8924), .ZN(n8931) );
  OAI22_X1 U10342 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(keyinput73), .B1(
        P1_REG0_REG_25__SCAN_IN), .B2(keyinput89), .ZN(n8925) );
  AOI221_X1 U10343 ( .B1(P1_REG3_REG_9__SCAN_IN), .B2(keyinput73), .C1(
        keyinput89), .C2(P1_REG0_REG_25__SCAN_IN), .A(n8925), .ZN(n8930) );
  OAI22_X1 U10344 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput72), .B1(
        P2_ADDR_REG_3__SCAN_IN), .B2(keyinput6), .ZN(n8926) );
  AOI221_X1 U10345 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput72), .C1(
        keyinput6), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n8926), .ZN(n8929) );
  OAI22_X1 U10346 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(keyinput125), .B1(
        keyinput87), .B2(P2_D_REG_15__SCAN_IN), .ZN(n8927) );
  AOI221_X1 U10347 ( .B1(P2_IR_REG_2__SCAN_IN), .B2(keyinput125), .C1(
        P2_D_REG_15__SCAN_IN), .C2(keyinput87), .A(n8927), .ZN(n8928) );
  NAND4_X1 U10348 ( .A1(n8931), .A2(n8930), .A3(n8929), .A4(n8928), .ZN(n8960)
         );
  OAI22_X1 U10349 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(keyinput67), .B1(
        P1_REG3_REG_5__SCAN_IN), .B2(keyinput21), .ZN(n8932) );
  AOI221_X1 U10350 ( .B1(P2_DATAO_REG_12__SCAN_IN), .B2(keyinput67), .C1(
        keyinput21), .C2(P1_REG3_REG_5__SCAN_IN), .A(n8932), .ZN(n8939) );
  OAI22_X1 U10351 ( .A1(P2_D_REG_24__SCAN_IN), .A2(keyinput28), .B1(
        P2_REG1_REG_19__SCAN_IN), .B2(keyinput92), .ZN(n8933) );
  AOI221_X1 U10352 ( .B1(P2_D_REG_24__SCAN_IN), .B2(keyinput28), .C1(
        keyinput92), .C2(P2_REG1_REG_19__SCAN_IN), .A(n8933), .ZN(n8938) );
  OAI22_X1 U10353 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(keyinput35), .B1(
        P2_IR_REG_19__SCAN_IN), .B2(keyinput39), .ZN(n8934) );
  AOI221_X1 U10354 ( .B1(P1_IR_REG_22__SCAN_IN), .B2(keyinput35), .C1(
        keyinput39), .C2(P2_IR_REG_19__SCAN_IN), .A(n8934), .ZN(n8937) );
  OAI22_X1 U10355 ( .A1(P1_D_REG_3__SCAN_IN), .A2(keyinput121), .B1(SI_13_), 
        .B2(keyinput18), .ZN(n8935) );
  AOI221_X1 U10356 ( .B1(P1_D_REG_3__SCAN_IN), .B2(keyinput121), .C1(
        keyinput18), .C2(SI_13_), .A(n8935), .ZN(n8936) );
  NAND4_X1 U10357 ( .A1(n8939), .A2(n8938), .A3(n8937), .A4(n8936), .ZN(n8959)
         );
  OAI22_X1 U10358 ( .A1(SI_12_), .A2(keyinput74), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(keyinput63), .ZN(n8940) );
  AOI221_X1 U10359 ( .B1(SI_12_), .B2(keyinput74), .C1(keyinput63), .C2(
        P2_REG3_REG_28__SCAN_IN), .A(n8940), .ZN(n8948) );
  OAI22_X1 U10360 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(keyinput117), .B1(keyinput0), .B2(P2_REG0_REG_0__SCAN_IN), .ZN(n8941) );
  AOI221_X1 U10361 ( .B1(P1_IR_REG_7__SCAN_IN), .B2(keyinput117), .C1(
        P2_REG0_REG_0__SCAN_IN), .C2(keyinput0), .A(n8941), .ZN(n8947) );
  INV_X1 U10362 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10096) );
  OAI22_X1 U10363 ( .A1(n9073), .A2(keyinput25), .B1(n10096), .B2(keyinput83), 
        .ZN(n8942) );
  AOI221_X1 U10364 ( .B1(n9073), .B2(keyinput25), .C1(keyinput83), .C2(n10096), 
        .A(n8942), .ZN(n8946) );
  INV_X1 U10365 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n8944) );
  OAI22_X1 U10366 ( .A1(n8944), .A2(keyinput3), .B1(n9210), .B2(keyinput7), 
        .ZN(n8943) );
  AOI221_X1 U10367 ( .B1(n8944), .B2(keyinput3), .C1(keyinput7), .C2(n9210), 
        .A(n8943), .ZN(n8945) );
  NAND4_X1 U10368 ( .A1(n8948), .A2(n8947), .A3(n8946), .A4(n8945), .ZN(n8958)
         );
  OAI22_X1 U10369 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(keyinput13), .B1(
        keyinput120), .B2(P1_REG3_REG_20__SCAN_IN), .ZN(n8949) );
  AOI221_X1 U10370 ( .B1(P1_IR_REG_10__SCAN_IN), .B2(keyinput13), .C1(
        P1_REG3_REG_20__SCAN_IN), .C2(keyinput120), .A(n8949), .ZN(n8956) );
  OAI22_X1 U10371 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput8), .B1(
        keyinput45), .B2(P2_REG1_REG_14__SCAN_IN), .ZN(n8950) );
  AOI221_X1 U10372 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput8), .C1(
        P2_REG1_REG_14__SCAN_IN), .C2(keyinput45), .A(n8950), .ZN(n8955) );
  OAI22_X1 U10373 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(keyinput111), .B1(
        keyinput9), .B2(P2_ADDR_REG_13__SCAN_IN), .ZN(n8951) );
  AOI221_X1 U10374 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(keyinput111), .C1(
        P2_ADDR_REG_13__SCAN_IN), .C2(keyinput9), .A(n8951), .ZN(n8954) );
  OAI22_X1 U10375 ( .A1(P1_REG2_REG_25__SCAN_IN), .A2(keyinput1), .B1(
        keyinput57), .B2(P2_REG0_REG_23__SCAN_IN), .ZN(n8952) );
  AOI221_X1 U10376 ( .B1(P1_REG2_REG_25__SCAN_IN), .B2(keyinput1), .C1(
        P2_REG0_REG_23__SCAN_IN), .C2(keyinput57), .A(n8952), .ZN(n8953) );
  NAND4_X1 U10377 ( .A1(n8956), .A2(n8955), .A3(n8954), .A4(n8953), .ZN(n8957)
         );
  NOR4_X1 U10378 ( .A1(n8960), .A2(n8959), .A3(n8958), .A4(n8957), .ZN(n9151)
         );
  AOI22_X1 U10379 ( .A1(n10291), .A2(keyinput222), .B1(keyinput224), .B2(n8962), .ZN(n8961) );
  OAI221_X1 U10380 ( .B1(n10291), .B2(keyinput222), .C1(n8962), .C2(
        keyinput224), .A(n8961), .ZN(n8963) );
  INV_X1 U10381 ( .A(n8963), .ZN(n8976) );
  INV_X1 U10382 ( .A(keyinput188), .ZN(n8964) );
  XNOR2_X1 U10383 ( .A(n8965), .B(n8964), .ZN(n8975) );
  XNOR2_X1 U10384 ( .A(keyinput152), .B(n8034), .ZN(n8968) );
  INV_X1 U10385 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n8966) );
  XNOR2_X1 U10386 ( .A(keyinput238), .B(n8966), .ZN(n8967) );
  NOR2_X1 U10387 ( .A1(n8968), .A2(n8967), .ZN(n8974) );
  AOI22_X1 U10388 ( .A1(n8971), .A2(keyinput170), .B1(n8970), .B2(keyinput149), 
        .ZN(n8969) );
  OAI221_X1 U10389 ( .B1(n8971), .B2(keyinput170), .C1(n8970), .C2(keyinput149), .A(n8969), .ZN(n8972) );
  INV_X1 U10390 ( .A(n8972), .ZN(n8973) );
  NAND4_X1 U10391 ( .A1(n8976), .A2(n8975), .A3(n8974), .A4(n8973), .ZN(n8992)
         );
  XNOR2_X1 U10392 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput159), .ZN(n8980) );
  XNOR2_X1 U10393 ( .A(SI_0_), .B(keyinput178), .ZN(n8979) );
  XNOR2_X1 U10394 ( .A(P2_REG2_REG_2__SCAN_IN), .B(keyinput190), .ZN(n8978) );
  XNOR2_X1 U10395 ( .A(P1_REG1_REG_13__SCAN_IN), .B(keyinput247), .ZN(n8977)
         );
  NAND4_X1 U10396 ( .A1(n8980), .A2(n8979), .A3(n8978), .A4(n8977), .ZN(n8986)
         );
  XNOR2_X1 U10397 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput237), .ZN(n8984) );
  XNOR2_X1 U10398 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(keyinput162), .ZN(n8983)
         );
  XNOR2_X1 U10399 ( .A(keyinput143), .B(P1_REG2_REG_23__SCAN_IN), .ZN(n8982)
         );
  XNOR2_X1 U10400 ( .A(keyinput184), .B(P1_RD_REG_SCAN_IN), .ZN(n8981) );
  NAND4_X1 U10401 ( .A1(n8984), .A2(n8983), .A3(n8982), .A4(n8981), .ZN(n8985)
         );
  NOR2_X1 U10402 ( .A1(n8986), .A2(n8985), .ZN(n8990) );
  INV_X1 U10403 ( .A(keyinput158), .ZN(n8987) );
  XNOR2_X1 U10404 ( .A(n8988), .B(n8987), .ZN(n8989) );
  NAND2_X1 U10405 ( .A1(n8990), .A2(n8989), .ZN(n8991) );
  NOR2_X1 U10406 ( .A1(n8992), .A2(n8991), .ZN(n9025) );
  AOI22_X1 U10407 ( .A1(n8994), .A2(keyinput132), .B1(keyinput166), .B2(n10286), .ZN(n8993) );
  OAI221_X1 U10408 ( .B1(n8994), .B2(keyinput132), .C1(n10286), .C2(
        keyinput166), .A(n8993), .ZN(n9001) );
  INV_X1 U10409 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10234) );
  AOI22_X1 U10410 ( .A1(n10234), .A2(keyinput249), .B1(keyinput176), .B2(n8996), .ZN(n8995) );
  OAI221_X1 U10411 ( .B1(n10234), .B2(keyinput249), .C1(n8996), .C2(
        keyinput176), .A(n8995), .ZN(n9000) );
  AOI22_X1 U10412 ( .A1(n5391), .A2(keyinput134), .B1(n8998), .B2(keyinput195), 
        .ZN(n8997) );
  OAI221_X1 U10413 ( .B1(n5391), .B2(keyinput134), .C1(n8998), .C2(keyinput195), .A(n8997), .ZN(n8999) );
  NOR3_X1 U10414 ( .A1(n9001), .A2(n9000), .A3(n8999), .ZN(n9024) );
  XNOR2_X1 U10415 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput251), .ZN(n9005)
         );
  XNOR2_X1 U10416 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(keyinput151), .ZN(n9004)
         );
  XNOR2_X1 U10417 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput160), .ZN(n9003) );
  XNOR2_X1 U10418 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput167), .ZN(n9002) );
  NAND4_X1 U10419 ( .A1(n9005), .A2(n9004), .A3(n9003), .A4(n9002), .ZN(n9011)
         );
  XNOR2_X1 U10420 ( .A(P1_REG0_REG_23__SCAN_IN), .B(keyinput189), .ZN(n9009)
         );
  XNOR2_X1 U10421 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(keyinput150), .ZN(n9008)
         );
  XNOR2_X1 U10422 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput141), .ZN(n9007) );
  XNOR2_X1 U10423 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput198), .ZN(n9006) );
  NAND4_X1 U10424 ( .A1(n9009), .A2(n9008), .A3(n9007), .A4(n9006), .ZN(n9010)
         );
  NOR2_X1 U10425 ( .A1(n9011), .A2(n9010), .ZN(n9023) );
  XNOR2_X1 U10426 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput163), .ZN(n9015) );
  XNOR2_X1 U10427 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput236), .ZN(n9014) );
  XNOR2_X1 U10428 ( .A(P2_REG1_REG_30__SCAN_IN), .B(keyinput203), .ZN(n9013)
         );
  XNOR2_X1 U10429 ( .A(P1_REG1_REG_29__SCAN_IN), .B(keyinput131), .ZN(n9012)
         );
  NAND4_X1 U10430 ( .A1(n9015), .A2(n9014), .A3(n9013), .A4(n9012), .ZN(n9021)
         );
  XNOR2_X1 U10431 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput171), .ZN(n9019) );
  XNOR2_X1 U10432 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput216), .ZN(n9018) );
  XNOR2_X1 U10433 ( .A(P1_REG2_REG_1__SCAN_IN), .B(keyinput148), .ZN(n9017) );
  XNOR2_X1 U10434 ( .A(P2_IR_REG_1__SCAN_IN), .B(keyinput210), .ZN(n9016) );
  NAND4_X1 U10435 ( .A1(n9019), .A2(n9018), .A3(n9017), .A4(n9016), .ZN(n9020)
         );
  NOR2_X1 U10436 ( .A1(n9021), .A2(n9020), .ZN(n9022) );
  NAND4_X1 U10437 ( .A1(n9025), .A2(n9024), .A3(n9023), .A4(n9022), .ZN(n9063)
         );
  AOI22_X1 U10438 ( .A1(P1_REG2_REG_25__SCAN_IN), .A2(keyinput129), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(keyinput204), .ZN(n9026) );
  OAI221_X1 U10439 ( .B1(P1_REG2_REG_25__SCAN_IN), .B2(keyinput129), .C1(
        P1_DATAO_REG_21__SCAN_IN), .C2(keyinput204), .A(n9026), .ZN(n9033) );
  AOI22_X1 U10440 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(keyinput183), .B1(
        P2_IR_REG_27__SCAN_IN), .B2(keyinput199), .ZN(n9027) );
  OAI221_X1 U10441 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(keyinput183), .C1(
        P2_IR_REG_27__SCAN_IN), .C2(keyinput199), .A(n9027), .ZN(n9032) );
  AOI22_X1 U10442 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput228), .B1(
        P1_REG1_REG_0__SCAN_IN), .B2(keyinput230), .ZN(n9028) );
  OAI221_X1 U10443 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput228), .C1(
        P1_REG1_REG_0__SCAN_IN), .C2(keyinput230), .A(n9028), .ZN(n9031) );
  AOI22_X1 U10444 ( .A1(P2_REG0_REG_20__SCAN_IN), .A2(keyinput233), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(keyinput235), .ZN(n9029) );
  OAI221_X1 U10445 ( .B1(P2_REG0_REG_20__SCAN_IN), .B2(keyinput233), .C1(
        P2_DATAO_REG_16__SCAN_IN), .C2(keyinput235), .A(n9029), .ZN(n9030) );
  NOR4_X1 U10446 ( .A1(n9033), .A2(n9032), .A3(n9031), .A4(n9030), .ZN(n9061)
         );
  AOI22_X1 U10447 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(keyinput174), .B1(
        P2_D_REG_3__SCAN_IN), .B2(keyinput181), .ZN(n9034) );
  OAI221_X1 U10448 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(keyinput174), .C1(
        P2_D_REG_3__SCAN_IN), .C2(keyinput181), .A(n9034), .ZN(n9041) );
  AOI22_X1 U10449 ( .A1(P1_REG0_REG_29__SCAN_IN), .A2(keyinput246), .B1(
        P1_IR_REG_7__SCAN_IN), .B2(keyinput245), .ZN(n9035) );
  OAI221_X1 U10450 ( .B1(P1_REG0_REG_29__SCAN_IN), .B2(keyinput246), .C1(
        P1_IR_REG_7__SCAN_IN), .C2(keyinput245), .A(n9035), .ZN(n9040) );
  AOI22_X1 U10451 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput191), .B1(
        P1_REG0_REG_11__SCAN_IN), .B2(keyinput133), .ZN(n9036) );
  OAI221_X1 U10452 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput191), .C1(
        P1_REG0_REG_11__SCAN_IN), .C2(keyinput133), .A(n9036), .ZN(n9039) );
  AOI22_X1 U10453 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(keyinput221), .B1(SI_20_), .B2(keyinput186), .ZN(n9037) );
  OAI221_X1 U10454 ( .B1(P1_REG3_REG_15__SCAN_IN), .B2(keyinput221), .C1(
        SI_20_), .C2(keyinput186), .A(n9037), .ZN(n9038) );
  NOR4_X1 U10455 ( .A1(n9041), .A2(n9040), .A3(n9039), .A4(n9038), .ZN(n9060)
         );
  AOI22_X1 U10456 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(keyinput177), .B1(
        P1_REG1_REG_18__SCAN_IN), .B2(keyinput208), .ZN(n9042) );
  OAI221_X1 U10457 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(keyinput177), .C1(
        P1_REG1_REG_18__SCAN_IN), .C2(keyinput208), .A(n9042), .ZN(n9049) );
  AOI22_X1 U10458 ( .A1(P2_REG0_REG_26__SCAN_IN), .A2(keyinput144), .B1(
        P1_IR_REG_27__SCAN_IN), .B2(keyinput197), .ZN(n9043) );
  OAI221_X1 U10459 ( .B1(P2_REG0_REG_26__SCAN_IN), .B2(keyinput144), .C1(
        P1_IR_REG_27__SCAN_IN), .C2(keyinput197), .A(n9043), .ZN(n9048) );
  AOI22_X1 U10460 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(keyinput205), .B1(
        P1_D_REG_12__SCAN_IN), .B2(keyinput138), .ZN(n9044) );
  OAI221_X1 U10461 ( .B1(P1_DATAO_REG_30__SCAN_IN), .B2(keyinput205), .C1(
        P1_D_REG_12__SCAN_IN), .C2(keyinput138), .A(n9044), .ZN(n9047) );
  AOI22_X1 U10462 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(keyinput187), .B1(
        P1_REG2_REG_9__SCAN_IN), .B2(keyinput226), .ZN(n9045) );
  OAI221_X1 U10463 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(keyinput187), .C1(
        P1_REG2_REG_9__SCAN_IN), .C2(keyinput226), .A(n9045), .ZN(n9046) );
  NOR4_X1 U10464 ( .A1(n9049), .A2(n9048), .A3(n9047), .A4(n9046), .ZN(n9059)
         );
  AOI22_X1 U10465 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(keyinput227), .B1(
        P2_REG1_REG_3__SCAN_IN), .B2(keyinput169), .ZN(n9050) );
  OAI221_X1 U10466 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(keyinput227), .C1(
        P2_REG1_REG_3__SCAN_IN), .C2(keyinput169), .A(n9050), .ZN(n9057) );
  AOI22_X1 U10467 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(keyinput253), .B1(
        P1_REG3_REG_17__SCAN_IN), .B2(keyinput243), .ZN(n9051) );
  OAI221_X1 U10468 ( .B1(P2_IR_REG_2__SCAN_IN), .B2(keyinput253), .C1(
        P1_REG3_REG_17__SCAN_IN), .C2(keyinput243), .A(n9051), .ZN(n9056) );
  AOI22_X1 U10469 ( .A1(P2_REG2_REG_31__SCAN_IN), .A2(keyinput192), .B1(
        P2_REG0_REG_0__SCAN_IN), .B2(keyinput128), .ZN(n9052) );
  OAI221_X1 U10470 ( .B1(P2_REG2_REG_31__SCAN_IN), .B2(keyinput192), .C1(
        P2_REG0_REG_0__SCAN_IN), .C2(keyinput128), .A(n9052), .ZN(n9055) );
  AOI22_X1 U10471 ( .A1(P2_D_REG_25__SCAN_IN), .A2(keyinput175), .B1(
        P1_IR_REG_31__SCAN_IN), .B2(keyinput179), .ZN(n9053) );
  OAI221_X1 U10472 ( .B1(P2_D_REG_25__SCAN_IN), .B2(keyinput175), .C1(
        P1_IR_REG_31__SCAN_IN), .C2(keyinput179), .A(n9053), .ZN(n9054) );
  NOR4_X1 U10473 ( .A1(n9057), .A2(n9056), .A3(n9055), .A4(n9054), .ZN(n9058)
         );
  NAND4_X1 U10474 ( .A1(n9061), .A2(n9060), .A3(n9059), .A4(n9058), .ZN(n9062)
         );
  NOR2_X1 U10475 ( .A1(n9063), .A2(n9062), .ZN(n9149) );
  INV_X1 U10476 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9066) );
  AOI22_X1 U10477 ( .A1(n9066), .A2(keyinput244), .B1(n9065), .B2(keyinput180), 
        .ZN(n9064) );
  OAI221_X1 U10478 ( .B1(n9066), .B2(keyinput244), .C1(n9065), .C2(keyinput180), .A(n9064), .ZN(n9077) );
  INV_X1 U10479 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9303) );
  AOI22_X1 U10480 ( .A1(n9068), .A2(keyinput232), .B1(keyinput248), .B2(n9303), 
        .ZN(n9067) );
  OAI221_X1 U10481 ( .B1(n9068), .B2(keyinput232), .C1(n9303), .C2(keyinput248), .A(n9067), .ZN(n9076) );
  AOI22_X1 U10482 ( .A1(n9071), .A2(keyinput234), .B1(keyinput136), .B2(n9070), 
        .ZN(n9069) );
  OAI221_X1 U10483 ( .B1(n9071), .B2(keyinput234), .C1(n9070), .C2(keyinput136), .A(n9069), .ZN(n9075) );
  AOI22_X1 U10484 ( .A1(n5852), .A2(keyinput239), .B1(n9073), .B2(keyinput153), 
        .ZN(n9072) );
  OAI221_X1 U10485 ( .B1(n5852), .B2(keyinput239), .C1(n9073), .C2(keyinput153), .A(n9072), .ZN(n9074) );
  NOR4_X1 U10486 ( .A1(n9077), .A2(n9076), .A3(n9075), .A4(n9074), .ZN(n9148)
         );
  AOI22_X1 U10487 ( .A1(n9079), .A2(keyinput207), .B1(keyinput250), .B2(n7051), 
        .ZN(n9078) );
  OAI221_X1 U10488 ( .B1(n9079), .B2(keyinput207), .C1(n7051), .C2(keyinput250), .A(n9078), .ZN(n9088) );
  AOI22_X1 U10489 ( .A1(n9082), .A2(keyinput202), .B1(keyinput220), .B2(n9081), 
        .ZN(n9080) );
  OAI221_X1 U10490 ( .B1(n9082), .B2(keyinput202), .C1(n9081), .C2(keyinput220), .A(n9080), .ZN(n9087) );
  AOI22_X1 U10491 ( .A1(n9085), .A2(keyinput214), .B1(n9084), .B2(keyinput130), 
        .ZN(n9083) );
  OAI221_X1 U10492 ( .B1(n9085), .B2(keyinput214), .C1(n9084), .C2(keyinput130), .A(n9083), .ZN(n9086) );
  NOR3_X1 U10493 ( .A1(n9088), .A2(n9087), .A3(n9086), .ZN(n9108) );
  AOI22_X1 U10494 ( .A1(n9090), .A2(keyinput252), .B1(n10209), .B2(keyinput161), .ZN(n9089) );
  OAI221_X1 U10495 ( .B1(n9090), .B2(keyinput252), .C1(n10209), .C2(
        keyinput161), .A(n9089), .ZN(n9095) );
  INV_X1 U10496 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n9092) );
  AOI22_X1 U10497 ( .A1(n9093), .A2(keyinput200), .B1(keyinput137), .B2(n9092), 
        .ZN(n9091) );
  OAI221_X1 U10498 ( .B1(n9093), .B2(keyinput200), .C1(n9092), .C2(keyinput137), .A(n9091), .ZN(n9094) );
  NOR2_X1 U10499 ( .A1(n9095), .A2(n9094), .ZN(n9107) );
  AOI22_X1 U10500 ( .A1(n9162), .A2(keyinput254), .B1(keyinput194), .B2(n5813), 
        .ZN(n9096) );
  OAI221_X1 U10501 ( .B1(n9162), .B2(keyinput254), .C1(n5813), .C2(keyinput194), .A(n9096), .ZN(n9099) );
  AOI22_X1 U10502 ( .A1(P1_REG0_REG_14__SCAN_IN), .A2(keyinput206), .B1(n10224), .B2(keyinput193), .ZN(n9097) );
  OAI221_X1 U10503 ( .B1(P1_REG0_REG_14__SCAN_IN), .B2(keyinput206), .C1(
        n10224), .C2(keyinput193), .A(n9097), .ZN(n9098) );
  NOR2_X1 U10504 ( .A1(n9099), .A2(n9098), .ZN(n9106) );
  AOI22_X1 U10505 ( .A1(n9101), .A2(keyinput164), .B1(n10228), .B2(keyinput155), .ZN(n9100) );
  OAI221_X1 U10506 ( .B1(n9101), .B2(keyinput164), .C1(n10228), .C2(
        keyinput155), .A(n9100), .ZN(n9104) );
  INV_X1 U10507 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10127) );
  AOI22_X1 U10508 ( .A1(n10127), .A2(keyinput139), .B1(n10222), .B2(
        keyinput209), .ZN(n9102) );
  OAI221_X1 U10509 ( .B1(n10127), .B2(keyinput139), .C1(n10222), .C2(
        keyinput209), .A(n9102), .ZN(n9103) );
  NOR2_X1 U10510 ( .A1(n9104), .A2(n9103), .ZN(n9105) );
  NAND4_X1 U10511 ( .A1(n9108), .A2(n9107), .A3(n9106), .A4(n9105), .ZN(n9146)
         );
  AOI22_X1 U10512 ( .A1(P2_REG0_REG_5__SCAN_IN), .A2(keyinput142), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(keyinput218), .ZN(n9109) );
  OAI221_X1 U10513 ( .B1(P2_REG0_REG_5__SCAN_IN), .B2(keyinput142), .C1(
        P1_DATAO_REG_22__SCAN_IN), .C2(keyinput218), .A(n9109), .ZN(n9116) );
  AOI22_X1 U10514 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(keyinput241), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(keyinput229), .ZN(n9110) );
  OAI221_X1 U10515 ( .B1(P1_DATAO_REG_14__SCAN_IN), .B2(keyinput241), .C1(
        P1_DATAO_REG_19__SCAN_IN), .C2(keyinput229), .A(n9110), .ZN(n9115) );
  AOI22_X1 U10516 ( .A1(P1_REG1_REG_27__SCAN_IN), .A2(keyinput172), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(keyinput223), .ZN(n9111) );
  OAI221_X1 U10517 ( .B1(P1_REG1_REG_27__SCAN_IN), .B2(keyinput172), .C1(
        P1_DATAO_REG_2__SCAN_IN), .C2(keyinput223), .A(n9111), .ZN(n9114) );
  AOI22_X1 U10518 ( .A1(P1_REG1_REG_20__SCAN_IN), .A2(keyinput231), .B1(
        P1_IR_REG_13__SCAN_IN), .B2(keyinput242), .ZN(n9112) );
  OAI221_X1 U10519 ( .B1(P1_REG1_REG_20__SCAN_IN), .B2(keyinput231), .C1(
        P1_IR_REG_13__SCAN_IN), .C2(keyinput242), .A(n9112), .ZN(n9113) );
  NOR4_X1 U10520 ( .A1(n9116), .A2(n9115), .A3(n9114), .A4(n9113), .ZN(n9144)
         );
  AOI22_X1 U10521 ( .A1(P2_B_REG_SCAN_IN), .A2(keyinput147), .B1(
        P1_REG3_REG_10__SCAN_IN), .B2(keyinput213), .ZN(n9117) );
  OAI221_X1 U10522 ( .B1(P2_B_REG_SCAN_IN), .B2(keyinput147), .C1(
        P1_REG3_REG_10__SCAN_IN), .C2(keyinput213), .A(n9117), .ZN(n9124) );
  AOI22_X1 U10523 ( .A1(P2_D_REG_15__SCAN_IN), .A2(keyinput215), .B1(
        P1_REG0_REG_25__SCAN_IN), .B2(keyinput217), .ZN(n9118) );
  OAI221_X1 U10524 ( .B1(P2_D_REG_15__SCAN_IN), .B2(keyinput215), .C1(
        P1_REG0_REG_25__SCAN_IN), .C2(keyinput217), .A(n9118), .ZN(n9123) );
  AOI22_X1 U10525 ( .A1(P2_REG0_REG_23__SCAN_IN), .A2(keyinput185), .B1(
        P2_REG1_REG_14__SCAN_IN), .B2(keyinput173), .ZN(n9119) );
  OAI221_X1 U10526 ( .B1(P2_REG0_REG_23__SCAN_IN), .B2(keyinput185), .C1(
        P2_REG1_REG_14__SCAN_IN), .C2(keyinput173), .A(n9119), .ZN(n9122) );
  AOI22_X1 U10527 ( .A1(P2_REG1_REG_24__SCAN_IN), .A2(keyinput157), .B1(
        P1_REG1_REG_19__SCAN_IN), .B2(keyinput211), .ZN(n9120) );
  OAI221_X1 U10528 ( .B1(P2_REG1_REG_24__SCAN_IN), .B2(keyinput157), .C1(
        P1_REG1_REG_19__SCAN_IN), .C2(keyinput211), .A(n9120), .ZN(n9121) );
  NOR4_X1 U10529 ( .A1(n9124), .A2(n9123), .A3(n9122), .A4(n9121), .ZN(n9143)
         );
  AOI22_X1 U10530 ( .A1(P2_D_REG_14__SCAN_IN), .A2(keyinput225), .B1(
        P2_D_REG_24__SCAN_IN), .B2(keyinput156), .ZN(n9125) );
  OAI221_X1 U10531 ( .B1(P2_D_REG_14__SCAN_IN), .B2(keyinput225), .C1(
        P2_D_REG_24__SCAN_IN), .C2(keyinput156), .A(n9125), .ZN(n9132) );
  AOI22_X1 U10532 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(keyinput240), .B1(
        P2_REG0_REG_18__SCAN_IN), .B2(keyinput135), .ZN(n9126) );
  OAI221_X1 U10533 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(keyinput240), .C1(
        P2_REG0_REG_18__SCAN_IN), .C2(keyinput135), .A(n9126), .ZN(n9131) );
  AOI22_X1 U10534 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(keyinput212), .B1(
        P1_REG1_REG_15__SCAN_IN), .B2(keyinput255), .ZN(n9127) );
  OAI221_X1 U10535 ( .B1(P2_IR_REG_17__SCAN_IN), .B2(keyinput212), .C1(
        P1_REG1_REG_15__SCAN_IN), .C2(keyinput255), .A(n9127), .ZN(n9130) );
  AOI22_X1 U10536 ( .A1(P2_D_REG_11__SCAN_IN), .A2(keyinput145), .B1(
        P1_REG0_REG_9__SCAN_IN), .B2(keyinput182), .ZN(n9128) );
  OAI221_X1 U10537 ( .B1(P2_D_REG_11__SCAN_IN), .B2(keyinput145), .C1(
        P1_REG0_REG_9__SCAN_IN), .C2(keyinput182), .A(n9128), .ZN(n9129) );
  NOR4_X1 U10538 ( .A1(n9132), .A2(n9131), .A3(n9130), .A4(n9129), .ZN(n9142)
         );
  AOI22_X1 U10539 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(keyinput140), .B1(
        P1_IR_REG_0__SCAN_IN), .B2(keyinput165), .ZN(n9133) );
  OAI221_X1 U10540 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(keyinput140), .C1(
        P1_IR_REG_0__SCAN_IN), .C2(keyinput165), .A(n9133), .ZN(n9140) );
  AOI22_X1 U10541 ( .A1(P1_REG2_REG_31__SCAN_IN), .A2(keyinput219), .B1(
        P2_REG0_REG_8__SCAN_IN), .B2(keyinput196), .ZN(n9134) );
  OAI221_X1 U10542 ( .B1(P1_REG2_REG_31__SCAN_IN), .B2(keyinput219), .C1(
        P2_REG0_REG_8__SCAN_IN), .C2(keyinput196), .A(n9134), .ZN(n9139) );
  AOI22_X1 U10543 ( .A1(P1_REG1_REG_26__SCAN_IN), .A2(keyinput168), .B1(SI_13_), .B2(keyinput146), .ZN(n9135) );
  OAI221_X1 U10544 ( .B1(P1_REG1_REG_26__SCAN_IN), .B2(keyinput168), .C1(
        SI_13_), .C2(keyinput146), .A(n9135), .ZN(n9138) );
  AOI22_X1 U10545 ( .A1(P2_REG0_REG_22__SCAN_IN), .A2(keyinput154), .B1(
        P1_REG3_REG_9__SCAN_IN), .B2(keyinput201), .ZN(n9136) );
  OAI221_X1 U10546 ( .B1(P2_REG0_REG_22__SCAN_IN), .B2(keyinput154), .C1(
        P1_REG3_REG_9__SCAN_IN), .C2(keyinput201), .A(n9136), .ZN(n9137) );
  NOR4_X1 U10547 ( .A1(n9140), .A2(n9139), .A3(n9138), .A4(n9137), .ZN(n9141)
         );
  NAND4_X1 U10548 ( .A1(n9144), .A2(n9143), .A3(n9142), .A4(n9141), .ZN(n9145)
         );
  NOR2_X1 U10549 ( .A1(n9146), .A2(n9145), .ZN(n9147) );
  NAND3_X1 U10550 ( .A1(n9149), .A2(n9148), .A3(n9147), .ZN(n9150) );
  NAND4_X1 U10551 ( .A1(n9153), .A2(n9152), .A3(n9151), .A4(n9150), .ZN(n9154)
         );
  XNOR2_X1 U10552 ( .A(n9155), .B(n9154), .ZN(P2_U3456) );
  MUX2_X1 U10553 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9156), .S(n10364), .Z(
        n9160) );
  OAI22_X1 U10554 ( .A1(n9158), .A2(n9212), .B1(n9157), .B2(n9178), .ZN(n9159)
         );
  OR2_X1 U10555 ( .A1(n9160), .A2(n9159), .ZN(P2_U3455) );
  MUX2_X1 U10556 ( .A(n9162), .B(n9161), .S(n10364), .Z(n9165) );
  NAND2_X1 U10557 ( .A1(n9163), .A2(n9204), .ZN(n9164) );
  OAI211_X1 U10558 ( .C1(n9166), .C2(n9212), .A(n9165), .B(n9164), .ZN(
        P2_U3454) );
  MUX2_X1 U10559 ( .A(n9168), .B(n9167), .S(n10364), .Z(n9169) );
  OAI21_X1 U10560 ( .B1(n9170), .B2(n9178), .A(n9169), .ZN(P2_U3453) );
  INV_X1 U10561 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9172) );
  MUX2_X1 U10562 ( .A(n9172), .B(n9171), .S(n10364), .Z(n9175) );
  NAND2_X1 U10563 ( .A1(n9173), .A2(n9204), .ZN(n9174) );
  OAI211_X1 U10564 ( .C1(n9176), .C2(n9212), .A(n9175), .B(n9174), .ZN(
        P2_U3452) );
  MUX2_X1 U10565 ( .A(n9177), .B(P2_REG0_REG_24__SCAN_IN), .S(n10366), .Z(
        n9182) );
  OAI22_X1 U10566 ( .A1(n9180), .A2(n9212), .B1(n9179), .B2(n9178), .ZN(n9181)
         );
  OR2_X1 U10567 ( .A1(n9182), .A2(n9181), .ZN(P2_U3451) );
  MUX2_X1 U10568 ( .A(n9184), .B(n9183), .S(n10364), .Z(n9187) );
  NAND2_X1 U10569 ( .A1(n9185), .A2(n9204), .ZN(n9186) );
  OAI211_X1 U10570 ( .C1(n9188), .C2(n9212), .A(n9187), .B(n9186), .ZN(
        P2_U3450) );
  MUX2_X1 U10571 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9189), .S(n10364), .Z(
        P2_U3449) );
  INV_X1 U10572 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9191) );
  MUX2_X1 U10573 ( .A(n9191), .B(n9190), .S(n10364), .Z(n9194) );
  NAND2_X1 U10574 ( .A1(n9192), .A2(n9204), .ZN(n9193) );
  OAI211_X1 U10575 ( .C1(n9195), .C2(n9212), .A(n9194), .B(n9193), .ZN(
        P2_U3448) );
  MUX2_X1 U10576 ( .A(n9197), .B(n9196), .S(n10364), .Z(n9200) );
  NAND2_X1 U10577 ( .A1(n9198), .A2(n9204), .ZN(n9199) );
  OAI211_X1 U10578 ( .C1(n9201), .C2(n9212), .A(n9200), .B(n9199), .ZN(
        P2_U3447) );
  INV_X1 U10579 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9203) );
  MUX2_X1 U10580 ( .A(n9203), .B(n9202), .S(n10364), .Z(n9207) );
  NAND2_X1 U10581 ( .A1(n9205), .A2(n9204), .ZN(n9206) );
  OAI211_X1 U10582 ( .C1(n9208), .C2(n9212), .A(n9207), .B(n9206), .ZN(
        P2_U3446) );
  MUX2_X1 U10583 ( .A(n9210), .B(n9209), .S(n10364), .Z(n9211) );
  OAI21_X1 U10584 ( .B1(n9213), .B2(n9212), .A(n9211), .ZN(P2_U3444) );
  INV_X1 U10585 ( .A(n9472), .ZN(n10174) );
  NOR4_X1 U10586 ( .A1(n9214), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n5314), .ZN(n9215) );
  AOI21_X1 U10587 ( .B1(n9216), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9215), .ZN(
        n9217) );
  OAI21_X1 U10588 ( .B1(n10174), .B2(n9220), .A(n9217), .ZN(P2_U3264) );
  OAI222_X1 U10589 ( .A1(n9222), .A2(n9221), .B1(n9220), .B2(n9219), .C1(
        P2_U3151), .C2(n9218), .ZN(P2_U3265) );
  INV_X1 U10590 ( .A(n9223), .ZN(n9224) );
  MUX2_X1 U10591 ( .A(n9224), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10592 ( .A(n9225), .ZN(n9230) );
  AOI21_X1 U10593 ( .B1(n9226), .B2(n9228), .A(n9227), .ZN(n9229) );
  OAI21_X1 U10594 ( .B1(n9230), .B2(n9229), .A(n9342), .ZN(n9234) );
  AOI22_X1 U10595 ( .A1(n9334), .A2(n9869), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n9233) );
  INV_X1 U10596 ( .A(n9845), .ZN(n9628) );
  AOI22_X1 U10597 ( .A1(n9357), .A2(n9847), .B1(n9355), .B2(n9628), .ZN(n9232)
         );
  NAND2_X1 U10598 ( .A1(n9846), .A2(n9363), .ZN(n9231) );
  NAND4_X1 U10599 ( .A1(n9234), .A2(n9233), .A3(n9232), .A4(n9231), .ZN(
        P1_U3214) );
  NAND2_X1 U10600 ( .A1(n9236), .A2(n9235), .ZN(n9238) );
  XNOR2_X1 U10601 ( .A(n9238), .B(n9237), .ZN(n9239) );
  NAND2_X1 U10602 ( .A1(n9239), .A2(n9342), .ZN(n9246) );
  NAND2_X1 U10603 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9709) );
  INV_X1 U10604 ( .A(n9709), .ZN(n9244) );
  INV_X1 U10605 ( .A(n9240), .ZN(n9242) );
  OAI22_X1 U10606 ( .A1(n9314), .A2(n9242), .B1(n9241), .B2(n9345), .ZN(n9243)
         );
  AOI211_X1 U10607 ( .C1(n9334), .C2(n9631), .A(n9244), .B(n9243), .ZN(n9245)
         );
  OAI211_X1 U10608 ( .C1(n9247), .C2(n9350), .A(n9246), .B(n9245), .ZN(
        P1_U3215) );
  XOR2_X1 U10609 ( .A(n9249), .B(n9248), .Z(n9253) );
  NAND2_X1 U10610 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9760) );
  OAI21_X1 U10611 ( .B1(n9941), .B2(n9345), .A(n9760), .ZN(n9251) );
  OAI22_X1 U10612 ( .A1(n9314), .A2(n9981), .B1(n10014), .B2(n9360), .ZN(n9250) );
  AOI211_X1 U10613 ( .C1(n9977), .C2(n9363), .A(n9251), .B(n9250), .ZN(n9252)
         );
  OAI21_X1 U10614 ( .B1(n9253), .B2(n9365), .A(n9252), .ZN(P1_U3219) );
  XNOR2_X1 U10615 ( .A(n9254), .B(n9255), .ZN(n9261) );
  OAI22_X1 U10616 ( .A1(n9941), .A2(n9360), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9256), .ZN(n9259) );
  INV_X1 U10617 ( .A(n9945), .ZN(n9257) );
  OAI22_X1 U10618 ( .A1(n9940), .A2(n9345), .B1(n9257), .B2(n9314), .ZN(n9258)
         );
  AOI211_X1 U10619 ( .C1(n9944), .C2(n9363), .A(n9259), .B(n9258), .ZN(n9260)
         );
  OAI21_X1 U10620 ( .B1(n9261), .B2(n9365), .A(n9260), .ZN(P1_U3223) );
  OAI21_X1 U10621 ( .B1(n9263), .B2(n9262), .A(n9339), .ZN(n9264) );
  NAND2_X1 U10622 ( .A1(n9264), .A2(n9342), .ZN(n9269) );
  OAI22_X1 U10623 ( .A1(n9345), .A2(n9842), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9265), .ZN(n9267) );
  OAI22_X1 U10624 ( .A1(n9443), .A2(n9360), .B1(n9879), .B2(n9314), .ZN(n9266)
         );
  AOI211_X1 U10625 ( .C1(n9877), .C2(n9363), .A(n9267), .B(n9266), .ZN(n9268)
         );
  NAND2_X1 U10626 ( .A1(n9269), .A2(n9268), .ZN(P1_U3225) );
  XNOR2_X1 U10627 ( .A(n9272), .B(n9271), .ZN(n9273) );
  XNOR2_X1 U10628 ( .A(n9270), .B(n9273), .ZN(n9279) );
  AOI22_X1 U10629 ( .A1(n9357), .A2(n9274), .B1(n9334), .B2(n9629), .ZN(n9276)
         );
  OAI211_X1 U10630 ( .C1(n9779), .C2(n9345), .A(n9276), .B(n9275), .ZN(n9277)
         );
  AOI21_X1 U10631 ( .B1(n10111), .B2(n9363), .A(n9277), .ZN(n9278) );
  OAI21_X1 U10632 ( .B1(n9279), .B2(n9365), .A(n9278), .ZN(P1_U3226) );
  NOR2_X1 U10633 ( .A1(n4584), .A2(n9281), .ZN(n9282) );
  XNOR2_X1 U10634 ( .A(n9283), .B(n9282), .ZN(n9288) );
  AOI22_X1 U10635 ( .A1(n9357), .A2(n10023), .B1(n9334), .B2(n9775), .ZN(n9285) );
  OAI211_X1 U10636 ( .C1(n10014), .C2(n9345), .A(n9285), .B(n9284), .ZN(n9286)
         );
  AOI21_X1 U10637 ( .B1(n10020), .B2(n9363), .A(n9286), .ZN(n9287) );
  OAI21_X1 U10638 ( .B1(n9288), .B2(n9365), .A(n9287), .ZN(P1_U3228) );
  INV_X1 U10639 ( .A(n9289), .ZN(n9291) );
  NOR3_X1 U10640 ( .A1(n4998), .A2(n9291), .A3(n9290), .ZN(n9294) );
  OAI21_X1 U10641 ( .B1(n9294), .B2(n4536), .A(n9342), .ZN(n9298) );
  AOI22_X1 U10642 ( .A1(n9891), .A2(n9334), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n9295) );
  OAI21_X1 U10643 ( .B1(n9897), .B2(n9314), .A(n9295), .ZN(n9296) );
  AOI21_X1 U10644 ( .B1(n9355), .B2(n9890), .A(n9296), .ZN(n9297) );
  OAI211_X1 U10645 ( .C1(n10145), .C2(n9350), .A(n9298), .B(n9297), .ZN(
        P1_U3229) );
  XNOR2_X1 U10646 ( .A(n9300), .B(n9299), .ZN(n9301) );
  XNOR2_X1 U10647 ( .A(n9302), .B(n9301), .ZN(n9308) );
  OAI22_X1 U10648 ( .A1(n9957), .A2(n9345), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9303), .ZN(n9306) );
  INV_X1 U10649 ( .A(n9963), .ZN(n9304) );
  OAI22_X1 U10650 ( .A1(n9314), .A2(n9304), .B1(n9956), .B2(n9360), .ZN(n9305)
         );
  AOI211_X1 U10651 ( .C1(n9962), .C2(n9363), .A(n9306), .B(n9305), .ZN(n9307)
         );
  OAI21_X1 U10652 ( .B1(n9308), .B2(n9365), .A(n9307), .ZN(P1_U3233) );
  XNOR2_X1 U10653 ( .A(n9310), .B(n9309), .ZN(n9311) );
  XNOR2_X1 U10654 ( .A(n9312), .B(n9311), .ZN(n9318) );
  OAI22_X1 U10655 ( .A1(n9957), .A2(n9360), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9313), .ZN(n9316) );
  OAI22_X1 U10656 ( .A1(n9924), .A2(n9345), .B1(n9314), .B2(n9927), .ZN(n9315)
         );
  AOI211_X1 U10657 ( .C1(n10079), .C2(n9363), .A(n9316), .B(n9315), .ZN(n9317)
         );
  OAI21_X1 U10658 ( .B1(n9318), .B2(n9365), .A(n9317), .ZN(P1_U3235) );
  INV_X1 U10659 ( .A(n9319), .ZN(n9324) );
  NOR3_X1 U10660 ( .A1(n9322), .A2(n9321), .A3(n9320), .ZN(n9323) );
  OAI21_X1 U10661 ( .B1(n9324), .B2(n9323), .A(n9342), .ZN(n9329) );
  AOI22_X1 U10662 ( .A1(n9334), .A2(n5593), .B1(n9325), .B2(n9363), .ZN(n9328)
         );
  AOI22_X1 U10663 ( .A1(P1_REG3_REG_2__SCAN_IN), .A2(n9326), .B1(n9355), .B2(
        n5739), .ZN(n9327) );
  NAND3_X1 U10664 ( .A1(n9329), .A2(n9328), .A3(n9327), .ZN(P1_U3237) );
  NAND2_X1 U10665 ( .A1(n9331), .A2(n9330), .ZN(n9333) );
  XNOR2_X1 U10666 ( .A(n9333), .B(n9332), .ZN(n9338) );
  AOI22_X1 U10667 ( .A1(n9357), .A2(n9991), .B1(n9334), .B2(n9998), .ZN(n9335)
         );
  NAND2_X1 U10668 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9724) );
  OAI211_X1 U10669 ( .C1(n9956), .C2(n9345), .A(n9335), .B(n9724), .ZN(n9336)
         );
  AOI21_X1 U10670 ( .B1(n10099), .B2(n9363), .A(n9336), .ZN(n9337) );
  OAI21_X1 U10671 ( .B1(n9338), .B2(n9365), .A(n9337), .ZN(P1_U3238) );
  NAND3_X1 U10672 ( .A1(n9343), .A2(n9342), .A3(n9226), .ZN(n9349) );
  OAI22_X1 U10673 ( .A1(n9345), .A2(n9859), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9344), .ZN(n9347) );
  INV_X1 U10674 ( .A(n9890), .ZN(n9858) );
  NOR2_X1 U10675 ( .A1(n9858), .A2(n9360), .ZN(n9346) );
  AOI211_X1 U10676 ( .C1(n9357), .C2(n9862), .A(n9347), .B(n9346), .ZN(n9348)
         );
  OAI211_X1 U10677 ( .C1(n4864), .C2(n9350), .A(n9349), .B(n9348), .ZN(
        P1_U3240) );
  XNOR2_X1 U10678 ( .A(n9353), .B(n9352), .ZN(n9354) );
  XNOR2_X1 U10679 ( .A(n9351), .B(n9354), .ZN(n9366) );
  AOI22_X1 U10680 ( .A1(n9357), .A2(n9356), .B1(n9355), .B2(n9775), .ZN(n9359)
         );
  OAI211_X1 U10681 ( .C1(n9361), .C2(n9360), .A(n9359), .B(n9358), .ZN(n9362)
         );
  AOI21_X1 U10682 ( .B1(n9418), .B2(n9363), .A(n9362), .ZN(n9364) );
  OAI21_X1 U10683 ( .B1(n9366), .B2(n9365), .A(n9364), .ZN(P1_U3241) );
  NAND2_X1 U10684 ( .A1(n9367), .A2(n9845), .ZN(n9483) );
  NAND2_X1 U10685 ( .A1(n9846), .A2(n9859), .ZN(n9484) );
  NAND2_X1 U10686 ( .A1(n9483), .A2(n9484), .ZN(n9528) );
  OAI21_X1 U10687 ( .B1(n9528), .B2(n9803), .A(n9804), .ZN(n9458) );
  NAND2_X1 U10688 ( .A1(n10058), .A2(n9842), .ZN(n9589) );
  INV_X1 U10689 ( .A(n9589), .ZN(n9839) );
  NOR3_X1 U10690 ( .A1(n9528), .A2(n9471), .A3(n9839), .ZN(n9368) );
  AOI21_X1 U10691 ( .B1(n9471), .B2(n9528), .A(n9368), .ZN(n9457) );
  INV_X1 U10692 ( .A(n9803), .ZN(n9369) );
  OR2_X1 U10693 ( .A1(n10058), .A2(n9842), .ZN(n9485) );
  OR2_X1 U10694 ( .A1(n9877), .A2(n9858), .ZN(n9800) );
  NAND2_X1 U10695 ( .A1(n9485), .A2(n9800), .ZN(n9519) );
  NOR3_X1 U10696 ( .A1(n9369), .A2(n4643), .A3(n9519), .ZN(n9451) );
  OR2_X1 U10697 ( .A1(n9944), .A2(n9957), .ZN(n9520) );
  NAND2_X1 U10698 ( .A1(n10155), .A2(n9972), .ZN(n9935) );
  AND2_X1 U10699 ( .A1(n9520), .A2(n9935), .ZN(n9588) );
  NAND2_X1 U10700 ( .A1(n9370), .A2(n9538), .ZN(n9372) );
  MUX2_X1 U10701 ( .A(n9372), .B(n9371), .S(n9471), .Z(n9376) );
  MUX2_X1 U10702 ( .A(n9534), .B(n9538), .S(n9471), .Z(n9373) );
  AND2_X1 U10703 ( .A1(n9373), .A2(n9494), .ZN(n9375) );
  INV_X1 U10704 ( .A(n9541), .ZN(n9374) );
  NAND2_X1 U10705 ( .A1(n9379), .A2(n9377), .ZN(n9540) );
  INV_X1 U10706 ( .A(n9540), .ZN(n9378) );
  INV_X1 U10707 ( .A(n9379), .ZN(n9380) );
  MUX2_X1 U10708 ( .A(n9384), .B(n9383), .S(n9471), .Z(n9385) );
  OAI21_X1 U10709 ( .B1(n9387), .B2(n9386), .A(n9385), .ZN(n9392) );
  MUX2_X1 U10710 ( .A(n9389), .B(n9388), .S(n4643), .Z(n9390) );
  INV_X1 U10711 ( .A(n9390), .ZN(n9391) );
  NAND2_X1 U10712 ( .A1(n9392), .A2(n9391), .ZN(n9397) );
  NAND2_X1 U10713 ( .A1(n9397), .A2(n9398), .ZN(n9393) );
  NAND2_X1 U10714 ( .A1(n9393), .A2(n9548), .ZN(n9394) );
  INV_X1 U10715 ( .A(n9554), .ZN(n9395) );
  NAND2_X1 U10716 ( .A1(n9397), .A2(n9396), .ZN(n9400) );
  NAND3_X1 U10717 ( .A1(n9400), .A2(n9399), .A3(n9398), .ZN(n9402) );
  AND2_X1 U10718 ( .A1(n9411), .A2(n9471), .ZN(n9408) );
  NAND3_X1 U10719 ( .A1(n9562), .A2(n9408), .A3(n9412), .ZN(n9406) );
  NAND3_X1 U10720 ( .A1(n9556), .A2(n4643), .A3(n9553), .ZN(n9405) );
  NAND2_X1 U10721 ( .A1(n9582), .A2(n9557), .ZN(n9407) );
  AND2_X1 U10722 ( .A1(n9407), .A2(n9562), .ZN(n9417) );
  NAND3_X1 U10723 ( .A1(n9412), .A2(n9408), .A3(n4848), .ZN(n9409) );
  OAI21_X1 U10724 ( .B1(n9556), .B2(n4643), .A(n9409), .ZN(n9410) );
  NAND2_X1 U10725 ( .A1(n9562), .A2(n9410), .ZN(n9415) );
  NAND2_X1 U10726 ( .A1(n9412), .A2(n9411), .ZN(n9559) );
  NAND3_X1 U10727 ( .A1(n9559), .A2(n4643), .A3(n9556), .ZN(n9413) );
  AND2_X1 U10728 ( .A1(n9561), .A2(n9413), .ZN(n9414) );
  OAI211_X1 U10729 ( .C1(n9562), .C2(n9471), .A(n9415), .B(n9414), .ZN(n9416)
         );
  NOR2_X1 U10730 ( .A1(n9417), .A2(n9416), .ZN(n9423) );
  INV_X1 U10731 ( .A(n9417), .ZN(n9421) );
  OR2_X1 U10732 ( .A1(n9418), .A2(n4643), .ZN(n9420) );
  NAND2_X1 U10733 ( .A1(n9582), .A2(n9629), .ZN(n9419) );
  AOI22_X1 U10734 ( .A1(n9421), .A2(n9420), .B1(n9471), .B2(n9419), .ZN(n9422)
         );
  AOI21_X1 U10735 ( .B1(n9424), .B2(n9423), .A(n9422), .ZN(n9425) );
  XNOR2_X1 U10736 ( .A(n10165), .B(n9998), .ZN(n10006) );
  OR2_X1 U10737 ( .A1(n9425), .A2(n10006), .ZN(n9433) );
  OR2_X1 U10738 ( .A1(n10099), .A2(n10014), .ZN(n9585) );
  OR2_X1 U10739 ( .A1(n10020), .A2(n9779), .ZN(n9583) );
  NAND2_X1 U10740 ( .A1(n9585), .A2(n9583), .ZN(n9563) );
  INV_X1 U10741 ( .A(n9563), .ZN(n9426) );
  NAND2_X1 U10742 ( .A1(n9433), .A2(n9426), .ZN(n9427) );
  NAND2_X1 U10743 ( .A1(n9977), .A2(n9956), .ZN(n9587) );
  NAND2_X1 U10744 ( .A1(n10099), .A2(n10014), .ZN(n9586) );
  NAND3_X1 U10745 ( .A1(n9427), .A2(n9587), .A3(n9586), .ZN(n9428) );
  OR2_X1 U10746 ( .A1(n9977), .A2(n9956), .ZN(n9487) );
  NAND3_X1 U10747 ( .A1(n9428), .A2(n9487), .A3(n9935), .ZN(n9430) );
  NAND2_X1 U10748 ( .A1(n9962), .A2(n9941), .ZN(n9434) );
  NAND2_X1 U10749 ( .A1(n9434), .A2(n9587), .ZN(n9429) );
  NAND2_X1 U10750 ( .A1(n10020), .A2(n9779), .ZN(n9584) );
  NAND2_X1 U10751 ( .A1(n9586), .A2(n9584), .ZN(n9566) );
  INV_X1 U10752 ( .A(n9566), .ZN(n9432) );
  AND2_X1 U10753 ( .A1(n9487), .A2(n9585), .ZN(n9565) );
  NAND2_X1 U10754 ( .A1(n9565), .A2(n4643), .ZN(n9431) );
  AOI21_X1 U10755 ( .B1(n9433), .B2(n9432), .A(n9431), .ZN(n9435) );
  NAND2_X1 U10756 ( .A1(n9944), .A2(n9957), .ZN(n9436) );
  NAND2_X1 U10757 ( .A1(n9436), .A2(n9434), .ZN(n9521) );
  XNOR2_X1 U10758 ( .A(n10079), .B(n9940), .ZN(n9921) );
  NAND2_X1 U10759 ( .A1(n10071), .A2(n9924), .ZN(n9889) );
  NAND2_X1 U10760 ( .A1(n10079), .A2(n9940), .ZN(n9522) );
  OAI211_X1 U10761 ( .C1(n9921), .C2(n9436), .A(n9889), .B(n9522), .ZN(n9437)
         );
  NAND2_X1 U10762 ( .A1(n9437), .A2(n4643), .ZN(n9438) );
  NAND2_X1 U10763 ( .A1(n9439), .A2(n9438), .ZN(n9440) );
  NAND2_X1 U10764 ( .A1(n9440), .A2(n9486), .ZN(n9442) );
  OR2_X1 U10765 ( .A1(n10079), .A2(n9940), .ZN(n9796) );
  NAND2_X1 U10766 ( .A1(n9486), .A2(n9796), .ZN(n9515) );
  NAND2_X1 U10767 ( .A1(n9515), .A2(n9471), .ZN(n9441) );
  NAND2_X1 U10768 ( .A1(n9442), .A2(n9441), .ZN(n9449) );
  OR2_X1 U10769 ( .A1(n9786), .A2(n9443), .ZN(n9799) );
  NAND2_X1 U10770 ( .A1(n9786), .A2(n9443), .ZN(n9523) );
  NAND2_X1 U10771 ( .A1(n9799), .A2(n9523), .ZN(n9887) );
  NOR2_X1 U10772 ( .A1(n9889), .A2(n4643), .ZN(n9444) );
  NOR2_X1 U10773 ( .A1(n9887), .A2(n9444), .ZN(n9448) );
  INV_X1 U10774 ( .A(n9523), .ZN(n9446) );
  INV_X1 U10775 ( .A(n9799), .ZN(n9445) );
  MUX2_X1 U10776 ( .A(n9446), .B(n9445), .S(n9471), .Z(n9447) );
  NOR2_X1 U10777 ( .A1(n10141), .A2(n9890), .ZN(n9452) );
  NAND2_X1 U10778 ( .A1(n9452), .A2(n9485), .ZN(n9526) );
  AOI21_X1 U10779 ( .B1(n9526), .B2(n9589), .A(n4643), .ZN(n9450) );
  AOI22_X1 U10780 ( .A1(n9451), .A2(n9454), .B1(n9450), .B2(n9803), .ZN(n9456)
         );
  INV_X1 U10781 ( .A(n9804), .ZN(n9455) );
  INV_X1 U10782 ( .A(n9452), .ZN(n9453) );
  NAND2_X1 U10783 ( .A1(n9459), .A2(n9467), .ZN(n9461) );
  NAND2_X1 U10784 ( .A1(n9473), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n9460) );
  NOR2_X1 U10785 ( .A1(n9814), .A2(n9820), .ZN(n9598) );
  NOR2_X1 U10786 ( .A1(n10042), .A2(n9462), .ZN(n9463) );
  NOR2_X1 U10787 ( .A1(n9598), .A2(n9463), .ZN(n9793) );
  INV_X1 U10788 ( .A(n9793), .ZN(n9805) );
  INV_X1 U10789 ( .A(n9463), .ZN(n9570) );
  INV_X1 U10790 ( .A(n9598), .ZN(n9464) );
  MUX2_X1 U10791 ( .A(n9570), .B(n9464), .S(n9471), .Z(n9465) );
  OAI21_X1 U10792 ( .B1(n9466), .B2(n9805), .A(n9465), .ZN(n9481) );
  NAND2_X1 U10793 ( .A1(n9468), .A2(n9467), .ZN(n9470) );
  NAND2_X1 U10794 ( .A1(n9473), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n9469) );
  NAND2_X1 U10795 ( .A1(n9472), .A2(n9467), .ZN(n9475) );
  NAND2_X1 U10796 ( .A1(n9473), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n9474) );
  NOR2_X1 U10797 ( .A1(n9766), .A2(n9482), .ZN(n9513) );
  INV_X1 U10798 ( .A(n9513), .ZN(n9622) );
  NAND2_X1 U10799 ( .A1(n9476), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n9480) );
  NAND2_X1 U10800 ( .A1(n9477), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9479) );
  NAND2_X1 U10801 ( .A1(n4492), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9478) );
  AND3_X1 U10802 ( .A1(n9480), .A2(n9479), .A3(n9478), .ZN(n9806) );
  INV_X1 U10803 ( .A(n9806), .ZN(n9627) );
  NAND2_X1 U10804 ( .A1(n9627), .A2(n9765), .ZN(n9597) );
  AND2_X1 U10805 ( .A1(n9766), .A2(n9482), .ZN(n9574) );
  INV_X1 U10806 ( .A(n5280), .ZN(n9615) );
  AOI21_X1 U10807 ( .B1(n9616), .B2(n9615), .A(n5514), .ZN(n9626) );
  NAND2_X1 U10808 ( .A1(n4661), .A2(n9627), .ZN(n9572) );
  INV_X1 U10809 ( .A(n9572), .ZN(n9512) );
  INV_X1 U10810 ( .A(n9824), .ZN(n9511) );
  NAND2_X1 U10811 ( .A1(n9485), .A2(n9589), .ZN(n9856) );
  NAND2_X1 U10812 ( .A1(n9486), .A2(n9889), .ZN(n9909) );
  XNOR2_X1 U10813 ( .A(n10151), .B(n9957), .ZN(n9936) );
  INV_X1 U10814 ( .A(n9777), .ZN(n9580) );
  INV_X1 U10815 ( .A(n9488), .ZN(n9504) );
  NOR4_X1 U10816 ( .A1(n9491), .A2(n9490), .A3(n9489), .A4(n9531), .ZN(n9495)
         );
  NAND4_X1 U10817 ( .A1(n9495), .A2(n9494), .A3(n9493), .A4(n9492), .ZN(n9496)
         );
  OR4_X1 U10818 ( .A1(n9544), .A2(n9498), .A3(n9497), .A4(n9496), .ZN(n9499)
         );
  NOR4_X1 U10819 ( .A1(n9502), .A2(n9501), .A3(n9500), .A4(n9499), .ZN(n9503)
         );
  NAND4_X1 U10820 ( .A1(n9580), .A2(n9505), .A3(n9504), .A4(n9503), .ZN(n9506)
         );
  NOR3_X1 U10821 ( .A1(n9563), .A2(n9566), .A3(n9506), .ZN(n9507) );
  XNOR2_X1 U10822 ( .A(n10155), .B(n9941), .ZN(n9953) );
  NAND4_X1 U10823 ( .A1(n9936), .A2(n9975), .A3(n9507), .A4(n9953), .ZN(n9508)
         );
  NOR4_X1 U10824 ( .A1(n9887), .A2(n9909), .A3(n9921), .A4(n9508), .ZN(n9509)
         );
  XNOR2_X1 U10825 ( .A(n9877), .B(n9890), .ZN(n9873) );
  NAND4_X1 U10826 ( .A1(n9836), .A2(n9801), .A3(n9509), .A4(n9873), .ZN(n9510)
         );
  NOR4_X1 U10827 ( .A1(n9805), .A2(n9512), .A3(n9511), .A4(n9510), .ZN(n9514)
         );
  AOI21_X1 U10828 ( .B1(n9806), .B2(n9596), .A(n9513), .ZN(n9576) );
  NAND3_X1 U10829 ( .A1(n9514), .A2(n9576), .A3(n9614), .ZN(n9607) );
  NAND4_X1 U10830 ( .A1(n9607), .A2(n9604), .A3(n5281), .A4(n9610), .ZN(n9625)
         );
  NAND2_X1 U10831 ( .A1(n9515), .A2(n9889), .ZN(n9516) );
  NAND2_X1 U10832 ( .A1(n9799), .A2(n9516), .ZN(n9517) );
  AND2_X1 U10833 ( .A1(n9517), .A2(n9523), .ZN(n9518) );
  OR2_X1 U10834 ( .A1(n9519), .A2(n9518), .ZN(n9590) );
  INV_X1 U10835 ( .A(n9590), .ZN(n9525) );
  NAND2_X1 U10836 ( .A1(n9521), .A2(n9520), .ZN(n9794) );
  NAND4_X1 U10837 ( .A1(n9523), .A2(n9889), .A3(n9522), .A4(n9794), .ZN(n9524)
         );
  NAND2_X1 U10838 ( .A1(n9525), .A2(n9524), .ZN(n9527) );
  NAND2_X1 U10839 ( .A1(n9527), .A2(n9526), .ZN(n9529) );
  AOI21_X1 U10840 ( .B1(n9803), .B2(n9529), .A(n9528), .ZN(n9591) );
  NAND2_X1 U10841 ( .A1(n5594), .A2(n9530), .ZN(n9533) );
  NAND2_X1 U10842 ( .A1(n5593), .A2(n5597), .ZN(n9532) );
  AND3_X1 U10843 ( .A1(n9533), .A2(n9532), .A3(n9531), .ZN(n9536) );
  OAI211_X1 U10844 ( .C1(n9537), .C2(n9536), .A(n9535), .B(n9534), .ZN(n9539)
         );
  NAND2_X1 U10845 ( .A1(n9539), .A2(n9538), .ZN(n9542) );
  AOI21_X1 U10846 ( .B1(n9542), .B2(n9541), .A(n9540), .ZN(n9546) );
  INV_X1 U10847 ( .A(n9544), .ZN(n9545) );
  OAI21_X1 U10848 ( .B1(n9546), .B2(n4684), .A(n9545), .ZN(n9549) );
  NAND4_X1 U10849 ( .A1(n9549), .A2(n9551), .A3(n9548), .A4(n9547), .ZN(n9555)
         );
  NAND2_X1 U10850 ( .A1(n9551), .A2(n4642), .ZN(n9552) );
  AND4_X1 U10851 ( .A1(n9555), .A2(n9554), .A3(n9553), .A4(n9552), .ZN(n9558)
         );
  OAI211_X1 U10852 ( .C1(n9559), .C2(n9558), .A(n9557), .B(n9556), .ZN(n9560)
         );
  NAND3_X1 U10853 ( .A1(n9562), .A2(n9561), .A3(n9560), .ZN(n9564) );
  AOI21_X1 U10854 ( .B1(n9582), .B2(n9564), .A(n9563), .ZN(n9567) );
  OAI21_X1 U10855 ( .B1(n9567), .B2(n9566), .A(n9565), .ZN(n9568) );
  AOI211_X1 U10856 ( .C1(n9587), .C2(n9568), .A(n4828), .B(n9590), .ZN(n9569)
         );
  OAI21_X1 U10857 ( .B1(n9569), .B2(n9839), .A(n9803), .ZN(n9571) );
  NAND2_X1 U10858 ( .A1(n9570), .A2(n9804), .ZN(n9595) );
  AOI21_X1 U10859 ( .B1(n9591), .B2(n9571), .A(n9595), .ZN(n9573) );
  OAI21_X1 U10860 ( .B1(n9573), .B2(n9598), .A(n9572), .ZN(n9575) );
  AOI21_X1 U10861 ( .B1(n9576), .B2(n9575), .A(n9574), .ZN(n9579) );
  AOI21_X1 U10862 ( .B1(n5281), .B2(n9577), .A(n9579), .ZN(n9578) );
  AOI211_X1 U10863 ( .C1(n9579), .C2(n5516), .A(n9618), .B(n9578), .ZN(n9613)
         );
  INV_X1 U10864 ( .A(n9597), .ZN(n9601) );
  NAND2_X1 U10865 ( .A1(n9995), .A2(n9996), .ZN(n9994) );
  NAND2_X1 U10866 ( .A1(n9994), .A2(n9586), .ZN(n9970) );
  NAND2_X1 U10867 ( .A1(n9970), .A2(n9975), .ZN(n9969) );
  OAI21_X1 U10868 ( .B1(n9590), .B2(n9795), .A(n9589), .ZN(n9593) );
  INV_X1 U10869 ( .A(n9591), .ZN(n9592) );
  AOI21_X1 U10870 ( .B1(n9803), .B2(n9593), .A(n9592), .ZN(n9594) );
  NOR2_X1 U10871 ( .A1(n9595), .A2(n9594), .ZN(n9599) );
  OAI22_X1 U10872 ( .A1(n9599), .A2(n9598), .B1(n9597), .B2(n9596), .ZN(n9600)
         );
  OAI211_X1 U10873 ( .C1(n4661), .C2(n9601), .A(n9600), .B(n9622), .ZN(n9603)
         );
  NAND3_X1 U10874 ( .A1(n9603), .A2(n9602), .A3(n9614), .ZN(n9606) );
  NAND2_X1 U10875 ( .A1(n9604), .A2(n9621), .ZN(n9605) );
  AOI211_X1 U10876 ( .C1(n9607), .C2(n9606), .A(n9618), .B(n9605), .ZN(n9612)
         );
  INV_X1 U10877 ( .A(P1_B_REG_SCAN_IN), .ZN(n9609) );
  NOR4_X1 U10878 ( .A1(n10011), .A2(n10239), .A3(n5175), .A4(n5516), .ZN(n9608) );
  AOI211_X1 U10879 ( .C1(n9610), .C2(n5280), .A(n9609), .B(n9608), .ZN(n9611)
         );
  NOR3_X1 U10880 ( .A1(n9613), .A2(n9612), .A3(n9611), .ZN(n9624) );
  NOR2_X1 U10881 ( .A1(n9618), .A2(n9617), .ZN(n9619) );
  OAI211_X1 U10882 ( .C1(n9622), .C2(n9621), .A(n9620), .B(n9619), .ZN(n9623)
         );
  OAI211_X1 U10883 ( .C1(n9626), .C2(n9625), .A(n9624), .B(n9623), .ZN(
        P1_U3242) );
  MUX2_X1 U10884 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9627), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10885 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9820), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10886 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9628), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10887 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9821), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10888 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9869), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10889 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9890), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10890 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9913), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10891 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9891), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10892 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9914), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10893 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9784), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10894 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9972), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10895 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n10000), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10896 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9971), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10897 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9998), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10898 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9775), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10899 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9629), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10900 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9630), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10901 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9631), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10902 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9632), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10903 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9633), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10904 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9634), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10905 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n4836), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10906 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9635), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10907 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9636), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10908 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9637), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10909 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9638), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10910 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n5742), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10911 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n5739), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10912 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n5735), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10913 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n5593), .S(P1_U3973), .Z(
        P1_U3555) );
  MUX2_X1 U10914 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n5594), .S(P1_U3973), .Z(
        P1_U3554) );
  OAI211_X1 U10915 ( .C1(n9651), .C2(n9640), .A(n9740), .B(n9639), .ZN(n9649)
         );
  OAI211_X1 U10916 ( .C1(n9643), .C2(n9642), .A(n9756), .B(n9641), .ZN(n9648)
         );
  AOI22_X1 U10917 ( .A1(n9644), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9647) );
  NAND2_X1 U10918 ( .A1(n9755), .A2(n9645), .ZN(n9646) );
  NAND4_X1 U10919 ( .A1(n9649), .A2(n9648), .A3(n9647), .A4(n9646), .ZN(
        P1_U3244) );
  MUX2_X1 U10920 ( .A(n9651), .B(n9650), .S(n5175), .Z(n9653) );
  NAND2_X1 U10921 ( .A1(n9653), .A2(n9652), .ZN(n9654) );
  OAI211_X1 U10922 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n9655), .A(n9654), .B(
        P1_U3973), .ZN(n9695) );
  OAI22_X1 U10923 ( .A1(n9761), .A2(n8966), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9656), .ZN(n9657) );
  AOI21_X1 U10924 ( .B1(n9755), .B2(n9658), .A(n9657), .ZN(n9667) );
  OAI211_X1 U10925 ( .C1(n9661), .C2(n9660), .A(n9756), .B(n9659), .ZN(n9666)
         );
  OAI211_X1 U10926 ( .C1(n9664), .C2(n9663), .A(n9740), .B(n9662), .ZN(n9665)
         );
  NAND4_X1 U10927 ( .A1(n9695), .A2(n9667), .A3(n9666), .A4(n9665), .ZN(
        P1_U3245) );
  INV_X1 U10928 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9669) );
  OAI21_X1 U10929 ( .B1(n9761), .B2(n9669), .A(n9668), .ZN(n9670) );
  AOI21_X1 U10930 ( .B1(n9755), .B2(n9671), .A(n9670), .ZN(n9680) );
  OAI211_X1 U10931 ( .C1(n9674), .C2(n9673), .A(n9756), .B(n9672), .ZN(n9679)
         );
  OAI211_X1 U10932 ( .C1(n9677), .C2(n9676), .A(n9740), .B(n9675), .ZN(n9678)
         );
  NAND3_X1 U10933 ( .A1(n9680), .A2(n9679), .A3(n9678), .ZN(P1_U3246) );
  INV_X1 U10934 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9683) );
  INV_X1 U10935 ( .A(n9681), .ZN(n9682) );
  OAI21_X1 U10936 ( .B1(n9761), .B2(n9683), .A(n9682), .ZN(n9684) );
  AOI21_X1 U10937 ( .B1(n9755), .B2(n9685), .A(n9684), .ZN(n9694) );
  OAI211_X1 U10938 ( .C1(n9688), .C2(n9687), .A(n9740), .B(n9686), .ZN(n9693)
         );
  OAI211_X1 U10939 ( .C1(n9691), .C2(n9690), .A(n9756), .B(n9689), .ZN(n9692)
         );
  NAND4_X1 U10940 ( .A1(n9695), .A2(n9694), .A3(n9693), .A4(n9692), .ZN(
        P1_U3247) );
  INV_X1 U10941 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9697) );
  OAI21_X1 U10942 ( .B1(n9761), .B2(n9697), .A(n9696), .ZN(n9698) );
  AOI21_X1 U10943 ( .B1(n9755), .B2(n9699), .A(n9698), .ZN(n9708) );
  OAI211_X1 U10944 ( .C1(n9702), .C2(n9701), .A(n9740), .B(n9700), .ZN(n9707)
         );
  OAI211_X1 U10945 ( .C1(n9705), .C2(n9704), .A(n9756), .B(n9703), .ZN(n9706)
         );
  NAND3_X1 U10946 ( .A1(n9708), .A2(n9707), .A3(n9706), .ZN(P1_U3256) );
  INV_X1 U10947 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9710) );
  OAI21_X1 U10948 ( .B1(n9761), .B2(n9710), .A(n9709), .ZN(n9711) );
  AOI21_X1 U10949 ( .B1(n9755), .B2(n9712), .A(n9711), .ZN(n9723) );
  INV_X1 U10950 ( .A(n9713), .ZN(n9714) );
  OAI211_X1 U10951 ( .C1(n9716), .C2(n9715), .A(n9756), .B(n9714), .ZN(n9722)
         );
  INV_X1 U10952 ( .A(n9717), .ZN(n9718) );
  OAI211_X1 U10953 ( .C1(n9720), .C2(n9719), .A(n9740), .B(n9718), .ZN(n9721)
         );
  NAND3_X1 U10954 ( .A1(n9723), .A2(n9722), .A3(n9721), .ZN(P1_U3257) );
  OAI21_X1 U10955 ( .B1(n9761), .B2(n10388), .A(n9724), .ZN(n9734) );
  NAND2_X1 U10956 ( .A1(n9738), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9748) );
  OR2_X1 U10957 ( .A1(n9738), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9725) );
  NAND2_X1 U10958 ( .A1(n9748), .A2(n9725), .ZN(n9732) );
  NAND2_X1 U10959 ( .A1(n9727), .A2(n9726), .ZN(n9729) );
  OR2_X1 U10960 ( .A1(n9735), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9728) );
  NAND2_X1 U10961 ( .A1(n9729), .A2(n9728), .ZN(n9731) );
  INV_X1 U10962 ( .A(n9749), .ZN(n9730) );
  AOI211_X1 U10963 ( .C1(n9732), .C2(n9731), .A(n9751), .B(n9730), .ZN(n9733)
         );
  AOI211_X1 U10964 ( .C1(n9755), .C2(n9738), .A(n9734), .B(n9733), .ZN(n9744)
         );
  OR2_X1 U10965 ( .A1(n9735), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9736) );
  AND2_X1 U10966 ( .A1(n9737), .A2(n9736), .ZN(n9742) );
  NAND2_X1 U10967 ( .A1(n9738), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9745) );
  OR2_X1 U10968 ( .A1(n9738), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9739) );
  AND2_X1 U10969 ( .A1(n9745), .A2(n9739), .ZN(n9741) );
  NAND2_X1 U10970 ( .A1(n9742), .A2(n9741), .ZN(n9746) );
  OAI211_X1 U10971 ( .C1(n9742), .C2(n9741), .A(n9746), .B(n9740), .ZN(n9743)
         );
  NAND2_X1 U10972 ( .A1(n9744), .A2(n9743), .ZN(P1_U3261) );
  NAND2_X1 U10973 ( .A1(n9746), .A2(n9745), .ZN(n9747) );
  XNOR2_X1 U10974 ( .A(n9747), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9754) );
  NAND2_X1 U10975 ( .A1(n9749), .A2(n9748), .ZN(n9750) );
  XNOR2_X1 U10976 ( .A(n9750), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9757) );
  NAND3_X1 U10977 ( .A1(n9754), .A2(n9762), .A3(n9753), .ZN(n9759) );
  AOI21_X1 U10978 ( .B1(n9757), .B2(n9756), .A(n9755), .ZN(n9758) );
  NOR2_X4 U10979 ( .A1(n10019), .A2(n10020), .ZN(n10018) );
  OR2_X2 U10980 ( .A1(n10079), .A2(n9942), .ZN(n9925) );
  NOR2_X2 U10981 ( .A1(n10042), .A2(n9828), .ZN(n9810) );
  NAND2_X1 U10982 ( .A1(n4661), .A2(n9810), .ZN(n9770) );
  XNOR2_X1 U10983 ( .A(n9770), .B(n9766), .ZN(n10032) );
  NAND2_X1 U10984 ( .A1(n9762), .A2(P1_B_REG_SCAN_IN), .ZN(n9763) );
  NAND2_X1 U10985 ( .A1(n9999), .A2(n9763), .ZN(n9807) );
  INV_X1 U10986 ( .A(n9807), .ZN(n9764) );
  NAND2_X1 U10987 ( .A1(n9765), .A2(n9764), .ZN(n10035) );
  NOR2_X1 U10988 ( .A1(n9986), .A2(n10035), .ZN(n9772) );
  NOR2_X1 U10989 ( .A1(n10125), .A2(n10026), .ZN(n9767) );
  AOI211_X1 U10990 ( .C1(n9986), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9772), .B(
        n9767), .ZN(n9768) );
  OAI21_X1 U10991 ( .B1(n10032), .B2(n9769), .A(n9768), .ZN(P1_U3263) );
  OAI211_X1 U10992 ( .C1(n4661), .C2(n9810), .A(n10072), .B(n9770), .ZN(n10036) );
  NOR2_X1 U10993 ( .A1(n4661), .A2(n10026), .ZN(n9771) );
  AOI211_X1 U10994 ( .C1(n9986), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9772), .B(
        n9771), .ZN(n9773) );
  OAI21_X1 U10995 ( .B1(n9774), .B2(n10036), .A(n9773), .ZN(P1_U3264) );
  AOI21_X1 U10996 ( .B1(n9778), .B2(n9777), .A(n9776), .ZN(n10005) );
  AOI21_X1 U10997 ( .B1(n9941), .B2(n10155), .A(n9952), .ZN(n9783) );
  NAND2_X1 U10998 ( .A1(n10079), .A2(n9914), .ZN(n9785) );
  NAND2_X1 U10999 ( .A1(n9877), .A2(n9890), .ZN(n9787) );
  NAND2_X1 U11000 ( .A1(n9788), .A2(n9787), .ZN(n9853) );
  NAND2_X1 U11001 ( .A1(n9853), .A2(n9856), .ZN(n9790) );
  NAND2_X1 U11002 ( .A1(n10058), .A2(n9869), .ZN(n9789) );
  NAND2_X1 U11003 ( .A1(n9790), .A2(n9789), .ZN(n9835) );
  NAND2_X1 U11004 ( .A1(n4863), .A2(n9859), .ZN(n9791) );
  INV_X1 U11005 ( .A(n10039), .ZN(n9817) );
  OR2_X1 U11006 ( .A1(n9908), .A2(n9909), .ZN(n9910) );
  INV_X1 U11007 ( .A(n9889), .ZN(n9797) );
  NOR2_X1 U11008 ( .A1(n9887), .A2(n9797), .ZN(n9798) );
  NAND2_X1 U11009 ( .A1(n9910), .A2(n9798), .ZN(n9886) );
  NAND2_X1 U11010 ( .A1(n9886), .A2(n9799), .ZN(n9868) );
  INV_X1 U11011 ( .A(n9836), .ZN(n9838) );
  NOR2_X1 U11012 ( .A1(n9838), .A2(n9839), .ZN(n9802) );
  NAND2_X1 U11013 ( .A1(n9837), .A2(n9802), .ZN(n9840) );
  NAND2_X1 U11014 ( .A1(n9840), .A2(n9803), .ZN(n9819) );
  NAND2_X1 U11015 ( .A1(n9819), .A2(n9824), .ZN(n9818) );
  INV_X1 U11016 ( .A(n9808), .ZN(n9809) );
  AOI211_X1 U11017 ( .C1(n10042), .C2(n9828), .A(n10266), .B(n9810), .ZN(
        n10041) );
  NAND2_X1 U11018 ( .A1(n10041), .A2(n10021), .ZN(n9813) );
  AOI22_X1 U11019 ( .A1(n9986), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n10022), 
        .B2(n9811), .ZN(n9812) );
  OAI211_X1 U11020 ( .C1(n9814), .C2(n10026), .A(n9813), .B(n9812), .ZN(n9815)
         );
  AOI21_X1 U11021 ( .B1(n10040), .B2(n10028), .A(n9815), .ZN(n9816) );
  OAI21_X1 U11022 ( .B1(n9817), .B2(n10030), .A(n9816), .ZN(P1_U3356) );
  OAI211_X1 U11023 ( .C1(n9819), .C2(n9824), .A(n9818), .B(n10009), .ZN(n9823)
         );
  AOI22_X1 U11024 ( .A1(n9821), .A2(n9997), .B1(n9999), .B2(n9820), .ZN(n9822)
         );
  AND2_X1 U11025 ( .A1(n9823), .A2(n9822), .ZN(n10046) );
  NAND2_X1 U11026 ( .A1(n9825), .A2(n9824), .ZN(n9826) );
  NAND2_X1 U11027 ( .A1(n10048), .A2(n9976), .ZN(n9834) );
  OAI211_X1 U11028 ( .C1(n10133), .C2(n4505), .A(n10072), .B(n9828), .ZN(
        n10045) );
  INV_X1 U11029 ( .A(n10045), .ZN(n9832) );
  AOI22_X1 U11030 ( .A1(n9986), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9829), .B2(
        n10022), .ZN(n9830) );
  OAI21_X1 U11031 ( .B1(n10133), .B2(n10026), .A(n9830), .ZN(n9831) );
  AOI21_X1 U11032 ( .B1(n9832), .B2(n10021), .A(n9831), .ZN(n9833) );
  OAI211_X1 U11033 ( .C1(n10046), .C2(n9986), .A(n9834), .B(n9833), .ZN(
        P1_U3265) );
  XNOR2_X1 U11034 ( .A(n9835), .B(n9836), .ZN(n10053) );
  INV_X1 U11035 ( .A(n10053), .ZN(n9852) );
  INV_X1 U11036 ( .A(n9837), .ZN(n9854) );
  OAI21_X1 U11037 ( .B1(n9854), .B2(n9839), .A(n9838), .ZN(n9841) );
  NAND3_X1 U11038 ( .A1(n9841), .A2(n10009), .A3(n9840), .ZN(n9844) );
  OR2_X1 U11039 ( .A1(n9842), .A2(n10011), .ZN(n9843) );
  OAI211_X1 U11040 ( .C1(n9845), .C2(n10013), .A(n9844), .B(n9843), .ZN(n10051) );
  AOI211_X1 U11041 ( .C1(n9846), .C2(n9860), .A(n10266), .B(n4505), .ZN(n10052) );
  NAND2_X1 U11042 ( .A1(n10052), .A2(n10021), .ZN(n9849) );
  AOI22_X1 U11043 ( .A1(n9986), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n10022), 
        .B2(n9847), .ZN(n9848) );
  OAI211_X1 U11044 ( .C1(n4863), .C2(n10026), .A(n9849), .B(n9848), .ZN(n9850)
         );
  AOI21_X1 U11045 ( .B1(n10051), .B2(n10028), .A(n9850), .ZN(n9851) );
  OAI21_X1 U11046 ( .B1(n9852), .B2(n10030), .A(n9851), .ZN(P1_U3266) );
  XNOR2_X1 U11047 ( .A(n9853), .B(n9856), .ZN(n10060) );
  AOI21_X1 U11048 ( .B1(n9856), .B2(n9855), .A(n9854), .ZN(n9857) );
  OAI222_X1 U11049 ( .A1(n10013), .A2(n9859), .B1(n10011), .B2(n9858), .C1(
        n9938), .C2(n9857), .ZN(n10056) );
  INV_X1 U11050 ( .A(n9860), .ZN(n9861) );
  AOI211_X1 U11051 ( .C1(n10058), .C2(n9874), .A(n10266), .B(n9861), .ZN(
        n10057) );
  NAND2_X1 U11052 ( .A1(n10057), .A2(n10021), .ZN(n9864) );
  AOI22_X1 U11053 ( .A1(n9986), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9862), .B2(
        n10022), .ZN(n9863) );
  OAI211_X1 U11054 ( .C1(n4864), .C2(n10026), .A(n9864), .B(n9863), .ZN(n9865)
         );
  AOI21_X1 U11055 ( .B1(n10056), .B2(n10028), .A(n9865), .ZN(n9866) );
  OAI21_X1 U11056 ( .B1(n10060), .B2(n10030), .A(n9866), .ZN(P1_U3267) );
  OAI211_X1 U11057 ( .C1(n9868), .C2(n9873), .A(n9867), .B(n10009), .ZN(n9871)
         );
  AOI22_X1 U11058 ( .A1(n9913), .A2(n9997), .B1(n9999), .B2(n9869), .ZN(n9870)
         );
  NAND2_X1 U11059 ( .A1(n9871), .A2(n9870), .ZN(n10061) );
  INV_X1 U11060 ( .A(n10061), .ZN(n9884) );
  XNOR2_X1 U11061 ( .A(n9872), .B(n9873), .ZN(n10063) );
  NAND2_X1 U11062 ( .A1(n10063), .A2(n9976), .ZN(n9883) );
  INV_X1 U11063 ( .A(n9895), .ZN(n9876) );
  INV_X1 U11064 ( .A(n9874), .ZN(n9875) );
  AOI211_X1 U11065 ( .C1(n9877), .C2(n9876), .A(n10266), .B(n9875), .ZN(n10062) );
  NOR2_X1 U11066 ( .A1(n10141), .A2(n10026), .ZN(n9881) );
  INV_X1 U11067 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9878) );
  OAI22_X1 U11068 ( .A1(n9879), .A2(n9980), .B1(n9878), .B2(n10028), .ZN(n9880) );
  AOI211_X1 U11069 ( .C1(n10062), .C2(n10021), .A(n9881), .B(n9880), .ZN(n9882) );
  OAI211_X1 U11070 ( .C1(n9986), .C2(n9884), .A(n9883), .B(n9882), .ZN(
        P1_U3268) );
  XNOR2_X1 U11071 ( .A(n9885), .B(n9887), .ZN(n10068) );
  INV_X1 U11072 ( .A(n10068), .ZN(n9903) );
  NAND2_X1 U11073 ( .A1(n9886), .A2(n10009), .ZN(n9894) );
  INV_X1 U11074 ( .A(n9887), .ZN(n9888) );
  AOI21_X1 U11075 ( .B1(n9910), .B2(n9889), .A(n9888), .ZN(n9893) );
  AOI22_X1 U11076 ( .A1(n9891), .A2(n9997), .B1(n9890), .B2(n9999), .ZN(n9892)
         );
  OAI21_X1 U11077 ( .B1(n9894), .B2(n9893), .A(n9892), .ZN(n10066) );
  OAI21_X1 U11078 ( .B1(n10145), .B2(n9904), .A(n10072), .ZN(n9896) );
  NOR2_X1 U11079 ( .A1(n9896), .A2(n9895), .ZN(n10067) );
  NAND2_X1 U11080 ( .A1(n10067), .A2(n10021), .ZN(n9900) );
  INV_X1 U11081 ( .A(n9897), .ZN(n9898) );
  AOI22_X1 U11082 ( .A1(n9898), .A2(n10022), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n9986), .ZN(n9899) );
  OAI211_X1 U11083 ( .C1(n10145), .C2(n10026), .A(n9900), .B(n9899), .ZN(n9901) );
  AOI21_X1 U11084 ( .B1(n10066), .B2(n10028), .A(n9901), .ZN(n9902) );
  OAI21_X1 U11085 ( .B1(n9903), .B2(n10030), .A(n9902), .ZN(P1_U3269) );
  XNOR2_X1 U11086 ( .A(n4547), .B(n9909), .ZN(n10076) );
  AOI21_X1 U11087 ( .B1(n10071), .B2(n9925), .A(n9904), .ZN(n10073) );
  AOI22_X1 U11088 ( .A1(n9905), .A2(n10022), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n9986), .ZN(n9906) );
  OAI21_X1 U11089 ( .B1(n9907), .B2(n10026), .A(n9906), .ZN(n9917) );
  INV_X1 U11090 ( .A(n9908), .ZN(n9912) );
  INV_X1 U11091 ( .A(n9909), .ZN(n9911) );
  OAI21_X1 U11092 ( .B1(n9912), .B2(n9911), .A(n9910), .ZN(n9915) );
  AOI222_X1 U11093 ( .A1(n10009), .A2(n9915), .B1(n9914), .B2(n9997), .C1(
        n9913), .C2(n9999), .ZN(n10075) );
  NOR2_X1 U11094 ( .A1(n10075), .A2(n9986), .ZN(n9916) );
  AOI211_X1 U11095 ( .C1(n10073), .C2(n9918), .A(n9917), .B(n9916), .ZN(n9919)
         );
  OAI21_X1 U11096 ( .B1(n10076), .B2(n10030), .A(n9919), .ZN(P1_U3270) );
  XNOR2_X1 U11097 ( .A(n9920), .B(n4823), .ZN(n10081) );
  XNOR2_X1 U11098 ( .A(n9922), .B(n9921), .ZN(n9923) );
  OAI222_X1 U11099 ( .A1(n10013), .A2(n9924), .B1(n10011), .B2(n9957), .C1(
        n9938), .C2(n9923), .ZN(n10077) );
  INV_X1 U11100 ( .A(n9925), .ZN(n9926) );
  AOI211_X1 U11101 ( .C1(n10079), .C2(n9942), .A(n10266), .B(n9926), .ZN(
        n10078) );
  NAND2_X1 U11102 ( .A1(n10078), .A2(n10021), .ZN(n9930) );
  INV_X1 U11103 ( .A(n9927), .ZN(n9928) );
  AOI22_X1 U11104 ( .A1(n9928), .A2(n10022), .B1(n9986), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n9929) );
  OAI211_X1 U11105 ( .C1(n9931), .C2(n10026), .A(n9930), .B(n9929), .ZN(n9932)
         );
  AOI21_X1 U11106 ( .B1(n10077), .B2(n10028), .A(n9932), .ZN(n9933) );
  OAI21_X1 U11107 ( .B1(n10081), .B2(n10030), .A(n9933), .ZN(P1_U3271) );
  XOR2_X1 U11108 ( .A(n9934), .B(n9936), .Z(n10084) );
  INV_X1 U11109 ( .A(n10084), .ZN(n9950) );
  INV_X1 U11110 ( .A(n9953), .ZN(n9951) );
  OAI21_X1 U11111 ( .B1(n9954), .B2(n9951), .A(n9935), .ZN(n9937) );
  XNOR2_X1 U11112 ( .A(n9937), .B(n9936), .ZN(n9939) );
  OAI222_X1 U11113 ( .A1(n10011), .A2(n9941), .B1(n10013), .B2(n9940), .C1(
        n9939), .C2(n9938), .ZN(n10082) );
  INV_X1 U11114 ( .A(n9942), .ZN(n9943) );
  AOI211_X1 U11115 ( .C1(n9944), .C2(n4860), .A(n10266), .B(n9943), .ZN(n10083) );
  NAND2_X1 U11116 ( .A1(n10083), .A2(n10021), .ZN(n9947) );
  AOI22_X1 U11117 ( .A1(n9986), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9945), .B2(
        n10022), .ZN(n9946) );
  OAI211_X1 U11118 ( .C1(n10151), .C2(n10026), .A(n9947), .B(n9946), .ZN(n9948) );
  AOI21_X1 U11119 ( .B1(n10082), .B2(n10028), .A(n9948), .ZN(n9949) );
  OAI21_X1 U11120 ( .B1(n9950), .B2(n10030), .A(n9949), .ZN(P1_U3272) );
  XNOR2_X1 U11121 ( .A(n9952), .B(n9951), .ZN(n10089) );
  INV_X1 U11122 ( .A(n10089), .ZN(n9968) );
  XNOR2_X1 U11123 ( .A(n9954), .B(n9953), .ZN(n9955) );
  NAND2_X1 U11124 ( .A1(n9955), .A2(n10009), .ZN(n9960) );
  OAI22_X1 U11125 ( .A1(n9957), .A2(n10013), .B1(n9956), .B2(n10011), .ZN(
        n9958) );
  INV_X1 U11126 ( .A(n9958), .ZN(n9959) );
  NAND2_X1 U11127 ( .A1(n9960), .A2(n9959), .ZN(n10087) );
  AOI211_X1 U11128 ( .C1(n9962), .C2(n9979), .A(n10266), .B(n9961), .ZN(n10088) );
  NAND2_X1 U11129 ( .A1(n10088), .A2(n10021), .ZN(n9965) );
  AOI22_X1 U11130 ( .A1(n9986), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9963), .B2(
        n10022), .ZN(n9964) );
  OAI211_X1 U11131 ( .C1(n10155), .C2(n10026), .A(n9965), .B(n9964), .ZN(n9966) );
  AOI21_X1 U11132 ( .B1(n10087), .B2(n10028), .A(n9966), .ZN(n9967) );
  OAI21_X1 U11133 ( .B1(n9968), .B2(n10030), .A(n9967), .ZN(P1_U3273) );
  OAI21_X1 U11134 ( .B1(n9975), .B2(n9970), .A(n9969), .ZN(n9973) );
  AOI222_X1 U11135 ( .A1(n10009), .A2(n9973), .B1(n9972), .B2(n9999), .C1(
        n9971), .C2(n9997), .ZN(n10092) );
  XOR2_X1 U11136 ( .A(n9975), .B(n9974), .Z(n10095) );
  NAND2_X1 U11137 ( .A1(n10095), .A2(n9976), .ZN(n9985) );
  NAND2_X1 U11138 ( .A1(n9977), .A2(n9988), .ZN(n9978) );
  NOR2_X1 U11139 ( .A1(n10159), .A2(n10026), .ZN(n9983) );
  OAI22_X1 U11140 ( .A1(n10028), .A2(n9066), .B1(n9981), .B2(n9980), .ZN(n9982) );
  AOI211_X1 U11141 ( .C1(n10094), .C2(n10021), .A(n9983), .B(n9982), .ZN(n9984) );
  OAI211_X1 U11142 ( .C1(n9986), .C2(n10092), .A(n9985), .B(n9984), .ZN(
        P1_U3274) );
  XNOR2_X1 U11143 ( .A(n9987), .B(n9996), .ZN(n10102) );
  INV_X1 U11144 ( .A(n10018), .ZN(n9990) );
  INV_X1 U11145 ( .A(n9988), .ZN(n9989) );
  AOI211_X1 U11146 ( .C1(n10099), .C2(n9990), .A(n10266), .B(n9989), .ZN(
        n10098) );
  AOI22_X1 U11147 ( .A1(n9986), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9991), .B2(
        n10022), .ZN(n9992) );
  OAI21_X1 U11148 ( .B1(n9993), .B2(n10026), .A(n9992), .ZN(n10003) );
  OAI21_X1 U11149 ( .B1(n9996), .B2(n9995), .A(n9994), .ZN(n10001) );
  AOI222_X1 U11150 ( .A1(n10009), .A2(n10001), .B1(n10000), .B2(n9999), .C1(
        n9998), .C2(n9997), .ZN(n10101) );
  NOR2_X1 U11151 ( .A1(n10101), .A2(n9986), .ZN(n10002) );
  AOI211_X1 U11152 ( .C1(n10098), .C2(n10021), .A(n10003), .B(n10002), .ZN(
        n10004) );
  OAI21_X1 U11153 ( .B1(n10102), .B2(n10030), .A(n10004), .ZN(P1_U3275) );
  XNOR2_X1 U11154 ( .A(n10005), .B(n10006), .ZN(n10105) );
  INV_X1 U11155 ( .A(n10105), .ZN(n10031) );
  INV_X1 U11156 ( .A(n10006), .ZN(n10007) );
  XNOR2_X1 U11157 ( .A(n10008), .B(n10007), .ZN(n10010) );
  NAND2_X1 U11158 ( .A1(n10010), .A2(n10009), .ZN(n10017) );
  OAI22_X1 U11159 ( .A1(n10014), .A2(n10013), .B1(n10012), .B2(n10011), .ZN(
        n10015) );
  INV_X1 U11160 ( .A(n10015), .ZN(n10016) );
  NAND2_X1 U11161 ( .A1(n10017), .A2(n10016), .ZN(n10103) );
  AOI211_X1 U11162 ( .C1(n10020), .C2(n10019), .A(n10266), .B(n10018), .ZN(
        n10104) );
  NAND2_X1 U11163 ( .A1(n10104), .A2(n10021), .ZN(n10025) );
  AOI22_X1 U11164 ( .A1(n9986), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n10023), 
        .B2(n10022), .ZN(n10024) );
  OAI211_X1 U11165 ( .C1(n10165), .C2(n10026), .A(n10025), .B(n10024), .ZN(
        n10027) );
  AOI21_X1 U11166 ( .B1(n10028), .B2(n10103), .A(n10027), .ZN(n10029) );
  OAI21_X1 U11167 ( .B1(n10031), .B2(n10030), .A(n10029), .ZN(P1_U3276) );
  INV_X1 U11168 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n10033) );
  MUX2_X1 U11169 ( .A(n10033), .B(n10123), .S(n10293), .Z(n10034) );
  OAI21_X1 U11170 ( .B1(n10125), .B2(n10108), .A(n10034), .ZN(P1_U3553) );
  INV_X1 U11171 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10037) );
  AND2_X1 U11172 ( .A1(n10036), .A2(n10035), .ZN(n10126) );
  MUX2_X1 U11173 ( .A(n10037), .B(n10126), .S(n10293), .Z(n10038) );
  OAI21_X1 U11174 ( .B1(n4661), .B2(n10108), .A(n10038), .ZN(P1_U3552) );
  NAND2_X1 U11175 ( .A1(n10039), .A2(n10276), .ZN(n10044) );
  NAND2_X1 U11176 ( .A1(n10044), .A2(n10043), .ZN(n10129) );
  MUX2_X1 U11177 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n10129), .S(n10293), .Z(
        P1_U3551) );
  INV_X1 U11178 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n10049) );
  NAND2_X1 U11179 ( .A1(n10046), .A2(n10045), .ZN(n10047) );
  AOI21_X1 U11180 ( .B1(n10048), .B2(n10276), .A(n10047), .ZN(n10130) );
  MUX2_X1 U11181 ( .A(n10049), .B(n10130), .S(n10293), .Z(n10050) );
  OAI21_X1 U11182 ( .B1(n10133), .B2(n10108), .A(n10050), .ZN(P1_U3550) );
  AOI211_X1 U11183 ( .C1(n10053), .C2(n10276), .A(n10052), .B(n10051), .ZN(
        n10134) );
  MUX2_X1 U11184 ( .A(n10054), .B(n10134), .S(n10293), .Z(n10055) );
  OAI21_X1 U11185 ( .B1(n4863), .B2(n10108), .A(n10055), .ZN(P1_U3549) );
  AOI211_X1 U11186 ( .C1(n10117), .C2(n10058), .A(n10057), .B(n10056), .ZN(
        n10059) );
  OAI21_X1 U11187 ( .B1(n10060), .B2(n10113), .A(n10059), .ZN(n10137) );
  MUX2_X1 U11188 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10137), .S(n10293), .Z(
        P1_U3548) );
  INV_X1 U11189 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n10064) );
  AOI211_X1 U11190 ( .C1(n10063), .C2(n10276), .A(n10062), .B(n10061), .ZN(
        n10138) );
  MUX2_X1 U11191 ( .A(n10064), .B(n10138), .S(n10293), .Z(n10065) );
  OAI21_X1 U11192 ( .B1(n10141), .B2(n10108), .A(n10065), .ZN(P1_U3547) );
  INV_X1 U11193 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n10069) );
  AOI211_X1 U11194 ( .C1(n10068), .C2(n10276), .A(n10067), .B(n10066), .ZN(
        n10142) );
  MUX2_X1 U11195 ( .A(n10069), .B(n10142), .S(n10293), .Z(n10070) );
  OAI21_X1 U11196 ( .B1(n10145), .B2(n10108), .A(n10070), .ZN(P1_U3546) );
  AOI22_X1 U11197 ( .A1(n10073), .A2(n10072), .B1(n10117), .B2(n10071), .ZN(
        n10074) );
  OAI211_X1 U11198 ( .C1(n10076), .C2(n10113), .A(n10075), .B(n10074), .ZN(
        n10146) );
  MUX2_X1 U11199 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10146), .S(n10293), .Z(
        P1_U3545) );
  AOI211_X1 U11200 ( .C1(n10117), .C2(n10079), .A(n10078), .B(n10077), .ZN(
        n10080) );
  OAI21_X1 U11201 ( .B1(n10081), .B2(n10113), .A(n10080), .ZN(n10147) );
  MUX2_X1 U11202 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10147), .S(n10293), .Z(
        P1_U3544) );
  INV_X1 U11203 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10085) );
  AOI211_X1 U11204 ( .C1(n10084), .C2(n10276), .A(n10083), .B(n10082), .ZN(
        n10148) );
  MUX2_X1 U11205 ( .A(n10085), .B(n10148), .S(n10293), .Z(n10086) );
  OAI21_X1 U11206 ( .B1(n10151), .B2(n10108), .A(n10086), .ZN(P1_U3543) );
  AOI211_X1 U11207 ( .C1(n10089), .C2(n10276), .A(n10088), .B(n10087), .ZN(
        n10152) );
  MUX2_X1 U11208 ( .A(n10090), .B(n10152), .S(n10293), .Z(n10091) );
  OAI21_X1 U11209 ( .B1(n10155), .B2(n10108), .A(n10091), .ZN(P1_U3542) );
  INV_X1 U11210 ( .A(n10092), .ZN(n10093) );
  AOI211_X1 U11211 ( .C1(n10095), .C2(n10276), .A(n10094), .B(n10093), .ZN(
        n10156) );
  MUX2_X1 U11212 ( .A(n10096), .B(n10156), .S(n10293), .Z(n10097) );
  OAI21_X1 U11213 ( .B1(n10159), .B2(n10108), .A(n10097), .ZN(P1_U3541) );
  AOI21_X1 U11214 ( .B1(n10117), .B2(n10099), .A(n10098), .ZN(n10100) );
  OAI211_X1 U11215 ( .C1(n10102), .C2(n10113), .A(n10101), .B(n10100), .ZN(
        n10160) );
  MUX2_X1 U11216 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10160), .S(n10293), .Z(
        P1_U3540) );
  AOI211_X1 U11217 ( .C1(n10105), .C2(n10276), .A(n10104), .B(n10103), .ZN(
        n10161) );
  MUX2_X1 U11218 ( .A(n10106), .B(n10161), .S(n10293), .Z(n10107) );
  OAI21_X1 U11219 ( .B1(n10165), .B2(n10108), .A(n10107), .ZN(P1_U3539) );
  AOI211_X1 U11220 ( .C1(n10117), .C2(n10111), .A(n10110), .B(n10109), .ZN(
        n10112) );
  OAI21_X1 U11221 ( .B1(n10114), .B2(n10113), .A(n10112), .ZN(n10166) );
  MUX2_X1 U11222 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10166), .S(n10293), .Z(
        P1_U3538) );
  AOI21_X1 U11223 ( .B1(n10117), .B2(n10116), .A(n10115), .ZN(n10118) );
  OAI211_X1 U11224 ( .C1(n10121), .C2(n10120), .A(n10119), .B(n10118), .ZN(
        n10167) );
  MUX2_X1 U11225 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10167), .S(n10293), .Z(
        P1_U3536) );
  MUX2_X1 U11226 ( .A(n10122), .B(P1_REG1_REG_0__SCAN_IN), .S(n10290), .Z(
        P1_U3522) );
  INV_X1 U11227 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n10124) );
  MUX2_X1 U11228 ( .A(n10127), .B(n10126), .S(n10280), .Z(n10128) );
  OAI21_X1 U11229 ( .B1(n4661), .B2(n10164), .A(n10128), .ZN(P1_U3520) );
  MUX2_X1 U11230 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10129), .S(n10280), .Z(
        P1_U3519) );
  INV_X1 U11231 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n10131) );
  MUX2_X1 U11232 ( .A(n10131), .B(n10130), .S(n10280), .Z(n10132) );
  OAI21_X1 U11233 ( .B1(n10133), .B2(n10164), .A(n10132), .ZN(P1_U3518) );
  INV_X1 U11234 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10135) );
  MUX2_X1 U11235 ( .A(n10135), .B(n10134), .S(n10280), .Z(n10136) );
  OAI21_X1 U11236 ( .B1(n4863), .B2(n10164), .A(n10136), .ZN(P1_U3517) );
  MUX2_X1 U11237 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10137), .S(n10280), .Z(
        P1_U3516) );
  MUX2_X1 U11238 ( .A(n10139), .B(n10138), .S(n10280), .Z(n10140) );
  OAI21_X1 U11239 ( .B1(n10141), .B2(n10164), .A(n10140), .ZN(P1_U3515) );
  MUX2_X1 U11240 ( .A(n10143), .B(n10142), .S(n10280), .Z(n10144) );
  OAI21_X1 U11241 ( .B1(n10145), .B2(n10164), .A(n10144), .ZN(P1_U3514) );
  MUX2_X1 U11242 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10146), .S(n10280), .Z(
        P1_U3513) );
  MUX2_X1 U11243 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10147), .S(n10280), .Z(
        P1_U3512) );
  INV_X1 U11244 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10149) );
  MUX2_X1 U11245 ( .A(n10149), .B(n10148), .S(n10280), .Z(n10150) );
  OAI21_X1 U11246 ( .B1(n10151), .B2(n10164), .A(n10150), .ZN(P1_U3511) );
  INV_X1 U11247 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10153) );
  MUX2_X1 U11248 ( .A(n10153), .B(n10152), .S(n10280), .Z(n10154) );
  OAI21_X1 U11249 ( .B1(n10155), .B2(n10164), .A(n10154), .ZN(P1_U3510) );
  INV_X1 U11250 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n10157) );
  MUX2_X1 U11251 ( .A(n10157), .B(n10156), .S(n10280), .Z(n10158) );
  OAI21_X1 U11252 ( .B1(n10159), .B2(n10164), .A(n10158), .ZN(P1_U3509) );
  MUX2_X1 U11253 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10160), .S(n10280), .Z(
        P1_U3507) );
  INV_X1 U11254 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n10162) );
  MUX2_X1 U11255 ( .A(n10162), .B(n10161), .S(n10280), .Z(n10163) );
  OAI21_X1 U11256 ( .B1(n10165), .B2(n10164), .A(n10163), .ZN(P1_U3504) );
  MUX2_X1 U11257 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10166), .S(n10280), .Z(
        P1_U3501) );
  MUX2_X1 U11258 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10167), .S(n10280), .Z(
        P1_U3495) );
  MUX2_X1 U11259 ( .A(n10168), .B(P1_D_REG_0__SCAN_IN), .S(n10239), .Z(
        P1_U3439) );
  NOR4_X1 U11260 ( .A1(n5291), .A2(P1_IR_REG_30__SCAN_IN), .A3(n10169), .A4(
        P1_U3086), .ZN(n10170) );
  AOI21_X1 U11261 ( .B1(n10171), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10170), 
        .ZN(n10172) );
  OAI21_X1 U11262 ( .B1(n10174), .B2(n10173), .A(n10172), .ZN(P1_U3324) );
  MUX2_X1 U11263 ( .A(n10175), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  NAND2_X1 U11264 ( .A1(n10359), .A2(n10176), .ZN(n10178) );
  NAND2_X1 U11265 ( .A1(n10178), .A2(n10189), .ZN(n10177) );
  OAI21_X1 U11266 ( .B1(n10178), .B2(n10189), .A(n10177), .ZN(n10179) );
  INV_X1 U11267 ( .A(n10179), .ZN(n10202) );
  INV_X1 U11268 ( .A(n10180), .ZN(n10199) );
  OAI22_X1 U11269 ( .A1(n10199), .A2(n10183), .B1(n10182), .B2(n10181), .ZN(
        n10195) );
  NAND2_X1 U11270 ( .A1(n10185), .A2(n10184), .ZN(n10187) );
  NAND2_X1 U11271 ( .A1(n10187), .A2(n10186), .ZN(n10188) );
  XOR2_X1 U11272 ( .A(n10189), .B(n10188), .Z(n10190) );
  OAI222_X1 U11273 ( .A1(n10194), .A2(n10193), .B1(n10192), .B2(n10191), .C1(
        n10296), .C2(n10190), .ZN(n10200) );
  AOI211_X1 U11274 ( .C1(n10202), .C2(n10196), .A(n10195), .B(n10200), .ZN(
        n10197) );
  AOI22_X1 U11275 ( .A1(n10198), .A2(n7051), .B1(n10197), .B2(n8724), .ZN(
        P2_U3220) );
  NOR2_X1 U11276 ( .A1(n10199), .A2(n10352), .ZN(n10201) );
  AOI211_X1 U11277 ( .C1(n10202), .C2(n10358), .A(n10201), .B(n10200), .ZN(
        n10203) );
  AOI22_X1 U11278 ( .A1(n10381), .A2(n10203), .B1(n7054), .B2(n10378), .ZN(
        P2_U3472) );
  INV_X1 U11279 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10204) );
  AOI22_X1 U11280 ( .A1(n10366), .A2(n10204), .B1(n10203), .B2(n10364), .ZN(
        P2_U3429) );
  XNOR2_X1 U11281 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XOR2_X1 U11282 ( .A(P2_RD_REG_SCAN_IN), .B(n4712), .Z(U126) );
  NOR2_X4 U11283 ( .A1(n10239), .A2(n10205), .ZN(n10236) );
  INV_X1 U11284 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10206) );
  NOR2_X1 U11285 ( .A1(n10236), .A2(n10206), .ZN(P1_U3294) );
  INV_X1 U11286 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10207) );
  NOR2_X1 U11287 ( .A1(n10236), .A2(n10207), .ZN(P1_U3295) );
  INV_X1 U11288 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10208) );
  NOR2_X1 U11289 ( .A1(n10236), .A2(n10208), .ZN(P1_U3296) );
  NOR2_X1 U11290 ( .A1(n10236), .A2(n10209), .ZN(P1_U3297) );
  INV_X1 U11291 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10210) );
  NOR2_X1 U11292 ( .A1(n10236), .A2(n10210), .ZN(P1_U3298) );
  INV_X1 U11293 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10211) );
  NOR2_X1 U11294 ( .A1(n10236), .A2(n10211), .ZN(P1_U3299) );
  INV_X1 U11295 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10212) );
  NOR2_X1 U11296 ( .A1(n10236), .A2(n10212), .ZN(P1_U3300) );
  INV_X1 U11297 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10213) );
  NOR2_X1 U11298 ( .A1(n10236), .A2(n10213), .ZN(P1_U3301) );
  INV_X1 U11299 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10214) );
  NOR2_X1 U11300 ( .A1(n10236), .A2(n10214), .ZN(P1_U3302) );
  INV_X1 U11301 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10215) );
  NOR2_X1 U11302 ( .A1(n10236), .A2(n10215), .ZN(P1_U3303) );
  INV_X1 U11303 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10216) );
  NOR2_X1 U11304 ( .A1(n10236), .A2(n10216), .ZN(P1_U3304) );
  INV_X1 U11305 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10217) );
  NOR2_X1 U11306 ( .A1(n10236), .A2(n10217), .ZN(P1_U3305) );
  INV_X1 U11307 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10218) );
  NOR2_X1 U11308 ( .A1(n10236), .A2(n10218), .ZN(P1_U3306) );
  INV_X1 U11309 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10219) );
  NOR2_X1 U11310 ( .A1(n10236), .A2(n10219), .ZN(P1_U3307) );
  INV_X1 U11311 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10220) );
  NOR2_X1 U11312 ( .A1(n10236), .A2(n10220), .ZN(P1_U3308) );
  INV_X1 U11313 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10221) );
  NOR2_X1 U11314 ( .A1(n10236), .A2(n10221), .ZN(P1_U3309) );
  NOR2_X1 U11315 ( .A1(n10236), .A2(n10222), .ZN(P1_U3310) );
  INV_X1 U11316 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10223) );
  NOR2_X1 U11317 ( .A1(n10236), .A2(n10223), .ZN(P1_U3311) );
  NOR2_X1 U11318 ( .A1(n10236), .A2(n10224), .ZN(P1_U3312) );
  INV_X1 U11319 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10225) );
  NOR2_X1 U11320 ( .A1(n10236), .A2(n10225), .ZN(P1_U3313) );
  INV_X1 U11321 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10226) );
  NOR2_X1 U11322 ( .A1(n10236), .A2(n10226), .ZN(P1_U3314) );
  INV_X1 U11323 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10227) );
  NOR2_X1 U11324 ( .A1(n10236), .A2(n10227), .ZN(P1_U3315) );
  NOR2_X1 U11325 ( .A1(n10236), .A2(n10228), .ZN(P1_U3316) );
  INV_X1 U11326 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10229) );
  NOR2_X1 U11327 ( .A1(n10236), .A2(n10229), .ZN(P1_U3317) );
  INV_X1 U11328 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10230) );
  NOR2_X1 U11329 ( .A1(n10236), .A2(n10230), .ZN(P1_U3318) );
  INV_X1 U11330 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10231) );
  NOR2_X1 U11331 ( .A1(n10236), .A2(n10231), .ZN(P1_U3319) );
  INV_X1 U11332 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10232) );
  NOR2_X1 U11333 ( .A1(n10236), .A2(n10232), .ZN(P1_U3320) );
  INV_X1 U11334 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10233) );
  NOR2_X1 U11335 ( .A1(n10236), .A2(n10233), .ZN(P1_U3321) );
  NOR2_X1 U11336 ( .A1(n10236), .A2(n10234), .ZN(P1_U3322) );
  INV_X1 U11337 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10235) );
  NOR2_X1 U11338 ( .A1(n10236), .A2(n10235), .ZN(P1_U3323) );
  AOI21_X1 U11339 ( .B1(n10239), .B2(n10238), .A(n10237), .ZN(P1_U3440) );
  OAI22_X1 U11340 ( .A1(n10240), .A2(n10266), .B1(n5736), .B2(n10274), .ZN(
        n10243) );
  INV_X1 U11341 ( .A(n10241), .ZN(n10242) );
  AOI211_X1 U11342 ( .C1(n10276), .C2(n10244), .A(n10243), .B(n10242), .ZN(
        n10282) );
  INV_X1 U11343 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10245) );
  AOI22_X1 U11344 ( .A1(n10280), .A2(n10282), .B1(n10245), .B2(n10278), .ZN(
        P1_U3459) );
  OAI21_X1 U11345 ( .B1(n10247), .B2(n10274), .A(n10246), .ZN(n10250) );
  INV_X1 U11346 ( .A(n10248), .ZN(n10249) );
  AOI211_X1 U11347 ( .C1(n10276), .C2(n10251), .A(n10250), .B(n10249), .ZN(
        n10283) );
  INV_X1 U11348 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10252) );
  AOI22_X1 U11349 ( .A1(n10280), .A2(n10283), .B1(n10252), .B2(n10278), .ZN(
        P1_U3465) );
  OAI21_X1 U11350 ( .B1(n10254), .B2(n10274), .A(n10253), .ZN(n10255) );
  AOI21_X1 U11351 ( .B1(n10256), .B2(n10276), .A(n10255), .ZN(n10257) );
  AND2_X1 U11352 ( .A1(n10258), .A2(n10257), .ZN(n10285) );
  INV_X1 U11353 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10259) );
  AOI22_X1 U11354 ( .A1(n10280), .A2(n10285), .B1(n10259), .B2(n10278), .ZN(
        P1_U3471) );
  OAI21_X1 U11355 ( .B1(n4837), .B2(n10274), .A(n10260), .ZN(n10262) );
  AOI211_X1 U11356 ( .C1(n10276), .C2(n10263), .A(n10262), .B(n10261), .ZN(
        n10287) );
  INV_X1 U11357 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10264) );
  AOI22_X1 U11358 ( .A1(n10280), .A2(n10287), .B1(n10264), .B2(n10278), .ZN(
        P1_U3480) );
  OAI22_X1 U11359 ( .A1(n10267), .A2(n10266), .B1(n10265), .B2(n10274), .ZN(
        n10268) );
  AOI211_X1 U11360 ( .C1(n10270), .C2(n10276), .A(n10269), .B(n10268), .ZN(
        n10289) );
  INV_X1 U11361 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10271) );
  AOI22_X1 U11362 ( .A1(n10280), .A2(n10289), .B1(n10271), .B2(n10278), .ZN(
        P1_U3483) );
  OAI211_X1 U11363 ( .C1(n4861), .C2(n10274), .A(n10273), .B(n10272), .ZN(
        n10275) );
  AOI21_X1 U11364 ( .B1(n10277), .B2(n10276), .A(n10275), .ZN(n10292) );
  INV_X1 U11365 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10279) );
  AOI22_X1 U11366 ( .A1(n10280), .A2(n10292), .B1(n10279), .B2(n10278), .ZN(
        P1_U3489) );
  AOI22_X1 U11367 ( .A1(n10293), .A2(n10282), .B1(n10281), .B2(n10290), .ZN(
        P1_U3524) );
  AOI22_X1 U11368 ( .A1(n10293), .A2(n10283), .B1(n5416), .B2(n10290), .ZN(
        P1_U3526) );
  INV_X1 U11369 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10284) );
  AOI22_X1 U11370 ( .A1(n10293), .A2(n10285), .B1(n10284), .B2(n10290), .ZN(
        P1_U3528) );
  AOI22_X1 U11371 ( .A1(n10293), .A2(n10287), .B1(n10286), .B2(n10290), .ZN(
        P1_U3531) );
  INV_X1 U11372 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10288) );
  AOI22_X1 U11373 ( .A1(n10293), .A2(n10289), .B1(n10288), .B2(n10290), .ZN(
        P1_U3532) );
  AOI22_X1 U11374 ( .A1(n10293), .A2(n10292), .B1(n10291), .B2(n10290), .ZN(
        P1_U3534) );
  INV_X1 U11375 ( .A(n10294), .ZN(n10298) );
  INV_X1 U11376 ( .A(n10358), .ZN(n10329) );
  AOI21_X1 U11377 ( .B1(n10296), .B2(n10329), .A(n10295), .ZN(n10297) );
  AOI211_X1 U11378 ( .C1(n10363), .C2(n10299), .A(n10298), .B(n10297), .ZN(
        n10367) );
  AOI22_X1 U11379 ( .A1(n10366), .A2(n5796), .B1(n10367), .B2(n10364), .ZN(
        P2_U3390) );
  INV_X1 U11380 ( .A(n10304), .ZN(n10301) );
  OAI22_X1 U11381 ( .A1(n10301), .A2(n10344), .B1(n10300), .B2(n10352), .ZN(
        n10302) );
  AOI211_X1 U11382 ( .C1(n10349), .C2(n10304), .A(n10303), .B(n10302), .ZN(
        n10368) );
  AOI22_X1 U11383 ( .A1(n10366), .A2(n5790), .B1(n10368), .B2(n10364), .ZN(
        P2_U3393) );
  OAI21_X1 U11384 ( .B1(n10306), .B2(n10352), .A(n10305), .ZN(n10307) );
  AOI21_X1 U11385 ( .B1(n10308), .B2(n10358), .A(n10307), .ZN(n10369) );
  AOI22_X1 U11386 ( .A1(n10366), .A2(n5822), .B1(n10369), .B2(n10364), .ZN(
        P2_U3399) );
  INV_X1 U11387 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10313) );
  NOR2_X1 U11388 ( .A1(n10309), .A2(n10352), .ZN(n10311) );
  AOI211_X1 U11389 ( .C1(n10312), .C2(n10358), .A(n10311), .B(n10310), .ZN(
        n10370) );
  AOI22_X1 U11390 ( .A1(n10366), .A2(n10313), .B1(n10370), .B2(n10364), .ZN(
        P2_U3402) );
  NOR2_X1 U11391 ( .A1(n10314), .A2(n10352), .ZN(n10316) );
  AOI211_X1 U11392 ( .C1(n10318), .C2(n10317), .A(n10316), .B(n10315), .ZN(
        n10371) );
  AOI22_X1 U11393 ( .A1(n10366), .A2(n6103), .B1(n10371), .B2(n10364), .ZN(
        P2_U3405) );
  INV_X1 U11394 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10323) );
  NOR2_X1 U11395 ( .A1(n10319), .A2(n10329), .ZN(n10321) );
  AOI211_X1 U11396 ( .C1(n10363), .C2(n10322), .A(n10321), .B(n10320), .ZN(
        n10372) );
  AOI22_X1 U11397 ( .A1(n10366), .A2(n10323), .B1(n10372), .B2(n10364), .ZN(
        P2_U3408) );
  INV_X1 U11398 ( .A(n10328), .ZN(n10325) );
  OAI22_X1 U11399 ( .A1(n10325), .A2(n10344), .B1(n10324), .B2(n10352), .ZN(
        n10326) );
  AOI211_X1 U11400 ( .C1(n10349), .C2(n10328), .A(n10327), .B(n10326), .ZN(
        n10373) );
  AOI22_X1 U11401 ( .A1(n10366), .A2(n6576), .B1(n10373), .B2(n10364), .ZN(
        P2_U3411) );
  NOR2_X1 U11402 ( .A1(n10330), .A2(n10329), .ZN(n10332) );
  AOI211_X1 U11403 ( .C1(n10363), .C2(n10333), .A(n10332), .B(n10331), .ZN(
        n10374) );
  AOI22_X1 U11404 ( .A1(n10366), .A2(n5322), .B1(n10374), .B2(n10364), .ZN(
        P2_U3414) );
  INV_X1 U11405 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10341) );
  INV_X1 U11406 ( .A(n10334), .ZN(n10335) );
  OAI22_X1 U11407 ( .A1(n10337), .A2(n10344), .B1(n10335), .B2(n10352), .ZN(
        n10339) );
  NOR2_X1 U11408 ( .A1(n10337), .A2(n10336), .ZN(n10338) );
  NOR3_X1 U11409 ( .A1(n10340), .A2(n10339), .A3(n10338), .ZN(n10375) );
  AOI22_X1 U11410 ( .A1(n10366), .A2(n10341), .B1(n10375), .B2(n10364), .ZN(
        P2_U3417) );
  INV_X1 U11411 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10350) );
  INV_X1 U11412 ( .A(n10342), .ZN(n10343) );
  OAI22_X1 U11413 ( .A1(n10345), .A2(n10344), .B1(n10343), .B2(n10352), .ZN(
        n10347) );
  AOI211_X1 U11414 ( .C1(n10349), .C2(n10348), .A(n10347), .B(n10346), .ZN(
        n10376) );
  AOI22_X1 U11415 ( .A1(n10366), .A2(n10350), .B1(n10376), .B2(n10364), .ZN(
        P2_U3420) );
  INV_X1 U11416 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10356) );
  OAI21_X1 U11417 ( .B1(n10353), .B2(n10352), .A(n10351), .ZN(n10354) );
  AOI21_X1 U11418 ( .B1(n10355), .B2(n10358), .A(n10354), .ZN(n10377) );
  AOI22_X1 U11419 ( .A1(n10366), .A2(n10356), .B1(n10377), .B2(n10364), .ZN(
        P2_U3423) );
  INV_X1 U11420 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10365) );
  AND3_X1 U11421 ( .A1(n10359), .A2(n10358), .A3(n10357), .ZN(n10361) );
  AOI211_X1 U11422 ( .C1(n10363), .C2(n10362), .A(n10361), .B(n10360), .ZN(
        n10380) );
  AOI22_X1 U11423 ( .A1(n10366), .A2(n10365), .B1(n10380), .B2(n10364), .ZN(
        P2_U3426) );
  AOI22_X1 U11424 ( .A1(n10381), .A2(n10367), .B1(n5795), .B2(n10378), .ZN(
        P2_U3459) );
  AOI22_X1 U11425 ( .A1(n10381), .A2(n10368), .B1(n5789), .B2(n10378), .ZN(
        P2_U3460) );
  AOI22_X1 U11426 ( .A1(n10381), .A2(n10369), .B1(n5824), .B2(n10378), .ZN(
        P2_U3462) );
  AOI22_X1 U11427 ( .A1(n10381), .A2(n10370), .B1(n6043), .B2(n10378), .ZN(
        P2_U3463) );
  AOI22_X1 U11428 ( .A1(n10381), .A2(n10371), .B1(n6107), .B2(n10378), .ZN(
        P2_U3464) );
  AOI22_X1 U11429 ( .A1(n10381), .A2(n10372), .B1(n6242), .B2(n10378), .ZN(
        P2_U3465) );
  AOI22_X1 U11430 ( .A1(n10381), .A2(n10373), .B1(n6580), .B2(n10378), .ZN(
        P2_U3466) );
  AOI22_X1 U11431 ( .A1(n10381), .A2(n10374), .B1(n6012), .B2(n10378), .ZN(
        P2_U3467) );
  AOI22_X1 U11432 ( .A1(n10381), .A2(n10375), .B1(n6123), .B2(n10378), .ZN(
        P2_U3468) );
  AOI22_X1 U11433 ( .A1(n10381), .A2(n10376), .B1(n6613), .B2(n10378), .ZN(
        P2_U3469) );
  AOI22_X1 U11434 ( .A1(n10381), .A2(n10377), .B1(n6382), .B2(n10378), .ZN(
        P2_U3470) );
  AOI22_X1 U11435 ( .A1(n10381), .A2(n10380), .B1(n10379), .B2(n10378), .ZN(
        P2_U3471) );
  OAI222_X1 U11436 ( .A1(n10386), .A2(n10385), .B1(n10386), .B2(n10384), .C1(
        n10383), .C2(n10382), .ZN(ADD_1068_U5) );
  XOR2_X1 U11437 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI21_X1 U11438 ( .B1(n10389), .B2(n10388), .A(n10387), .ZN(n10390) );
  XNOR2_X1 U11439 ( .A(n10390), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1068_U55)
         );
  OAI21_X1 U11440 ( .B1(n10393), .B2(n10392), .A(n10391), .ZN(ADD_1068_U56) );
  OAI21_X1 U11441 ( .B1(n10396), .B2(n10395), .A(n10394), .ZN(ADD_1068_U57) );
  OAI21_X1 U11442 ( .B1(n10399), .B2(n10398), .A(n10397), .ZN(ADD_1068_U58) );
  OAI21_X1 U11443 ( .B1(n10402), .B2(n10401), .A(n10400), .ZN(ADD_1068_U59) );
  OAI21_X1 U11444 ( .B1(n10405), .B2(n10404), .A(n10403), .ZN(ADD_1068_U60) );
  OAI21_X1 U11445 ( .B1(n10408), .B2(n10407), .A(n10406), .ZN(ADD_1068_U61) );
  OAI21_X1 U11446 ( .B1(n10411), .B2(n10410), .A(n10409), .ZN(ADD_1068_U62) );
  OAI21_X1 U11447 ( .B1(n10414), .B2(n10413), .A(n10412), .ZN(ADD_1068_U63) );
  OAI21_X1 U11448 ( .B1(n10417), .B2(n10416), .A(n10415), .ZN(ADD_1068_U50) );
  OAI21_X1 U11449 ( .B1(n10420), .B2(n10419), .A(n10418), .ZN(ADD_1068_U51) );
  OAI21_X1 U11450 ( .B1(n10423), .B2(n10422), .A(n10421), .ZN(ADD_1068_U47) );
  OAI21_X1 U11451 ( .B1(n10426), .B2(n10425), .A(n10424), .ZN(ADD_1068_U49) );
  OAI21_X1 U11452 ( .B1(n10429), .B2(n10428), .A(n10427), .ZN(ADD_1068_U48) );
  AOI21_X1 U11453 ( .B1(n10432), .B2(n10431), .A(n10430), .ZN(ADD_1068_U54) );
  AOI21_X1 U11454 ( .B1(n10435), .B2(n10434), .A(n10433), .ZN(ADD_1068_U53) );
  OAI21_X1 U11455 ( .B1(n10438), .B2(n10437), .A(n10436), .ZN(ADD_1068_U52) );
  OAI21_X2 U5961 ( .B1(n5156), .B2(n5155), .A(n5154), .ZN(n5280) );
  INV_X1 U4998 ( .A(n8097), .ZN(n8194) );
endmodule

