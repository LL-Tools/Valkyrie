

module b17_C_gen_AntiSAT_k_256_8 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput_f0, keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, 
        keyinput_f5, keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, 
        keyinput_f10, keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, 
        keyinput_f15, keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, 
        keyinput_f20, keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, 
        keyinput_f25, keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, 
        keyinput_f30, keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, 
        keyinput_f35, keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, 
        keyinput_f40, keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, 
        keyinput_f45, keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, 
        keyinput_f50, keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, 
        keyinput_f55, keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, 
        keyinput_f60, keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, 
        keyinput_f65, keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, 
        keyinput_f70, keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, 
        keyinput_f75, keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, 
        keyinput_f80, keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, 
        keyinput_f85, keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, 
        keyinput_f90, keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, 
        keyinput_f95, keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, 
        keyinput_f100, keyinput_f101, keyinput_f102, keyinput_f103, 
        keyinput_f104, keyinput_f105, keyinput_f106, keyinput_f107, 
        keyinput_f108, keyinput_f109, keyinput_f110, keyinput_f111, 
        keyinput_f112, keyinput_f113, keyinput_f114, keyinput_f115, 
        keyinput_f116, keyinput_f117, keyinput_f118, keyinput_f119, 
        keyinput_f120, keyinput_f121, keyinput_f122, keyinput_f123, 
        keyinput_f124, keyinput_f125, keyinput_f126, keyinput_f127, 
        keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3, keyinput_g4, 
        keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8, keyinput_g9, 
        keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13, keyinput_g14, 
        keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18, keyinput_g19, 
        keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23, keyinput_g24, 
        keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28, keyinput_g29, 
        keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33, keyinput_g34, 
        keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38, keyinput_g39, 
        keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43, keyinput_g44, 
        keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48, keyinput_g49, 
        keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53, keyinput_g54, 
        keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58, keyinput_g59, 
        keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63, keyinput_g64, 
        keyinput_g65, keyinput_g66, keyinput_g67, keyinput_g68, keyinput_g69, 
        keyinput_g70, keyinput_g71, keyinput_g72, keyinput_g73, keyinput_g74, 
        keyinput_g75, keyinput_g76, keyinput_g77, keyinput_g78, keyinput_g79, 
        keyinput_g80, keyinput_g81, keyinput_g82, keyinput_g83, keyinput_g84, 
        keyinput_g85, keyinput_g86, keyinput_g87, keyinput_g88, keyinput_g89, 
        keyinput_g90, keyinput_g91, keyinput_g92, keyinput_g93, keyinput_g94, 
        keyinput_g95, keyinput_g96, keyinput_g97, keyinput_g98, keyinput_g99, 
        keyinput_g100, keyinput_g101, keyinput_g102, keyinput_g103, 
        keyinput_g104, keyinput_g105, keyinput_g106, keyinput_g107, 
        keyinput_g108, keyinput_g109, keyinput_g110, keyinput_g111, 
        keyinput_g112, keyinput_g113, keyinput_g114, keyinput_g115, 
        keyinput_g116, keyinput_g117, keyinput_g118, keyinput_g119, 
        keyinput_g120, keyinput_g121, keyinput_g122, keyinput_g123, 
        keyinput_g124, keyinput_g125, keyinput_g126, keyinput_g127, U355, U356, 
        U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, U369, 
        U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, U352, 
        U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, U240, 
        U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, U228, 
        U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, U216, 
        U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, 
        U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, 
        U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, 
        P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, 
        P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, 
        P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, 
        P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, 
        P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, 
        P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, 
        P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, 
        P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, 
        P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, 
        P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, 
        P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, 
        P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, 
        P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, 
        P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, 
        P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, 
        P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, 
        P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, 
        P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, 
        P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, 
        P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, 
        P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, 
        P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, 
        P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, 
        P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, 
        P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, 
        P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, 
        P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, 
        P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, 
        P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, 
        P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, 
        P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, 
        P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, 
        P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, 
        P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, 
        P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, 
        P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, 
        P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, 
        P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, 
        P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, 
        P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, 
        P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, 
        P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, 
        P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, 
        P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, 
        P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, 
        P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, 
        P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, 
        P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, 
        P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, 
        P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, 
        P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, 
        P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, 
        P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, 
        P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, 
        P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, 
        P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, 
        P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, 
        P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, 
        P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, 
        P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, 
        P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, 
        P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, 
        P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, 
        P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, 
        P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, 
        P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, 
        P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, 
        P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, 
        P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, 
        P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, 
        P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, 
        P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, 
        P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, 
        P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, 
        P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, 
        P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, 
        P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, 
        P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, 
        P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, 
        P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, 
        P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, 
        P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, 
        P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, 
        P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, 
        P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, 
        P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, 
        P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, 
        P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, 
        P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, 
        P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, 
        P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, 
        P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, 
        P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, 
        P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, 
        P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, 
        P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, 
        P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, 
        P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, 
        P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, 
        P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, 
        P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, 
        P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, 
        P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, 
        P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, 
        P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, 
        P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, 
        P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, 
        P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, 
        P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, 
        P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, 
        P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, 
        P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, 
        P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, 
        P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, 
        P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, 
        P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, 
        P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, 
        P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, 
        P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, 
        P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, 
        P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, 
        P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, 
        P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, 
        P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, 
        P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, 
        P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, 
        P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, 
        P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, 
        P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, 
        P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, 
        P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, 
        P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, 
        P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, 
        P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, 
        P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, 
        P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, 
        P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, 
        P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, 
        P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, 
        P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, 
        P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, 
        P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, 
        P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, 
        P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, 
        P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, 
        P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, 
        P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, 
        P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, 
        P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, 
        P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, 
        P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, 
        P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, 
        P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, 
        P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, 
        P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, 
        P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, 
        P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, 
        P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, 
        P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, 
        P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, 
        P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, 
        P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, 
        P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, 
        P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, 
        P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, 
        P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, 
        P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, 
        P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, 
        P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, 
        P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, 
        P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, 
        P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, 
        P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, 
        P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, 
        P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, 
        P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, 
        P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, 
        P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, 
        P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, 
        P1_U2802, P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
         n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
         n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
         n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
         n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
         n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
         n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
         n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
         n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
         n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
         n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
         n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702,
         n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
         n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
         n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
         n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
         n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
         n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
         n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822,
         n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830,
         n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
         n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846,
         n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854,
         n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862,
         n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870,
         n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878,
         n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
         n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894,
         n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902,
         n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
         n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918,
         n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
         n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
         n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
         n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
         n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
         n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966,
         n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974,
         n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
         n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
         n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
         n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
         n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
         n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046,
         n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
         n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
         n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
         n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078,
         n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
         n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094,
         n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
         n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
         n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
         n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
         n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
         n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142,
         n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
         n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
         n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166,
         n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
         n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
         n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,
         n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
         n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
         n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
         n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,
         n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
         n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
         n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
         n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
         n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446,
         n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
         n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
         n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
         n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,
         n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486,
         n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,
         n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502,
         n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510,
         n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518,
         n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
         n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534,
         n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
         n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550,
         n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
         n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
         n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
         n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
         n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
         n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
         n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
         n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
         n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
         n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479,
         n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
         n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495,
         n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503,
         n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
         n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
         n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
         n16536, n16537, n16538, n16539, n16540, n16541, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,
         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
         n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
         n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,
         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,
         n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
         n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
         n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
         n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,
         n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,
         n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,
         n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256,
         n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
         n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,
         n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,
         n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
         n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296,
         n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304,
         n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,
         n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
         n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,
         n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,
         n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,
         n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,
         n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
         n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,
         n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376,
         n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,
         n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,
         n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,
         n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408,
         n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,
         n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424,
         n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
         n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440,
         n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448,
         n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,
         n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
         n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,
         n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,
         n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,
         n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,
         n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
         n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512,
         n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520,
         n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528,
         n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,
         n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544,
         n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,
         n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,
         n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,
         n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
         n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584,
         n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592,
         n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,
         n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,
         n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,
         n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,
         n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,
         n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,
         n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
         n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656,
         n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664,
         n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,
         n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,
         n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,
         n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,
         n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,
         n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,
         n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
         n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,
         n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,
         n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,
         n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
         n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,
         n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,
         n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,
         n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,
         n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
         n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800,
         n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808,
         n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,
         n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,
         n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832,
         n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,
         n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
         n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,
         n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
         n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872,
         n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,
         n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,
         n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,
         n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,
         n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,
         n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,
         n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,
         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
         n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,
         n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,
         n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960,
         n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,
         n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976,
         n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
         n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,
         n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,
         n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
         n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,
         n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024,
         n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032,
         n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040,
         n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,
         n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,
         n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,
         n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,
         n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
         n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088,
         n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096,
         n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104,
         n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,
         n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
         n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
         n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,
         n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
         n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160,
         n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168,
         n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176,
         n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,
         n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,
         n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,
         n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
         n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,
         n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
         n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232,
         n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240,
         n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,
         n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,
         n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,
         n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272,
         n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
         n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,
         n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,
         n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304,
         n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312,
         n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,
         n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
         n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
         n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,
         n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
         n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,
         n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,
         n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,
         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,
         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,
         n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
         n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,
         n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,
         n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,
         n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528,
         n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,
         n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,
         n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,
         n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560,
         n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
         n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576,
         n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584,
         n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592,
         n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600,
         n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,
         n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,
         n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
         n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632,
         n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,
         n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648,
         n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,
         n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,
         n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672,
         n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680,
         n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
         n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696,
         n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704,
         n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,
         n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720,
         n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,
         n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736,
         n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,
         n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752,
         n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,
         n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,
         n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776,
         n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,
         n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,
         n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,
         n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,
         n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816,
         n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,
         n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,
         n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840,
         n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848,
         n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,
         n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,
         n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,
         n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,
         n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888,
         n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896,
         n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,
         n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,
         n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920,
         n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,
         n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,
         n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944,
         n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952,
         n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960,
         n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968,
         n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
         n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984,
         n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992,
         n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,
         n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008,
         n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,
         n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024,
         n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032,
         n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040,
         n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048,
         n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056,
         n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064,
         n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,
         n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080,
         n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
         n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096,
         n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104,
         n19105, n19106, n19107, n19108, n19109, n19110, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304;

  AOI21_X1 U11258 ( .B1(n15139), .B2(n15136), .A(n15127), .ZN(n15131) );
  INV_X1 U11259 ( .A(n20069), .ZN(n20021) );
  NAND2_X1 U11260 ( .A1(n14892), .A2(n14894), .ZN(n14887) );
  NAND2_X1 U11261 ( .A1(n13312), .A2(n13311), .ZN(n13392) );
  NOR2_X1 U11263 ( .A1(n13719), .A2(n13718), .ZN(n18253) );
  INV_X1 U11264 ( .A(n13958), .ZN(n10795) );
  INV_X2 U11265 ( .A(n17798), .ZN(n17760) );
  AND2_X1 U11267 ( .A1(n11409), .A2(n10861), .ZN(n11254) );
  AND2_X1 U11268 ( .A1(n10861), .A2(n9839), .ZN(n9887) );
  AND2_X2 U11269 ( .A1(n11408), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11265) );
  AND2_X2 U11270 ( .A1(n10473), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10536) );
  AND2_X1 U11271 ( .A1(n9835), .A2(n10861), .ZN(n11256) );
  CLKBUF_X2 U11272 ( .A(n15581), .Z(n17208) );
  AND2_X1 U11273 ( .A1(n10478), .A2(n10479), .ZN(n11255) );
  CLKBUF_X2 U11274 ( .A(n15676), .Z(n16962) );
  INV_X1 U11275 ( .A(n17018), .ZN(n13703) );
  INV_X2 U11276 ( .A(n9871), .ZN(n17195) );
  CLKBUF_X2 U11277 ( .A(n10967), .Z(n13950) );
  CLKBUF_X1 U11278 ( .A(n13734), .Z(n17189) );
  CLKBUF_X1 U11279 ( .A(n13697), .Z(n17216) );
  BUF_X1 U11280 ( .A(n15603), .Z(n17146) );
  CLKBUF_X1 U11281 ( .A(n15676), .Z(n17217) );
  NOR2_X1 U11282 ( .A1(n10919), .A2(n10918), .ZN(n10960) );
  NOR2_X1 U11283 ( .A1(n13643), .A2(n18704), .ZN(n15713) );
  CLKBUF_X2 U11284 ( .A(n12147), .Z(n12111) );
  CLKBUF_X1 U11285 ( .A(n11561), .Z(n12229) );
  CLKBUF_X2 U11286 ( .A(n11654), .Z(n12284) );
  CLKBUF_X1 U11287 ( .A(n11632), .Z(n20263) );
  AND2_X1 U11288 ( .A1(n11632), .A2(n14328), .ZN(n12736) );
  NAND2_X2 U11289 ( .A1(n9884), .A2(n11576), .ZN(n11623) );
  INV_X1 U11290 ( .A(n11634), .ZN(n20248) );
  AND4_X1 U11291 ( .A1(n11499), .A2(n11498), .A3(n11497), .A4(n11496), .ZN(
        n11515) );
  AND2_X1 U11292 ( .A1(n12673), .A2(n19252), .ZN(n10909) );
  CLKBUF_X2 U11293 ( .A(n11765), .Z(n12146) );
  CLKBUF_X2 U11294 ( .A(n11770), .Z(n12134) );
  AND2_X1 U11295 ( .A1(n11495), .A2(n11505), .ZN(n11752) );
  AND2_X1 U11296 ( .A1(n11505), .A2(n13094), .ZN(n12147) );
  AND2_X1 U11297 ( .A1(n11495), .A2(n14735), .ZN(n11654) );
  CLKBUF_X1 U11298 ( .A(n18738), .Z(n9814) );
  NOR2_X1 U11299 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18863), .ZN(n18738) );
  INV_X1 U11300 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11488) );
  INV_X1 U11301 ( .A(n10433), .ZN(n9840) );
  AND3_X1 U11302 ( .A1(n9963), .A2(n9962), .A3(n9961), .ZN(n9902) );
  NAND2_X1 U11303 ( .A1(n11751), .A2(n11750), .ZN(n12334) );
  CLKBUF_X2 U11304 ( .A(n10843), .Z(n11420) );
  AND2_X1 U11305 ( .A1(n9842), .A2(n10861), .ZN(n11257) );
  AND2_X1 U11306 ( .A1(n11409), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10537) );
  XNOR2_X1 U11307 ( .A(n10960), .B(n10961), .ZN(n11121) );
  INV_X1 U11308 ( .A(n10902), .ZN(n12673) );
  INV_X2 U11309 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10861) );
  NOR2_X1 U11310 ( .A1(n18263), .A2(n18258), .ZN(n13750) );
  INV_X1 U11311 ( .A(n13435), .ZN(n11633) );
  AND2_X1 U11312 ( .A1(n13876), .A2(n13875), .ZN(n13878) );
  INV_X1 U11313 ( .A(n10774), .ZN(n13955) );
  OAI21_X1 U11314 ( .B1(n10240), .B2(n9982), .A(n9981), .ZN(n15118) );
  AND2_X1 U11315 ( .A1(n13395), .A2(n13394), .ZN(n13397) );
  NAND2_X1 U11317 ( .A1(n21304), .A2(n13193), .ZN(n13366) );
  BUF_X1 U11318 ( .A(n10855), .Z(n9837) );
  INV_X1 U11320 ( .A(n15711), .ZN(n17018) );
  INV_X1 U11321 ( .A(n15802), .ZN(n13758) );
  INV_X1 U11322 ( .A(n13498), .ZN(n16024) );
  NOR2_X2 U11323 ( .A1(n14502), .A2(n14425), .ZN(n14452) );
  BUF_X1 U11324 ( .A(n11637), .Z(n20231) );
  OR2_X1 U11325 ( .A1(n15067), .A2(n13908), .ZN(n9822) );
  INV_X1 U11326 ( .A(n10906), .ZN(n12679) );
  INV_X1 U11327 ( .A(n13535), .ZN(n10145) );
  NOR2_X1 U11328 ( .A1(n17611), .A2(n17612), .ZN(n16588) );
  INV_X1 U11329 ( .A(n18889), .ZN(n16578) );
  OR2_X1 U11330 ( .A1(n14309), .A2(n14308), .ZN(n14311) );
  XNOR2_X1 U11331 ( .A(n14448), .B(n14447), .ZN(n14617) );
  NAND2_X1 U11332 ( .A1(n11433), .A2(n10906), .ZN(n12667) );
  NOR2_X2 U11333 ( .A1(n13038), .A2(n11133), .ZN(n13129) );
  XNOR2_X1 U11334 ( .A(n11428), .B(n11427), .ZN(n12402) );
  NOR2_X1 U11335 ( .A1(n15066), .A2(n15060), .ZN(n15059) );
  AND2_X1 U11337 ( .A1(n10030), .A2(n9903), .ZN(n16436) );
  INV_X1 U11338 ( .A(n20079), .ZN(n20043) );
  XNOR2_X1 U11339 ( .A(n14073), .B(n14072), .ZN(n14594) );
  NOR2_X2 U11340 ( .A1(n17672), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17671) );
  NOR2_X2 U11341 ( .A1(n14871), .A2(n14874), .ZN(n14873) );
  NAND2_X2 U11342 ( .A1(n15076), .A2(n10327), .ZN(n9830) );
  NOR2_X2 U11343 ( .A1(n16171), .A2(n16170), .ZN(n16173) );
  NOR2_X2 U11344 ( .A1(n13249), .A2(n13238), .ZN(n13309) );
  NOR3_X2 U11345 ( .A1(n17787), .A2(n17750), .A3(n16812), .ZN(n17724) );
  INV_X1 U11346 ( .A(n10911), .ZN(n10855) );
  NAND2_X2 U11347 ( .A1(n14426), .A2(n15984), .ZN(n14502) );
  NOR2_X2 U11349 ( .A1(n17553), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17552) );
  INV_X4 U11350 ( .A(n11416), .ZN(n11408) );
  INV_X2 U11351 ( .A(n17800), .ZN(n17899) );
  XNOR2_X2 U11352 ( .A(n13611), .B(n13618), .ZN(n13610) );
  OAI21_X2 U11353 ( .B1(n13396), .B2(n13927), .A(n19107), .ZN(n13611) );
  NOR4_X4 U11354 ( .A1(n18237), .A2(n13758), .A3(n13757), .A4(n17271), .ZN(
        n17471) );
  NAND3_X1 U11355 ( .A1(n18244), .A2(n18253), .A3(n18263), .ZN(n13757) );
  NOR2_X2 U11356 ( .A1(n10183), .A2(n17579), .ZN(n17566) );
  CLKBUF_X1 U11357 ( .A(n14135), .Z(n14149) );
  NOR2_X1 U11358 ( .A1(n13897), .A2(n10100), .ZN(n10099) );
  OAI21_X2 U11359 ( .B1(n18971), .B2(n13941), .A(n15383), .ZN(n15149) );
  NAND2_X1 U11360 ( .A1(n11829), .A2(n11828), .ZN(n20766) );
  CLKBUF_X1 U11361 ( .A(n12848), .Z(n20631) );
  NAND2_X1 U11362 ( .A1(n13878), .A2(n10886), .ZN(n13872) );
  NOR2_X1 U11363 ( .A1(n16148), .A2(n16147), .ZN(n16150) );
  AND2_X1 U11364 ( .A1(n13838), .A2(n10885), .ZN(n13876) );
  AND2_X1 U11365 ( .A1(n13614), .A2(n13613), .ZN(n13819) );
  AND2_X1 U11366 ( .A1(n12661), .A2(n9980), .ZN(n10919) );
  AND3_X1 U11367 ( .A1(n10908), .A2(n10907), .A3(n12667), .ZN(n15521) );
  NOR2_X1 U11369 ( .A1(n11431), .A2(n19247), .ZN(n10916) );
  NAND3_X1 U11370 ( .A1(n13674), .A2(n13673), .A3(n13672), .ZN(n17415) );
  NAND2_X1 U11371 ( .A1(n10369), .A2(n10368), .ZN(n11634) );
  AND4_X1 U11372 ( .A1(n11493), .A2(n11492), .A3(n11491), .A4(n11490), .ZN(
        n11516) );
  CLKBUF_X2 U11373 ( .A(n11926), .Z(n12288) );
  BUF_X2 U11374 ( .A(n11578), .Z(n12230) );
  CLKBUF_X2 U11375 ( .A(n11607), .Z(n12129) );
  BUF_X2 U11376 ( .A(n15665), .Z(n17197) );
  BUF_X2 U11377 ( .A(n15604), .Z(n17196) );
  BUF_X1 U11378 ( .A(n15604), .Z(n17215) );
  BUF_X4 U11379 ( .A(n13698), .Z(n9817) );
  NOR2_X2 U11380 ( .A1(n11488), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11500) );
  INV_X2 U11381 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10320) );
  NOR2_X4 U11382 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15543) );
  INV_X4 U11383 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18851) );
  NAND2_X1 U11384 ( .A1(n9988), .A2(n9987), .ZN(n15116) );
  OAI21_X1 U11385 ( .B1(n15021), .B2(n10006), .A(n10005), .ZN(n15012) );
  NAND2_X1 U11386 ( .A1(n9815), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15066) );
  AND2_X1 U11387 ( .A1(n15380), .A2(n15379), .ZN(n15404) );
  NAND2_X1 U11388 ( .A1(n10245), .A2(n10246), .ZN(n10244) );
  AOI22_X1 U11389 ( .A1(n14843), .A2(n14844), .B1(n9899), .B2(n14833), .ZN(
        n14936) );
  NAND2_X1 U11390 ( .A1(n10349), .A2(n10353), .ZN(n14833) );
  XNOR2_X1 U11391 ( .A(n14086), .B(n12315), .ZN(n14433) );
  AOI21_X1 U11392 ( .B1(n14087), .B2(n14085), .A(n14086), .ZN(n14442) );
  AND2_X1 U11393 ( .A1(n14120), .A2(n10308), .ZN(n14086) );
  OR2_X1 U11394 ( .A1(n14850), .A2(n14852), .ZN(n9967) );
  NAND2_X1 U11395 ( .A1(n13939), .A2(n13938), .ZN(n16273) );
  NAND2_X1 U11396 ( .A1(n9995), .A2(n13814), .ZN(n15208) );
  AOI21_X1 U11397 ( .B1(n16457), .B2(n16456), .A(n16455), .ZN(n16459) );
  NAND2_X1 U11398 ( .A1(n10329), .A2(n10330), .ZN(n11319) );
  XNOR2_X1 U11399 ( .A(n13940), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16274) );
  CLKBUF_X1 U11400 ( .A(n14524), .Z(n16025) );
  XNOR2_X1 U11401 ( .A(n13942), .B(n13941), .ZN(n15206) );
  OR2_X1 U11402 ( .A1(n13942), .A2(n13941), .ZN(n13940) );
  OR3_X1 U11403 ( .A1(n13942), .A2(n13941), .A3(n11001), .ZN(n13943) );
  NAND2_X1 U11404 ( .A1(n13935), .A2(n13934), .ZN(n13942) );
  AND2_X1 U11405 ( .A1(n11273), .A2(n11296), .ZN(n11274) );
  NAND2_X1 U11406 ( .A1(n10011), .A2(n10012), .ZN(n14567) );
  AND2_X1 U11407 ( .A1(n14862), .A2(n14847), .ZN(n14849) );
  OR2_X2 U11408 ( .A1(n13379), .A2(n9997), .ZN(n13932) );
  NAND2_X1 U11409 ( .A1(n13313), .A2(n13315), .ZN(n13379) );
  AND2_X1 U11410 ( .A1(n16607), .A2(n16878), .ZN(n16601) );
  NAND2_X1 U11411 ( .A1(n13234), .A2(n13233), .ZN(n13237) );
  OR2_X1 U11412 ( .A1(n16609), .A2(n16610), .ZN(n16607) );
  AND2_X1 U11413 ( .A1(n13913), .A2(n10108), .ZN(n9824) );
  NOR3_X2 U11414 ( .A1(n14156), .A2(n10274), .A3(n14099), .ZN(n14098) );
  OR2_X1 U11415 ( .A1(n13375), .A2(n13374), .ZN(n13378) );
  NAND2_X1 U11416 ( .A1(n10098), .A2(n15089), .ZN(n10000) );
  AND2_X1 U11417 ( .A1(n10099), .A2(n15089), .ZN(n9998) );
  AND2_X1 U11418 ( .A1(n13220), .A2(n13219), .ZN(n10373) );
  AND2_X1 U11419 ( .A1(n15360), .A2(n14985), .ZN(n15341) );
  NAND2_X1 U11420 ( .A1(n17628), .A2(n10186), .ZN(n10185) );
  AND2_X1 U11421 ( .A1(n9958), .A2(n9957), .ZN(n9956) );
  AND2_X1 U11422 ( .A1(n9905), .A2(n9960), .ZN(n9959) );
  NAND2_X2 U11423 ( .A1(n15771), .A2(n17760), .ZN(n17628) );
  AND2_X1 U11424 ( .A1(n13205), .A2(n13193), .ZN(n19700) );
  AND2_X1 U11425 ( .A1(n13205), .A2(n13198), .ZN(n19747) );
  AND2_X1 U11426 ( .A1(n13205), .A2(n13199), .ZN(n19624) );
  CLKBUF_X1 U11427 ( .A(n12392), .Z(n14384) );
  CLKBUF_X1 U11428 ( .A(n14329), .Z(n14386) );
  NAND2_X2 U11429 ( .A1(n14391), .A2(n13081), .ZN(n14409) );
  AND2_X1 U11430 ( .A1(n12626), .A2(n11129), .ZN(n12692) );
  INV_X2 U11431 ( .A(n13021), .ZN(n20146) );
  NOR2_X1 U11432 ( .A1(n20395), .A2(n20249), .ZN(n20784) );
  NOR2_X1 U11433 ( .A1(n20395), .A2(n20242), .ZN(n20778) );
  NOR2_X1 U11434 ( .A1(n20395), .A2(n20289), .ZN(n20818) );
  NOR2_X1 U11435 ( .A1(n20395), .A2(n20232), .ZN(n20765) );
  NOR2_X1 U11436 ( .A1(n20395), .A2(n20257), .ZN(n20790) );
  NOR2_X1 U11437 ( .A1(n20395), .A2(n20272), .ZN(n20802) );
  AND2_X1 U11438 ( .A1(n12795), .A2(n14000), .ZN(n20193) );
  NOR2_X1 U11439 ( .A1(n20395), .A2(n20264), .ZN(n20796) );
  NOR2_X1 U11440 ( .A1(n20395), .A2(n20279), .ZN(n20810) );
  NAND2_X1 U11441 ( .A1(n11708), .A2(n10216), .ZN(n11829) );
  AND2_X1 U11442 ( .A1(n15374), .A2(n15377), .ZN(n15381) );
  AND2_X1 U11443 ( .A1(n14244), .A2(n14228), .ZN(n14230) );
  NAND2_X1 U11444 ( .A1(n9825), .A2(n10974), .ZN(n10034) );
  CLKBUF_X1 U11445 ( .A(n12739), .Z(n20323) );
  AND2_X1 U11446 ( .A1(n10026), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15767) );
  NAND2_X2 U11447 ( .A1(n12365), .A2(n12364), .ZN(n14003) );
  INV_X1 U11448 ( .A(n15525), .ZN(n16315) );
  NOR2_X2 U11449 ( .A1(n19253), .A2(n19665), .ZN(n19254) );
  NOR2_X2 U11450 ( .A1(n19248), .A2(n19665), .ZN(n19249) );
  NOR2_X1 U11451 ( .A1(n15916), .A2(n15915), .ZN(n17383) );
  NOR2_X2 U11452 ( .A1(n19239), .A2(n19665), .ZN(n19240) );
  NAND2_X1 U11453 ( .A1(n10977), .A2(n10976), .ZN(n10984) );
  NAND2_X1 U11454 ( .A1(n10971), .A2(n10970), .ZN(n11107) );
  NAND2_X1 U11455 ( .A1(n10982), .A2(n10981), .ZN(n10983) );
  OR2_X1 U11456 ( .A1(n11078), .A2(n13619), .ZN(n10982) );
  NOR2_X1 U11457 ( .A1(n12939), .A2(n12938), .ZN(n13120) );
  NOR3_X1 U11458 ( .A1(n16409), .A2(n16611), .A3(n10121), .ZN(n10117) );
  NOR2_X1 U11459 ( .A1(n13381), .A2(n13380), .ZN(n13614) );
  NOR2_X1 U11460 ( .A1(n17872), .A2(n15758), .ZN(n17864) );
  NOR2_X1 U11461 ( .A1(n17515), .A2(n18889), .ZN(n17521) );
  OR2_X1 U11462 ( .A1(n10937), .A2(n11431), .ZN(n10955) );
  CLKBUF_X1 U11463 ( .A(n12366), .Z(n13085) );
  OR2_X2 U11464 ( .A1(n12399), .A2(n10913), .ZN(n10967) );
  INV_X1 U11465 ( .A(n11742), .ZN(n10064) );
  NOR2_X1 U11466 ( .A1(n17890), .A2(n16413), .ZN(n16581) );
  NAND2_X1 U11467 ( .A1(n15521), .A2(n10909), .ZN(n10943) );
  NAND2_X2 U11468 ( .A1(n10468), .A2(n10522), .ZN(n13958) );
  OR2_X1 U11469 ( .A1(n12400), .A2(n18909), .ZN(n10913) );
  NAND2_X1 U11470 ( .A1(n10371), .A2(n11598), .ZN(n12831) );
  INV_X2 U11471 ( .A(n17415), .ZN(n18237) );
  AND2_X1 U11472 ( .A1(n15661), .A2(n10909), .ZN(n11469) );
  INV_X4 U11473 ( .A(n9837), .ZN(n19267) );
  OR2_X1 U11474 ( .A1(n10583), .A2(n10582), .ZN(n13315) );
  CLKBUF_X1 U11475 ( .A(n11645), .Z(n20278) );
  BUF_X2 U11476 ( .A(n11633), .Z(n20241) );
  NAND2_X1 U11477 ( .A1(n15716), .A2(n9851), .ZN(n17401) );
  AND2_X1 U11478 ( .A1(n15910), .A2(n14067), .ZN(n14062) );
  NAND4_X2 U11479 ( .A1(n10637), .A2(n10636), .A3(n10635), .A4(n10634), .ZN(
        n13927) );
  CLKBUF_X1 U11480 ( .A(n11634), .Z(n12837) );
  AOI211_X1 U11481 ( .C1(n17196), .C2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n13671), .B(n13670), .ZN(n13672) );
  NOR2_X2 U11482 ( .A1(n13654), .A2(n13653), .ZN(n18268) );
  NOR2_X2 U11483 ( .A1(n12740), .A2(n11634), .ZN(n13092) );
  CLKBUF_X1 U11484 ( .A(n13216), .Z(n14748) );
  INV_X1 U11485 ( .A(n14328), .ZN(n20271) );
  NOR2_X1 U11486 ( .A1(n17645), .A2(n17647), .ZN(n17632) );
  OR2_X2 U11487 ( .A1(n16507), .A2(n16463), .ZN(n16509) );
  NAND2_X1 U11488 ( .A1(n10455), .A2(n10454), .ZN(n10911) );
  NAND2_X2 U11489 ( .A1(n10440), .A2(n10439), .ZN(n13216) );
  NAND2_X2 U11490 ( .A1(n10854), .A2(n10853), .ZN(n10915) );
  NAND4_X2 U11491 ( .A1(n11536), .A2(n11535), .A3(n11534), .A4(n11533), .ZN(
        n14328) );
  NAND4_X2 U11492 ( .A1(n11556), .A2(n11555), .A3(n11554), .A4(n11553), .ZN(
        n12792) );
  AND4_X1 U11493 ( .A1(n11540), .A2(n11539), .A3(n11538), .A4(n11537), .ZN(
        n11556) );
  AND4_X1 U11494 ( .A1(n11602), .A2(n11601), .A3(n11600), .A4(n11599), .ZN(
        n11619) );
  NOR2_X1 U11495 ( .A1(n10367), .A2(n11548), .ZN(n11554) );
  NOR2_X1 U11496 ( .A1(n17682), .A2(n17686), .ZN(n17668) );
  NAND4_X1 U11497 ( .A1(n10453), .A2(n10452), .A3(n10451), .A4(n10450), .ZN(
        n10454) );
  NAND2_X2 U11498 ( .A1(n19868), .A2(n19856), .ZN(n19914) );
  NAND2_X2 U11499 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19868), .ZN(n19911) );
  AND4_X1 U11500 ( .A1(n11615), .A2(n11614), .A3(n11613), .A4(n11612), .ZN(
        n11616) );
  AND4_X1 U11501 ( .A1(n11611), .A2(n11610), .A3(n11609), .A4(n11608), .ZN(
        n11617) );
  AND4_X1 U11502 ( .A1(n11575), .A2(n11574), .A3(n11573), .A4(n11572), .ZN(
        n11576) );
  AND4_X1 U11503 ( .A1(n11512), .A2(n11511), .A3(n11510), .A4(n11509), .ZN(
        n11513) );
  AND2_X1 U11504 ( .A1(n10449), .A2(n10448), .ZN(n10453) );
  AND3_X1 U11505 ( .A1(n10824), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10823), .ZN(n10827) );
  INV_X2 U11506 ( .A(n20103), .ZN(n20132) );
  BUF_X2 U11507 ( .A(n11954), .Z(n12243) );
  NAND2_X1 U11508 ( .A1(n10033), .A2(n10032), .ZN(n16970) );
  CLKBUF_X1 U11509 ( .A(n11233), .Z(n11419) );
  INV_X2 U11510 ( .A(n18760), .ZN(n18823) );
  INV_X1 U11511 ( .A(n10096), .ZN(n9819) );
  BUF_X2 U11512 ( .A(n13697), .Z(n17174) );
  BUF_X2 U11513 ( .A(n15713), .Z(n17179) );
  AND2_X2 U11514 ( .A1(n12729), .A2(n20627), .ZN(n20158) );
  BUF_X2 U11515 ( .A(n12249), .Z(n12286) );
  BUF_X2 U11516 ( .A(n11752), .Z(n12296) );
  AND2_X1 U11517 ( .A1(n9844), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10442) );
  NAND2_X2 U11518 ( .A1(n18897), .A2(n18761), .ZN(n18815) );
  BUF_X2 U11519 ( .A(n13734), .Z(n17145) );
  AND2_X2 U11520 ( .A1(n11500), .A2(n13093), .ZN(n12244) );
  INV_X2 U11521 ( .A(n16548), .ZN(n16550) );
  INV_X1 U11522 ( .A(n16944), .ZN(n10033) );
  BUF_X4 U11523 ( .A(n15710), .Z(n9820) );
  OR2_X1 U11524 ( .A1(n13645), .A2(n13646), .ZN(n9883) );
  NAND4_X1 U11525 ( .A1(n10132), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A3(
        n10128), .A4(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17787) );
  INV_X2 U11526 ( .A(n20909), .ZN(n20876) );
  CLKBUF_X1 U11527 ( .A(n13091), .Z(n12112) );
  NOR2_X2 U11528 ( .A1(n18701), .A2(n18356), .ZN(n18409) );
  BUF_X2 U11530 ( .A(n11591), .Z(n12128) );
  BUF_X2 U11531 ( .A(n10846), .Z(n10473) );
  AND2_X2 U11532 ( .A1(n11506), .A2(n14735), .ZN(n12249) );
  OR2_X2 U11533 ( .A1(n18704), .A2(n13646), .ZN(n9871) );
  AND2_X1 U11534 ( .A1(n10273), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11506) );
  INV_X1 U11535 ( .A(n13646), .ZN(n10032) );
  AND2_X1 U11536 ( .A1(n12844), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11494) );
  NAND2_X1 U11537 ( .A1(n18861), .A2(n18869), .ZN(n16944) );
  CLKBUF_X1 U11538 ( .A(n11844), .Z(n12307) );
  AND2_X1 U11539 ( .A1(n11489), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11495) );
  AND2_X2 U11540 ( .A1(n12863), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9836) );
  AND2_X1 U11541 ( .A1(n10426), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15532) );
  AND2_X1 U11542 ( .A1(n12863), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9835) );
  AND2_X2 U11543 ( .A1(n15543), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10846) );
  AND2_X2 U11544 ( .A1(n10427), .A2(n15533), .ZN(n10845) );
  INV_X1 U11545 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16329) );
  AND2_X1 U11546 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12862) );
  AND2_X1 U11547 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12863) );
  NAND2_X1 U11548 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18704) );
  INV_X1 U11549 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18841) );
  INV_X1 U11551 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15533) );
  NOR2_X1 U11552 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11508) );
  AND2_X1 U11553 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13094) );
  AND2_X2 U11554 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14735) );
  OR2_X1 U11555 ( .A1(n10911), .A2(n10899), .ZN(n11461) );
  INV_X2 U11556 ( .A(n10899), .ZN(n11101) );
  AND2_X1 U11557 ( .A1(n12669), .A2(n10927), .ZN(n10950) );
  NAND2_X1 U11558 ( .A1(n9951), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9966) );
  NAND2_X2 U11559 ( .A1(n13216), .A2(n10915), .ZN(n10906) );
  NAND2_X1 U11560 ( .A1(n10901), .A2(n10900), .ZN(n9821) );
  NAND2_X1 U11561 ( .A1(n9827), .A2(n9977), .ZN(n10949) );
  NAND2_X1 U11562 ( .A1(n9966), .A2(n10955), .ZN(n9823) );
  NOR2_X2 U11563 ( .A1(n15450), .A2(n15452), .ZN(n15451) );
  NAND2_X1 U11564 ( .A1(n9966), .A2(n10955), .ZN(n10965) );
  NAND2_X1 U11565 ( .A1(n10110), .A2(n9824), .ZN(n15022) );
  AND2_X1 U11566 ( .A1(n10964), .A2(n10963), .ZN(n9825) );
  NOR2_X1 U11567 ( .A1(n10919), .A2(n10918), .ZN(n9826) );
  AND2_X1 U11568 ( .A1(n13186), .A2(n13189), .ZN(n13368) );
  AND2_X2 U11569 ( .A1(n12820), .A2(n13435), .ZN(n14067) );
  AND2_X1 U11570 ( .A1(n16588), .A2(n9926), .ZN(n16388) );
  INV_X2 U11571 ( .A(n10118), .ZN(n16911) );
  NAND2_X2 U11572 ( .A1(n10036), .A2(n13932), .ZN(n13396) );
  NAND2_X1 U11574 ( .A1(n9979), .A2(n9978), .ZN(n9827) );
  INV_X1 U11575 ( .A(n13313), .ZN(n9828) );
  CLKBUF_X1 U11576 ( .A(n13188), .Z(n9829) );
  OR2_X1 U11577 ( .A1(n9832), .A2(n15234), .ZN(n9831) );
  INV_X1 U11578 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n9832) );
  OAI211_X1 U11579 ( .C1(n13608), .C2(n13974), .A(n10321), .B(n13931), .ZN(
        n9833) );
  XNOR2_X1 U11580 ( .A(n9834), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13995) );
  NOR2_X1 U11581 ( .A1(n9830), .A2(n9831), .ZN(n9834) );
  OAI211_X1 U11582 ( .C1(n13608), .C2(n13974), .A(n10321), .B(n13931), .ZN(
        n15205) );
  AND2_X1 U11583 ( .A1(n12863), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12868) );
  AND2_X2 U11584 ( .A1(n13129), .A2(n11134), .ZN(n13173) );
  AOI21_X1 U11585 ( .B1(n9823), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10966), .ZN(n10973) );
  AND2_X1 U11586 ( .A1(n11115), .A2(n11118), .ZN(n15525) );
  INV_X2 U11587 ( .A(n11238), .ZN(n9844) );
  AND2_X2 U11588 ( .A1(n13186), .A2(n13198), .ZN(n13367) );
  INV_X1 U11589 ( .A(n10929), .ZN(n9979) );
  NAND2_X2 U11591 ( .A1(n15497), .A2(n9950), .ZN(n15175) );
  NAND2_X2 U11592 ( .A1(n13944), .A2(n13943), .ZN(n15497) );
  AND2_X1 U11593 ( .A1(n10427), .A2(n15533), .ZN(n9838) );
  AND2_X1 U11594 ( .A1(n10427), .A2(n15533), .ZN(n9842) );
  INV_X1 U11595 ( .A(n10433), .ZN(n9839) );
  NOR2_X1 U11597 ( .A1(n10042), .A2(n11058), .ZN(n15037) );
  INV_X2 U11598 ( .A(n10915), .ZN(n16347) );
  NAND2_X2 U11599 ( .A1(n10941), .A2(n10940), .ZN(n10961) );
  NAND2_X4 U11600 ( .A1(n10467), .A2(n10466), .ZN(n10930) );
  BUF_X2 U11601 ( .A(n13185), .Z(n13542) );
  AND2_X1 U11602 ( .A1(n10427), .A2(n15533), .ZN(n9841) );
  INV_X1 U11603 ( .A(n11238), .ZN(n9843) );
  INV_X1 U11604 ( .A(n11409), .ZN(n9845) );
  CLKBUF_X1 U11605 ( .A(n11699), .Z(n11713) );
  AND4_X1 U11606 ( .A1(n10622), .A2(n10621), .A3(n10620), .A4(n10619), .ZN(
        n10637) );
  OR2_X1 U11607 ( .A1(n11078), .A2(n13784), .ZN(n10971) );
  NAND2_X1 U11608 ( .A1(n10486), .A2(n9837), .ZN(n10748) );
  AND2_X1 U11609 ( .A1(n19247), .A2(n19938), .ZN(n10486) );
  NAND3_X1 U11610 ( .A1(n10902), .A2(n10930), .A3(n19252), .ZN(n10933) );
  NAND2_X1 U11611 ( .A1(n10438), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10439) );
  NAND2_X1 U11612 ( .A1(n10432), .A2(n10861), .ZN(n10440) );
  NAND2_X1 U11613 ( .A1(n11623), .A2(n13079), .ZN(n12763) );
  AND4_X1 U11614 ( .A1(n11606), .A2(n11605), .A3(n11604), .A4(n11603), .ZN(
        n11618) );
  AND2_X1 U11615 ( .A1(n14003), .A2(n14012), .ZN(n12765) );
  AND4_X1 U11616 ( .A1(n11504), .A2(n11503), .A3(n11502), .A4(n11501), .ZN(
        n11514) );
  NAND2_X1 U11617 ( .A1(n10185), .A2(n10184), .ZN(n10183) );
  INV_X1 U11618 ( .A(n17578), .ZN(n10184) );
  CLKBUF_X1 U11619 ( .A(n11938), .Z(n11987) );
  CLKBUF_X1 U11620 ( .A(n11954), .Z(n11939) );
  OR2_X1 U11621 ( .A1(n11689), .A2(n11688), .ZN(n12811) );
  NAND2_X1 U11622 ( .A1(n20231), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11750) );
  AND3_X1 U11623 ( .A1(n12792), .A2(n12820), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12355) );
  AND2_X1 U11624 ( .A1(n11631), .A2(n11647), .ZN(n12774) );
  NAND2_X1 U11625 ( .A1(n9827), .A2(n12673), .ZN(n10931) );
  NAND2_X1 U11626 ( .A1(n10912), .A2(n10911), .ZN(n10929) );
  NAND2_X1 U11627 ( .A1(n9826), .A2(n10962), .ZN(n10963) );
  NAND2_X1 U11628 ( .A1(n11639), .A2(n11638), .ZN(n11702) );
  AND4_X1 U11629 ( .A1(n11532), .A2(n11531), .A3(n11530), .A4(n11529), .ZN(
        n11533) );
  NOR2_X1 U11630 ( .A1(n11623), .A2(n20898), .ZN(n11996) );
  OAI21_X1 U11631 ( .B1(n10232), .B2(n10137), .A(n10227), .ZN(n10136) );
  NAND2_X1 U11632 ( .A1(n10228), .A2(n14519), .ZN(n10227) );
  NAND2_X1 U11633 ( .A1(n14519), .A2(n10138), .ZN(n10137) );
  INV_X1 U11634 ( .A(n10230), .ZN(n10228) );
  OR2_X1 U11635 ( .A1(n11865), .A2(n11864), .ZN(n13497) );
  AND4_X1 U11636 ( .A1(n11552), .A2(n11551), .A3(n11550), .A4(n11549), .ZN(
        n11553) );
  AND2_X1 U11637 ( .A1(n11702), .A2(n11701), .ZN(n11703) );
  OR2_X1 U11638 ( .A1(n11694), .A2(n11693), .ZN(n11709) );
  NAND2_X1 U11639 ( .A1(n20263), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11751) );
  OR2_X1 U11640 ( .A1(n11713), .A2(n11712), .ZN(n11726) );
  AOI21_X1 U11641 ( .B1(n11274), .B2(n10331), .A(n9938), .ZN(n10330) );
  NAND2_X1 U11642 ( .A1(n14873), .A2(n10331), .ZN(n10329) );
  NAND2_X1 U11643 ( .A1(n11102), .A2(n11101), .ZN(n11337) );
  AND2_X1 U11644 ( .A1(n13216), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11102) );
  NAND2_X1 U11645 ( .A1(n9837), .A2(n13816), .ZN(n13906) );
  AOI21_X1 U11646 ( .B1(n10106), .B2(n10103), .A(n10102), .ZN(n10101) );
  INV_X1 U11647 ( .A(n15183), .ZN(n10102) );
  AND3_X1 U11648 ( .A1(n10629), .A2(n10628), .A3(n10627), .ZN(n10635) );
  AND4_X1 U11649 ( .A1(n10633), .A2(n10632), .A3(n10631), .A4(n10630), .ZN(
        n10634) );
  AND4_X1 U11650 ( .A1(n10626), .A2(n10625), .A3(n10624), .A4(n10623), .ZN(
        n10636) );
  INV_X1 U11651 ( .A(n13932), .ZN(n13935) );
  INV_X1 U11652 ( .A(n10550), .ZN(n10235) );
  AND2_X1 U11653 ( .A1(n19247), .A2(n19267), .ZN(n10468) );
  NAND2_X1 U11654 ( .A1(n11097), .A2(n19938), .ZN(n11124) );
  NAND2_X1 U11655 ( .A1(n13542), .A2(n9910), .ZN(n9968) );
  NOR2_X1 U11656 ( .A1(n13645), .A2(n13644), .ZN(n13698) );
  NOR2_X1 U11657 ( .A1(n17390), .A2(n15760), .ZN(n15742) );
  INV_X1 U11658 ( .A(n13760), .ZN(n13769) );
  AOI21_X1 U11659 ( .B1(n18670), .B2(n9917), .A(n13776), .ZN(n15914) );
  INV_X1 U11660 ( .A(n14003), .ZN(n14007) );
  AND2_X1 U11661 ( .A1(n14000), .A2(n14007), .ZN(n12840) );
  NAND2_X2 U11662 ( .A1(n11633), .A2(n12820), .ZN(n15872) );
  INV_X1 U11663 ( .A(n11978), .ZN(n12308) );
  NAND2_X1 U11664 ( .A1(n10056), .A2(n13482), .ZN(n16035) );
  NAND2_X1 U11665 ( .A1(n11851), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11859) );
  INV_X2 U11666 ( .A(n15910), .ZN(n14082) );
  OAI21_X1 U11667 ( .B1(n14686), .B2(n14424), .A(n16024), .ZN(n15984) );
  NAND2_X1 U11668 ( .A1(n12767), .A2(n12766), .ZN(n12795) );
  OR2_X1 U11669 ( .A1(n19972), .A2(n12483), .ZN(n12497) );
  OR2_X1 U11670 ( .A1(n10145), .A2(n15062), .ZN(n10144) );
  OR2_X1 U11671 ( .A1(n12427), .A2(n10145), .ZN(n10143) );
  OAI21_X1 U11673 ( .B1(n13185), .B2(n9976), .A(n9910), .ZN(n11130) );
  INV_X1 U11674 ( .A(n11363), .ZN(n10349) );
  AND2_X1 U11675 ( .A1(n12418), .A2(n9941), .ZN(n14862) );
  INV_X1 U11676 ( .A(n14859), .ZN(n10204) );
  INV_X1 U11677 ( .A(n15117), .ZN(n9987) );
  NAND2_X1 U11678 ( .A1(n15169), .A2(n9847), .ZN(n10240) );
  NAND2_X1 U11679 ( .A1(n13401), .A2(n10616), .ZN(n13617) );
  INV_X1 U11680 ( .A(n13168), .ZN(n10238) );
  NAND2_X1 U11681 ( .A1(n10465), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10466) );
  NAND2_X1 U11682 ( .A1(n10460), .A2(n10861), .ZN(n10467) );
  INV_X1 U11683 ( .A(n18258), .ZN(n17271) );
  NAND2_X1 U11684 ( .A1(n10182), .A2(n10181), .ZN(n10180) );
  NAND2_X1 U11685 ( .A1(n17541), .A2(n17798), .ZN(n10182) );
  AND2_X1 U11686 ( .A1(n10180), .A2(n10179), .ZN(n17530) );
  NAND2_X1 U11687 ( .A1(n15742), .A2(n17815), .ZN(n16440) );
  NAND2_X1 U11688 ( .A1(n16436), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17541) );
  AND2_X1 U11689 ( .A1(n15777), .A2(n17581), .ZN(n10031) );
  INV_X1 U11690 ( .A(n16326), .ZN(n16301) );
  NAND2_X1 U11691 ( .A1(n13189), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n9954) );
  NAND2_X1 U11692 ( .A1(n13198), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n9955) );
  AOI21_X1 U11693 ( .B1(n9821), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10939), 
        .ZN(n10940) );
  NAND2_X1 U11694 ( .A1(n12319), .A2(n12318), .ZN(n12327) );
  CLKBUF_X1 U11695 ( .A(n12285), .Z(n12224) );
  NOR2_X1 U11696 ( .A1(n10084), .A2(n16078), .ZN(n10080) );
  NAND2_X1 U11697 ( .A1(n10135), .A2(n9918), .ZN(n11865) );
  INV_X1 U11698 ( .A(n12736), .ZN(n12775) );
  INV_X1 U11699 ( .A(n12812), .ZN(n11679) );
  OR2_X1 U11700 ( .A1(n11664), .A2(n11663), .ZN(n13487) );
  OR2_X1 U11701 ( .A1(n11762), .A2(n11761), .ZN(n13337) );
  INV_X1 U11702 ( .A(n10844), .ZN(n11416) );
  NAND2_X1 U11703 ( .A1(n10928), .A2(n10905), .ZN(n9993) );
  INV_X1 U11704 ( .A(n10905), .ZN(n12644) );
  AOI21_X1 U11705 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19935), .A(
        n10867), .ZN(n10870) );
  NOR2_X1 U11706 ( .A1(n17397), .A2(n15818), .ZN(n15743) );
  NOR2_X1 U11707 ( .A1(n12775), .A2(n12820), .ZN(n11628) );
  NOR2_X1 U11708 ( .A1(n10314), .A2(n10312), .ZN(n10311) );
  INV_X1 U11709 ( .A(n14097), .ZN(n10314) );
  OR2_X1 U11710 ( .A1(n14110), .A2(n10313), .ZN(n10312) );
  INV_X1 U11711 ( .A(n14121), .ZN(n10313) );
  NOR2_X1 U11712 ( .A1(n14176), .A2(n10318), .ZN(n10317) );
  INV_X1 U11713 ( .A(n14356), .ZN(n10318) );
  INV_X1 U11714 ( .A(n12311), .ZN(n12277) );
  NOR2_X1 U11715 ( .A1(n10305), .A2(n14307), .ZN(n10304) );
  INV_X1 U11716 ( .A(n14200), .ZN(n10305) );
  NAND2_X1 U11717 ( .A1(n20210), .A2(n12954), .ZN(n13060) );
  NAND2_X1 U11718 ( .A1(n10085), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10084) );
  NAND2_X1 U11719 ( .A1(n16012), .A2(n14422), .ZN(n10085) );
  OR2_X1 U11720 ( .A1(n14520), .A2(n14423), .ZN(n14686) );
  NOR2_X1 U11721 ( .A1(n9896), .A2(n10231), .ZN(n10230) );
  NOR2_X1 U11722 ( .A1(n16012), .A2(n14421), .ZN(n10231) );
  AND2_X1 U11723 ( .A1(n14541), .A2(n14543), .ZN(n14526) );
  NAND2_X1 U11724 ( .A1(n14567), .A2(n14412), .ZN(n14524) );
  NAND2_X1 U11725 ( .A1(n10075), .A2(n13494), .ZN(n10071) );
  INV_X1 U11726 ( .A(n14062), .ZN(n14041) );
  INV_X1 U11727 ( .A(n12579), .ZN(n12755) );
  NOR2_X1 U11728 ( .A1(n13920), .A2(n13918), .ZN(n13923) );
  INV_X1 U11729 ( .A(n10884), .ZN(n13376) );
  NOR2_X1 U11730 ( .A1(n10353), .A2(n10352), .ZN(n10351) );
  OR2_X1 U11731 ( .A1(n11362), .A2(n14844), .ZN(n10350) );
  INV_X1 U11732 ( .A(n12420), .ZN(n10270) );
  INV_X1 U11733 ( .A(n14913), .ZN(n10333) );
  INV_X1 U11734 ( .A(n12462), .ZN(n10206) );
  NOR2_X1 U11735 ( .A1(n19042), .A2(n10151), .ZN(n10150) );
  NAND2_X1 U11736 ( .A1(n10915), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11431) );
  INV_X1 U11737 ( .A(n10009), .ZN(n10008) );
  OAI21_X1 U11738 ( .B1(n13915), .B2(n9869), .A(n13921), .ZN(n10009) );
  INV_X1 U11739 ( .A(n15047), .ZN(n13913) );
  NAND2_X1 U11740 ( .A1(n13911), .A2(n9855), .ZN(n13917) );
  NOR2_X1 U11741 ( .A1(n14786), .A2(n10272), .ZN(n10271) );
  INV_X1 U11742 ( .A(n15340), .ZN(n10272) );
  AOI21_X1 U11743 ( .B1(n9986), .B2(n15149), .A(n9985), .ZN(n9984) );
  INV_X1 U11744 ( .A(n15101), .ZN(n9985) );
  NAND2_X1 U11745 ( .A1(n10241), .A2(n15148), .ZN(n9986) );
  INV_X1 U11746 ( .A(n15182), .ZN(n10107) );
  NAND2_X1 U11747 ( .A1(n10197), .A2(n10196), .ZN(n10195) );
  INV_X1 U11748 ( .A(n13035), .ZN(n10196) );
  INV_X1 U11749 ( .A(n10199), .ZN(n10197) );
  OR2_X1 U11750 ( .A1(n16279), .A2(n16275), .ZN(n10257) );
  NOR2_X1 U11751 ( .A1(n16298), .A2(n10261), .ZN(n10260) );
  INV_X1 U11752 ( .A(n15513), .ZN(n10261) );
  NAND2_X1 U11753 ( .A1(n10487), .A2(n10768), .ZN(n10503) );
  AND2_X1 U11754 ( .A1(n10930), .A2(n19938), .ZN(n10522) );
  AND2_X1 U11755 ( .A1(n16347), .A2(n10912), .ZN(n10856) );
  NAND2_X1 U11756 ( .A1(n13191), .A2(n16315), .ZN(n13202) );
  INV_X1 U11757 ( .A(n19949), .ZN(n19375) );
  NAND2_X1 U11758 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13646) );
  NAND2_X1 U11759 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18861), .ZN(
        n13647) );
  NOR2_X1 U11760 ( .A1(n18704), .A2(n13644), .ZN(n13697) );
  NOR2_X1 U11761 ( .A1(n13647), .A2(n13644), .ZN(n15603) );
  NOR2_X1 U11762 ( .A1(n18268), .A2(n18248), .ZN(n15802) );
  NAND2_X1 U11763 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n10121) );
  OAI21_X1 U11764 ( .B1(n16611), .B2(n10122), .A(n10123), .ZN(n10120) );
  NOR2_X1 U11765 ( .A1(n17680), .A2(n18013), .ZN(n17622) );
  AND2_X1 U11766 ( .A1(n10054), .A2(n10052), .ZN(n13773) );
  NOR2_X1 U11767 ( .A1(n10055), .A2(n13752), .ZN(n10054) );
  AOI21_X1 U11768 ( .B1(n13753), .B2(n18237), .A(n10053), .ZN(n10052) );
  AOI22_X1 U11769 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13662) );
  NAND2_X1 U11770 ( .A1(n11637), .A2(n11633), .ZN(n14010) );
  OR2_X1 U11771 ( .A1(n11723), .A2(n11724), .ZN(n11721) );
  INV_X1 U11772 ( .A(n20059), .ZN(n20019) );
  NAND2_X1 U11773 ( .A1(n10288), .A2(n14067), .ZN(n10287) );
  INV_X1 U11774 ( .A(n12926), .ZN(n10288) );
  XNOR2_X1 U11775 ( .A(n11702), .B(n11653), .ZN(n11838) );
  AND4_X1 U11776 ( .A1(n11528), .A2(n11527), .A3(n11526), .A4(n11525), .ZN(
        n11534) );
  AND4_X1 U11777 ( .A1(n11524), .A2(n11523), .A3(n11522), .A4(n11521), .ZN(
        n11535) );
  AND4_X1 U11778 ( .A1(n11520), .A2(n11519), .A3(n11518), .A4(n11517), .ZN(
        n11536) );
  INV_X1 U11779 ( .A(n14227), .ZN(n11984) );
  AND2_X1 U11780 ( .A1(n11966), .A2(n10307), .ZN(n10306) );
  OR2_X1 U11781 ( .A1(n14238), .A2(n14403), .ZN(n10307) );
  NAND2_X1 U11782 ( .A1(n11857), .A2(n11856), .ZN(n10290) );
  NAND2_X1 U11783 ( .A1(n11820), .A2(n11819), .ZN(n13075) );
  NAND2_X1 U11784 ( .A1(n14046), .A2(n14082), .ZN(n14071) );
  NAND2_X1 U11785 ( .A1(n14452), .A2(n9893), .ZN(n14435) );
  OR2_X1 U11786 ( .A1(n10014), .A2(n10013), .ZN(n9850) );
  INV_X1 U11787 ( .A(n10015), .ZN(n10013) );
  INV_X1 U11788 ( .A(n14452), .ZN(n10014) );
  NAND2_X1 U11789 ( .A1(n14437), .A2(n16012), .ZN(n10215) );
  NAND2_X1 U11790 ( .A1(n16035), .A2(n10219), .ZN(n10223) );
  INV_X1 U11791 ( .A(n13493), .ZN(n10220) );
  INV_X1 U11792 ( .A(n10222), .ZN(n10221) );
  NAND2_X1 U11793 ( .A1(n16036), .A2(n13493), .ZN(n10224) );
  INV_X1 U11794 ( .A(n13334), .ZN(n10211) );
  INV_X1 U11795 ( .A(n16049), .ZN(n10208) );
  NOR2_X1 U11796 ( .A1(n12781), .A2(n12779), .ZN(n14000) );
  NAND2_X1 U11797 ( .A1(n12743), .A2(n12742), .ZN(n12744) );
  OR2_X1 U11798 ( .A1(n12739), .A2(n13064), .ZN(n12743) );
  NAND2_X1 U11799 ( .A1(n10217), .A2(n11707), .ZN(n12810) );
  NAND2_X1 U11800 ( .A1(n10218), .A2(n20297), .ZN(n10217) );
  AND2_X1 U11801 ( .A1(n11728), .A2(n20902), .ZN(n10218) );
  NAND2_X1 U11802 ( .A1(n11709), .A2(n11695), .ZN(n11827) );
  NAND2_X1 U11803 ( .A1(n11829), .A2(n11709), .ZN(n11822) );
  INV_X1 U11804 ( .A(n20534), .ZN(n20692) );
  NOR2_X1 U11805 ( .A1(n20395), .A2(n20633), .ZN(n20563) );
  NOR2_X1 U11806 ( .A1(n20561), .A2(n20395), .ZN(n20729) );
  INV_X1 U11807 ( .A(n20556), .ZN(n20719) );
  NAND2_X1 U11808 ( .A1(n20902), .A2(n20230), .ZN(n20395) );
  OR2_X1 U11809 ( .A1(n12352), .A2(n12323), .ZN(n12365) );
  NOR2_X1 U11810 ( .A1(n12768), .A2(n14007), .ZN(n15867) );
  AND2_X1 U11811 ( .A1(n10143), .A2(n9864), .ZN(n16213) );
  NAND2_X1 U11812 ( .A1(n13911), .A2(n13910), .ZN(n16207) );
  NAND2_X1 U11813 ( .A1(n10892), .A2(n10092), .ZN(n16221) );
  AND2_X1 U11814 ( .A1(n9868), .A2(n16222), .ZN(n10092) );
  NOR2_X1 U11815 ( .A1(n12455), .A2(n10095), .ZN(n10094) );
  OAI21_X1 U11816 ( .B1(n10145), .B2(n15092), .A(n10390), .ZN(n10156) );
  AOI21_X1 U11817 ( .B1(n11032), .B2(P2_EBX_REG_0__SCAN_IN), .A(n10956), .ZN(
        n10957) );
  NAND2_X1 U11818 ( .A1(n10335), .A2(n9920), .ZN(n13038) );
  XNOR2_X1 U11819 ( .A(n11319), .B(n11317), .ZN(n14855) );
  NAND2_X1 U11820 ( .A1(n10341), .A2(n11296), .ZN(n10340) );
  NAND2_X1 U11821 ( .A1(n10338), .A2(n10345), .ZN(n10339) );
  AND2_X1 U11822 ( .A1(n19160), .A2(n11482), .ZN(n12630) );
  INV_X1 U11823 ( .A(n11431), .ZN(n14747) );
  XNOR2_X1 U11824 ( .A(n10377), .B(n10376), .ZN(n13992) );
  OR2_X1 U11825 ( .A1(n14902), .A2(n14895), .ZN(n14897) );
  AND2_X1 U11826 ( .A1(n11050), .A2(n11049), .ZN(n14886) );
  AND2_X1 U11827 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10406) );
  INV_X1 U11828 ( .A(n13951), .ZN(n10201) );
  NAND2_X1 U11829 ( .A1(n10004), .A2(n10002), .ZN(n14997) );
  AOI21_X1 U11830 ( .B1(n10006), .B2(n10005), .A(n10003), .ZN(n10002) );
  NAND2_X1 U11831 ( .A1(n15021), .A2(n10005), .ZN(n10004) );
  INV_X1 U11832 ( .A(n15010), .ZN(n10003) );
  NOR2_X2 U11833 ( .A1(n9830), .A2(n15234), .ZN(n15014) );
  AND2_X1 U11834 ( .A1(n15381), .A2(n16316), .ZN(n15473) );
  OR3_X1 U11835 ( .A1(n13900), .A2(n13941), .A3(n13899), .ZN(n15088) );
  NAND2_X1 U11836 ( .A1(n15468), .A2(n10099), .ZN(n10001) );
  OR2_X1 U11837 ( .A1(n15362), .A2(n13970), .ZN(n15325) );
  NAND2_X1 U11838 ( .A1(n10038), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10037) );
  INV_X1 U11839 ( .A(n10039), .ZN(n10038) );
  NAND2_X1 U11840 ( .A1(n10263), .A2(n13468), .ZN(n10262) );
  INV_X1 U11841 ( .A(n15393), .ZN(n10263) );
  AOI21_X1 U11842 ( .B1(n9847), .B2(n10243), .A(n10242), .ZN(n10241) );
  INV_X1 U11843 ( .A(n15099), .ZN(n10242) );
  INV_X1 U11844 ( .A(n10246), .ZN(n10243) );
  NOR2_X1 U11845 ( .A1(n15174), .A2(n10247), .ZN(n10246) );
  INV_X1 U11846 ( .A(n15405), .ZN(n10247) );
  NAND2_X2 U11847 ( .A1(n9964), .A2(n10251), .ZN(n15468) );
  AND2_X1 U11848 ( .A1(n10252), .A2(n13834), .ZN(n10251) );
  NAND2_X1 U11849 ( .A1(n15208), .A2(n10253), .ZN(n9964) );
  AND2_X1 U11850 ( .A1(n15193), .A2(n15505), .ZN(n13834) );
  AND3_X1 U11851 ( .A1(n10686), .A2(n10685), .A3(n10684), .ZN(n15483) );
  NAND2_X1 U11852 ( .A1(n10234), .A2(n9897), .ZN(n13401) );
  NOR2_X1 U11853 ( .A1(n10237), .A2(n10239), .ZN(n10233) );
  NAND2_X1 U11854 ( .A1(n13306), .A2(n13305), .ZN(n9991) );
  AND3_X1 U11855 ( .A1(n10586), .A2(n10585), .A3(n10584), .ZN(n13168) );
  NAND2_X1 U11856 ( .A1(n9990), .A2(n13619), .ZN(n13307) );
  NAND2_X1 U11857 ( .A1(n11120), .A2(n11119), .ZN(n11127) );
  NAND2_X1 U11858 ( .A1(n15525), .A2(n12597), .ZN(n11120) );
  AOI21_X1 U11859 ( .B1(n13191), .B2(n12597), .A(n11126), .ZN(n12623) );
  OR2_X1 U11860 ( .A1(n9976), .A2(n11114), .ZN(n9974) );
  AOI21_X1 U11861 ( .B1(n9910), .B2(n9976), .A(n9971), .ZN(n9970) );
  OR2_X1 U11862 ( .A1(n19936), .A2(n19375), .ZN(n19414) );
  OR2_X1 U11863 ( .A1(n19936), .A2(n19949), .ZN(n13156) );
  NOR2_X2 U11864 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19923) );
  AND2_X1 U11865 ( .A1(n19936), .A2(n19375), .ZN(n19922) );
  NAND2_X2 U11866 ( .A1(n10822), .A2(n10821), .ZN(n19252) );
  NAND4_X1 U11867 ( .A1(n10818), .A2(n9885), .A3(n10819), .A4(n10820), .ZN(
        n10821) );
  NAND2_X1 U11868 ( .A1(n10365), .A2(n10361), .ZN(n10822) );
  INV_X1 U11869 ( .A(n19414), .ZN(n19669) );
  INV_X1 U11870 ( .A(n19758), .ZN(n19665) );
  NOR2_X1 U11871 ( .A1(n19522), .A2(n19958), .ZN(n19670) );
  NOR2_X2 U11872 ( .A1(n13155), .A2(n13154), .ZN(n19273) );
  NOR2_X2 U11873 ( .A1(n13153), .A2(n13154), .ZN(n19274) );
  NOR2_X1 U11874 ( .A1(n18244), .A2(n13759), .ZN(n13774) );
  OAI21_X1 U11875 ( .B1(n13766), .B2(n15786), .A(n13765), .ZN(n18673) );
  AOI21_X1 U11876 ( .B1(n17597), .B2(n16733), .A(n16911), .ZN(n16708) );
  INV_X1 U11877 ( .A(n9873), .ZN(n17188) );
  NOR2_X1 U11878 ( .A1(n13648), .A2(n13647), .ZN(n15710) );
  OAI21_X1 U11879 ( .B1(n15914), .B2(n15913), .A(n18882), .ZN(n15915) );
  INV_X1 U11880 ( .A(n17671), .ZN(n15771) );
  INV_X1 U11881 ( .A(n15778), .ZN(n17680) );
  INV_X1 U11882 ( .A(n17382), .ZN(n16392) );
  INV_X1 U11883 ( .A(n10025), .ZN(n10022) );
  XNOR2_X1 U11884 ( .A(n15744), .B(n18171), .ZN(n17854) );
  NAND2_X1 U11885 ( .A1(n10023), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10019) );
  INV_X1 U11886 ( .A(n17865), .ZN(n10023) );
  NOR2_X1 U11887 ( .A1(n16578), .A2(n18132), .ZN(n18037) );
  NAND2_X1 U11888 ( .A1(n13761), .A2(n18671), .ZN(n15806) );
  NOR2_X2 U11889 ( .A1(n13729), .A2(n13728), .ZN(n18263) );
  NAND2_X1 U11890 ( .A1(n9997), .A2(n13379), .ZN(n10036) );
  INV_X1 U11891 ( .A(n20075), .ZN(n20064) );
  AND2_X1 U11892 ( .A1(n13021), .A2(n20241), .ZN(n20147) );
  AND2_X1 U11893 ( .A1(n16041), .A2(n12808), .ZN(n16037) );
  AND2_X1 U11894 ( .A1(n15867), .A2(n14012), .ZN(n20159) );
  XNOR2_X1 U11895 ( .A(n14456), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14633) );
  XNOR2_X1 U11896 ( .A(n10066), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14636) );
  NAND2_X1 U11897 ( .A1(n10068), .A2(n10067), .ZN(n10066) );
  OR2_X1 U11898 ( .A1(n14465), .A2(n16024), .ZN(n10067) );
  NAND2_X1 U11899 ( .A1(n14466), .A2(n16024), .ZN(n10068) );
  AND2_X1 U11900 ( .A1(n12795), .A2(n12771), .ZN(n20208) );
  OR2_X1 U11901 ( .A1(n12738), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20207) );
  NAND2_X1 U11902 ( .A1(n20297), .A2(n11728), .ZN(n20558) );
  NAND2_X1 U11903 ( .A1(n12647), .A2(n12498), .ZN(n12596) );
  NOR2_X1 U11904 ( .A1(n15072), .A2(n12428), .ZN(n12427) );
  AND2_X1 U11905 ( .A1(n14906), .A2(n10930), .ZN(n14901) );
  INV_X2 U11906 ( .A(n14906), .ZN(n14919) );
  AND2_X2 U11907 ( .A1(n12401), .A2(n16362), .ZN(n14906) );
  NAND2_X1 U11908 ( .A1(n14828), .A2(n11405), .ZN(n11428) );
  NAND2_X1 U11909 ( .A1(n14833), .A2(n10354), .ZN(n14843) );
  NAND2_X1 U11910 ( .A1(n11363), .A2(n11362), .ZN(n10354) );
  NAND2_X1 U11911 ( .A1(n19160), .A2(n11481), .ZN(n14988) );
  OR2_X1 U11912 ( .A1(n12881), .A2(n11470), .ZN(n11471) );
  INV_X1 U11913 ( .A(n19958), .ZN(n19488) );
  XNOR2_X1 U11914 ( .A(n14768), .B(n13951), .ZN(n15223) );
  OR2_X1 U11915 ( .A1(n14838), .A2(n12444), .ZN(n15260) );
  NAND2_X1 U11916 ( .A1(n15116), .A2(n10250), .ZN(n10249) );
  OR2_X1 U11917 ( .A1(n12681), .A2(n12666), .ZN(n16326) );
  OR2_X1 U11918 ( .A1(n12681), .A2(n12662), .ZN(n16314) );
  INV_X1 U11919 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19938) );
  INV_X1 U11920 ( .A(n19923), .ZN(n19931) );
  NAND2_X1 U11921 ( .A1(n15916), .A2(n17406), .ZN(n17405) );
  NAND2_X1 U11922 ( .A1(n17351), .A2(n17264), .ZN(n17400) );
  INV_X1 U11923 ( .A(n17383), .ZN(n17411) );
  INV_X1 U11924 ( .A(n17400), .ZN(n17406) );
  INV_X1 U11925 ( .A(n15915), .ZN(n17264) );
  INV_X1 U11926 ( .A(n17405), .ZN(n17409) );
  OR2_X1 U11927 ( .A1(n17532), .A2(n10175), .ZN(n10174) );
  AND2_X1 U11928 ( .A1(n17610), .A2(n17533), .ZN(n10175) );
  INV_X1 U11929 ( .A(n10177), .ZN(n10176) );
  OAI21_X1 U11930 ( .B1(n10180), .B2(n10179), .A(n17799), .ZN(n10177) );
  INV_X1 U11931 ( .A(n17530), .ZN(n10178) );
  INV_X1 U11932 ( .A(n17728), .ZN(n17735) );
  NAND2_X1 U11933 ( .A1(n16449), .A2(n16448), .ZN(n16457) );
  INV_X1 U11934 ( .A(n16447), .ZN(n16449) );
  OAI21_X1 U11935 ( .B1(n17530), .B2(n16446), .A(n16445), .ZN(n16447) );
  INV_X1 U11936 ( .A(n16436), .ZN(n15782) );
  NAND2_X1 U11937 ( .A1(n13601), .A2(n13600), .ZN(n13933) );
  OR2_X1 U11938 ( .A1(n13597), .A2(n13596), .ZN(n13601) );
  NOR2_X1 U11939 ( .A1(n15538), .A2(n18909), .ZN(n9980) );
  AOI22_X1 U11940 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20271), .B1(n13435), 
        .B2(n12334), .ZN(n12340) );
  OR2_X1 U11941 ( .A1(n10543), .A2(n10542), .ZN(n10881) );
  NOR2_X1 U11942 ( .A1(n10865), .A2(n10864), .ZN(n10867) );
  OR2_X1 U11943 ( .A1(n13683), .A2(n13684), .ZN(n13676) );
  NAND2_X1 U11944 ( .A1(n12757), .A2(n14730), .ZN(n11641) );
  INV_X1 U11945 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11489) );
  NOR2_X1 U11946 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11844) );
  NOR2_X1 U11947 ( .A1(n10073), .A2(n13064), .ZN(n10070) );
  NOR2_X1 U11948 ( .A1(n9915), .A2(n10074), .ZN(n10073) );
  NAND2_X1 U11949 ( .A1(n10076), .A2(n10078), .ZN(n10075) );
  OR2_X1 U11950 ( .A1(n11776), .A2(n11775), .ZN(n13336) );
  INV_X1 U11951 ( .A(n11835), .ZN(n10296) );
  INV_X1 U11952 ( .A(n20902), .ZN(n10297) );
  NAND2_X1 U11953 ( .A1(n11741), .A2(n10061), .ZN(n10060) );
  INV_X1 U11954 ( .A(n11750), .ZN(n11741) );
  OR2_X1 U11955 ( .A1(n11739), .A2(n11738), .ZN(n11740) );
  AOI21_X1 U11956 ( .B1(n12327), .B2(n12326), .A(n12320), .ZN(n12325) );
  NOR2_X1 U11957 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n12321), .ZN(
        n12324) );
  NAND2_X1 U11958 ( .A1(n10096), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11328) );
  NAND2_X1 U11959 ( .A1(n10096), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11321) );
  AOI21_X1 U11960 ( .B1(n11408), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n9946), .ZN(n11398) );
  NAND2_X1 U11961 ( .A1(n10096), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11351) );
  NAND2_X1 U11962 ( .A1(n10096), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11344) );
  INV_X1 U11963 ( .A(n14866), .ZN(n10331) );
  NAND2_X1 U11964 ( .A1(n10096), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11305) );
  NAND2_X1 U11965 ( .A1(n10096), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11298) );
  NAND2_X1 U11966 ( .A1(n10096), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11283) );
  NAND2_X1 U11967 ( .A1(n10096), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11276) );
  NAND2_X1 U11968 ( .A1(n10096), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11235) );
  NAND2_X1 U11969 ( .A1(n13367), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n9960) );
  NAND2_X1 U11970 ( .A1(n13205), .A2(n9894), .ZN(n9961) );
  NAND2_X1 U11971 ( .A1(n19566), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n9962) );
  NAND2_X1 U11972 ( .A1(n19242), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n9957) );
  NAND2_X1 U11973 ( .A1(n13365), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n9958) );
  AND2_X1 U11974 ( .A1(n13211), .A2(n13210), .ZN(n13215) );
  NOR2_X1 U11975 ( .A1(n19247), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10469) );
  INV_X1 U11976 ( .A(n10881), .ZN(n13262) );
  AND2_X1 U11977 ( .A1(n10929), .A2(n10930), .ZN(n9992) );
  AOI22_X1 U11978 ( .A1(n11233), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9844), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10803) );
  AOI22_X1 U11979 ( .A1(n9835), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9840), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10495) );
  INV_X1 U11980 ( .A(n11435), .ZN(n10857) );
  AOI22_X1 U11981 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10845), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10445) );
  NAND2_X1 U11982 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18869), .ZN(
        n13645) );
  NAND2_X1 U11983 ( .A1(n18851), .A2(n18841), .ZN(n13643) );
  NAND2_X1 U11984 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18851), .ZN(
        n13644) );
  NOR2_X1 U11985 ( .A1(n13751), .A2(n18253), .ZN(n10053) );
  AOI21_X1 U11986 ( .B1(n13760), .B2(n18244), .A(n13750), .ZN(n10055) );
  NAND2_X1 U11987 ( .A1(n16578), .A2(n18237), .ZN(n13760) );
  AOI22_X1 U11988 ( .A1(n9836), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9840), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10434) );
  NAND2_X1 U11989 ( .A1(n13091), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11526) );
  BUF_X1 U11990 ( .A(n11629), .Z(n13080) );
  NAND2_X1 U11991 ( .A1(n10077), .A2(n11858), .ZN(n10076) );
  INV_X1 U11992 ( .A(n11849), .ZN(n10077) );
  INV_X1 U11993 ( .A(n11858), .ZN(n10078) );
  NAND2_X1 U11994 ( .A1(n13092), .A2(n20271), .ZN(n12378) );
  NAND2_X1 U11995 ( .A1(n12285), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11613) );
  AND2_X1 U11996 ( .A1(n10316), .A2(n10317), .ZN(n10315) );
  INV_X1 U11997 ( .A(n14161), .ZN(n10316) );
  AOI21_X1 U11998 ( .B1(n14539), .B2(n14526), .A(n10139), .ZN(n14527) );
  NAND2_X1 U11999 ( .A1(n14694), .A2(n14691), .ZN(n10139) );
  OR2_X1 U12000 ( .A1(n13498), .A2(n14419), .ZN(n14525) );
  INV_X1 U12001 ( .A(n13475), .ZN(n10291) );
  NOR2_X1 U12002 ( .A1(n9875), .A2(n10211), .ZN(n10210) );
  XNOR2_X1 U12003 ( .A(n13497), .B(n11802), .ZN(n13483) );
  AND2_X1 U12004 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n11860), .ZN(
        n11804) );
  NOR2_X1 U12005 ( .A1(n11859), .A2(n20036), .ZN(n11860) );
  NAND2_X1 U12006 ( .A1(n12816), .A2(n12815), .ZN(n12951) );
  OR2_X1 U12007 ( .A1(n12810), .A2(n20241), .ZN(n12816) );
  NOR2_X1 U12008 ( .A1(n10016), .A2(n10017), .ZN(n10015) );
  NAND2_X1 U12009 ( .A1(n14644), .A2(n14627), .ZN(n10017) );
  INV_X1 U12010 ( .A(n14427), .ZN(n10016) );
  NAND2_X1 U12011 ( .A1(n14122), .A2(n10277), .ZN(n10276) );
  INV_X1 U12012 ( .A(n14132), .ZN(n10277) );
  NAND2_X1 U12013 ( .A1(n10275), .A2(n14107), .ZN(n10274) );
  INV_X1 U12014 ( .A(n10276), .ZN(n10275) );
  NAND2_X1 U12015 ( .A1(n10079), .A2(n10082), .ZN(n14481) );
  INV_X1 U12016 ( .A(n10083), .ZN(n10082) );
  NAND2_X1 U12017 ( .A1(n10280), .A2(n14189), .ZN(n10279) );
  INV_X1 U12018 ( .A(n14201), .ZN(n10280) );
  INV_X1 U12019 ( .A(n15970), .ZN(n10284) );
  OR2_X1 U12020 ( .A1(n11800), .A2(n11799), .ZN(n13485) );
  NAND2_X1 U12021 ( .A1(n14067), .A2(n14082), .ZN(n14059) );
  OR2_X1 U12022 ( .A1(n11674), .A2(n11673), .ZN(n12812) );
  INV_X1 U12023 ( .A(n12811), .ZN(n11706) );
  NAND2_X1 U12024 ( .A1(n10293), .A2(n10292), .ZN(n11694) );
  AOI21_X1 U12025 ( .B1(n10295), .B2(n11675), .A(n13495), .ZN(n10292) );
  NAND2_X1 U12026 ( .A1(n11838), .A2(n10295), .ZN(n10293) );
  AOI21_X1 U12027 ( .B1(n11676), .B2(n10297), .A(n10296), .ZN(n10295) );
  INV_X1 U12028 ( .A(n11740), .ZN(n13065) );
  INV_X1 U12029 ( .A(n11822), .ZN(n10289) );
  NAND2_X1 U12030 ( .A1(n11640), .A2(n9895), .ZN(n12366) );
  INV_X2 U12031 ( .A(n12820), .ZN(n11637) );
  INV_X1 U12032 ( .A(n11623), .ZN(n11645) );
  INV_X1 U12033 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20325) );
  NAND2_X1 U12034 ( .A1(n11764), .A2(n11763), .ZN(n13121) );
  NAND2_X1 U12035 ( .A1(n20500), .A2(n20902), .ZN(n11764) );
  NAND2_X1 U12036 ( .A1(n12355), .A2(n13494), .ZN(n12352) );
  NOR3_X1 U12037 ( .A1(n13872), .A2(n10086), .A3(n10087), .ZN(n13847) );
  OR2_X1 U12038 ( .A1(n10890), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10086) );
  AND2_X1 U12039 ( .A1(n12416), .A2(n13906), .ZN(n13850) );
  NAND2_X1 U12040 ( .A1(n10088), .A2(n13851), .ZN(n10087) );
  INV_X1 U12041 ( .A(n13855), .ZN(n10088) );
  AND2_X1 U12042 ( .A1(n19267), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n13855) );
  OR2_X1 U12043 ( .A1(n13872), .A2(n10890), .ZN(n13863) );
  AND2_X1 U12044 ( .A1(n13819), .A2(n10089), .ZN(n13835) );
  AND2_X1 U12045 ( .A1(n9853), .A2(n19056), .ZN(n10089) );
  AND2_X1 U12046 ( .A1(n13817), .A2(n13815), .ZN(n10090) );
  AND2_X1 U12047 ( .A1(n19247), .A2(n11461), .ZN(n9977) );
  INV_X1 U12048 ( .A(n10950), .ZN(n10951) );
  INV_X1 U12049 ( .A(n11257), .ZN(n10756) );
  NAND2_X1 U12050 ( .A1(n10268), .A2(n10267), .ZN(n10266) );
  INV_X1 U12051 ( .A(n14943), .ZN(n10268) );
  NOR2_X1 U12052 ( .A1(n14929), .A2(n10269), .ZN(n10267) );
  NAND2_X1 U12053 ( .A1(n10096), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11372) );
  NAND2_X1 U12054 ( .A1(n10096), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11365) );
  NAND2_X1 U12055 ( .A1(n11319), .A2(n11318), .ZN(n11320) );
  INV_X1 U12056 ( .A(n11362), .ZN(n10353) );
  INV_X1 U12057 ( .A(n11337), .ZN(n11360) );
  INV_X1 U12058 ( .A(n14889), .ZN(n10342) );
  NOR2_X1 U12059 ( .A1(n10344), .A2(n14879), .ZN(n10343) );
  INV_X1 U12060 ( .A(n14884), .ZN(n10344) );
  INV_X1 U12061 ( .A(n14900), .ZN(n10332) );
  NOR2_X1 U12062 ( .A1(n15070), .A2(n10164), .ZN(n10163) );
  NOR2_X1 U12063 ( .A1(n18982), .A2(n10142), .ZN(n10141) );
  INV_X1 U12064 ( .A(n14916), .ZN(n10192) );
  INV_X1 U12065 ( .A(n13418), .ZN(n11031) );
  NOR2_X1 U12066 ( .A1(n13298), .A2(n13299), .ZN(n13300) );
  NOR2_X1 U12067 ( .A1(n16295), .A2(n10168), .ZN(n10167) );
  INV_X1 U12068 ( .A(n10407), .ZN(n10166) );
  NOR3_X1 U12069 ( .A1(n14952), .A2(n14769), .A3(n10266), .ZN(n10799) );
  INV_X1 U12070 ( .A(n14766), .ZN(n10202) );
  AND2_X1 U12071 ( .A1(n12443), .A2(n14837), .ZN(n10203) );
  AND2_X1 U12072 ( .A1(n13981), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10328) );
  INV_X1 U12073 ( .A(n12429), .ZN(n10205) );
  INV_X1 U12074 ( .A(n10101), .ZN(n10100) );
  OR2_X1 U12075 ( .A1(n10324), .A2(n10040), .ZN(n10039) );
  NAND2_X1 U12076 ( .A1(n10325), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10324) );
  NAND2_X1 U12077 ( .A1(n10265), .A2(n15411), .ZN(n10264) );
  INV_X1 U12078 ( .A(n15422), .ZN(n10265) );
  NOR2_X1 U12079 ( .A1(n15195), .A2(n10255), .ZN(n10253) );
  NAND2_X1 U12080 ( .A1(n10253), .A2(n10257), .ZN(n10252) );
  NOR2_X1 U12081 ( .A1(n15488), .A2(n13826), .ZN(n10323) );
  NAND2_X1 U12082 ( .A1(n10200), .A2(n12918), .ZN(n10199) );
  INV_X1 U12083 ( .A(n12945), .ZN(n10200) );
  OR2_X1 U12084 ( .A1(n10600), .A2(n10599), .ZN(n10884) );
  NAND2_X1 U12085 ( .A1(n10238), .A2(n13402), .ZN(n10237) );
  NAND2_X1 U12086 ( .A1(n13392), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13391) );
  INV_X1 U12087 ( .A(n11078), .ZN(n11086) );
  OAI21_X1 U12088 ( .B1(n13241), .B2(n13927), .A(n13528), .ZN(n13242) );
  OR2_X1 U12089 ( .A1(n10521), .A2(n10520), .ZN(n13226) );
  NOR2_X1 U12090 ( .A1(n10528), .A2(n10527), .ZN(n10549) );
  NAND2_X1 U12091 ( .A1(n10901), .A2(n10900), .ZN(n10938) );
  NOR2_X1 U12092 ( .A1(n11114), .A2(n9972), .ZN(n9971) );
  NAND2_X1 U12093 ( .A1(n11113), .A2(n9973), .ZN(n9972) );
  NAND2_X1 U12094 ( .A1(n11113), .A2(n9973), .ZN(n9975) );
  AOI22_X1 U12095 ( .A1(n9835), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(n9840), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10813) );
  NAND2_X1 U12096 ( .A1(n9840), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10035) );
  AOI21_X1 U12097 ( .B1(n9836), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n10861), .ZN(n10817) );
  AOI22_X1 U12098 ( .A1(n11233), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9844), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10809) );
  AOI21_X1 U12099 ( .B1(n9836), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10829) );
  AND2_X1 U12100 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19691), .ZN(
        n11109) );
  INV_X1 U12101 ( .A(n10883), .ZN(n11429) );
  NOR2_X1 U12102 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18869), .ZN(
        n13764) );
  NAND2_X1 U12103 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18841), .ZN(
        n13648) );
  NOR2_X1 U12104 ( .A1(n13643), .A2(n13645), .ZN(n15604) );
  INV_X1 U12105 ( .A(n17724), .ZN(n16778) );
  INV_X1 U12106 ( .A(n17622), .ZN(n10186) );
  AOI21_X1 U12107 ( .B1(n18143), .B2(n10172), .A(n10171), .ZN(n15772) );
  INV_X1 U12108 ( .A(n15767), .ZN(n10172) );
  OAI21_X1 U12109 ( .B1(n15767), .B2(n17760), .A(n10173), .ZN(n10171) );
  NOR2_X1 U12110 ( .A1(n17816), .A2(n17817), .ZN(n15829) );
  OR2_X1 U12111 ( .A1(n17393), .A2(n15812), .ZN(n15810) );
  AOI21_X1 U12112 ( .B1(n10020), .B2(n10024), .A(n15759), .ZN(n15761) );
  NOR2_X1 U12113 ( .A1(n17854), .A2(n10022), .ZN(n10020) );
  XNOR2_X1 U12114 ( .A(n15819), .B(n17401), .ZN(n15757) );
  NOR2_X1 U12115 ( .A1(n18268), .A2(n17415), .ZN(n13756) );
  AND2_X1 U12116 ( .A1(n13205), .A2(n13189), .ZN(n19662) );
  AND2_X1 U12117 ( .A1(n11640), .A2(n11628), .ZN(n12579) );
  OR2_X1 U12118 ( .A1(n20021), .A2(n20020), .ZN(n20038) );
  OR3_X1 U12119 ( .A1(n20904), .A2(n13428), .A3(n13427), .ZN(n20059) );
  NOR2_X1 U12120 ( .A1(n14156), .A2(n14132), .ZN(n14133) );
  AND2_X1 U12121 ( .A1(n12798), .A2(n12797), .ZN(n12926) );
  AND2_X1 U12122 ( .A1(n14487), .A2(n12307), .ZN(n12198) );
  AND2_X1 U12123 ( .A1(n12127), .A2(n12126), .ZN(n14356) );
  OAI211_X1 U12124 ( .C1(n11978), .C2(n20122), .A(n11871), .B(n11870), .ZN(
        n13164) );
  AND2_X1 U12125 ( .A1(n12283), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13429) );
  AND2_X1 U12126 ( .A1(n10311), .A2(n10309), .ZN(n10308) );
  INV_X1 U12127 ( .A(n14087), .ZN(n10309) );
  AND2_X1 U12128 ( .A1(n12259), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12260) );
  NAND2_X1 U12129 ( .A1(n12260), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12282) );
  INV_X1 U12130 ( .A(n10312), .ZN(n10310) );
  AND2_X1 U12131 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n12178), .ZN(
        n12179) );
  INV_X1 U12132 ( .A(n12177), .ZN(n12178) );
  AND2_X1 U12133 ( .A1(n14357), .A2(n10315), .ZN(n14160) );
  NAND2_X1 U12134 ( .A1(n14357), .A2(n10317), .ZN(n14174) );
  NOR2_X1 U12135 ( .A1(n12124), .A2(n12123), .ZN(n12125) );
  NAND2_X1 U12136 ( .A1(n12125), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12177) );
  AND2_X1 U12137 ( .A1(n12105), .A2(n12104), .ZN(n14361) );
  NOR2_X1 U12138 ( .A1(n12086), .A2(n14513), .ZN(n12087) );
  NAND2_X1 U12139 ( .A1(n12054), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12086) );
  NOR2_X1 U12140 ( .A1(n10302), .A2(n14296), .ZN(n10301) );
  INV_X1 U12141 ( .A(n10304), .ZN(n10302) );
  NAND2_X1 U12142 ( .A1(n10303), .A2(n10304), .ZN(n14199) );
  NOR2_X1 U12143 ( .A1(n12019), .A2(n12018), .ZN(n12020) );
  NAND2_X1 U12144 ( .A1(n11986), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12019) );
  INV_X1 U12145 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12018) );
  AND2_X1 U12146 ( .A1(n16008), .A2(n14417), .ZN(n14541) );
  OR2_X1 U12147 ( .A1(n13498), .A2(n16118), .ZN(n16008) );
  NOR2_X1 U12148 ( .A1(n11962), .A2(n11961), .ZN(n11967) );
  AND2_X1 U12149 ( .A1(n11918), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11919) );
  NOR2_X1 U12150 ( .A1(n11914), .A2(n20006), .ZN(n11918) );
  NAND2_X1 U12151 ( .A1(n11888), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11914) );
  INV_X1 U12152 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20006) );
  CLKBUF_X1 U12153 ( .A(n13476), .Z(n13477) );
  CLKBUF_X1 U12154 ( .A(n13162), .Z(n13163) );
  NOR2_X1 U12155 ( .A1(n11813), .A2(n11803), .ZN(n11851) );
  XNOR2_X1 U12156 ( .A(n13060), .B(n20203), .ZN(n12962) );
  AOI21_X1 U12157 ( .B1(n11826), .B2(n10300), .A(n10299), .ZN(n10298) );
  INV_X1 U12158 ( .A(n11848), .ZN(n10299) );
  AND2_X1 U12159 ( .A1(n15879), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n14012) );
  NOR2_X1 U12160 ( .A1(n14156), .A2(n10276), .ZN(n14124) );
  NAND2_X1 U12161 ( .A1(n14452), .A2(n14427), .ZN(n14466) );
  NOR2_X1 U12162 ( .A1(n14427), .A2(n14653), .ZN(n14465) );
  INV_X1 U12163 ( .A(n10081), .ZN(n14426) );
  AOI21_X1 U12164 ( .B1(n14685), .B2(n16012), .A(n10084), .ZN(n10081) );
  NOR2_X1 U12165 ( .A1(n15926), .A2(n14049), .ZN(n14182) );
  OR2_X1 U12166 ( .A1(n9848), .A2(n15889), .ZN(n15926) );
  OAI21_X1 U12167 ( .B1(n10232), .B2(n14524), .A(n10230), .ZN(n14520) );
  INV_X1 U12168 ( .A(n10232), .ZN(n10226) );
  AOI21_X1 U12169 ( .B1(n14524), .B2(n10230), .A(n10229), .ZN(n10225) );
  NOR3_X1 U12170 ( .A1(n14311), .A2(n10281), .A3(n14201), .ZN(n14301) );
  NOR2_X1 U12171 ( .A1(n14311), .A2(n14201), .ZN(n14299) );
  XNOR2_X1 U12172 ( .A(n16024), .B(n16090), .ZN(n14694) );
  NAND2_X1 U12173 ( .A1(n14230), .A2(n14024), .ZN(n14309) );
  NOR2_X1 U12174 ( .A1(n14322), .A2(n14245), .ZN(n14244) );
  NAND2_X1 U12175 ( .A1(n16150), .A2(n10282), .ZN(n14322) );
  AND2_X1 U12176 ( .A1(n9913), .A2(n10283), .ZN(n10282) );
  INV_X1 U12177 ( .A(n14320), .ZN(n10283) );
  NAND2_X1 U12178 ( .A1(n16150), .A2(n9913), .ZN(n15973) );
  NAND2_X1 U12179 ( .A1(n16150), .A2(n13570), .ZN(n15971) );
  OR2_X1 U12180 ( .A1(n16012), .A2(n16156), .ZN(n10012) );
  AND2_X1 U12181 ( .A1(n10223), .A2(n10221), .ZN(n10011) );
  AND2_X1 U12182 ( .A1(n13443), .A2(n13442), .ZN(n13444) );
  NAND2_X1 U12183 ( .A1(n16173), .A2(n10285), .ZN(n16148) );
  AND2_X1 U12184 ( .A1(n9889), .A2(n10286), .ZN(n10285) );
  INV_X1 U12185 ( .A(n13444), .ZN(n10286) );
  OR2_X1 U12186 ( .A1(n16035), .A2(n16036), .ZN(n16033) );
  NAND2_X1 U12187 ( .A1(n16173), .A2(n9889), .ZN(n16161) );
  AND2_X1 U12188 ( .A1(n16173), .A2(n13183), .ZN(n16159) );
  AND2_X1 U12189 ( .A1(n13053), .A2(n13052), .ZN(n13054) );
  OR2_X1 U12190 ( .A1(n13118), .A2(n13054), .ZN(n16171) );
  AND4_X1 U12191 ( .A1(n11544), .A2(n11543), .A3(n11542), .A4(n11541), .ZN(
        n11555) );
  AND2_X1 U12192 ( .A1(n16117), .A2(n13506), .ZN(n14582) );
  NAND2_X1 U12193 ( .A1(n10294), .A2(n11676), .ZN(n11836) );
  INV_X1 U12194 ( .A(n12810), .ZN(n10216) );
  NAND2_X1 U12195 ( .A1(n11744), .A2(n11729), .ZN(n12848) );
  INV_X1 U12196 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12844) );
  AND3_X1 U12197 ( .A1(n12843), .A2(n12842), .A3(n12841), .ZN(n15853) );
  NAND2_X1 U12198 ( .A1(n13063), .A2(n20221), .ZN(n20368) );
  OR2_X1 U12199 ( .A1(n20471), .A2(n20692), .ZN(n20441) );
  AND2_X1 U12200 ( .A1(n20766), .A2(n20323), .ZN(n20556) );
  NAND2_X1 U12201 ( .A1(n20766), .A2(n20625), .ZN(n20588) );
  NAND3_X1 U12202 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20902), .A3(n20230), 
        .ZN(n20287) );
  NAND2_X1 U12203 ( .A1(n13909), .A2(n10893), .ZN(n13920) );
  OR2_X1 U12204 ( .A1(n12427), .A2(n10145), .ZN(n10146) );
  NAND2_X1 U12205 ( .A1(n15341), .A2(n9936), .ZN(n12465) );
  INV_X1 U12206 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10093) );
  INV_X1 U12207 ( .A(n13850), .ZN(n10892) );
  NAND2_X1 U12208 ( .A1(n13847), .A2(n10891), .ZN(n12416) );
  NOR2_X1 U12209 ( .A1(n10145), .A2(n18936), .ZN(n14780) );
  AND2_X1 U12210 ( .A1(n13860), .A2(n13862), .ZN(n18986) );
  NAND2_X1 U12211 ( .A1(n13819), .A2(n10090), .ZN(n13823) );
  AND2_X1 U12212 ( .A1(n11046), .A2(n11045), .ZN(n14895) );
  OR2_X1 U12213 ( .A1(n10669), .A2(n10668), .ZN(n13043) );
  AND2_X1 U12214 ( .A1(n11006), .A2(n11005), .ZN(n13035) );
  NAND2_X1 U12215 ( .A1(n11402), .A2(n11401), .ZN(n11405) );
  AOI21_X1 U12216 ( .B1(n11408), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n9949), .ZN(n11411) );
  NOR3_X1 U12217 ( .A1(n11418), .A2(n11417), .A3(n9948), .ZN(n11423) );
  NAND2_X1 U12218 ( .A1(n10348), .A2(n10346), .ZN(n14829) );
  AOI21_X1 U12219 ( .B1(n10351), .B2(n10350), .A(n10347), .ZN(n10346) );
  INV_X1 U12220 ( .A(n14835), .ZN(n10347) );
  AND2_X1 U12221 ( .A1(n10782), .A2(n10781), .ZN(n12420) );
  NAND2_X1 U12222 ( .A1(n14883), .A2(n14884), .ZN(n14878) );
  CLKBUF_X1 U12223 ( .A(n14887), .Z(n14888) );
  CLKBUF_X1 U12224 ( .A(n14892), .Z(n14893) );
  INV_X1 U12225 ( .A(n9827), .ZN(n10920) );
  CLKBUF_X1 U12226 ( .A(n10928), .Z(n10499) );
  OAI21_X1 U12227 ( .B1(n11480), .B2(n11479), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12570) );
  INV_X1 U12228 ( .A(n12570), .ZN(n13155) );
  NOR2_X1 U12229 ( .A1(n10384), .A2(n10380), .ZN(n10379) );
  OR2_X1 U12230 ( .A1(n10387), .A2(n15039), .ZN(n10384) );
  NAND2_X1 U12231 ( .A1(n10388), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10389) );
  NAND2_X1 U12232 ( .A1(n12418), .A2(n9931), .ZN(n12459) );
  AND2_X1 U12233 ( .A1(n10398), .A2(n10141), .ZN(n10419) );
  NAND2_X1 U12234 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10326) );
  AND2_X1 U12235 ( .A1(n13300), .A2(n9861), .ZN(n14909) );
  NAND2_X1 U12236 ( .A1(n10041), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10040) );
  NAND2_X1 U12237 ( .A1(n10398), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10420) );
  NAND2_X1 U12238 ( .A1(n13300), .A2(n11031), .ZN(n14917) );
  NOR2_X1 U12239 ( .A1(n9857), .A2(n10149), .ZN(n10148) );
  NOR2_X1 U12240 ( .A1(n13284), .A2(n13283), .ZN(n13286) );
  NOR2_X1 U12241 ( .A1(n10415), .A2(n19042), .ZN(n10414) );
  OR2_X1 U12242 ( .A1(n13145), .A2(n13130), .ZN(n13284) );
  NAND2_X1 U12243 ( .A1(n13143), .A2(n13142), .ZN(n13145) );
  NOR2_X1 U12244 ( .A1(n10407), .A2(n10165), .ZN(n10411) );
  NAND2_X1 U12245 ( .A1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n9849), .ZN(
        n10165) );
  NAND2_X1 U12246 ( .A1(n10166), .A2(n10167), .ZN(n10409) );
  NAND2_X1 U12247 ( .A1(n10408), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10407) );
  NAND2_X1 U12248 ( .A1(n10406), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10405) );
  NOR2_X1 U12249 ( .A1(n10405), .A2(n19235), .ZN(n10408) );
  AND2_X1 U12250 ( .A1(n10799), .A2(n10798), .ZN(n13960) );
  OR3_X1 U12251 ( .A1(n13925), .A2(n13941), .A3(n9832), .ZN(n14998) );
  AOI21_X1 U12252 ( .B1(n10008), .B2(n9869), .A(n10007), .ZN(n10005) );
  INV_X1 U12253 ( .A(n9892), .ZN(n10007) );
  NOR2_X1 U12254 ( .A1(n10008), .A2(n9846), .ZN(n10006) );
  AND2_X1 U12255 ( .A1(n10328), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10327) );
  OR2_X1 U12256 ( .A1(n13914), .A2(n13941), .ZN(n15023) );
  NAND2_X1 U12257 ( .A1(n13912), .A2(n13917), .ZN(n15047) );
  NAND2_X1 U12258 ( .A1(n12418), .A2(n9932), .ZN(n14860) );
  OR2_X1 U12259 ( .A1(n13903), .A2(n13902), .ZN(n13904) );
  NAND2_X1 U12260 ( .A1(n12418), .A2(n12419), .ZN(n12461) );
  NOR2_X1 U12261 ( .A1(n14897), .A2(n14886), .ZN(n14784) );
  NAND2_X1 U12262 ( .A1(n15341), .A2(n15340), .ZN(n15339) );
  NAND2_X1 U12263 ( .A1(n15341), .A2(n10271), .ZN(n14788) );
  NAND2_X1 U12264 ( .A1(n15149), .A2(n9989), .ZN(n9982) );
  OR2_X1 U12265 ( .A1(n9984), .A2(n15100), .ZN(n9981) );
  NOR2_X1 U12266 ( .A1(n10326), .A2(n15366), .ZN(n10325) );
  NOR2_X1 U12267 ( .A1(n9870), .A2(n15361), .ZN(n15360) );
  NAND2_X1 U12268 ( .A1(n9965), .A2(n15149), .ZN(n15139) );
  NAND2_X1 U12269 ( .A1(n10240), .A2(n9983), .ZN(n9965) );
  INV_X1 U12270 ( .A(n9986), .ZN(n9983) );
  AND2_X1 U12271 ( .A1(n10772), .A2(n10771), .ZN(n15393) );
  NOR3_X1 U12272 ( .A1(n15438), .A2(n10264), .A3(n15393), .ZN(n15394) );
  NOR2_X1 U12273 ( .A1(n15438), .A2(n15422), .ZN(n15421) );
  OAI21_X1 U12274 ( .B1(n15468), .B2(n10104), .A(n10101), .ZN(n15436) );
  NAND2_X1 U12275 ( .A1(n15451), .A2(n15439), .ZN(n15438) );
  AND2_X1 U12276 ( .A1(n15514), .A2(n10258), .ZN(n15470) );
  AND2_X1 U12277 ( .A1(n9914), .A2(n10259), .ZN(n10258) );
  INV_X1 U12278 ( .A(n15483), .ZN(n10259) );
  OR2_X1 U12279 ( .A1(n13831), .A2(n13830), .ZN(n15193) );
  NAND2_X1 U12280 ( .A1(n10256), .A2(n10254), .ZN(n15192) );
  NOR2_X1 U12281 ( .A1(n12944), .A2(n10193), .ZN(n13143) );
  NAND2_X1 U12282 ( .A1(n10194), .A2(n13044), .ZN(n10193) );
  INV_X1 U12283 ( .A(n10195), .ZN(n10194) );
  OR2_X1 U12284 ( .A1(n15208), .A2(n10257), .ZN(n10256) );
  AND3_X1 U12285 ( .A1(n10657), .A2(n10656), .A3(n10655), .ZN(n16298) );
  AND2_X1 U12286 ( .A1(n15514), .A2(n10260), .ZN(n16296) );
  NAND2_X1 U12287 ( .A1(n15514), .A2(n15513), .ZN(n16297) );
  OR2_X1 U12288 ( .A1(n12944), .A2(n10199), .ZN(n13036) );
  AND2_X1 U12289 ( .A1(n19082), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16275) );
  NAND2_X1 U12290 ( .A1(n9996), .A2(n13612), .ZN(n13812) );
  OAI22_X1 U12291 ( .A1(n11096), .A2(n11095), .B1(n10984), .B2(n10983), .ZN(
        n12896) );
  NOR2_X1 U12292 ( .A1(n12896), .A2(n12895), .ZN(n12912) );
  NAND2_X1 U12293 ( .A1(n13237), .A2(n9828), .ZN(n13241) );
  NAND2_X1 U12294 ( .A1(n10034), .A2(n11106), .ZN(n11108) );
  INV_X1 U12295 ( .A(n11122), .ZN(n13187) );
  OAI21_X1 U12296 ( .B1(n13958), .B2(n18926), .A(n10506), .ZN(n12634) );
  AND2_X1 U12297 ( .A1(n12633), .A2(n12634), .ZN(n12632) );
  AND4_X1 U12298 ( .A1(n12652), .A2(n12673), .A3(n10930), .A4(n10855), .ZN(
        n10925) );
  AND2_X2 U12299 ( .A1(n13186), .A2(n13199), .ZN(n19242) );
  NAND2_X1 U12300 ( .A1(n10842), .A2(n10861), .ZN(n10854) );
  NAND2_X1 U12301 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19758), .ZN(n19266) );
  NOR2_X1 U12302 ( .A1(n19522), .A2(n19488), .ZN(n19690) );
  AND2_X1 U12303 ( .A1(n11109), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19760) );
  INV_X1 U12304 ( .A(n13156), .ZN(n19753) );
  NAND3_X1 U12305 ( .A1(n10934), .A2(n10912), .A3(n9818), .ZN(n16346) );
  AND2_X1 U12306 ( .A1(n11449), .A2(n14747), .ZN(n11450) );
  NOR2_X2 U12307 ( .A1(n10933), .A2(n10837), .ZN(n10914) );
  AND2_X1 U12308 ( .A1(n10911), .A2(n10905), .ZN(n10836) );
  INV_X1 U12309 ( .A(n16376), .ZN(n18678) );
  NOR2_X1 U12310 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16793), .ZN(n16775) );
  NAND2_X1 U12311 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n10027) );
  NOR2_X1 U12312 ( .A1(n15718), .A2(n10029), .ZN(n10028) );
  INV_X1 U12313 ( .A(n15717), .ZN(n10029) );
  NOR2_X1 U12314 ( .A1(n17496), .A2(n10049), .ZN(n10048) );
  NOR2_X1 U12315 ( .A1(n17414), .A2(n17413), .ZN(n17442) );
  NOR2_X1 U12316 ( .A1(n18732), .A2(n18673), .ZN(n17473) );
  INV_X1 U12317 ( .A(n10120), .ZN(n10119) );
  NOR2_X1 U12318 ( .A1(n16409), .A2(n16611), .ZN(n16408) );
  INV_X1 U12319 ( .A(n17531), .ZN(n10179) );
  NAND2_X1 U12320 ( .A1(n16588), .A2(n9858), .ZN(n17534) );
  NOR2_X1 U12321 ( .A1(n17570), .A2(n10126), .ZN(n10125) );
  NAND2_X1 U12322 ( .A1(n16588), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17569) );
  NAND2_X1 U12323 ( .A1(n17632), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17611) );
  INV_X1 U12324 ( .A(n17725), .ZN(n16779) );
  NOR2_X1 U12325 ( .A1(n17541), .A2(n16437), .ZN(n15896) );
  AOI21_X1 U12326 ( .B1(n18100), .B2(n16444), .A(n16443), .ZN(n16445) );
  NOR2_X1 U12327 ( .A1(n16442), .A2(n18677), .ZN(n16443) );
  INV_X1 U12328 ( .A(n10185), .ZN(n17665) );
  INV_X1 U12329 ( .A(n18036), .ZN(n17964) );
  NAND2_X1 U12330 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17699), .ZN(
        n18099) );
  NOR2_X1 U12331 ( .A1(n18143), .A2(n17798), .ZN(n17797) );
  NOR2_X1 U12332 ( .A1(n17811), .A2(n18146), .ZN(n17810) );
  OR2_X1 U12333 ( .A1(n17836), .A2(n10189), .ZN(n10018) );
  OR2_X1 U12334 ( .A1(n17824), .A2(n17837), .ZN(n10189) );
  NAND2_X1 U12335 ( .A1(n15763), .A2(n10188), .ZN(n10187) );
  INV_X1 U12336 ( .A(n17824), .ZN(n10188) );
  OR2_X1 U12337 ( .A1(n17836), .A2(n17837), .ZN(n10191) );
  XNOR2_X1 U12338 ( .A(n15819), .B(n18845), .ZN(n17883) );
  NOR2_X1 U12339 ( .A1(n15804), .A2(n13759), .ZN(n15800) );
  NAND2_X1 U12340 ( .A1(n15801), .A2(n18902), .ZN(n18709) );
  INV_X1 U12341 ( .A(n18709), .ZN(n18684) );
  NAND2_X1 U12342 ( .A1(n13762), .A2(n15800), .ZN(n18670) );
  INV_X1 U12343 ( .A(n15806), .ZN(n13762) );
  NOR2_X2 U12344 ( .A1(n13664), .A2(n13663), .ZN(n18889) );
  NOR2_X1 U12345 ( .A1(n13696), .A2(n13695), .ZN(n18248) );
  NOR2_X1 U12346 ( .A1(n13740), .A2(n13739), .ZN(n18258) );
  NOR2_X1 U12347 ( .A1(n18735), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n16574) );
  INV_X1 U12348 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18735) );
  INV_X1 U12349 ( .A(n18732), .ZN(n18882) );
  OR2_X1 U12350 ( .A1(n10615), .A2(n10614), .ZN(n13598) );
  INV_X1 U12351 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20036) );
  INV_X1 U12352 ( .A(n20080), .ZN(n20060) );
  AND2_X1 U12353 ( .A1(n13450), .A2(n13437), .ZN(n20077) );
  AND2_X1 U12354 ( .A1(n20059), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20080) );
  AND2_X1 U12355 ( .A1(n13450), .A2(n13448), .ZN(n20069) );
  XNOR2_X1 U12356 ( .A(n12932), .B(n12926), .ZN(n20072) );
  CLKBUF_X1 U12357 ( .A(n11838), .Z(n11839) );
  AND2_X1 U12358 ( .A1(n13450), .A2(n13449), .ZN(n20075) );
  AND2_X1 U12359 ( .A1(n15937), .A2(n14254), .ZN(n20087) );
  INV_X1 U12360 ( .A(n14316), .ZN(n20097) );
  INV_X1 U12361 ( .A(n14362), .ZN(n14383) );
  INV_X1 U12362 ( .A(n14391), .ZN(n14405) );
  NOR2_X1 U12363 ( .A1(n14405), .A2(n13081), .ZN(n14407) );
  INV_X1 U12364 ( .A(n14407), .ZN(n14393) );
  AND2_X1 U12365 ( .A1(n12698), .A2(n12697), .ZN(n20105) );
  AND2_X1 U12366 ( .A1(n12765), .A2(n15873), .ZN(n12697) );
  AND2_X1 U12367 ( .A1(n15872), .A2(n20835), .ZN(n12966) );
  INV_X1 U12368 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14533) );
  INV_X1 U12369 ( .A(n10290), .ZN(n13057) );
  NAND2_X1 U12370 ( .A1(n13074), .A2(n13075), .ZN(n13058) );
  INV_X1 U12371 ( .A(n20159), .ZN(n19988) );
  NAND2_X1 U12372 ( .A1(n10213), .A2(n10212), .ZN(n14429) );
  OR2_X1 U12373 ( .A1(n14435), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10213) );
  NAND2_X1 U12374 ( .A1(n10215), .A2(n9850), .ZN(n14448) );
  OAI21_X1 U12375 ( .B1(n14685), .B2(n14422), .A(n13498), .ZN(n15985) );
  NAND2_X1 U12376 ( .A1(n10223), .A2(n10221), .ZN(n14411) );
  OAI21_X1 U12377 ( .B1(n20155), .B2(n10208), .A(n10207), .ZN(n13480) );
  AOI21_X1 U12378 ( .B1(n16049), .B2(n10211), .A(n9875), .ZN(n10207) );
  NAND2_X1 U12379 ( .A1(n16050), .A2(n16049), .ZN(n16048) );
  NAND2_X1 U12380 ( .A1(n20155), .A2(n13334), .ZN(n16050) );
  INV_X1 U12381 ( .A(n14582), .ZN(n20206) );
  NAND2_X1 U12382 ( .A1(n12795), .A2(n14734), .ZN(n16117) );
  INV_X1 U12383 ( .A(n20171), .ZN(n20214) );
  AOI21_X1 U12384 ( .B1(n13111), .B2(n13110), .A(n13109), .ZN(n14728) );
  INV_X1 U12385 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20634) );
  INV_X1 U12386 ( .A(n14728), .ZN(n20219) );
  NOR2_X1 U12387 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n16181) );
  OAI21_X1 U12388 ( .B1(n20411), .B2(n20396), .A(n20729), .ZN(n20414) );
  INV_X1 U12389 ( .A(n20441), .ZN(n20464) );
  NOR2_X1 U12390 ( .A1(n20686), .A2(n20470), .ZN(n20492) );
  OAI211_X1 U12391 ( .C1(n20523), .C2(n20641), .A(n20563), .B(n20508), .ZN(
        n20526) );
  INV_X1 U12392 ( .A(n20567), .ZN(n20584) );
  OAI21_X1 U12393 ( .B1(n20604), .B2(n20603), .A(n20602), .ZN(n20622) );
  OAI211_X1 U12394 ( .C1(n20646), .C2(n20641), .A(n20729), .B(n20640), .ZN(
        n20681) );
  OAI211_X1 U12395 ( .C1(n20753), .C2(n20730), .A(n20729), .B(n20728), .ZN(
        n20757) );
  NOR2_X1 U12396 ( .A1(n20686), .A2(n20763), .ZN(n20815) );
  INV_X1 U12397 ( .A(n20807), .ZN(n20820) );
  AND2_X1 U12398 ( .A1(n16192), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15879) );
  INV_X1 U12399 ( .A(n15879), .ZN(n20826) );
  INV_X2 U12400 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20898) );
  NOR2_X1 U12401 ( .A1(n10901), .A2(n12471), .ZN(n18911) );
  AOI21_X1 U12402 ( .B1(n10423), .B2(n15006), .A(n19831), .ZN(n10424) );
  NAND2_X1 U12403 ( .A1(n10160), .A2(n10158), .ZN(n14775) );
  NAND2_X1 U12404 ( .A1(n10159), .A2(n10162), .ZN(n10158) );
  INV_X1 U12405 ( .A(n10161), .ZN(n10159) );
  NAND2_X1 U12406 ( .A1(n12439), .A2(n15031), .ZN(n10157) );
  NOR2_X1 U12407 ( .A1(n15041), .A2(n12440), .ZN(n12439) );
  NAND2_X1 U12408 ( .A1(n10143), .A2(n10144), .ZN(n16214) );
  AND2_X1 U12409 ( .A1(n10146), .A2(n15062), .ZN(n16225) );
  INV_X1 U12410 ( .A(n10146), .ZN(n16227) );
  INV_X1 U12411 ( .A(n10155), .ZN(n12428) );
  NAND2_X1 U12412 ( .A1(n10892), .A2(n10094), .ZN(n12458) );
  NOR2_X1 U12413 ( .A1(n12412), .A2(n10145), .ZN(n12453) );
  NOR2_X1 U12414 ( .A1(n10145), .A2(n14779), .ZN(n12413) );
  NOR2_X1 U12415 ( .A1(n12413), .A2(n12414), .ZN(n12412) );
  AND2_X1 U12416 ( .A1(n18911), .A2(n16367), .ZN(n19036) );
  NAND2_X1 U12417 ( .A1(n19122), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19105) );
  INV_X1 U12418 ( .A(n19085), .ZN(n19109) );
  INV_X1 U12419 ( .A(n19036), .ZN(n19116) );
  NAND2_X1 U12420 ( .A1(n11137), .A2(n11136), .ZN(n14914) );
  OR2_X1 U12421 ( .A1(n10731), .A2(n10730), .ZN(n13294) );
  OR2_X1 U12422 ( .A1(n10700), .A2(n10699), .ZN(n13281) );
  AND2_X1 U12423 ( .A1(n9860), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10334) );
  INV_X1 U12424 ( .A(n11131), .ZN(n10336) );
  CLKBUF_X1 U12425 ( .A(n13038), .Z(n13039) );
  NAND2_X1 U12426 ( .A1(n12751), .A2(n12750), .ZN(n19522) );
  OR2_X1 U12427 ( .A1(n12748), .A2(n12749), .ZN(n12751) );
  INV_X1 U12428 ( .A(n14901), .ZN(n14921) );
  AND2_X1 U12429 ( .A1(n9879), .A2(n14930), .ZN(n16204) );
  CLKBUF_X1 U12430 ( .A(n14855), .Z(n14856) );
  CLKBUF_X1 U12431 ( .A(n14871), .Z(n14872) );
  AND2_X1 U12432 ( .A1(n12630), .A2(n13155), .ZN(n19129) );
  NOR2_X1 U12433 ( .A1(n19137), .A2(n19177), .ZN(n19169) );
  NAND2_X1 U12434 ( .A1(n12631), .A2(n14988), .ZN(n19162) );
  AND2_X1 U12435 ( .A1(n19160), .A2(n9978), .ZN(n19177) );
  AND2_X1 U12436 ( .A1(n19160), .A2(n10499), .ZN(n19137) );
  INV_X1 U12437 ( .A(n19162), .ZN(n19185) );
  NOR2_X1 U12438 ( .A1(n19186), .A2(n19218), .ZN(n19204) );
  BUF_X1 U12440 ( .A(n12719), .Z(n19218) );
  INV_X1 U12441 ( .A(n12614), .ZN(n12567) );
  OR2_X1 U12442 ( .A1(n12500), .A2(n14748), .ZN(n12614) );
  INV_X1 U12443 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n19042) );
  INV_X1 U12444 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n16295) );
  INV_X1 U12445 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19235) );
  NAND2_X1 U12446 ( .A1(n12596), .A2(n12595), .ZN(n19234) );
  CLKBUF_X1 U12447 ( .A(n13192), .Z(n13532) );
  INV_X1 U12448 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10404) );
  INV_X1 U12449 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14806) );
  AND2_X1 U12450 ( .A1(n19234), .A2(n12608), .ZN(n19222) );
  NAND2_X1 U12451 ( .A1(n12590), .A2(n19247), .ZN(n19225) );
  INV_X1 U12452 ( .A(n19234), .ZN(n15162) );
  XOR2_X1 U12453 ( .A(n13953), .B(n13952), .Z(n14825) );
  AND2_X1 U12454 ( .A1(n14849), .A2(n9942), .ZN(n13952) );
  AND2_X1 U12455 ( .A1(n15254), .A2(n15232), .ZN(n15253) );
  OR2_X1 U12456 ( .A1(n15313), .A2(n13980), .ZN(n15297) );
  NAND2_X1 U12457 ( .A1(n10001), .A2(n10097), .ZN(n15091) );
  NAND2_X1 U12458 ( .A1(n10240), .A2(n10241), .ZN(n15151) );
  NAND2_X1 U12459 ( .A1(n10244), .A2(n9847), .ZN(n15159) );
  NOR2_X1 U12460 ( .A1(n15169), .A2(n15174), .ZN(n15407) );
  NAND2_X1 U12461 ( .A1(n10105), .A2(n15465), .ZN(n15185) );
  OR2_X1 U12462 ( .A1(n15468), .A2(n15466), .ZN(n10105) );
  NAND2_X1 U12463 ( .A1(n15514), .A2(n9914), .ZN(n15484) );
  NOR2_X1 U12464 ( .A1(n13974), .A2(n13973), .ZN(n16307) );
  NOR2_X1 U12465 ( .A1(n12902), .A2(n10236), .ZN(n13403) );
  NAND2_X1 U12466 ( .A1(n9945), .A2(n10238), .ZN(n10236) );
  NAND2_X1 U12467 ( .A1(n9991), .A2(n13307), .ZN(n13384) );
  NAND2_X1 U12468 ( .A1(n13241), .A2(n9994), .ZN(n13276) );
  INV_X1 U12469 ( .A(n13269), .ZN(n9994) );
  OR2_X1 U12470 ( .A1(n12681), .A2(n16353), .ZN(n15374) );
  INV_X1 U12471 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13784) );
  INV_X1 U12472 ( .A(n16314), .ZN(n16304) );
  OR2_X1 U12473 ( .A1(n12681), .A2(n12663), .ZN(n16313) );
  INV_X1 U12474 ( .A(n15495), .ZN(n16322) );
  INV_X1 U12475 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19964) );
  NAND2_X1 U12476 ( .A1(n15527), .A2(n12584), .ZN(n19958) );
  INV_X1 U12477 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19955) );
  INV_X1 U12478 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19946) );
  INV_X1 U12479 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16340) );
  INV_X1 U12480 ( .A(n11127), .ZN(n15527) );
  AND2_X1 U12481 ( .A1(n12626), .A2(n12625), .ZN(n19949) );
  INV_X1 U12482 ( .A(n11433), .ZN(n15661) );
  INV_X1 U12483 ( .A(n19374), .ZN(n19365) );
  INV_X1 U12484 ( .A(n19384), .ZN(n19402) );
  AND2_X1 U12485 ( .A1(n19376), .A2(n19669), .ZN(n19429) );
  INV_X1 U12486 ( .A(n19447), .ZN(n19465) );
  AOI22_X1 U12487 ( .A1(n19496), .A2(n19495), .B1(n19494), .B2(n19825), .ZN(
        n19517) );
  INV_X1 U12488 ( .A(n19548), .ZN(n19551) );
  INV_X1 U12489 ( .A(n19574), .ZN(n19588) );
  INV_X1 U12490 ( .A(n19771), .ZN(n19637) );
  INV_X1 U12491 ( .A(n19778), .ZN(n19641) );
  INV_X1 U12492 ( .A(n19628), .ZN(n19657) );
  AND2_X1 U12493 ( .A1(n10915), .A2(n19275), .ZN(n19692) );
  INV_X1 U12494 ( .A(n19792), .ZN(n19720) );
  OAI22_X1 U12495 ( .A1(n20273), .A2(n19265), .B1(n19264), .B2(n19263), .ZN(
        n19726) );
  OAI21_X1 U12496 ( .B1(n19703), .B2(n19702), .A(n19701), .ZN(n19740) );
  AND2_X1 U12497 ( .A1(n19758), .A2(n19277), .ZN(n19741) );
  INV_X1 U12498 ( .A(n19735), .ZN(n19739) );
  INV_X1 U12499 ( .A(n19820), .ZN(n19738) );
  INV_X1 U12500 ( .A(n19706), .ZN(n19761) );
  INV_X1 U12501 ( .A(n19819), .ZN(n19797) );
  INV_X1 U12502 ( .A(n19730), .ZN(n19796) );
  NAND2_X1 U12503 ( .A1(n19690), .A2(n19753), .ZN(n19819) );
  AND2_X1 U12504 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19829), .ZN(n16362) );
  INV_X1 U12505 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n19832) );
  INV_X1 U12506 ( .A(n18886), .ZN(n18901) );
  INV_X1 U12507 ( .A(n17473), .ZN(n17414) );
  XNOR2_X1 U12508 ( .A(n16601), .B(n10116), .ZN(n10115) );
  INV_X1 U12509 ( .A(n16602), .ZN(n10116) );
  INV_X1 U12510 ( .A(n16606), .ZN(n10112) );
  NOR2_X1 U12511 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16747), .ZN(n16730) );
  INV_X1 U12512 ( .A(n16939), .ZN(n16915) );
  NOR2_X1 U12513 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16818), .ZN(n16799) );
  NOR2_X2 U12514 ( .A1(n18863), .A2(n16947), .ZN(n16873) );
  NOR2_X2 U12515 ( .A1(n18724), .A2(n16580), .ZN(n16939) );
  INV_X1 U12516 ( .A(n16952), .ZN(n16940) );
  NAND4_X1 U12517 ( .A1(n18201), .A2(n18901), .A3(n16902), .A4(n18730), .ZN(
        n16955) );
  INV_X1 U12518 ( .A(n17257), .ZN(n17260) );
  NOR2_X2 U12519 ( .A1(n17260), .A2(n18268), .ZN(n17261) );
  NAND2_X1 U12520 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(P3_EAX_REG_29__SCAN_IN), 
        .ZN(n10044) );
  NOR3_X1 U12521 ( .A1(n17290), .A2(n17489), .A3(n10045), .ZN(n17276) );
  NOR2_X1 U12522 ( .A1(n17290), .A2(n17489), .ZN(n17284) );
  NAND2_X1 U12523 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17294), .ZN(n17290) );
  NOR2_X1 U12524 ( .A1(n17424), .A2(n17301), .ZN(n17294) );
  OR2_X1 U12525 ( .A1(n17485), .A2(n17300), .ZN(n17301) );
  NOR2_X1 U12526 ( .A1(n17483), .A2(n9890), .ZN(n17305) );
  NOR2_X1 U12527 ( .A1(n17434), .A2(n17330), .ZN(n17325) );
  INV_X1 U12528 ( .A(n17335), .ZN(n17331) );
  NOR3_X1 U12529 ( .A1(n17351), .A2(n17346), .A3(n17441), .ZN(n17336) );
  NOR2_X1 U12530 ( .A1(n17400), .A2(n18263), .ZN(n17340) );
  NAND2_X1 U12531 ( .A1(n17355), .A2(P3_EAX_REG_15__SCAN_IN), .ZN(n17346) );
  NOR2_X1 U12532 ( .A1(n17350), .A2(n17445), .ZN(n17355) );
  INV_X1 U12533 ( .A(n18268), .ZN(n17351) );
  NAND2_X1 U12534 ( .A1(n17264), .A2(n10046), .ZN(n17377) );
  NOR2_X1 U12535 ( .A1(n10050), .A2(n10047), .ZN(n10046) );
  NAND2_X1 U12536 ( .A1(n10048), .A2(P3_EAX_REG_7__SCAN_IN), .ZN(n10047) );
  INV_X1 U12537 ( .A(n17381), .ZN(n10050) );
  NOR2_X1 U12538 ( .A1(n17377), .A2(n17504), .ZN(n17376) );
  NOR2_X1 U12539 ( .A1(n15686), .A2(n15685), .ZN(n17390) );
  NOR2_X1 U12540 ( .A1(n17468), .A2(n17442), .ZN(n17438) );
  CLKBUF_X1 U12541 ( .A(n17438), .Z(n17467) );
  CLKBUF_X1 U12542 ( .A(n17520), .Z(n17515) );
  INV_X1 U12543 ( .A(n17523), .ZN(n17516) );
  INV_X1 U12544 ( .A(n17803), .ZN(n17745) );
  NOR2_X1 U12545 ( .A1(n17827), .A2(n17859), .ZN(n10130) );
  NAND2_X1 U12546 ( .A1(n10131), .A2(n10132), .ZN(n17826) );
  NOR2_X1 U12547 ( .A1(n10133), .A2(n17859), .ZN(n10131) );
  NOR2_X1 U12548 ( .A1(n17845), .A2(n17859), .ZN(n17838) );
  INV_X1 U12549 ( .A(n18575), .ZN(n18616) );
  INV_X1 U12550 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17890) );
  NOR2_X1 U12551 ( .A1(n17844), .A2(n17846), .ZN(n17889) );
  INV_X1 U12552 ( .A(n17855), .ZN(n17891) );
  INV_X1 U12553 ( .A(n9816), .ZN(n17898) );
  INV_X1 U12554 ( .A(n16454), .ZN(n16455) );
  AOI21_X1 U12555 ( .B1(n17981), .B2(n17533), .A(n16453), .ZN(n16454) );
  AND2_X1 U12556 ( .A1(n17798), .A2(n17906), .ZN(n15779) );
  NAND2_X1 U12557 ( .A1(n17628), .A2(n15777), .ZN(n17580) );
  INV_X1 U12558 ( .A(n17628), .ZN(n17605) );
  INV_X2 U12559 ( .A(n18694), .ZN(n18104) );
  NAND2_X1 U12560 ( .A1(n10024), .A2(n10025), .ZN(n17853) );
  AND2_X1 U12561 ( .A1(n10021), .A2(n10024), .ZN(n17852) );
  NOR2_X1 U12562 ( .A1(n17854), .A2(n10022), .ZN(n10021) );
  NAND2_X1 U12563 ( .A1(n17864), .A2(n17865), .ZN(n17863) );
  AOI21_X2 U12564 ( .B1(n15797), .B2(n15796), .A(n18732), .ZN(n18214) );
  AOI211_X1 U12565 ( .C1(n15799), .C2(n15790), .A(n15789), .B(n15788), .ZN(
        n15797) );
  INV_X1 U12566 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18712) );
  INV_X1 U12567 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18716) );
  AND2_X1 U12568 ( .A1(n12391), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20227)
         );
  CLKBUF_X1 U12569 ( .A(n16538), .Z(n16544) );
  NAND2_X1 U12570 ( .A1(n14636), .A2(n20159), .ZN(n14467) );
  OAI21_X1 U12571 ( .B1(n14633), .B2(n20196), .A(n10140), .ZN(P1_U3003) );
  AOI21_X1 U12572 ( .B1(n14635), .B2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14634), .ZN(n10140) );
  OAI21_X1 U12573 ( .B1(n15223), .B2(n14919), .A(n12403), .ZN(n12404) );
  NAND2_X1 U12574 ( .A1(n14936), .A2(n14901), .ZN(n14846) );
  NAND2_X1 U12575 ( .A1(n10249), .A2(n16282), .ZN(n10248) );
  INV_X1 U12576 ( .A(n10249), .ZN(n15349) );
  NAND2_X1 U12577 ( .A1(n10114), .A2(n10111), .ZN(P3_U2641) );
  NOR4_X1 U12578 ( .A1(n9882), .A2(n16604), .A3(n10113), .A4(n10112), .ZN(
        n10111) );
  NAND2_X1 U12579 ( .A1(n10115), .A2(n18741), .ZN(n10114) );
  AND2_X1 U12580 ( .A1(n16614), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n10113) );
  NAND2_X1 U12581 ( .A1(n17264), .A2(P3_EAX_REG_0__SCAN_IN), .ZN(n17407) );
  AOI21_X1 U12582 ( .B1(n10178), .B2(n10176), .A(n10174), .ZN(n17538) );
  NAND2_X1 U12583 ( .A1(n13607), .A2(n13933), .ZN(n13608) );
  NOR2_X1 U12585 ( .A1(n18704), .A2(n13648), .ZN(n15581) );
  BUF_X1 U12586 ( .A(n15581), .Z(n17143) );
  AND2_X1 U12587 ( .A1(n13915), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9846) );
  NAND2_X1 U12588 ( .A1(n10398), .A2(n9856), .ZN(n10397) );
  OAI21_X2 U12589 ( .B1(n13992), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n13945), 
        .ZN(n13535) );
  NAND2_X1 U12590 ( .A1(n10388), .A2(n9867), .ZN(n10385) );
  AND2_X1 U12591 ( .A1(n15160), .A2(n15406), .ZN(n9847) );
  NAND2_X1 U12592 ( .A1(n15409), .A2(n10325), .ZN(n15125) );
  OR3_X1 U12593 ( .A1(n14311), .A2(n10279), .A3(n9919), .ZN(n9848) );
  NAND2_X1 U12594 ( .A1(n13186), .A2(n13193), .ZN(n13588) );
  NAND2_X1 U12595 ( .A1(n13560), .A2(n14238), .ZN(n14237) );
  NOR2_X1 U12596 ( .A1(n13648), .A2(n16944), .ZN(n13734) );
  NOR2_X1 U12597 ( .A1(n14887), .A2(n10338), .ZN(n11273) );
  NAND2_X1 U12598 ( .A1(n15497), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15198) );
  INV_X1 U12599 ( .A(n10930), .ZN(n9978) );
  AND2_X1 U12600 ( .A1(n10167), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9849) );
  AND4_X1 U12601 ( .A1(n10028), .A2(n15720), .A3(n15715), .A4(n9900), .ZN(
        n9851) );
  OR2_X1 U12602 ( .A1(n9875), .A2(n16049), .ZN(n9852) );
  XNOR2_X1 U12603 ( .A(n11342), .B(n10366), .ZN(n14850) );
  AND2_X1 U12604 ( .A1(n10090), .A2(n11008), .ZN(n9853) );
  NOR2_X1 U12605 ( .A1(n14865), .A2(n14866), .ZN(n9854) );
  OR2_X1 U12606 ( .A1(n13216), .A2(n10915), .ZN(n11433) );
  AND2_X1 U12607 ( .A1(n13910), .A2(n9947), .ZN(n9855) );
  NAND2_X1 U12608 ( .A1(n10335), .A2(n12890), .ZN(n12893) );
  INV_X4 U12609 ( .A(n13216), .ZN(n19247) );
  NAND2_X1 U12610 ( .A1(n10147), .A2(n10150), .ZN(n10402) );
  AND2_X1 U12611 ( .A1(n10141), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9856) );
  NAND2_X1 U12612 ( .A1(n10150), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9857) );
  AND2_X1 U12613 ( .A1(n10125), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9858) );
  AND2_X1 U12614 ( .A1(n11031), .A2(n10192), .ZN(n9859) );
  AND2_X1 U12615 ( .A1(n12890), .A2(n9935), .ZN(n9860) );
  AND2_X1 U12616 ( .A1(n9859), .A2(n14907), .ZN(n9861) );
  AND2_X1 U12617 ( .A1(n9916), .A2(n13466), .ZN(n9862) );
  AND2_X1 U12618 ( .A1(n10271), .A2(n10270), .ZN(n9863) );
  AND2_X1 U12619 ( .A1(n10144), .A2(n15050), .ZN(n9864) );
  AND2_X1 U12620 ( .A1(n9856), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9865) );
  INV_X1 U12621 ( .A(n12902), .ZN(n10234) );
  AND2_X1 U12622 ( .A1(n10234), .A2(n9945), .ZN(n9866) );
  AND2_X1 U12623 ( .A1(n10163), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9867) );
  AND2_X1 U12624 ( .A1(n10094), .A2(n10093), .ZN(n9868) );
  OR2_X1 U12625 ( .A1(n10569), .A2(n10568), .ZN(n13166) );
  NAND2_X1 U12626 ( .A1(n10010), .A2(n15255), .ZN(n9869) );
  AND2_X2 U12627 ( .A1(n11419), .A2(n10861), .ZN(n10603) );
  OR3_X1 U12628 ( .A1(n15438), .A2(n10262), .A3(n10264), .ZN(n9870) );
  CLKBUF_X3 U12629 ( .A(n15700), .Z(n17214) );
  OR3_X1 U12630 ( .A1(n17290), .A2(n17489), .A3(n10044), .ZN(n9872) );
  INV_X1 U12631 ( .A(n10026), .ZN(n15836) );
  OR2_X1 U12632 ( .A1(n17810), .A2(n15766), .ZN(n10026) );
  OR2_X1 U12633 ( .A1(n13643), .A2(n16944), .ZN(n9873) );
  OR2_X1 U12634 ( .A1(n12465), .A2(n12431), .ZN(n9874) );
  NOR2_X1 U12635 ( .A1(n15165), .A2(n15403), .ZN(n15152) );
  NAND2_X1 U12636 ( .A1(n9822), .A2(n13907), .ZN(n15046) );
  AND2_X1 U12637 ( .A1(n13342), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9875) );
  OR3_X1 U12638 ( .A1(n13872), .A2(n10087), .A3(n10890), .ZN(n9876) );
  NAND2_X1 U12639 ( .A1(n14357), .A2(n14356), .ZN(n14173) );
  NOR2_X1 U12640 ( .A1(n15175), .A2(n15425), .ZN(n15176) );
  NOR2_X1 U12641 ( .A1(n15165), .A2(n10326), .ZN(n15144) );
  NOR2_X1 U12642 ( .A1(n14213), .A2(n14307), .ZN(n14198) );
  OR2_X1 U12643 ( .A1(n15175), .A2(n10039), .ZN(n9877) );
  OR2_X1 U12644 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n16221), .ZN(n9878) );
  OR2_X1 U12645 ( .A1(n14952), .A2(n10266), .ZN(n9879) );
  AND2_X1 U12646 ( .A1(n14420), .A2(n16012), .ZN(n10232) );
  OR3_X1 U12647 ( .A1(n13872), .A2(n13855), .A3(n10890), .ZN(n9880) );
  NOR2_X1 U12648 ( .A1(n11132), .A2(n10336), .ZN(n9881) );
  NOR2_X1 U12649 ( .A1(n16617), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n9882) );
  INV_X1 U12650 ( .A(n10106), .ZN(n10104) );
  AOI21_X1 U12651 ( .B1(n15466), .B2(n15465), .A(n10107), .ZN(n10106) );
  AND4_X1 U12652 ( .A1(n11571), .A2(n11570), .A3(n11569), .A4(n11568), .ZN(
        n9884) );
  AND2_X1 U12653 ( .A1(n10817), .A2(n10035), .ZN(n9885) );
  AND2_X1 U12654 ( .A1(n15497), .A2(n10323), .ZN(n15199) );
  AND2_X1 U12655 ( .A1(n15341), .A2(n9863), .ZN(n9886) );
  NAND2_X1 U12656 ( .A1(n13378), .A2(n13377), .ZN(n9997) );
  OR2_X1 U12657 ( .A1(n14156), .A2(n10274), .ZN(n9888) );
  AND2_X1 U12658 ( .A1(n13183), .A2(n16158), .ZN(n9889) );
  OR3_X1 U12659 ( .A1(n17346), .A2(n17266), .A3(n10043), .ZN(n9890) );
  INV_X1 U12660 ( .A(n17799), .ZN(n17773) );
  NOR2_X1 U12661 ( .A1(n17898), .A2(n16392), .ZN(n17799) );
  OAI21_X1 U12662 ( .B1(n10226), .B2(n10228), .A(n10225), .ZN(n14509) );
  XNOR2_X1 U12663 ( .A(n10065), .B(n10064), .ZN(n11743) );
  INV_X1 U12664 ( .A(n11743), .ZN(n11821) );
  INV_X1 U12665 ( .A(n14519), .ZN(n10229) );
  AND2_X1 U12666 ( .A1(n12892), .A2(n11105), .ZN(n12749) );
  OR2_X1 U12667 ( .A1(n15525), .A2(n13191), .ZN(n13203) );
  INV_X1 U12668 ( .A(n13203), .ZN(n13199) );
  AND2_X1 U12669 ( .A1(n10157), .A2(n10161), .ZN(n9891) );
  NOR2_X2 U12670 ( .A1(n13709), .A2(n13708), .ZN(n18244) );
  INV_X1 U12671 ( .A(n9967), .ZN(n14851) );
  AND2_X1 U12672 ( .A1(n13917), .A2(n15056), .ZN(n9892) );
  AND2_X1 U12673 ( .A1(n10015), .A2(n10214), .ZN(n9893) );
  AND2_X1 U12674 ( .A1(n13189), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n9894) );
  NAND2_X1 U12675 ( .A1(n15086), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10042) );
  AND2_X1 U12676 ( .A1(n11628), .A2(n20241), .ZN(n9895) );
  INV_X1 U12677 ( .A(n14213), .ZN(n10303) );
  NAND2_X1 U12678 ( .A1(n14526), .A2(n14525), .ZN(n9896) );
  AND2_X1 U12679 ( .A1(n10235), .A2(n10233), .ZN(n9897) );
  AND2_X1 U12680 ( .A1(n15782), .A2(n15781), .ZN(n17540) );
  INV_X1 U12681 ( .A(n17540), .ZN(n10181) );
  OR2_X1 U12682 ( .A1(n15175), .A2(n10040), .ZN(n15165) );
  INV_X1 U12683 ( .A(n10255), .ZN(n10254) );
  NAND2_X1 U12684 ( .A1(n15506), .A2(n13822), .ZN(n10255) );
  INV_X1 U12685 ( .A(n13166), .ZN(n10239) );
  AOI21_X1 U12686 ( .B1(n15023), .B2(n15255), .A(n15055), .ZN(n13915) );
  OR2_X1 U12687 ( .A1(n10100), .A2(n10106), .ZN(n9898) );
  AND2_X1 U12688 ( .A1(n15173), .A2(n15170), .ZN(n15169) );
  INV_X1 U12689 ( .A(n15169), .ZN(n10245) );
  NAND2_X1 U12690 ( .A1(n15076), .A2(n10328), .ZN(n15029) );
  OAI21_X1 U12691 ( .B1(n13897), .B2(n9898), .A(n13896), .ZN(n10098) );
  INV_X1 U12692 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17827) );
  AND2_X1 U12693 ( .A1(n10354), .A2(n10352), .ZN(n9899) );
  AND3_X1 U12694 ( .A1(n15714), .A2(n15719), .A3(n10027), .ZN(n9900) );
  AND2_X1 U12695 ( .A1(n10256), .A2(n13822), .ZN(n9901) );
  NOR2_X1 U12696 ( .A1(n15780), .A2(n15779), .ZN(n9903) );
  NAND2_X1 U12697 ( .A1(n14120), .A2(n10311), .ZN(n14085) );
  NOR2_X1 U12698 ( .A1(n16194), .A2(n16195), .ZN(n9904) );
  OR2_X1 U12699 ( .A1(n10319), .A2(n9953), .ZN(n9905) );
  NAND2_X1 U12700 ( .A1(n14857), .A2(n11320), .ZN(n11342) );
  NAND2_X1 U12701 ( .A1(n11342), .A2(n10366), .ZN(n9906) );
  AND2_X1 U12702 ( .A1(n11636), .A2(n20241), .ZN(n9907) );
  INV_X1 U12703 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10426) );
  OR2_X1 U12704 ( .A1(n13481), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9908) );
  NAND2_X1 U12705 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15764), .ZN(
        n9909) );
  INV_X1 U12706 ( .A(n10507), .ZN(n10774) );
  AND2_X1 U12707 ( .A1(n11114), .A2(n9975), .ZN(n9910) );
  INV_X1 U12708 ( .A(n11996), .ZN(n10300) );
  NAND2_X1 U12709 ( .A1(n12750), .A2(n9881), .ZN(n10335) );
  INV_X1 U12710 ( .A(n11113), .ZN(n9976) );
  NOR2_X1 U12711 ( .A1(n14887), .A2(n14889), .ZN(n14883) );
  NAND2_X1 U12712 ( .A1(n11137), .A2(n9862), .ZN(n13464) );
  NOR2_X1 U12713 ( .A1(n10415), .A2(n9857), .ZN(n10400) );
  NOR2_X1 U12714 ( .A1(n10407), .A2(n16295), .ZN(n10403) );
  NOR2_X1 U12715 ( .A1(n14164), .A2(n14157), .ZN(n14055) );
  AND2_X1 U12716 ( .A1(n10892), .A2(n9868), .ZN(n9911) );
  INV_X1 U12717 ( .A(n14730), .ZN(n10058) );
  NOR2_X1 U12718 ( .A1(n10401), .A2(n18995), .ZN(n10398) );
  OR2_X1 U12719 ( .A1(n10654), .A2(n10653), .ZN(n13040) );
  NAND2_X1 U12720 ( .A1(n11873), .A2(n11872), .ZN(n13289) );
  BUF_X1 U12721 ( .A(n13050), .Z(n14046) );
  AND2_X1 U12722 ( .A1(n13300), .A2(n9859), .ZN(n9912) );
  AND2_X1 U12723 ( .A1(n13570), .A2(n10284), .ZN(n9913) );
  AND2_X1 U12724 ( .A1(n10260), .A2(n14793), .ZN(n9914) );
  AND2_X1 U12725 ( .A1(n10078), .A2(n11849), .ZN(n9915) );
  NAND2_X1 U12726 ( .A1(n12928), .A2(n11848), .ZN(n13074) );
  NOR2_X1 U12727 ( .A1(n12902), .A2(n10550), .ZN(n13165) );
  NAND2_X1 U12728 ( .A1(n16033), .A2(n13493), .ZN(n13633) );
  AND2_X1 U12729 ( .A1(n10333), .A2(n11136), .ZN(n9916) );
  AND2_X1 U12730 ( .A1(n11137), .A2(n9916), .ZN(n13465) );
  INV_X1 U12731 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11811) );
  OR2_X1 U12732 ( .A1(n13767), .A2(n18889), .ZN(n9917) );
  INV_X1 U12733 ( .A(n15465), .ZN(n10103) );
  NOR2_X1 U12734 ( .A1(n14873), .A2(n11274), .ZN(n14865) );
  NAND2_X1 U12735 ( .A1(n10856), .A2(n10925), .ZN(n11452) );
  AND2_X1 U12736 ( .A1(n11858), .A2(n11849), .ZN(n9918) );
  INV_X1 U12737 ( .A(n10278), .ZN(n14291) );
  NOR3_X1 U12738 ( .A1(n14311), .A2(n10279), .A3(n10281), .ZN(n10278) );
  AND2_X1 U12739 ( .A1(n14784), .A2(n14783), .ZN(n12418) );
  NAND2_X1 U12740 ( .A1(n10166), .A2(n9849), .ZN(n10169) );
  OR2_X1 U12741 ( .A1(n14038), .A2(n10281), .ZN(n9919) );
  NAND2_X1 U12742 ( .A1(n13397), .A2(n13398), .ZN(n13604) );
  AND2_X1 U12743 ( .A1(n10334), .A2(n13040), .ZN(n9920) );
  AND2_X1 U12744 ( .A1(n9993), .A2(n10929), .ZN(n11451) );
  NOR2_X1 U12745 ( .A1(n17797), .A2(n15767), .ZN(n9921) );
  INV_X1 U12746 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n19017) );
  INV_X1 U12747 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n18909) );
  NAND2_X1 U12748 ( .A1(n13819), .A2(n9853), .ZN(n10091) );
  OR2_X1 U12749 ( .A1(n15438), .A2(n10264), .ZN(n9922) );
  AND3_X1 U12750 ( .A1(n13498), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n9923) );
  AND2_X1 U12751 ( .A1(n10315), .A2(n14150), .ZN(n9924) );
  AND2_X1 U12752 ( .A1(n11887), .A2(n10291), .ZN(n9925) );
  AND2_X1 U12753 ( .A1(n9858), .A2(n10124), .ZN(n9926) );
  AND2_X1 U12754 ( .A1(n9862), .A2(n10332), .ZN(n9927) );
  AOI21_X1 U12755 ( .B1(n12413), .B2(n13535), .A(n10156), .ZN(n10154) );
  AND2_X1 U12756 ( .A1(n9861), .A2(n14903), .ZN(n9928) );
  INV_X2 U12757 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20902) );
  AND2_X1 U12758 ( .A1(n11494), .A2(n11495), .ZN(n11954) );
  AND2_X1 U12759 ( .A1(n17264), .A2(n10048), .ZN(n9929) );
  INV_X1 U12760 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n10170) );
  AND2_X1 U12761 ( .A1(n16588), .A2(n10125), .ZN(n9930) );
  AND2_X1 U12762 ( .A1(n10335), .A2(n9860), .ZN(n12917) );
  INV_X1 U12763 ( .A(n11137), .ZN(n13295) );
  AND2_X1 U12764 ( .A1(n10391), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10388) );
  NOR2_X1 U12765 ( .A1(n10395), .A2(n15110), .ZN(n10391) );
  AND2_X1 U12766 ( .A1(n10398), .A2(n9865), .ZN(n10396) );
  AND2_X1 U12767 ( .A1(n10206), .A2(n12419), .ZN(n9931) );
  AND2_X1 U12768 ( .A1(n9931), .A2(n10205), .ZN(n9932) );
  NAND3_X2 U12769 ( .A1(n10426), .A2(n10320), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11238) );
  INV_X2 U12770 ( .A(n11238), .ZN(n11409) );
  AND2_X1 U12771 ( .A1(n10203), .A2(n10202), .ZN(n9933) );
  INV_X1 U12772 ( .A(n13927), .ZN(n13941) );
  INV_X1 U12773 ( .A(n16450), .ZN(n10173) );
  INV_X1 U12774 ( .A(n12415), .ZN(n10095) );
  AND2_X1 U12775 ( .A1(n10388), .A2(n10163), .ZN(n9934) );
  INV_X1 U12776 ( .A(n11296), .ZN(n10345) );
  NAND2_X1 U12777 ( .A1(n12750), .A2(n11131), .ZN(n12889) );
  AND2_X1 U12778 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n9935) );
  AND2_X1 U12779 ( .A1(n9863), .A2(n12463), .ZN(n9936) );
  AND2_X1 U12780 ( .A1(n10335), .A2(n10334), .ZN(n9937) );
  AND2_X1 U12781 ( .A1(n11296), .A2(n11295), .ZN(n9938) );
  NOR2_X1 U12782 ( .A1(n12944), .A2(n10195), .ZN(n9939) );
  AND2_X1 U12783 ( .A1(n10343), .A2(n10342), .ZN(n10341) );
  INV_X1 U12784 ( .A(n10341), .ZN(n10338) );
  AND2_X1 U12785 ( .A1(n10162), .A2(n15031), .ZN(n9940) );
  INV_X1 U12786 ( .A(n10198), .ZN(n12946) );
  OR2_X1 U12787 ( .A1(n12944), .A2(n12945), .ZN(n10198) );
  AND2_X1 U12788 ( .A1(n9932), .A2(n10204), .ZN(n9941) );
  AND2_X1 U12789 ( .A1(n9933), .A2(n10201), .ZN(n9942) );
  AND2_X1 U12790 ( .A1(n10191), .A2(n10190), .ZN(n9943) );
  AND2_X1 U12791 ( .A1(n9867), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9944) );
  AND2_X1 U12792 ( .A1(n10235), .A2(n13166), .ZN(n9945) );
  NOR2_X1 U12793 ( .A1(n13645), .A2(n13648), .ZN(n15676) );
  INV_X1 U12794 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10164) );
  NAND2_X1 U12795 ( .A1(n17864), .A2(n10019), .ZN(n10024) );
  INV_X1 U12796 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10126) );
  NAND2_X1 U12797 ( .A1(n12590), .A2(n14748), .ZN(n19227) );
  INV_X1 U12798 ( .A(n19227), .ZN(n16282) );
  NAND2_X1 U12799 ( .A1(n10912), .A2(n10925), .ZN(n15657) );
  AND2_X1 U12800 ( .A1(n10096), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n9946) );
  AND2_X1 U12801 ( .A1(n13927), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9947) );
  INV_X1 U12802 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10142) );
  INV_X1 U12803 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18982) );
  INV_X1 U12804 ( .A(n14844), .ZN(n10352) );
  NAND2_X1 U12805 ( .A1(n19247), .A2(n11364), .ZN(n14844) );
  INV_X1 U12806 ( .A(n17845), .ZN(n10132) );
  INV_X1 U12807 ( .A(n12597), .ZN(n9973) );
  AND2_X1 U12808 ( .A1(n10096), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n9948) );
  AND2_X1 U12809 ( .A1(n10096), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n9949) );
  INV_X1 U12810 ( .A(n15425), .ZN(n10041) );
  INV_X1 U12811 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10127) );
  AND2_X1 U12812 ( .A1(n10323), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9950) );
  INV_X1 U12813 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10122) );
  INV_X1 U12814 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10129) );
  INV_X1 U12815 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n10051) );
  INV_X1 U12816 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n10049) );
  INV_X1 U12817 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n10123) );
  INV_X1 U12818 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10149) );
  INV_X1 U12819 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10151) );
  INV_X1 U12820 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10168) );
  INV_X1 U12821 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10133) );
  INV_X1 U12822 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n10045) );
  INV_X1 U12823 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10010) );
  INV_X1 U12824 ( .A(n14326), .ZN(n20098) );
  INV_X1 U12825 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18863) );
  NOR2_X2 U12826 ( .A1(n18256), .A2(n18575), .ZN(n18594) );
  OR2_X1 U12827 ( .A1(n18426), .A2(n18473), .ZN(n18575) );
  NOR3_X2 U12828 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n9814), .A3(
        n18272), .ZN(n18288) );
  NOR3_X2 U12829 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n9814), .A3(
        n18356), .ZN(n18374) );
  NOR3_X2 U12830 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n9814), .A3(
        n18496), .ZN(n18467) );
  OAI22_X2 U12831 ( .A1(n14335), .A2(n20291), .B1(n21274), .B2(n20290), .ZN(
        n20743) );
  OAI22_X2 U12832 ( .A1(n20285), .A2(n20290), .B1(n20284), .B2(n20291), .ZN(
        n20755) );
  NOR4_X2 U12833 ( .A1(n17679), .A2(n17760), .A3(n18135), .A4(n18146), .ZN(
        n17774) );
  AND3_X1 U12834 ( .A1(n10018), .A2(n10187), .A3(n9909), .ZN(n17679) );
  NOR3_X2 U12835 ( .A1(n9814), .A2(n18522), .A3(n18496), .ZN(n18491) );
  NOR3_X4 U12836 ( .A1(n12500), .A2(n19247), .A3(n19851), .ZN(n12572) );
  OAI22_X2 U12837 ( .A1(n20255), .A2(n20291), .B1(n21104), .B2(n20290), .ZN(
        n20739) );
  OAI22_X2 U12838 ( .A1(n20277), .A2(n20291), .B1(n21251), .B2(n20290), .ZN(
        n20749) );
  NAND2_X1 U12839 ( .A1(n20158), .A2(n20228), .ZN(n20290) );
  NAND2_X1 U12840 ( .A1(n20158), .A2(n20227), .ZN(n20291) );
  NAND2_X1 U12841 ( .A1(n9952), .A2(n10950), .ZN(n9951) );
  NAND3_X1 U12842 ( .A1(n10926), .A2(n16347), .A3(n15657), .ZN(n12669) );
  NAND2_X1 U12843 ( .A1(n10948), .A2(n12679), .ZN(n9952) );
  NAND2_X1 U12844 ( .A1(n10932), .A2(n10931), .ZN(n10948) );
  AND2_X1 U12845 ( .A1(n9954), .A2(n9955), .ZN(n9953) );
  NOR2_X2 U12846 ( .A1(n10319), .A2(n13204), .ZN(n13356) );
  NOR2_X2 U12847 ( .A1(n10319), .A2(n13206), .ZN(n13579) );
  AND3_X2 U12848 ( .A1(n9902), .A2(n9959), .A3(n9956), .ZN(n13208) );
  NAND2_X1 U12849 ( .A1(n19593), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n9963) );
  INV_X1 U12850 ( .A(n11461), .ZN(n10928) );
  NAND3_X1 U12851 ( .A1(n9992), .A2(n9993), .A3(n11453), .ZN(n12672) );
  NAND2_X1 U12852 ( .A1(n12644), .A2(n11461), .ZN(n11453) );
  NAND2_X1 U12853 ( .A1(n10965), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10941) );
  AND2_X2 U12854 ( .A1(n9967), .A2(n9906), .ZN(n11363) );
  OAI211_X1 U12855 ( .C1(n13185), .C2(n9974), .A(n9968), .B(n9970), .ZN(n9969)
         );
  INV_X1 U12856 ( .A(n9969), .ZN(n12690) );
  AND2_X2 U12857 ( .A1(n10905), .A2(n10899), .ZN(n10912) );
  AND2_X2 U12858 ( .A1(n11137), .A2(n9927), .ZN(n14892) );
  AND2_X2 U12859 ( .A1(n13173), .A2(n11135), .ZN(n11137) );
  AND2_X2 U12860 ( .A1(n12661), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10952) );
  INV_X2 U12861 ( .A(n10952), .ZN(n11078) );
  NOR2_X2 U12862 ( .A1(n13542), .A2(n13192), .ZN(n13186) );
  INV_X1 U12863 ( .A(n15118), .ZN(n9988) );
  INV_X1 U12864 ( .A(n15100), .ZN(n9989) );
  NAND3_X1 U12865 ( .A1(n9991), .A2(n13386), .A3(n13307), .ZN(n13389) );
  INV_X1 U12866 ( .A(n13242), .ZN(n9990) );
  NAND2_X1 U12867 ( .A1(n12672), .A2(n10902), .ZN(n10932) );
  AOI21_X2 U12868 ( .B1(n15436), .B2(n15433), .A(n15097), .ZN(n15173) );
  NAND2_X1 U12869 ( .A1(n13812), .A2(n13811), .ZN(n9995) );
  NAND2_X1 U12870 ( .A1(n13610), .A2(n13609), .ZN(n9996) );
  NAND2_X1 U12871 ( .A1(n15468), .A2(n9998), .ZN(n9999) );
  NAND3_X1 U12872 ( .A1(n10000), .A2(n9999), .A3(n15088), .ZN(n15083) );
  INV_X1 U12873 ( .A(n14524), .ZN(n10138) );
  NAND2_X4 U12874 ( .A1(n13497), .A2(n13496), .ZN(n13498) );
  INV_X2 U12875 ( .A(n11850), .ZN(n10135) );
  NAND2_X1 U12876 ( .A1(n10018), .A2(n10187), .ZN(n17823) );
  NAND2_X1 U12877 ( .A1(n17865), .A2(n10170), .ZN(n10025) );
  XNOR2_X1 U12878 ( .A(n15743), .B(n15813), .ZN(n15744) );
  INV_X1 U12879 ( .A(n17552), .ZN(n10030) );
  AND2_X2 U12880 ( .A1(n17628), .A2(n10031), .ZN(n17579) );
  INV_X2 U12881 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18869) );
  NAND2_X1 U12882 ( .A1(n10975), .A2(n10034), .ZN(n11096) );
  OR2_X2 U12883 ( .A1(n13396), .A2(n13618), .ZN(n13606) );
  OR2_X2 U12884 ( .A1(n15175), .A2(n10037), .ZN(n15108) );
  INV_X2 U12885 ( .A(n10042), .ZN(n15076) );
  INV_X2 U12886 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18861) );
  NAND3_X1 U12887 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(P3_EAX_REG_16__SCAN_IN), 
        .A3(P3_EAX_REG_21__SCAN_IN), .ZN(n10043) );
  INV_X1 U12888 ( .A(n17276), .ZN(n17281) );
  NAND3_X1 U12889 ( .A1(n9852), .A2(n10209), .A3(n9908), .ZN(n10056) );
  OAI21_X1 U12890 ( .B1(n12757), .B2(n10059), .A(n10057), .ZN(n10063) );
  AOI21_X1 U12891 ( .B1(n11635), .B2(n10058), .A(n20902), .ZN(n10057) );
  INV_X1 U12892 ( .A(n11635), .ZN(n10059) );
  AND3_X2 U12893 ( .A1(n11626), .A2(n10370), .A3(n11627), .ZN(n11640) );
  NAND3_X1 U12894 ( .A1(n10063), .A2(n11699), .A3(n10060), .ZN(n11714) );
  NAND2_X1 U12895 ( .A1(n11640), .A2(n9907), .ZN(n10061) );
  NAND2_X1 U12896 ( .A1(n10062), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11699) );
  NAND3_X1 U12897 ( .A1(n12366), .A2(n12793), .A3(n11622), .ZN(n10062) );
  OAI22_X2 U12898 ( .A1(n12848), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n13065), 
        .B2(n11751), .ZN(n10065) );
  NAND2_X1 U12899 ( .A1(n10135), .A2(n10070), .ZN(n10069) );
  OAI211_X1 U12900 ( .C1(n10135), .C2(n10071), .A(n13341), .B(n10069), .ZN(
        n13342) );
  OAI211_X1 U12901 ( .C1(n10135), .C2(n10078), .A(n10076), .B(n10072), .ZN(
        n13335) );
  NAND2_X1 U12902 ( .A1(n10135), .A2(n9915), .ZN(n10072) );
  INV_X1 U12903 ( .A(n10076), .ZN(n10074) );
  NAND2_X1 U12904 ( .A1(n10136), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14685) );
  NAND2_X1 U12905 ( .A1(n10136), .A2(n10080), .ZN(n10079) );
  OAI21_X1 U12906 ( .B1(n10084), .B2(n16012), .A(n16012), .ZN(n10083) );
  AND2_X1 U12907 ( .A1(n13819), .A2(n13817), .ZN(n13816) );
  INV_X1 U12908 ( .A(n10091), .ZN(n13827) );
  NAND2_X1 U12909 ( .A1(n10892), .A2(n12415), .ZN(n12456) );
  CLKBUF_X1 U12910 ( .A(n9839), .Z(n10096) );
  INV_X1 U12911 ( .A(n10098), .ZN(n10097) );
  NAND3_X1 U12912 ( .A1(n9822), .A2(n13913), .A3(n13907), .ZN(n15021) );
  OR2_X2 U12913 ( .A1(n15067), .A2(n13908), .ZN(n10110) );
  NOR2_X1 U12914 ( .A1(n15055), .A2(n10109), .ZN(n10108) );
  INV_X1 U12915 ( .A(n13907), .ZN(n10109) );
  AOI211_X1 U12916 ( .C1(n16409), .C2(n10123), .A(n10117), .B(n10119), .ZN(
        n10118) );
  INV_X1 U12917 ( .A(n16911), .ZN(n16878) );
  INV_X1 U12918 ( .A(n17535), .ZN(n10124) );
  NOR2_X1 U12919 ( .A1(n17859), .A2(n10129), .ZN(n10128) );
  NAND3_X1 U12920 ( .A1(n10132), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A3(
        n10130), .ZN(n10134) );
  INV_X1 U12921 ( .A(n10134), .ZN(n17788) );
  INV_X2 U12922 ( .A(n16024), .ZN(n16012) );
  INV_X1 U12923 ( .A(n10415), .ZN(n10147) );
  NAND2_X1 U12924 ( .A1(n10147), .A2(n10148), .ZN(n10401) );
  OAI21_X1 U12925 ( .B1(n12413), .B2(n10156), .A(n10152), .ZN(n10155) );
  INV_X1 U12926 ( .A(n10153), .ZN(n10152) );
  OAI21_X1 U12927 ( .B1(n10156), .B2(n13535), .A(n13535), .ZN(n10153) );
  NAND2_X1 U12928 ( .A1(n12439), .A2(n9940), .ZN(n10160) );
  NOR2_X1 U12929 ( .A1(n12439), .A2(n10145), .ZN(n16194) );
  AOI21_X1 U12930 ( .B1(n10145), .B2(n15031), .A(n10145), .ZN(n10161) );
  INV_X1 U12931 ( .A(n15017), .ZN(n10162) );
  NAND2_X1 U12932 ( .A1(n10388), .A2(n9944), .ZN(n10387) );
  INV_X1 U12933 ( .A(n10169), .ZN(n10410) );
  XNOR2_X2 U12934 ( .A(n10026), .B(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18143) );
  INV_X1 U12935 ( .A(n10191), .ZN(n17835) );
  INV_X1 U12936 ( .A(n15763), .ZN(n10190) );
  NAND2_X1 U12937 ( .A1(n13300), .A2(n9928), .ZN(n14902) );
  NAND2_X1 U12938 ( .A1(n14849), .A2(n9933), .ZN(n14768) );
  NAND2_X1 U12939 ( .A1(n14849), .A2(n10203), .ZN(n14840) );
  AND2_X1 U12940 ( .A1(n14849), .A2(n12443), .ZN(n14838) );
  AND2_X2 U12941 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13096) );
  NOR2_X4 U12942 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11505) );
  INV_X1 U12943 ( .A(n12955), .ZN(n20221) );
  NAND2_X1 U12944 ( .A1(n12955), .A2(n13494), .ZN(n12960) );
  NAND2_X1 U12945 ( .A1(n12955), .A2(n13121), .ZN(n20769) );
  NAND2_X1 U12946 ( .A1(n12955), .A2(n13123), .ZN(n20471) );
  NOR2_X1 U12947 ( .A1(n13063), .A2(n12955), .ZN(n20590) );
  MUX2_X1 U12948 ( .A(n14725), .B(n20472), .S(n12955), .Z(n14726) );
  NAND2_X1 U12949 ( .A1(n20155), .A2(n10210), .ZN(n10209) );
  NAND3_X1 U12950 ( .A1(n10215), .A2(n9850), .A3(n9923), .ZN(n10212) );
  NOR2_X1 U12951 ( .A1(n16012), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10214) );
  NAND2_X1 U12952 ( .A1(n14465), .A2(n14428), .ZN(n14437) );
  NOR2_X1 U12953 ( .A1(n13632), .A2(n10220), .ZN(n10219) );
  OAI21_X1 U12954 ( .B1(n10224), .B2(n13632), .A(n13631), .ZN(n10222) );
  AND2_X1 U12955 ( .A1(n10244), .A2(n15406), .ZN(n15161) );
  NAND2_X1 U12956 ( .A1(n10248), .A2(n15124), .ZN(P2_U2994) );
  NAND2_X1 U12957 ( .A1(n15118), .A2(n15117), .ZN(n10250) );
  OR3_X1 U12958 ( .A1(n14952), .A2(n10269), .A3(n14943), .ZN(n12446) );
  NOR2_X1 U12959 ( .A1(n14952), .A2(n14943), .ZN(n14945) );
  INV_X1 U12960 ( .A(n12445), .ZN(n10269) );
  INV_X1 U12961 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10273) );
  INV_X1 U12962 ( .A(n14298), .ZN(n10281) );
  NAND2_X1 U12963 ( .A1(n12932), .A2(n10287), .ZN(n12939) );
  NAND2_X1 U12964 ( .A1(n11821), .A2(n10289), .ZN(n11809) );
  NAND3_X1 U12965 ( .A1(n10289), .A2(n11821), .A3(n13121), .ZN(n11850) );
  NAND3_X1 U12966 ( .A1(n13074), .A2(n13075), .A3(n10290), .ZN(n13056) );
  NOR2_X2 U12967 ( .A1(n13056), .A2(n13135), .ZN(n13134) );
  NAND3_X1 U12968 ( .A1(n11873), .A2(n11872), .A3(n11887), .ZN(n13413) );
  AND3_X2 U12969 ( .A1(n11873), .A2(n11872), .A3(n9925), .ZN(n13476) );
  NAND2_X1 U12970 ( .A1(n11838), .A2(n20902), .ZN(n10294) );
  OAI21_X1 U12971 ( .B1(n12955), .B2(n11825), .A(n10298), .ZN(n12931) );
  XNOR2_X2 U12972 ( .A(n11822), .B(n11821), .ZN(n12955) );
  NAND2_X1 U12973 ( .A1(n10303), .A2(n10301), .ZN(n14188) );
  NAND2_X1 U12974 ( .A1(n13560), .A2(n10306), .ZN(n14226) );
  INV_X1 U12975 ( .A(n14226), .ZN(n11985) );
  AND2_X1 U12976 ( .A1(n14120), .A2(n10310), .ZN(n14096) );
  NAND2_X1 U12977 ( .A1(n14120), .A2(n14121), .ZN(n14109) );
  NAND2_X1 U12978 ( .A1(n14357), .A2(n9924), .ZN(n14135) );
  NOR2_X2 U12979 ( .A1(n10319), .A2(n13203), .ZN(n19380) );
  NOR2_X2 U12980 ( .A1(n10319), .A2(n13202), .ZN(n19443) );
  OR2_X2 U12981 ( .A1(n13188), .A2(n13192), .ZN(n10319) );
  NAND2_X1 U12983 ( .A1(n13605), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10321) );
  NAND2_X1 U12984 ( .A1(n10322), .A2(n13608), .ZN(n13930) );
  NAND2_X1 U12985 ( .A1(n13931), .A2(n13605), .ZN(n10322) );
  NAND3_X1 U12986 ( .A1(n13237), .A2(n13314), .A3(n13269), .ZN(n13312) );
  NAND2_X1 U12987 ( .A1(n14887), .A2(n10345), .ZN(n10337) );
  OAI211_X1 U12988 ( .C1(n14887), .C2(n10340), .A(n10337), .B(n10339), .ZN(
        n14871) );
  NAND2_X1 U12989 ( .A1(n11363), .A2(n10350), .ZN(n10348) );
  INV_X1 U12990 ( .A(n12792), .ZN(n11632) );
  CLKBUF_X1 U12992 ( .A(n14213), .Z(n14306) );
  NAND2_X1 U12993 ( .A1(n11698), .A2(n11697), .ZN(n11700) );
  INV_X1 U12994 ( .A(n12931), .ZN(n11847) );
  NAND2_X1 U12995 ( .A1(n14730), .A2(n12740), .ZN(n11626) );
  AOI22_X1 U12996 ( .A1(n11578), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12147), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11568) );
  NAND2_X1 U12997 ( .A1(n13604), .A2(n13615), .ZN(n13605) );
  NAND2_X1 U12998 ( .A1(n20101), .A2(n13079), .ZN(n14326) );
  AOI22_X1 U12999 ( .A1(n11233), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10846), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10494) );
  AND2_X1 U13000 ( .A1(n11233), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10443) );
  NAND2_X1 U13001 ( .A1(n14433), .A2(n10356), .ZN(n12398) );
  OAI22_X1 U13002 ( .A1(n9823), .A2(n10942), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n11032), .ZN(n10947) );
  INV_X1 U13003 ( .A(n12868), .ZN(n12869) );
  NOR2_X1 U13004 ( .A1(n20559), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10355) );
  AND2_X1 U13005 ( .A1(n14391), .A2(n20286), .ZN(n10356) );
  OR2_X1 U13006 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15235), .ZN(
        n10357) );
  AND2_X1 U13007 ( .A1(n13207), .A2(n19247), .ZN(n10358) );
  INV_X1 U13008 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19935) );
  INV_X1 U13009 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15663) );
  AND2_X1 U13010 ( .A1(n10489), .A2(n10488), .ZN(n10359) );
  NOR2_X1 U13011 ( .A1(n13643), .A2(n13647), .ZN(n15665) );
  OR3_X1 U13012 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n17606), .ZN(n10360) );
  INV_X1 U13013 ( .A(n19912), .ZN(n19978) );
  AND2_X1 U13014 ( .A1(n10816), .A2(n10815), .ZN(n10361) );
  AND2_X1 U13015 ( .A1(n10826), .A2(n10825), .ZN(n10362) );
  AND2_X1 U13016 ( .A1(n10493), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10363) );
  NAND2_X1 U13017 ( .A1(n17722), .A2(n17894), .ZN(n17633) );
  INV_X1 U13018 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11710) );
  INV_X2 U13019 ( .A(n17261), .ZN(n17246) );
  OR2_X1 U13020 ( .A1(n19040), .A2(n19909), .ZN(n10364) );
  INV_X1 U13021 ( .A(n13204), .ZN(n13189) );
  AND3_X1 U13022 ( .A1(n10814), .A2(n10861), .A3(n10813), .ZN(n10365) );
  AND2_X1 U13023 ( .A1(n11339), .A2(n11343), .ZN(n10366) );
  INV_X1 U13024 ( .A(n11136), .ZN(n13417) );
  OR2_X1 U13025 ( .A1(n10767), .A2(n10766), .ZN(n11136) );
  INV_X1 U13026 ( .A(n13154), .ZN(n19231) );
  NAND3_X2 U13027 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19923), .A3(n19758), 
        .ZN(n13154) );
  INV_X1 U13028 ( .A(n10469), .ZN(n10773) );
  AND2_X1 U13029 ( .A1(n13091), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10367) );
  AND4_X1 U13030 ( .A1(n11586), .A2(n11585), .A3(n11584), .A4(n11583), .ZN(
        n10368) );
  AND4_X1 U13031 ( .A1(n11582), .A2(n11581), .A3(n11580), .A4(n11579), .ZN(
        n10369) );
  NAND2_X1 U13032 ( .A1(n11625), .A2(n12763), .ZN(n10370) );
  AND3_X1 U13033 ( .A1(n11577), .A2(n13079), .A3(n11645), .ZN(n10371) );
  NAND2_X1 U13034 ( .A1(n20101), .A2(n20286), .ZN(n14316) );
  AND2_X1 U13035 ( .A1(n16363), .A2(n10953), .ZN(n10372) );
  AOI21_X1 U13036 ( .B1(n9836), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10489) );
  NAND2_X1 U13037 ( .A1(n13367), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n13211) );
  OR3_X1 U13038 ( .A1(n12348), .A2(n12347), .A3(n12368), .ZN(n12349) );
  AOI22_X1 U13039 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11571) );
  INV_X1 U13040 ( .A(n11317), .ZN(n11318) );
  OAI22_X1 U13041 ( .A1(n10863), .A2(n10860), .B1(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n19946), .ZN(n10865) );
  OR2_X1 U13042 ( .A1(n11788), .A2(n11787), .ZN(n13345) );
  OAI21_X1 U13043 ( .B1(n20263), .B2(n15872), .A(n12825), .ZN(n11648) );
  NAND2_X1 U13044 ( .A1(n10902), .A2(n9818), .ZN(n10903) );
  AOI22_X1 U13045 ( .A1(n13368), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13190), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13196) );
  AOI22_X1 U13046 ( .A1(n9839), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(n9836), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10431) );
  OAI21_X1 U13047 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18851), .A(
        n13676), .ZN(n13677) );
  INV_X1 U13048 ( .A(n12332), .ZN(n12329) );
  NOR2_X1 U13049 ( .A1(n11751), .A2(n13499), .ZN(n13495) );
  AND2_X1 U13050 ( .A1(n14324), .A2(n14240), .ZN(n11966) );
  INV_X1 U13051 ( .A(n13415), .ZN(n11887) );
  INV_X1 U13052 ( .A(n13290), .ZN(n11873) );
  INV_X1 U13053 ( .A(n13487), .ZN(n13499) );
  AND2_X1 U13054 ( .A1(n11720), .A2(n20233), .ZN(n11724) );
  INV_X1 U13055 ( .A(n10558), .ZN(n10723) );
  INV_X1 U13056 ( .A(n13615), .ZN(n13602) );
  INV_X1 U13057 ( .A(n19252), .ZN(n12652) );
  AND2_X1 U13058 ( .A1(n10829), .A2(n10828), .ZN(n10833) );
  NAND2_X1 U13059 ( .A1(n10859), .A2(n10858), .ZN(n10863) );
  AND2_X1 U13060 ( .A1(n13763), .A2(n13764), .ZN(n13675) );
  AOI22_X1 U13061 ( .A1(n12249), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11561), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11595) );
  AND2_X1 U13062 ( .A1(n12325), .A2(n12324), .ZN(n12370) );
  INV_X1 U13063 ( .A(n11812), .ZN(n11978) );
  INV_X1 U13064 ( .A(n14214), .ZN(n12002) );
  INV_X1 U13065 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11961) );
  INV_X1 U13066 ( .A(n12930), .ZN(n11846) );
  INV_X1 U13067 ( .A(n12378), .ZN(n11620) );
  NAND2_X1 U13068 ( .A1(n10379), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10374) );
  NAND2_X1 U13069 ( .A1(n19041), .A2(n13835), .ZN(n13841) );
  INV_X1 U13070 ( .A(n13947), .ZN(n11079) );
  AND2_X1 U13071 ( .A1(n13296), .A2(n13294), .ZN(n11135) );
  AND2_X1 U13072 ( .A1(n13280), .A2(n13281), .ZN(n11134) );
  NAND2_X1 U13073 ( .A1(n10920), .A2(n12679), .ZN(n12399) );
  OR2_X1 U13074 ( .A1(n11338), .A2(n11340), .ZN(n11343) );
  AOI221_X1 U13075 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n10870), 
        .C1(n15663), .C2(n10870), .A(n10869), .ZN(n11449) );
  NAND2_X1 U13076 ( .A1(n10852), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10853) );
  AOI21_X1 U13077 ( .B1(n18699), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n13675), .ZN(n13684) );
  AOI21_X1 U13078 ( .B1(n12325), .B2(n12322), .A(n12324), .ZN(n12372) );
  NAND2_X1 U13079 ( .A1(n20059), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14253) );
  OR2_X1 U13080 ( .A1(n14288), .A2(n14287), .ZN(n12090) );
  NAND2_X1 U13081 ( .A1(n10058), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12311) );
  NOR2_X1 U13082 ( .A1(n13079), .A2(n20898), .ZN(n11812) );
  AND2_X1 U13083 ( .A1(n20898), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12314) );
  NOR2_X1 U13084 ( .A1(n12201), .A2(n14485), .ZN(n12202) );
  INV_X1 U13085 ( .A(n11844), .ZN(n13425) );
  NOR2_X1 U13086 ( .A1(n12053), .A2(n14533), .ZN(n12054) );
  AND2_X1 U13087 ( .A1(n14328), .A2(n13435), .ZN(n13494) );
  INV_X1 U13088 ( .A(n14601), .ZN(n14428) );
  OR2_X1 U13089 ( .A1(n12782), .A2(n12778), .ZN(n12779) );
  NAND2_X1 U13090 ( .A1(n11645), .A2(n14328), .ZN(n11629) );
  INV_X1 U13091 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n15858) );
  XNOR2_X1 U13092 ( .A(n11836), .B(n11835), .ZN(n12739) );
  OAI211_X1 U13093 ( .C1(n16192), .C2(P1_STATE2_REG_2__SCAN_IN), .A(n15882), 
        .B(n20826), .ZN(n20230) );
  NAND2_X1 U13094 ( .A1(n13308), .A2(n13309), .ZN(n13381) );
  AND2_X1 U13095 ( .A1(n11035), .A2(n11034), .ZN(n14916) );
  AND2_X1 U13096 ( .A1(n11275), .A2(n11293), .ZN(n11291) );
  INV_X1 U13097 ( .A(n10603), .ZN(n11225) );
  INV_X1 U13098 ( .A(n13300), .ZN(n13419) );
  AND2_X1 U13099 ( .A1(n10995), .A2(n10994), .ZN(n12945) );
  AND2_X1 U13100 ( .A1(n18909), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12597) );
  INV_X1 U13101 ( .A(n15473), .ZN(n15316) );
  NOR2_X1 U13103 ( .A1(n13826), .A2(n15501), .ZN(n15485) );
  INV_X1 U13104 ( .A(n17685), .ZN(n16387) );
  NAND2_X1 U13105 ( .A1(n15778), .A2(n15837), .ZN(n15776) );
  INV_X1 U13106 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n15756) );
  OAI21_X2 U13107 ( .B1(n18687), .B2(n15806), .A(n18686), .ZN(n18694) );
  AOI21_X1 U13108 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n18716), .A(
        n13678), .ZN(n13765) );
  AND2_X1 U13109 ( .A1(n14028), .A2(n14027), .ZN(n14308) );
  AND2_X1 U13110 ( .A1(n11804), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11888) );
  NAND2_X1 U13111 ( .A1(n11749), .A2(n11748), .ZN(n20389) );
  NOR2_X1 U13112 ( .A1(n14253), .A2(n20231), .ZN(n13450) );
  NAND2_X1 U13113 ( .A1(n12202), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12258) );
  NAND2_X1 U13114 ( .A1(n12179), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12201) );
  INV_X1 U13115 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14513) );
  AND2_X1 U13116 ( .A1(n11967), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11986) );
  AND2_X1 U13117 ( .A1(n11996), .A2(n11933), .ZN(n14403) );
  AND3_X1 U13118 ( .A1(n11886), .A2(n11885), .A3(n11884), .ZN(n13415) );
  NOR2_X1 U13119 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20627) );
  AND2_X1 U13120 ( .A1(n14017), .A2(n14016), .ZN(n14320) );
  NAND2_X1 U13121 ( .A1(n11705), .A2(n11704), .ZN(n20297) );
  AND2_X1 U13122 ( .A1(n20361), .A2(n20360), .ZN(n20363) );
  OR2_X1 U13123 ( .A1(n20471), .A2(n20719), .ZN(n20448) );
  NOR2_X1 U13124 ( .A1(n20766), .A2(n20323), .ZN(n20534) );
  AOI21_X1 U13125 ( .B1(n20686), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20395), 
        .ZN(n20770) );
  AND2_X1 U13126 ( .A1(n10871), .A2(n12492), .ZN(n16348) );
  INV_X1 U13127 ( .A(n19115), .ZN(n11089) );
  OR2_X1 U13128 ( .A1(n10714), .A2(n10713), .ZN(n13280) );
  OAI21_X1 U13129 ( .B1(n11426), .B2(n11425), .A(n11424), .ZN(n11427) );
  INV_X1 U13130 ( .A(n19222), .ZN(n15211) );
  OR2_X1 U13131 ( .A1(n15458), .A2(n13978), .ZN(n15354) );
  INV_X1 U13132 ( .A(n15176), .ZN(n15410) );
  AND3_X1 U13133 ( .A1(n10717), .A2(n10716), .A3(n10715), .ZN(n15452) );
  OR2_X1 U13134 ( .A1(n18908), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19083) );
  AND2_X1 U13135 ( .A1(n12903), .A2(n10234), .ZN(n19939) );
  OR2_X1 U13136 ( .A1(n16365), .A2(n12587), .ZN(n12588) );
  NOR2_X1 U13137 ( .A1(n12645), .A2(n11450), .ZN(n12612) );
  NAND2_X1 U13138 ( .A1(n19522), .A2(n19488), .ZN(n19415) );
  INV_X1 U13139 ( .A(n19922), .ZN(n19598) );
  NAND2_X1 U13140 ( .A1(n18909), .A2(n19832), .ZN(n16363) );
  NOR2_X1 U13141 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16678), .ZN(n16662) );
  NOR2_X1 U13142 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16718), .ZN(n16703) );
  INV_X1 U13143 ( .A(n16953), .ZN(n16724) );
  NOR2_X1 U13144 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16868), .ZN(n16852) );
  INV_X1 U13145 ( .A(n16576), .ZN(n16580) );
  INV_X1 U13146 ( .A(n16926), .ZN(n16951) );
  NOR2_X1 U13147 ( .A1(n13768), .A2(n18688), .ZN(n15801) );
  NAND2_X1 U13148 ( .A1(n17724), .A2(n16387), .ZN(n17682) );
  NOR2_X1 U13149 ( .A1(n15810), .A2(n17390), .ZN(n17819) );
  INV_X1 U13150 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15781) );
  XNOR2_X1 U13151 ( .A(n15757), .B(n15756), .ZN(n17873) );
  INV_X1 U13152 ( .A(n18214), .ZN(n18207) );
  INV_X1 U13153 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18699) );
  INV_X1 U13154 ( .A(n17895), .ZN(n17722) );
  NAND2_X1 U13155 ( .A1(n12087), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12124) );
  AND2_X1 U13156 ( .A1(n20059), .A2(n13431), .ZN(n20031) );
  AND2_X1 U13157 ( .A1(n20059), .A2(n13434), .ZN(n20079) );
  INV_X1 U13158 ( .A(n20558), .ZN(n20726) );
  NAND2_X1 U13159 ( .A1(n12840), .A2(n14012), .ZN(n12823) );
  OR2_X1 U13160 ( .A1(n12841), .A2(n19982), .ZN(n12380) );
  AND2_X1 U13161 ( .A1(n14188), .A2(n14297), .ZN(n15950) );
  NAND2_X1 U13162 ( .A1(n12020), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12053) );
  NAND2_X1 U13163 ( .A1(n11919), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11962) );
  INV_X1 U13164 ( .A(n16041), .ZN(n20151) );
  OR2_X1 U13165 ( .A1(n14669), .A2(n14595), .ZN(n16091) );
  INV_X1 U13166 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12859) );
  NOR2_X2 U13167 ( .A1(n20368), .A2(n20498), .ZN(n20319) );
  OAI21_X1 U13168 ( .B1(n20330), .B2(n20329), .A(n20328), .ZN(n20353) );
  NOR2_X2 U13169 ( .A1(n20368), .A2(n20719), .ZN(n20384) );
  NOR2_X2 U13170 ( .A1(n20368), .A2(n20588), .ZN(n20413) );
  OR2_X1 U13171 ( .A1(n20766), .A2(n20625), .ZN(n20498) );
  INV_X1 U13172 ( .A(n20448), .ZN(n20494) );
  INV_X1 U13173 ( .A(n20504), .ZN(n20525) );
  AND2_X1 U13174 ( .A1(n20590), .A2(n20534), .ZN(n20583) );
  AND2_X1 U13175 ( .A1(n20590), .A2(n20556), .ZN(n20621) );
  INV_X1 U13176 ( .A(n20642), .ZN(n20680) );
  INV_X1 U13177 ( .A(n20323), .ZN(n20625) );
  INV_X1 U13178 ( .A(n20724), .ZN(n20756) );
  NAND2_X1 U13179 ( .A1(n14003), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n15882) );
  INV_X1 U13180 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20843) );
  INV_X1 U13181 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20834) );
  NAND2_X1 U13182 ( .A1(n11090), .A2(n11089), .ZN(n11091) );
  OR2_X1 U13183 ( .A1(n12500), .A2(n10878), .ZN(n19085) );
  INV_X1 U13184 ( .A(n19122), .ZN(n19080) );
  INV_X1 U13185 ( .A(n19105), .ZN(n19089) );
  OR2_X1 U13186 ( .A1(n10746), .A2(n10745), .ZN(n13296) );
  OR2_X1 U13187 ( .A1(n10683), .A2(n10682), .ZN(n13140) );
  AND2_X1 U13188 ( .A1(n12630), .A2(n12570), .ZN(n19128) );
  INV_X1 U13189 ( .A(n19160), .ZN(n19176) );
  INV_X1 U13190 ( .A(n12522), .ZN(n12576) );
  INV_X1 U13191 ( .A(n19225), .ZN(n16283) );
  OAI211_X1 U13192 ( .C1(n14997), .C2(n15000), .A(n14998), .B(n15011), .ZN(
        n13929) );
  AND2_X1 U13193 ( .A1(n13886), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15174) );
  INV_X1 U13194 ( .A(n16313), .ZN(n16299) );
  NAND2_X1 U13195 ( .A1(n12660), .A2(n16362), .ZN(n12681) );
  AND2_X1 U13196 ( .A1(n12588), .A2(n18909), .ZN(n19758) );
  NOR2_X1 U13197 ( .A1(n12612), .A2(n19938), .ZN(n16365) );
  NOR2_X2 U13198 ( .A1(n19292), .A2(n19415), .ZN(n19341) );
  INV_X1 U13199 ( .A(n19422), .ZN(n19436) );
  AND2_X1 U13200 ( .A1(n19522), .A2(n19958), .ZN(n19376) );
  NOR2_X2 U13201 ( .A1(n13156), .A2(n19415), .ZN(n19516) );
  AND2_X1 U13202 ( .A1(n19936), .A2(n19949), .ZN(n19530) );
  AND2_X1 U13203 ( .A1(n19670), .A2(n19530), .ZN(n19587) );
  NOR2_X1 U13204 ( .A1(n19556), .A2(n19598), .ZN(n19619) );
  INV_X1 U13205 ( .A(n19808), .ZN(n19651) );
  NOR2_X1 U13206 ( .A1(n19664), .A2(n19663), .ZN(n19685) );
  AND2_X1 U13207 ( .A1(n10902), .A2(n19275), .ZN(n19713) );
  AND2_X1 U13208 ( .A1(n10930), .A2(n19275), .ZN(n19737) );
  INV_X1 U13209 ( .A(n19718), .ZN(n19782) );
  INV_X1 U13210 ( .A(n19800), .ZN(n19815) );
  NOR2_X1 U13211 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n18909), .ZN(n19829) );
  INV_X1 U13212 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19848) );
  INV_X1 U13213 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19856) );
  INV_X1 U13214 ( .A(n18037), .ZN(n18677) );
  NOR2_X1 U13215 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16765), .ZN(n16756) );
  NOR4_X1 U13216 ( .A1(n16915), .A2(n18788), .A3(n18785), .A4(n16786), .ZN(
        n16763) );
  NOR2_X1 U13217 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16839), .ZN(n16828) );
  NOR2_X1 U13218 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16893), .ZN(n16879) );
  INV_X1 U13219 ( .A(n18201), .ZN(n17990) );
  INV_X1 U13220 ( .A(n16955), .ZN(n16947) );
  AOI21_X1 U13221 ( .B1(n18671), .B2(n18670), .A(n17414), .ZN(n18886) );
  INV_X1 U13222 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17235) );
  INV_X1 U13223 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17241) );
  NAND2_X1 U13224 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17331), .ZN(n17330) );
  NOR2_X1 U13225 ( .A1(n18013), .A2(n17693), .ZN(n17610) );
  NOR2_X1 U13226 ( .A1(n15835), .A2(n17795), .ZN(n17744) );
  INV_X1 U13227 ( .A(n17894), .ZN(n17844) );
  NOR2_X1 U13228 ( .A1(n18889), .A2(n16558), .ZN(n17887) );
  NAND2_X1 U13229 ( .A1(n18112), .A2(n18104), .ZN(n18132) );
  NOR2_X1 U13230 ( .A1(n18099), .A2(n18058), .ZN(n17707) );
  NOR2_X1 U13231 ( .A1(n17990), .A2(n18214), .ZN(n18209) );
  NOR2_X1 U13232 ( .A1(n16441), .A2(n18207), .ZN(n18205) );
  INV_X1 U13233 ( .A(n18333), .ZN(n18326) );
  INV_X1 U13234 ( .A(n18355), .ZN(n18346) );
  INV_X1 U13235 ( .A(n18378), .ZN(n18371) );
  INV_X1 U13236 ( .A(n18449), .ZN(n18441) );
  INV_X1 U13237 ( .A(n18444), .ZN(n18468) );
  INV_X1 U13238 ( .A(n18517), .ZN(n18510) );
  INV_X1 U13239 ( .A(n18560), .ZN(n18569) );
  INV_X1 U13240 ( .A(n18601), .ZN(n18603) );
  INV_X1 U13241 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18847) );
  INV_X1 U13242 ( .A(n13155), .ZN(n13153) );
  NOR2_X1 U13243 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12411), .ZN(n16538)
         );
  NAND2_X1 U13244 ( .A1(n12765), .A2(n14005), .ZN(n13423) );
  NAND2_X1 U13245 ( .A1(n13424), .A2(n13423), .ZN(n20904) );
  INV_X1 U13246 ( .A(n20031), .ZN(n15937) );
  INV_X1 U13247 ( .A(n20077), .ZN(n20073) );
  NAND2_X2 U13248 ( .A1(n12823), .A2(n12822), .ZN(n20101) );
  OAI211_X2 U13249 ( .C1(n12381), .C2(n13423), .A(n12380), .B(n12379), .ZN(
        n14391) );
  INV_X1 U13250 ( .A(n20105), .ZN(n20134) );
  NOR2_X1 U13251 ( .A1(n13423), .A2(n12966), .ZN(n13021) );
  INV_X1 U13252 ( .A(n20147), .ZN(n13034) );
  OR2_X1 U13253 ( .A1(n20159), .A2(n12737), .ZN(n16041) );
  INV_X1 U13254 ( .A(n16037), .ZN(n20164) );
  NAND2_X1 U13255 ( .A1(n12795), .A2(n12794), .ZN(n20171) );
  INV_X1 U13256 ( .A(n20208), .ZN(n20196) );
  INV_X1 U13257 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20686) );
  AOI211_X2 U13258 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20391), .A(n20327), 
        .B(n20226), .ZN(n20296) );
  OR2_X1 U13259 ( .A1(n20368), .A2(n20692), .ZN(n20351) );
  AOI22_X1 U13260 ( .A1(n20326), .A2(n20329), .B1(n10355), .B2(n20561), .ZN(
        n20356) );
  INV_X1 U13261 ( .A(n20362), .ZN(n20388) );
  OR2_X1 U13262 ( .A1(n20471), .A2(n20498), .ZN(n20440) );
  AOI22_X1 U13263 ( .A1(n20446), .A2(n20443), .B1(n20633), .B2(n10355), .ZN(
        n20468) );
  OR2_X1 U13264 ( .A1(n20471), .A2(n20588), .ZN(n20504) );
  NAND2_X1 U13265 ( .A1(n20590), .A2(n20499), .ZN(n20554) );
  AOI22_X1 U13266 ( .A1(n20566), .A2(n20562), .B1(n20561), .B2(n20560), .ZN(
        n20587) );
  NAND2_X1 U13267 ( .A1(n20590), .A2(n20589), .ZN(n20642) );
  AOI22_X1 U13268 ( .A1(n20639), .A2(n20636), .B1(n20633), .B2(n20632), .ZN(
        n20685) );
  OR2_X1 U13269 ( .A1(n20626), .A2(n20625), .ZN(n20718) );
  OR2_X1 U13270 ( .A1(n20769), .A2(n20588), .ZN(n20807) );
  OR2_X1 U13271 ( .A1(n20769), .A2(n20719), .ZN(n20824) );
  INV_X1 U13272 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n16192) );
  INV_X1 U13273 ( .A(n20888), .ZN(n20829) );
  OR2_X1 U13274 ( .A1(n10874), .A2(n12471), .ZN(n12500) );
  INV_X1 U13275 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19924) );
  AND2_X1 U13276 ( .A1(n11092), .A2(n11091), .ZN(n11093) );
  INV_X1 U13277 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18959) );
  OR3_X1 U13278 ( .A1(n18911), .A2(n19223), .A3(n10873), .ZN(n19122) );
  OAI21_X1 U13279 ( .B1(n12690), .B2(n12692), .A(n12691), .ZN(n19936) );
  AND2_X1 U13280 ( .A1(n11471), .A2(n16362), .ZN(n19160) );
  INV_X1 U13281 ( .A(n19137), .ZN(n19181) );
  INV_X1 U13282 ( .A(n19186), .ZN(n19220) );
  INV_X1 U13283 ( .A(n12502), .ZN(n12522) );
  INV_X1 U13284 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18995) );
  INV_X1 U13285 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16288) );
  AOI211_X1 U13286 ( .C1(n15242), .C2(n16301), .A(n15241), .B(n15240), .ZN(
        n15243) );
  OR2_X1 U13287 ( .A1(n12681), .A2(n19967), .ZN(n15495) );
  NAND2_X1 U13288 ( .A1(n19530), .A2(n19376), .ZN(n19319) );
  NAND2_X1 U13289 ( .A1(n19376), .A2(n19922), .ZN(n19374) );
  AND2_X1 U13290 ( .A1(n19410), .A2(n19409), .ZN(n19422) );
  INV_X1 U13291 ( .A(n19429), .ZN(n19439) );
  NAND2_X1 U13292 ( .A1(n19376), .A2(n19753), .ZN(n19487) );
  AOI211_X2 U13293 ( .C1(n19493), .C2(n19494), .A(n19492), .B(n19665), .ZN(
        n19521) );
  INV_X1 U13294 ( .A(n19587), .ZN(n19557) );
  INV_X1 U13295 ( .A(n19619), .ZN(n19614) );
  NAND2_X1 U13296 ( .A1(n19690), .A2(n19669), .ZN(n19689) );
  NAND2_X1 U13297 ( .A1(n19670), .A2(n19669), .ZN(n19735) );
  INV_X1 U13298 ( .A(n19726), .ZN(n19801) );
  INV_X1 U13299 ( .A(n19921), .ZN(n19834) );
  INV_X1 U13300 ( .A(n19978), .ZN(n19868) );
  NAND2_X1 U13301 ( .A1(n18882), .A2(n18722), .ZN(n16558) );
  NOR2_X1 U13302 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16696), .ZN(n16693) );
  INV_X1 U13303 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17750) );
  INV_X1 U13304 ( .A(n16873), .ZN(n16942) );
  AND2_X1 U13305 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17138), .ZN(n17140) );
  NOR2_X1 U13306 ( .A1(n15649), .A2(n17236), .ZN(n17226) );
  NOR2_X1 U13307 ( .A1(n17260), .A2(n15648), .ZN(n17244) );
  INV_X1 U13308 ( .A(n17340), .ZN(n17316) );
  NOR2_X1 U13309 ( .A1(n17453), .A2(n17371), .ZN(n17375) );
  NOR2_X1 U13310 ( .A1(n15697), .A2(n15696), .ZN(n17397) );
  INV_X1 U13311 ( .A(n17442), .ZN(n17470) );
  INV_X1 U13312 ( .A(n17521), .ZN(n17518) );
  NAND2_X1 U13313 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17889), .ZN(n17728) );
  INV_X1 U13314 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17758) );
  NAND2_X1 U13315 ( .A1(n16392), .A2(n9816), .ZN(n17803) );
  OAI21_X1 U13316 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18881), .A(n16558), 
        .ZN(n17894) );
  INV_X1 U13317 ( .A(n18209), .ZN(n18194) );
  INV_X1 U13318 ( .A(n18138), .ZN(n18124) );
  INV_X1 U13319 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18518) );
  INV_X1 U13320 ( .A(n18393), .ZN(n18400) );
  INV_X1 U13321 ( .A(n18649), .ZN(n18597) );
  NAND2_X1 U13322 ( .A1(n16574), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18732) );
  INV_X1 U13323 ( .A(n18833), .ZN(n18830) );
  INV_X1 U13324 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18758) );
  NAND2_X1 U13325 ( .A1(n12398), .A2(n12397), .ZN(P1_U2873) );
  INV_X1 U13326 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16272) );
  NAND2_X1 U13327 ( .A1(n10411), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10415) );
  NAND2_X1 U13328 ( .A1(n10396), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10395) );
  INV_X1 U13329 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15110) );
  INV_X1 U13330 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15070) );
  INV_X1 U13331 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16206) );
  INV_X1 U13332 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15039) );
  INV_X1 U13333 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10380) );
  XNOR2_X1 U13334 ( .A(n10374), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15006) );
  INV_X1 U13335 ( .A(n10374), .ZN(n10375) );
  NAND2_X1 U13336 ( .A1(n10375), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10377) );
  INV_X1 U13337 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n10376) );
  NAND2_X1 U13338 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13945) );
  OR2_X1 U13339 ( .A1(n10379), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10378) );
  AND2_X1 U13340 ( .A1(n10378), .A2(n10374), .ZN(n15017) );
  INV_X1 U13341 ( .A(n10379), .ZN(n10382) );
  NAND2_X1 U13342 ( .A1(n10384), .A2(n10380), .ZN(n10381) );
  NAND2_X1 U13343 ( .A1(n10382), .A2(n10381), .ZN(n15031) );
  INV_X1 U13344 ( .A(n15031), .ZN(n16195) );
  NAND2_X1 U13345 ( .A1(n10387), .A2(n15039), .ZN(n10383) );
  AND2_X1 U13346 ( .A1(n10384), .A2(n10383), .ZN(n15041) );
  NAND2_X1 U13347 ( .A1(n10385), .A2(n16206), .ZN(n10386) );
  NAND2_X1 U13348 ( .A1(n10387), .A2(n10386), .ZN(n15050) );
  INV_X1 U13349 ( .A(n15050), .ZN(n16215) );
  OAI21_X1 U13350 ( .B1(n9934), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n10385), .ZN(n15062) );
  INV_X1 U13351 ( .A(n15062), .ZN(n16226) );
  AOI21_X1 U13352 ( .B1(n15070), .B2(n10389), .A(n9934), .ZN(n15072) );
  OAI21_X1 U13353 ( .B1(n10388), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n10389), .ZN(n10390) );
  INV_X1 U13354 ( .A(n10390), .ZN(n15079) );
  INV_X1 U13355 ( .A(n10388), .ZN(n10394) );
  INV_X1 U13356 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11054) );
  INV_X1 U13357 ( .A(n10391), .ZN(n10392) );
  NAND2_X1 U13358 ( .A1(n11054), .A2(n10392), .ZN(n10393) );
  NAND2_X1 U13359 ( .A1(n10394), .A2(n10393), .ZN(n15092) );
  INV_X1 U13360 ( .A(n15092), .ZN(n12414) );
  AOI21_X1 U13361 ( .B1(n15110), .B2(n10395), .A(n10391), .ZN(n15112) );
  OAI21_X1 U13362 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n10396), .A(
        n10395), .ZN(n15120) );
  INV_X1 U13363 ( .A(n15120), .ZN(n18938) );
  OAI21_X1 U13364 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n10419), .A(
        n10397), .ZN(n15140) );
  INV_X1 U13365 ( .A(n15140), .ZN(n18962) );
  OR2_X1 U13366 ( .A1(n10398), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10399) );
  NAND2_X1 U13367 ( .A1(n10399), .A2(n10420), .ZN(n15164) );
  INV_X1 U13368 ( .A(n15164), .ZN(n18985) );
  OAI21_X1 U13369 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n10400), .A(
        n10401), .ZN(n15178) );
  INV_X1 U13370 ( .A(n15178), .ZN(n19008) );
  OAI21_X1 U13371 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n10414), .A(
        n10402), .ZN(n15187) );
  INV_X1 U13372 ( .A(n15187), .ZN(n19031) );
  OAI21_X1 U13373 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n10411), .A(
        n10415), .ZN(n19060) );
  INV_X1 U13374 ( .A(n19060), .ZN(n10413) );
  AOI21_X1 U13375 ( .B1(n16288), .B2(n10409), .A(n10410), .ZN(n19067) );
  AOI21_X1 U13376 ( .B1(n16295), .B2(n10407), .A(n10403), .ZN(n19099) );
  AOI21_X1 U13377 ( .B1(n19235), .B2(n10405), .A(n10408), .ZN(n19221) );
  AOI21_X1 U13378 ( .B1(n14806), .B2(n10404), .A(n10406), .ZN(n13806) );
  AOI22_X1 U13379 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18909), .ZN(n14815) );
  AOI22_X1 U13380 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n14806), .B2(n18909), .ZN(
        n14805) );
  NAND2_X1 U13381 ( .A1(n14815), .A2(n14805), .ZN(n14804) );
  NOR2_X1 U13382 ( .A1(n13806), .A2(n14804), .ZN(n13522) );
  OAI21_X1 U13383 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n10406), .A(
        n10405), .ZN(n13523) );
  NAND2_X1 U13384 ( .A1(n13522), .A2(n13523), .ZN(n13548) );
  NOR2_X1 U13385 ( .A1(n19221), .A2(n13548), .ZN(n19110) );
  OAI21_X1 U13386 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n10408), .A(
        n10407), .ZN(n19113) );
  NAND2_X1 U13387 ( .A1(n19110), .A2(n19113), .ZN(n19097) );
  NOR2_X1 U13388 ( .A1(n19099), .A2(n19097), .ZN(n19077) );
  OAI21_X1 U13389 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n10403), .A(
        n10409), .ZN(n19079) );
  NAND2_X1 U13390 ( .A1(n19077), .A2(n19079), .ZN(n19065) );
  NOR2_X1 U13391 ( .A1(n19067), .A2(n19065), .ZN(n14794) );
  AOI21_X1 U13392 ( .B1(n16272), .B2(n10169), .A(n10411), .ZN(n16263) );
  INV_X1 U13393 ( .A(n16263), .ZN(n10412) );
  NAND2_X1 U13394 ( .A1(n14794), .A2(n10412), .ZN(n19058) );
  NOR2_X1 U13395 ( .A1(n10413), .A2(n19058), .ZN(n19046) );
  AOI21_X1 U13396 ( .B1(n19042), .B2(n10415), .A(n10414), .ZN(n19047) );
  INV_X1 U13397 ( .A(n19047), .ZN(n10416) );
  NAND2_X1 U13398 ( .A1(n19046), .A2(n10416), .ZN(n19029) );
  NOR2_X1 U13399 ( .A1(n19031), .A2(n19029), .ZN(n19021) );
  AOI21_X1 U13400 ( .B1(n19017), .B2(n10402), .A(n10400), .ZN(n19022) );
  INV_X1 U13401 ( .A(n19022), .ZN(n10417) );
  NAND2_X1 U13402 ( .A1(n19021), .A2(n10417), .ZN(n19006) );
  NOR2_X1 U13403 ( .A1(n19008), .A2(n19006), .ZN(n18998) );
  AOI21_X1 U13404 ( .B1(n18995), .B2(n10401), .A(n10398), .ZN(n19000) );
  INV_X1 U13405 ( .A(n19000), .ZN(n10418) );
  NAND2_X1 U13406 ( .A1(n18998), .A2(n10418), .ZN(n18983) );
  NOR2_X1 U13407 ( .A1(n18985), .A2(n18983), .ZN(n18973) );
  AOI21_X1 U13408 ( .B1(n18982), .B2(n10420), .A(n10419), .ZN(n10421) );
  INV_X1 U13409 ( .A(n10421), .ZN(n18975) );
  NAND2_X1 U13410 ( .A1(n18973), .A2(n18975), .ZN(n18960) );
  NOR2_X1 U13411 ( .A1(n18962), .A2(n18960), .ZN(n18950) );
  AOI21_X1 U13412 ( .B1(n10397), .B2(n18959), .A(n10396), .ZN(n18952) );
  INV_X1 U13413 ( .A(n18952), .ZN(n10422) );
  NAND2_X1 U13414 ( .A1(n18950), .A2(n10422), .ZN(n18937) );
  NOR2_X1 U13415 ( .A1(n18938), .A2(n18937), .ZN(n18936) );
  NOR2_X1 U13416 ( .A1(n15112), .A2(n14780), .ZN(n14779) );
  NOR2_X1 U13417 ( .A1(n10145), .A2(n16213), .ZN(n12440) );
  NOR2_X1 U13418 ( .A1(n10145), .A2(n14775), .ZN(n10423) );
  NOR2_X1 U13419 ( .A1(n15006), .A2(n10423), .ZN(n14756) );
  INV_X1 U13420 ( .A(n14756), .ZN(n10425) );
  INV_X1 U13421 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19825) );
  NAND4_X1 U13422 ( .A1(n19825), .A2(n18909), .A3(n19924), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19831) );
  NAND2_X1 U13423 ( .A1(n10425), .A2(n10424), .ZN(n11094) );
  AND2_X4 U13424 ( .A1(n15532), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11233) );
  AOI22_X1 U13425 ( .A1(n11233), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9844), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10430) );
  AND2_X4 U13426 ( .A1(n10478), .A2(n16329), .ZN(n10844) );
  AND2_X4 U13427 ( .A1(n12862), .A2(n16329), .ZN(n10843) );
  AOI22_X1 U13428 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10843), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10429) );
  NOR2_X2 U13429 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10427) );
  AOI22_X1 U13430 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10845), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10428) );
  NAND4_X1 U13431 ( .A1(n10431), .A2(n10430), .A3(n10429), .A4(n10428), .ZN(
        n10432) );
  AOI22_X1 U13432 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n10843), .ZN(n10437) );
  AOI22_X1 U13433 ( .A1(n11233), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9844), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10436) );
  AOI22_X1 U13434 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10845), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10435) );
  NAND4_X1 U13435 ( .A1(n10437), .A2(n10436), .A3(n10435), .A4(n10434), .ZN(
        n10438) );
  AOI22_X1 U13436 ( .A1(n9836), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(n9839), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10441) );
  AND2_X1 U13437 ( .A1(n10441), .A2(n10861), .ZN(n10447) );
  NOR2_X1 U13438 ( .A1(n10443), .A2(n10442), .ZN(n10446) );
  AOI22_X1 U13439 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10843), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10444) );
  NAND4_X1 U13440 ( .A1(n10447), .A2(n10446), .A3(n10445), .A4(n10444), .ZN(
        n10455) );
  AOI21_X1 U13441 ( .B1(n9836), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n10861), .ZN(n10449) );
  NAND2_X1 U13442 ( .A1(n9839), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10448) );
  AOI22_X1 U13443 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9838), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10452) );
  AOI22_X1 U13444 ( .A1(n11233), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9844), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10451) );
  AOI22_X1 U13445 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10843), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10450) );
  AOI22_X1 U13446 ( .A1(n9844), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11233), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10459) );
  AOI22_X1 U13447 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10843), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10458) );
  AOI22_X1 U13448 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n9836), .B1(n9840), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10457) );
  AOI22_X1 U13449 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10846), .B1(
        n10845), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10456) );
  NAND4_X1 U13450 ( .A1(n10459), .A2(n10458), .A3(n10457), .A4(n10456), .ZN(
        n10460) );
  AOI22_X1 U13451 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10843), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10464) );
  AOI22_X1 U13452 ( .A1(n11233), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9843), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10463) );
  AOI22_X1 U13453 ( .A1(n9836), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9840), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10462) );
  AOI22_X1 U13454 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10845), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10461) );
  NAND4_X1 U13455 ( .A1(n10464), .A2(n10463), .A3(n10462), .A4(n10461), .ZN(
        n10465) );
  INV_X1 U13456 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n15003) );
  NAND2_X1 U13457 ( .A1(n13954), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10471) );
  NOR2_X1 U13458 ( .A1(n10930), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10507) );
  NAND2_X1 U13459 ( .A1(n13955), .A2(P2_EAX_REG_30__SCAN_IN), .ZN(n10470) );
  OAI211_X1 U13460 ( .C1(n13958), .C2(n15003), .A(n10471), .B(n10470), .ZN(
        n10798) );
  INV_X1 U13461 ( .A(n10798), .ZN(n10800) );
  NAND3_X1 U13462 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12481) );
  INV_X1 U13463 ( .A(n12481), .ZN(n10472) );
  AOI22_X1 U13464 ( .A1(n10537), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10558), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10477) );
  AND2_X2 U13465 ( .A1(n10473), .A2(n10861), .ZN(n11253) );
  AOI22_X1 U13466 ( .A1(n11265), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11253), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10476) );
  AOI22_X1 U13467 ( .A1(n10603), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9887), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10475) );
  AND2_X2 U13468 ( .A1(n11420), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10594) );
  AOI22_X1 U13469 ( .A1(n10594), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10536), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10474) );
  NAND4_X1 U13470 ( .A1(n10477), .A2(n10476), .A3(n10475), .A4(n10474), .ZN(
        n10485) );
  AND2_X2 U13471 ( .A1(n11408), .A2(n10861), .ZN(n11264) );
  AND2_X2 U13472 ( .A1(n11420), .A2(n10861), .ZN(n10553) );
  AOI22_X1 U13473 ( .A1(n11264), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10553), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10483) );
  NAND2_X1 U13474 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11234) );
  INV_X1 U13475 ( .A(n11234), .ZN(n10479) );
  AOI22_X1 U13476 ( .A1(n11257), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11255), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10482) );
  AND2_X2 U13477 ( .A1(n10845), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10648) );
  AOI22_X1 U13478 ( .A1(n11254), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10481) );
  AND2_X2 U13479 ( .A1(n11419), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11166) );
  AOI22_X1 U13480 ( .A1(n11166), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11256), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10480) );
  NAND4_X1 U13481 ( .A1(n10483), .A2(n10482), .A3(n10481), .A4(n10480), .ZN(
        n10484) );
  NOR2_X1 U13482 ( .A1(n10485), .A2(n10484), .ZN(n13228) );
  INV_X1 U13483 ( .A(n13228), .ZN(n10487) );
  NAND2_X1 U13484 ( .A1(n9839), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10488) );
  AOI22_X1 U13485 ( .A1(n11233), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9844), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10492) );
  AOI22_X1 U13486 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10843), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10491) );
  AOI22_X1 U13487 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10845), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10490) );
  NAND4_X1 U13488 ( .A1(n10359), .A2(n10492), .A3(n10491), .A4(n10490), .ZN(
        n10498) );
  AOI22_X1 U13489 ( .A1(n9842), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(n9843), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10493) );
  AOI22_X1 U13490 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10843), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10496) );
  NAND4_X1 U13491 ( .A1(n10363), .A2(n10496), .A3(n10495), .A4(n10494), .ZN(
        n10497) );
  AND2_X2 U13492 ( .A1(n10498), .A2(n10497), .ZN(n10899) );
  NAND2_X1 U13493 ( .A1(n10469), .A2(n10499), .ZN(n10544) );
  INV_X1 U13494 ( .A(n10522), .ZN(n10500) );
  NAND2_X1 U13495 ( .A1(n19964), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19956) );
  NAND2_X1 U13496 ( .A1(n10500), .A2(n19956), .ZN(n10501) );
  AND2_X1 U13497 ( .A1(n10544), .A2(n10501), .ZN(n10502) );
  NAND2_X1 U13498 ( .A1(n10503), .A2(n10502), .ZN(n12633) );
  INV_X1 U13499 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18926) );
  INV_X1 U13500 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12592) );
  NAND2_X1 U13501 ( .A1(n9978), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n10504) );
  OAI211_X1 U13502 ( .C1(n19247), .C2(n12592), .A(n10504), .B(n19938), .ZN(
        n10505) );
  INV_X1 U13503 ( .A(n10505), .ZN(n10506) );
  INV_X1 U13504 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19857) );
  INV_X1 U13505 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15538) );
  NAND2_X1 U13506 ( .A1(n10469), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10509) );
  NAND2_X1 U13507 ( .A1(n10507), .A2(P2_EAX_REG_1__SCAN_IN), .ZN(n10508) );
  OAI211_X1 U13508 ( .C1(n13958), .C2(n19857), .A(n10509), .B(n10508), .ZN(
        n10526) );
  XNOR2_X1 U13509 ( .A(n12632), .B(n10526), .ZN(n12665) );
  AOI22_X1 U13510 ( .A1(n11166), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n11253), .ZN(n10515) );
  AOI22_X1 U13511 ( .A1(n10603), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n11254), .ZN(n10514) );
  AOI22_X1 U13512 ( .A1(n11255), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10558), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10511) );
  NAND2_X1 U13513 ( .A1(n11257), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10510) );
  AND2_X1 U13514 ( .A1(n10511), .A2(n10510), .ZN(n10513) );
  NAND2_X1 U13515 ( .A1(n11256), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10512) );
  NAND4_X1 U13516 ( .A1(n10515), .A2(n10514), .A3(n10513), .A4(n10512), .ZN(
        n10521) );
  AOI22_X1 U13517 ( .A1(n11264), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n10594), .ZN(n10519) );
  AOI22_X1 U13518 ( .A1(n11265), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9887), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10518) );
  AOI22_X1 U13519 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n10536), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10517) );
  AOI22_X1 U13520 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10553), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10516) );
  NAND4_X1 U13521 ( .A1(n10519), .A2(n10518), .A3(n10517), .A4(n10516), .ZN(
        n10520) );
  INV_X1 U13522 ( .A(n13226), .ZN(n10525) );
  NAND2_X1 U13523 ( .A1(n11461), .A2(n10522), .ZN(n10524) );
  NAND2_X1 U13524 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10523) );
  OAI211_X1 U13525 ( .C1(n10748), .C2(n10525), .A(n10524), .B(n10523), .ZN(
        n12664) );
  NOR2_X1 U13526 ( .A1(n12665), .A2(n12664), .ZN(n10528) );
  NOR2_X1 U13527 ( .A1(n12632), .A2(n10526), .ZN(n10527) );
  AOI22_X1 U13528 ( .A1(n11255), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10558), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10531) );
  NAND2_X1 U13529 ( .A1(n11256), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n10530) );
  NAND2_X1 U13530 ( .A1(n11257), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n10529) );
  AND3_X1 U13531 ( .A1(n10531), .A2(n10530), .A3(n10529), .ZN(n10535) );
  AOI22_X1 U13532 ( .A1(n11253), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10534) );
  NAND2_X1 U13533 ( .A1(n10603), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n10533) );
  NAND2_X1 U13534 ( .A1(n11166), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10532) );
  NAND4_X1 U13535 ( .A1(n10535), .A2(n10534), .A3(n10533), .A4(n10532), .ZN(
        n10543) );
  AOI22_X1 U13536 ( .A1(n11264), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10541) );
  AOI22_X1 U13537 ( .A1(n11265), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9887), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10540) );
  AOI22_X1 U13538 ( .A1(n11254), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10536), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10539) );
  AOI22_X1 U13539 ( .A1(n10553), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10538) );
  NAND4_X1 U13540 ( .A1(n10541), .A2(n10540), .A3(n10539), .A4(n10538), .ZN(
        n10542) );
  NAND2_X1 U13541 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10545) );
  OAI211_X1 U13542 ( .C1(n10748), .C2(n13262), .A(n10545), .B(n10544), .ZN(
        n10548) );
  XNOR2_X1 U13543 ( .A(n10549), .B(n10548), .ZN(n12901) );
  INV_X1 U13544 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19860) );
  INV_X2 U13545 ( .A(n10773), .ZN(n13954) );
  NAND2_X1 U13546 ( .A1(n13954), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10547) );
  NAND2_X1 U13547 ( .A1(n13955), .A2(P2_EAX_REG_2__SCAN_IN), .ZN(n10546) );
  OAI211_X1 U13548 ( .C1(n13958), .C2(n19860), .A(n10547), .B(n10546), .ZN(
        n12900) );
  NOR2_X1 U13549 ( .A1(n12901), .A2(n12900), .ZN(n12902) );
  NOR2_X1 U13550 ( .A1(n10549), .A2(n10548), .ZN(n10550) );
  INV_X1 U13551 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n13272) );
  NAND2_X1 U13552 ( .A1(n13954), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10552) );
  NAND2_X1 U13553 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10551) );
  OAI211_X1 U13554 ( .C1(n13958), .C2(n13272), .A(n10552), .B(n10551), .ZN(
        n10569) );
  AOI22_X1 U13555 ( .A1(n11264), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10557) );
  AOI22_X1 U13556 ( .A1(n11265), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9887), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10556) );
  AOI22_X1 U13557 ( .A1(n10603), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11253), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10555) );
  AOI22_X1 U13558 ( .A1(n10553), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10554) );
  NAND4_X1 U13559 ( .A1(n10557), .A2(n10556), .A3(n10555), .A4(n10554), .ZN(
        n10566) );
  AOI22_X1 U13560 ( .A1(n11166), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10536), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10564) );
  AOI22_X1 U13561 ( .A1(n11255), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10558), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10560) );
  NAND2_X1 U13562 ( .A1(n11257), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n10559) );
  AND2_X1 U13563 ( .A1(n10560), .A2(n10559), .ZN(n10563) );
  AOI22_X1 U13564 ( .A1(n11254), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10562) );
  NAND2_X1 U13565 ( .A1(n11256), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n10561) );
  NAND4_X1 U13566 ( .A1(n10564), .A2(n10563), .A3(n10562), .A4(n10561), .ZN(
        n10565) );
  NOR2_X1 U13567 ( .A1(n10566), .A2(n10565), .ZN(n13207) );
  NAND2_X1 U13568 ( .A1(n13955), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n10567) );
  OAI21_X1 U13569 ( .B1(n10748), .B2(n13207), .A(n10567), .ZN(n10568) );
  AOI22_X1 U13570 ( .A1(n13954), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n13955), .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n10586) );
  NAND2_X1 U13571 ( .A1(n10795), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n10585) );
  AOI22_X1 U13572 ( .A1(n11264), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10573) );
  AOI22_X1 U13573 ( .A1(n11265), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9887), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10572) );
  AOI22_X1 U13574 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10536), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10571) );
  AOI22_X1 U13575 ( .A1(n10553), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10570) );
  NAND4_X1 U13576 ( .A1(n10573), .A2(n10572), .A3(n10571), .A4(n10570), .ZN(
        n10583) );
  AOI22_X1 U13577 ( .A1(n11166), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11253), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10581) );
  AOI22_X1 U13578 ( .A1(n10603), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11254), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10580) );
  INV_X1 U13579 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11345) );
  NOR2_X1 U13580 ( .A1(n10756), .A2(n11345), .ZN(n10577) );
  INV_X1 U13581 ( .A(n11255), .ZN(n10752) );
  INV_X1 U13582 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10575) );
  INV_X1 U13583 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10574) );
  OAI22_X1 U13584 ( .A1(n10752), .A2(n10575), .B1(n10574), .B2(n10723), .ZN(
        n10576) );
  NOR2_X1 U13585 ( .A1(n10577), .A2(n10576), .ZN(n10579) );
  NAND2_X1 U13586 ( .A1(n11256), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10578) );
  NAND4_X1 U13587 ( .A1(n10581), .A2(n10580), .A3(n10579), .A4(n10578), .ZN(
        n10582) );
  NAND2_X1 U13588 ( .A1(n10768), .A2(n13315), .ZN(n10584) );
  AOI22_X1 U13589 ( .A1(n10795), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n13954), 
        .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10602) );
  AOI22_X1 U13590 ( .A1(n11255), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10558), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10589) );
  NAND2_X1 U13591 ( .A1(n11256), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10588) );
  NAND2_X1 U13592 ( .A1(n11257), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n10587) );
  AND3_X1 U13593 ( .A1(n10589), .A2(n10588), .A3(n10587), .ZN(n10593) );
  AOI22_X1 U13594 ( .A1(n11253), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10592) );
  NAND2_X1 U13595 ( .A1(n10603), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10591) );
  NAND2_X1 U13596 ( .A1(n11166), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10590) );
  NAND4_X1 U13597 ( .A1(n10593), .A2(n10592), .A3(n10591), .A4(n10590), .ZN(
        n10600) );
  AOI22_X1 U13598 ( .A1(n11264), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10598) );
  AOI22_X1 U13599 ( .A1(n11265), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9887), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10597) );
  AOI22_X1 U13600 ( .A1(n11254), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10536), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10596) );
  AOI22_X1 U13601 ( .A1(n10553), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10595) );
  NAND4_X1 U13602 ( .A1(n10598), .A2(n10597), .A3(n10596), .A4(n10595), .ZN(
        n10599) );
  AOI22_X1 U13603 ( .A1(n10768), .A2(n10884), .B1(n13955), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n10601) );
  NAND2_X1 U13604 ( .A1(n10602), .A2(n10601), .ZN(n13402) );
  AOI22_X1 U13605 ( .A1(n11166), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n11253), .ZN(n10609) );
  AOI22_X1 U13606 ( .A1(n10603), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__6__SCAN_IN), .B2(n11254), .ZN(n10608) );
  AOI22_X1 U13607 ( .A1(n11255), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n10558), .ZN(n10605) );
  NAND2_X1 U13608 ( .A1(n11257), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10604) );
  AND2_X1 U13609 ( .A1(n10605), .A2(n10604), .ZN(n10607) );
  NAND2_X1 U13610 ( .A1(n11256), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n10606) );
  NAND4_X1 U13611 ( .A1(n10609), .A2(n10608), .A3(n10607), .A4(n10606), .ZN(
        n10615) );
  AOI22_X1 U13612 ( .A1(n11264), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_12__6__SCAN_IN), .B2(n10594), .ZN(n10613) );
  AOI22_X1 U13613 ( .A1(n11265), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9887), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10612) );
  AOI22_X1 U13614 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n10648), .B1(
        n10536), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10611) );
  AOI22_X1 U13615 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10553), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10610) );
  NAND4_X1 U13616 ( .A1(n10613), .A2(n10612), .A3(n10611), .A4(n10610), .ZN(
        n10614) );
  NAND2_X1 U13617 ( .A1(n10768), .A2(n13598), .ZN(n10616) );
  INV_X1 U13618 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19865) );
  NAND2_X1 U13619 ( .A1(n13954), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10618) );
  NAND2_X1 U13620 ( .A1(n13955), .A2(P2_EAX_REG_6__SCAN_IN), .ZN(n10617) );
  OAI211_X1 U13621 ( .C1(n13958), .C2(n19865), .A(n10618), .B(n10617), .ZN(
        n13616) );
  NAND2_X1 U13622 ( .A1(n13617), .A2(n13616), .ZN(n10639) );
  NAND2_X1 U13623 ( .A1(n11264), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10622) );
  NAND2_X1 U13624 ( .A1(n11265), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10621) );
  NAND2_X1 U13625 ( .A1(n10594), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10620) );
  NAND2_X1 U13626 ( .A1(n9887), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10619) );
  NAND2_X1 U13627 ( .A1(n10603), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10626) );
  NAND2_X1 U13628 ( .A1(n11166), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10625) );
  NAND2_X1 U13629 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10624) );
  NAND2_X1 U13630 ( .A1(n10536), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10623) );
  AOI22_X1 U13631 ( .A1(n11255), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n10558), .ZN(n10629) );
  NAND2_X1 U13632 ( .A1(n11256), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10628) );
  NAND2_X1 U13633 ( .A1(n11257), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10627) );
  NAND2_X1 U13634 ( .A1(n11253), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10633) );
  NAND2_X1 U13635 ( .A1(n10553), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10632) );
  NAND2_X1 U13636 ( .A1(n11254), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10631) );
  NAND2_X1 U13637 ( .A1(n10537), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10630) );
  NAND2_X1 U13638 ( .A1(n10768), .A2(n13927), .ZN(n10638) );
  NAND2_X1 U13639 ( .A1(n10639), .A2(n10638), .ZN(n15514) );
  INV_X1 U13640 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19867) );
  NAND2_X1 U13641 ( .A1(n13954), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10641) );
  NAND2_X1 U13642 ( .A1(n13955), .A2(P2_EAX_REG_7__SCAN_IN), .ZN(n10640) );
  OAI211_X1 U13643 ( .C1(n13958), .C2(n19867), .A(n10641), .B(n10640), .ZN(
        n15513) );
  AOI22_X1 U13644 ( .A1(n13954), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n13955), .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n10657) );
  NAND2_X1 U13645 ( .A1(n10795), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n10656) );
  AOI22_X1 U13646 ( .A1(n11166), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11254), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10647) );
  AOI22_X1 U13647 ( .A1(n10603), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11253), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10646) );
  AOI22_X1 U13648 ( .A1(n11255), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10558), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10644) );
  NAND2_X1 U13649 ( .A1(n9887), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10643) );
  NAND2_X1 U13650 ( .A1(n11257), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10642) );
  AND3_X1 U13651 ( .A1(n10644), .A2(n10643), .A3(n10642), .ZN(n10645) );
  NAND3_X1 U13652 ( .A1(n10647), .A2(n10646), .A3(n10645), .ZN(n10654) );
  AOI22_X1 U13653 ( .A1(n11264), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10652) );
  AOI22_X1 U13654 ( .A1(n11265), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11256), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10651) );
  AOI22_X1 U13655 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10536), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10650) );
  AOI22_X1 U13656 ( .A1(n10553), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10649) );
  NAND4_X1 U13657 ( .A1(n10652), .A2(n10651), .A3(n10650), .A4(n10649), .ZN(
        n10653) );
  NAND2_X1 U13658 ( .A1(n10768), .A2(n13040), .ZN(n10655) );
  AOI22_X1 U13659 ( .A1(n10795), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n13954), .ZN(n10671) );
  AOI22_X1 U13660 ( .A1(n11166), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n11253), .ZN(n10663) );
  AOI22_X1 U13661 ( .A1(n10603), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n11254), .ZN(n10662) );
  AOI22_X1 U13662 ( .A1(n11255), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n10558), .ZN(n10660) );
  NAND2_X1 U13663 ( .A1(n11256), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10659) );
  NAND2_X1 U13664 ( .A1(n11257), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10658) );
  AND3_X1 U13665 ( .A1(n10660), .A2(n10659), .A3(n10658), .ZN(n10661) );
  NAND3_X1 U13666 ( .A1(n10663), .A2(n10662), .A3(n10661), .ZN(n10669) );
  AOI22_X1 U13667 ( .A1(n11264), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10667) );
  AOI22_X1 U13668 ( .A1(n11265), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9887), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10666) );
  AOI22_X1 U13669 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n10536), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10665) );
  AOI22_X1 U13670 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10553), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10664) );
  NAND4_X1 U13671 ( .A1(n10667), .A2(n10666), .A3(n10665), .A4(n10664), .ZN(
        n10668) );
  AOI22_X1 U13672 ( .A1(n10768), .A2(n13043), .B1(P2_EAX_REG_9__SCAN_IN), .B2(
        n13955), .ZN(n10670) );
  NAND2_X1 U13673 ( .A1(n10671), .A2(n10670), .ZN(n14793) );
  AOI22_X1 U13674 ( .A1(n13954), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n10507), .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n10686) );
  NAND2_X1 U13675 ( .A1(n10795), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n10685) );
  AOI22_X1 U13676 ( .A1(n11166), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10677) );
  AOI22_X1 U13677 ( .A1(n10603), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11253), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10676) );
  AOI22_X1 U13678 ( .A1(n11255), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10558), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10674) );
  NAND2_X1 U13679 ( .A1(n11256), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10673) );
  NAND2_X1 U13680 ( .A1(n11257), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n10672) );
  AND3_X1 U13681 ( .A1(n10674), .A2(n10673), .A3(n10672), .ZN(n10675) );
  NAND3_X1 U13682 ( .A1(n10677), .A2(n10676), .A3(n10675), .ZN(n10683) );
  AOI22_X1 U13683 ( .A1(n11264), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10681) );
  AOI22_X1 U13684 ( .A1(n11265), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9887), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10680) );
  AOI22_X1 U13685 ( .A1(n11254), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10679) );
  AOI22_X1 U13686 ( .A1(n10553), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10536), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10678) );
  NAND4_X1 U13687 ( .A1(n10681), .A2(n10680), .A3(n10679), .A4(n10678), .ZN(
        n10682) );
  NAND2_X1 U13688 ( .A1(n10768), .A2(n13140), .ZN(n10684) );
  AOI22_X1 U13689 ( .A1(n11264), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10690) );
  AOI22_X1 U13690 ( .A1(n11265), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9887), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10689) );
  AOI22_X1 U13691 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10536), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10688) );
  AOI22_X1 U13692 ( .A1(n10553), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10687) );
  NAND4_X1 U13693 ( .A1(n10690), .A2(n10689), .A3(n10688), .A4(n10687), .ZN(
        n10700) );
  AOI22_X1 U13694 ( .A1(n11166), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11253), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10698) );
  AOI22_X1 U13695 ( .A1(n10603), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11254), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10697) );
  INV_X1 U13696 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10691) );
  NOR2_X1 U13697 ( .A1(n10756), .A2(n10691), .ZN(n10694) );
  INV_X1 U13698 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10692) );
  INV_X1 U13699 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11322) );
  OAI22_X1 U13700 ( .A1(n10752), .A2(n10692), .B1(n10723), .B2(n11322), .ZN(
        n10693) );
  NOR2_X1 U13701 ( .A1(n10694), .A2(n10693), .ZN(n10696) );
  NAND2_X1 U13702 ( .A1(n11256), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n10695) );
  NAND4_X1 U13703 ( .A1(n10698), .A2(n10697), .A3(n10696), .A4(n10695), .ZN(
        n10699) );
  AOI22_X1 U13704 ( .A1(n10795), .A2(P2_REIP_REG_11__SCAN_IN), .B1(n10768), 
        .B2(n13281), .ZN(n10702) );
  AOI22_X1 U13705 ( .A1(n13954), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(
        n10507), .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n10701) );
  NAND2_X1 U13706 ( .A1(n10702), .A2(n10701), .ZN(n15469) );
  NAND2_X1 U13707 ( .A1(n15470), .A2(n15469), .ZN(n15450) );
  AOI22_X1 U13708 ( .A1(n13954), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n10507), .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n10717) );
  NAND2_X1 U13709 ( .A1(n10795), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n10716) );
  AOI22_X1 U13710 ( .A1(n11166), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10708) );
  AOI22_X1 U13711 ( .A1(n11255), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10558), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10705) );
  NAND2_X1 U13712 ( .A1(n11256), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10704) );
  NAND2_X1 U13713 ( .A1(n11257), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10703) );
  AND3_X1 U13714 ( .A1(n10705), .A2(n10704), .A3(n10703), .ZN(n10707) );
  AOI22_X1 U13715 ( .A1(n11253), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10706) );
  NAND3_X1 U13716 ( .A1(n10708), .A2(n10707), .A3(n10706), .ZN(n10714) );
  AOI22_X1 U13717 ( .A1(n11264), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10712) );
  AOI22_X1 U13718 ( .A1(n11265), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9887), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10711) );
  AOI22_X1 U13719 ( .A1(n10603), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11254), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10710) );
  AOI22_X1 U13720 ( .A1(n10553), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10536), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10709) );
  NAND4_X1 U13721 ( .A1(n10712), .A2(n10711), .A3(n10710), .A4(n10709), .ZN(
        n10713) );
  NAND2_X1 U13722 ( .A1(n10768), .A2(n13280), .ZN(n10715) );
  AOI22_X1 U13723 ( .A1(n10795), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n13954), .ZN(n10733) );
  AOI22_X1 U13724 ( .A1(n11264), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10721) );
  AOI22_X1 U13725 ( .A1(n11265), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9887), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10720) );
  AOI22_X1 U13726 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10536), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10719) );
  AOI22_X1 U13727 ( .A1(n10553), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10718) );
  NAND4_X1 U13728 ( .A1(n10721), .A2(n10720), .A3(n10719), .A4(n10718), .ZN(
        n10731) );
  AOI22_X1 U13729 ( .A1(n11166), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11253), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10729) );
  AOI22_X1 U13730 ( .A1(n10603), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11254), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10728) );
  INV_X1 U13731 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10722) );
  NOR2_X1 U13732 ( .A1(n10756), .A2(n10722), .ZN(n10725) );
  INV_X1 U13733 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11210) );
  INV_X1 U13734 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11366) );
  OAI22_X1 U13735 ( .A1(n10752), .A2(n11210), .B1(n10723), .B2(n11366), .ZN(
        n10724) );
  NOR2_X1 U13736 ( .A1(n10725), .A2(n10724), .ZN(n10727) );
  NAND2_X1 U13737 ( .A1(n11256), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10726) );
  NAND4_X1 U13738 ( .A1(n10729), .A2(n10728), .A3(n10727), .A4(n10726), .ZN(
        n10730) );
  AOI22_X1 U13739 ( .A1(n10768), .A2(n13294), .B1(P2_EAX_REG_13__SCAN_IN), 
        .B2(n13955), .ZN(n10732) );
  NAND2_X1 U13740 ( .A1(n10733), .A2(n10732), .ZN(n15439) );
  AOI22_X1 U13741 ( .A1(n11255), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n10558), .ZN(n10736) );
  NAND2_X1 U13742 ( .A1(n9887), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n10735) );
  NAND2_X1 U13743 ( .A1(n11257), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n10734) );
  AND3_X1 U13744 ( .A1(n10736), .A2(n10735), .A3(n10734), .ZN(n10740) );
  AOI22_X1 U13745 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n11253), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10739) );
  NAND2_X1 U13746 ( .A1(n10603), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n10738) );
  NAND2_X1 U13747 ( .A1(n11166), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n10737) );
  NAND4_X1 U13748 ( .A1(n10740), .A2(n10739), .A3(n10738), .A4(n10737), .ZN(
        n10746) );
  AOI22_X1 U13749 ( .A1(n11264), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10744) );
  AOI22_X1 U13750 ( .A1(n11265), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11256), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10743) );
  AOI22_X1 U13751 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n11254), .B1(
        n10536), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10742) );
  AOI22_X1 U13752 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10553), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10741) );
  NAND4_X1 U13753 ( .A1(n10744), .A2(n10743), .A3(n10742), .A4(n10741), .ZN(
        n10745) );
  INV_X1 U13754 ( .A(n13296), .ZN(n10749) );
  AOI22_X1 U13755 ( .A1(n13954), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n10507), .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n10747) );
  OAI21_X1 U13756 ( .B1(n10749), .B2(n10748), .A(n10747), .ZN(n10750) );
  AOI21_X1 U13757 ( .B1(P2_REIP_REG_14__SCAN_IN), .B2(n10795), .A(n10750), 
        .ZN(n15422) );
  AOI22_X1 U13758 ( .A1(n11166), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n11253), .ZN(n10761) );
  AOI22_X1 U13759 ( .A1(n10603), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n11254), .ZN(n10760) );
  INV_X1 U13760 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10755) );
  INV_X1 U13761 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10751) );
  OR2_X1 U13762 ( .A1(n10752), .A2(n10751), .ZN(n10754) );
  NAND2_X1 U13763 ( .A1(n10558), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10753) );
  OAI211_X1 U13764 ( .C1(n10756), .C2(n10755), .A(n10754), .B(n10753), .ZN(
        n10757) );
  INV_X1 U13765 ( .A(n10757), .ZN(n10759) );
  NAND2_X1 U13766 ( .A1(n11256), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10758) );
  NAND4_X1 U13767 ( .A1(n10761), .A2(n10760), .A3(n10759), .A4(n10758), .ZN(
        n10767) );
  AOI22_X1 U13768 ( .A1(n11264), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10765) );
  AOI22_X1 U13769 ( .A1(n11265), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9887), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10764) );
  AOI22_X1 U13770 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n10648), .B1(
        n10536), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10763) );
  AOI22_X1 U13771 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10553), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10762) );
  NAND4_X1 U13772 ( .A1(n10765), .A2(n10764), .A3(n10763), .A4(n10762), .ZN(
        n10766) );
  AOI22_X1 U13773 ( .A1(n10795), .A2(P2_REIP_REG_15__SCAN_IN), .B1(n10768), 
        .B2(n11136), .ZN(n10770) );
  AOI22_X1 U13774 ( .A1(n13954), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(
        n10507), .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n10769) );
  NAND2_X1 U13775 ( .A1(n10770), .A2(n10769), .ZN(n15411) );
  AOI22_X1 U13776 ( .A1(n13954), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n10507), .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n10772) );
  NAND2_X1 U13777 ( .A1(n10795), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n10771) );
  INV_X1 U13778 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19887) );
  INV_X1 U13779 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13469) );
  INV_X1 U13780 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15383) );
  OAI222_X1 U13781 ( .A1(n13958), .A2(n19887), .B1(n10774), .B2(n13469), .C1(
        n15383), .C2(n10773), .ZN(n13468) );
  AOI222_X1 U13782 ( .A1(P2_REIP_REG_18__SCAN_IN), .A2(n10795), .B1(n13954), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .C1(n10507), .C2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n15361) );
  INV_X1 U13783 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19891) );
  NAND2_X1 U13784 ( .A1(n13954), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10776) );
  NAND2_X1 U13785 ( .A1(n13955), .A2(P2_EAX_REG_19__SCAN_IN), .ZN(n10775) );
  OAI211_X1 U13786 ( .C1(n13958), .C2(n19891), .A(n10776), .B(n10775), .ZN(
        n14985) );
  INV_X1 U13787 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19893) );
  NAND2_X1 U13788 ( .A1(n13954), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10778) );
  NAND2_X1 U13789 ( .A1(n13955), .A2(P2_EAX_REG_20__SCAN_IN), .ZN(n10777) );
  OAI211_X1 U13790 ( .C1(n13958), .C2(n19893), .A(n10778), .B(n10777), .ZN(
        n15340) );
  AOI22_X1 U13791 ( .A1(n13954), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(
        n10507), .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n10780) );
  NAND2_X1 U13792 ( .A1(n10795), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n10779) );
  AND2_X1 U13793 ( .A1(n10780), .A2(n10779), .ZN(n14786) );
  AOI22_X1 U13794 ( .A1(n13954), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B1(
        n13955), .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n10782) );
  NAND2_X1 U13795 ( .A1(n10795), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n10781) );
  INV_X1 U13796 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19899) );
  NAND2_X1 U13797 ( .A1(n13954), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10784) );
  NAND2_X1 U13798 ( .A1(n13955), .A2(P2_EAX_REG_23__SCAN_IN), .ZN(n10783) );
  OAI211_X1 U13799 ( .C1(n13958), .C2(n19899), .A(n10784), .B(n10783), .ZN(
        n12463) );
  AOI22_X1 U13800 ( .A1(n13954), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B1(
        n13955), .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n10786) );
  NAND2_X1 U13801 ( .A1(n10795), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n10785) );
  AND2_X1 U13802 ( .A1(n10786), .A2(n10785), .ZN(n12431) );
  AOI22_X1 U13803 ( .A1(n13954), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n13955), .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n10788) );
  NAND2_X1 U13804 ( .A1(n10795), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n10787) );
  AND2_X1 U13805 ( .A1(n10788), .A2(n10787), .ZN(n14950) );
  OR2_X2 U13806 ( .A1(n9874), .A2(n14950), .ZN(n14952) );
  AOI22_X1 U13807 ( .A1(n13954), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B1(
        n13955), .B2(P2_EAX_REG_26__SCAN_IN), .ZN(n10790) );
  NAND2_X1 U13808 ( .A1(n10795), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n10789) );
  AND2_X1 U13809 ( .A1(n10790), .A2(n10789), .ZN(n14943) );
  INV_X1 U13810 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19907) );
  NAND2_X1 U13811 ( .A1(n13954), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10792) );
  NAND2_X1 U13812 ( .A1(n13955), .A2(P2_EAX_REG_27__SCAN_IN), .ZN(n10791) );
  OAI211_X1 U13813 ( .C1(n13958), .C2(n19907), .A(n10792), .B(n10791), .ZN(
        n12445) );
  AOI22_X1 U13814 ( .A1(n13954), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        n13955), .B2(P2_EAX_REG_28__SCAN_IN), .ZN(n10794) );
  NAND2_X1 U13815 ( .A1(n10795), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n10793) );
  AND2_X1 U13816 ( .A1(n10794), .A2(n10793), .ZN(n14929) );
  AOI22_X1 U13817 ( .A1(n13954), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        n13955), .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n10797) );
  NAND2_X1 U13818 ( .A1(n10795), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n10796) );
  AND2_X1 U13819 ( .A1(n10797), .A2(n10796), .ZN(n14769) );
  INV_X1 U13820 ( .A(n10799), .ZN(n14771) );
  AOI21_X1 U13821 ( .B1(n10800), .B2(n14771), .A(n13960), .ZN(n15221) );
  AOI22_X1 U13822 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10843), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10804) );
  AOI22_X1 U13823 ( .A1(n9836), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(n9839), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10802) );
  AOI22_X1 U13824 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10845), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10801) );
  NAND4_X1 U13825 ( .A1(n10804), .A2(n10803), .A3(n10802), .A4(n10801), .ZN(
        n10805) );
  NAND2_X1 U13826 ( .A1(n10805), .A2(n10861), .ZN(n10812) );
  AOI22_X1 U13827 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10843), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10808) );
  AOI22_X1 U13828 ( .A1(n9836), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9839), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10807) );
  AOI22_X1 U13829 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10845), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10806) );
  NAND4_X1 U13830 ( .A1(n10809), .A2(n10808), .A3(n10807), .A4(n10806), .ZN(
        n10810) );
  NAND2_X1 U13831 ( .A1(n10810), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10811) );
  NAND2_X2 U13832 ( .A1(n10812), .A2(n10811), .ZN(n10902) );
  AOI22_X1 U13833 ( .A1(n11233), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9844), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10814) );
  AOI22_X1 U13834 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10843), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10816) );
  AOI22_X1 U13835 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10845), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10815) );
  AOI22_X1 U13836 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10843), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10820) );
  AOI22_X1 U13837 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9838), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10819) );
  AOI22_X1 U13838 ( .A1(n11233), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9843), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10818) );
  AOI22_X1 U13839 ( .A1(n9835), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9840), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10824) );
  AOI22_X1 U13840 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9838), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10823) );
  AOI22_X1 U13841 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10843), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10826) );
  AOI22_X1 U13842 ( .A1(n11233), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9844), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10825) );
  NAND2_X1 U13843 ( .A1(n10827), .A2(n10362), .ZN(n10835) );
  NAND2_X1 U13844 ( .A1(n9839), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10828) );
  AOI22_X1 U13845 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10843), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10832) );
  AOI22_X1 U13846 ( .A1(n11233), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9843), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10831) );
  AOI22_X1 U13847 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10845), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10830) );
  NAND4_X1 U13848 ( .A1(n10833), .A2(n10832), .A3(n10831), .A4(n10830), .ZN(
        n10834) );
  NAND2_X2 U13849 ( .A1(n10835), .A2(n10834), .ZN(n10905) );
  NAND2_X1 U13850 ( .A1(n10836), .A2(n11101), .ZN(n10837) );
  AOI22_X1 U13851 ( .A1(n9835), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(n9840), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10841) );
  AOI22_X1 U13852 ( .A1(n11233), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9844), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10840) );
  AOI22_X1 U13853 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10843), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10839) );
  AOI22_X1 U13854 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9838), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10838) );
  NAND4_X1 U13855 ( .A1(n10841), .A2(n10840), .A3(n10839), .A4(n10838), .ZN(
        n10842) );
  AOI22_X1 U13856 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10843), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10851) );
  AOI22_X1 U13857 ( .A1(n11233), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9844), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10850) );
  AOI22_X1 U13858 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10845), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10849) );
  AOI22_X1 U13859 ( .A1(n9840), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9835), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10848) );
  NAND4_X1 U13860 ( .A1(n10851), .A2(n10850), .A3(n10849), .A4(n10848), .ZN(
        n10852) );
  NAND2_X1 U13861 ( .A1(n10914), .A2(n10915), .ZN(n10874) );
  AND2_X2 U13862 ( .A1(n10874), .A2(n11452), .ZN(n10901) );
  NAND2_X1 U13863 ( .A1(n19964), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11435) );
  XNOR2_X1 U13864 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12485) );
  INV_X1 U13865 ( .A(n12485), .ZN(n11438) );
  XNOR2_X1 U13866 ( .A(n10857), .B(n11438), .ZN(n11436) );
  NAND2_X1 U13867 ( .A1(n10857), .A2(n12485), .ZN(n10859) );
  NAND2_X1 U13868 ( .A1(n19955), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10858) );
  NOR2_X1 U13869 ( .A1(n16329), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10860) );
  MUX2_X1 U13870 ( .A(n19935), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        n10861), .Z(n10864) );
  NAND3_X1 U13871 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n10870), .A3(
        n15663), .ZN(n11430) );
  XNOR2_X1 U13872 ( .A(n16329), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10862) );
  XNOR2_X1 U13873 ( .A(n10863), .B(n10862), .ZN(n11434) );
  AND2_X1 U13874 ( .A1(n10865), .A2(n10864), .ZN(n10866) );
  OR2_X1 U13875 ( .A1(n10867), .A2(n10866), .ZN(n10883) );
  NAND3_X1 U13876 ( .A1(n11430), .A2(n11434), .A3(n11429), .ZN(n12479) );
  INV_X1 U13877 ( .A(n12479), .ZN(n10868) );
  NAND2_X1 U13878 ( .A1(n11436), .A2(n10868), .ZN(n10871) );
  NOR2_X1 U13879 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16340), .ZN(
        n10869) );
  INV_X1 U13880 ( .A(n11449), .ZN(n12492) );
  NAND2_X1 U13881 ( .A1(n16348), .A2(n16362), .ZN(n12471) );
  INV_X1 U13882 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19837) );
  NAND2_X1 U13883 ( .A1(n19848), .A2(n19856), .ZN(n19836) );
  OAI211_X1 U13884 ( .C1(n19848), .C2(n19856), .A(n19837), .B(n19836), .ZN(
        n19841) );
  NAND2_X1 U13885 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19835) );
  INV_X1 U13886 ( .A(n19835), .ZN(n19851) );
  NOR2_X1 U13887 ( .A1(n19841), .A2(n19851), .ZN(n12649) );
  INV_X1 U13888 ( .A(n12649), .ZN(n12475) );
  NOR2_X1 U13889 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n12475), .ZN(n10875) );
  AND3_X1 U13890 ( .A1(n19247), .A2(n10875), .A3(n10915), .ZN(n16367) );
  NAND2_X1 U13891 ( .A1(n19923), .A2(n19832), .ZN(n18908) );
  AND3_X1 U13892 ( .A1(n19825), .A2(n19829), .A3(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n16361) );
  INV_X1 U13893 ( .A(n16361), .ZN(n10872) );
  NAND2_X1 U13894 ( .A1(n19831), .A2(n10872), .ZN(n10873) );
  NAND2_X1 U13895 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19089), .ZN(
        n10880) );
  NAND2_X1 U13896 ( .A1(n19924), .A2(n19835), .ZN(n11087) );
  INV_X1 U13897 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n14827) );
  AND2_X1 U13898 ( .A1(n11087), .A2(n14827), .ZN(n10877) );
  INV_X1 U13899 ( .A(n10875), .ZN(n10876) );
  OAI21_X1 U13900 ( .B1(n19247), .B2(n10877), .A(n10876), .ZN(n10878) );
  NAND2_X1 U13901 ( .A1(n19109), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10879) );
  OAI211_X1 U13902 ( .C1(n19122), .C2(n15003), .A(n10880), .B(n10879), .ZN(
        n10898) );
  MUX2_X1 U13903 ( .A(n11430), .B(n13315), .S(n12679), .Z(n12490) );
  INV_X1 U13904 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n12897) );
  MUX2_X1 U13905 ( .A(n12490), .B(n12897), .S(n19267), .Z(n13308) );
  MUX2_X1 U13906 ( .A(n10881), .B(n11434), .S(n10906), .Z(n12486) );
  INV_X1 U13907 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13537) );
  MUX2_X1 U13908 ( .A(n12486), .B(n13537), .S(n19267), .Z(n13247) );
  NOR2_X1 U13909 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n10882) );
  MUX2_X1 U13910 ( .A(n13226), .B(n10882), .S(n19267), .Z(n13246) );
  NAND2_X1 U13911 ( .A1(n13247), .A2(n13246), .ZN(n13249) );
  MUX2_X1 U13912 ( .A(n13207), .B(n10883), .S(n10906), .Z(n12488) );
  MUX2_X1 U13913 ( .A(n12488), .B(P2_EBX_REG_3__SCAN_IN), .S(n19267), .Z(
        n13238) );
  MUX2_X1 U13914 ( .A(n13376), .B(P2_EBX_REG_5__SCAN_IN), .S(n19267), .Z(
        n13380) );
  INV_X1 U13915 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n12950) );
  MUX2_X1 U13916 ( .A(n13598), .B(n12950), .S(n19267), .Z(n13613) );
  INV_X1 U13917 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n10997) );
  MUX2_X1 U13918 ( .A(n13927), .B(n10997), .S(n19267), .Z(n13817) );
  INV_X1 U13919 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n19041) );
  NAND2_X1 U13920 ( .A1(n19267), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13815) );
  INV_X1 U13921 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n19056) );
  NAND2_X1 U13922 ( .A1(n13906), .A2(n13841), .ZN(n13838) );
  NAND2_X1 U13923 ( .A1(n19267), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10885) );
  NAND2_X1 U13924 ( .A1(n19267), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n13875) );
  OAI21_X1 U13925 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(P2_EBX_REG_14__SCAN_IN), 
        .A(n19267), .ZN(n10886) );
  INV_X1 U13926 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n10888) );
  INV_X1 U13927 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n10887) );
  NAND2_X1 U13928 ( .A1(n10888), .A2(n10887), .ZN(n10889) );
  AND2_X1 U13929 ( .A1(n19267), .A2(n10889), .ZN(n10890) );
  NAND2_X1 U13930 ( .A1(n19267), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n13851) );
  INV_X1 U13931 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n10891) );
  NAND2_X1 U13932 ( .A1(n19267), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12415) );
  AND2_X1 U13933 ( .A1(n19267), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12455) );
  INV_X1 U13934 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n16222) );
  NAND2_X1 U13935 ( .A1(n13906), .A2(n9878), .ZN(n13909) );
  NAND2_X1 U13936 ( .A1(n19267), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10893) );
  AND2_X1 U13937 ( .A1(n19267), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n13918) );
  NAND2_X1 U13938 ( .A1(n19267), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n13922) );
  NAND2_X1 U13939 ( .A1(n13923), .A2(n13922), .ZN(n14760) );
  AND2_X1 U13940 ( .A1(n19267), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10894) );
  XNOR2_X1 U13941 ( .A(n14760), .B(n10894), .ZN(n13925) );
  NAND2_X1 U13942 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n11087), .ZN(n10895) );
  NOR2_X1 U13943 ( .A1(n10906), .A2(n10895), .ZN(n10896) );
  NAND2_X2 U13944 ( .A1(n18911), .A2(n10896), .ZN(n19106) );
  NOR2_X1 U13945 ( .A1(n13925), .A2(n19106), .ZN(n10897) );
  AOI211_X1 U13946 ( .C1(n15221), .C2(n19036), .A(n10898), .B(n10897), .ZN(
        n11092) );
  AND2_X1 U13947 ( .A1(n10911), .A2(n10899), .ZN(n11459) );
  NAND3_X1 U13948 ( .A1(n11469), .A2(n11459), .A3(n10930), .ZN(n10900) );
  NAND2_X1 U13949 ( .A1(n10938), .A2(n19247), .ZN(n10910) );
  NAND3_X1 U13950 ( .A1(n12673), .A2(n10911), .A3(n19247), .ZN(n10904) );
  NAND2_X1 U13951 ( .A1(n10904), .A2(n10903), .ZN(n10908) );
  NAND2_X1 U13952 ( .A1(n12644), .A2(n10930), .ZN(n11455) );
  NOR2_X1 U13953 ( .A1(n11455), .A2(n10899), .ZN(n10907) );
  INV_X1 U13954 ( .A(n10909), .ZN(n12400) );
  NAND2_X2 U13955 ( .A1(n10910), .A2(n10943), .ZN(n12661) );
  BUF_X2 U13956 ( .A(n10914), .Z(n12648) );
  AND2_X4 U13957 ( .A1(n12648), .A2(n10916), .ZN(n13947) );
  AOI22_X1 U13958 ( .A1(n13947), .A2(P2_REIP_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10917) );
  OAI21_X1 U13959 ( .B1(n10967), .B2(n12627), .A(n10917), .ZN(n10918) );
  NAND2_X1 U13960 ( .A1(n10949), .A2(n16347), .ZN(n10927) );
  INV_X1 U13961 ( .A(n10912), .ZN(n10924) );
  NAND2_X1 U13962 ( .A1(n10924), .A2(n11455), .ZN(n10923) );
  NAND2_X1 U13963 ( .A1(n11461), .A2(n10902), .ZN(n10922) );
  AOI21_X1 U13964 ( .B1(n9818), .B2(n10899), .A(n12652), .ZN(n10921) );
  NAND3_X1 U13965 ( .A1(n10923), .A2(n10922), .A3(n10921), .ZN(n10926) );
  INV_X1 U13966 ( .A(n12648), .ZN(n10936) );
  INV_X1 U13967 ( .A(n10933), .ZN(n10934) );
  NAND3_X1 U13968 ( .A1(n16346), .A2(n19252), .A3(n13216), .ZN(n10935) );
  NAND2_X1 U13969 ( .A1(n10936), .A2(n10935), .ZN(n10937) );
  NOR2_X1 U13970 ( .A1(n16363), .A2(n19955), .ZN(n10939) );
  AND3_X1 U13971 ( .A1(n10909), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n12679), 
        .ZN(n10942) );
  INV_X4 U13972 ( .A(n10967), .ZN(n11032) );
  INV_X1 U13973 ( .A(n10943), .ZN(n10945) );
  NOR2_X1 U13974 ( .A1(n16363), .A2(n19964), .ZN(n10944) );
  AOI21_X1 U13975 ( .B1(n10945), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10944), 
        .ZN(n10946) );
  NAND2_X1 U13976 ( .A1(n10947), .A2(n10946), .ZN(n11116) );
  AOI21_X1 U13977 ( .B1(n10948), .B2(n10949), .A(n10951), .ZN(n10959) );
  NAND2_X1 U13978 ( .A1(n10952), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10958) );
  NAND2_X1 U13979 ( .A1(n13947), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10954) );
  NAND2_X1 U13980 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10953) );
  NAND3_X1 U13981 ( .A1(n10955), .A2(n10954), .A3(n10372), .ZN(n10956) );
  OAI211_X1 U13982 ( .C1(n10959), .C2(n18909), .A(n10958), .B(n10957), .ZN(
        n11117) );
  NAND2_X1 U13983 ( .A1(n11116), .A2(n11117), .ZN(n11115) );
  NAND2_X1 U13984 ( .A1(n11121), .A2(n11115), .ZN(n10964) );
  INV_X1 U13985 ( .A(n10961), .ZN(n10962) );
  NAND2_X1 U13986 ( .A1(n10964), .A2(n10963), .ZN(n10972) );
  OAI21_X1 U13987 ( .B1(n19946), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n19832), 
        .ZN(n10966) );
  NAND2_X1 U13988 ( .A1(n10972), .A2(n10973), .ZN(n11106) );
  AOI22_X1 U13989 ( .A1(n13947), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10968) );
  OAI21_X1 U13990 ( .B1(n13950), .B2(n13537), .A(n10968), .ZN(n10969) );
  INV_X1 U13991 ( .A(n10969), .ZN(n10970) );
  NAND2_X1 U13992 ( .A1(n11106), .A2(n11107), .ZN(n10975) );
  INV_X1 U13993 ( .A(n10973), .ZN(n10974) );
  NAND2_X1 U13994 ( .A1(n9823), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10977) );
  OR2_X1 U13995 ( .A1(n16363), .A2(n19935), .ZN(n10976) );
  INV_X1 U13996 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13619) );
  INV_X1 U13997 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n10979) );
  AOI22_X1 U13998 ( .A1(n13947), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10978) );
  OAI21_X1 U13999 ( .B1(n13950), .B2(n10979), .A(n10978), .ZN(n10980) );
  INV_X1 U14000 ( .A(n10980), .ZN(n10981) );
  XNOR2_X2 U14001 ( .A(n10984), .B(n10983), .ZN(n11095) );
  AOI22_X1 U14002 ( .A1(n13947), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10985) );
  OAI21_X1 U14003 ( .B1(n13950), .B2(n12897), .A(n10985), .ZN(n10986) );
  AOI21_X1 U14004 ( .B1(n11086), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n10986), .ZN(n12895) );
  INV_X1 U14005 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13618) );
  OR2_X1 U14006 ( .A1(n11078), .A2(n13618), .ZN(n10991) );
  INV_X1 U14007 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n10988) );
  AOI22_X1 U14008 ( .A1(n13947), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10987) );
  OAI21_X1 U14009 ( .B1(n13950), .B2(n10988), .A(n10987), .ZN(n10989) );
  INV_X1 U14010 ( .A(n10989), .ZN(n10990) );
  NAND2_X1 U14011 ( .A1(n10991), .A2(n10990), .ZN(n12913) );
  NAND2_X1 U14012 ( .A1(n12912), .A2(n12913), .ZN(n12944) );
  INV_X1 U14013 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13974) );
  OR2_X1 U14014 ( .A1(n11078), .A2(n13974), .ZN(n10995) );
  AOI22_X1 U14015 ( .A1(n13947), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10992) );
  OAI21_X1 U14016 ( .B1(n13950), .B2(n12950), .A(n10992), .ZN(n10993) );
  INV_X1 U14017 ( .A(n10993), .ZN(n10994) );
  INV_X1 U14018 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15511) );
  OR2_X1 U14019 ( .A1(n11078), .A2(n15511), .ZN(n11000) );
  AOI22_X1 U14020 ( .A1(n13947), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10996) );
  OAI21_X1 U14021 ( .B1(n13950), .B2(n10997), .A(n10996), .ZN(n10998) );
  INV_X1 U14022 ( .A(n10998), .ZN(n10999) );
  NAND2_X1 U14023 ( .A1(n11000), .A2(n10999), .ZN(n12918) );
  INV_X1 U14024 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11001) );
  OR2_X1 U14025 ( .A1(n11078), .A2(n11001), .ZN(n11006) );
  INV_X1 U14026 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n11003) );
  AOI22_X1 U14027 ( .A1(n13947), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11002) );
  OAI21_X1 U14028 ( .B1(n13950), .B2(n11003), .A(n11002), .ZN(n11004) );
  INV_X1 U14029 ( .A(n11004), .ZN(n11005) );
  INV_X1 U14030 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n13826) );
  OR2_X1 U14031 ( .A1(n11078), .A2(n13826), .ZN(n11011) );
  INV_X1 U14032 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n11008) );
  AOI22_X1 U14033 ( .A1(n13947), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11007) );
  OAI21_X1 U14034 ( .B1(n13950), .B2(n11008), .A(n11007), .ZN(n11009) );
  INV_X1 U14035 ( .A(n11009), .ZN(n11010) );
  NAND2_X1 U14036 ( .A1(n11011), .A2(n11010), .ZN(n13044) );
  INV_X1 U14037 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15488) );
  OR2_X1 U14038 ( .A1(n11078), .A2(n15488), .ZN(n11015) );
  AOI22_X1 U14039 ( .A1(n13947), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11012) );
  OAI21_X1 U14040 ( .B1(n13950), .B2(n19056), .A(n11012), .ZN(n11013) );
  INV_X1 U14041 ( .A(n11013), .ZN(n11014) );
  NAND2_X1 U14042 ( .A1(n11015), .A2(n11014), .ZN(n13142) );
  AOI22_X1 U14043 ( .A1(n13947), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11016) );
  OAI21_X1 U14044 ( .B1(n13950), .B2(n19041), .A(n11016), .ZN(n11017) );
  AOI21_X1 U14045 ( .B1(n11086), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n11017), .ZN(n13130) );
  INV_X1 U14046 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n11019) );
  AOI22_X1 U14047 ( .A1(n13947), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11018) );
  OAI21_X1 U14048 ( .B1(n13950), .B2(n11019), .A(n11018), .ZN(n11020) );
  AOI21_X1 U14049 ( .B1(n11086), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n11020), .ZN(n13283) );
  INV_X1 U14050 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15437) );
  OR2_X1 U14051 ( .A1(n11078), .A2(n15437), .ZN(n11025) );
  INV_X1 U14052 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n11022) );
  AOI22_X1 U14053 ( .A1(n13947), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n11021) );
  OAI21_X1 U14054 ( .B1(n13950), .B2(n11022), .A(n11021), .ZN(n11023) );
  INV_X1 U14055 ( .A(n11023), .ZN(n11024) );
  NAND2_X1 U14056 ( .A1(n11025), .A2(n11024), .ZN(n13174) );
  NAND2_X1 U14057 ( .A1(n13286), .A2(n13174), .ZN(n13298) );
  INV_X1 U14058 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n13866) );
  AOI22_X1 U14059 ( .A1(n13947), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11026) );
  OAI21_X1 U14060 ( .B1(n13950), .B2(n13866), .A(n11026), .ZN(n11027) );
  AOI21_X1 U14061 ( .B1(n11086), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n11027), .ZN(n13299) );
  INV_X1 U14062 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n11029) );
  AOI22_X1 U14063 ( .A1(n13947), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11028) );
  OAI21_X1 U14064 ( .B1(n13950), .B2(n11029), .A(n11028), .ZN(n11030) );
  AOI21_X1 U14065 ( .B1(n11086), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n11030), .ZN(n13418) );
  INV_X1 U14066 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15403) );
  OR2_X1 U14067 ( .A1(n11078), .A2(n15403), .ZN(n11035) );
  INV_X1 U14068 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19885) );
  OAI22_X1 U14069 ( .A1(n11079), .A2(n19885), .B1(n19832), .B2(n10142), .ZN(
        n11033) );
  AOI21_X1 U14070 ( .B1(n11032), .B2(P2_EBX_REG_16__SCAN_IN), .A(n11033), .ZN(
        n11034) );
  OR2_X1 U14071 ( .A1(n11078), .A2(n15383), .ZN(n11038) );
  OAI22_X1 U14072 ( .A1(n11079), .A2(n19887), .B1(n19832), .B2(n18982), .ZN(
        n11036) );
  AOI21_X1 U14073 ( .B1(n11032), .B2(P2_EBX_REG_17__SCAN_IN), .A(n11036), .ZN(
        n11037) );
  NAND2_X1 U14074 ( .A1(n11038), .A2(n11037), .ZN(n14907) );
  INV_X1 U14075 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15366) );
  OR2_X1 U14076 ( .A1(n11078), .A2(n15366), .ZN(n11043) );
  INV_X1 U14077 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n11040) );
  AOI22_X1 U14078 ( .A1(n13947), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11039) );
  OAI21_X1 U14079 ( .B1(n13950), .B2(n11040), .A(n11039), .ZN(n11041) );
  INV_X1 U14080 ( .A(n11041), .ZN(n11042) );
  NAND2_X1 U14081 ( .A1(n11043), .A2(n11042), .ZN(n14903) );
  INV_X1 U14082 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15337) );
  OR2_X1 U14083 ( .A1(n11078), .A2(n15337), .ZN(n11046) );
  OAI22_X1 U14084 ( .A1(n11079), .A2(n19891), .B1(n19832), .B2(n18959), .ZN(
        n11044) );
  AOI21_X1 U14085 ( .B1(n11032), .B2(P2_EBX_REG_19__SCAN_IN), .A(n11044), .ZN(
        n11045) );
  INV_X1 U14086 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15338) );
  OR2_X1 U14087 ( .A1(n11078), .A2(n15338), .ZN(n11050) );
  INV_X1 U14088 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11047) );
  OAI22_X1 U14089 ( .A1(n11079), .A2(n19893), .B1(n19832), .B2(n11047), .ZN(
        n11048) );
  AOI21_X1 U14090 ( .B1(n11032), .B2(P2_EBX_REG_20__SCAN_IN), .A(n11048), .ZN(
        n11049) );
  INV_X1 U14091 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15109) );
  OR2_X1 U14092 ( .A1(n11078), .A2(n15109), .ZN(n11053) );
  INV_X1 U14093 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19895) );
  OAI22_X1 U14094 ( .A1(n11079), .A2(n19895), .B1(n19832), .B2(n15110), .ZN(
        n11051) );
  AOI21_X1 U14095 ( .B1(n11032), .B2(P2_EBX_REG_21__SCAN_IN), .A(n11051), .ZN(
        n11052) );
  NAND2_X1 U14096 ( .A1(n11053), .A2(n11052), .ZN(n14783) );
  INV_X1 U14097 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n13899) );
  OR2_X1 U14098 ( .A1(n11078), .A2(n13899), .ZN(n11057) );
  INV_X1 U14099 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19897) );
  OAI22_X1 U14100 ( .A1(n11079), .A2(n19897), .B1(n19832), .B2(n11054), .ZN(
        n11055) );
  AOI21_X1 U14101 ( .B1(n11032), .B2(P2_EBX_REG_22__SCAN_IN), .A(n11055), .ZN(
        n11056) );
  NAND2_X1 U14102 ( .A1(n11057), .A2(n11056), .ZN(n12419) );
  INV_X1 U14103 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11058) );
  OR2_X1 U14104 ( .A1(n11078), .A2(n11058), .ZN(n11061) );
  OAI22_X1 U14105 ( .A1(n11079), .A2(n19899), .B1(n19832), .B2(n10164), .ZN(
        n11059) );
  AOI21_X1 U14106 ( .B1(n11032), .B2(P2_EBX_REG_23__SCAN_IN), .A(n11059), .ZN(
        n11060) );
  AND2_X1 U14107 ( .A1(n11061), .A2(n11060), .ZN(n12462) );
  INV_X1 U14108 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15289) );
  OR2_X1 U14109 ( .A1(n11078), .A2(n15289), .ZN(n11064) );
  INV_X1 U14110 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19901) );
  OAI22_X1 U14111 ( .A1(n11079), .A2(n19901), .B1(n19832), .B2(n15070), .ZN(
        n11062) );
  AOI21_X1 U14112 ( .B1(n11032), .B2(P2_EBX_REG_24__SCAN_IN), .A(n11062), .ZN(
        n11063) );
  AND2_X1 U14113 ( .A1(n11064), .A2(n11063), .ZN(n12429) );
  AOI22_X1 U14114 ( .A1(n13947), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n11065) );
  OAI21_X1 U14115 ( .B1(n13950), .B2(n16222), .A(n11065), .ZN(n11066) );
  AOI21_X1 U14116 ( .B1(n11086), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n11066), .ZN(n14859) );
  INV_X1 U14117 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15272) );
  OR2_X1 U14118 ( .A1(n11078), .A2(n15272), .ZN(n11069) );
  INV_X1 U14119 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n15049) );
  OAI22_X1 U14120 ( .A1(n11079), .A2(n15049), .B1(n19832), .B2(n16206), .ZN(
        n11067) );
  AOI21_X1 U14121 ( .B1(n11032), .B2(P2_EBX_REG_26__SCAN_IN), .A(n11067), .ZN(
        n11068) );
  NAND2_X1 U14122 ( .A1(n11069), .A2(n11068), .ZN(n14847) );
  INV_X1 U14123 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15255) );
  OR2_X1 U14124 ( .A1(n11078), .A2(n15255), .ZN(n11072) );
  OAI22_X1 U14125 ( .A1(n11079), .A2(n19907), .B1(n19832), .B2(n15039), .ZN(
        n11070) );
  AOI21_X1 U14126 ( .B1(n11032), .B2(P2_EBX_REG_27__SCAN_IN), .A(n11070), .ZN(
        n11071) );
  NAND2_X1 U14127 ( .A1(n11072), .A2(n11071), .ZN(n12443) );
  OR2_X1 U14128 ( .A1(n11078), .A2(n10010), .ZN(n11077) );
  INV_X1 U14129 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n11074) );
  AOI22_X1 U14130 ( .A1(n13947), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n11073) );
  OAI21_X1 U14131 ( .B1(n13950), .B2(n11074), .A(n11073), .ZN(n11075) );
  INV_X1 U14132 ( .A(n11075), .ZN(n11076) );
  NAND2_X1 U14133 ( .A1(n11077), .A2(n11076), .ZN(n14837) );
  INV_X1 U14134 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15234) );
  OR2_X1 U14135 ( .A1(n11078), .A2(n15234), .ZN(n11082) );
  INV_X1 U14136 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19909) );
  INV_X1 U14137 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15015) );
  OAI22_X1 U14138 ( .A1(n11079), .A2(n19909), .B1(n19832), .B2(n15015), .ZN(
        n11080) );
  AOI21_X1 U14139 ( .B1(n11032), .B2(P2_EBX_REG_29__SCAN_IN), .A(n11080), .ZN(
        n11081) );
  AND2_X1 U14140 ( .A1(n11082), .A2(n11081), .ZN(n14766) );
  INV_X1 U14141 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n11084) );
  AOI22_X1 U14142 ( .A1(n13947), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11083) );
  OAI21_X1 U14143 ( .B1(n13950), .B2(n11084), .A(n11083), .ZN(n11085) );
  AOI21_X1 U14144 ( .B1(n11086), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n11085), .ZN(n13951) );
  INV_X1 U14145 ( .A(n15223), .ZN(n11090) );
  NOR2_X1 U14146 ( .A1(n10906), .A2(n11087), .ZN(n11088) );
  NAND2_X1 U14147 ( .A1(n18911), .A2(n11088), .ZN(n19115) );
  NAND2_X1 U14148 ( .A1(n11094), .A2(n11093), .ZN(P2_U2825) );
  XNOR2_X2 U14149 ( .A(n11096), .B(n11095), .ZN(n13192) );
  NAND2_X1 U14150 ( .A1(n13192), .A2(n12597), .ZN(n11100) );
  NAND2_X1 U14151 ( .A1(n10899), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11097) );
  NOR2_X1 U14152 ( .A1(n19946), .A2(n19955), .ZN(n19691) );
  OAI21_X1 U14153 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n11109), .A(
        n19923), .ZN(n11098) );
  NOR2_X1 U14154 ( .A1(n11098), .A2(n19760), .ZN(n19623) );
  AOI21_X1 U14155 ( .B1(n11124), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19623), .ZN(n11099) );
  NAND2_X1 U14156 ( .A1(n11100), .A2(n11099), .ZN(n11104) );
  NOR2_X1 U14157 ( .A1(n11337), .A2(n10692), .ZN(n11103) );
  NAND2_X1 U14158 ( .A1(n11104), .A2(n11103), .ZN(n12892) );
  OR2_X1 U14159 ( .A1(n11104), .A2(n11103), .ZN(n11105) );
  XNOR2_X2 U14160 ( .A(n11108), .B(n11107), .ZN(n13185) );
  INV_X1 U14161 ( .A(n11109), .ZN(n11111) );
  NAND2_X1 U14162 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19592) );
  NAND2_X1 U14163 ( .A1(n19592), .A2(n19946), .ZN(n11110) );
  NAND2_X1 U14164 ( .A1(n11111), .A2(n11110), .ZN(n19378) );
  NOR2_X1 U14165 ( .A1(n19931), .A2(n19378), .ZN(n11112) );
  AOI21_X1 U14166 ( .B1(n11124), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11112), .ZN(n11113) );
  INV_X1 U14167 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11168) );
  NOR2_X1 U14168 ( .A1(n11337), .A2(n11168), .ZN(n11114) );
  OR2_X1 U14169 ( .A1(n11117), .A2(n11116), .ZN(n11118) );
  AOI22_X1 U14170 ( .A1(n11124), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19923), .B2(n19964), .ZN(n11119) );
  NAND2_X1 U14171 ( .A1(n11360), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11128) );
  XNOR2_X1 U14172 ( .A(n11127), .B(n11128), .ZN(n12624) );
  INV_X1 U14173 ( .A(n11115), .ZN(n11123) );
  XNOR2_X2 U14174 ( .A(n13187), .B(n11123), .ZN(n13191) );
  NAND2_X1 U14175 ( .A1(n11124), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11125) );
  NAND2_X1 U14176 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19964), .ZN(
        n19563) );
  NAND2_X1 U14177 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19955), .ZN(
        n19525) );
  NAND2_X1 U14178 ( .A1(n19563), .A2(n19525), .ZN(n19377) );
  NAND2_X1 U14179 ( .A1(n19923), .A2(n19377), .ZN(n19568) );
  NAND2_X1 U14180 ( .A1(n11125), .A2(n19568), .ZN(n11126) );
  NAND2_X1 U14181 ( .A1(n12624), .A2(n12623), .ZN(n12626) );
  NAND2_X1 U14182 ( .A1(n15527), .A2(n11128), .ZN(n11129) );
  NAND2_X1 U14183 ( .A1(n12690), .A2(n12692), .ZN(n12691) );
  NAND2_X1 U14184 ( .A1(n12691), .A2(n11130), .ZN(n12748) );
  NAND2_X1 U14185 ( .A1(n12749), .A2(n12748), .ZN(n12750) );
  NAND2_X1 U14186 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n10899), .ZN(
        n11131) );
  AND2_X1 U14187 ( .A1(n11104), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11132) );
  NOR2_X1 U14188 ( .A1(n11337), .A2(n10574), .ZN(n12890) );
  NAND2_X1 U14189 ( .A1(n13043), .A2(n13140), .ZN(n11133) );
  AOI22_X1 U14190 ( .A1(n11166), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11253), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11143) );
  AOI22_X1 U14191 ( .A1(n10603), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11254), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11142) );
  AOI22_X1 U14192 ( .A1(n11255), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10558), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11140) );
  NAND2_X1 U14193 ( .A1(n11256), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11139) );
  NAND2_X1 U14194 ( .A1(n11257), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11138) );
  AND3_X1 U14195 ( .A1(n11140), .A2(n11139), .A3(n11138), .ZN(n11141) );
  NAND3_X1 U14196 ( .A1(n11143), .A2(n11142), .A3(n11141), .ZN(n11149) );
  AOI22_X1 U14197 ( .A1(n11264), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11147) );
  AOI22_X1 U14198 ( .A1(n11265), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9887), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11146) );
  AOI22_X1 U14199 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10536), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11145) );
  AOI22_X1 U14200 ( .A1(n10553), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11144) );
  NAND4_X1 U14201 ( .A1(n11147), .A2(n11146), .A3(n11145), .A4(n11144), .ZN(
        n11148) );
  NOR2_X1 U14202 ( .A1(n11149), .A2(n11148), .ZN(n14913) );
  AOI22_X1 U14203 ( .A1(n11166), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n11253), .ZN(n11155) );
  AOI22_X1 U14204 ( .A1(n10603), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n11254), .ZN(n11154) );
  AOI22_X1 U14205 ( .A1(n11255), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n10558), .ZN(n11152) );
  NAND2_X1 U14206 ( .A1(n11256), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11151) );
  NAND2_X1 U14207 ( .A1(n11257), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11150) );
  AND3_X1 U14208 ( .A1(n11152), .A2(n11151), .A3(n11150), .ZN(n11153) );
  NAND3_X1 U14209 ( .A1(n11155), .A2(n11154), .A3(n11153), .ZN(n11161) );
  AOI22_X1 U14210 ( .A1(n11264), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11159) );
  AOI22_X1 U14211 ( .A1(n11265), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9887), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11158) );
  AOI22_X1 U14212 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10536), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11157) );
  AOI22_X1 U14213 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10553), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11156) );
  NAND4_X1 U14214 ( .A1(n11159), .A2(n11158), .A3(n11157), .A4(n11156), .ZN(
        n11160) );
  OR2_X1 U14215 ( .A1(n11161), .A2(n11160), .ZN(n13466) );
  AOI22_X1 U14216 ( .A1(n11264), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11165) );
  AOI22_X1 U14217 ( .A1(n11265), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9887), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11164) );
  AOI22_X1 U14218 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10536), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11163) );
  AOI22_X1 U14219 ( .A1(n10553), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11162) );
  NAND4_X1 U14220 ( .A1(n11165), .A2(n11164), .A3(n11163), .A4(n11162), .ZN(
        n11177) );
  INV_X1 U14221 ( .A(n11166), .ZN(n11223) );
  INV_X1 U14222 ( .A(n11253), .ZN(n11221) );
  INV_X1 U14223 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11167) );
  OAI22_X1 U14224 ( .A1(n11223), .A2(n11168), .B1(n11221), .B2(n11167), .ZN(
        n11176) );
  INV_X1 U14225 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11170) );
  INV_X1 U14226 ( .A(n11254), .ZN(n11224) );
  INV_X1 U14227 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11169) );
  OAI22_X1 U14228 ( .A1(n11225), .A2(n11170), .B1(n11224), .B2(n11169), .ZN(
        n11175) );
  AOI22_X1 U14229 ( .A1(n11255), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10558), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11173) );
  NAND2_X1 U14230 ( .A1(n11256), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11172) );
  NAND2_X1 U14231 ( .A1(n11257), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11171) );
  NAND3_X1 U14232 ( .A1(n11173), .A2(n11172), .A3(n11171), .ZN(n11174) );
  NOR4_X1 U14233 ( .A1(n11177), .A2(n11176), .A3(n11175), .A4(n11174), .ZN(
        n14900) );
  AOI22_X1 U14234 ( .A1(n11166), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11253), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11183) );
  AOI22_X1 U14235 ( .A1(n10603), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11254), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11182) );
  AOI22_X1 U14236 ( .A1(n11255), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10558), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11180) );
  NAND2_X1 U14237 ( .A1(n11256), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11179) );
  NAND2_X1 U14238 ( .A1(n11257), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11178) );
  AND3_X1 U14239 ( .A1(n11180), .A2(n11179), .A3(n11178), .ZN(n11181) );
  NAND3_X1 U14240 ( .A1(n11183), .A2(n11182), .A3(n11181), .ZN(n11189) );
  AOI22_X1 U14241 ( .A1(n11264), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11187) );
  AOI22_X1 U14242 ( .A1(n11265), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9887), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11186) );
  AOI22_X1 U14243 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10536), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11185) );
  AOI22_X1 U14244 ( .A1(n10553), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11184) );
  NAND4_X1 U14245 ( .A1(n11187), .A2(n11186), .A3(n11185), .A4(n11184), .ZN(
        n11188) );
  OR2_X1 U14246 ( .A1(n11189), .A2(n11188), .ZN(n14894) );
  AOI22_X1 U14247 ( .A1(n11166), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11253), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11195) );
  AOI22_X1 U14248 ( .A1(n10603), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11254), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11194) );
  AOI22_X1 U14249 ( .A1(n11255), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10558), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11192) );
  NAND2_X1 U14250 ( .A1(n11256), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11191) );
  NAND2_X1 U14251 ( .A1(n11257), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11190) );
  AND3_X1 U14252 ( .A1(n11192), .A2(n11191), .A3(n11190), .ZN(n11193) );
  NAND3_X1 U14253 ( .A1(n11195), .A2(n11194), .A3(n11193), .ZN(n11201) );
  AOI22_X1 U14254 ( .A1(n11264), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11199) );
  AOI22_X1 U14255 ( .A1(n11265), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9887), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11198) );
  AOI22_X1 U14256 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10536), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11197) );
  AOI22_X1 U14257 ( .A1(n10553), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11196) );
  NAND4_X1 U14258 ( .A1(n11199), .A2(n11198), .A3(n11197), .A4(n11196), .ZN(
        n11200) );
  NOR2_X1 U14259 ( .A1(n11201), .A2(n11200), .ZN(n14889) );
  AOI22_X1 U14260 ( .A1(n11264), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11205) );
  AOI22_X1 U14261 ( .A1(n11265), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9887), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11204) );
  AOI22_X1 U14262 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10536), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11203) );
  AOI22_X1 U14263 ( .A1(n10553), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11202) );
  NAND4_X1 U14264 ( .A1(n11205), .A2(n11204), .A3(n11203), .A4(n11202), .ZN(
        n11216) );
  AOI22_X1 U14265 ( .A1(n11255), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10558), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11208) );
  NAND2_X1 U14266 ( .A1(n11256), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11207) );
  NAND2_X1 U14267 ( .A1(n11257), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11206) );
  NAND3_X1 U14268 ( .A1(n11208), .A2(n11207), .A3(n11206), .ZN(n11215) );
  INV_X1 U14269 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11209) );
  OAI22_X1 U14270 ( .A1(n11223), .A2(n11210), .B1(n11221), .B2(n11209), .ZN(
        n11214) );
  INV_X1 U14271 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11212) );
  INV_X1 U14272 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11211) );
  OAI22_X1 U14273 ( .A1(n11225), .A2(n11212), .B1(n11224), .B2(n11211), .ZN(
        n11213) );
  OR4_X1 U14274 ( .A1(n11216), .A2(n11215), .A3(n11214), .A4(n11213), .ZN(
        n14884) );
  AOI22_X1 U14275 ( .A1(n11264), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11220) );
  AOI22_X1 U14276 ( .A1(n11265), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9887), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11219) );
  AOI22_X1 U14277 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n10536), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11218) );
  AOI22_X1 U14278 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10553), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11217) );
  NAND4_X1 U14279 ( .A1(n11220), .A2(n11219), .A3(n11218), .A4(n11217), .ZN(
        n11232) );
  INV_X1 U14280 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11383) );
  INV_X1 U14281 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11222) );
  OAI22_X1 U14282 ( .A1(n11223), .A2(n11383), .B1(n11222), .B2(n11221), .ZN(
        n11231) );
  INV_X1 U14283 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13582) );
  INV_X1 U14284 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13161) );
  OAI22_X1 U14285 ( .A1(n11225), .A2(n13582), .B1(n13161), .B2(n11224), .ZN(
        n11230) );
  AOI22_X1 U14286 ( .A1(n11255), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n10558), .ZN(n11228) );
  NAND2_X1 U14287 ( .A1(n11256), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11227) );
  NAND2_X1 U14288 ( .A1(n11257), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11226) );
  NAND3_X1 U14289 ( .A1(n11228), .A2(n11227), .A3(n11226), .ZN(n11229) );
  NOR4_X1 U14290 ( .A1(n11232), .A2(n11231), .A3(n11230), .A4(n11229), .ZN(
        n14879) );
  INV_X1 U14291 ( .A(n11233), .ZN(n11373) );
  INV_X1 U14292 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11236) );
  OAI21_X1 U14293 ( .B1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n11234), .ZN(n11413) );
  OAI211_X1 U14294 ( .C1(n11373), .C2(n11236), .A(n11235), .B(n11413), .ZN(
        n11237) );
  INV_X1 U14295 ( .A(n11237), .ZN(n11242) );
  AOI22_X1 U14296 ( .A1(n11408), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12868), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11241) );
  AOI22_X1 U14297 ( .A1(n9841), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11409), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11240) );
  AOI22_X1 U14298 ( .A1(n11420), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10473), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11239) );
  NAND4_X1 U14299 ( .A1(n11242), .A2(n11241), .A3(n11240), .A4(n11239), .ZN(
        n11252) );
  AOI22_X1 U14300 ( .A1(n11408), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12868), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11250) );
  AOI22_X1 U14301 ( .A1(n11419), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11420), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11249) );
  AOI22_X1 U14302 ( .A1(n9841), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11409), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11248) );
  INV_X1 U14303 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11245) );
  INV_X1 U14304 ( .A(n10473), .ZN(n11391) );
  INV_X1 U14305 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11243) );
  OR2_X1 U14306 ( .A1(n11391), .A2(n11243), .ZN(n11244) );
  INV_X1 U14307 ( .A(n11413), .ZN(n11392) );
  OAI211_X1 U14308 ( .C1(n9819), .C2(n11245), .A(n11244), .B(n11392), .ZN(
        n11246) );
  INV_X1 U14309 ( .A(n11246), .ZN(n11247) );
  NAND4_X1 U14310 ( .A1(n11250), .A2(n11249), .A3(n11248), .A4(n11247), .ZN(
        n11251) );
  AND2_X1 U14311 ( .A1(n11252), .A2(n11251), .ZN(n11293) );
  NAND2_X1 U14312 ( .A1(n14748), .A2(n11293), .ZN(n11272) );
  AOI22_X1 U14313 ( .A1(n11166), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n11253), .ZN(n11263) );
  AOI22_X1 U14314 ( .A1(n10603), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n11254), .ZN(n11262) );
  AOI22_X1 U14315 ( .A1(n11255), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n10558), .ZN(n11260) );
  NAND2_X1 U14316 ( .A1(n11256), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11259) );
  NAND2_X1 U14317 ( .A1(n11257), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11258) );
  AND3_X1 U14318 ( .A1(n11260), .A2(n11259), .A3(n11258), .ZN(n11261) );
  NAND3_X1 U14319 ( .A1(n11263), .A2(n11262), .A3(n11261), .ZN(n11271) );
  AOI22_X1 U14320 ( .A1(n11264), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11269) );
  AOI22_X1 U14321 ( .A1(n11265), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9887), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11268) );
  AOI22_X1 U14322 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n10536), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11267) );
  AOI22_X1 U14323 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10553), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11266) );
  NAND4_X1 U14324 ( .A1(n11269), .A2(n11268), .A3(n11267), .A4(n11266), .ZN(
        n11270) );
  OR2_X1 U14325 ( .A1(n11271), .A2(n11270), .ZN(n11275) );
  XNOR2_X1 U14326 ( .A(n11272), .B(n11275), .ZN(n11296) );
  NAND2_X1 U14327 ( .A1(n19247), .A2(n11293), .ZN(n14874) );
  INV_X1 U14328 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11277) );
  OAI211_X1 U14329 ( .C1(n11373), .C2(n11277), .A(n11276), .B(n11413), .ZN(
        n11278) );
  INV_X1 U14330 ( .A(n11278), .ZN(n11282) );
  AOI22_X1 U14331 ( .A1(n11408), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12868), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11281) );
  AOI22_X1 U14332 ( .A1(n10473), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11409), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11280) );
  AOI22_X1 U14333 ( .A1(n11420), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9841), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11279) );
  NAND4_X1 U14334 ( .A1(n11282), .A2(n11281), .A3(n11280), .A4(n11279), .ZN(
        n11290) );
  INV_X1 U14335 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13217) );
  OAI211_X1 U14336 ( .C1(n11373), .C2(n13217), .A(n11392), .B(n11283), .ZN(
        n11284) );
  INV_X1 U14337 ( .A(n11284), .ZN(n11288) );
  AOI22_X1 U14338 ( .A1(n11408), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12868), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11287) );
  AOI22_X1 U14339 ( .A1(n10473), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11409), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11286) );
  AOI22_X1 U14340 ( .A1(n11420), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9841), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11285) );
  NAND4_X1 U14341 ( .A1(n11288), .A2(n11287), .A3(n11286), .A4(n11285), .ZN(
        n11289) );
  AND2_X1 U14342 ( .A1(n11290), .A2(n11289), .ZN(n11292) );
  NAND2_X1 U14343 ( .A1(n11291), .A2(n11292), .ZN(n11297) );
  OAI211_X1 U14344 ( .C1(n11291), .C2(n11292), .A(n11297), .B(n11360), .ZN(
        n14866) );
  NAND2_X1 U14345 ( .A1(n19247), .A2(n11292), .ZN(n14868) );
  INV_X1 U14346 ( .A(n11293), .ZN(n11294) );
  NOR2_X1 U14347 ( .A1(n14868), .A2(n11294), .ZN(n11295) );
  INV_X1 U14348 ( .A(n11297), .ZN(n11314) );
  INV_X1 U14349 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11299) );
  OAI211_X1 U14350 ( .C1(n11373), .C2(n11299), .A(n11298), .B(n11413), .ZN(
        n11300) );
  INV_X1 U14351 ( .A(n11300), .ZN(n11304) );
  AOI22_X1 U14352 ( .A1(n11408), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12868), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11303) );
  AOI22_X1 U14353 ( .A1(n10473), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11409), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11302) );
  AOI22_X1 U14354 ( .A1(n11420), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9841), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11301) );
  NAND4_X1 U14355 ( .A1(n11304), .A2(n11303), .A3(n11302), .A4(n11301), .ZN(
        n11313) );
  INV_X1 U14356 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11306) );
  OAI211_X1 U14357 ( .C1(n11373), .C2(n11306), .A(n11392), .B(n11305), .ZN(
        n11307) );
  INV_X1 U14358 ( .A(n11307), .ZN(n11311) );
  AOI22_X1 U14359 ( .A1(n11408), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12868), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11310) );
  AOI22_X1 U14360 ( .A1(n10473), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11409), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11309) );
  AOI22_X1 U14361 ( .A1(n11420), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9841), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11308) );
  NAND4_X1 U14362 ( .A1(n11311), .A2(n11310), .A3(n11309), .A4(n11308), .ZN(
        n11312) );
  AND2_X1 U14363 ( .A1(n11313), .A2(n11312), .ZN(n11315) );
  NAND2_X1 U14364 ( .A1(n11314), .A2(n11315), .ZN(n11338) );
  OAI211_X1 U14365 ( .C1(n11314), .C2(n11315), .A(n11360), .B(n11338), .ZN(
        n11317) );
  INV_X1 U14366 ( .A(n11315), .ZN(n11316) );
  NOR2_X1 U14367 ( .A1(n14748), .A2(n11316), .ZN(n14858) );
  NAND2_X1 U14368 ( .A1(n14855), .A2(n14858), .ZN(n14857) );
  OAI211_X1 U14369 ( .C1(n11373), .C2(n11322), .A(n11321), .B(n11413), .ZN(
        n11323) );
  INV_X1 U14370 ( .A(n11323), .ZN(n11327) );
  AOI22_X1 U14371 ( .A1(n11408), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12868), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11326) );
  AOI22_X1 U14372 ( .A1(n10473), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11409), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11325) );
  AOI22_X1 U14373 ( .A1(n11420), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9841), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11324) );
  NAND4_X1 U14374 ( .A1(n11327), .A2(n11326), .A3(n11325), .A4(n11324), .ZN(
        n11336) );
  INV_X1 U14375 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11329) );
  OAI211_X1 U14376 ( .C1(n11373), .C2(n11329), .A(n11392), .B(n11328), .ZN(
        n11330) );
  INV_X1 U14377 ( .A(n11330), .ZN(n11334) );
  AOI22_X1 U14378 ( .A1(n11408), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12868), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11333) );
  AOI22_X1 U14379 ( .A1(n10473), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11409), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11332) );
  AOI22_X1 U14380 ( .A1(n11420), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9841), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11331) );
  NAND4_X1 U14381 ( .A1(n11334), .A2(n11333), .A3(n11332), .A4(n11331), .ZN(
        n11335) );
  NAND2_X1 U14382 ( .A1(n11336), .A2(n11335), .ZN(n11340) );
  AOI21_X1 U14383 ( .B1(n11338), .B2(n11340), .A(n11337), .ZN(n11339) );
  INV_X1 U14384 ( .A(n11340), .ZN(n11341) );
  NAND2_X1 U14385 ( .A1(n19247), .A2(n11341), .ZN(n14852) );
  INV_X1 U14386 ( .A(n11343), .ZN(n11361) );
  OAI211_X1 U14387 ( .C1(n11373), .C2(n11345), .A(n11344), .B(n11413), .ZN(
        n11346) );
  INV_X1 U14388 ( .A(n11346), .ZN(n11350) );
  AOI22_X1 U14389 ( .A1(n11408), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12868), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11349) );
  AOI22_X1 U14390 ( .A1(n10473), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11409), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11348) );
  AOI22_X1 U14391 ( .A1(n11420), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9841), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11347) );
  NAND4_X1 U14392 ( .A1(n11350), .A2(n11349), .A3(n11348), .A4(n11347), .ZN(
        n11359) );
  INV_X1 U14393 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11352) );
  OAI211_X1 U14394 ( .C1(n11373), .C2(n11352), .A(n11392), .B(n11351), .ZN(
        n11353) );
  INV_X1 U14395 ( .A(n11353), .ZN(n11357) );
  AOI22_X1 U14396 ( .A1(n11408), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12868), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11356) );
  AOI22_X1 U14397 ( .A1(n10473), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11409), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11355) );
  AOI22_X1 U14398 ( .A1(n11420), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9841), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11354) );
  NAND4_X1 U14399 ( .A1(n11357), .A2(n11356), .A3(n11355), .A4(n11354), .ZN(
        n11358) );
  AND2_X1 U14400 ( .A1(n11359), .A2(n11358), .ZN(n11364) );
  NAND2_X1 U14401 ( .A1(n11361), .A2(n11364), .ZN(n14834) );
  OAI211_X1 U14402 ( .C1(n11361), .C2(n11364), .A(n14834), .B(n11360), .ZN(
        n11362) );
  OAI211_X1 U14403 ( .C1(n11373), .C2(n11366), .A(n11365), .B(n11413), .ZN(
        n11367) );
  INV_X1 U14404 ( .A(n11367), .ZN(n11371) );
  AOI22_X1 U14405 ( .A1(n11408), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12868), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11370) );
  AOI22_X1 U14406 ( .A1(n10473), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11409), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11369) );
  AOI22_X1 U14407 ( .A1(n11420), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9841), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11368) );
  NAND4_X1 U14408 ( .A1(n11371), .A2(n11370), .A3(n11369), .A4(n11368), .ZN(
        n11380) );
  INV_X1 U14409 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13359) );
  OAI211_X1 U14410 ( .C1(n11373), .C2(n13359), .A(n11392), .B(n11372), .ZN(
        n11374) );
  INV_X1 U14411 ( .A(n11374), .ZN(n11378) );
  AOI22_X1 U14412 ( .A1(n11408), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12868), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11377) );
  AOI22_X1 U14413 ( .A1(n10473), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11409), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11376) );
  AOI22_X1 U14414 ( .A1(n11420), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9841), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11375) );
  NAND4_X1 U14415 ( .A1(n11378), .A2(n11377), .A3(n11376), .A4(n11375), .ZN(
        n11379) );
  AND2_X1 U14416 ( .A1(n11380), .A2(n11379), .ZN(n14835) );
  INV_X1 U14417 ( .A(n14829), .ZN(n11404) );
  INV_X1 U14418 ( .A(n14834), .ZN(n11382) );
  AND2_X1 U14419 ( .A1(n14748), .A2(n14835), .ZN(n11381) );
  AND2_X1 U14420 ( .A1(n11382), .A2(n11381), .ZN(n11402) );
  AOI22_X1 U14421 ( .A1(n11408), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12868), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11389) );
  AOI22_X1 U14422 ( .A1(n11419), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10473), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11388) );
  AOI22_X1 U14423 ( .A1(n11420), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9841), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11387) );
  INV_X1 U14424 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13590) );
  OR2_X1 U14425 ( .A1(n9845), .A2(n11383), .ZN(n11384) );
  OAI211_X1 U14426 ( .C1(n9819), .C2(n13590), .A(n11384), .B(n11413), .ZN(
        n11385) );
  INV_X1 U14427 ( .A(n11385), .ZN(n11386) );
  NAND4_X1 U14428 ( .A1(n11389), .A2(n11388), .A3(n11387), .A4(n11386), .ZN(
        n11400) );
  AOI22_X1 U14429 ( .A1(n11419), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11409), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11397) );
  AOI22_X1 U14430 ( .A1(n11420), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9841), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11396) );
  INV_X1 U14431 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13589) );
  INV_X1 U14432 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11390) );
  OR2_X1 U14433 ( .A1(n11391), .A2(n11390), .ZN(n11393) );
  OAI211_X1 U14434 ( .C1(n12869), .C2(n13589), .A(n11393), .B(n11392), .ZN(
        n11394) );
  INV_X1 U14435 ( .A(n11394), .ZN(n11395) );
  NAND4_X1 U14436 ( .A1(n11398), .A2(n11397), .A3(n11396), .A4(n11395), .ZN(
        n11399) );
  AND2_X1 U14437 ( .A1(n11400), .A2(n11399), .ZN(n11401) );
  OAI21_X1 U14438 ( .B1(n11402), .B2(n11401), .A(n11405), .ZN(n14830) );
  INV_X1 U14439 ( .A(n14830), .ZN(n11403) );
  NAND2_X1 U14440 ( .A1(n11404), .A2(n11403), .ZN(n14828) );
  AOI22_X1 U14441 ( .A1(n11419), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10473), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11407) );
  AOI22_X1 U14442 ( .A1(n11420), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9841), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11406) );
  NAND2_X1 U14443 ( .A1(n11407), .A2(n11406), .ZN(n11426) );
  INV_X1 U14444 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11412) );
  AOI21_X1 U14445 ( .B1(n11409), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n11413), .ZN(n11410) );
  OAI211_X1 U14446 ( .C1(n12869), .C2(n11412), .A(n11411), .B(n11410), .ZN(
        n11425) );
  OAI21_X1 U14447 ( .B1(n9845), .B2(n10751), .A(n11413), .ZN(n11418) );
  INV_X1 U14448 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11415) );
  INV_X1 U14449 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11414) );
  OAI22_X1 U14450 ( .A1(n11416), .A2(n11415), .B1(n12869), .B2(n11414), .ZN(
        n11417) );
  AOI22_X1 U14451 ( .A1(n11419), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10473), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11422) );
  AOI22_X1 U14452 ( .A1(n11420), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9841), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11421) );
  NAND3_X1 U14453 ( .A1(n11423), .A2(n11422), .A3(n11421), .ZN(n11424) );
  NAND2_X1 U14454 ( .A1(n12490), .A2(n11429), .ZN(n11446) );
  AND2_X1 U14455 ( .A1(n11430), .A2(n11429), .ZN(n11445) );
  NAND2_X1 U14456 ( .A1(n11431), .A2(n13216), .ZN(n11432) );
  MUX2_X1 U14457 ( .A(n11432), .B(n10906), .S(n11434), .Z(n11443) );
  INV_X1 U14458 ( .A(n11434), .ZN(n11441) );
  OAI21_X1 U14459 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19964), .A(
        n11435), .ZN(n12484) );
  INV_X1 U14460 ( .A(n12484), .ZN(n11437) );
  OAI211_X1 U14461 ( .C1(n13216), .C2(n11437), .A(n16347), .B(n11436), .ZN(
        n11440) );
  OAI21_X1 U14462 ( .B1(n11438), .B2(n12484), .A(n12679), .ZN(n11439) );
  OAI211_X1 U14463 ( .C1(n11433), .C2(n11441), .A(n11440), .B(n11439), .ZN(
        n11442) );
  NAND2_X1 U14464 ( .A1(n11443), .A2(n11442), .ZN(n11444) );
  AOI22_X1 U14465 ( .A1(n11446), .A2(n10906), .B1(n11445), .B2(n11444), .ZN(
        n11447) );
  NOR2_X1 U14466 ( .A1(n11447), .A2(n11449), .ZN(n11448) );
  MUX2_X1 U14467 ( .A(n11448), .B(n15663), .S(n18909), .Z(n12645) );
  NAND2_X1 U14468 ( .A1(n11453), .A2(n19252), .ZN(n11454) );
  NAND2_X1 U14469 ( .A1(n11452), .A2(n11454), .ZN(n11464) );
  INV_X1 U14470 ( .A(n11455), .ZN(n11456) );
  NAND2_X1 U14471 ( .A1(n11456), .A2(n19247), .ZN(n11465) );
  NAND2_X1 U14472 ( .A1(n10915), .A2(n10930), .ZN(n11457) );
  AND2_X1 U14473 ( .A1(n11457), .A2(n19252), .ZN(n11458) );
  AOI21_X1 U14474 ( .B1(n11465), .B2(n11458), .A(n10909), .ZN(n11463) );
  INV_X1 U14475 ( .A(n11459), .ZN(n11460) );
  NAND3_X1 U14476 ( .A1(n11461), .A2(n11460), .A3(n10930), .ZN(n11462) );
  AND2_X1 U14477 ( .A1(n19247), .A2(n10915), .ZN(n12494) );
  NAND2_X1 U14478 ( .A1(n11462), .A2(n12494), .ZN(n12674) );
  NAND4_X1 U14479 ( .A1(n11451), .A2(n11464), .A3(n11463), .A4(n12674), .ZN(
        n12651) );
  INV_X1 U14480 ( .A(n12651), .ZN(n11467) );
  INV_X1 U14481 ( .A(n11465), .ZN(n11466) );
  NAND2_X1 U14482 ( .A1(n11467), .A2(n11466), .ZN(n16353) );
  INV_X1 U14483 ( .A(n10901), .ZN(n16350) );
  NAND4_X1 U14484 ( .A1(n16350), .A2(n16348), .A3(n12667), .A4(n19835), .ZN(
        n11468) );
  OAI21_X1 U14485 ( .B1(n12612), .B2(n16353), .A(n11468), .ZN(n12881) );
  AND2_X1 U14486 ( .A1(n11469), .A2(n10920), .ZN(n11470) );
  NAND2_X1 U14487 ( .A1(n12402), .A2(n19137), .ZN(n11487) );
  NOR4_X1 U14488 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n11475) );
  NOR4_X1 U14489 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n11474) );
  NOR4_X1 U14490 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n11473) );
  NOR4_X1 U14491 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n11472) );
  NAND4_X1 U14492 ( .A1(n11475), .A2(n11474), .A3(n11473), .A4(n11472), .ZN(
        n11480) );
  NOR4_X1 U14493 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n11478) );
  NOR4_X1 U14494 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n11477) );
  NOR4_X1 U14495 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n11476) );
  INV_X1 U14496 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19861) );
  NAND4_X1 U14497 ( .A1(n11478), .A2(n11477), .A3(n11476), .A4(n19861), .ZN(
        n11479) );
  AOI22_X1 U14498 ( .A1(n13155), .A2(BUF1_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n13153), .ZN(n19140) );
  AND2_X1 U14499 ( .A1(n19267), .A2(n10930), .ZN(n11481) );
  AOI22_X1 U14500 ( .A1(n15221), .A2(n19177), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n19176), .ZN(n11484) );
  NOR2_X1 U14501 ( .A1(n9978), .A2(n11101), .ZN(n11482) );
  AOI22_X1 U14502 ( .A1(n19128), .A2(BUF2_REG_30__SCAN_IN), .B1(n19129), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n11483) );
  OAI211_X1 U14503 ( .C1(n19140), .C2(n14988), .A(n11484), .B(n11483), .ZN(
        n11485) );
  INV_X1 U14504 ( .A(n11485), .ZN(n11486) );
  NAND2_X1 U14505 ( .A1(n11487), .A2(n11486), .ZN(P2_U2889) );
  XNOR2_X1 U14506 ( .A(n20843), .B(P1_STATE_REG_1__SCAN_IN), .ZN(n12696) );
  NOR2_X4 U14507 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13093) );
  NAND2_X1 U14508 ( .A1(n12244), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11493) );
  AND2_X2 U14509 ( .A1(n11494), .A2(n13093), .ZN(n11770) );
  BUF_X4 U14510 ( .A(n11770), .Z(n12042) );
  NAND2_X1 U14511 ( .A1(n12042), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11492) );
  AND2_X2 U14512 ( .A1(n11506), .A2(n11500), .ZN(n11765) );
  BUF_X4 U14513 ( .A(n11765), .Z(n12106) );
  NAND2_X1 U14514 ( .A1(n12106), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11491) );
  NAND2_X1 U14515 ( .A1(n11654), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11490) );
  NAND2_X1 U14516 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11499) );
  AND2_X2 U14517 ( .A1(n11500), .A2(n11495), .ZN(n11578) );
  NAND2_X1 U14518 ( .A1(n11578), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11498) );
  NAND2_X1 U14519 ( .A1(n11752), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11497) );
  AND2_X2 U14520 ( .A1(n13093), .A2(n11505), .ZN(n11561) );
  NAND2_X1 U14521 ( .A1(n11561), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11496) );
  NAND2_X1 U14522 ( .A1(n12249), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11504) );
  AND2_X2 U14523 ( .A1(n11500), .A2(n13094), .ZN(n11607) );
  NAND2_X1 U14524 ( .A1(n11607), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11503) );
  NAND2_X1 U14525 ( .A1(n12147), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11502) );
  AND2_X4 U14526 ( .A1(n14735), .A2(n13094), .ZN(n13091) );
  NAND2_X1 U14527 ( .A1(n13091), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11501) );
  AND2_X2 U14528 ( .A1(n11506), .A2(n11505), .ZN(n11938) );
  NAND2_X1 U14529 ( .A1(n11938), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11512) );
  NOR2_X1 U14530 ( .A1(n11811), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11507) );
  AND2_X2 U14531 ( .A1(n11507), .A2(n13096), .ZN(n11926) );
  NAND2_X1 U14532 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11511) );
  AND2_X4 U14533 ( .A1(n13093), .A2(n14735), .ZN(n12285) );
  NAND2_X1 U14534 ( .A1(n12285), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11510) );
  AND2_X2 U14535 ( .A1(n13096), .A2(n11508), .ZN(n11591) );
  NAND2_X1 U14536 ( .A1(n12128), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11509) );
  NAND4_X4 U14537 ( .A1(n11516), .A2(n11515), .A3(n11514), .A4(n11513), .ZN(
        n13435) );
  NAND2_X1 U14538 ( .A1(n12106), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11520) );
  NAND2_X1 U14539 ( .A1(n11938), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11519) );
  NAND2_X1 U14540 ( .A1(n12249), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11518) );
  NAND2_X1 U14541 ( .A1(n11578), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11517) );
  NAND2_X1 U14542 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11524) );
  NAND2_X1 U14543 ( .A1(n11607), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11523) );
  NAND2_X1 U14544 ( .A1(n12134), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11522) );
  NAND2_X1 U14545 ( .A1(n12244), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11521) );
  NAND2_X1 U14546 ( .A1(n11752), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11528) );
  NAND2_X1 U14547 ( .A1(n11654), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11527) );
  NAND2_X1 U14548 ( .A1(n12147), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11525) );
  NAND2_X1 U14549 ( .A1(n11561), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11532) );
  NAND2_X1 U14550 ( .A1(n12285), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11531) );
  NAND2_X1 U14551 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11530) );
  NAND2_X1 U14552 ( .A1(n12128), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11529) );
  NAND2_X1 U14553 ( .A1(n12042), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11540) );
  NAND2_X1 U14554 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11539) );
  NAND2_X1 U14555 ( .A1(n12106), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11538) );
  NAND2_X1 U14556 ( .A1(n12244), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11537) );
  NAND2_X1 U14557 ( .A1(n11654), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11544) );
  NAND2_X1 U14558 ( .A1(n11578), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11543) );
  NAND2_X1 U14559 ( .A1(n11752), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11542) );
  NAND2_X1 U14560 ( .A1(n12147), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11541) );
  NAND2_X1 U14561 ( .A1(n11561), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11547) );
  NAND2_X1 U14562 ( .A1(n11607), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11546) );
  NAND2_X1 U14563 ( .A1(n12249), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11545) );
  NAND3_X1 U14564 ( .A1(n11547), .A2(n11546), .A3(n11545), .ZN(n11548) );
  NAND2_X1 U14565 ( .A1(n11938), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11552) );
  NAND2_X1 U14566 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11551) );
  NAND2_X1 U14567 ( .A1(n12285), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11550) );
  NAND2_X1 U14568 ( .A1(n12128), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11549) );
  NOR2_X1 U14569 ( .A1(n14328), .A2(n12792), .ZN(n11577) );
  BUF_X2 U14570 ( .A(n11954), .Z(n12294) );
  BUF_X2 U14571 ( .A(n11770), .Z(n12293) );
  AOI22_X1 U14572 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11560) );
  BUF_X2 U14573 ( .A(n11765), .Z(n12295) );
  AOI22_X1 U14574 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12244), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11559) );
  AOI22_X1 U14575 ( .A1(n11654), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11752), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11558) );
  AOI22_X1 U14576 ( .A1(n11578), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12147), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11557) );
  NAND4_X1 U14577 ( .A1(n11560), .A2(n11559), .A3(n11558), .A4(n11557), .ZN(
        n11567) );
  AOI22_X1 U14578 ( .A1(n12249), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11561), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11565) );
  AOI22_X1 U14579 ( .A1(n11938), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12285), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11564) );
  BUF_X4 U14580 ( .A(n11591), .Z(n12287) );
  AOI22_X1 U14581 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11563) );
  AOI22_X1 U14582 ( .A1(n11607), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13091), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11562) );
  NAND4_X1 U14583 ( .A1(n11565), .A2(n11564), .A3(n11563), .A4(n11562), .ZN(
        n11566) );
  OR2_X2 U14584 ( .A1(n11567), .A2(n11566), .ZN(n13079) );
  AOI22_X1 U14585 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12244), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11570) );
  AOI22_X1 U14586 ( .A1(n11654), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11752), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11569) );
  AOI22_X1 U14587 ( .A1(n12249), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11561), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11575) );
  AOI22_X1 U14588 ( .A1(n11938), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12285), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11574) );
  AOI22_X1 U14589 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11573) );
  AOI22_X1 U14590 ( .A1(n11607), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13091), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11572) );
  AOI22_X1 U14591 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11582) );
  AOI22_X1 U14592 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12244), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11581) );
  AOI22_X1 U14593 ( .A1(n11654), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11752), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11580) );
  AOI22_X1 U14594 ( .A1(n11578), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12147), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11579) );
  AOI22_X1 U14595 ( .A1(n12249), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11561), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11586) );
  AOI22_X1 U14596 ( .A1(n11938), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12285), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11585) );
  AOI22_X1 U14597 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11591), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11584) );
  AOI22_X1 U14598 ( .A1(n11607), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13091), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11583) );
  AOI22_X1 U14599 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11590) );
  AOI22_X1 U14600 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12244), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11589) );
  AOI22_X1 U14601 ( .A1(n11654), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11752), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11588) );
  AOI22_X1 U14602 ( .A1(n11578), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12147), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11587) );
  NAND4_X1 U14603 ( .A1(n11590), .A2(n11589), .A3(n11588), .A4(n11587), .ZN(
        n11597) );
  AOI22_X1 U14604 ( .A1(n11938), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12285), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11594) );
  AOI22_X1 U14605 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11591), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11593) );
  AOI22_X1 U14606 ( .A1(n11607), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13091), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11592) );
  NAND4_X1 U14607 ( .A1(n11595), .A2(n11594), .A3(n11593), .A4(n11592), .ZN(
        n11596) );
  OR2_X2 U14608 ( .A1(n11597), .A2(n11596), .ZN(n12740) );
  NAND2_X1 U14609 ( .A1(n20248), .A2(n12740), .ZN(n12375) );
  INV_X1 U14610 ( .A(n12375), .ZN(n11598) );
  NAND2_X1 U14611 ( .A1(n12042), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11602) );
  NAND2_X1 U14612 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11601) );
  NAND2_X1 U14613 ( .A1(n12106), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11600) );
  NAND2_X1 U14614 ( .A1(n12244), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11599) );
  NAND2_X1 U14615 ( .A1(n11654), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11606) );
  NAND2_X1 U14616 ( .A1(n11578), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11605) );
  NAND2_X1 U14617 ( .A1(n11752), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11604) );
  NAND2_X1 U14618 ( .A1(n12147), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11603) );
  NAND2_X1 U14619 ( .A1(n12249), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11611) );
  NAND2_X1 U14620 ( .A1(n11607), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11610) );
  NAND2_X1 U14621 ( .A1(n11561), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11609) );
  NAND2_X1 U14622 ( .A1(n13091), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11608) );
  NAND2_X1 U14623 ( .A1(n11938), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11615) );
  NAND2_X1 U14624 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11614) );
  NAND2_X1 U14625 ( .A1(n12128), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11612) );
  NAND4_X4 U14626 ( .A1(n11619), .A2(n11618), .A3(n11617), .A4(n11616), .ZN(
        n12820) );
  NOR2_X4 U14627 ( .A1(n12831), .A2(n11637), .ZN(n14005) );
  OAI21_X1 U14628 ( .B1(n12696), .B2(n13435), .A(n14005), .ZN(n11622) );
  INV_X2 U14629 ( .A(n14010), .ZN(n11621) );
  NAND2_X1 U14630 ( .A1(n11621), .A2(n11620), .ZN(n12826) );
  OR2_X2 U14631 ( .A1(n12826), .A2(n12763), .ZN(n12793) );
  NAND2_X1 U14632 ( .A1(n13079), .A2(n12792), .ZN(n11625) );
  NAND2_X1 U14633 ( .A1(n11623), .A2(n14328), .ZN(n11624) );
  MUX2_X2 U14634 ( .A(n12736), .B(n11624), .S(n20248), .Z(n11627) );
  OR2_X2 U14635 ( .A1(n11629), .A2(n11625), .ZN(n14730) );
  OR2_X1 U14636 ( .A1(n13080), .A2(n12792), .ZN(n11631) );
  NAND2_X1 U14637 ( .A1(n20271), .A2(n11623), .ZN(n11630) );
  AND2_X1 U14638 ( .A1(n11630), .A2(n13079), .ZN(n11647) );
  NAND2_X1 U14639 ( .A1(n12774), .A2(n20263), .ZN(n12757) );
  AND2_X2 U14640 ( .A1(n12740), .A2(n13435), .ZN(n15910) );
  NAND2_X1 U14641 ( .A1(n12736), .A2(n15910), .ZN(n12825) );
  INV_X1 U14642 ( .A(n12740), .ZN(n20256) );
  NAND2_X1 U14643 ( .A1(n20256), .A2(n12820), .ZN(n13050) );
  NAND2_X1 U14644 ( .A1(n12837), .A2(n12820), .ZN(n11644) );
  NAND2_X1 U14645 ( .A1(n13050), .A2(n11644), .ZN(n12772) );
  NOR2_X1 U14646 ( .A1(n11648), .A2(n12772), .ZN(n11635) );
  INV_X1 U14647 ( .A(n13092), .ZN(n11636) );
  NAND2_X1 U14648 ( .A1(n11714), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11639) );
  NAND2_X1 U14649 ( .A1(n16181), .A2(n20902), .ZN(n12738) );
  MUX2_X1 U14650 ( .A(n12738), .B(n15879), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n11638) );
  AND3_X1 U14651 ( .A1(n13080), .A2(n14010), .A3(n12740), .ZN(n11652) );
  NAND2_X1 U14652 ( .A1(n11641), .A2(n12820), .ZN(n11642) );
  NAND2_X1 U14653 ( .A1(n11642), .A2(n13435), .ZN(n11651) );
  INV_X1 U14654 ( .A(n16181), .ZN(n14744) );
  NOR2_X1 U14655 ( .A1(n14744), .A2(n20902), .ZN(n11643) );
  AND2_X1 U14656 ( .A1(n11644), .A2(n11643), .ZN(n11646) );
  NAND2_X1 U14657 ( .A1(n13092), .A2(n20278), .ZN(n12787) );
  OAI211_X1 U14658 ( .C1(n11647), .C2(n15872), .A(n11646), .B(n12787), .ZN(
        n11649) );
  NOR2_X1 U14659 ( .A1(n11649), .A2(n11648), .ZN(n11650) );
  OAI211_X1 U14660 ( .C1(n11640), .C2(n11652), .A(n11651), .B(n11650), .ZN(
        n11701) );
  INV_X1 U14661 ( .A(n11701), .ZN(n11653) );
  AOI22_X1 U14662 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11658) );
  AOI22_X1 U14663 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11657) );
  AOI22_X1 U14664 ( .A1(n11578), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12244), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11656) );
  AOI22_X1 U14665 ( .A1(n12129), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13091), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11655) );
  NAND4_X1 U14666 ( .A1(n11658), .A2(n11657), .A3(n11656), .A4(n11655), .ZN(
        n11664) );
  AOI22_X1 U14667 ( .A1(n11938), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12285), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11662) );
  AOI22_X1 U14668 ( .A1(n12296), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12229), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11661) );
  AOI22_X1 U14669 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11660) );
  AOI22_X1 U14670 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11659) );
  NAND4_X1 U14671 ( .A1(n11662), .A2(n11661), .A3(n11660), .A4(n11659), .ZN(
        n11663) );
  NOR2_X1 U14672 ( .A1(n11751), .A2(n13487), .ZN(n11690) );
  AOI22_X1 U14673 ( .A1(n12129), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11668) );
  AOI22_X1 U14674 ( .A1(n12230), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11667) );
  AOI22_X1 U14675 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12285), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11666) );
  AOI22_X1 U14676 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13091), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11665) );
  NAND4_X1 U14677 ( .A1(n11668), .A2(n11667), .A3(n11666), .A4(n11665), .ZN(
        n11674) );
  AOI22_X1 U14678 ( .A1(n11938), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11672) );
  AOI22_X1 U14679 ( .A1(n12042), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12229), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11671) );
  AOI22_X1 U14680 ( .A1(n12135), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11670) );
  AOI22_X1 U14681 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11669) );
  NAND4_X1 U14682 ( .A1(n11672), .A2(n11671), .A3(n11670), .A4(n11669), .ZN(
        n11673) );
  MUX2_X1 U14683 ( .A(n11690), .B(n13495), .S(n11679), .Z(n11675) );
  INV_X1 U14684 ( .A(n11675), .ZN(n11676) );
  NAND2_X1 U14685 ( .A1(n12355), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11678) );
  AOI21_X1 U14686 ( .B1(n20263), .B2(n13487), .A(n20902), .ZN(n11677) );
  OAI211_X1 U14687 ( .C1(n11679), .C2(n12820), .A(n11678), .B(n11677), .ZN(
        n11835) );
  AOI22_X1 U14688 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11683) );
  AOI22_X1 U14689 ( .A1(n12042), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11682) );
  AOI22_X1 U14690 ( .A1(n12230), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11681) );
  AOI22_X1 U14691 ( .A1(n12285), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13091), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11680) );
  NAND4_X1 U14692 ( .A1(n11683), .A2(n11682), .A3(n11681), .A4(n11680), .ZN(
        n11689) );
  BUF_X1 U14693 ( .A(n12244), .Z(n12135) );
  AOI22_X1 U14694 ( .A1(n11938), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11687) );
  AOI22_X1 U14695 ( .A1(n12129), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12229), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11686) );
  AOI22_X1 U14696 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11685) );
  AOI22_X1 U14697 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11684) );
  NAND4_X1 U14698 ( .A1(n11687), .A2(n11686), .A3(n11685), .A4(n11684), .ZN(
        n11688) );
  INV_X1 U14699 ( .A(n11690), .ZN(n11692) );
  NAND2_X1 U14700 ( .A1(n12355), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11691) );
  OAI211_X1 U14701 ( .C1(n11750), .C2(n11706), .A(n11692), .B(n11691), .ZN(
        n11693) );
  NAND2_X1 U14702 ( .A1(n11694), .A2(n11693), .ZN(n11695) );
  INV_X1 U14703 ( .A(n11827), .ZN(n11708) );
  NAND2_X1 U14704 ( .A1(n11714), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11698) );
  NAND2_X1 U14705 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11718) );
  OAI21_X1 U14706 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n11718), .ZN(n20559) );
  OR2_X1 U14707 ( .A1(n15879), .A2(n20325), .ZN(n11711) );
  OAI21_X1 U14708 ( .B1(n12738), .B2(n20559), .A(n11711), .ZN(n11696) );
  INV_X1 U14709 ( .A(n11696), .ZN(n11697) );
  XNOR2_X2 U14710 ( .A(n11700), .B(n11713), .ZN(n20358) );
  NAND2_X2 U14711 ( .A1(n20358), .A2(n11703), .ZN(n11728) );
  INV_X1 U14712 ( .A(n20358), .ZN(n11705) );
  INV_X1 U14713 ( .A(n11703), .ZN(n11704) );
  OR2_X1 U14714 ( .A1(n11751), .A2(n11706), .ZN(n11707) );
  AND2_X1 U14715 ( .A1(n11711), .A2(n11710), .ZN(n11712) );
  NAND2_X1 U14716 ( .A1(n11728), .A2(n11726), .ZN(n11722) );
  NAND2_X1 U14717 ( .A1(n11745), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11716) );
  NAND2_X1 U14718 ( .A1(n20826), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11715) );
  NAND2_X1 U14719 ( .A1(n11716), .A2(n11715), .ZN(n11723) );
  INV_X1 U14720 ( .A(n12738), .ZN(n11720) );
  INV_X1 U14721 ( .A(n11718), .ZN(n11717) );
  NAND2_X1 U14722 ( .A1(n11717), .A2(n15858), .ZN(n20591) );
  NAND2_X1 U14723 ( .A1(n11718), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11719) );
  NAND2_X1 U14724 ( .A1(n20591), .A2(n11719), .ZN(n20233) );
  NAND2_X2 U14725 ( .A1(n11722), .A2(n11721), .ZN(n11744) );
  INV_X1 U14726 ( .A(n11723), .ZN(n11727) );
  INV_X1 U14727 ( .A(n11724), .ZN(n11725) );
  NAND4_X1 U14728 ( .A1(n11728), .A2(n11727), .A3(n11726), .A4(n11725), .ZN(
        n11729) );
  AOI22_X1 U14729 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11733) );
  AOI22_X1 U14730 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11732) );
  AOI22_X1 U14731 ( .A1(n12284), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11731) );
  AOI22_X1 U14732 ( .A1(n12230), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11730) );
  NAND4_X1 U14733 ( .A1(n11733), .A2(n11732), .A3(n11731), .A4(n11730), .ZN(
        n11739) );
  AOI22_X1 U14734 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12229), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11737) );
  AOI22_X1 U14735 ( .A1(n11987), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12285), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11736) );
  AOI22_X1 U14736 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11735) );
  AOI22_X1 U14737 ( .A1(n12129), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13091), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11734) );
  NAND4_X1 U14738 ( .A1(n11737), .A2(n11736), .A3(n11735), .A4(n11734), .ZN(
        n11738) );
  AOI22_X1 U14739 ( .A1(n11741), .A2(n11740), .B1(n12355), .B2(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11742) );
  NAND2_X1 U14740 ( .A1(n11745), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11749) );
  NAND3_X1 U14741 ( .A1(n20634), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20470) );
  NOR3_X1 U14742 ( .A1(n20634), .A2(n15858), .A3(n20325), .ZN(n20772) );
  INV_X1 U14743 ( .A(n20772), .ZN(n20763) );
  INV_X1 U14744 ( .A(n20815), .ZN(n11746) );
  OAI21_X1 U14745 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20492), .A(
        n11746), .ZN(n20501) );
  OAI22_X1 U14746 ( .A1(n12738), .A2(n20501), .B1(n15879), .B2(n20634), .ZN(
        n11747) );
  INV_X1 U14747 ( .A(n11747), .ZN(n11748) );
  XNOR2_X2 U14748 ( .A(n11744), .B(n20389), .ZN(n20500) );
  AOI22_X1 U14749 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12134), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11756) );
  AOI22_X1 U14750 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11755) );
  AOI22_X1 U14751 ( .A1(n12284), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11754) );
  AOI22_X1 U14752 ( .A1(n12230), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11753) );
  NAND4_X1 U14753 ( .A1(n11756), .A2(n11755), .A3(n11754), .A4(n11753), .ZN(
        n11762) );
  AOI22_X1 U14754 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12229), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11760) );
  AOI22_X1 U14755 ( .A1(n11987), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12285), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11759) );
  AOI22_X1 U14756 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11758) );
  AOI22_X1 U14757 ( .A1(n12129), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13091), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11757) );
  NAND4_X1 U14758 ( .A1(n11760), .A2(n11759), .A3(n11758), .A4(n11757), .ZN(
        n11761) );
  AOI22_X1 U14759 ( .A1(n12334), .A2(n13337), .B1(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n12355), .ZN(n11763) );
  AOI22_X1 U14760 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12106), .B1(
        n12230), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11769) );
  AOI22_X1 U14761 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n12129), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11768) );
  AOI22_X1 U14762 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11767) );
  AOI22_X1 U14763 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12135), .B1(
        n12285), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11766) );
  NAND4_X1 U14764 ( .A1(n11769), .A2(n11768), .A3(n11767), .A4(n11766), .ZN(
        n11776) );
  AOI22_X1 U14765 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12042), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11774) );
  AOI22_X1 U14766 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12229), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11773) );
  AOI22_X1 U14767 ( .A1(n11987), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11772) );
  AOI22_X1 U14768 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12112), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11771) );
  NAND4_X1 U14769 ( .A1(n11774), .A2(n11773), .A3(n11772), .A4(n11771), .ZN(
        n11775) );
  NAND2_X1 U14770 ( .A1(n12334), .A2(n13336), .ZN(n11778) );
  NAND2_X1 U14771 ( .A1(n12355), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11777) );
  NAND2_X1 U14772 ( .A1(n11778), .A2(n11777), .ZN(n11849) );
  AOI22_X1 U14773 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12134), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11782) );
  AOI22_X1 U14774 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11781) );
  AOI22_X1 U14775 ( .A1(n12284), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11780) );
  AOI22_X1 U14776 ( .A1(n12230), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11779) );
  NAND4_X1 U14777 ( .A1(n11782), .A2(n11781), .A3(n11780), .A4(n11779), .ZN(
        n11788) );
  AOI22_X1 U14778 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12229), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11786) );
  AOI22_X1 U14779 ( .A1(n11987), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12285), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11785) );
  AOI22_X1 U14780 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11784) );
  INV_X1 U14781 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n20276) );
  AOI22_X1 U14782 ( .A1(n12129), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12112), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11783) );
  NAND4_X1 U14783 ( .A1(n11786), .A2(n11785), .A3(n11784), .A4(n11783), .ZN(
        n11787) );
  NAND2_X1 U14784 ( .A1(n12334), .A2(n13345), .ZN(n11790) );
  NAND2_X1 U14785 ( .A1(n12355), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11789) );
  NAND2_X1 U14786 ( .A1(n11790), .A2(n11789), .ZN(n11858) );
  AOI22_X1 U14787 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12134), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11794) );
  AOI22_X1 U14788 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12129), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11793) );
  AOI22_X1 U14789 ( .A1(n11987), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12229), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11792) );
  AOI22_X1 U14790 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11791) );
  NAND4_X1 U14791 ( .A1(n11794), .A2(n11793), .A3(n11792), .A4(n11791), .ZN(
        n11800) );
  AOI22_X1 U14792 ( .A1(n12230), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11798) );
  AOI22_X1 U14793 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11797) );
  AOI22_X1 U14794 ( .A1(n12284), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11796) );
  AOI22_X1 U14795 ( .A1(n12135), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12112), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11795) );
  NAND4_X1 U14796 ( .A1(n11798), .A2(n11797), .A3(n11796), .A4(n11795), .ZN(
        n11799) );
  AOI22_X1 U14797 ( .A1(n12334), .A2(n13485), .B1(n12355), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11864) );
  INV_X1 U14798 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n20295) );
  INV_X1 U14799 ( .A(n12355), .ZN(n12351) );
  NAND2_X1 U14800 ( .A1(n12334), .A2(n13487), .ZN(n11801) );
  OAI21_X1 U14801 ( .B1(n20295), .B2(n12351), .A(n11801), .ZN(n11802) );
  INV_X1 U14802 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n13292) );
  NAND2_X1 U14803 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11813) );
  INV_X1 U14804 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11803) );
  INV_X1 U14805 ( .A(n11888), .ZN(n11806) );
  INV_X1 U14806 ( .A(n11804), .ZN(n11869) );
  INV_X1 U14807 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16042) );
  NAND2_X1 U14808 ( .A1(n11869), .A2(n16042), .ZN(n11805) );
  NAND2_X1 U14809 ( .A1(n11806), .A2(n11805), .ZN(n20025) );
  AOI22_X1 U14810 ( .A1(n20025), .A2(n12307), .B1(n12314), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11807) );
  OAI21_X1 U14811 ( .B1(n11978), .B2(n13292), .A(n11807), .ZN(n11808) );
  AOI21_X1 U14812 ( .B1(n13483), .B2(n11996), .A(n11808), .ZN(n13290) );
  INV_X1 U14813 ( .A(n13121), .ZN(n13123) );
  NAND2_X1 U14814 ( .A1(n11809), .A2(n13123), .ZN(n11810) );
  NAND2_X1 U14815 ( .A1(n11810), .A2(n11850), .ZN(n13063) );
  OR2_X1 U14816 ( .A1(n13063), .A2(n10300), .ZN(n11820) );
  OR2_X1 U14817 ( .A1(n12763), .A2(n20898), .ZN(n11854) );
  NAND2_X1 U14818 ( .A1(n12308), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11817) );
  INV_X1 U14819 ( .A(n11813), .ZN(n11815) );
  INV_X1 U14820 ( .A(n11851), .ZN(n11814) );
  OAI21_X1 U14821 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11815), .A(
        n11814), .ZN(n14260) );
  AOI22_X1 U14822 ( .A1(n12307), .A2(n14260), .B1(n12314), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11816) );
  OAI211_X1 U14823 ( .C1(n11854), .C2(n11811), .A(n11817), .B(n11816), .ZN(
        n11818) );
  INV_X1 U14824 ( .A(n11818), .ZN(n11819) );
  NAND2_X1 U14825 ( .A1(n11812), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11824) );
  XNOR2_X1 U14826 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14269) );
  AOI21_X1 U14827 ( .B1(n11844), .B2(n14269), .A(n12314), .ZN(n11823) );
  OAI211_X1 U14828 ( .C1(n11854), .C2(n12859), .A(n11824), .B(n11823), .ZN(
        n11825) );
  INV_X1 U14829 ( .A(n11825), .ZN(n11826) );
  NAND2_X1 U14830 ( .A1(n12314), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11848) );
  NAND2_X1 U14831 ( .A1(n11827), .A2(n12810), .ZN(n11828) );
  NAND2_X1 U14832 ( .A1(n20766), .A2(n11996), .ZN(n11834) );
  NAND2_X1 U14833 ( .A1(n11812), .A2(P1_EAX_REG_1__SCAN_IN), .ZN(n11831) );
  NAND2_X1 U14834 ( .A1(n20898), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11830) );
  OAI211_X1 U14835 ( .C1(n11854), .C2(n11710), .A(n11831), .B(n11830), .ZN(
        n11832) );
  INV_X1 U14836 ( .A(n11832), .ZN(n11833) );
  NAND2_X1 U14837 ( .A1(n11834), .A2(n11833), .ZN(n12805) );
  NAND2_X1 U14838 ( .A1(n20323), .A2(n20278), .ZN(n11837) );
  NAND2_X1 U14839 ( .A1(n11837), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12730) );
  NAND2_X1 U14840 ( .A1(n11812), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11841) );
  NAND2_X1 U14841 ( .A1(n20898), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11840) );
  OAI211_X1 U14842 ( .C1(n11854), .C2(n12844), .A(n11841), .B(n11840), .ZN(
        n11842) );
  AOI21_X1 U14843 ( .B1(n11839), .B2(n11996), .A(n11842), .ZN(n11843) );
  OR2_X1 U14844 ( .A1(n12730), .A2(n11843), .ZN(n12731) );
  INV_X1 U14845 ( .A(n11843), .ZN(n12732) );
  OR2_X1 U14846 ( .A1(n12732), .A2(n13425), .ZN(n11845) );
  NAND2_X1 U14847 ( .A1(n12731), .A2(n11845), .ZN(n12804) );
  NAND2_X1 U14848 ( .A1(n12805), .A2(n12804), .ZN(n12930) );
  NAND2_X1 U14849 ( .A1(n11847), .A2(n11846), .ZN(n12928) );
  XNOR2_X1 U14850 ( .A(n11850), .B(n11849), .ZN(n13328) );
  NAND2_X1 U14851 ( .A1(n13328), .A2(n11996), .ZN(n11857) );
  OAI21_X1 U14852 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n11851), .A(
        n11859), .ZN(n20163) );
  INV_X1 U14853 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16184) );
  NAND2_X1 U14854 ( .A1(n12308), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11853) );
  INV_X1 U14855 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21280) );
  OAI21_X1 U14856 ( .B1(n21280), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20898), .ZN(n11852) );
  OAI211_X1 U14857 ( .C1(n11854), .C2(n16184), .A(n11853), .B(n11852), .ZN(
        n11855) );
  OAI21_X1 U14858 ( .B1(n13425), .B2(n20163), .A(n11855), .ZN(n11856) );
  INV_X1 U14859 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n13137) );
  INV_X1 U14860 ( .A(n11859), .ZN(n11861) );
  INV_X1 U14861 ( .A(n11860), .ZN(n11866) );
  OAI21_X1 U14862 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n11861), .A(
        n11866), .ZN(n20044) );
  AOI22_X1 U14863 ( .A1(n12307), .A2(n20044), .B1(n12314), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11862) );
  OAI21_X1 U14864 ( .B1(n11978), .B2(n13137), .A(n11862), .ZN(n11863) );
  AOI21_X1 U14865 ( .B1(n13335), .B2(n11996), .A(n11863), .ZN(n13135) );
  INV_X1 U14866 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n20122) );
  NAND2_X1 U14867 ( .A1(n11865), .A2(n11864), .ZN(n13343) );
  NAND2_X1 U14868 ( .A1(n13343), .A2(n11996), .ZN(n11871) );
  INV_X1 U14869 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11867) );
  NAND2_X1 U14870 ( .A1(n11867), .A2(n11866), .ZN(n11868) );
  NAND2_X1 U14871 ( .A1(n11869), .A2(n11868), .ZN(n20035) );
  AOI22_X1 U14872 ( .A1(n20035), .A2(n12307), .B1(n12314), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11870) );
  NAND2_X1 U14873 ( .A1(n13134), .A2(n13164), .ZN(n13162) );
  INV_X1 U14874 ( .A(n13162), .ZN(n11872) );
  AOI22_X1 U14875 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12129), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11877) );
  AOI22_X1 U14876 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11876) );
  AOI22_X1 U14877 ( .A1(n11987), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12229), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11875) );
  AOI22_X1 U14878 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11874) );
  NAND4_X1 U14879 ( .A1(n11877), .A2(n11876), .A3(n11875), .A4(n11874), .ZN(
        n11883) );
  AOI22_X1 U14880 ( .A1(n12230), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11881) );
  AOI22_X1 U14881 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11880) );
  AOI22_X1 U14882 ( .A1(n12284), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11879) );
  AOI22_X1 U14883 ( .A1(n12042), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12112), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11878) );
  NAND4_X1 U14884 ( .A1(n11881), .A2(n11880), .A3(n11879), .A4(n11878), .ZN(
        n11882) );
  OAI21_X1 U14885 ( .B1(n11883), .B2(n11882), .A(n11996), .ZN(n11886) );
  XNOR2_X1 U14886 ( .A(n11888), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13517) );
  AOI22_X1 U14887 ( .A1(n13517), .A2(n12307), .B1(n12314), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11885) );
  NAND2_X1 U14888 ( .A1(n12308), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11884) );
  XOR2_X1 U14889 ( .A(n20006), .B(n11914), .Z(n20009) );
  INV_X1 U14890 ( .A(n20009), .ZN(n11903) );
  AOI22_X1 U14891 ( .A1(n11987), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11892) );
  AOI22_X1 U14892 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U14893 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11890) );
  AOI22_X1 U14894 ( .A1(n12129), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11889) );
  NAND4_X1 U14895 ( .A1(n11892), .A2(n11891), .A3(n11890), .A4(n11889), .ZN(
        n11898) );
  AOI22_X1 U14896 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11896) );
  AOI22_X1 U14897 ( .A1(n12042), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11895) );
  AOI22_X1 U14898 ( .A1(n11561), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12112), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11894) );
  AOI22_X1 U14899 ( .A1(n12230), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11893) );
  NAND4_X1 U14900 ( .A1(n11896), .A2(n11895), .A3(n11894), .A4(n11893), .ZN(
        n11897) );
  OAI21_X1 U14901 ( .B1(n11898), .B2(n11897), .A(n11996), .ZN(n11901) );
  NAND2_X1 U14902 ( .A1(n12308), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11900) );
  NAND2_X1 U14903 ( .A1(n12314), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11899) );
  NAND3_X1 U14904 ( .A1(n11901), .A2(n11900), .A3(n11899), .ZN(n11902) );
  AOI21_X1 U14905 ( .B1(n11903), .B2(n12307), .A(n11902), .ZN(n13475) );
  AOI22_X1 U14906 ( .A1(n11987), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12286), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11907) );
  AOI22_X1 U14907 ( .A1(n12230), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12134), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11906) );
  AOI22_X1 U14908 ( .A1(n12284), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11905) );
  AOI22_X1 U14909 ( .A1(n12129), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12112), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11904) );
  NAND4_X1 U14910 ( .A1(n11907), .A2(n11906), .A3(n11905), .A4(n11904), .ZN(
        n11913) );
  AOI22_X1 U14911 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11911) );
  AOI22_X1 U14912 ( .A1(n12106), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11910) );
  AOI22_X1 U14913 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11909) );
  AOI22_X1 U14914 ( .A1(n11561), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11908) );
  NAND4_X1 U14915 ( .A1(n11911), .A2(n11910), .A3(n11909), .A4(n11908), .ZN(
        n11912) );
  NOR2_X1 U14916 ( .A1(n11913), .A2(n11912), .ZN(n11917) );
  XNOR2_X1 U14917 ( .A(n11918), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14572) );
  NAND2_X1 U14918 ( .A1(n14572), .A2(n12307), .ZN(n11916) );
  AOI22_X1 U14919 ( .A1(n12308), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n12314), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11915) );
  OAI211_X1 U14920 ( .C1(n11917), .C2(n10300), .A(n11916), .B(n11915), .ZN(
        n13559) );
  AND2_X2 U14921 ( .A1(n13476), .A2(n13559), .ZN(n13560) );
  NAND2_X1 U14922 ( .A1(n12308), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n11921) );
  OAI21_X1 U14923 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11919), .A(
        n11962), .ZN(n16032) );
  AOI22_X1 U14924 ( .A1(n12307), .A2(n16032), .B1(n12314), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11920) );
  NAND2_X1 U14925 ( .A1(n11921), .A2(n11920), .ZN(n14238) );
  AOI22_X1 U14926 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11925) );
  AOI22_X1 U14927 ( .A1(n12106), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12230), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11924) );
  AOI22_X1 U14928 ( .A1(n12042), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11923) );
  AOI22_X1 U14929 ( .A1(n11987), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12112), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11922) );
  NAND4_X1 U14930 ( .A1(n11925), .A2(n11924), .A3(n11923), .A4(n11922), .ZN(
        n11932) );
  AOI22_X1 U14931 ( .A1(n12129), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11930) );
  AOI22_X1 U14932 ( .A1(n12296), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12229), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11929) );
  AOI22_X1 U14933 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11928) );
  AOI22_X1 U14934 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11927) );
  NAND4_X1 U14935 ( .A1(n11930), .A2(n11929), .A3(n11928), .A4(n11927), .ZN(
        n11931) );
  OR2_X1 U14936 ( .A1(n11932), .A2(n11931), .ZN(n11933) );
  AOI22_X1 U14937 ( .A1(n12129), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11937) );
  AOI22_X1 U14938 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n12230), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11936) );
  AOI22_X1 U14939 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11935) );
  AOI22_X1 U14940 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12042), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11934) );
  NAND4_X1 U14941 ( .A1(n11937), .A2(n11936), .A3(n11935), .A4(n11934), .ZN(
        n11945) );
  AOI22_X1 U14942 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12106), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11943) );
  AOI22_X1 U14943 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12229), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11942) );
  AOI22_X1 U14944 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11987), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11941) );
  AOI22_X1 U14945 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12112), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11940) );
  NAND4_X1 U14946 ( .A1(n11943), .A2(n11942), .A3(n11941), .A4(n11940), .ZN(
        n11944) );
  NOR2_X1 U14947 ( .A1(n11945), .A2(n11944), .ZN(n11949) );
  XNOR2_X1 U14948 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n11962), .ZN(
        n16020) );
  INV_X1 U14949 ( .A(n12314), .ZN(n12034) );
  OAI22_X1 U14950 ( .A1(n16020), .A2(n13425), .B1(n12034), .B2(n11961), .ZN(
        n11946) );
  INV_X1 U14951 ( .A(n11946), .ZN(n11948) );
  NAND2_X1 U14952 ( .A1(n12308), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n11947) );
  OAI211_X1 U14953 ( .C1(n10300), .C2(n11949), .A(n11948), .B(n11947), .ZN(
        n14324) );
  AOI22_X1 U14954 ( .A1(n12042), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11953) );
  AOI22_X1 U14955 ( .A1(n12106), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11952) );
  AOI22_X1 U14956 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11951) );
  AOI22_X1 U14957 ( .A1(n12129), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11950) );
  NAND4_X1 U14958 ( .A1(n11953), .A2(n11952), .A3(n11951), .A4(n11950), .ZN(
        n11960) );
  AOI22_X1 U14959 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11958) );
  AOI22_X1 U14960 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12229), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11957) );
  AOI22_X1 U14961 ( .A1(n12230), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11956) );
  AOI22_X1 U14962 ( .A1(n11987), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12112), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11955) );
  NAND4_X1 U14963 ( .A1(n11958), .A2(n11957), .A3(n11956), .A4(n11955), .ZN(
        n11959) );
  NOR2_X1 U14964 ( .A1(n11960), .A2(n11959), .ZN(n11965) );
  XNOR2_X1 U14965 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n11967), .ZN(
        n14559) );
  AOI22_X1 U14966 ( .A1(n12307), .A2(n14559), .B1(n12314), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11964) );
  NAND2_X1 U14967 ( .A1(n12308), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11963) );
  OAI211_X1 U14968 ( .C1(n10300), .C2(n11965), .A(n11964), .B(n11963), .ZN(
        n14240) );
  XOR2_X1 U14969 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n11986), .Z(
        n16015) );
  INV_X1 U14970 ( .A(n16015), .ZN(n11983) );
  AOI22_X1 U14971 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12134), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11971) );
  AOI22_X1 U14972 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11970) );
  AOI22_X1 U14973 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11969) );
  AOI22_X1 U14974 ( .A1(n12129), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11968) );
  NAND4_X1 U14975 ( .A1(n11971), .A2(n11970), .A3(n11969), .A4(n11968), .ZN(
        n11977) );
  AOI22_X1 U14976 ( .A1(n12284), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11975) );
  AOI22_X1 U14977 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12229), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11974) );
  AOI22_X1 U14978 ( .A1(n12230), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11973) );
  AOI22_X1 U14979 ( .A1(n11987), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12112), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11972) );
  NAND4_X1 U14980 ( .A1(n11975), .A2(n11974), .A3(n11973), .A4(n11972), .ZN(
        n11976) );
  OAI21_X1 U14981 ( .B1(n11977), .B2(n11976), .A(n11996), .ZN(n11981) );
  NAND2_X1 U14982 ( .A1(n12308), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11980) );
  NAND2_X1 U14983 ( .A1(n12314), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11979) );
  NAND3_X1 U14984 ( .A1(n11981), .A2(n11980), .A3(n11979), .ZN(n11982) );
  AOI21_X1 U14985 ( .B1(n11983), .B2(n12307), .A(n11982), .ZN(n14227) );
  NAND2_X1 U14986 ( .A1(n11985), .A2(n11984), .ZN(n14212) );
  INV_X1 U14987 ( .A(n14212), .ZN(n12003) );
  XNOR2_X1 U14988 ( .A(n12019), .B(n12018), .ZN(n14547) );
  AOI22_X1 U14989 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12134), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11991) );
  AOI22_X1 U14990 ( .A1(n11987), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12129), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11990) );
  AOI22_X1 U14991 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12128), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11989) );
  AOI22_X1 U14992 ( .A1(n11561), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11988) );
  NAND4_X1 U14993 ( .A1(n11991), .A2(n11990), .A3(n11989), .A4(n11988), .ZN(
        n11998) );
  AOI22_X1 U14994 ( .A1(n12284), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11995) );
  AOI22_X1 U14995 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11994) );
  AOI22_X1 U14996 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13091), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11993) );
  AOI22_X1 U14997 ( .A1(n12230), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11992) );
  NAND4_X1 U14998 ( .A1(n11995), .A2(n11994), .A3(n11993), .A4(n11992), .ZN(
        n11997) );
  OAI21_X1 U14999 ( .B1(n11998), .B2(n11997), .A(n11996), .ZN(n12000) );
  NAND2_X1 U15000 ( .A1(n12308), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11999) );
  OAI211_X1 U15001 ( .C1(n12034), .C2(n12018), .A(n12000), .B(n11999), .ZN(
        n12001) );
  AOI21_X1 U15002 ( .B1(n14547), .B2(n12307), .A(n12001), .ZN(n14214) );
  NAND2_X1 U15003 ( .A1(n12003), .A2(n12002), .ZN(n14213) );
  AOI22_X1 U15004 ( .A1(n12042), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12129), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12007) );
  AOI22_X1 U15005 ( .A1(n12135), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12006) );
  AOI22_X1 U15006 ( .A1(n11987), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12229), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12005) );
  AOI22_X1 U15007 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12128), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12004) );
  NAND4_X1 U15008 ( .A1(n12007), .A2(n12006), .A3(n12005), .A4(n12004), .ZN(
        n12013) );
  AOI22_X1 U15009 ( .A1(n12106), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12230), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12011) );
  AOI22_X1 U15010 ( .A1(n12284), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12010) );
  AOI22_X1 U15011 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12009) );
  AOI22_X1 U15012 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12112), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12008) );
  NAND4_X1 U15013 ( .A1(n12011), .A2(n12010), .A3(n12009), .A4(n12008), .ZN(
        n12012) );
  NOR2_X1 U15014 ( .A1(n12013), .A2(n12012), .ZN(n12017) );
  NAND2_X1 U15015 ( .A1(n20898), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12014) );
  NAND2_X1 U15016 ( .A1(n13425), .A2(n12014), .ZN(n12015) );
  AOI21_X1 U15017 ( .B1(n12308), .B2(P1_EAX_REG_16__SCAN_IN), .A(n12015), .ZN(
        n12016) );
  OAI21_X1 U15018 ( .B1(n12311), .B2(n12017), .A(n12016), .ZN(n12022) );
  OAI21_X1 U15019 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12020), .A(
        n12053), .ZN(n16007) );
  OR2_X1 U15020 ( .A1(n13425), .A2(n16007), .ZN(n12021) );
  NAND2_X1 U15021 ( .A1(n12022), .A2(n12021), .ZN(n14307) );
  AOI22_X1 U15022 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12134), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12026) );
  AOI22_X1 U15023 ( .A1(n12135), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12025) );
  AOI22_X1 U15024 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12128), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12024) );
  AOI22_X1 U15025 ( .A1(n11561), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12023) );
  NAND4_X1 U15026 ( .A1(n12026), .A2(n12025), .A3(n12024), .A4(n12023), .ZN(
        n12032) );
  AOI22_X1 U15027 ( .A1(n11987), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12286), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12030) );
  AOI22_X1 U15028 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12029) );
  AOI22_X1 U15029 ( .A1(n12230), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12028) );
  AOI22_X1 U15030 ( .A1(n12129), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13091), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12027) );
  NAND4_X1 U15031 ( .A1(n12030), .A2(n12029), .A3(n12028), .A4(n12027), .ZN(
        n12031) );
  OR2_X1 U15032 ( .A1(n12032), .A2(n12031), .ZN(n12033) );
  NAND2_X1 U15033 ( .A1(n12277), .A2(n12033), .ZN(n12037) );
  XNOR2_X1 U15034 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n12053), .ZN(
        n14537) );
  OAI22_X1 U15035 ( .A1(n13425), .A2(n14537), .B1(n12034), .B2(n14533), .ZN(
        n12035) );
  AOI21_X1 U15036 ( .B1(n12308), .B2(P1_EAX_REG_17__SCAN_IN), .A(n12035), .ZN(
        n12036) );
  NAND2_X1 U15037 ( .A1(n12037), .A2(n12036), .ZN(n14200) );
  AOI22_X1 U15038 ( .A1(n11987), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12041) );
  AOI22_X1 U15039 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12040) );
  AOI22_X1 U15040 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12128), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12039) );
  AOI22_X1 U15041 ( .A1(n12129), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12285), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12038) );
  NAND4_X1 U15042 ( .A1(n12041), .A2(n12040), .A3(n12039), .A4(n12038), .ZN(
        n12048) );
  AOI22_X1 U15043 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12046) );
  AOI22_X1 U15044 ( .A1(n12042), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12045) );
  AOI22_X1 U15045 ( .A1(n11561), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13091), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12044) );
  AOI22_X1 U15046 ( .A1(n12230), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12043) );
  NAND4_X1 U15047 ( .A1(n12046), .A2(n12045), .A3(n12044), .A4(n12043), .ZN(
        n12047) );
  NOR2_X1 U15048 ( .A1(n12048), .A2(n12047), .ZN(n12052) );
  NAND2_X1 U15049 ( .A1(n20898), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12049) );
  NAND2_X1 U15050 ( .A1(n13425), .A2(n12049), .ZN(n12050) );
  AOI21_X1 U15051 ( .B1(n12308), .B2(P1_EAX_REG_18__SCAN_IN), .A(n12050), .ZN(
        n12051) );
  OAI21_X1 U15052 ( .B1(n12311), .B2(n12052), .A(n12051), .ZN(n12056) );
  OAI21_X1 U15053 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n12054), .A(
        n12086), .ZN(n15948) );
  OR2_X1 U15054 ( .A1(n13425), .A2(n15948), .ZN(n12055) );
  NAND2_X1 U15055 ( .A1(n12056), .A2(n12055), .ZN(n14296) );
  AOI22_X1 U15056 ( .A1(n11987), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12129), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12060) );
  AOI22_X1 U15057 ( .A1(n12042), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12059) );
  AOI22_X1 U15058 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12128), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12058) );
  AOI22_X1 U15059 ( .A1(n11561), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12285), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12057) );
  NAND4_X1 U15060 ( .A1(n12060), .A2(n12059), .A3(n12058), .A4(n12057), .ZN(
        n12066) );
  AOI22_X1 U15061 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12064) );
  AOI22_X1 U15062 ( .A1(n12230), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12063) );
  AOI22_X1 U15063 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13091), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12062) );
  AOI22_X1 U15064 ( .A1(n12284), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12061) );
  NAND4_X1 U15065 ( .A1(n12064), .A2(n12063), .A3(n12062), .A4(n12061), .ZN(
        n12065) );
  NOR2_X1 U15066 ( .A1(n12066), .A2(n12065), .ZN(n12069) );
  OAI21_X1 U15067 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14513), .A(n13425), 
        .ZN(n12067) );
  AOI21_X1 U15068 ( .B1(n12308), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12067), .ZN(
        n12068) );
  OAI21_X1 U15069 ( .B1(n12311), .B2(n12069), .A(n12068), .ZN(n12071) );
  XNOR2_X1 U15070 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n12086), .ZN(
        n14517) );
  NAND2_X1 U15071 ( .A1(n12307), .A2(n14517), .ZN(n12070) );
  NAND2_X1 U15072 ( .A1(n12071), .A2(n12070), .ZN(n14288) );
  AOI22_X1 U15073 ( .A1(n11987), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12075) );
  AOI22_X1 U15074 ( .A1(n12230), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12074) );
  AOI22_X1 U15075 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12128), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12073) );
  AOI22_X1 U15076 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n11939), .B1(
        n12285), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12072) );
  NAND4_X1 U15077 ( .A1(n12075), .A2(n12074), .A3(n12073), .A4(n12072), .ZN(
        n12081) );
  AOI22_X1 U15078 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n12284), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12079) );
  AOI22_X1 U15079 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12229), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12078) );
  AOI22_X1 U15080 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12129), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12077) );
  AOI22_X1 U15081 ( .A1(n12042), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13091), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12076) );
  NAND4_X1 U15082 ( .A1(n12079), .A2(n12078), .A3(n12077), .A4(n12076), .ZN(
        n12080) );
  NOR2_X1 U15083 ( .A1(n12081), .A2(n12080), .ZN(n12085) );
  NAND2_X1 U15084 ( .A1(n20898), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12082) );
  NAND2_X1 U15085 ( .A1(n13425), .A2(n12082), .ZN(n12083) );
  AOI21_X1 U15086 ( .B1(n12308), .B2(P1_EAX_REG_20__SCAN_IN), .A(n12083), .ZN(
        n12084) );
  OAI21_X1 U15087 ( .B1(n12311), .B2(n12085), .A(n12084), .ZN(n12089) );
  OAI21_X1 U15088 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12087), .A(
        n12124), .ZN(n15996) );
  OR2_X1 U15089 ( .A1(n13425), .A2(n15996), .ZN(n12088) );
  NAND2_X1 U15090 ( .A1(n12089), .A2(n12088), .ZN(n14287) );
  NOR2_X2 U15091 ( .A1(n14188), .A2(n12090), .ZN(n14286) );
  AOI22_X1 U15092 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12129), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12094) );
  AOI22_X1 U15093 ( .A1(n12134), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12093) );
  AOI22_X1 U15094 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12229), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12092) );
  AOI22_X1 U15095 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12128), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12091) );
  NAND4_X1 U15096 ( .A1(n12094), .A2(n12093), .A3(n12092), .A4(n12091), .ZN(
        n12100) );
  AOI22_X1 U15097 ( .A1(n11938), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12098) );
  AOI22_X1 U15098 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12285), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12097) );
  AOI22_X1 U15099 ( .A1(n12230), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12096) );
  AOI22_X1 U15100 ( .A1(n12244), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13091), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12095) );
  NAND4_X1 U15101 ( .A1(n12098), .A2(n12097), .A3(n12096), .A4(n12095), .ZN(
        n12099) );
  NOR2_X1 U15102 ( .A1(n12100), .A2(n12099), .ZN(n12103) );
  INV_X1 U15103 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12123) );
  OAI21_X1 U15104 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n12123), .A(n13425), 
        .ZN(n12101) );
  AOI21_X1 U15105 ( .B1(n12308), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12101), .ZN(
        n12102) );
  OAI21_X1 U15106 ( .B1(n12311), .B2(n12103), .A(n12102), .ZN(n12105) );
  XNOR2_X1 U15107 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n12124), .ZN(
        n15991) );
  NAND2_X1 U15108 ( .A1(n15991), .A2(n12307), .ZN(n12104) );
  AND2_X2 U15109 ( .A1(n14286), .A2(n14361), .ZN(n14357) );
  AOI22_X1 U15110 ( .A1(n11938), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12110) );
  AOI22_X1 U15111 ( .A1(n12230), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12134), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12109) );
  AOI22_X1 U15112 ( .A1(n11926), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12108) );
  AOI22_X1 U15113 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12229), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12107) );
  NAND4_X1 U15114 ( .A1(n12110), .A2(n12109), .A3(n12108), .A4(n12107), .ZN(
        n12118) );
  AOI22_X1 U15115 ( .A1(n12129), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12116) );
  AOI22_X1 U15116 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12115) );
  AOI22_X1 U15117 ( .A1(n12284), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12114) );
  AOI22_X1 U15118 ( .A1(n12244), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12112), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12113) );
  NAND4_X1 U15119 ( .A1(n12116), .A2(n12115), .A3(n12114), .A4(n12113), .ZN(
        n12117) );
  NOR2_X1 U15120 ( .A1(n12118), .A2(n12117), .ZN(n12122) );
  NAND2_X1 U15121 ( .A1(n20898), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12119) );
  NAND2_X1 U15122 ( .A1(n13425), .A2(n12119), .ZN(n12120) );
  AOI21_X1 U15123 ( .B1(n12308), .B2(P1_EAX_REG_22__SCAN_IN), .A(n12120), .ZN(
        n12121) );
  OAI21_X1 U15124 ( .B1(n12311), .B2(n12122), .A(n12121), .ZN(n12127) );
  OAI21_X1 U15125 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n12125), .A(
        n12177), .ZN(n15990) );
  OR2_X1 U15126 ( .A1(n13425), .A2(n15990), .ZN(n12126) );
  AOI22_X1 U15127 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12229), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12133) );
  AOI22_X1 U15128 ( .A1(n11987), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12285), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12132) );
  AOI22_X1 U15129 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12128), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12131) );
  AOI22_X1 U15130 ( .A1(n12129), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13091), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12130) );
  NAND4_X1 U15131 ( .A1(n12133), .A2(n12132), .A3(n12131), .A4(n12130), .ZN(
        n12141) );
  AOI22_X1 U15132 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12134), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12139) );
  AOI22_X1 U15133 ( .A1(n12106), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12138) );
  AOI22_X1 U15134 ( .A1(n12284), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12137) );
  AOI22_X1 U15135 ( .A1(n12230), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12136) );
  NAND4_X1 U15136 ( .A1(n12139), .A2(n12138), .A3(n12137), .A4(n12136), .ZN(
        n12140) );
  NOR2_X1 U15137 ( .A1(n12141), .A2(n12140), .ZN(n12161) );
  AOI22_X1 U15138 ( .A1(n12284), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12145) );
  AOI22_X1 U15139 ( .A1(n12249), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12144) );
  AOI22_X1 U15140 ( .A1(n11561), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12143) );
  AOI22_X1 U15141 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12112), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12142) );
  NAND4_X1 U15142 ( .A1(n12145), .A2(n12144), .A3(n12143), .A4(n12142), .ZN(
        n12153) );
  AOI22_X1 U15143 ( .A1(n12042), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12129), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12151) );
  AOI22_X1 U15144 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12150) );
  AOI22_X1 U15145 ( .A1(n11987), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12149) );
  AOI22_X1 U15146 ( .A1(n11578), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12148) );
  NAND4_X1 U15147 ( .A1(n12151), .A2(n12150), .A3(n12149), .A4(n12148), .ZN(
        n12152) );
  NOR2_X1 U15148 ( .A1(n12153), .A2(n12152), .ZN(n12162) );
  XOR2_X1 U15149 ( .A(n12161), .B(n12162), .Z(n12154) );
  NAND2_X1 U15150 ( .A1(n12154), .A2(n12277), .ZN(n12158) );
  NAND2_X1 U15151 ( .A1(n20898), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12155) );
  NAND2_X1 U15152 ( .A1(n13425), .A2(n12155), .ZN(n12156) );
  AOI21_X1 U15153 ( .B1(n12308), .B2(P1_EAX_REG_23__SCAN_IN), .A(n12156), .ZN(
        n12157) );
  NAND2_X1 U15154 ( .A1(n12158), .A2(n12157), .ZN(n12160) );
  XNOR2_X1 U15155 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B(n12177), .ZN(
        n14503) );
  NAND2_X1 U15156 ( .A1(n12307), .A2(n14503), .ZN(n12159) );
  NAND2_X1 U15157 ( .A1(n12160), .A2(n12159), .ZN(n14176) );
  NOR2_X1 U15158 ( .A1(n12162), .A2(n12161), .ZN(n12185) );
  AOI22_X1 U15159 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12166) );
  AOI22_X1 U15160 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12165) );
  AOI22_X1 U15161 ( .A1(n12284), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12164) );
  INV_X1 U15162 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n20246) );
  AOI22_X1 U15163 ( .A1(n12230), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12163) );
  NAND4_X1 U15164 ( .A1(n12166), .A2(n12165), .A3(n12164), .A4(n12163), .ZN(
        n12172) );
  AOI22_X1 U15165 ( .A1(n12249), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12229), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12170) );
  AOI22_X1 U15166 ( .A1(n11987), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12169) );
  AOI22_X1 U15167 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12168) );
  AOI22_X1 U15168 ( .A1(n11607), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12112), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12167) );
  NAND4_X1 U15169 ( .A1(n12170), .A2(n12169), .A3(n12168), .A4(n12167), .ZN(
        n12171) );
  OR2_X1 U15170 ( .A1(n12172), .A2(n12171), .ZN(n12184) );
  XNOR2_X1 U15171 ( .A(n12185), .B(n12184), .ZN(n12176) );
  NAND2_X1 U15172 ( .A1(n20898), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12173) );
  NAND2_X1 U15173 ( .A1(n13425), .A2(n12173), .ZN(n12174) );
  AOI21_X1 U15174 ( .B1(n12308), .B2(P1_EAX_REG_24__SCAN_IN), .A(n12174), .ZN(
        n12175) );
  OAI21_X1 U15175 ( .B1(n12176), .B2(n12311), .A(n12175), .ZN(n12183) );
  INV_X1 U15176 ( .A(n12179), .ZN(n12180) );
  INV_X1 U15177 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14495) );
  NAND2_X1 U15178 ( .A1(n12180), .A2(n14495), .ZN(n12181) );
  AND2_X1 U15179 ( .A1(n12201), .A2(n12181), .ZN(n14497) );
  NAND2_X1 U15180 ( .A1(n14497), .A2(n12307), .ZN(n12182) );
  NAND2_X1 U15181 ( .A1(n12183), .A2(n12182), .ZN(n14161) );
  NAND2_X1 U15182 ( .A1(n12185), .A2(n12184), .ZN(n12206) );
  AOI22_X1 U15183 ( .A1(n11987), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12286), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12189) );
  AOI22_X1 U15184 ( .A1(n12244), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12188) );
  AOI22_X1 U15185 ( .A1(n11607), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12187) );
  AOI22_X1 U15186 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12112), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12186) );
  NAND4_X1 U15187 ( .A1(n12189), .A2(n12188), .A3(n12187), .A4(n12186), .ZN(
        n12195) );
  AOI22_X1 U15188 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12193) );
  AOI22_X1 U15189 ( .A1(n12042), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12229), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12192) );
  AOI22_X1 U15190 ( .A1(n12230), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12191) );
  AOI22_X1 U15191 ( .A1(n12285), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12190) );
  NAND4_X1 U15192 ( .A1(n12193), .A2(n12192), .A3(n12191), .A4(n12190), .ZN(
        n12194) );
  NOR2_X1 U15193 ( .A1(n12195), .A2(n12194), .ZN(n12207) );
  XOR2_X1 U15194 ( .A(n12206), .B(n12207), .Z(n12196) );
  NAND2_X1 U15195 ( .A1(n12196), .A2(n12277), .ZN(n12200) );
  INV_X1 U15196 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14485) );
  AOI21_X1 U15197 ( .B1(n14485), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12197) );
  AOI21_X1 U15198 ( .B1(n12308), .B2(P1_EAX_REG_25__SCAN_IN), .A(n12197), .ZN(
        n12199) );
  XNOR2_X1 U15199 ( .A(n12201), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14487) );
  AOI21_X1 U15200 ( .B1(n12200), .B2(n12199), .A(n12198), .ZN(n14150) );
  INV_X1 U15201 ( .A(n12202), .ZN(n12204) );
  INV_X1 U15202 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12203) );
  NAND2_X1 U15203 ( .A1(n12204), .A2(n12203), .ZN(n12205) );
  NAND2_X1 U15204 ( .A1(n12258), .A2(n12205), .ZN(n14475) );
  NOR2_X1 U15205 ( .A1(n12207), .A2(n12206), .ZN(n12223) );
  AOI22_X1 U15206 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12211) );
  AOI22_X1 U15207 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12244), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12210) );
  AOI22_X1 U15208 ( .A1(n12284), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12209) );
  AOI22_X1 U15209 ( .A1(n12230), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12208) );
  NAND4_X1 U15210 ( .A1(n12211), .A2(n12210), .A3(n12209), .A4(n12208), .ZN(
        n12217) );
  AOI22_X1 U15211 ( .A1(n12249), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12229), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12215) );
  AOI22_X1 U15212 ( .A1(n11987), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12214) );
  AOI22_X1 U15213 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12213) );
  AOI22_X1 U15214 ( .A1(n11607), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12112), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12212) );
  NAND4_X1 U15215 ( .A1(n12215), .A2(n12214), .A3(n12213), .A4(n12212), .ZN(
        n12216) );
  OR2_X1 U15216 ( .A1(n12217), .A2(n12216), .ZN(n12222) );
  XNOR2_X1 U15217 ( .A(n12223), .B(n12222), .ZN(n12220) );
  AOI21_X1 U15218 ( .B1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n20898), .A(
        n12307), .ZN(n12219) );
  NAND2_X1 U15219 ( .A1(n12308), .A2(P1_EAX_REG_26__SCAN_IN), .ZN(n12218) );
  OAI211_X1 U15220 ( .C1(n12220), .C2(n12311), .A(n12219), .B(n12218), .ZN(
        n12221) );
  OAI21_X1 U15221 ( .B1(n13425), .B2(n14475), .A(n12221), .ZN(n14136) );
  NOR2_X2 U15222 ( .A1(n14135), .A2(n14136), .ZN(n14120) );
  NAND2_X1 U15223 ( .A1(n12223), .A2(n12222), .ZN(n12241) );
  AOI22_X1 U15224 ( .A1(n11987), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12286), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12228) );
  AOI22_X1 U15225 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12227) );
  AOI22_X1 U15226 ( .A1(n11607), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12226) );
  AOI22_X1 U15227 ( .A1(n12134), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12112), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12225) );
  NAND4_X1 U15228 ( .A1(n12228), .A2(n12227), .A3(n12226), .A4(n12225), .ZN(
        n12236) );
  AOI22_X1 U15229 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12244), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12234) );
  AOI22_X1 U15230 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n12284), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12233) );
  AOI22_X1 U15231 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n11939), .B1(
        n12229), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12232) );
  AOI22_X1 U15232 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12230), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12231) );
  NAND4_X1 U15233 ( .A1(n12234), .A2(n12233), .A3(n12232), .A4(n12231), .ZN(
        n12235) );
  NOR2_X1 U15234 ( .A1(n12236), .A2(n12235), .ZN(n12242) );
  XOR2_X1 U15235 ( .A(n12241), .B(n12242), .Z(n12237) );
  NAND2_X1 U15236 ( .A1(n12237), .A2(n12277), .ZN(n12240) );
  INV_X1 U15237 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14462) );
  AOI21_X1 U15238 ( .B1(n14462), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12238) );
  AOI21_X1 U15239 ( .B1(n12308), .B2(P1_EAX_REG_27__SCAN_IN), .A(n12238), .ZN(
        n12239) );
  XNOR2_X1 U15240 ( .A(n12258), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14464) );
  AOI22_X1 U15241 ( .A1(n12240), .A2(n12239), .B1(n12307), .B2(n14464), .ZN(
        n14121) );
  NOR2_X1 U15242 ( .A1(n12242), .A2(n12241), .ZN(n12266) );
  AOI22_X1 U15243 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12248) );
  AOI22_X1 U15244 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12244), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12247) );
  AOI22_X1 U15245 ( .A1(n12284), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12246) );
  AOI22_X1 U15246 ( .A1(n11578), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12245) );
  NAND4_X1 U15247 ( .A1(n12248), .A2(n12247), .A3(n12246), .A4(n12245), .ZN(
        n12255) );
  AOI22_X1 U15248 ( .A1(n12249), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12229), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12253) );
  AOI22_X1 U15249 ( .A1(n11938), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12285), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12252) );
  AOI22_X1 U15250 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12251) );
  AOI22_X1 U15251 ( .A1(n11607), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13091), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12250) );
  NAND4_X1 U15252 ( .A1(n12253), .A2(n12252), .A3(n12251), .A4(n12250), .ZN(
        n12254) );
  OR2_X1 U15253 ( .A1(n12255), .A2(n12254), .ZN(n12265) );
  XNOR2_X1 U15254 ( .A(n12266), .B(n12265), .ZN(n12256) );
  NOR2_X1 U15255 ( .A1(n12256), .A2(n12311), .ZN(n12264) );
  INV_X1 U15256 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n21275) );
  NOR2_X1 U15257 ( .A1(n21280), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12257) );
  OAI22_X1 U15258 ( .A1(n11978), .A2(n21275), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n12257), .ZN(n12263) );
  INV_X1 U15259 ( .A(n12258), .ZN(n12259) );
  INV_X1 U15260 ( .A(n12260), .ZN(n12261) );
  INV_X1 U15261 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14111) );
  NAND2_X1 U15262 ( .A1(n12261), .A2(n14111), .ZN(n12262) );
  NAND2_X1 U15263 ( .A1(n12282), .A2(n12262), .ZN(n14458) );
  OAI22_X1 U15264 ( .A1(n12264), .A2(n12263), .B1(n13425), .B2(n14458), .ZN(
        n14110) );
  NAND2_X1 U15265 ( .A1(n12266), .A2(n12265), .ZN(n12303) );
  AOI22_X1 U15266 ( .A1(n12244), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12270) );
  AOI22_X1 U15267 ( .A1(n11578), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12269) );
  AOI22_X1 U15268 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12268) );
  AOI22_X1 U15269 ( .A1(n12042), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13091), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12267) );
  NAND4_X1 U15270 ( .A1(n12270), .A2(n12269), .A3(n12268), .A4(n12267), .ZN(
        n12276) );
  AOI22_X1 U15271 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12129), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12274) );
  AOI22_X1 U15272 ( .A1(n11938), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12229), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12273) );
  AOI22_X1 U15273 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12272) );
  AOI22_X1 U15274 ( .A1(n12285), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12271) );
  NAND4_X1 U15275 ( .A1(n12274), .A2(n12273), .A3(n12272), .A4(n12271), .ZN(
        n12275) );
  NOR2_X1 U15276 ( .A1(n12276), .A2(n12275), .ZN(n12304) );
  XOR2_X1 U15277 ( .A(n12303), .B(n12304), .Z(n12278) );
  NAND2_X1 U15278 ( .A1(n12278), .A2(n12277), .ZN(n12281) );
  INV_X1 U15279 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14444) );
  AOI21_X1 U15280 ( .B1(n14444), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12279) );
  AOI21_X1 U15281 ( .B1(n12308), .B2(P1_EAX_REG_29__SCAN_IN), .A(n12279), .ZN(
        n12280) );
  XNOR2_X1 U15282 ( .A(n12282), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14446) );
  AOI22_X1 U15283 ( .A1(n12281), .A2(n12280), .B1(n12307), .B2(n14446), .ZN(
        n14097) );
  INV_X1 U15284 ( .A(n12282), .ZN(n12283) );
  XNOR2_X1 U15285 ( .A(n13429), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14440) );
  AOI22_X1 U15286 ( .A1(n11578), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12292) );
  AOI22_X1 U15287 ( .A1(n12286), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12285), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12291) );
  AOI22_X1 U15288 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12290) );
  AOI22_X1 U15289 ( .A1(n11561), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13091), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12289) );
  NAND4_X1 U15290 ( .A1(n12292), .A2(n12291), .A3(n12290), .A4(n12289), .ZN(
        n12302) );
  AOI22_X1 U15291 ( .A1(n11938), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12129), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12300) );
  AOI22_X1 U15292 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12299) );
  AOI22_X1 U15293 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12298) );
  AOI22_X1 U15294 ( .A1(n12296), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12297) );
  NAND4_X1 U15295 ( .A1(n12300), .A2(n12299), .A3(n12298), .A4(n12297), .ZN(
        n12301) );
  NOR2_X1 U15296 ( .A1(n12302), .A2(n12301), .ZN(n12306) );
  NOR2_X1 U15297 ( .A1(n12304), .A2(n12303), .ZN(n12305) );
  XOR2_X1 U15298 ( .A(n12306), .B(n12305), .Z(n12312) );
  AOI21_X1 U15299 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20898), .A(
        n12307), .ZN(n12310) );
  NAND2_X1 U15300 ( .A1(n12308), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n12309) );
  OAI211_X1 U15301 ( .C1(n12312), .C2(n12311), .A(n12310), .B(n12309), .ZN(
        n12313) );
  OAI21_X1 U15302 ( .B1(n13425), .B2(n14440), .A(n12313), .ZN(n14087) );
  AOI22_X1 U15303 ( .A1(n12308), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n12314), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12315) );
  NAND2_X1 U15304 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20906) );
  NAND2_X1 U15305 ( .A1(n13435), .A2(n20906), .ZN(n12381) );
  XNOR2_X1 U15306 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12328) );
  NAND2_X1 U15307 ( .A1(n20686), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12332) );
  NAND2_X1 U15308 ( .A1(n12328), .A2(n12329), .ZN(n12317) );
  NAND2_X1 U15309 ( .A1(n20325), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12316) );
  NAND2_X1 U15310 ( .A1(n12317), .A2(n12316), .ZN(n12342) );
  MUX2_X1 U15311 ( .A(n15858), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n12341) );
  NAND2_X1 U15312 ( .A1(n12342), .A2(n12341), .ZN(n12319) );
  NAND2_X1 U15313 ( .A1(n15858), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12318) );
  XNOR2_X1 U15314 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12326) );
  NOR2_X1 U15315 ( .A1(n10273), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12320) );
  INV_X1 U15316 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n12321) );
  NAND2_X1 U15317 ( .A1(n12321), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12322) );
  INV_X1 U15318 ( .A(n12372), .ZN(n12323) );
  NAND2_X1 U15319 ( .A1(n12372), .A2(n12334), .ZN(n12363) );
  NAND2_X1 U15320 ( .A1(n12340), .A2(n13435), .ZN(n12360) );
  NAND2_X1 U15321 ( .A1(n12355), .A2(n12370), .ZN(n12359) );
  XNOR2_X1 U15322 ( .A(n12327), .B(n12326), .ZN(n12367) );
  XNOR2_X1 U15323 ( .A(n12329), .B(n12328), .ZN(n12369) );
  INV_X1 U15324 ( .A(n12340), .ZN(n12330) );
  NOR2_X1 U15325 ( .A1(n12369), .A2(n12330), .ZN(n12338) );
  NAND2_X1 U15326 ( .A1(n20271), .A2(n12820), .ZN(n12331) );
  NAND2_X1 U15327 ( .A1(n12331), .A2(n20241), .ZN(n12347) );
  OAI21_X1 U15328 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20686), .A(
        n12332), .ZN(n12335) );
  INV_X1 U15329 ( .A(n12335), .ZN(n12333) );
  OAI211_X1 U15330 ( .C1(n20231), .C2(n12775), .A(n12347), .B(n12333), .ZN(
        n12337) );
  INV_X1 U15331 ( .A(n12334), .ZN(n12348) );
  OAI21_X1 U15332 ( .B1(n12348), .B2(n12335), .A(n12352), .ZN(n12336) );
  NAND2_X1 U15333 ( .A1(n12337), .A2(n12336), .ZN(n12339) );
  NAND2_X1 U15334 ( .A1(n12338), .A2(n12339), .ZN(n12346) );
  OAI211_X1 U15335 ( .C1(n12340), .C2(n12339), .A(n12369), .B(n12360), .ZN(
        n12345) );
  XNOR2_X1 U15336 ( .A(n12342), .B(n12341), .ZN(n12368) );
  NAND2_X1 U15337 ( .A1(n12355), .A2(n12368), .ZN(n12343) );
  OAI211_X1 U15338 ( .C1(n12348), .C2(n12368), .A(n12343), .B(n12347), .ZN(
        n12344) );
  NAND3_X1 U15339 ( .A1(n12346), .A2(n12345), .A3(n12344), .ZN(n12350) );
  AOI22_X1 U15340 ( .A1(n12351), .A2(n12367), .B1(n12350), .B2(n12349), .ZN(
        n12357) );
  INV_X1 U15341 ( .A(n12367), .ZN(n12353) );
  NOR2_X1 U15342 ( .A1(n12353), .A2(n12352), .ZN(n12356) );
  INV_X1 U15343 ( .A(n12370), .ZN(n12354) );
  OAI22_X1 U15344 ( .A1(n12357), .A2(n12356), .B1(n12355), .B2(n12354), .ZN(
        n12358) );
  OAI21_X1 U15345 ( .B1(n12360), .B2(n12359), .A(n12358), .ZN(n12361) );
  AOI21_X1 U15346 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20902), .A(
        n12361), .ZN(n12362) );
  NAND2_X1 U15347 ( .A1(n12363), .A2(n12362), .ZN(n12364) );
  INV_X1 U15348 ( .A(n13085), .ZN(n12374) );
  NOR4_X1 U15349 ( .A1(n12370), .A2(n12369), .A3(n12368), .A4(n12367), .ZN(
        n12371) );
  OR2_X1 U15350 ( .A1(n12372), .A2(n12371), .ZN(n13999) );
  INV_X1 U15351 ( .A(n20906), .ZN(n20835) );
  NOR2_X1 U15352 ( .A1(n13999), .A2(n20835), .ZN(n12373) );
  NAND2_X1 U15353 ( .A1(n12374), .A2(n12373), .ZN(n12841) );
  INV_X1 U15354 ( .A(n14012), .ZN(n19982) );
  AOI21_X1 U15355 ( .B1(n14730), .B2(n20231), .A(n12375), .ZN(n12753) );
  AND2_X1 U15356 ( .A1(n12753), .A2(n11621), .ZN(n12849) );
  INV_X1 U15357 ( .A(n13079), .ZN(n20286) );
  NAND4_X1 U15358 ( .A1(n20286), .A2(n20263), .A3(n14012), .A4(n11623), .ZN(
        n12377) );
  NOR2_X1 U15359 ( .A1(n12378), .A2(n12377), .ZN(n12821) );
  AOI22_X1 U15360 ( .A1(n12849), .A2(n12765), .B1(n11621), .B2(n12821), .ZN(
        n12379) );
  NOR4_X1 U15361 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12385) );
  NOR4_X1 U15362 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12384) );
  NOR4_X1 U15363 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12383) );
  NOR4_X1 U15364 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12382) );
  AND4_X1 U15365 ( .A1(n12385), .A2(n12384), .A3(n12383), .A4(n12382), .ZN(
        n12390) );
  NOR4_X1 U15366 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n12388) );
  NOR4_X1 U15367 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12387) );
  NOR4_X1 U15368 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12386) );
  INV_X1 U15369 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20847) );
  AND4_X1 U15370 ( .A1(n12388), .A2(n12387), .A3(n12386), .A4(n20847), .ZN(
        n12389) );
  NAND2_X1 U15371 ( .A1(n12390), .A2(n12389), .ZN(n12391) );
  NOR3_X1 U15372 ( .A1(n14405), .A2(n20227), .A3(n12763), .ZN(n12392) );
  AOI22_X1 U15373 ( .A1(n14384), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14405), .ZN(n12393) );
  INV_X1 U15374 ( .A(n12393), .ZN(n12396) );
  INV_X1 U15375 ( .A(n20227), .ZN(n20228) );
  NOR2_X1 U15376 ( .A1(n12763), .A2(n20228), .ZN(n12394) );
  NAND2_X1 U15377 ( .A1(n14391), .A2(n12394), .ZN(n14362) );
  INV_X1 U15378 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20284) );
  NOR2_X1 U15379 ( .A1(n14362), .A2(n20284), .ZN(n12395) );
  NOR2_X1 U15380 ( .A1(n12396), .A2(n12395), .ZN(n12397) );
  AND2_X1 U15381 ( .A1(n10937), .A2(n15521), .ZN(n16351) );
  NAND2_X1 U15382 ( .A1(n12612), .A2(n16351), .ZN(n12879) );
  OR2_X1 U15383 ( .A1(n12399), .A2(n12400), .ZN(n12867) );
  NAND2_X1 U15384 ( .A1(n12879), .A2(n12867), .ZN(n12401) );
  NAND2_X1 U15385 ( .A1(n12402), .A2(n14901), .ZN(n12406) );
  NAND2_X1 U15386 ( .A1(n14919), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12403) );
  INV_X1 U15387 ( .A(n12404), .ZN(n12405) );
  NAND2_X1 U15388 ( .A1(n12406), .A2(n12405), .ZN(P2_U2857) );
  NOR2_X1 U15389 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12408) );
  NOR4_X1 U15390 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12407) );
  NAND4_X1 U15391 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12408), .A4(n12407), .ZN(n12411) );
  INV_X1 U15392 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n21241) );
  NOR3_X1 U15393 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(P1_ADS_N_REG_SCAN_IN), .A3(
        n21241), .ZN(n12410) );
  NOR4_X1 U15394 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(P1_BE_N_REG_2__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n12409)
         );
  NAND4_X1 U15395 ( .A1(n20227), .A2(P1_W_R_N_REG_SCAN_IN), .A3(n12410), .A4(
        n12409), .ZN(U214) );
  NOR2_X1 U15396 ( .A1(n13153), .A2(n12411), .ZN(n16463) );
  NAND2_X1 U15397 ( .A1(n16463), .A2(U214), .ZN(U212) );
  AOI211_X1 U15398 ( .C1(n12414), .C2(n12413), .A(n12412), .B(n19831), .ZN(
        n12426) );
  INV_X1 U15399 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n14881) );
  OAI22_X1 U15400 ( .A1(n19897), .A2(n19122), .B1(n14881), .B2(n19085), .ZN(
        n12425) );
  NAND2_X1 U15401 ( .A1(n12416), .A2(n10095), .ZN(n12417) );
  NAND2_X1 U15402 ( .A1(n12456), .A2(n12417), .ZN(n13900) );
  OAI22_X1 U15403 ( .A1(n13900), .A2(n19106), .B1(n19105), .B2(n11054), .ZN(
        n12424) );
  OAI21_X1 U15404 ( .B1(n12418), .B2(n12419), .A(n12461), .ZN(n15319) );
  AND2_X1 U15405 ( .A1(n14788), .A2(n12420), .ZN(n12421) );
  NOR2_X1 U15406 ( .A1(n9886), .A2(n12421), .ZN(n15315) );
  INV_X1 U15407 ( .A(n15315), .ZN(n12422) );
  OAI22_X1 U15408 ( .A1(n15319), .A2(n19115), .B1(n19116), .B2(n12422), .ZN(
        n12423) );
  OR4_X1 U15409 ( .A1(n12426), .A2(n12425), .A3(n12424), .A4(n12423), .ZN(
        P2_U2833) );
  AOI211_X1 U15410 ( .C1(n15072), .C2(n12428), .A(n12427), .B(n19831), .ZN(
        n12438) );
  AOI211_X1 U15411 ( .C1(P2_EBX_REG_24__SCAN_IN), .C2(n12458), .A(n19106), .B(
        n9911), .ZN(n12437) );
  NAND2_X1 U15412 ( .A1(n12459), .A2(n12429), .ZN(n12430) );
  NAND2_X1 U15413 ( .A1(n14860), .A2(n12430), .ZN(n15288) );
  NOR2_X1 U15414 ( .A1(n15288), .A2(n19115), .ZN(n12436) );
  NAND2_X1 U15415 ( .A1(n12465), .A2(n12431), .ZN(n12432) );
  NAND2_X1 U15416 ( .A1(n9874), .A2(n12432), .ZN(n15292) );
  AOI22_X1 U15417 ( .A1(P2_REIP_REG_24__SCAN_IN), .A2(n19080), .B1(
        P2_EBX_REG_24__SCAN_IN), .B2(n19109), .ZN(n12434) );
  NAND2_X1 U15418 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19089), .ZN(
        n12433) );
  OAI211_X1 U15419 ( .C1(n15292), .C2(n19116), .A(n12434), .B(n12433), .ZN(
        n12435) );
  OR4_X1 U15420 ( .A1(n12438), .A2(n12437), .A3(n12436), .A4(n12435), .ZN(
        P2_U2831) );
  AOI211_X1 U15421 ( .C1(n15041), .C2(n12440), .A(n12439), .B(n19831), .ZN(
        n12452) );
  INV_X1 U15422 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n12441) );
  OAI22_X1 U15423 ( .A1(n19907), .A2(n19122), .B1(n12441), .B2(n19085), .ZN(
        n12451) );
  NAND3_X1 U15424 ( .A1(n19267), .A2(P2_EBX_REG_27__SCAN_IN), .A3(n9878), .ZN(
        n12442) );
  NAND2_X1 U15425 ( .A1(n13920), .A2(n12442), .ZN(n13914) );
  OAI22_X1 U15426 ( .A1(n13914), .A2(n19106), .B1(n19105), .B2(n15039), .ZN(
        n12450) );
  NOR2_X1 U15427 ( .A1(n14849), .A2(n12443), .ZN(n12444) );
  OR2_X1 U15428 ( .A1(n14945), .A2(n12445), .ZN(n12447) );
  AND2_X1 U15429 ( .A1(n12447), .A2(n12446), .ZN(n15258) );
  INV_X1 U15430 ( .A(n15258), .ZN(n12448) );
  OAI22_X1 U15431 ( .A1(n15260), .A2(n19115), .B1(n12448), .B2(n19116), .ZN(
        n12449) );
  OR4_X1 U15432 ( .A1(n12452), .A2(n12451), .A3(n12450), .A4(n12449), .ZN(
        P2_U2828) );
  AOI211_X1 U15433 ( .C1(n15079), .C2(n12453), .A(n10154), .B(n19831), .ZN(
        n12470) );
  AOI22_X1 U15434 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n19080), .B1(
        P2_EBX_REG_23__SCAN_IN), .B2(n19109), .ZN(n12454) );
  INV_X1 U15435 ( .A(n12454), .ZN(n12469) );
  NAND2_X1 U15436 ( .A1(n12456), .A2(n12455), .ZN(n12457) );
  NAND2_X1 U15437 ( .A1(n12458), .A2(n12457), .ZN(n13903) );
  OAI22_X1 U15438 ( .A1(n13903), .A2(n19106), .B1(n19105), .B2(n10164), .ZN(
        n12468) );
  INV_X1 U15439 ( .A(n12459), .ZN(n12460) );
  AOI21_X1 U15440 ( .B1(n12462), .B2(n12461), .A(n12460), .ZN(n15306) );
  INV_X1 U15441 ( .A(n15306), .ZN(n12466) );
  OR2_X1 U15442 ( .A1(n9886), .A2(n12463), .ZN(n12464) );
  NAND2_X1 U15443 ( .A1(n12465), .A2(n12464), .ZN(n15304) );
  OAI22_X1 U15444 ( .A1(n12466), .A2(n19115), .B1(n19116), .B2(n15304), .ZN(
        n12467) );
  OR4_X1 U15445 ( .A1(n12470), .A2(n12469), .A3(n12468), .A4(n12467), .ZN(
        P2_U2832) );
  INV_X1 U15446 ( .A(n11452), .ZN(n12613) );
  INV_X1 U15447 ( .A(n12471), .ZN(n12472) );
  NAND2_X1 U15448 ( .A1(n12613), .A2(n12472), .ZN(n14824) );
  INV_X1 U15449 ( .A(n14824), .ZN(n12474) );
  INV_X1 U15450 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n12473) );
  OAI211_X1 U15451 ( .C1(n12474), .C2(n12473), .A(n18908), .B(n12500), .ZN(
        P2_U2814) );
  INV_X1 U15452 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12885) );
  NAND2_X1 U15453 ( .A1(n12667), .A2(n19835), .ZN(n12476) );
  NAND3_X1 U15454 ( .A1(n12476), .A2(n16348), .A3(n12475), .ZN(n12477) );
  NOR2_X1 U15455 ( .A1(n10901), .A2(n12477), .ZN(n16342) );
  INV_X1 U15456 ( .A(n16362), .ZN(n12478) );
  OR2_X1 U15457 ( .A1(n16342), .A2(n12478), .ZN(n19976) );
  INV_X1 U15458 ( .A(n19976), .ZN(n12499) );
  OAI21_X1 U15459 ( .B1(n12484), .B2(n12479), .A(n16348), .ZN(n12480) );
  NAND2_X1 U15460 ( .A1(n12480), .A2(n19832), .ZN(n12482) );
  NAND2_X1 U15461 ( .A1(n15663), .A2(n12481), .ZN(n15658) );
  OAI211_X1 U15462 ( .C1(n11166), .C2(n15658), .A(P2_STATE2_REG_1__SCAN_IN), 
        .B(n12885), .ZN(n19960) );
  NAND2_X1 U15463 ( .A1(n12482), .A2(n19960), .ZN(n19972) );
  INV_X1 U15464 ( .A(n16346), .ZN(n12680) );
  NAND2_X1 U15465 ( .A1(n12680), .A2(n13216), .ZN(n12483) );
  MUX2_X1 U15466 ( .A(n13228), .B(n12484), .S(n10906), .Z(n12589) );
  INV_X1 U15467 ( .A(n12486), .ZN(n12487) );
  OAI21_X1 U15468 ( .B1(n12589), .B2(n11438), .A(n12487), .ZN(n12491) );
  INV_X1 U15469 ( .A(n12488), .ZN(n12489) );
  NAND3_X1 U15470 ( .A1(n12491), .A2(n12490), .A3(n12489), .ZN(n12493) );
  AND2_X1 U15471 ( .A1(n12493), .A2(n12492), .ZN(n19968) );
  INV_X1 U15472 ( .A(n12494), .ZN(n12495) );
  NOR2_X1 U15473 ( .A1(n16346), .A2(n12495), .ZN(n19969) );
  NAND2_X1 U15474 ( .A1(n19968), .A2(n19969), .ZN(n12496) );
  NAND2_X1 U15475 ( .A1(n12497), .A2(n12496), .ZN(n12647) );
  AND2_X1 U15476 ( .A1(n10915), .A2(n16362), .ZN(n12498) );
  OAI21_X1 U15477 ( .B1(n12885), .B2(n12499), .A(n12596), .ZN(P2_U2819) );
  INV_X1 U15478 ( .A(n12572), .ZN(n12510) );
  OAI22_X1 U15479 ( .A1(n12570), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n13155), .ZN(n19239) );
  INV_X1 U15480 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n12725) );
  INV_X1 U15481 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n12503) );
  INV_X1 U15482 ( .A(n12500), .ZN(n12501) );
  OAI21_X1 U15483 ( .B1(n19247), .B2(n19835), .A(n12501), .ZN(n12502) );
  OAI222_X1 U15484 ( .A1(n12510), .A2(n19239), .B1(n12614), .B2(n12725), .C1(
        n12503), .C2(n12522), .ZN(P2_U2952) );
  INV_X1 U15485 ( .A(n12667), .ZN(n12507) );
  INV_X1 U15486 ( .A(n18911), .ZN(n12506) );
  INV_X1 U15487 ( .A(n18908), .ZN(n12504) );
  OAI21_X1 U15488 ( .B1(n12504), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n12506), 
        .ZN(n12505) );
  OAI21_X1 U15489 ( .B1(n12507), .B2(n12506), .A(n12505), .ZN(P2_U3612) );
  INV_X1 U15490 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n12509) );
  INV_X1 U15491 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n12508) );
  AOI22_X1 U15492 ( .A1(n13155), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n13153), .ZN(n19138) );
  OAI222_X1 U15493 ( .A1(n12509), .A2(n12614), .B1(n12508), .B2(n12522), .C1(
        n12510), .C2(n19138), .ZN(P2_U2982) );
  INV_X1 U15494 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n12512) );
  INV_X1 U15495 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n12511) );
  OAI222_X1 U15496 ( .A1(n12614), .A2(n12512), .B1(n12511), .B2(n12522), .C1(
        n12510), .C2(n19239), .ZN(P2_U2967) );
  AOI22_X1 U15497 ( .A1(P2_UWORD_REG_14__SCAN_IN), .A2(n12502), .B1(n12567), 
        .B2(P2_EAX_REG_30__SCAN_IN), .ZN(n12514) );
  INV_X1 U15498 ( .A(n19140), .ZN(n12513) );
  NAND2_X1 U15499 ( .A1(n12572), .A2(n12513), .ZN(n12552) );
  NAND2_X1 U15500 ( .A1(n12514), .A2(n12552), .ZN(P2_U2966) );
  AOI22_X1 U15501 ( .A1(P2_UWORD_REG_8__SCAN_IN), .A2(n12502), .B1(n12567), 
        .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n12516) );
  AOI22_X1 U15502 ( .A1(n13155), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n13153), .ZN(n19155) );
  INV_X1 U15503 ( .A(n19155), .ZN(n12515) );
  NAND2_X1 U15504 ( .A1(n12572), .A2(n12515), .ZN(n12538) );
  NAND2_X1 U15505 ( .A1(n12516), .A2(n12538), .ZN(P2_U2960) );
  AOI22_X1 U15506 ( .A1(P2_UWORD_REG_9__SCAN_IN), .A2(n12502), .B1(n12567), 
        .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n12521) );
  INV_X1 U15507 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n12517) );
  OR2_X1 U15508 ( .A1(n12570), .A2(n12517), .ZN(n12519) );
  NAND2_X1 U15509 ( .A1(n13153), .A2(BUF2_REG_9__SCAN_IN), .ZN(n12518) );
  AND2_X1 U15510 ( .A1(n12519), .A2(n12518), .ZN(n19153) );
  INV_X1 U15511 ( .A(n19153), .ZN(n12520) );
  NAND2_X1 U15512 ( .A1(n12572), .A2(n12520), .ZN(n12523) );
  NAND2_X1 U15513 ( .A1(n12521), .A2(n12523), .ZN(P2_U2961) );
  AOI22_X1 U15514 ( .A1(P2_LWORD_REG_9__SCAN_IN), .A2(n12576), .B1(n12567), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n12524) );
  NAND2_X1 U15515 ( .A1(n12524), .A2(n12523), .ZN(P2_U2976) );
  AOI22_X1 U15516 ( .A1(P2_LWORD_REG_3__SCAN_IN), .A2(n12576), .B1(n12567), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n12526) );
  AOI22_X1 U15517 ( .A1(n13155), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13153), .ZN(n19257) );
  INV_X1 U15518 ( .A(n19257), .ZN(n12525) );
  NAND2_X1 U15519 ( .A1(n12572), .A2(n12525), .ZN(n12565) );
  NAND2_X1 U15520 ( .A1(n12526), .A2(n12565), .ZN(P2_U2970) );
  AOI22_X1 U15521 ( .A1(P2_LWORD_REG_4__SCAN_IN), .A2(n12576), .B1(n12567), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n12527) );
  OAI22_X1 U15522 ( .A1(n12570), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n13155), .ZN(n19260) );
  INV_X1 U15523 ( .A(n19260), .ZN(n16233) );
  NAND2_X1 U15524 ( .A1(n12572), .A2(n16233), .ZN(n12541) );
  NAND2_X1 U15525 ( .A1(n12527), .A2(n12541), .ZN(P2_U2971) );
  AOI22_X1 U15526 ( .A1(P2_UWORD_REG_13__SCAN_IN), .A2(n12502), .B1(n12567), 
        .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n12531) );
  INV_X1 U15527 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16484) );
  OR2_X1 U15528 ( .A1(n12570), .A2(n16484), .ZN(n12529) );
  NAND2_X1 U15529 ( .A1(n13153), .A2(BUF2_REG_13__SCAN_IN), .ZN(n12528) );
  AND2_X1 U15530 ( .A1(n12529), .A2(n12528), .ZN(n19142) );
  INV_X1 U15531 ( .A(n19142), .ZN(n12530) );
  NAND2_X1 U15532 ( .A1(n12572), .A2(n12530), .ZN(n12550) );
  NAND2_X1 U15533 ( .A1(n12531), .A2(n12550), .ZN(P2_U2965) );
  AOI22_X1 U15534 ( .A1(P2_LWORD_REG_1__SCAN_IN), .A2(n12576), .B1(n12567), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n12533) );
  AOI22_X1 U15535 ( .A1(n13155), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13153), .ZN(n19248) );
  INV_X1 U15536 ( .A(n19248), .ZN(n12532) );
  NAND2_X1 U15537 ( .A1(n12572), .A2(n12532), .ZN(n12561) );
  NAND2_X1 U15538 ( .A1(n12533), .A2(n12561), .ZN(P2_U2968) );
  AOI22_X1 U15539 ( .A1(P2_LWORD_REG_7__SCAN_IN), .A2(n12576), .B1(n12567), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n12537) );
  INV_X1 U15540 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n12534) );
  OR2_X1 U15541 ( .A1(n12570), .A2(n12534), .ZN(n12536) );
  NAND2_X1 U15542 ( .A1(n12570), .A2(BUF2_REG_7__SCAN_IN), .ZN(n12535) );
  AND2_X1 U15543 ( .A1(n12536), .A2(n12535), .ZN(n19157) );
  INV_X1 U15544 ( .A(n19157), .ZN(n19277) );
  NAND2_X1 U15545 ( .A1(n12572), .A2(n19277), .ZN(n12563) );
  NAND2_X1 U15546 ( .A1(n12537), .A2(n12563), .ZN(P2_U2974) );
  AOI22_X1 U15547 ( .A1(P2_LWORD_REG_8__SCAN_IN), .A2(n12576), .B1(n12567), 
        .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n12539) );
  NAND2_X1 U15548 ( .A1(n12539), .A2(n12538), .ZN(P2_U2975) );
  AOI22_X1 U15549 ( .A1(P2_UWORD_REG_5__SCAN_IN), .A2(n12502), .B1(n12567), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n12540) );
  INV_X1 U15550 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16497) );
  INV_X1 U15551 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18257) );
  OAI22_X1 U15552 ( .A1(n12570), .A2(n16497), .B1(n18257), .B2(n13155), .ZN(
        n19163) );
  NAND2_X1 U15553 ( .A1(n12572), .A2(n19163), .ZN(n12559) );
  NAND2_X1 U15554 ( .A1(n12540), .A2(n12559), .ZN(P2_U2957) );
  AOI22_X1 U15555 ( .A1(P2_UWORD_REG_4__SCAN_IN), .A2(n12502), .B1(n12567), 
        .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n12542) );
  NAND2_X1 U15556 ( .A1(n12542), .A2(n12541), .ZN(P2_U2956) );
  AOI22_X1 U15557 ( .A1(P2_LWORD_REG_11__SCAN_IN), .A2(n12576), .B1(n12567), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n12547) );
  INV_X1 U15558 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n12543) );
  OR2_X1 U15559 ( .A1(n12570), .A2(n12543), .ZN(n12545) );
  NAND2_X1 U15560 ( .A1(n13153), .A2(BUF2_REG_11__SCAN_IN), .ZN(n12544) );
  AND2_X1 U15561 ( .A1(n12545), .A2(n12544), .ZN(n19148) );
  INV_X1 U15562 ( .A(n19148), .ZN(n12546) );
  NAND2_X1 U15563 ( .A1(n12572), .A2(n12546), .ZN(n12548) );
  NAND2_X1 U15564 ( .A1(n12547), .A2(n12548), .ZN(P2_U2978) );
  AOI22_X1 U15565 ( .A1(P2_UWORD_REG_11__SCAN_IN), .A2(n12502), .B1(n12567), 
        .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n12549) );
  NAND2_X1 U15566 ( .A1(n12549), .A2(n12548), .ZN(P2_U2963) );
  AOI22_X1 U15567 ( .A1(P2_LWORD_REG_13__SCAN_IN), .A2(n12576), .B1(n12567), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n12551) );
  NAND2_X1 U15568 ( .A1(n12551), .A2(n12550), .ZN(P2_U2980) );
  AOI22_X1 U15569 ( .A1(P2_LWORD_REG_14__SCAN_IN), .A2(n12502), .B1(n12567), 
        .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n12553) );
  NAND2_X1 U15570 ( .A1(n12553), .A2(n12552), .ZN(P2_U2981) );
  AOI22_X1 U15571 ( .A1(P2_LWORD_REG_2__SCAN_IN), .A2(n12576), .B1(n12567), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n12554) );
  OAI22_X1 U15572 ( .A1(n12570), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n13155), .ZN(n19253) );
  INV_X1 U15573 ( .A(n19253), .ZN(n16239) );
  NAND2_X1 U15574 ( .A1(n12572), .A2(n16239), .ZN(n12568) );
  NAND2_X1 U15575 ( .A1(n12554), .A2(n12568), .ZN(P2_U2969) );
  AOI22_X1 U15576 ( .A1(P2_UWORD_REG_6__SCAN_IN), .A2(n12502), .B1(n12567), 
        .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n12556) );
  AOI22_X1 U15577 ( .A1(n13155), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n13153), .ZN(n19159) );
  INV_X1 U15578 ( .A(n19159), .ZN(n12555) );
  NAND2_X1 U15579 ( .A1(n12572), .A2(n12555), .ZN(n12557) );
  NAND2_X1 U15580 ( .A1(n12556), .A2(n12557), .ZN(P2_U2958) );
  AOI22_X1 U15581 ( .A1(P2_LWORD_REG_6__SCAN_IN), .A2(n12576), .B1(n12567), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n12558) );
  NAND2_X1 U15582 ( .A1(n12558), .A2(n12557), .ZN(P2_U2973) );
  AOI22_X1 U15583 ( .A1(P2_LWORD_REG_5__SCAN_IN), .A2(n12576), .B1(n12567), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n12560) );
  NAND2_X1 U15584 ( .A1(n12560), .A2(n12559), .ZN(P2_U2972) );
  AOI22_X1 U15585 ( .A1(P2_UWORD_REG_1__SCAN_IN), .A2(n12576), .B1(n12567), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n12562) );
  NAND2_X1 U15586 ( .A1(n12562), .A2(n12561), .ZN(P2_U2953) );
  AOI22_X1 U15587 ( .A1(P2_UWORD_REG_7__SCAN_IN), .A2(n12502), .B1(n12567), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n12564) );
  NAND2_X1 U15588 ( .A1(n12564), .A2(n12563), .ZN(P2_U2959) );
  AOI22_X1 U15589 ( .A1(P2_UWORD_REG_3__SCAN_IN), .A2(n12576), .B1(n12567), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n12566) );
  NAND2_X1 U15590 ( .A1(n12566), .A2(n12565), .ZN(P2_U2955) );
  AOI22_X1 U15591 ( .A1(P2_UWORD_REG_2__SCAN_IN), .A2(n12576), .B1(n12567), 
        .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n12569) );
  NAND2_X1 U15592 ( .A1(n12569), .A2(n12568), .ZN(P2_U2954) );
  INV_X1 U15593 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19193) );
  MUX2_X1 U15594 ( .A(BUF1_REG_12__SCAN_IN), .B(BUF2_REG_12__SCAN_IN), .S(
        n12570), .Z(n19145) );
  NAND2_X1 U15595 ( .A1(n12572), .A2(n19145), .ZN(n12575) );
  NAND2_X1 U15596 ( .A1(n12576), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n12571) );
  OAI211_X1 U15597 ( .C1(n19193), .C2(n12614), .A(n12575), .B(n12571), .ZN(
        P2_U2979) );
  INV_X1 U15598 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n12716) );
  MUX2_X1 U15599 ( .A(BUF1_REG_10__SCAN_IN), .B(BUF2_REG_10__SCAN_IN), .S(
        n13153), .Z(n19150) );
  NAND2_X1 U15600 ( .A1(n12572), .A2(n19150), .ZN(n12578) );
  NAND2_X1 U15601 ( .A1(n12576), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n12573) );
  OAI211_X1 U15602 ( .C1(n12716), .C2(n12614), .A(n12578), .B(n12573), .ZN(
        P2_U2962) );
  INV_X1 U15603 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n12723) );
  NAND2_X1 U15604 ( .A1(n12576), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n12574) );
  OAI211_X1 U15605 ( .C1(n12723), .C2(n12614), .A(n12575), .B(n12574), .ZN(
        P2_U2964) );
  INV_X1 U15606 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19197) );
  NAND2_X1 U15607 ( .A1(n12576), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n12577) );
  OAI211_X1 U15608 ( .C1(n19197), .C2(n12614), .A(n12578), .B(n12577), .ZN(
        P2_U2977) );
  NOR2_X1 U15609 ( .A1(n12755), .A2(n13999), .ZN(n14006) );
  NAND2_X1 U15610 ( .A1(n14006), .A2(n14012), .ZN(n13424) );
  INV_X1 U15611 ( .A(n13424), .ZN(n12581) );
  INV_X1 U15612 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n21181) );
  INV_X1 U15613 ( .A(n20627), .ZN(n12580) );
  INV_X1 U15614 ( .A(n12580), .ZN(n20598) );
  NAND2_X1 U15615 ( .A1(n20598), .A2(n16192), .ZN(n19985) );
  OAI211_X1 U15616 ( .C1(n12581), .C2(n21181), .A(n13423), .B(n19985), .ZN(
        P1_U2801) );
  INV_X1 U15617 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12583) );
  AND2_X1 U15618 ( .A1(n19938), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12582) );
  OAI211_X1 U15619 ( .C1(n19247), .C2(n12583), .A(n11101), .B(n12582), .ZN(
        n12584) );
  INV_X1 U15620 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n12585) );
  MUX2_X1 U15621 ( .A(n12585), .B(n16315), .S(n14906), .Z(n12586) );
  OAI21_X1 U15622 ( .B1(n14921), .B2(n19958), .A(n12586), .ZN(P2_U2887) );
  NAND2_X1 U15623 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n12884) );
  INV_X1 U15624 ( .A(n12884), .ZN(n19961) );
  NOR2_X1 U15625 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16364) );
  NOR2_X1 U15626 ( .A1(n19961), .A2(n16364), .ZN(n12587) );
  INV_X1 U15627 ( .A(n12596), .ZN(n12590) );
  MUX2_X1 U15628 ( .A(n12589), .B(n12585), .S(n19267), .Z(n14821) );
  NOR2_X1 U15629 ( .A1(n14821), .A2(n12592), .ZN(n12606) );
  AOI21_X1 U15630 ( .B1(n12592), .B2(n14821), .A(n12606), .ZN(n16321) );
  OR2_X1 U15631 ( .A1(n13228), .A2(n13216), .ZN(n12591) );
  NAND2_X1 U15632 ( .A1(n12591), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13264) );
  OR2_X1 U15633 ( .A1(n13228), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12593) );
  NAND2_X1 U15634 ( .A1(n13264), .A2(n12593), .ZN(n16325) );
  INV_X2 U15635 ( .A(n19083), .ZN(n19223) );
  INV_X2 U15636 ( .A(n19223), .ZN(n19040) );
  OR2_X1 U15637 ( .A1(n19040), .A2(n18926), .ZN(n16323) );
  OAI21_X1 U15638 ( .B1(n19225), .B2(n16325), .A(n16323), .ZN(n12594) );
  AOI21_X1 U15639 ( .B1(n16282), .B2(n16321), .A(n12594), .ZN(n12600) );
  NOR2_X1 U15640 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15553) );
  OR2_X1 U15641 ( .A1(n19923), .A2(n15553), .ZN(n19947) );
  NAND2_X1 U15642 ( .A1(n19947), .A2(n18909), .ZN(n12595) );
  NAND2_X1 U15643 ( .A1(n19924), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12598) );
  NAND2_X1 U15644 ( .A1(n9973), .A2(n12598), .ZN(n12608) );
  OAI21_X1 U15645 ( .B1(n15162), .B2(n12608), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12599) );
  OAI211_X1 U15646 ( .C1(n13154), .C2(n16315), .A(n12600), .B(n12599), .ZN(
        P2_U3014) );
  INV_X1 U15647 ( .A(n13191), .ZN(n12611) );
  AND2_X1 U15648 ( .A1(n19223), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n12682) );
  XOR2_X1 U15649 ( .A(n13228), .B(n13226), .Z(n13263) );
  XNOR2_X1 U15650 ( .A(n13264), .B(n13263), .ZN(n12601) );
  NOR2_X1 U15651 ( .A1(n15538), .A2(n12601), .ZN(n13265) );
  AOI21_X1 U15652 ( .B1(n15538), .B2(n12601), .A(n13265), .ZN(n12602) );
  INV_X1 U15653 ( .A(n12602), .ZN(n12686) );
  NOR2_X1 U15654 ( .A1(n19225), .A2(n12686), .ZN(n12603) );
  AOI211_X1 U15655 ( .C1(n15162), .C2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n12682), .B(n12603), .ZN(n12610) );
  INV_X1 U15656 ( .A(n13246), .ZN(n12605) );
  INV_X1 U15657 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n12627) );
  NAND3_X1 U15658 ( .A1(n19267), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n12604) );
  NAND2_X1 U15659 ( .A1(n12605), .A2(n12604), .ZN(n14807) );
  INV_X1 U15660 ( .A(n12606), .ZN(n13243) );
  NAND2_X1 U15661 ( .A1(n13243), .A2(n14807), .ZN(n13244) );
  OAI21_X1 U15662 ( .B1(n14807), .B2(n13243), .A(n13244), .ZN(n12607) );
  XOR2_X1 U15663 ( .A(n12607), .B(n15538), .Z(n12683) );
  AOI22_X1 U15664 ( .A1(n16282), .A2(n12683), .B1(n19222), .B2(n14806), .ZN(
        n12609) );
  OAI211_X1 U15665 ( .C1(n12611), .C2(n13154), .A(n12610), .B(n12609), .ZN(
        P2_U3013) );
  INV_X1 U15666 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n12619) );
  INV_X1 U15667 ( .A(n12612), .ZN(n16354) );
  NAND2_X1 U15668 ( .A1(n16354), .A2(n14748), .ZN(n12658) );
  NAND2_X1 U15669 ( .A1(n12613), .A2(n16362), .ZN(n12615) );
  OAI21_X1 U15670 ( .B1(n12658), .B2(n12615), .A(n12614), .ZN(n12617) );
  INV_X1 U15671 ( .A(n19841), .ZN(n12616) );
  AND2_X1 U15672 ( .A1(n12617), .A2(n12616), .ZN(n19186) );
  NAND2_X1 U15673 ( .A1(n19186), .A2(n14747), .ZN(n12728) );
  NOR2_X1 U15674 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n12884), .ZN(n12719) );
  AOI22_X1 U15675 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n19204), .B1(n19218), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n12618) );
  OAI21_X1 U15676 ( .B1(n12619), .B2(n12728), .A(n12618), .ZN(P2_U2921) );
  INV_X1 U15677 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n14965) );
  AOI22_X1 U15678 ( .A1(n12719), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19204), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n12620) );
  OAI21_X1 U15679 ( .B1(n14965), .B2(n12728), .A(n12620), .ZN(P2_U2928) );
  INV_X1 U15680 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14953) );
  AOI22_X1 U15681 ( .A1(n12719), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19204), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n12621) );
  OAI21_X1 U15682 ( .B1(n14953), .B2(n12728), .A(n12621), .ZN(P2_U2926) );
  INV_X1 U15683 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14937) );
  AOI22_X1 U15684 ( .A1(n12719), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19204), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n12622) );
  OAI21_X1 U15685 ( .B1(n14937), .B2(n12728), .A(n12622), .ZN(P2_U2924) );
  OR2_X1 U15686 ( .A1(n12624), .A2(n12623), .ZN(n12625) );
  NOR2_X1 U15687 ( .A1(n14906), .A2(n12627), .ZN(n12628) );
  AOI21_X1 U15688 ( .B1(n14906), .B2(n13191), .A(n12628), .ZN(n12629) );
  OAI21_X1 U15689 ( .B1(n19949), .B2(n14921), .A(n12629), .ZN(P2_U2886) );
  INV_X1 U15690 ( .A(n12630), .ZN(n12631) );
  INV_X1 U15691 ( .A(n12632), .ZN(n12638) );
  INV_X1 U15692 ( .A(n12633), .ZN(n12636) );
  INV_X1 U15693 ( .A(n12634), .ZN(n12635) );
  NAND2_X1 U15694 ( .A1(n12636), .A2(n12635), .ZN(n12637) );
  NAND2_X1 U15695 ( .A1(n12638), .A2(n12637), .ZN(n16312) );
  INV_X1 U15696 ( .A(n16312), .ZN(n12640) );
  AOI22_X1 U15697 ( .A1(n19177), .A2(n12640), .B1(n19176), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n12642) );
  NOR2_X1 U15698 ( .A1(n19958), .A2(n16312), .ZN(n19180) );
  INV_X1 U15699 ( .A(n19180), .ZN(n12639) );
  OAI211_X1 U15700 ( .C1(n19488), .C2(n12640), .A(n12639), .B(n19137), .ZN(
        n12641) );
  OAI211_X1 U15701 ( .C1(n19185), .C2(n19239), .A(n12642), .B(n12641), .ZN(
        P2_U2919) );
  INV_X1 U15702 ( .A(n12658), .ZN(n12643) );
  NAND2_X1 U15703 ( .A1(n12643), .A2(n12649), .ZN(n12877) );
  OAI21_X1 U15704 ( .B1(n12645), .B2(n10915), .A(n12644), .ZN(n12646) );
  INV_X1 U15705 ( .A(n12646), .ZN(n12657) );
  INV_X1 U15706 ( .A(n12647), .ZN(n12655) );
  AND3_X1 U15707 ( .A1(n10914), .A2(n16348), .A3(n12649), .ZN(n12650) );
  NOR2_X1 U15708 ( .A1(n12651), .A2(n12650), .ZN(n12878) );
  MUX2_X1 U15709 ( .A(n12648), .B(n12652), .S(n19247), .Z(n12653) );
  NAND3_X1 U15710 ( .A1(n12653), .A2(n16348), .A3(n19835), .ZN(n12654) );
  NAND3_X1 U15711 ( .A1(n12655), .A2(n12878), .A3(n12654), .ZN(n12656) );
  AOI21_X1 U15712 ( .B1(n12658), .B2(n12657), .A(n12656), .ZN(n12659) );
  OAI21_X1 U15713 ( .B1(n12877), .B2(n19252), .A(n12659), .ZN(n12660) );
  INV_X1 U15714 ( .A(n12661), .ZN(n12662) );
  AOI21_X1 U15715 ( .B1(n14748), .B2(n16350), .A(n16351), .ZN(n12663) );
  XNOR2_X1 U15716 ( .A(n12665), .B(n12664), .ZN(n19953) );
  INV_X1 U15717 ( .A(n19953), .ZN(n12904) );
  NAND2_X1 U15718 ( .A1(n12681), .A2(n19083), .ZN(n16316) );
  OAI22_X1 U15719 ( .A1(n16313), .A2(n12904), .B1(n16316), .B2(n15538), .ZN(
        n12688) );
  INV_X1 U15720 ( .A(n19969), .ZN(n12666) );
  OAI211_X1 U15721 ( .C1(n10949), .C2(n10915), .A(n10909), .B(n12399), .ZN(
        n12671) );
  OAI22_X1 U15722 ( .A1(n12667), .A2(n10905), .B1(n16347), .B2(n19252), .ZN(
        n12668) );
  INV_X1 U15723 ( .A(n12668), .ZN(n12670) );
  NAND3_X1 U15724 ( .A1(n12671), .A2(n12670), .A3(n12669), .ZN(n12676) );
  NAND2_X1 U15725 ( .A1(n12672), .A2(n14748), .ZN(n15523) );
  AOI21_X1 U15726 ( .B1(n15523), .B2(n12674), .A(n12673), .ZN(n12675) );
  OR2_X1 U15727 ( .A1(n12676), .A2(n12675), .ZN(n15550) );
  INV_X1 U15728 ( .A(n12867), .ZN(n12677) );
  NOR2_X1 U15729 ( .A1(n15550), .A2(n12677), .ZN(n12678) );
  OR2_X1 U15730 ( .A1(n12681), .A2(n12678), .ZN(n15377) );
  INV_X1 U15731 ( .A(n15381), .ZN(n16318) );
  NAND2_X1 U15732 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13254) );
  OAI211_X1 U15733 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n16318), .B(n13254), .ZN(n12685) );
  NAND2_X1 U15734 ( .A1(n12680), .A2(n12679), .ZN(n19967) );
  AOI21_X1 U15735 ( .B1(n16322), .B2(n12683), .A(n12682), .ZN(n12684) );
  OAI211_X1 U15736 ( .C1(n16326), .C2(n12686), .A(n12685), .B(n12684), .ZN(
        n12687) );
  AOI211_X1 U15737 ( .C1(n13191), .C2(n16304), .A(n12688), .B(n12687), .ZN(
        n12689) );
  INV_X1 U15738 ( .A(n12689), .ZN(P2_U3045) );
  INV_X1 U15739 ( .A(n13185), .ZN(n13188) );
  MUX2_X1 U15740 ( .A(n9829), .B(n13537), .S(n14919), .Z(n12693) );
  OAI21_X1 U15741 ( .B1(n19936), .B2(n14921), .A(n12693), .ZN(P2_U2885) );
  INV_X1 U15742 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n21256) );
  NOR2_X1 U15743 ( .A1(n12755), .A2(n20241), .ZN(n14734) );
  NAND2_X1 U15744 ( .A1(n14005), .A2(n20241), .ZN(n12791) );
  INV_X1 U15745 ( .A(n12791), .ZN(n12694) );
  OR2_X1 U15746 ( .A1(n14734), .A2(n12694), .ZN(n12698) );
  INV_X1 U15747 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n12695) );
  NAND2_X1 U15748 ( .A1(n12696), .A2(n12695), .ZN(n15906) );
  INV_X1 U15749 ( .A(n15906), .ZN(n15873) );
  NAND2_X1 U15750 ( .A1(n20105), .A2(n12820), .ZN(n13017) );
  NAND2_X1 U15751 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16188) );
  INV_X1 U15752 ( .A(n16188), .ZN(n13113) );
  NAND2_X1 U15753 ( .A1(n20902), .A2(n13113), .ZN(n20103) );
  NOR2_X4 U15754 ( .A1(n20105), .A2(n20132), .ZN(n15908) );
  AOI22_X1 U15755 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n12699) );
  OAI21_X1 U15756 ( .B1(n21256), .B2(n13017), .A(n12699), .ZN(P1_U2916) );
  INV_X1 U15757 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n21247) );
  AOI22_X1 U15758 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n12700) );
  OAI21_X1 U15759 ( .B1(n21247), .B2(n13017), .A(n12700), .ZN(P1_U2913) );
  INV_X1 U15760 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n12702) );
  AOI22_X1 U15761 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n12701) );
  OAI21_X1 U15762 ( .B1(n12702), .B2(n13017), .A(n12701), .ZN(P1_U2917) );
  INV_X1 U15763 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n21244) );
  AOI22_X1 U15764 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n12703) );
  OAI21_X1 U15765 ( .B1(n21244), .B2(n13017), .A(n12703), .ZN(P1_U2914) );
  AOI22_X1 U15766 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n12704) );
  OAI21_X1 U15767 ( .B1(n21275), .B2(n13017), .A(n12704), .ZN(P1_U2908) );
  INV_X1 U15768 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n20953) );
  AOI22_X1 U15769 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12705) );
  OAI21_X1 U15770 ( .B1(n20953), .B2(n13017), .A(n12705), .ZN(P1_U2907) );
  INV_X1 U15771 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n20984) );
  AOI22_X1 U15772 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n12706) );
  OAI21_X1 U15773 ( .B1(n20984), .B2(n13017), .A(n12706), .ZN(P1_U2915) );
  INV_X1 U15774 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n21279) );
  AOI22_X1 U15775 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n12707) );
  OAI21_X1 U15776 ( .B1(n21279), .B2(n13017), .A(n12707), .ZN(P1_U2911) );
  INV_X1 U15777 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13026) );
  AOI22_X1 U15778 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n12708) );
  OAI21_X1 U15779 ( .B1(n13026), .B2(n13017), .A(n12708), .ZN(P1_U2909) );
  INV_X1 U15780 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n21187) );
  AOI22_X1 U15781 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n12709) );
  OAI21_X1 U15782 ( .B1(n21187), .B2(n13017), .A(n12709), .ZN(P1_U2912) );
  INV_X1 U15783 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n14959) );
  AOI22_X1 U15784 ( .A1(n12719), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19217), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n12710) );
  OAI21_X1 U15785 ( .B1(n14959), .B2(n12728), .A(n12710), .ZN(P2_U2927) );
  INV_X1 U15786 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n14973) );
  AOI22_X1 U15787 ( .A1(n12719), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19217), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n12711) );
  OAI21_X1 U15788 ( .B1(n14973), .B2(n12728), .A(n12711), .ZN(P2_U2929) );
  INV_X1 U15789 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n14987) );
  AOI22_X1 U15790 ( .A1(n12719), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19217), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n12712) );
  OAI21_X1 U15791 ( .B1(n14987), .B2(n12728), .A(n12712), .ZN(P2_U2932) );
  INV_X1 U15792 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n12714) );
  AOI22_X1 U15793 ( .A1(n12719), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19217), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n12713) );
  OAI21_X1 U15794 ( .B1(n12714), .B2(n12728), .A(n12713), .ZN(P2_U2933) );
  AOI22_X1 U15795 ( .A1(n12719), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19217), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n12715) );
  OAI21_X1 U15796 ( .B1(n12716), .B2(n12728), .A(n12715), .ZN(P2_U2925) );
  INV_X1 U15797 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n12718) );
  AOI22_X1 U15798 ( .A1(n12719), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19217), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n12717) );
  OAI21_X1 U15799 ( .B1(n12718), .B2(n12728), .A(n12717), .ZN(P2_U2930) );
  INV_X1 U15800 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n12721) );
  AOI22_X1 U15801 ( .A1(n12719), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19217), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n12720) );
  OAI21_X1 U15802 ( .B1(n12721), .B2(n12728), .A(n12720), .ZN(P2_U2931) );
  AOI22_X1 U15803 ( .A1(n19218), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19217), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12722) );
  OAI21_X1 U15804 ( .B1(n12723), .B2(n12728), .A(n12722), .ZN(P2_U2923) );
  AOI22_X1 U15805 ( .A1(n19218), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19217), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n12724) );
  OAI21_X1 U15806 ( .B1(n12725), .B2(n12728), .A(n12724), .ZN(P2_U2935) );
  AOI22_X1 U15807 ( .A1(n19218), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19217), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n12726) );
  OAI21_X1 U15808 ( .B1(n13469), .B2(n12728), .A(n12726), .ZN(P2_U2934) );
  INV_X1 U15809 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14923) );
  AOI22_X1 U15810 ( .A1(n19218), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19217), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12727) );
  OAI21_X1 U15811 ( .B1(n14923), .B2(n12728), .A(n12727), .ZN(P2_U2922) );
  NAND3_X1 U15812 ( .A1(n20902), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16187) );
  INV_X1 U15813 ( .A(n16187), .ZN(n12729) );
  INV_X1 U15814 ( .A(n20158), .ZN(n15997) );
  INV_X1 U15815 ( .A(n12730), .ZN(n12733) );
  OAI21_X1 U15816 ( .B1(n12733), .B2(n12732), .A(n12731), .ZN(n20086) );
  NAND2_X1 U15817 ( .A1(n20902), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12735) );
  NAND2_X1 U15818 ( .A1(n21280), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12734) );
  AND2_X1 U15819 ( .A1(n12735), .A2(n12734), .ZN(n12807) );
  NAND3_X1 U15820 ( .A1(n12753), .A2(n12736), .A3(n12774), .ZN(n12768) );
  NAND2_X1 U15821 ( .A1(n12580), .A2(n12738), .ZN(n20905) );
  AND2_X1 U15822 ( .A1(n20905), .A2(n20902), .ZN(n12737) );
  NAND2_X1 U15823 ( .A1(n12807), .A2(n16041), .ZN(n12746) );
  NOR2_X1 U15824 ( .A1(n20207), .A2(n21162), .ZN(n12800) );
  INV_X1 U15825 ( .A(n13494), .ZN(n13064) );
  NAND2_X1 U15826 ( .A1(n20231), .A2(n12740), .ZN(n12956) );
  OAI21_X1 U15827 ( .B1(n15872), .B2(n12812), .A(n12956), .ZN(n12741) );
  INV_X1 U15828 ( .A(n12741), .ZN(n12742) );
  NAND2_X1 U15829 ( .A1(n12744), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12953) );
  OAI21_X1 U15830 ( .B1(n12744), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12953), .ZN(n12803) );
  NOR2_X1 U15831 ( .A1(n12803), .A2(n19988), .ZN(n12745) );
  AOI211_X1 U15832 ( .C1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n12746), .A(
        n12800), .B(n12745), .ZN(n12747) );
  OAI21_X1 U15833 ( .B1(n15997), .B2(n20086), .A(n12747), .ZN(P1_U2999) );
  INV_X1 U15834 ( .A(n13532), .ZN(n13253) );
  MUX2_X1 U15835 ( .A(n10979), .B(n13253), .S(n14906), .Z(n12752) );
  OAI21_X1 U15836 ( .B1(n19522), .B2(n14921), .A(n12752), .ZN(P2_U2884) );
  NAND2_X1 U15837 ( .A1(n12753), .A2(n12774), .ZN(n12754) );
  NAND2_X1 U15838 ( .A1(n12755), .A2(n12754), .ZN(n12758) );
  OR2_X1 U15839 ( .A1(n13080), .A2(n20241), .ZN(n12778) );
  AND2_X1 U15840 ( .A1(n12778), .A2(n12820), .ZN(n12756) );
  NAND2_X1 U15841 ( .A1(n12757), .A2(n12756), .ZN(n12784) );
  NAND2_X1 U15842 ( .A1(n12758), .A2(n12784), .ZN(n12838) );
  NAND2_X1 U15843 ( .A1(n10058), .A2(n13435), .ZN(n12761) );
  NAND2_X1 U15844 ( .A1(n13435), .A2(n15906), .ZN(n12759) );
  NAND3_X1 U15845 ( .A1(n12759), .A2(n12837), .A3(n20906), .ZN(n12760) );
  OAI22_X1 U15846 ( .A1(n14003), .A2(n12761), .B1(n13999), .B2(n12760), .ZN(
        n12762) );
  OAI21_X1 U15847 ( .B1(n12838), .B2(n12762), .A(n14012), .ZN(n12767) );
  OAI21_X1 U15848 ( .B1(n13435), .B2(n15873), .A(n20906), .ZN(n13432) );
  OAI211_X1 U15849 ( .C1(n12831), .C2(n13432), .A(n12820), .B(n12763), .ZN(
        n12764) );
  NAND3_X1 U15850 ( .A1(n12765), .A2(n20248), .A3(n12764), .ZN(n12766) );
  INV_X1 U15851 ( .A(n12849), .ZN(n12834) );
  AND2_X1 U15852 ( .A1(n12834), .A2(n12768), .ZN(n14004) );
  INV_X1 U15853 ( .A(n12793), .ZN(n12769) );
  AOI22_X1 U15854 ( .A1(n12769), .A2(n12792), .B1(n14005), .B2(n13435), .ZN(
        n12770) );
  NAND3_X1 U15855 ( .A1(n14004), .A2(n13085), .A3(n12770), .ZN(n12771) );
  INV_X1 U15856 ( .A(n12772), .ZN(n12773) );
  OAI21_X1 U15857 ( .B1(n12774), .B2(n14082), .A(n12773), .ZN(n12781) );
  OAI21_X1 U15858 ( .B1(n12775), .B2(n13092), .A(n20231), .ZN(n12777) );
  AOI21_X1 U15859 ( .B1(n20278), .B2(n12837), .A(n20286), .ZN(n12776) );
  NAND2_X1 U15860 ( .A1(n12777), .A2(n12776), .ZN(n12782) );
  INV_X1 U15861 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20190) );
  INV_X2 U15862 ( .A(n20207), .ZN(n20150) );
  INV_X1 U15863 ( .A(n11640), .ZN(n12780) );
  NAND2_X1 U15864 ( .A1(n12780), .A2(n11621), .ZN(n12786) );
  INV_X1 U15865 ( .A(n12781), .ZN(n12785) );
  NAND2_X1 U15866 ( .A1(n12782), .A2(n13435), .ZN(n12783) );
  NAND4_X1 U15867 ( .A1(n12786), .A2(n12785), .A3(n12784), .A4(n12783), .ZN(
        n12828) );
  INV_X1 U15868 ( .A(n12828), .ZN(n12788) );
  OAI211_X1 U15869 ( .C1(n14082), .C2(n12820), .A(n12788), .B(n12787), .ZN(
        n12789) );
  NAND2_X1 U15870 ( .A1(n12795), .A2(n12789), .ZN(n14680) );
  OAI22_X1 U15871 ( .A1(n20150), .A2(n12795), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n14680), .ZN(n14696) );
  AOI21_X1 U15872 ( .B1(n20193), .B2(n20190), .A(n14696), .ZN(n20216) );
  INV_X2 U15873 ( .A(n20193), .ZN(n20195) );
  AND2_X1 U15874 ( .A1(n20195), .A2(n14680), .ZN(n13506) );
  AOI22_X1 U15875 ( .A1(n20216), .A2(n16117), .B1(n20190), .B2(n13506), .ZN(
        n12790) );
  INV_X1 U15876 ( .A(n12790), .ZN(n12802) );
  OAI21_X1 U15877 ( .B1(n12793), .B2(n12792), .A(n12791), .ZN(n12794) );
  NAND2_X1 U15878 ( .A1(n14046), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12798) );
  INV_X1 U15879 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n12796) );
  NAND2_X1 U15880 ( .A1(n14082), .A2(n12796), .ZN(n12797) );
  NOR2_X1 U15881 ( .A1(n14071), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12799) );
  OR2_X1 U15882 ( .A1(n12926), .A2(n12799), .ZN(n12824) );
  INV_X1 U15883 ( .A(n12824), .ZN(n20076) );
  AOI21_X1 U15884 ( .B1(n20214), .B2(n20076), .A(n12800), .ZN(n12801) );
  OAI211_X1 U15885 ( .C1(n20196), .C2(n12803), .A(n12802), .B(n12801), .ZN(
        P1_U3031) );
  OR2_X1 U15886 ( .A1(n12805), .A2(n12804), .ZN(n12806) );
  NAND2_X1 U15887 ( .A1(n12930), .A2(n12806), .ZN(n20066) );
  INV_X1 U15888 ( .A(n12807), .ZN(n12808) );
  INV_X1 U15889 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20062) );
  OAI22_X1 U15890 ( .A1(n16041), .A2(n20062), .B1(n20207), .B2(n20889), .ZN(
        n12809) );
  AOI21_X1 U15891 ( .B1(n16037), .B2(n20062), .A(n12809), .ZN(n12819) );
  NAND2_X1 U15892 ( .A1(n12811), .A2(n12812), .ZN(n13066) );
  OAI21_X1 U15893 ( .B1(n12812), .B2(n12811), .A(n13066), .ZN(n12813) );
  OAI211_X1 U15894 ( .C1(n12813), .C2(n15872), .A(n20248), .B(n14328), .ZN(
        n12814) );
  INV_X1 U15895 ( .A(n12814), .ZN(n12815) );
  XNOR2_X1 U15896 ( .A(n12951), .B(n12953), .ZN(n12817) );
  OR2_X1 U15897 ( .A1(n12817), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20209) );
  NAND2_X1 U15898 ( .A1(n12817), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20210) );
  NAND3_X1 U15899 ( .A1(n20209), .A2(n20210), .A3(n20159), .ZN(n12818) );
  OAI211_X1 U15900 ( .C1(n20066), .C2(n15997), .A(n12819), .B(n12818), .ZN(
        P1_U2998) );
  NAND2_X1 U15901 ( .A1(n12821), .A2(n14067), .ZN(n12822) );
  OAI222_X1 U15902 ( .A1(n20086), .A2(n14326), .B1(n20101), .B2(n12796), .C1(
        n12824), .C2(n14316), .ZN(P1_U2872) );
  INV_X1 U15903 ( .A(n11839), .ZN(n13114) );
  NAND3_X1 U15904 ( .A1(n12826), .A2(n12831), .A3(n12825), .ZN(n12827) );
  NOR2_X1 U15905 ( .A1(n12828), .A2(n12827), .ZN(n12829) );
  AND2_X1 U15906 ( .A1(n12829), .A2(n13085), .ZN(n14731) );
  OAI22_X1 U15907 ( .A1(n13114), .A2(n14731), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14730), .ZN(n15852) );
  OAI22_X1 U15908 ( .A1(n16192), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15882), .ZN(n12830) );
  AOI21_X1 U15909 ( .B1(n15852), .B2(n16181), .A(n12830), .ZN(n12847) );
  INV_X1 U15910 ( .A(n12831), .ZN(n15874) );
  INV_X1 U15911 ( .A(n14005), .ZN(n12832) );
  AOI21_X1 U15912 ( .B1(n12832), .B2(n15906), .A(n13432), .ZN(n12833) );
  OAI21_X1 U15913 ( .B1(n14734), .B2(n15874), .A(n12833), .ZN(n12835) );
  NAND2_X1 U15914 ( .A1(n12835), .A2(n12834), .ZN(n12836) );
  NAND2_X1 U15915 ( .A1(n12836), .A2(n14003), .ZN(n12843) );
  NAND2_X1 U15916 ( .A1(n20231), .A2(n13435), .ZN(n14255) );
  NOR2_X1 U15917 ( .A1(n14255), .A2(n12837), .ZN(n12839) );
  NOR3_X1 U15918 ( .A1(n12840), .A2(n12839), .A3(n12838), .ZN(n12842) );
  NAND2_X1 U15919 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n13113), .ZN(n16193) );
  INV_X1 U15920 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n21022) );
  OAI22_X1 U15921 ( .A1(n15853), .A2(n19982), .B1(n16193), .B2(n21022), .ZN(
        n16180) );
  AOI21_X1 U15922 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20902), .A(n16180), 
        .ZN(n12857) );
  INV_X1 U15923 ( .A(n14734), .ZN(n12845) );
  NOR2_X1 U15924 ( .A1(n12845), .A2(n12844), .ZN(n15851) );
  AOI22_X1 U15925 ( .A1(n15851), .A2(n16181), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n12857), .ZN(n12846) );
  OAI21_X1 U15926 ( .B1(n12847), .B2(n12857), .A(n12846), .ZN(P1_U3474) );
  OR2_X1 U15927 ( .A1(n14000), .A2(n12849), .ZN(n13099) );
  XNOR2_X1 U15928 ( .A(n14735), .B(n12859), .ZN(n12854) );
  INV_X1 U15929 ( .A(n12854), .ZN(n12851) );
  XNOR2_X1 U15930 ( .A(n11710), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12850) );
  AOI22_X1 U15931 ( .A1(n13099), .A2(n12851), .B1(n14734), .B2(n12850), .ZN(
        n12853) );
  NAND3_X1 U15932 ( .A1(n14731), .A2(n13092), .A3(n12854), .ZN(n12852) );
  OAI211_X1 U15933 ( .C1(n20631), .C2(n14731), .A(n12853), .B(n12852), .ZN(
        n13088) );
  INV_X1 U15934 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14602) );
  INV_X1 U15935 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20217) );
  OAI22_X1 U15936 ( .A1(n14602), .A2(n20217), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14738) );
  INV_X1 U15937 ( .A(n14738), .ZN(n12856) );
  NOR2_X1 U15938 ( .A1(n16192), .A2(n20190), .ZN(n14737) );
  INV_X1 U15939 ( .A(n15882), .ZN(n12855) );
  AOI222_X1 U15940 ( .A1(n13088), .A2(n16181), .B1(n12856), .B2(n14737), .C1(
        n12855), .C2(n12854), .ZN(n12858) );
  INV_X1 U15941 ( .A(n12857), .ZN(n16185) );
  MUX2_X1 U15942 ( .A(n12859), .B(n12858), .S(n16185), .Z(n12860) );
  INV_X1 U15943 ( .A(n12860), .ZN(P1_U3472) );
  INV_X1 U15944 ( .A(n19522), .ZN(n19928) );
  NAND2_X1 U15945 ( .A1(n13532), .A2(n15550), .ZN(n12876) );
  INV_X1 U15946 ( .A(n16351), .ZN(n12861) );
  NAND2_X1 U15947 ( .A1(n16353), .A2(n12861), .ZN(n15542) );
  NOR2_X1 U15948 ( .A1(n12862), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15548) );
  INV_X1 U15949 ( .A(n15548), .ZN(n12866) );
  NAND2_X1 U15950 ( .A1(n9821), .A2(n12863), .ZN(n12864) );
  NAND2_X1 U15951 ( .A1(n12864), .A2(n12869), .ZN(n12865) );
  AOI21_X1 U15952 ( .B1(n15542), .B2(n12866), .A(n12865), .ZN(n12874) );
  NAND2_X1 U15953 ( .A1(n12867), .A2(n10943), .ZN(n12870) );
  NAND2_X1 U15954 ( .A1(n12870), .A2(n12869), .ZN(n15547) );
  INV_X1 U15955 ( .A(n12863), .ZN(n12871) );
  NAND2_X1 U15956 ( .A1(n9821), .A2(n12871), .ZN(n15544) );
  NAND2_X1 U15957 ( .A1(n15547), .A2(n15544), .ZN(n12872) );
  AOI21_X1 U15958 ( .B1(n15548), .B2(n15542), .A(n12872), .ZN(n12873) );
  MUX2_X1 U15959 ( .A(n12874), .B(n12873), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12875) );
  NAND2_X1 U15960 ( .A1(n12876), .A2(n12875), .ZN(n16327) );
  AOI22_X1 U15961 ( .A1(n19928), .A2(n16365), .B1(n16327), .B2(n15553), .ZN(
        n12888) );
  OR2_X1 U15962 ( .A1(n12877), .A2(n11452), .ZN(n12883) );
  NAND2_X1 U15963 ( .A1(n12879), .A2(n12878), .ZN(n12880) );
  NOR2_X1 U15964 ( .A1(n12881), .A2(n12880), .ZN(n12882) );
  NAND2_X1 U15965 ( .A1(n12883), .A2(n12882), .ZN(n16330) );
  NOR2_X1 U15966 ( .A1(n18909), .A2(n12884), .ZN(n16373) );
  INV_X1 U15967 ( .A(n16373), .ZN(n16372) );
  OAI22_X1 U15968 ( .A1(n16372), .A2(n12885), .B1(P2_STATE2_REG_0__SCAN_IN), 
        .B2(n19938), .ZN(n12886) );
  AOI21_X1 U15969 ( .B1(n16330), .B2(n16362), .A(n12886), .ZN(n15557) );
  NAND2_X1 U15970 ( .A1(n15557), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12887) );
  OAI21_X1 U15971 ( .B1(n12888), .B2(n15557), .A(n12887), .ZN(P2_U3596) );
  INV_X1 U15972 ( .A(n12890), .ZN(n12891) );
  NAND2_X1 U15973 ( .A1(n12892), .A2(n12891), .ZN(n12894) );
  OAI21_X1 U15974 ( .B1(n12889), .B2(n12894), .A(n12893), .ZN(n19164) );
  AOI21_X1 U15975 ( .B1(n12896), .B2(n12895), .A(n12912), .ZN(n19230) );
  NOR2_X1 U15976 ( .A1(n14906), .A2(n12897), .ZN(n12898) );
  AOI21_X1 U15977 ( .B1(n19230), .B2(n14906), .A(n12898), .ZN(n12899) );
  OAI21_X1 U15978 ( .B1(n19164), .B2(n14921), .A(n12899), .ZN(P2_U2883) );
  NAND2_X1 U15979 ( .A1(n12901), .A2(n12900), .ZN(n12903) );
  XNOR2_X1 U15980 ( .A(n19936), .B(n19939), .ZN(n12908) );
  NAND2_X1 U15981 ( .A1(n19949), .A2(n12904), .ZN(n12905) );
  OAI21_X1 U15982 ( .B1(n19949), .B2(n12904), .A(n12905), .ZN(n19179) );
  NOR2_X1 U15983 ( .A1(n19179), .A2(n19180), .ZN(n19178) );
  INV_X1 U15984 ( .A(n12905), .ZN(n12906) );
  NOR2_X1 U15985 ( .A1(n19178), .A2(n12906), .ZN(n12907) );
  NOR2_X1 U15986 ( .A1(n12908), .A2(n12907), .ZN(n13167) );
  AOI21_X1 U15987 ( .B1(n12908), .B2(n12907), .A(n13167), .ZN(n12911) );
  AOI22_X1 U15988 ( .A1(n19162), .A2(n16239), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19176), .ZN(n12910) );
  INV_X1 U15989 ( .A(n19939), .ZN(n13798) );
  NAND2_X1 U15990 ( .A1(n13798), .A2(n19177), .ZN(n12909) );
  OAI211_X1 U15991 ( .C1(n12911), .C2(n19181), .A(n12910), .B(n12909), .ZN(
        P2_U2917) );
  XOR2_X1 U15992 ( .A(n12893), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n12916)
         );
  OR2_X1 U15993 ( .A1(n12913), .A2(n12912), .ZN(n12914) );
  NAND2_X1 U15994 ( .A1(n12914), .A2(n12944), .ZN(n19114) );
  MUX2_X1 U15995 ( .A(n10988), .B(n19114), .S(n14906), .Z(n12915) );
  OAI21_X1 U15996 ( .B1(n12916), .B2(n14921), .A(n12915), .ZN(P2_U2882) );
  XNOR2_X1 U15997 ( .A(n12917), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12921) );
  OR2_X1 U15998 ( .A1(n12918), .A2(n12946), .ZN(n12919) );
  NAND2_X1 U15999 ( .A1(n12919), .A2(n13036), .ZN(n19086) );
  MUX2_X1 U16000 ( .A(n10997), .B(n19086), .S(n14906), .Z(n12920) );
  OAI21_X1 U16001 ( .B1(n12921), .B2(n14921), .A(n12920), .ZN(P2_U2880) );
  INV_X1 U16002 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n20065) );
  NAND2_X1 U16003 ( .A1(n14062), .A2(n20065), .ZN(n12925) );
  NAND2_X1 U16004 ( .A1(n14046), .A2(n20217), .ZN(n12923) );
  NAND2_X1 U16005 ( .A1(n14067), .A2(n20065), .ZN(n12922) );
  NAND3_X1 U16006 ( .A1(n12923), .A2(n14082), .A3(n12922), .ZN(n12924) );
  NAND2_X1 U16007 ( .A1(n12925), .A2(n12924), .ZN(n12932) );
  XNOR2_X1 U16008 ( .A(n20072), .B(n14070), .ZN(n20213) );
  INV_X1 U16009 ( .A(n20101), .ZN(n14304) );
  AOI22_X1 U16010 ( .A1(n20097), .A2(n20213), .B1(n14304), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n12927) );
  OAI21_X1 U16011 ( .B1(n20066), .B2(n14326), .A(n12927), .ZN(P1_U2871) );
  INV_X1 U16012 ( .A(n12928), .ZN(n12929) );
  AOI21_X1 U16013 ( .B1(n12931), .B2(n12930), .A(n12929), .ZN(n14276) );
  INV_X1 U16014 ( .A(n14276), .ZN(n13083) );
  INV_X1 U16015 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n12933) );
  NAND2_X1 U16016 ( .A1(n14062), .A2(n12933), .ZN(n12937) );
  INV_X1 U16017 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20203) );
  NAND2_X1 U16018 ( .A1(n14046), .A2(n20203), .ZN(n12935) );
  NAND2_X1 U16019 ( .A1(n14067), .A2(n12933), .ZN(n12934) );
  NAND3_X1 U16020 ( .A1(n12935), .A2(n14082), .A3(n12934), .ZN(n12936) );
  AND2_X1 U16021 ( .A1(n12937), .A2(n12936), .ZN(n12938) );
  AND2_X1 U16022 ( .A1(n12939), .A2(n12938), .ZN(n12940) );
  OR2_X1 U16023 ( .A1(n12940), .A2(n13120), .ZN(n14272) );
  INV_X1 U16024 ( .A(n14272), .ZN(n20200) );
  AOI22_X1 U16025 ( .A1(n20097), .A2(n20200), .B1(n14304), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n12941) );
  OAI21_X1 U16026 ( .B1(n13083), .B2(n14326), .A(n12941), .ZN(P1_U2870) );
  NOR2_X1 U16027 ( .A1(n12893), .A2(n11210), .ZN(n12943) );
  INV_X1 U16028 ( .A(n12917), .ZN(n12942) );
  OAI211_X1 U16029 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n12943), .A(
        n12942), .B(n14901), .ZN(n12949) );
  NAND2_X1 U16030 ( .A1(n12945), .A2(n12944), .ZN(n12947) );
  AND2_X1 U16031 ( .A1(n12947), .A2(n10198), .ZN(n19100) );
  NAND2_X1 U16032 ( .A1(n14906), .A2(n19100), .ZN(n12948) );
  OAI211_X1 U16033 ( .C1(n14906), .C2(n12950), .A(n12949), .B(n12948), .ZN(
        P2_U2881) );
  INV_X1 U16034 ( .A(n12951), .ZN(n12952) );
  OR2_X1 U16035 ( .A1(n12953), .A2(n12952), .ZN(n12954) );
  XNOR2_X1 U16036 ( .A(n13066), .B(n13065), .ZN(n12958) );
  INV_X1 U16037 ( .A(n15872), .ZN(n13488) );
  INV_X1 U16038 ( .A(n12956), .ZN(n12957) );
  AOI21_X1 U16039 ( .B1(n12958), .B2(n13488), .A(n12957), .ZN(n12959) );
  NAND2_X1 U16040 ( .A1(n12960), .A2(n12959), .ZN(n12961) );
  NAND2_X1 U16041 ( .A1(n12962), .A2(n12961), .ZN(n13062) );
  OAI21_X1 U16042 ( .B1(n12962), .B2(n12961), .A(n13062), .ZN(n20197) );
  AOI22_X1 U16043 ( .A1(n20151), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20150), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n12963) );
  OAI21_X1 U16044 ( .B1(n20164), .B2(n14269), .A(n12963), .ZN(n12964) );
  AOI21_X1 U16045 ( .B1(n14276), .B2(n20158), .A(n12964), .ZN(n12965) );
  OAI21_X1 U16046 ( .B1(n19988), .B2(n20197), .A(n12965), .ZN(P1_U2997) );
  NOR2_X2 U16047 ( .A1(n20146), .A2(n20241), .ZN(n13030) );
  MUX2_X1 U16048 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n20227), .Z(
        n14401) );
  NAND2_X1 U16049 ( .A1(n13030), .A2(n14401), .ZN(n20142) );
  AOI22_X1 U16050 ( .A1(n20147), .A2(P1_EAX_REG_28__SCAN_IN), .B1(n20146), 
        .B2(P1_UWORD_REG_12__SCAN_IN), .ZN(n12967) );
  NAND2_X1 U16051 ( .A1(n20142), .A2(n12967), .ZN(P1_U2949) );
  NAND2_X1 U16052 ( .A1(n20228), .A2(DATAI_6_), .ZN(n12969) );
  NAND2_X1 U16053 ( .A1(n20227), .A2(BUF1_REG_6__SCAN_IN), .ZN(n12968) );
  AND2_X1 U16054 ( .A1(n12969), .A2(n12968), .ZN(n20279) );
  INV_X1 U16055 ( .A(n20279), .ZN(n12970) );
  NAND2_X1 U16056 ( .A1(n13030), .A2(n12970), .ZN(n12992) );
  AOI22_X1 U16057 ( .A1(n20147), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n20146), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n12971) );
  NAND2_X1 U16058 ( .A1(n12992), .A2(n12971), .ZN(P1_U2958) );
  NAND2_X1 U16059 ( .A1(n20228), .A2(DATAI_0_), .ZN(n12973) );
  NAND2_X1 U16060 ( .A1(n20227), .A2(BUF1_REG_0__SCAN_IN), .ZN(n12972) );
  AND2_X1 U16061 ( .A1(n12973), .A2(n12972), .ZN(n20232) );
  INV_X1 U16062 ( .A(n20232), .ZN(n14385) );
  NAND2_X1 U16063 ( .A1(n13030), .A2(n14385), .ZN(n13001) );
  AOI22_X1 U16064 ( .A1(n20147), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n20146), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n12974) );
  NAND2_X1 U16065 ( .A1(n13001), .A2(n12974), .ZN(P1_U2937) );
  NAND2_X1 U16066 ( .A1(n20228), .A2(DATAI_5_), .ZN(n12976) );
  NAND2_X1 U16067 ( .A1(n20227), .A2(BUF1_REG_5__SCAN_IN), .ZN(n12975) );
  AND2_X1 U16068 ( .A1(n12976), .A2(n12975), .ZN(n20272) );
  INV_X1 U16069 ( .A(n20272), .ZN(n12977) );
  NAND2_X1 U16070 ( .A1(n13030), .A2(n12977), .ZN(n12999) );
  AOI22_X1 U16071 ( .A1(n20147), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n20146), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n12978) );
  NAND2_X1 U16072 ( .A1(n12999), .A2(n12978), .ZN(P1_U2942) );
  NAND2_X1 U16073 ( .A1(n20228), .A2(DATAI_1_), .ZN(n12980) );
  NAND2_X1 U16074 ( .A1(n20227), .A2(BUF1_REG_1__SCAN_IN), .ZN(n12979) );
  AND2_X1 U16075 ( .A1(n12980), .A2(n12979), .ZN(n20242) );
  INV_X1 U16076 ( .A(n20242), .ZN(n14380) );
  NAND2_X1 U16077 ( .A1(n13030), .A2(n14380), .ZN(n13009) );
  AOI22_X1 U16078 ( .A1(n20147), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n20146), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n12981) );
  NAND2_X1 U16079 ( .A1(n13009), .A2(n12981), .ZN(P1_U2953) );
  NAND2_X1 U16080 ( .A1(n20228), .A2(DATAI_3_), .ZN(n12983) );
  NAND2_X1 U16081 ( .A1(n20227), .A2(BUF1_REG_3__SCAN_IN), .ZN(n12982) );
  AND2_X1 U16082 ( .A1(n12983), .A2(n12982), .ZN(n20257) );
  INV_X1 U16083 ( .A(n20257), .ZN(n14373) );
  NAND2_X1 U16084 ( .A1(n13030), .A2(n14373), .ZN(n13007) );
  AOI22_X1 U16085 ( .A1(n20147), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n20146), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n12984) );
  NAND2_X1 U16086 ( .A1(n13007), .A2(n12984), .ZN(P1_U2940) );
  NAND2_X1 U16087 ( .A1(n20228), .A2(DATAI_4_), .ZN(n12986) );
  NAND2_X1 U16088 ( .A1(n20227), .A2(BUF1_REG_4__SCAN_IN), .ZN(n12985) );
  AND2_X1 U16089 ( .A1(n12986), .A2(n12985), .ZN(n20264) );
  INV_X1 U16090 ( .A(n20264), .ZN(n14370) );
  NAND2_X1 U16091 ( .A1(n13030), .A2(n14370), .ZN(n13005) );
  AOI22_X1 U16092 ( .A1(n20147), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n20146), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n12987) );
  NAND2_X1 U16093 ( .A1(n13005), .A2(n12987), .ZN(P1_U2941) );
  NAND2_X1 U16094 ( .A1(n20228), .A2(DATAI_7_), .ZN(n12989) );
  NAND2_X1 U16095 ( .A1(n20227), .A2(BUF1_REG_7__SCAN_IN), .ZN(n12988) );
  AND2_X1 U16096 ( .A1(n12989), .A2(n12988), .ZN(n20289) );
  INV_X1 U16097 ( .A(n20289), .ZN(n14352) );
  NAND2_X1 U16098 ( .A1(n13030), .A2(n14352), .ZN(n12994) );
  AOI22_X1 U16099 ( .A1(n20147), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n20146), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n12990) );
  NAND2_X1 U16100 ( .A1(n12994), .A2(n12990), .ZN(P1_U2944) );
  AOI22_X1 U16101 ( .A1(n20147), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n20146), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n12991) );
  NAND2_X1 U16102 ( .A1(n12992), .A2(n12991), .ZN(P1_U2943) );
  AOI22_X1 U16103 ( .A1(n20147), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n20146), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n12993) );
  NAND2_X1 U16104 ( .A1(n12994), .A2(n12993), .ZN(P1_U2959) );
  NAND2_X1 U16105 ( .A1(n20228), .A2(DATAI_2_), .ZN(n12996) );
  NAND2_X1 U16106 ( .A1(n20227), .A2(BUF1_REG_2__SCAN_IN), .ZN(n12995) );
  AND2_X1 U16107 ( .A1(n12996), .A2(n12995), .ZN(n20249) );
  INV_X1 U16108 ( .A(n20249), .ZN(n14376) );
  NAND2_X1 U16109 ( .A1(n13030), .A2(n14376), .ZN(n13003) );
  AOI22_X1 U16110 ( .A1(n20147), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n20146), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n12997) );
  NAND2_X1 U16111 ( .A1(n13003), .A2(n12997), .ZN(P1_U2954) );
  AOI22_X1 U16112 ( .A1(n20147), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n20146), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n12998) );
  NAND2_X1 U16113 ( .A1(n12999), .A2(n12998), .ZN(P1_U2957) );
  AOI22_X1 U16114 ( .A1(n20147), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n20146), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n13000) );
  NAND2_X1 U16115 ( .A1(n13001), .A2(n13000), .ZN(P1_U2952) );
  AOI22_X1 U16116 ( .A1(n20147), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n20146), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n13002) );
  NAND2_X1 U16117 ( .A1(n13003), .A2(n13002), .ZN(P1_U2939) );
  AOI22_X1 U16118 ( .A1(n20147), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20146), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n13004) );
  NAND2_X1 U16119 ( .A1(n13005), .A2(n13004), .ZN(P1_U2956) );
  AOI22_X1 U16120 ( .A1(n20147), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n20146), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n13006) );
  NAND2_X1 U16121 ( .A1(n13007), .A2(n13006), .ZN(P1_U2955) );
  AOI22_X1 U16122 ( .A1(n20147), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n20146), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13008) );
  NAND2_X1 U16123 ( .A1(n13009), .A2(n13008), .ZN(P1_U2938) );
  INV_X1 U16124 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n20975) );
  AOI22_X1 U16125 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20132), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n15908), .ZN(n13010) );
  OAI21_X1 U16126 ( .B1(n20975), .B2(n13017), .A(n13010), .ZN(P1_U2906) );
  INV_X1 U16127 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n21215) );
  AOI22_X1 U16128 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13011) );
  OAI21_X1 U16129 ( .B1(n21215), .B2(n13017), .A(n13011), .ZN(P1_U2910) );
  INV_X1 U16130 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13013) );
  AOI22_X1 U16131 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13012) );
  OAI21_X1 U16132 ( .B1(n13013), .B2(n13017), .A(n13012), .ZN(P1_U2919) );
  INV_X1 U16133 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13015) );
  AOI22_X1 U16134 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13014) );
  OAI21_X1 U16135 ( .B1(n13015), .B2(n13017), .A(n13014), .ZN(P1_U2920) );
  INV_X1 U16136 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13018) );
  AOI22_X1 U16137 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13016) );
  OAI21_X1 U16138 ( .B1(n13018), .B2(n13017), .A(n13016), .ZN(P1_U2918) );
  INV_X1 U16139 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14390) );
  INV_X1 U16140 ( .A(n13030), .ZN(n13022) );
  INV_X1 U16141 ( .A(DATAI_15_), .ZN(n13019) );
  NOR2_X1 U16142 ( .A1(n20227), .A2(n13019), .ZN(n13020) );
  AOI21_X1 U16143 ( .B1(n20227), .B2(BUF1_REG_15__SCAN_IN), .A(n13020), .ZN(
        n14392) );
  INV_X1 U16144 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20104) );
  OAI222_X1 U16145 ( .A1(n13034), .A2(n14390), .B1(n13022), .B2(n14392), .C1(
        n13021), .C2(n20104), .ZN(P1_U2967) );
  NOR2_X1 U16146 ( .A1(n20227), .A2(DATAI_9_), .ZN(n13023) );
  AOI21_X1 U16147 ( .B1(n20227), .B2(n12517), .A(n13023), .ZN(n14346) );
  NAND2_X1 U16148 ( .A1(n13030), .A2(n14346), .ZN(n20136) );
  NAND2_X1 U16149 ( .A1(n20146), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n13024) );
  OAI211_X1 U16150 ( .C1(n21279), .C2(n13034), .A(n20136), .B(n13024), .ZN(
        P1_U2946) );
  MUX2_X1 U16151 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n20227), .Z(
        n14406) );
  NAND2_X1 U16152 ( .A1(n13030), .A2(n14406), .ZN(n20140) );
  NAND2_X1 U16153 ( .A1(n20146), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n13025) );
  OAI211_X1 U16154 ( .C1(n13026), .C2(n13034), .A(n20140), .B(n13025), .ZN(
        P1_U2948) );
  INV_X1 U16155 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20119) );
  MUX2_X1 U16156 ( .A(DATAI_8_), .B(BUF1_REG_8__SCAN_IN), .S(n20227), .Z(
        n14349) );
  NAND2_X1 U16157 ( .A1(n13030), .A2(n14349), .ZN(n13033) );
  NAND2_X1 U16158 ( .A1(n20146), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n13027) );
  OAI211_X1 U16159 ( .C1(n20119), .C2(n13034), .A(n13033), .B(n13027), .ZN(
        P1_U2960) );
  MUX2_X1 U16160 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n20227), .Z(
        n14342) );
  NAND2_X1 U16161 ( .A1(n13030), .A2(n14342), .ZN(n20138) );
  NAND2_X1 U16162 ( .A1(n20146), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n13028) );
  OAI211_X1 U16163 ( .C1(n21215), .C2(n13034), .A(n20138), .B(n13028), .ZN(
        P1_U2947) );
  MUX2_X1 U16164 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n20227), .Z(
        n14395) );
  NAND2_X1 U16165 ( .A1(n13030), .A2(n14395), .ZN(n20148) );
  NAND2_X1 U16166 ( .A1(n20146), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13029) );
  OAI211_X1 U16167 ( .C1(n20975), .C2(n13034), .A(n20148), .B(n13029), .ZN(
        P1_U2951) );
  MUX2_X1 U16168 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n20227), .Z(
        n14398) );
  NAND2_X1 U16169 ( .A1(n13030), .A2(n14398), .ZN(n20144) );
  NAND2_X1 U16170 ( .A1(n20146), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n13031) );
  OAI211_X1 U16171 ( .C1(n20953), .C2(n13034), .A(n20144), .B(n13031), .ZN(
        P1_U2950) );
  NAND2_X1 U16172 ( .A1(n20146), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n13032) );
  OAI211_X1 U16173 ( .C1(n21187), .C2(n13034), .A(n13033), .B(n13032), .ZN(
        P1_U2945) );
  AND2_X1 U16174 ( .A1(n13036), .A2(n13035), .ZN(n13037) );
  OR2_X1 U16175 ( .A1(n13037), .A2(n9939), .ZN(n19072) );
  OAI211_X1 U16176 ( .C1(n9937), .C2(n13040), .A(n14901), .B(n13039), .ZN(
        n13042) );
  NAND2_X1 U16177 ( .A1(n14919), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13041) );
  OAI211_X1 U16178 ( .C1(n19072), .C2(n14919), .A(n13042), .B(n13041), .ZN(
        P2_U2879) );
  INV_X1 U16179 ( .A(n13043), .ZN(n13138) );
  XNOR2_X1 U16180 ( .A(n13039), .B(n13138), .ZN(n13047) );
  NOR2_X1 U16181 ( .A1(n9939), .A2(n13044), .ZN(n13045) );
  OR2_X1 U16182 ( .A1(n13143), .A2(n13045), .ZN(n15499) );
  MUX2_X1 U16183 ( .A(n11008), .B(n15499), .S(n14906), .Z(n13046) );
  OAI21_X1 U16184 ( .B1(n13047), .B2(n14921), .A(n13046), .ZN(P2_U2878) );
  MUX2_X1 U16185 ( .A(n14059), .B(n14082), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n13048) );
  OAI21_X1 U16186 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14071), .A(
        n13048), .ZN(n13049) );
  INV_X1 U16187 ( .A(n13049), .ZN(n13119) );
  NAND2_X1 U16188 ( .A1(n13120), .A2(n13119), .ZN(n13118) );
  MUX2_X1 U16189 ( .A(n14041), .B(n14046), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n13053) );
  INV_X1 U16190 ( .A(n13050), .ZN(n14056) );
  NAND2_X1 U16191 ( .A1(n14056), .A2(n14070), .ZN(n14015) );
  NAND2_X1 U16192 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n14070), .ZN(
        n13051) );
  AND2_X1 U16193 ( .A1(n14015), .A2(n13051), .ZN(n13052) );
  NAND2_X1 U16194 ( .A1(n13118), .A2(n13054), .ZN(n13055) );
  NAND2_X1 U16195 ( .A1(n16171), .A2(n13055), .ZN(n20172) );
  INV_X1 U16196 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n20058) );
  NAND2_X1 U16197 ( .A1(n13058), .A2(n13057), .ZN(n13059) );
  NAND2_X1 U16198 ( .A1(n13056), .A2(n13059), .ZN(n20156) );
  OAI222_X1 U16199 ( .A1(n20172), .A2(n14316), .B1(n20101), .B2(n20058), .C1(
        n14326), .C2(n20156), .ZN(P1_U2868) );
  NAND2_X1 U16200 ( .A1(n13060), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13061) );
  NAND2_X1 U16201 ( .A1(n13062), .A2(n13061), .ZN(n13325) );
  INV_X1 U16202 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20187) );
  XNOR2_X1 U16203 ( .A(n13325), .B(n20187), .ZN(n13072) );
  OR2_X1 U16204 ( .A1(n13063), .A2(n13064), .ZN(n13070) );
  NAND2_X1 U16205 ( .A1(n13066), .A2(n13065), .ZN(n13339) );
  INV_X1 U16206 ( .A(n13337), .ZN(n13067) );
  XNOR2_X1 U16207 ( .A(n13339), .B(n13067), .ZN(n13068) );
  NAND2_X1 U16208 ( .A1(n13068), .A2(n13488), .ZN(n13069) );
  NAND2_X1 U16209 ( .A1(n13070), .A2(n13069), .ZN(n13071) );
  NAND2_X1 U16210 ( .A1(n13072), .A2(n13071), .ZN(n13327) );
  OR2_X1 U16211 ( .A1(n13072), .A2(n13071), .ZN(n13073) );
  NAND2_X1 U16212 ( .A1(n13327), .A2(n13073), .ZN(n20182) );
  XOR2_X1 U16213 ( .A(n13074), .B(n13075), .Z(n13082) );
  NAND2_X1 U16214 ( .A1(n20150), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n20179) );
  NAND2_X1 U16215 ( .A1(n20151), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13076) );
  OAI211_X1 U16216 ( .C1(n20164), .C2(n14260), .A(n20179), .B(n13076), .ZN(
        n13077) );
  AOI21_X1 U16217 ( .B1(n13082), .B2(n20158), .A(n13077), .ZN(n13078) );
  OAI21_X1 U16218 ( .B1(n19988), .B2(n20182), .A(n13078), .ZN(P1_U2996) );
  NAND2_X1 U16219 ( .A1(n13080), .A2(n13079), .ZN(n13081) );
  INV_X1 U16220 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20131) );
  OAI222_X1 U16221 ( .A1(n20066), .A2(n14409), .B1(n14393), .B2(n20242), .C1(
        n14391), .C2(n20131), .ZN(P1_U2903) );
  INV_X1 U16222 ( .A(n13082), .ZN(n14266) );
  INV_X1 U16223 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20127) );
  OAI222_X1 U16224 ( .A1(n14266), .A2(n14409), .B1(n14393), .B2(n20257), .C1(
        n14391), .C2(n20127), .ZN(P1_U2901) );
  INV_X1 U16225 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20129) );
  OAI222_X1 U16226 ( .A1(n13083), .A2(n14409), .B1(n14393), .B2(n20249), .C1(
        n14391), .C2(n20129), .ZN(P1_U2902) );
  INV_X1 U16227 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20135) );
  OAI222_X1 U16228 ( .A1(n20086), .A2(n14409), .B1(n14393), .B2(n20232), .C1(
        n14391), .C2(n20135), .ZN(P1_U2904) );
  INV_X1 U16229 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20125) );
  OAI222_X1 U16230 ( .A1(n20156), .A2(n14409), .B1(n14393), .B2(n20264), .C1(
        n20125), .C2(n14391), .ZN(P1_U2900) );
  NOR2_X1 U16231 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n16192), .ZN(n13105) );
  INV_X1 U16232 ( .A(n20389), .ZN(n20630) );
  NOR2_X1 U16233 ( .A1(n11744), .A2(n20630), .ZN(n13084) );
  XNOR2_X1 U16234 ( .A(n13084), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20046) );
  NOR2_X1 U16235 ( .A1(n20046), .A2(n13085), .ZN(n16182) );
  OAI21_X1 U16236 ( .B1(n16182), .B2(n15853), .A(n16192), .ZN(n13086) );
  AOI21_X1 U16237 ( .B1(n15853), .B2(n16184), .A(n13086), .ZN(n13087) );
  AOI21_X1 U16238 ( .B1(n13105), .B2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n13087), .ZN(n15870) );
  MUX2_X1 U16239 ( .A(n13088), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15853), .Z(n15859) );
  AOI22_X1 U16240 ( .A1(n15859), .A2(n16192), .B1(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n13105), .ZN(n13107) );
  INV_X1 U16241 ( .A(n14731), .ZN(n13089) );
  NAND2_X1 U16242 ( .A1(n20500), .A2(n13089), .ZN(n13103) );
  AOI21_X1 U16243 ( .B1(n14735), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13090) );
  NOR2_X1 U16244 ( .A1(n13091), .A2(n13090), .ZN(n14742) );
  NAND3_X1 U16245 ( .A1(n14731), .A2(n13092), .A3(n14742), .ZN(n13101) );
  MUX2_X1 U16246 ( .A(n13093), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n14735), .Z(n13095) );
  NOR2_X1 U16247 ( .A1(n13095), .A2(n13094), .ZN(n13098) );
  XNOR2_X1 U16248 ( .A(n13096), .B(n11811), .ZN(n13097) );
  AOI22_X1 U16249 ( .A1(n13099), .A2(n13098), .B1(n14734), .B2(n13097), .ZN(
        n13100) );
  AND2_X1 U16250 ( .A1(n13101), .A2(n13100), .ZN(n13102) );
  NAND2_X1 U16251 ( .A1(n13103), .A2(n13102), .ZN(n14741) );
  INV_X1 U16252 ( .A(n15853), .ZN(n13104) );
  MUX2_X1 U16253 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14741), .S(
        n13104), .Z(n15862) );
  AOI22_X1 U16254 ( .A1(n13105), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n16192), .B2(n15862), .ZN(n13106) );
  NOR2_X1 U16255 ( .A1(n13107), .A2(n13106), .ZN(n15868) );
  INV_X1 U16256 ( .A(n11505), .ZN(n13108) );
  NAND2_X1 U16257 ( .A1(n15868), .A2(n13108), .ZN(n13112) );
  NAND3_X1 U16258 ( .A1(n15870), .A2(n21022), .A3(n13112), .ZN(n13111) );
  INV_X1 U16259 ( .A(n16193), .ZN(n13110) );
  INV_X1 U16260 ( .A(n20395), .ZN(n13109) );
  NAND3_X1 U16261 ( .A1(n15870), .A2(n13113), .A3(n13112), .ZN(n15884) );
  INV_X1 U16262 ( .A(n15884), .ZN(n13116) );
  INV_X1 U16263 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20641) );
  AND2_X1 U16264 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20641), .ZN(n14727) );
  OAI22_X1 U16265 ( .A1(n20323), .A2(n12580), .B1(n13114), .B2(n14727), .ZN(
        n13115) );
  OAI21_X1 U16266 ( .B1(n13116), .B2(n13115), .A(n20219), .ZN(n13117) );
  OAI21_X1 U16267 ( .B1(n20219), .B2(n20686), .A(n13117), .ZN(P1_U3478) );
  OAI21_X1 U16268 ( .B1(n13120), .B2(n13119), .A(n13118), .ZN(n20178) );
  INV_X1 U16269 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n21248) );
  OAI222_X1 U16270 ( .A1(n20178), .A2(n14316), .B1(n20101), .B2(n21248), .C1(
        n14326), .C2(n14266), .ZN(P1_U2869) );
  OR2_X1 U16271 ( .A1(n20769), .A2(n20766), .ZN(n20626) );
  NAND2_X1 U16272 ( .A1(n20627), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14721) );
  NOR2_X1 U16273 ( .A1(n20626), .A2(n14721), .ZN(n20690) );
  INV_X1 U16274 ( .A(n14721), .ZN(n13122) );
  NAND2_X1 U16275 ( .A1(n20766), .A2(n13122), .ZN(n14725) );
  NAND2_X1 U16276 ( .A1(n20598), .A2(n21280), .ZN(n20628) );
  INV_X1 U16277 ( .A(n20500), .ZN(n13124) );
  OAI22_X1 U16278 ( .A1(n13063), .A2(n20628), .B1(n13124), .B2(n14727), .ZN(
        n13125) );
  AOI21_X1 U16279 ( .B1(n20590), .B2(n20627), .A(n13125), .ZN(n13126) );
  OAI21_X1 U16280 ( .B1(n14725), .B2(n20471), .A(n13126), .ZN(n13127) );
  OAI21_X1 U16281 ( .B1(n20690), .B2(n13127), .A(n20219), .ZN(n13128) );
  OAI21_X1 U16282 ( .B1(n20219), .B2(n20634), .A(n13128), .ZN(P1_U3475) );
  XNOR2_X1 U16283 ( .A(n13129), .B(n13281), .ZN(n13133) );
  NAND2_X1 U16284 ( .A1(n13145), .A2(n13130), .ZN(n13131) );
  NAND2_X1 U16285 ( .A1(n13284), .A2(n13131), .ZN(n19049) );
  MUX2_X1 U16286 ( .A(n19041), .B(n19049), .S(n14906), .Z(n13132) );
  OAI21_X1 U16287 ( .B1(n13133), .B2(n14921), .A(n13132), .ZN(P2_U2876) );
  AND2_X1 U16288 ( .A1(n13056), .A2(n13135), .ZN(n13136) );
  OR2_X1 U16289 ( .A1(n13134), .A2(n13136), .ZN(n16052) );
  OAI222_X1 U16290 ( .A1(n16052), .A2(n14409), .B1(n14393), .B2(n20272), .C1(
        n13137), .C2(n14391), .ZN(P1_U2899) );
  NOR2_X1 U16291 ( .A1(n13039), .A2(n13138), .ZN(n13141) );
  INV_X1 U16292 ( .A(n13129), .ZN(n13139) );
  OAI211_X1 U16293 ( .C1(n13141), .C2(n13140), .A(n13139), .B(n14901), .ZN(
        n13147) );
  OR2_X1 U16294 ( .A1(n13143), .A2(n13142), .ZN(n13144) );
  NAND2_X1 U16295 ( .A1(n13145), .A2(n13144), .ZN(n15201) );
  INV_X1 U16296 ( .A(n15201), .ZN(n19061) );
  NAND2_X1 U16297 ( .A1(n19061), .A2(n14906), .ZN(n13146) );
  OAI211_X1 U16298 ( .C1(n14906), .C2(n19056), .A(n13147), .B(n13146), .ZN(
        P2_U2877) );
  NAND2_X1 U16299 ( .A1(n19522), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19405) );
  INV_X1 U16300 ( .A(n19405), .ZN(n19286) );
  NAND2_X1 U16301 ( .A1(n19286), .A2(n19753), .ZN(n19932) );
  NAND2_X1 U16302 ( .A1(n19691), .A2(n19935), .ZN(n19440) );
  NAND2_X1 U16303 ( .A1(n19932), .A2(n19440), .ZN(n13151) );
  NAND2_X1 U16304 ( .A1(n15525), .A2(n11122), .ZN(n13206) );
  NAND2_X1 U16305 ( .A1(n13579), .A2(n19938), .ZN(n13149) );
  NOR2_X1 U16306 ( .A1(n19964), .A2(n19440), .ZN(n19491) );
  NOR2_X1 U16307 ( .A1(n19923), .A2(n19491), .ZN(n13148) );
  AOI21_X1 U16308 ( .B1(n13149), .B2(n13148), .A(n19665), .ZN(n13150) );
  NAND2_X1 U16309 ( .A1(n13151), .A2(n13150), .ZN(n19484) );
  INV_X1 U16310 ( .A(n19484), .ZN(n19476) );
  OAI21_X1 U16311 ( .B1(n13579), .B2(n19491), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13152) );
  OAI21_X1 U16312 ( .B1(n19440), .B2(n19931), .A(n13152), .ZN(n19483) );
  NOR2_X2 U16313 ( .A1(n19159), .A2(n19665), .ZN(n19732) );
  NOR2_X2 U16314 ( .A1(n11101), .A2(n19266), .ZN(n19731) );
  INV_X1 U16315 ( .A(n19731), .ZN(n19802) );
  INV_X1 U16316 ( .A(n19491), .ZN(n13158) );
  INV_X1 U16317 ( .A(n19487), .ZN(n19473) );
  AOI22_X1 U16318 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19274), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19273), .ZN(n19808) );
  AOI22_X1 U16319 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19274), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19273), .ZN(n19654) );
  INV_X1 U16320 ( .A(n19654), .ZN(n19805) );
  AOI22_X1 U16321 ( .A1(n19473), .A2(n19651), .B1(n19516), .B2(n19805), .ZN(
        n13157) );
  OAI21_X1 U16322 ( .B1(n19802), .B2(n13158), .A(n13157), .ZN(n13159) );
  AOI21_X1 U16323 ( .B1(n19483), .B2(n19732), .A(n13159), .ZN(n13160) );
  OAI21_X1 U16324 ( .B1(n19476), .B2(n13161), .A(n13160), .ZN(P2_U3110) );
  OAI21_X1 U16325 ( .B1(n13134), .B2(n13164), .A(n13163), .ZN(n16044) );
  OAI222_X1 U16326 ( .A1(n16044), .A2(n14409), .B1(n14393), .B2(n20279), .C1(
        n20122), .C2(n14391), .ZN(P1_U2898) );
  XNOR2_X1 U16327 ( .A(n13165), .B(n13166), .ZN(n13529) );
  AOI21_X1 U16328 ( .B1(n19939), .B2(n19936), .A(n13167), .ZN(n19171) );
  XNOR2_X1 U16329 ( .A(n19522), .B(n13529), .ZN(n19172) );
  NOR2_X1 U16330 ( .A1(n19171), .A2(n19172), .ZN(n19170) );
  AOI21_X1 U16331 ( .B1(n13529), .B2(n19522), .A(n19170), .ZN(n13169) );
  XNOR2_X1 U16332 ( .A(n13168), .B(n9866), .ZN(n13553) );
  NOR2_X1 U16333 ( .A1(n13169), .A2(n13553), .ZN(n19165) );
  XNOR2_X1 U16334 ( .A(n19165), .B(n19164), .ZN(n13172) );
  AOI22_X1 U16335 ( .A1(n19177), .A2(n13553), .B1(n19176), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n13171) );
  NAND2_X1 U16336 ( .A1(n19162), .A2(n16233), .ZN(n13170) );
  OAI211_X1 U16337 ( .C1(n13172), .C2(n19181), .A(n13171), .B(n13170), .ZN(
        P2_U2915) );
  XNOR2_X1 U16338 ( .A(n13173), .B(n13294), .ZN(n13177) );
  OR2_X1 U16339 ( .A1(n13286), .A2(n13174), .ZN(n13175) );
  NAND2_X1 U16340 ( .A1(n13298), .A2(n13175), .ZN(n19024) );
  MUX2_X1 U16341 ( .A(n11022), .B(n19024), .S(n14906), .Z(n13176) );
  OAI21_X1 U16342 ( .B1(n13177), .B2(n14921), .A(n13176), .ZN(P2_U2874) );
  NAND2_X1 U16343 ( .A1(n14082), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13178) );
  OAI211_X1 U16344 ( .C1(n14070), .C2(P1_EBX_REG_5__SCAN_IN), .A(n14046), .B(
        n13178), .ZN(n13179) );
  OAI21_X1 U16345 ( .B1(n14059), .B2(P1_EBX_REG_5__SCAN_IN), .A(n13179), .ZN(
        n16170) );
  MUX2_X1 U16346 ( .A(n14041), .B(n14046), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n13182) );
  NAND2_X1 U16347 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14070), .ZN(
        n13180) );
  AND2_X1 U16348 ( .A1(n14015), .A2(n13180), .ZN(n13181) );
  NAND2_X1 U16349 ( .A1(n13182), .A2(n13181), .ZN(n13183) );
  NOR2_X1 U16350 ( .A1(n16173), .A2(n13183), .ZN(n13184) );
  OR2_X1 U16351 ( .A1(n16159), .A2(n13184), .ZN(n20028) );
  INV_X1 U16352 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n20948) );
  OAI222_X1 U16353 ( .A1(n20028), .A2(n14316), .B1(n20101), .B2(n20948), .C1(
        n14326), .C2(n16044), .ZN(P1_U2866) );
  INV_X1 U16354 ( .A(n13202), .ZN(n13193) );
  INV_X1 U16355 ( .A(n13588), .ZN(n13369) );
  AOI22_X1 U16356 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19443), .B1(
        n13369), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13197) );
  NAND2_X1 U16357 ( .A1(n13187), .A2(n15525), .ZN(n13204) );
  NAND2_X2 U16359 ( .A1(n21304), .A2(n13189), .ZN(n13357) );
  INV_X1 U16360 ( .A(n13357), .ZN(n13190) );
  AND2_X1 U16361 ( .A1(n13192), .A2(n13185), .ZN(n13205) );
  AOI22_X1 U16362 ( .A1(n19380), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n19624), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13195) );
  INV_X1 U16363 ( .A(n13206), .ZN(n13198) );
  AOI22_X1 U16364 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19747), .B1(
        n19700), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13194) );
  AND4_X2 U16365 ( .A1(n13197), .A2(n13196), .A3(n13195), .A4(n13194), .ZN(
        n13209) );
  AND2_X2 U16367 ( .A1(n21304), .A2(n13199), .ZN(n13365) );
  AOI21_X2 U16368 ( .B1(n13209), .B2(n13208), .A(n10358), .ZN(n13236) );
  INV_X1 U16369 ( .A(n13236), .ZN(n13234) );
  NAND2_X1 U16370 ( .A1(n13368), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n13210) );
  AOI22_X1 U16371 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19593), .B1(
        n19662), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13214) );
  AOI22_X1 U16372 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n13365), .B1(
        n19747), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13213) );
  AOI22_X1 U16373 ( .A1(n13356), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n19700), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13212) );
  NAND4_X1 U16374 ( .A1(n13215), .A2(n13214), .A3(n13213), .A4(n13212), .ZN(
        n13231) );
  AOI22_X1 U16375 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19380), .B1(
        n19443), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13225) );
  OAI21_X1 U16376 ( .B1(n13357), .B2(n13217), .A(n13216), .ZN(n13218) );
  INV_X1 U16377 ( .A(n13218), .ZN(n13220) );
  NAND2_X1 U16378 ( .A1(n19242), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13219) );
  INV_X1 U16379 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13221) );
  INV_X1 U16380 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n19573) );
  OAI22_X1 U16381 ( .A1(n13588), .A2(n13221), .B1(n13366), .B2(n19573), .ZN(
        n13222) );
  INV_X1 U16382 ( .A(n13222), .ZN(n13224) );
  AOI22_X1 U16383 ( .A1(n13579), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n19624), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13223) );
  NAND4_X1 U16384 ( .A1(n13225), .A2(n10373), .A3(n13224), .A4(n13223), .ZN(
        n13230) );
  NAND2_X1 U16385 ( .A1(n19247), .A2(n13226), .ZN(n13227) );
  OR2_X1 U16386 ( .A1(n13228), .A2(n13227), .ZN(n13261) );
  NAND2_X1 U16387 ( .A1(n13261), .A2(n13262), .ZN(n13229) );
  OAI21_X1 U16388 ( .B1(n13231), .B2(n13230), .A(n13229), .ZN(n13232) );
  INV_X1 U16389 ( .A(n13232), .ZN(n13235) );
  INV_X1 U16390 ( .A(n13235), .ZN(n13233) );
  NAND2_X1 U16391 ( .A1(n13236), .A2(n13235), .ZN(n13314) );
  INV_X1 U16392 ( .A(n13309), .ZN(n13240) );
  NAND2_X1 U16393 ( .A1(n13249), .A2(n13238), .ZN(n13239) );
  NAND2_X1 U16394 ( .A1(n13240), .A2(n13239), .ZN(n13528) );
  NAND2_X1 U16395 ( .A1(n13242), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13306) );
  NAND2_X1 U16396 ( .A1(n13307), .A2(n13306), .ZN(n13252) );
  NOR2_X1 U16397 ( .A1(n13243), .A2(n14807), .ZN(n13245) );
  OAI21_X1 U16398 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13245), .A(
        n13244), .ZN(n13790) );
  OR2_X1 U16399 ( .A1(n13247), .A2(n13246), .ZN(n13248) );
  NAND2_X1 U16400 ( .A1(n13249), .A2(n13248), .ZN(n13540) );
  XNOR2_X1 U16401 ( .A(n13540), .B(n13784), .ZN(n13789) );
  OR2_X1 U16402 ( .A1(n13790), .A2(n13789), .ZN(n13808) );
  INV_X1 U16403 ( .A(n13540), .ZN(n13250) );
  NAND2_X1 U16404 ( .A1(n13250), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13251) );
  AND2_X1 U16405 ( .A1(n13808), .A2(n13251), .ZN(n13305) );
  XNOR2_X1 U16406 ( .A(n13252), .B(n13305), .ZN(n13279) );
  INV_X1 U16407 ( .A(n13529), .ZN(n19927) );
  OAI22_X1 U16408 ( .A1(n13253), .A2(n16314), .B1(n13272), .B2(n19083), .ZN(
        n13260) );
  INV_X1 U16409 ( .A(n15374), .ZN(n13256) );
  NAND2_X1 U16410 ( .A1(n13784), .A2(n13254), .ZN(n13961) );
  NAND3_X1 U16411 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13785) );
  INV_X1 U16412 ( .A(n13785), .ZN(n13255) );
  AOI21_X1 U16413 ( .B1(n13256), .B2(n13961), .A(n13255), .ZN(n13319) );
  NAND2_X1 U16414 ( .A1(n13619), .A2(n16318), .ZN(n13258) );
  NOR2_X1 U16415 ( .A1(n15374), .A2(n13961), .ZN(n13799) );
  INV_X1 U16416 ( .A(n15377), .ZN(n13257) );
  NAND2_X1 U16417 ( .A1(n13257), .A2(n13785), .ZN(n13794) );
  NAND2_X1 U16418 ( .A1(n16316), .A2(n13794), .ZN(n13964) );
  NOR2_X1 U16419 ( .A1(n13799), .A2(n13964), .ZN(n13624) );
  OAI22_X1 U16420 ( .A1(n13319), .A2(n13258), .B1(n13624), .B2(n13619), .ZN(
        n13259) );
  AOI211_X1 U16421 ( .C1(n16299), .C2(n19927), .A(n13260), .B(n13259), .ZN(
        n13271) );
  XOR2_X1 U16422 ( .A(n13262), .B(n13261), .Z(n13788) );
  NOR2_X1 U16423 ( .A1(n13264), .A2(n13263), .ZN(n13266) );
  NOR2_X1 U16424 ( .A1(n13266), .A2(n13265), .ZN(n13267) );
  XOR2_X1 U16425 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n13267), .Z(
        n13787) );
  NOR2_X1 U16426 ( .A1(n13788), .A2(n13787), .ZN(n13786) );
  NOR2_X1 U16427 ( .A1(n13267), .A2(n13784), .ZN(n13268) );
  OR2_X1 U16428 ( .A1(n13786), .A2(n13268), .ZN(n13310) );
  XNOR2_X1 U16429 ( .A(n13310), .B(n13619), .ZN(n13269) );
  NAND3_X1 U16430 ( .A1(n13276), .A2(n16301), .A3(n13312), .ZN(n13270) );
  OAI211_X1 U16431 ( .C1(n13279), .C2(n15495), .A(n13271), .B(n13270), .ZN(
        P2_U3043) );
  NOR2_X1 U16432 ( .A1(n19040), .A2(n13272), .ZN(n13275) );
  INV_X1 U16433 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13273) );
  OAI22_X1 U16434 ( .A1(n13273), .A2(n19234), .B1(n15211), .B2(n13523), .ZN(
        n13274) );
  AOI211_X1 U16435 ( .C1(n19231), .C2(n13532), .A(n13275), .B(n13274), .ZN(
        n13278) );
  NAND3_X1 U16436 ( .A1(n13276), .A2(n16283), .A3(n13312), .ZN(n13277) );
  OAI211_X1 U16437 ( .C1(n13279), .C2(n19227), .A(n13278), .B(n13277), .ZN(
        P2_U3011) );
  AOI21_X1 U16438 ( .B1(n13129), .B2(n13281), .A(n13280), .ZN(n13282) );
  OR3_X1 U16439 ( .A1(n13173), .A2(n13282), .A3(n14921), .ZN(n13288) );
  AND2_X1 U16440 ( .A1(n13284), .A2(n13283), .ZN(n13285) );
  OR2_X1 U16441 ( .A1(n13286), .A2(n13285), .ZN(n15454) );
  INV_X1 U16442 ( .A(n15454), .ZN(n19035) );
  NAND2_X1 U16443 ( .A1(n19035), .A2(n14906), .ZN(n13287) );
  OAI211_X1 U16444 ( .C1(n14906), .C2(n11019), .A(n13288), .B(n13287), .ZN(
        P2_U2875) );
  NAND2_X1 U16445 ( .A1(n13163), .A2(n13290), .ZN(n13291) );
  AND2_X1 U16446 ( .A1(n13289), .A2(n13291), .ZN(n20094) );
  INV_X1 U16447 ( .A(n20094), .ZN(n13293) );
  OAI222_X1 U16448 ( .A1(n13293), .A2(n14409), .B1(n14393), .B2(n20289), .C1(
        n13292), .C2(n14391), .ZN(P1_U2897) );
  AND2_X1 U16449 ( .A1(n13173), .A2(n13294), .ZN(n13297) );
  OAI211_X1 U16450 ( .C1(n13297), .C2(n13296), .A(n14901), .B(n13295), .ZN(
        n13304) );
  INV_X1 U16451 ( .A(n13298), .ZN(n13302) );
  INV_X1 U16452 ( .A(n13299), .ZN(n13301) );
  OAI21_X1 U16453 ( .B1(n13302), .B2(n13301), .A(n13419), .ZN(n15423) );
  INV_X1 U16454 ( .A(n15423), .ZN(n19012) );
  NAND2_X1 U16455 ( .A1(n19012), .A2(n14906), .ZN(n13303) );
  OAI211_X1 U16456 ( .C1(n14906), .C2(n13866), .A(n13304), .B(n13303), .ZN(
        P2_U2873) );
  OAI21_X1 U16457 ( .B1(n13309), .B2(n13308), .A(n13381), .ZN(n13555) );
  INV_X1 U16458 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13620) );
  XNOR2_X1 U16459 ( .A(n13555), .B(n13620), .ZN(n13385) );
  XOR2_X1 U16460 ( .A(n13384), .B(n13385), .Z(n19224) );
  NAND2_X1 U16461 ( .A1(n13310), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13311) );
  INV_X1 U16462 ( .A(n13314), .ZN(n13313) );
  INV_X1 U16463 ( .A(n13315), .ZN(n13316) );
  NAND2_X1 U16464 ( .A1(n13314), .A2(n13316), .ZN(n13317) );
  NAND2_X1 U16465 ( .A1(n13379), .A2(n13317), .ZN(n13390) );
  XNOR2_X1 U16466 ( .A(n13390), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13318) );
  XNOR2_X1 U16467 ( .A(n13392), .B(n13318), .ZN(n19226) );
  NOR2_X1 U16468 ( .A1(n15381), .A2(n13319), .ZN(n13621) );
  AND2_X1 U16469 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13621), .ZN(
        n13408) );
  OAI21_X1 U16470 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n15381), .A(
        n13624), .ZN(n13407) );
  INV_X1 U16471 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n19862) );
  NOR2_X1 U16472 ( .A1(n19862), .A2(n19040), .ZN(n13320) );
  AOI221_X1 U16473 ( .B1(n13408), .B2(n13620), .C1(n13407), .C2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n13320), .ZN(n13322) );
  AOI22_X1 U16474 ( .A1(n19230), .A2(n16304), .B1(n16299), .B2(n13553), .ZN(
        n13321) );
  OAI211_X1 U16475 ( .C1(n19226), .C2(n16326), .A(n13322), .B(n13321), .ZN(
        n13323) );
  AOI21_X1 U16476 ( .B1(n19224), .B2(n16322), .A(n13323), .ZN(n13324) );
  INV_X1 U16477 ( .A(n13324), .ZN(P2_U3042) );
  NAND2_X1 U16478 ( .A1(n13325), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13326) );
  NAND2_X1 U16479 ( .A1(n13327), .A2(n13326), .ZN(n20153) );
  NAND2_X1 U16480 ( .A1(n13328), .A2(n13494), .ZN(n13332) );
  NAND2_X1 U16481 ( .A1(n13339), .A2(n13337), .ZN(n13329) );
  XNOR2_X1 U16482 ( .A(n13329), .B(n13336), .ZN(n13330) );
  NAND2_X1 U16483 ( .A1(n13330), .A2(n13488), .ZN(n13331) );
  NAND2_X1 U16484 ( .A1(n13332), .A2(n13331), .ZN(n13333) );
  INV_X1 U16485 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20177) );
  XNOR2_X1 U16486 ( .A(n13333), .B(n20177), .ZN(n20152) );
  NAND2_X1 U16487 ( .A1(n20153), .A2(n20152), .ZN(n20155) );
  NAND2_X1 U16488 ( .A1(n13333), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13334) );
  AND2_X1 U16489 ( .A1(n13337), .A2(n13336), .ZN(n13338) );
  NAND2_X1 U16490 ( .A1(n13339), .A2(n13338), .ZN(n13344) );
  XNOR2_X1 U16491 ( .A(n13344), .B(n13345), .ZN(n13340) );
  NAND2_X1 U16492 ( .A1(n13340), .A2(n13488), .ZN(n13341) );
  INV_X1 U16493 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14578) );
  XNOR2_X1 U16494 ( .A(n13342), .B(n14578), .ZN(n16049) );
  NAND3_X1 U16495 ( .A1(n13497), .A2(n13343), .A3(n13494), .ZN(n13349) );
  INV_X1 U16496 ( .A(n13344), .ZN(n13346) );
  NAND2_X1 U16497 ( .A1(n13346), .A2(n13345), .ZN(n13484) );
  XNOR2_X1 U16498 ( .A(n13484), .B(n13485), .ZN(n13347) );
  NAND2_X1 U16499 ( .A1(n13347), .A2(n13488), .ZN(n13348) );
  NAND2_X1 U16500 ( .A1(n13349), .A2(n13348), .ZN(n13481) );
  XOR2_X1 U16501 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n13481), .Z(
        n13350) );
  XNOR2_X1 U16502 ( .A(n13480), .B(n13350), .ZN(n16043) );
  NOR2_X1 U16503 ( .A1(n20177), .A2(n20187), .ZN(n20169) );
  INV_X1 U16504 ( .A(n20169), .ZN(n13351) );
  OAI21_X1 U16505 ( .B1(n20190), .B2(n20217), .A(n20203), .ZN(n20194) );
  NAND2_X1 U16506 ( .A1(n16117), .A2(n14680), .ZN(n14705) );
  NAND2_X1 U16507 ( .A1(n20190), .A2(n16117), .ZN(n20205) );
  NAND2_X1 U16508 ( .A1(n14705), .A2(n20205), .ZN(n14708) );
  NOR2_X1 U16509 ( .A1(n20217), .A2(n14708), .ZN(n20189) );
  NAND2_X1 U16510 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n20189), .ZN(
        n13352) );
  NAND2_X1 U16511 ( .A1(n20195), .A2(n13352), .ZN(n16108) );
  NAND2_X1 U16512 ( .A1(n20194), .A2(n16108), .ZN(n20183) );
  NOR3_X1 U16513 ( .A1(n14578), .A2(n13351), .A3(n20183), .ZN(n14714) );
  INV_X1 U16514 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13508) );
  NAND2_X1 U16515 ( .A1(n14714), .A2(n13508), .ZN(n13355) );
  NAND2_X1 U16516 ( .A1(n20169), .A2(n14578), .ZN(n16179) );
  NAND3_X1 U16517 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n20169), .ZN(n14577) );
  INV_X1 U16518 ( .A(n20194), .ZN(n20168) );
  NOR3_X1 U16519 ( .A1(n20168), .A2(n13351), .A3(n14578), .ZN(n14579) );
  INV_X1 U16520 ( .A(n14696), .ZN(n20165) );
  OAI21_X1 U16521 ( .B1(n14579), .B2(n20195), .A(n20165), .ZN(n16138) );
  AOI21_X1 U16522 ( .B1(n14705), .B2(n14577), .A(n16138), .ZN(n16174) );
  OAI21_X1 U16523 ( .B1(n13352), .B2(n16179), .A(n16174), .ZN(n13507) );
  INV_X1 U16524 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21235) );
  OAI22_X1 U16525 ( .A1(n20028), .A2(n20171), .B1(n21235), .B2(n20207), .ZN(
        n13353) );
  AOI21_X1 U16526 ( .B1(n13507), .B2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n13353), .ZN(n13354) );
  OAI211_X1 U16527 ( .C1(n16043), .C2(n20196), .A(n13355), .B(n13354), .ZN(
        P1_U3025) );
  AOI22_X1 U16528 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n13356), .B1(
        n13579), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13364) );
  AOI22_X1 U16529 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19593), .B1(
        n19662), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13363) );
  AOI22_X1 U16530 ( .A1(n19443), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n19700), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13362) );
  INV_X1 U16531 ( .A(n19624), .ZN(n19630) );
  INV_X1 U16532 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13358) );
  OAI22_X1 U16533 ( .A1(n13359), .A2(n13357), .B1(n19630), .B2(n13358), .ZN(
        n13360) );
  INV_X1 U16534 ( .A(n13360), .ZN(n13361) );
  NAND4_X1 U16535 ( .A1(n13364), .A2(n13363), .A3(n13362), .A4(n13361), .ZN(
        n13375) );
  AOI22_X1 U16536 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n13365), .B1(
        n19242), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13373) );
  AOI22_X1 U16537 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19566), .B1(
        n13367), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13372) );
  AOI22_X1 U16538 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19380), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13371) );
  AOI22_X1 U16539 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n13369), .B1(
        n19747), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13370) );
  NAND4_X1 U16540 ( .A1(n13373), .A2(n13372), .A3(n13371), .A4(n13370), .ZN(
        n13374) );
  NAND2_X1 U16541 ( .A1(n13376), .A2(n19247), .ZN(n13377) );
  INV_X1 U16542 ( .A(n13614), .ZN(n13383) );
  NAND2_X1 U16543 ( .A1(n13381), .A2(n13380), .ZN(n13382) );
  NAND2_X1 U16544 ( .A1(n13383), .A2(n13382), .ZN(n19107) );
  INV_X1 U16545 ( .A(n13385), .ZN(n13386) );
  INV_X1 U16546 ( .A(n13555), .ZN(n13387) );
  NAND2_X1 U16547 ( .A1(n13387), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13388) );
  NAND2_X1 U16548 ( .A1(n13389), .A2(n13388), .ZN(n13609) );
  XNOR2_X1 U16549 ( .A(n13610), .B(n13609), .ZN(n13461) );
  NAND2_X1 U16550 ( .A1(n13391), .A2(n13390), .ZN(n13395) );
  INV_X1 U16551 ( .A(n13392), .ZN(n13393) );
  NAND2_X1 U16552 ( .A1(n13393), .A2(n13620), .ZN(n13394) );
  NAND2_X1 U16553 ( .A1(n13396), .A2(n13618), .ZN(n13398) );
  INV_X1 U16554 ( .A(n13604), .ZN(n13400) );
  AOI21_X1 U16555 ( .B1(n13606), .B2(n13398), .A(n13397), .ZN(n13399) );
  AOI21_X1 U16556 ( .B1(n13400), .B2(n13606), .A(n13399), .ZN(n13459) );
  OAI21_X1 U16557 ( .B1(n13403), .B2(n13402), .A(n13401), .ZN(n19168) );
  INV_X1 U16558 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n13404) );
  OR2_X1 U16559 ( .A1(n19040), .A2(n13404), .ZN(n13456) );
  INV_X1 U16560 ( .A(n13456), .ZN(n13406) );
  NOR2_X1 U16561 ( .A1(n16314), .A2(n19114), .ZN(n13405) );
  AOI211_X1 U16562 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n13407), .A(
        n13406), .B(n13405), .ZN(n13410) );
  OAI221_X1 U16563 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C1(n13620), .C2(n13618), .A(
        n13408), .ZN(n13409) );
  OAI211_X1 U16564 ( .C1(n19168), .C2(n16313), .A(n13410), .B(n13409), .ZN(
        n13411) );
  AOI21_X1 U16565 ( .B1(n13459), .B2(n16301), .A(n13411), .ZN(n13412) );
  OAI21_X1 U16566 ( .B1(n15495), .B2(n13461), .A(n13412), .ZN(P2_U3041) );
  INV_X1 U16567 ( .A(n13413), .ZN(n13414) );
  AOI21_X1 U16568 ( .B1(n13415), .B2(n13289), .A(n13414), .ZN(n13519) );
  INV_X1 U16569 ( .A(n13519), .ZN(n13462) );
  AOI22_X1 U16570 ( .A1(n14407), .A2(n14349), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n14405), .ZN(n13416) );
  OAI21_X1 U16571 ( .B1(n13462), .B2(n14409), .A(n13416), .ZN(P1_U2896) );
  XNOR2_X1 U16572 ( .A(n13295), .B(n13417), .ZN(n13422) );
  NAND2_X1 U16573 ( .A1(n13419), .A2(n13418), .ZN(n13420) );
  AND2_X1 U16574 ( .A1(n14917), .A2(n13420), .ZN(n16245) );
  INV_X1 U16575 ( .A(n16245), .ZN(n19001) );
  MUX2_X1 U16576 ( .A(n19001), .B(n11029), .S(n14919), .Z(n13421) );
  OAI21_X1 U16577 ( .B1(n13422), .B2(n14921), .A(n13421), .ZN(P2_U2872) );
  NAND2_X1 U16578 ( .A1(n20898), .A2(n16192), .ZN(n20901) );
  OR2_X1 U16579 ( .A1(n20641), .A2(n20901), .ZN(n15877) );
  NOR2_X1 U16580 ( .A1(n15877), .A2(n20902), .ZN(n13428) );
  NAND2_X1 U16581 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20902), .ZN(n13426) );
  OAI21_X1 U16582 ( .B1(n13426), .B2(n13425), .A(n20207), .ZN(n13427) );
  NAND2_X1 U16583 ( .A1(n13429), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13430) );
  INV_X1 U16584 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14076) );
  XNOR2_X1 U16585 ( .A(n13430), .B(n14076), .ZN(n14431) );
  NOR2_X1 U16586 ( .A1(n14431), .A2(n16192), .ZN(n13431) );
  INV_X1 U16587 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n21208) );
  NAND4_X1 U16588 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n20020)
         );
  NAND3_X1 U16589 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n20003) );
  NOR3_X1 U16590 ( .A1(n21208), .A2(n20020), .A3(n20003), .ZN(n13563) );
  NOR2_X1 U16591 ( .A1(n13432), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13448) );
  OAI21_X1 U16592 ( .B1(n13563), .B2(n20021), .A(n20059), .ZN(n20005) );
  NOR2_X1 U16593 ( .A1(n20003), .A2(n20038), .ZN(n13433) );
  AOI22_X1 U16594 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20005), .B1(n13433), 
        .B2(n21208), .ZN(n13455) );
  AND2_X1 U16595 ( .A1(n14431), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13434) );
  INV_X1 U16596 ( .A(n13517), .ZN(n13453) );
  NOR2_X2 U16597 ( .A1(n20019), .A2(n19985), .ZN(n20048) );
  NAND2_X1 U16598 ( .A1(n13435), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13446) );
  AND2_X1 U16599 ( .A1(n20906), .A2(n21280), .ZN(n13436) );
  NOR2_X1 U16600 ( .A1(n13446), .A2(n13436), .ZN(n13437) );
  INV_X1 U16601 ( .A(n14059), .ZN(n14044) );
  INV_X1 U16602 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n21201) );
  NAND2_X1 U16603 ( .A1(n14044), .A2(n21201), .ZN(n13440) );
  NAND2_X1 U16604 ( .A1(n14082), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13438) );
  OAI211_X1 U16605 ( .C1(n14070), .C2(P1_EBX_REG_7__SCAN_IN), .A(n14046), .B(
        n13438), .ZN(n13439) );
  AND2_X1 U16606 ( .A1(n13440), .A2(n13439), .ZN(n16158) );
  MUX2_X1 U16607 ( .A(n14041), .B(n14046), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n13443) );
  NAND2_X1 U16608 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n14070), .ZN(
        n13441) );
  AND2_X1 U16609 ( .A1(n14015), .A2(n13441), .ZN(n13442) );
  NAND2_X1 U16610 ( .A1(n16161), .A2(n13444), .ZN(n13445) );
  NAND2_X1 U16611 ( .A1(n16148), .A2(n13445), .ZN(n13505) );
  INV_X1 U16612 ( .A(n13446), .ZN(n13447) );
  NOR2_X1 U16613 ( .A1(n13448), .A2(n13447), .ZN(n13449) );
  AOI22_X1 U16614 ( .A1(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n20080), .B1(
        P1_EBX_REG_8__SCAN_IN), .B2(n20075), .ZN(n13451) );
  OAI21_X1 U16615 ( .B1(n20073), .B2(n13505), .A(n13451), .ZN(n13452) );
  AOI211_X1 U16616 ( .C1(n20079), .C2(n13453), .A(n20048), .B(n13452), .ZN(
        n13454) );
  OAI211_X1 U16617 ( .C1(n13462), .C2(n15937), .A(n13455), .B(n13454), .ZN(
        P1_U2832) );
  INV_X1 U16618 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19104) );
  OAI22_X1 U16619 ( .A1(n19104), .A2(n19234), .B1(n15211), .B2(n19113), .ZN(
        n13458) );
  OAI21_X1 U16620 ( .B1(n13154), .B2(n19114), .A(n13456), .ZN(n13457) );
  AOI211_X1 U16621 ( .C1(n13459), .C2(n16283), .A(n13458), .B(n13457), .ZN(
        n13460) );
  OAI21_X1 U16622 ( .B1(n19227), .B2(n13461), .A(n13460), .ZN(P2_U3009) );
  INV_X1 U16623 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13463) );
  OAI222_X1 U16624 ( .A1(n13505), .A2(n14316), .B1(n20101), .B2(n13463), .C1(
        n14326), .C2(n13462), .ZN(P1_U2864) );
  OR2_X1 U16625 ( .A1(n13465), .A2(n13466), .ZN(n13467) );
  NAND2_X1 U16626 ( .A1(n13464), .A2(n13467), .ZN(n14912) );
  OAI21_X1 U16627 ( .B1(n15394), .B2(n13468), .A(n9870), .ZN(n18977) );
  INV_X1 U16628 ( .A(n19177), .ZN(n19131) );
  OAI22_X1 U16629 ( .A1(n14988), .A2(n19248), .B1(n19160), .B2(n13469), .ZN(
        n13470) );
  AOI21_X1 U16630 ( .B1(n19129), .B2(BUF1_REG_17__SCAN_IN), .A(n13470), .ZN(
        n13472) );
  NAND2_X1 U16631 ( .A1(n19128), .A2(BUF2_REG_17__SCAN_IN), .ZN(n13471) );
  OAI211_X1 U16632 ( .C1(n18977), .C2(n19131), .A(n13472), .B(n13471), .ZN(
        n13473) );
  INV_X1 U16633 ( .A(n13473), .ZN(n13474) );
  OAI21_X1 U16634 ( .B1(n19181), .B2(n14912), .A(n13474), .ZN(P2_U2902) );
  AND2_X1 U16635 ( .A1(n13413), .A2(n13475), .ZN(n13478) );
  OR2_X1 U16636 ( .A1(n13478), .A2(n13477), .ZN(n20089) );
  AOI22_X1 U16637 ( .A1(n14407), .A2(n14346), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n14405), .ZN(n13479) );
  OAI21_X1 U16638 ( .B1(n20089), .B2(n14409), .A(n13479), .ZN(P1_U2895) );
  NAND2_X1 U16639 ( .A1(n13481), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13482) );
  NAND2_X1 U16640 ( .A1(n13483), .A2(n13494), .ZN(n13491) );
  INV_X1 U16641 ( .A(n13484), .ZN(n13486) );
  NAND2_X1 U16642 ( .A1(n13486), .A2(n13485), .ZN(n13500) );
  XNOR2_X1 U16643 ( .A(n13500), .B(n13487), .ZN(n13489) );
  NAND2_X1 U16644 ( .A1(n13489), .A2(n13488), .ZN(n13490) );
  NAND2_X1 U16645 ( .A1(n13491), .A2(n13490), .ZN(n13492) );
  XNOR2_X1 U16646 ( .A(n13492), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16036) );
  OR2_X1 U16647 ( .A1(n13492), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13493) );
  AND2_X1 U16648 ( .A1(n13495), .A2(n13494), .ZN(n13496) );
  OR3_X1 U16649 ( .A1(n13500), .A2(n13499), .A3(n15872), .ZN(n13501) );
  NAND2_X1 U16650 ( .A1(n13498), .A2(n13501), .ZN(n13502) );
  NOR2_X1 U16651 ( .A1(n13502), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13632) );
  INV_X1 U16652 ( .A(n13632), .ZN(n13503) );
  NAND2_X1 U16653 ( .A1(n13502), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13631) );
  NAND2_X1 U16654 ( .A1(n13503), .A2(n13631), .ZN(n13504) );
  XNOR2_X1 U16655 ( .A(n13633), .B(n13504), .ZN(n13521) );
  INV_X1 U16656 ( .A(n13505), .ZN(n13513) );
  NAND2_X1 U16657 ( .A1(n20150), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n13516) );
  INV_X1 U16658 ( .A(n13516), .ZN(n13512) );
  AOI21_X1 U16659 ( .B1(n13508), .B2(n20206), .A(n13507), .ZN(n16169) );
  INV_X1 U16660 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n13510) );
  NAND2_X1 U16661 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14714), .ZN(
        n16163) );
  NAND2_X1 U16662 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16130) );
  OAI21_X1 U16663 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16130), .ZN(n13509) );
  OAI22_X1 U16664 ( .A1(n16169), .A2(n13510), .B1(n16163), .B2(n13509), .ZN(
        n13511) );
  AOI211_X1 U16665 ( .C1(n20214), .C2(n13513), .A(n13512), .B(n13511), .ZN(
        n13514) );
  OAI21_X1 U16666 ( .B1(n13521), .B2(n20196), .A(n13514), .ZN(P1_U3023) );
  NAND2_X1 U16667 ( .A1(n20151), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13515) );
  OAI211_X1 U16668 ( .C1(n20164), .C2(n13517), .A(n13516), .B(n13515), .ZN(
        n13518) );
  AOI21_X1 U16669 ( .B1(n13519), .B2(n20158), .A(n13518), .ZN(n13520) );
  OAI21_X1 U16670 ( .B1(n13521), .B2(n19988), .A(n13520), .ZN(P1_U2991) );
  NOR2_X1 U16671 ( .A1(n10145), .A2(n13522), .ZN(n13524) );
  XNOR2_X1 U16672 ( .A(n13524), .B(n13523), .ZN(n13525) );
  INV_X1 U16673 ( .A(n19831), .ZN(n19118) );
  NAND2_X1 U16674 ( .A1(n13525), .A2(n19118), .ZN(n13534) );
  OAI22_X1 U16675 ( .A1(n13272), .A2(n19122), .B1(n10979), .B2(n19085), .ZN(
        n13526) );
  AOI21_X1 U16676 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n19089), .A(
        n13526), .ZN(n13527) );
  OAI21_X1 U16677 ( .B1(n13528), .B2(n19106), .A(n13527), .ZN(n13531) );
  NOR2_X1 U16678 ( .A1(n13529), .A2(n19116), .ZN(n13530) );
  AOI211_X1 U16679 ( .C1(n11089), .C2(n13532), .A(n13531), .B(n13530), .ZN(
        n13533) );
  OAI211_X1 U16680 ( .C1(n14824), .C2(n19522), .A(n13534), .B(n13533), .ZN(
        P2_U2852) );
  NAND2_X1 U16681 ( .A1(n13535), .A2(n14804), .ZN(n13536) );
  XNOR2_X1 U16682 ( .A(n13806), .B(n13536), .ZN(n13546) );
  OAI22_X1 U16683 ( .A1(n19860), .A2(n19122), .B1(n13537), .B2(n19085), .ZN(
        n13538) );
  AOI21_X1 U16684 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19089), .A(
        n13538), .ZN(n13539) );
  OAI21_X1 U16685 ( .B1(n19106), .B2(n13540), .A(n13539), .ZN(n13541) );
  AOI21_X1 U16686 ( .B1(n13798), .B2(n19036), .A(n13541), .ZN(n13544) );
  NAND2_X1 U16687 ( .A1(n13542), .A2(n11089), .ZN(n13543) );
  OAI211_X1 U16688 ( .C1(n19936), .C2(n14824), .A(n13544), .B(n13543), .ZN(
        n13545) );
  AOI21_X1 U16689 ( .B1(n13546), .B2(n19118), .A(n13545), .ZN(n13547) );
  INV_X1 U16690 ( .A(n13547), .ZN(P2_U2853) );
  AND2_X1 U16691 ( .A1(n13535), .A2(n13548), .ZN(n13550) );
  AOI21_X1 U16692 ( .B1(n19221), .B2(n13550), .A(n19831), .ZN(n13549) );
  OAI21_X1 U16693 ( .B1(n19221), .B2(n13550), .A(n13549), .ZN(n13558) );
  AOI22_X1 U16694 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19080), .B1(
        P2_EBX_REG_4__SCAN_IN), .B2(n19109), .ZN(n13551) );
  OAI211_X1 U16695 ( .C1(n19105), .C2(n19235), .A(n19083), .B(n13551), .ZN(
        n13552) );
  AOI21_X1 U16696 ( .B1(n19036), .B2(n13553), .A(n13552), .ZN(n13554) );
  OAI21_X1 U16697 ( .B1(n13555), .B2(n19106), .A(n13554), .ZN(n13556) );
  AOI21_X1 U16698 ( .B1(n19230), .B2(n11089), .A(n13556), .ZN(n13557) );
  OAI211_X1 U16699 ( .C1(n19164), .C2(n14824), .A(n13558), .B(n13557), .ZN(
        P2_U2851) );
  INV_X1 U16700 ( .A(n13559), .ZN(n13562) );
  INV_X1 U16701 ( .A(n13477), .ZN(n13561) );
  AOI21_X1 U16702 ( .B1(n13562), .B2(n13561), .A(n13560), .ZN(n14574) );
  INV_X1 U16703 ( .A(n14574), .ZN(n13630) );
  INV_X1 U16704 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n21026) );
  NAND2_X1 U16705 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n13563), .ZN(n13572) );
  NOR2_X1 U16706 ( .A1(n21026), .A2(n13572), .ZN(n14205) );
  OAI21_X1 U16707 ( .B1(n20021), .B2(n14205), .A(n20059), .ZN(n15974) );
  INV_X1 U16708 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n13564) );
  OAI22_X1 U16709 ( .A1(n20064), .A2(n13564), .B1(n14572), .B2(n20043), .ZN(
        n13576) );
  NAND2_X1 U16710 ( .A1(n14082), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13565) );
  OAI211_X1 U16711 ( .C1(n14070), .C2(P1_EBX_REG_9__SCAN_IN), .A(n14046), .B(
        n13565), .ZN(n13566) );
  OAI21_X1 U16712 ( .B1(n14059), .B2(P1_EBX_REG_9__SCAN_IN), .A(n13566), .ZN(
        n16147) );
  MUX2_X1 U16713 ( .A(n14041), .B(n14046), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n13569) );
  NAND2_X1 U16714 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n14070), .ZN(
        n13567) );
  AND2_X1 U16715 ( .A1(n14015), .A2(n13567), .ZN(n13568) );
  NAND2_X1 U16716 ( .A1(n13569), .A2(n13568), .ZN(n13570) );
  OR2_X1 U16717 ( .A1(n16150), .A2(n13570), .ZN(n13571) );
  NAND2_X1 U16718 ( .A1(n15971), .A2(n13571), .ZN(n16141) );
  NOR3_X1 U16719 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n20021), .A3(n13572), 
        .ZN(n13573) );
  AOI211_X1 U16720 ( .C1(n20080), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n20048), .B(n13573), .ZN(n13574) );
  OAI21_X1 U16721 ( .B1(n20073), .B2(n16141), .A(n13574), .ZN(n13575) );
  AOI211_X1 U16722 ( .C1(P1_REIP_REG_10__SCAN_IN), .C2(n15974), .A(n13576), 
        .B(n13575), .ZN(n13577) );
  OAI21_X1 U16723 ( .B1(n13630), .B2(n15937), .A(n13577), .ZN(P1_U2830) );
  AOI22_X1 U16724 ( .A1(n14407), .A2(n14342), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n14405), .ZN(n13578) );
  OAI21_X1 U16725 ( .B1(n13630), .B2(n14409), .A(n13578), .ZN(P1_U2894) );
  NAND2_X1 U16726 ( .A1(n13604), .A2(n13606), .ZN(n13603) );
  AOI22_X1 U16727 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n13579), .B1(
        n19443), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13587) );
  INV_X1 U16728 ( .A(n13365), .ZN(n13581) );
  INV_X1 U16729 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13580) );
  OAI22_X1 U16730 ( .A1(n13582), .A2(n13581), .B1(n13366), .B2(n13580), .ZN(
        n13583) );
  INV_X1 U16731 ( .A(n13583), .ZN(n13586) );
  AOI22_X1 U16732 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n13356), .B1(
        n13367), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13585) );
  AOI22_X1 U16733 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n13190), .B1(
        n19624), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13584) );
  NAND4_X1 U16734 ( .A1(n13587), .A2(n13586), .A3(n13585), .A4(n13584), .ZN(
        n13597) );
  AOI22_X1 U16735 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19380), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13595) );
  AOI22_X1 U16736 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19242), .B1(
        n19662), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13594) );
  AOI22_X1 U16737 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19747), .B1(
        n19700), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13593) );
  INV_X1 U16738 ( .A(n19593), .ZN(n19596) );
  OAI22_X1 U16739 ( .A1(n13588), .A2(n13590), .B1(n19596), .B2(n13589), .ZN(
        n13591) );
  INV_X1 U16740 ( .A(n13591), .ZN(n13592) );
  NAND4_X1 U16741 ( .A1(n13595), .A2(n13594), .A3(n13593), .A4(n13592), .ZN(
        n13596) );
  INV_X1 U16742 ( .A(n13598), .ZN(n13599) );
  NAND2_X1 U16743 ( .A1(n13599), .A2(n19247), .ZN(n13600) );
  XNOR2_X2 U16744 ( .A(n13932), .B(n13933), .ZN(n13615) );
  NAND2_X1 U16745 ( .A1(n13603), .A2(n13602), .ZN(n13931) );
  INV_X1 U16746 ( .A(n13606), .ZN(n13607) );
  XNOR2_X1 U16747 ( .A(n13930), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16290) );
  NAND2_X1 U16748 ( .A1(n13611), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13612) );
  XNOR2_X1 U16749 ( .A(n13614), .B(n13613), .ZN(n19092) );
  OAI21_X2 U16750 ( .B1(n13615), .B2(n13927), .A(n19092), .ZN(n13813) );
  XNOR2_X1 U16751 ( .A(n13813), .B(n13974), .ZN(n13811) );
  XOR2_X1 U16752 ( .A(n13812), .B(n13811), .Z(n16289) );
  XNOR2_X1 U16753 ( .A(n13617), .B(n13616), .ZN(n19161) );
  NOR2_X1 U16754 ( .A1(n19161), .A2(n16313), .ZN(n13628) );
  NOR3_X1 U16755 ( .A1(n13620), .A2(n13619), .A3(n13618), .ZN(n13623) );
  NAND2_X1 U16756 ( .A1(n13621), .A2(n13623), .ZN(n13973) );
  NOR2_X1 U16757 ( .A1(n19865), .A2(n19040), .ZN(n13622) );
  AOI21_X1 U16758 ( .B1(n16304), .B2(n19100), .A(n13622), .ZN(n13626) );
  AND2_X1 U16759 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13623), .ZN(
        n13962) );
  OAI21_X1 U16760 ( .B1(n15381), .B2(n13962), .A(n13624), .ZN(n16300) );
  NAND2_X1 U16761 ( .A1(n16300), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13625) );
  OAI211_X1 U16762 ( .C1(n13973), .C2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n13626), .B(n13625), .ZN(n13627) );
  AOI211_X1 U16763 ( .C1(n16289), .C2(n16322), .A(n13628), .B(n13627), .ZN(
        n13629) );
  OAI21_X1 U16764 ( .B1(n16290), .B2(n16326), .A(n13629), .ZN(P2_U3040) );
  OAI222_X1 U16765 ( .A1(n16141), .A2(n14316), .B1(n20101), .B2(n13564), .C1(
        n14326), .C2(n13630), .ZN(P1_U2862) );
  INV_X1 U16766 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16156) );
  XNOR2_X1 U16767 ( .A(n16012), .B(n16156), .ZN(n13634) );
  XNOR2_X1 U16768 ( .A(n14411), .B(n13634), .ZN(n16153) );
  NAND2_X1 U16769 ( .A1(n16153), .A2(n20159), .ZN(n13638) );
  INV_X1 U16770 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n13635) );
  NOR2_X1 U16771 ( .A1(n20207), .A2(n13635), .ZN(n16151) );
  AND2_X1 U16772 ( .A1(n20151), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13636) );
  AOI211_X1 U16773 ( .C1(n20009), .C2(n16037), .A(n16151), .B(n13636), .ZN(
        n13637) );
  OAI211_X1 U16774 ( .C1(n15997), .C2(n20089), .A(n13638), .B(n13637), .ZN(
        P1_U2990) );
  INV_X2 U16775 ( .A(n16970), .ZN(n17213) );
  AOI22_X1 U16776 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n17194), .B1(
        P3_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n17213), .ZN(n13642) );
  AOI22_X1 U16777 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13641) );
  AOI22_X1 U16778 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n17019), .ZN(n13640) );
  NOR2_X2 U16779 ( .A1(n16944), .A2(n13644), .ZN(n15700) );
  NOR2_X2 U16780 ( .A1(n13646), .A2(n13647), .ZN(n15711) );
  AOI22_X1 U16781 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13703), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13639) );
  NAND4_X1 U16782 ( .A1(n13642), .A2(n13641), .A3(n13640), .A4(n13639), .ZN(
        n13654) );
  AOI22_X1 U16783 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17188), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13652) );
  AOI22_X1 U16784 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n16962), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n17143), .ZN(n13651) );
  AOI22_X1 U16785 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n17179), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n9817), .ZN(n13650) );
  AOI22_X1 U16786 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9820), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13649) );
  NAND4_X1 U16787 ( .A1(n13652), .A2(n13651), .A3(n13650), .A4(n13649), .ZN(
        n13653) );
  INV_X1 U16788 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n17042) );
  INV_X1 U16789 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17084) );
  AOI22_X1 U16790 ( .A1(n17208), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13658) );
  AOI22_X1 U16791 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13703), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13657) );
  AOI22_X1 U16792 ( .A1(n17197), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17019), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13656) );
  AOI22_X1 U16793 ( .A1(n9820), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17179), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13655) );
  NAND4_X1 U16794 ( .A1(n13658), .A2(n13657), .A3(n13656), .A4(n13655), .ZN(
        n13664) );
  AOI22_X1 U16795 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13661) );
  AOI22_X1 U16796 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13660) );
  AOI22_X1 U16797 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13659) );
  NAND4_X1 U16798 ( .A1(n13662), .A2(n13661), .A3(n13660), .A4(n13659), .ZN(
        n13663) );
  AOI22_X1 U16799 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13674) );
  AOI22_X1 U16800 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n16962), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13673) );
  INV_X1 U16801 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15746) );
  AOI22_X1 U16802 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9820), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13665) );
  OAI21_X1 U16803 ( .B1(n9873), .B2(n15746), .A(n13665), .ZN(n13671) );
  AOI22_X1 U16804 ( .A1(n17197), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13669) );
  INV_X2 U16805 ( .A(n17018), .ZN(n17144) );
  INV_X2 U16806 ( .A(n9883), .ZN(n17019) );
  AOI22_X1 U16807 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17019), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13668) );
  AOI22_X1 U16808 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17179), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13667) );
  AOI22_X1 U16809 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13666) );
  NAND4_X1 U16810 ( .A1(n13669), .A2(n13668), .A3(n13667), .A4(n13666), .ZN(
        n13670) );
  OAI22_X1 U16811 ( .A1(n18851), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18712), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13683) );
  AOI22_X1 U16812 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18699), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18861), .ZN(n13763) );
  NAND2_X1 U16813 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13677), .ZN(
        n13679) );
  OAI22_X1 U16814 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18716), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13677), .ZN(n13681) );
  AOI21_X1 U16815 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n13679), .A(
        n13681), .ZN(n13678) );
  NOR2_X1 U16816 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18716), .ZN(
        n13680) );
  AOI22_X1 U16817 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13681), .B1(
        n13680), .B2(n13679), .ZN(n13685) );
  NAND2_X1 U16818 ( .A1(n13684), .A2(n13683), .ZN(n13682) );
  OAI211_X1 U16819 ( .C1(n13684), .C2(n13683), .A(n13685), .B(n13682), .ZN(
        n15786) );
  AOI21_X1 U16820 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n18869), .A(
        n13764), .ZN(n15784) );
  NAND3_X1 U16821 ( .A1(n13763), .A2(n13685), .A3(n15784), .ZN(n13686) );
  NAND3_X1 U16822 ( .A1(n13765), .A2(n15786), .A3(n13686), .ZN(n16376) );
  AOI22_X1 U16823 ( .A1(n9820), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13690) );
  AOI22_X1 U16824 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13689) );
  AOI22_X1 U16825 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17019), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13688) );
  AOI22_X1 U16826 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n15691), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13687) );
  NAND4_X1 U16827 ( .A1(n13690), .A2(n13689), .A3(n13688), .A4(n13687), .ZN(
        n13696) );
  AOI22_X1 U16828 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17179), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13694) );
  AOI22_X1 U16829 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13693) );
  AOI22_X1 U16830 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n16962), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13692) );
  AOI22_X1 U16831 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13691) );
  NAND4_X1 U16832 ( .A1(n13694), .A2(n13693), .A3(n13692), .A4(n13691), .ZN(
        n13695) );
  AOI22_X1 U16833 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13702) );
  AOI22_X1 U16834 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13701) );
  AOI22_X1 U16835 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17019), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13700) );
  AOI22_X1 U16836 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13699) );
  NAND4_X1 U16837 ( .A1(n13702), .A2(n13701), .A3(n13700), .A4(n13699), .ZN(
        n13709) );
  AOI22_X1 U16838 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13707) );
  AOI22_X1 U16839 ( .A1(n17197), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n15691), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13706) );
  AOI22_X1 U16840 ( .A1(n9820), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17179), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13705) );
  AOI22_X1 U16841 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13703), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13704) );
  NAND4_X1 U16842 ( .A1(n13707), .A2(n13706), .A3(n13705), .A4(n13704), .ZN(
        n13708) );
  AOI22_X1 U16843 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13703), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13713) );
  AOI22_X1 U16844 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13712) );
  AOI22_X1 U16845 ( .A1(n17197), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n16962), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13711) );
  AOI22_X1 U16846 ( .A1(n17179), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17019), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13710) );
  NAND4_X1 U16847 ( .A1(n13713), .A2(n13712), .A3(n13711), .A4(n13710), .ZN(
        n13719) );
  BUF_X2 U16848 ( .A(n15603), .Z(n17194) );
  AOI22_X1 U16849 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13717) );
  AOI22_X1 U16850 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n15691), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13716) );
  AOI22_X1 U16851 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13715) );
  AOI22_X1 U16852 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9820), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13714) );
  NAND4_X1 U16853 ( .A1(n13717), .A2(n13716), .A3(n13715), .A4(n13714), .ZN(
        n13718) );
  AOI22_X1 U16854 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13723) );
  AOI22_X1 U16855 ( .A1(n9820), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13722) );
  AOI22_X1 U16856 ( .A1(n17197), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13721) );
  AOI22_X1 U16857 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17019), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13720) );
  NAND4_X1 U16858 ( .A1(n13723), .A2(n13722), .A3(n13721), .A4(n13720), .ZN(
        n13729) );
  AOI22_X1 U16859 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13727) );
  AOI22_X1 U16860 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17179), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13726) );
  AOI22_X1 U16861 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13725) );
  INV_X2 U16862 ( .A(n9873), .ZN(n15691) );
  AOI22_X1 U16863 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n15691), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13724) );
  NAND4_X1 U16864 ( .A1(n13727), .A2(n13726), .A3(n13725), .A4(n13724), .ZN(
        n13728) );
  BUF_X2 U16865 ( .A(n15713), .Z(n15699) );
  AOI22_X1 U16866 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15699), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13733) );
  AOI22_X1 U16867 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17019), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13732) );
  AOI22_X1 U16868 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13731) );
  AOI22_X1 U16869 ( .A1(n17208), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13730) );
  NAND4_X1 U16870 ( .A1(n13733), .A2(n13732), .A3(n13731), .A4(n13730), .ZN(
        n13740) );
  AOI22_X1 U16871 ( .A1(n9820), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17197), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13738) );
  AOI22_X1 U16872 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13737) );
  AOI22_X1 U16873 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n15691), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13736) );
  AOI22_X1 U16874 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13735) );
  NAND4_X1 U16875 ( .A1(n13738), .A2(n13737), .A3(n13736), .A4(n13735), .ZN(
        n13739) );
  NAND2_X1 U16876 ( .A1(n18244), .A2(n17271), .ZN(n15794) );
  NAND2_X1 U16877 ( .A1(n13757), .A2(n15794), .ZN(n13754) );
  NAND2_X1 U16878 ( .A1(n15802), .A2(n13754), .ZN(n13768) );
  INV_X1 U16879 ( .A(n18253), .ZN(n13771) );
  NAND2_X1 U16880 ( .A1(n18263), .A2(n13771), .ZN(n18688) );
  NAND2_X1 U16881 ( .A1(n18248), .A2(n18244), .ZN(n18687) );
  NOR3_X1 U16882 ( .A1(n18263), .A2(n17271), .A3(n18687), .ZN(n13755) );
  NOR2_X1 U16883 ( .A1(n17351), .A2(n13771), .ZN(n13741) );
  AOI22_X1 U16884 ( .A1(n18678), .A2(n15801), .B1(n13755), .B2(n13741), .ZN(
        n15912) );
  NOR4_X2 U16885 ( .A1(n18889), .A2(n18237), .A3(n15912), .A4(n18732), .ZN(
        n17257) );
  INV_X1 U16886 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17250) );
  NAND2_X1 U16887 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17251) );
  NOR2_X1 U16888 ( .A1(n17250), .A2(n17251), .ZN(n17240) );
  NAND3_X1 U16889 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n17240), .ZN(n15648) );
  NAND4_X1 U16890 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .A3(P3_EBX_REG_6__SCAN_IN), .A4(P3_EBX_REG_5__SCAN_IN), .ZN(n15649) );
  INV_X1 U16891 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16794) );
  NAND4_X1 U16892 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(P3_EBX_REG_11__SCAN_IN), 
        .A3(P3_EBX_REG_10__SCAN_IN), .A4(P3_EBX_REG_9__SCAN_IN), .ZN(n13742)
         );
  NOR2_X1 U16893 ( .A1(n16794), .A2(n13742), .ZN(n15650) );
  NAND4_X1 U16894 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_15__SCAN_IN), 
        .A3(P3_EBX_REG_14__SCAN_IN), .A4(n15650), .ZN(n13743) );
  NOR3_X1 U16895 ( .A1(n15648), .A2(n15649), .A3(n13743), .ZN(n17097) );
  NAND3_X1 U16896 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17257), .A3(n17097), 
        .ZN(n17073) );
  NOR2_X1 U16897 ( .A1(n17084), .A2(n17073), .ZN(n17071) );
  NAND2_X1 U16898 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17071), .ZN(n17070) );
  INV_X1 U16899 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16653) );
  INV_X1 U16900 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16679) );
  NOR2_X1 U16901 ( .A1(n16653), .A2(n16679), .ZN(n13744) );
  NAND4_X1 U16902 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(P3_EBX_REG_21__SCAN_IN), .A4(n13744), .ZN(n15560) );
  NAND4_X1 U16903 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_28__SCAN_IN), 
        .A3(P3_EBX_REG_27__SCAN_IN), .A4(P3_EBX_REG_26__SCAN_IN), .ZN(n13745)
         );
  NOR4_X1 U16904 ( .A1(n17042), .A2(n17070), .A3(n15560), .A4(n13745), .ZN(
        n16981) );
  NAND2_X1 U16905 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16981), .ZN(n13746) );
  NOR2_X1 U16906 ( .A1(n17351), .A2(n13746), .ZN(n13748) );
  NAND2_X1 U16907 ( .A1(n17246), .A2(n13746), .ZN(n16982) );
  INV_X1 U16908 ( .A(n16982), .ZN(n13747) );
  MUX2_X1 U16909 ( .A(n13748), .B(n13747), .S(P3_EBX_REG_31__SCAN_IN), .Z(
        P3_U2672) );
  NAND2_X1 U16910 ( .A1(n18847), .A2(n18863), .ZN(n18900) );
  NAND4_X1 U16911 ( .A1(n18248), .A2(n18253), .A3(n13756), .A4(n13750), .ZN(
        n13759) );
  NAND2_X1 U16912 ( .A1(n17271), .A2(n18263), .ZN(n15916) );
  INV_X1 U16913 ( .A(n15916), .ZN(n18695) );
  OAI211_X1 U16914 ( .C1(n18268), .C2(n18695), .A(n18889), .B(n17415), .ZN(
        n13772) );
  NAND2_X1 U16915 ( .A1(n18244), .A2(n13750), .ZN(n15787) );
  NAND2_X1 U16916 ( .A1(n13757), .A2(n15787), .ZN(n13753) );
  INV_X1 U16917 ( .A(n18248), .ZN(n13749) );
  OAI22_X1 U16918 ( .A1(n13756), .A2(n13749), .B1(n13771), .B2(n15916), .ZN(
        n13752) );
  NOR2_X1 U16919 ( .A1(n18268), .A2(n13750), .ZN(n13751) );
  INV_X1 U16920 ( .A(n18244), .ZN(n15791) );
  OAI211_X1 U16921 ( .C1(n18248), .C2(n13754), .A(n13772), .B(n13773), .ZN(
        n15804) );
  NAND3_X1 U16922 ( .A1(n13756), .A2(n13755), .A3(n18889), .ZN(n13761) );
  NOR2_X2 U16923 ( .A1(n17471), .A2(n13774), .ZN(n16557) );
  NOR2_X2 U16924 ( .A1(n16557), .A2(n13760), .ZN(n15803) );
  NOR2_X2 U16925 ( .A1(n17471), .A2(n15803), .ZN(n18671) );
  NOR2_X1 U16926 ( .A1(n18851), .A2(n18861), .ZN(n18690) );
  AOI21_X1 U16927 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18690), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13779) );
  OR2_X1 U16928 ( .A1(n18670), .A2(n13779), .ZN(n18681) );
  NOR2_X1 U16929 ( .A1(n18900), .A2(n18681), .ZN(n13778) );
  XNOR2_X1 U16930 ( .A(n13764), .B(n13763), .ZN(n13766) );
  INV_X1 U16931 ( .A(n18673), .ZN(n15795) );
  NAND2_X1 U16932 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n18890) );
  NAND2_X1 U16933 ( .A1(n15795), .A2(n18890), .ZN(n13776) );
  NAND2_X1 U16934 ( .A1(n18889), .A2(n17471), .ZN(n18725) );
  INV_X1 U16935 ( .A(n18725), .ZN(n17472) );
  NAND2_X1 U16936 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18758), .ZN(n18898) );
  INV_X1 U16937 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18761) );
  NOR2_X1 U16938 ( .A1(n18898), .A2(n18761), .ZN(n18760) );
  NOR2_X1 U16939 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18745) );
  NOR3_X1 U16940 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18760), .A3(n18745), 
        .ZN(n18751) );
  OAI21_X1 U16941 ( .B1(n15803), .B2(n17472), .A(n18751), .ZN(n17413) );
  INV_X1 U16942 ( .A(n17471), .ZN(n13767) );
  INV_X1 U16943 ( .A(n18263), .ZN(n13770) );
  AOI211_X1 U16944 ( .C1(n13771), .C2(n13770), .A(n13769), .B(n13768), .ZN(
        n15798) );
  OAI211_X1 U16945 ( .C1(n13774), .C2(n15798), .A(n13773), .B(n13772), .ZN(
        n15788) );
  AOI211_X1 U16946 ( .C1(n15801), .C2(n18678), .A(n15914), .B(n15788), .ZN(
        n13775) );
  OAI21_X1 U16947 ( .B1(n13776), .B2(n17413), .A(n13775), .ZN(n18710) );
  NOR2_X1 U16948 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18863), .ZN(n18236) );
  INV_X1 U16949 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18224) );
  INV_X1 U16950 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18726) );
  NOR3_X1 U16951 ( .A1(n18847), .A2(n18735), .A3(n18726), .ZN(n18742) );
  INV_X1 U16952 ( .A(n18742), .ZN(n18834) );
  NOR2_X1 U16953 ( .A1(n18224), .A2(n18834), .ZN(n13777) );
  AOI211_X2 U16954 ( .C1(n18882), .C2(n18710), .A(n18236), .B(n13777), .ZN(
        n18868) );
  MUX2_X1 U16955 ( .A(n13778), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n18868), .Z(P3_U3284) );
  NAND2_X1 U16956 ( .A1(n13779), .A2(n17018), .ZN(n18223) );
  NOR2_X1 U16957 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18223), .ZN(n13780) );
  INV_X1 U16958 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18682) );
  NAND2_X1 U16959 ( .A1(n18682), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18854) );
  OAI221_X1 U16960 ( .B1(n18726), .B2(P3_STATE2_REG_1__SCAN_IN), .C1(
        P3_STATE2_REG_2__SCAN_IN), .C2(n18847), .A(n18854), .ZN(n18235) );
  NAND2_X1 U16961 ( .A1(n18735), .A2(n18235), .ZN(n18426) );
  OAI21_X1 U16962 ( .B1(n13780), .B2(n18834), .A(n18426), .ZN(n18229) );
  INV_X1 U16963 ( .A(n18229), .ZN(n13781) );
  NAND2_X1 U16964 ( .A1(n18726), .A2(n18863), .ZN(n16554) );
  AND2_X1 U16965 ( .A1(n18900), .A2(n16554), .ZN(n18881) );
  INV_X1 U16966 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18888) );
  NOR2_X1 U16967 ( .A1(n18847), .A2(n18888), .ZN(n17846) );
  NOR2_X1 U16968 ( .A1(n18881), .A2(n17846), .ZN(n15654) );
  AOI21_X1 U16969 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n15654), .ZN(n15655) );
  NOR2_X1 U16970 ( .A1(n13781), .A2(n15655), .ZN(n13783) );
  NAND3_X1 U16971 ( .A1(n18726), .A2(n18863), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18473) );
  INV_X1 U16972 ( .A(n18473), .ZN(n18520) );
  NOR2_X1 U16973 ( .A1(n18863), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18273) );
  OR2_X1 U16974 ( .A1(n18273), .A2(n13781), .ZN(n15653) );
  OR2_X1 U16975 ( .A1(n18520), .A2(n15653), .ZN(n13782) );
  MUX2_X1 U16976 ( .A(n13783), .B(n13782), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  OAI22_X1 U16977 ( .A1(n13785), .A2(n15374), .B1(n16316), .B2(n13784), .ZN(
        n13797) );
  INV_X1 U16978 ( .A(n13961), .ZN(n13795) );
  AOI21_X1 U16979 ( .B1(n13788), .B2(n13787), .A(n13786), .ZN(n13802) );
  NOR2_X1 U16980 ( .A1(n19860), .A2(n19040), .ZN(n13792) );
  NAND2_X1 U16981 ( .A1(n13790), .A2(n13789), .ZN(n13807) );
  AND3_X1 U16982 ( .A1(n16322), .A2(n13808), .A3(n13807), .ZN(n13791) );
  AOI211_X1 U16983 ( .C1(n13802), .C2(n16301), .A(n13792), .B(n13791), .ZN(
        n13793) );
  OAI21_X1 U16984 ( .B1(n13795), .B2(n13794), .A(n13793), .ZN(n13796) );
  AOI211_X1 U16985 ( .C1(n16299), .C2(n13798), .A(n13797), .B(n13796), .ZN(
        n13801) );
  INV_X1 U16986 ( .A(n13799), .ZN(n13800) );
  OAI211_X1 U16987 ( .C1(n9829), .C2(n16314), .A(n13801), .B(n13800), .ZN(
        P2_U3044) );
  INV_X1 U16988 ( .A(n13802), .ZN(n13804) );
  AOI22_X1 U16989 ( .A1(n15162), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        P2_REIP_REG_2__SCAN_IN), .B2(n19223), .ZN(n13803) );
  OAI21_X1 U16990 ( .B1(n13804), .B2(n19225), .A(n13803), .ZN(n13805) );
  AOI21_X1 U16991 ( .B1(n19222), .B2(n13806), .A(n13805), .ZN(n13810) );
  NAND3_X1 U16992 ( .A1(n13808), .A2(n16282), .A3(n13807), .ZN(n13809) );
  OAI211_X1 U16993 ( .C1(n9829), .C2(n13154), .A(n13810), .B(n13809), .ZN(
        P2_U3012) );
  NAND2_X1 U16994 ( .A1(n13813), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13814) );
  OAI21_X1 U16995 ( .B1(n13816), .B2(n13815), .A(n13823), .ZN(n19069) );
  OR2_X1 U16996 ( .A1(n19069), .A2(n13941), .ZN(n13820) );
  NOR2_X1 U16997 ( .A1(n13820), .A2(n11001), .ZN(n16279) );
  INV_X1 U16998 ( .A(n13817), .ZN(n13818) );
  XNOR2_X1 U16999 ( .A(n13819), .B(n13818), .ZN(n19082) );
  NAND2_X1 U17000 ( .A1(n13820), .A2(n11001), .ZN(n16277) );
  INV_X1 U17001 ( .A(n19082), .ZN(n13821) );
  NAND2_X1 U17002 ( .A1(n13821), .A2(n15511), .ZN(n16276) );
  AND2_X1 U17003 ( .A1(n16277), .A2(n16276), .ZN(n13822) );
  NAND2_X1 U17004 ( .A1(n19267), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n13824) );
  MUX2_X1 U17005 ( .A(n19267), .B(n13824), .S(n13823), .Z(n13825) );
  NAND2_X1 U17006 ( .A1(n10091), .A2(n13825), .ZN(n14803) );
  OAI21_X1 U17007 ( .B1(n14803), .B2(n13941), .A(n13826), .ZN(n15506) );
  NAND2_X1 U17008 ( .A1(n19267), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n13828) );
  MUX2_X1 U17009 ( .A(n13828), .B(P2_EBX_REG_10__SCAN_IN), .S(n13827), .Z(
        n13829) );
  AND2_X1 U17010 ( .A1(n13829), .A2(n13906), .ZN(n19054) );
  AOI21_X1 U17011 ( .B1(n19054), .B2(n13927), .A(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15195) );
  INV_X1 U17012 ( .A(n19054), .ZN(n13831) );
  NAND2_X1 U17013 ( .A1(n13927), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13830) );
  INV_X1 U17014 ( .A(n14803), .ZN(n13833) );
  AND2_X1 U17015 ( .A1(n13927), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13832) );
  NAND2_X1 U17016 ( .A1(n13833), .A2(n13832), .ZN(n15505) );
  INV_X1 U17017 ( .A(n13835), .ZN(n13836) );
  AND3_X1 U17018 ( .A1(n19267), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n13836), .ZN(
        n13837) );
  OR2_X1 U17019 ( .A1(n13838), .A2(n13837), .ZN(n19043) );
  NOR2_X1 U17020 ( .A1(n19043), .A2(n13941), .ZN(n13839) );
  AND2_X1 U17021 ( .A1(n13839), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15466) );
  INV_X1 U17022 ( .A(n13839), .ZN(n13840) );
  INV_X1 U17023 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15471) );
  NAND2_X1 U17024 ( .A1(n13840), .A2(n15471), .ZN(n15465) );
  INV_X1 U17025 ( .A(n13841), .ZN(n13842) );
  NOR2_X1 U17026 ( .A1(n13842), .A2(n11019), .ZN(n13843) );
  AND2_X1 U17027 ( .A1(n19267), .A2(n13843), .ZN(n13844) );
  NOR2_X1 U17028 ( .A1(n13876), .A2(n13844), .ZN(n19032) );
  AND2_X1 U17029 ( .A1(n13927), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13845) );
  NAND2_X1 U17030 ( .A1(n19032), .A2(n13845), .ZN(n15182) );
  INV_X1 U17031 ( .A(n19032), .ZN(n13846) );
  INV_X1 U17032 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15441) );
  OAI21_X1 U17033 ( .B1(n13846), .B2(n13941), .A(n15441), .ZN(n15183) );
  INV_X1 U17034 ( .A(n13847), .ZN(n13848) );
  NAND3_X1 U17035 ( .A1(n13848), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n19267), 
        .ZN(n13849) );
  AND2_X1 U17036 ( .A1(n13850), .A2(n13849), .ZN(n13884) );
  INV_X1 U17037 ( .A(n13884), .ZN(n14792) );
  OAI21_X1 U17038 ( .B1(n14792), .B2(n13941), .A(n15109), .ZN(n15105) );
  INV_X1 U17039 ( .A(n13851), .ZN(n13852) );
  NAND2_X1 U17040 ( .A1(n9880), .A2(n13852), .ZN(n13853) );
  NAND2_X1 U17041 ( .A1(n9876), .A2(n13853), .ZN(n18948) );
  OR2_X1 U17042 ( .A1(n18948), .A2(n13941), .ZN(n13854) );
  NAND2_X1 U17043 ( .A1(n13854), .A2(n15337), .ZN(n15129) );
  NAND2_X1 U17044 ( .A1(n13863), .A2(n13855), .ZN(n13856) );
  NAND2_X1 U17045 ( .A1(n9880), .A2(n13856), .ZN(n18963) );
  OR2_X1 U17046 ( .A1(n18963), .A2(n13941), .ZN(n13857) );
  NAND2_X1 U17047 ( .A1(n13857), .A2(n15366), .ZN(n15137) );
  NAND2_X1 U17048 ( .A1(n15129), .A2(n15137), .ZN(n15100) );
  AND2_X1 U17049 ( .A1(n19267), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n13859) );
  INV_X1 U17050 ( .A(n13906), .ZN(n13858) );
  AOI21_X1 U17051 ( .B1(n13872), .B2(n13859), .A(n13858), .ZN(n13860) );
  OR2_X1 U17052 ( .A1(n13872), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n13862) );
  NAND2_X1 U17053 ( .A1(n18986), .A2(n13927), .ZN(n13861) );
  XNOR2_X1 U17054 ( .A(n13861), .B(n15403), .ZN(n15098) );
  NAND3_X1 U17055 ( .A1(n13862), .A2(P2_EBX_REG_17__SCAN_IN), .A3(n19267), 
        .ZN(n13864) );
  AND2_X1 U17056 ( .A1(n13864), .A2(n13863), .ZN(n13888) );
  INV_X1 U17057 ( .A(n13888), .ZN(n18971) );
  NAND2_X1 U17058 ( .A1(n19267), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n13865) );
  MUX2_X1 U17059 ( .A(n13865), .B(n19267), .S(n13878), .Z(n13867) );
  NAND2_X1 U17060 ( .A1(n13878), .A2(n13866), .ZN(n13871) );
  NAND2_X1 U17061 ( .A1(n13867), .A2(n13871), .ZN(n19010) );
  NOR2_X1 U17062 ( .A1(n19010), .A2(n13941), .ZN(n13886) );
  INV_X1 U17063 ( .A(n13886), .ZN(n13869) );
  INV_X1 U17064 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n13868) );
  NAND2_X1 U17065 ( .A1(n13869), .A2(n13868), .ZN(n15170) );
  AND2_X1 U17066 ( .A1(n19267), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n13870) );
  NAND2_X1 U17067 ( .A1(n13871), .A2(n13870), .ZN(n13873) );
  NAND2_X1 U17068 ( .A1(n13873), .A2(n13872), .ZN(n18996) );
  OR2_X1 U17069 ( .A1(n18996), .A2(n13941), .ZN(n13874) );
  INV_X1 U17070 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15415) );
  NAND2_X1 U17071 ( .A1(n13874), .A2(n15415), .ZN(n15406) );
  NOR2_X1 U17072 ( .A1(n13876), .A2(n13875), .ZN(n13877) );
  OR2_X1 U17073 ( .A1(n13878), .A2(n13877), .ZN(n19018) );
  OAI21_X1 U17074 ( .B1(n19018), .B2(n13941), .A(n15437), .ZN(n15434) );
  NAND4_X1 U17075 ( .A1(n15149), .A2(n15170), .A3(n15406), .A4(n15434), .ZN(
        n13879) );
  NOR3_X1 U17076 ( .A1(n15100), .A2(n15098), .A3(n13879), .ZN(n13882) );
  AND2_X1 U17077 ( .A1(n19267), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n13880) );
  XNOR2_X1 U17078 ( .A(n9876), .B(n13880), .ZN(n13894) );
  INV_X1 U17079 ( .A(n13894), .ZN(n18935) );
  NAND2_X1 U17080 ( .A1(n18935), .A2(n13927), .ZN(n13881) );
  NAND2_X1 U17081 ( .A1(n13881), .A2(n15338), .ZN(n15103) );
  NAND3_X1 U17082 ( .A1(n15105), .A2(n13882), .A3(n15103), .ZN(n13897) );
  AND2_X1 U17083 ( .A1(n13927), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13883) );
  NAND2_X1 U17084 ( .A1(n13884), .A2(n13883), .ZN(n15104) );
  OR3_X1 U17085 ( .A1(n18948), .A2(n13941), .A3(n15337), .ZN(n15128) );
  NAND2_X1 U17086 ( .A1(n13927), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13885) );
  OR2_X1 U17087 ( .A1(n18963), .A2(n13885), .ZN(n15136) );
  AND2_X1 U17088 ( .A1(n15128), .A2(n15136), .ZN(n15101) );
  AND2_X1 U17089 ( .A1(n13927), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13887) );
  NAND2_X1 U17090 ( .A1(n13888), .A2(n13887), .ZN(n15148) );
  AND2_X1 U17091 ( .A1(n13927), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13889) );
  NAND2_X1 U17092 ( .A1(n18986), .A2(n13889), .ZN(n15099) );
  NAND2_X1 U17093 ( .A1(n13927), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13890) );
  OR2_X1 U17094 ( .A1(n18996), .A2(n13890), .ZN(n15405) );
  INV_X1 U17095 ( .A(n19018), .ZN(n13892) );
  AND2_X1 U17096 ( .A1(n13927), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13891) );
  NAND2_X1 U17097 ( .A1(n13892), .A2(n13891), .ZN(n15433) );
  NAND4_X1 U17098 ( .A1(n15148), .A2(n15099), .A3(n15405), .A4(n15433), .ZN(
        n13893) );
  NOR2_X1 U17099 ( .A1(n15174), .A2(n13893), .ZN(n13895) );
  OR3_X1 U17100 ( .A1(n13894), .A2(n13941), .A3(n15338), .ZN(n15102) );
  AND4_X1 U17101 ( .A1(n15104), .A2(n15101), .A3(n13895), .A4(n15102), .ZN(
        n13896) );
  OR2_X1 U17102 ( .A1(n13900), .A2(n13941), .ZN(n13898) );
  NAND2_X1 U17103 ( .A1(n13898), .A2(n13899), .ZN(n15089) );
  OR2_X1 U17104 ( .A1(n13903), .A2(n13941), .ZN(n13901) );
  XNOR2_X1 U17105 ( .A(n13901), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15082) );
  NAND2_X1 U17106 ( .A1(n15083), .A2(n15082), .ZN(n13905) );
  NAND2_X1 U17107 ( .A1(n13927), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13902) );
  NAND2_X1 U17108 ( .A1(n13905), .A2(n13904), .ZN(n15067) );
  NAND2_X1 U17109 ( .A1(n13906), .A2(n13927), .ZN(n15068) );
  NOR2_X1 U17110 ( .A1(n15068), .A2(n15289), .ZN(n13908) );
  NAND2_X1 U17111 ( .A1(n15068), .A2(n15289), .ZN(n13907) );
  INV_X1 U17112 ( .A(n13909), .ZN(n13911) );
  NAND3_X1 U17113 ( .A1(n19267), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n16221), 
        .ZN(n13910) );
  OAI21_X1 U17114 ( .B1(n16207), .B2(n13941), .A(n15272), .ZN(n13912) );
  INV_X1 U17115 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15060) );
  AND2_X1 U17116 ( .A1(n15068), .A2(n15060), .ZN(n15055) );
  INV_X1 U17117 ( .A(n15068), .ZN(n13916) );
  NAND2_X1 U17118 ( .A1(n13916), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15056) );
  INV_X1 U17119 ( .A(n13918), .ZN(n13919) );
  XNOR2_X1 U17120 ( .A(n13920), .B(n13919), .ZN(n16199) );
  NAND2_X1 U17121 ( .A1(n16199), .A2(n13927), .ZN(n15026) );
  INV_X1 U17122 ( .A(n15026), .ZN(n13921) );
  XNOR2_X1 U17123 ( .A(n13923), .B(n13922), .ZN(n13926) );
  OAI21_X1 U17124 ( .B1(n13926), .B2(n13941), .A(n15234), .ZN(n15010) );
  INV_X1 U17125 ( .A(n13925), .ZN(n13924) );
  AOI21_X1 U17126 ( .B1(n13924), .B2(n13927), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15000) );
  INV_X1 U17127 ( .A(n13926), .ZN(n14772) );
  NAND3_X1 U17128 ( .A1(n14772), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n13927), .ZN(n15011) );
  XOR2_X1 U17129 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n13916), .Z(
        n13928) );
  XNOR2_X1 U17130 ( .A(n13929), .B(n13928), .ZN(n13998) );
  INV_X1 U17131 ( .A(n13933), .ZN(n13934) );
  NAND2_X1 U17132 ( .A1(n15206), .A2(n15511), .ZN(n13936) );
  NAND2_X1 U17133 ( .A1(n15205), .A2(n13936), .ZN(n13939) );
  INV_X1 U17134 ( .A(n15206), .ZN(n13937) );
  NAND2_X1 U17135 ( .A1(n13937), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13938) );
  NAND2_X1 U17136 ( .A1(n16273), .A2(n16274), .ZN(n13944) );
  AND2_X1 U17137 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15440) );
  NAND2_X1 U17138 ( .A1(n15440), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15425) );
  NOR2_X2 U17139 ( .A1(n15108), .A2(n15109), .ZN(n15086) );
  AND2_X1 U17140 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15268) );
  NAND2_X1 U17141 ( .A1(n15268), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15228) );
  NOR2_X1 U17142 ( .A1(n15228), .A2(n15255), .ZN(n13981) );
  INV_X1 U17143 ( .A(n13945), .ZN(n13946) );
  NAND2_X1 U17144 ( .A1(n12661), .A2(n13946), .ZN(n13949) );
  AOI22_X1 U17145 ( .A1(n13947), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n13948) );
  OAI211_X1 U17146 ( .C1(n13950), .C2(n14827), .A(n13949), .B(n13948), .ZN(
        n13953) );
  INV_X1 U17147 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n14759) );
  NAND2_X1 U17148 ( .A1(n13954), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13957) );
  NAND2_X1 U17149 ( .A1(n13955), .A2(P2_EAX_REG_31__SCAN_IN), .ZN(n13956) );
  OAI211_X1 U17150 ( .C1(n13958), .C2(n14759), .A(n13957), .B(n13956), .ZN(
        n13959) );
  XNOR2_X1 U17151 ( .A(n13960), .B(n13959), .ZN(n14757) );
  NAND2_X1 U17152 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16306) );
  INV_X1 U17153 ( .A(n16306), .ZN(n13975) );
  AND3_X1 U17154 ( .A1(n13975), .A2(n13962), .A3(n13961), .ZN(n13963) );
  OR2_X1 U17155 ( .A1(n15381), .A2(n13963), .ZN(n13966) );
  NOR2_X1 U17156 ( .A1(n13964), .A2(n13826), .ZN(n13965) );
  AND2_X1 U17157 ( .A1(n13966), .A2(n13965), .ZN(n15500) );
  AND2_X1 U17158 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n13976) );
  NAND2_X1 U17159 ( .A1(n15500), .A2(n13976), .ZN(n13967) );
  NAND2_X1 U17160 ( .A1(n13967), .A2(n15316), .ZN(n15445) );
  NAND3_X1 U17161 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n13968) );
  NOR2_X1 U17162 ( .A1(n15425), .A2(n13968), .ZN(n15363) );
  AND2_X1 U17163 ( .A1(n15363), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13977) );
  OR2_X1 U17164 ( .A1(n15381), .A2(n13977), .ZN(n13969) );
  NAND2_X1 U17165 ( .A1(n15445), .A2(n13969), .ZN(n15362) );
  NAND2_X1 U17166 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n13979) );
  INV_X1 U17167 ( .A(n13979), .ZN(n15336) );
  OAI21_X1 U17168 ( .B1(n15381), .B2(n15336), .A(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n13970) );
  NAND2_X1 U17169 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n13980) );
  NOR2_X1 U17170 ( .A1(n15325), .A2(n13980), .ZN(n15290) );
  NAND4_X1 U17171 ( .A1(n15290), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A4(n13981), .ZN(n13971) );
  NAND2_X1 U17172 ( .A1(n13971), .A2(n15316), .ZN(n15218) );
  OAI21_X1 U17173 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15381), .A(
        n15218), .ZN(n13972) );
  NAND2_X1 U17174 ( .A1(n13972), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13985) );
  NAND2_X1 U17175 ( .A1(n16307), .A2(n13975), .ZN(n15501) );
  NAND2_X1 U17176 ( .A1(n15485), .A2(n13976), .ZN(n15458) );
  INV_X1 U17177 ( .A(n13977), .ZN(n13978) );
  NOR2_X1 U17178 ( .A1(n15354), .A2(n13979), .ZN(n15326) );
  NAND2_X1 U17179 ( .A1(n15326), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15313) );
  INV_X1 U17180 ( .A(n13981), .ZN(n13982) );
  NOR2_X1 U17181 ( .A1(n15297), .A2(n13982), .ZN(n15233) );
  NAND2_X1 U17182 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n15233), .ZN(
        n15235) );
  NOR2_X1 U17183 ( .A1(n15234), .A2(n15235), .ZN(n15215) );
  NOR2_X1 U17184 ( .A1(n9832), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13983) );
  NOR2_X1 U17185 ( .A1(n19083), .A2(n14759), .ZN(n13990) );
  AOI21_X1 U17186 ( .B1(n15215), .B2(n13983), .A(n13990), .ZN(n13984) );
  OAI211_X1 U17187 ( .C1(n14757), .C2(n16313), .A(n13985), .B(n13984), .ZN(
        n13986) );
  AOI21_X1 U17188 ( .B1(n14825), .B2(n16304), .A(n13986), .ZN(n13987) );
  OAI21_X1 U17189 ( .B1(n13995), .B2(n16326), .A(n13987), .ZN(n13988) );
  INV_X1 U17190 ( .A(n13988), .ZN(n13989) );
  OAI21_X1 U17191 ( .B1(n13998), .B2(n15495), .A(n13989), .ZN(P2_U3015) );
  AOI21_X1 U17192 ( .B1(n15162), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n13990), .ZN(n13991) );
  OAI21_X1 U17193 ( .B1(n15211), .B2(n13992), .A(n13991), .ZN(n13993) );
  AOI21_X1 U17194 ( .B1(n14825), .B2(n19231), .A(n13993), .ZN(n13994) );
  OAI21_X1 U17195 ( .B1(n13995), .B2(n19225), .A(n13994), .ZN(n13996) );
  INV_X1 U17196 ( .A(n13996), .ZN(n13997) );
  OAI21_X1 U17197 ( .B1(n13998), .B2(n19227), .A(n13997), .ZN(P2_U2983) );
  AOI22_X1 U17198 ( .A1(n12579), .A2(n13999), .B1(n14005), .B2(n14007), .ZN(
        n14002) );
  NAND2_X1 U17199 ( .A1(n14000), .A2(n14003), .ZN(n14001) );
  OAI211_X1 U17200 ( .C1(n14004), .C2(n14003), .A(n14002), .B(n14001), .ZN(
        n15865) );
  OR2_X1 U17201 ( .A1(n14006), .A2(n14005), .ZN(n14009) );
  NAND2_X1 U17202 ( .A1(n14007), .A2(n14010), .ZN(n14008) );
  AND2_X1 U17203 ( .A1(n14009), .A2(n14008), .ZN(n19981) );
  NAND3_X1 U17204 ( .A1(n14070), .A2(n14010), .A3(n15906), .ZN(n14011) );
  NAND2_X1 U17205 ( .A1(n14011), .A2(n20906), .ZN(n20900) );
  NAND2_X1 U17206 ( .A1(n19981), .A2(n20900), .ZN(n15864) );
  AND2_X1 U17207 ( .A1(n15864), .A2(n14012), .ZN(n19989) );
  MUX2_X1 U17208 ( .A(P1_MORE_REG_SCAN_IN), .B(n15865), .S(n19989), .Z(
        P1_U3484) );
  AOI22_X1 U17209 ( .A1(n14071), .A2(P1_EBX_REG_30__SCAN_IN), .B1(n14070), 
        .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14084) );
  MUX2_X1 U17210 ( .A(n14059), .B(n14082), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n14013) );
  OAI21_X1 U17211 ( .B1(n14071), .B2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n14013), .ZN(n15970) );
  MUX2_X1 U17212 ( .A(n14041), .B(n14046), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n14017) );
  NAND2_X1 U17213 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14070), .ZN(
        n14014) );
  AND2_X1 U17214 ( .A1(n14015), .A2(n14014), .ZN(n14016) );
  MUX2_X1 U17215 ( .A(n14059), .B(n14082), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n14018) );
  OAI21_X1 U17216 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n14071), .A(
        n14018), .ZN(n14245) );
  INV_X1 U17217 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16110) );
  NAND2_X1 U17218 ( .A1(n14046), .A2(n16110), .ZN(n14020) );
  INV_X1 U17219 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n21236) );
  NAND2_X1 U17220 ( .A1(n14067), .A2(n21236), .ZN(n14019) );
  NAND3_X1 U17221 ( .A1(n14020), .A2(n14082), .A3(n14019), .ZN(n14021) );
  OAI21_X1 U17222 ( .B1(n14041), .B2(P1_EBX_REG_14__SCAN_IN), .A(n14021), .ZN(
        n14228) );
  MUX2_X1 U17223 ( .A(n14059), .B(n14082), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n14023) );
  OR2_X1 U17224 ( .A1(n14071), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14022) );
  NAND2_X1 U17225 ( .A1(n14023), .A2(n14022), .ZN(n14220) );
  INV_X1 U17226 ( .A(n14220), .ZN(n14024) );
  INV_X1 U17227 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n15953) );
  NAND2_X1 U17228 ( .A1(n14062), .A2(n15953), .ZN(n14028) );
  INV_X1 U17229 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16090) );
  NAND2_X1 U17230 ( .A1(n14046), .A2(n16090), .ZN(n14026) );
  NAND2_X1 U17231 ( .A1(n14067), .A2(n15953), .ZN(n14025) );
  NAND3_X1 U17232 ( .A1(n14026), .A2(n14082), .A3(n14025), .ZN(n14027) );
  MUX2_X1 U17233 ( .A(n14059), .B(n14082), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n14029) );
  OAI21_X1 U17234 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n14071), .A(
        n14029), .ZN(n14201) );
  INV_X1 U17235 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16089) );
  NAND2_X1 U17236 ( .A1(n14046), .A2(n16089), .ZN(n14031) );
  INV_X1 U17237 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n20959) );
  NAND2_X1 U17238 ( .A1(n14067), .A2(n20959), .ZN(n14030) );
  NAND3_X1 U17239 ( .A1(n14031), .A2(n14082), .A3(n14030), .ZN(n14032) );
  OAI21_X1 U17240 ( .B1(n14041), .B2(P1_EBX_REG_18__SCAN_IN), .A(n14032), .ZN(
        n14298) );
  INV_X1 U17241 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n21034) );
  NAND2_X1 U17242 ( .A1(n14044), .A2(n21034), .ZN(n14035) );
  NAND2_X1 U17243 ( .A1(n14082), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14033) );
  OAI211_X1 U17244 ( .C1(n14070), .C2(P1_EBX_REG_19__SCAN_IN), .A(n14046), .B(
        n14033), .ZN(n14034) );
  AND2_X1 U17245 ( .A1(n14035), .A2(n14034), .ZN(n14189) );
  MUX2_X1 U17246 ( .A(n14041), .B(n14046), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n14037) );
  NAND2_X1 U17247 ( .A1(n14070), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14036) );
  NAND2_X1 U17248 ( .A1(n14037), .A2(n14036), .ZN(n14292) );
  INV_X1 U17249 ( .A(n14292), .ZN(n14038) );
  INV_X1 U17250 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14039) );
  MUX2_X1 U17251 ( .A(n14082), .B(n14059), .S(n14039), .Z(n14040) );
  OAI21_X1 U17252 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n14071), .A(
        n14040), .ZN(n15889) );
  MUX2_X1 U17253 ( .A(n14041), .B(n14046), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n14043) );
  NAND2_X1 U17254 ( .A1(n14070), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14042) );
  NAND2_X1 U17255 ( .A1(n14043), .A2(n14042), .ZN(n15925) );
  INV_X1 U17256 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n21168) );
  NAND2_X1 U17257 ( .A1(n14044), .A2(n21168), .ZN(n14048) );
  INV_X1 U17258 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16062) );
  NAND2_X1 U17259 ( .A1(n14067), .A2(n21168), .ZN(n14045) );
  OAI211_X1 U17260 ( .C1(n15910), .C2(n16062), .A(n14046), .B(n14045), .ZN(
        n14047) );
  AND2_X1 U17261 ( .A1(n14048), .A2(n14047), .ZN(n14180) );
  NAND2_X1 U17262 ( .A1(n15925), .A2(n14180), .ZN(n14049) );
  INV_X1 U17263 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14677) );
  NAND2_X1 U17264 ( .A1(n14046), .A2(n14677), .ZN(n14050) );
  OAI211_X1 U17265 ( .C1(n14070), .C2(P1_EBX_REG_24__SCAN_IN), .A(n14082), .B(
        n14050), .ZN(n14052) );
  INV_X1 U17266 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n20999) );
  NAND2_X1 U17267 ( .A1(n14062), .A2(n20999), .ZN(n14051) );
  NAND2_X1 U17268 ( .A1(n14052), .A2(n14051), .ZN(n14163) );
  NAND2_X1 U17269 ( .A1(n14182), .A2(n14163), .ZN(n14164) );
  INV_X1 U17270 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14649) );
  INV_X1 U17271 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n21193) );
  NAND2_X1 U17272 ( .A1(n14067), .A2(n21193), .ZN(n14053) );
  OAI211_X1 U17273 ( .C1(n15910), .C2(n14649), .A(n14046), .B(n14053), .ZN(
        n14054) );
  OAI21_X1 U17274 ( .B1(n14059), .B2(P1_EBX_REG_25__SCAN_IN), .A(n14054), .ZN(
        n14157) );
  INV_X1 U17275 ( .A(n14055), .ZN(n14156) );
  MUX2_X1 U17276 ( .A(n14062), .B(n14056), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n14058) );
  INV_X1 U17277 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14652) );
  NOR2_X1 U17278 ( .A1(n14067), .A2(n14652), .ZN(n14057) );
  NOR2_X1 U17279 ( .A1(n14058), .A2(n14057), .ZN(n14132) );
  MUX2_X1 U17280 ( .A(n14059), .B(n14082), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n14060) );
  OAI21_X1 U17281 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14071), .A(
        n14060), .ZN(n14061) );
  INV_X1 U17282 ( .A(n14061), .ZN(n14122) );
  INV_X1 U17283 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14279) );
  NAND2_X1 U17284 ( .A1(n14062), .A2(n14279), .ZN(n14066) );
  INV_X1 U17285 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14627) );
  NAND2_X1 U17286 ( .A1(n14046), .A2(n14627), .ZN(n14064) );
  NAND2_X1 U17287 ( .A1(n14067), .A2(n14279), .ZN(n14063) );
  NAND3_X1 U17288 ( .A1(n14064), .A2(n14082), .A3(n14063), .ZN(n14065) );
  NAND2_X1 U17289 ( .A1(n14066), .A2(n14065), .ZN(n14107) );
  OR2_X1 U17290 ( .A1(n14071), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14069) );
  INV_X1 U17291 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14103) );
  NAND2_X1 U17292 ( .A1(n14067), .A2(n14103), .ZN(n14068) );
  NAND2_X1 U17293 ( .A1(n14069), .A2(n14068), .ZN(n14081) );
  MUX2_X1 U17294 ( .A(n14081), .B(P1_EBX_REG_29__SCAN_IN), .S(n15910), .Z(
        n14099) );
  MUX2_X1 U17295 ( .A(n14082), .B(n14084), .S(n14098), .Z(n14073) );
  AOI22_X1 U17296 ( .A1(n14071), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n14070), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14072) );
  NAND2_X1 U17297 ( .A1(n14433), .A2(n20031), .ZN(n14080) );
  INV_X1 U17298 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n21227) );
  INV_X1 U17299 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n14473) );
  INV_X1 U17300 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21198) );
  INV_X1 U17301 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n15920) );
  INV_X1 U17302 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n15945) );
  INV_X1 U17303 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n21171) );
  NAND4_X1 U17304 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(P1_REIP_REG_12__SCAN_IN), .A4(P1_REIP_REG_11__SCAN_IN), .ZN(n14216) );
  INV_X1 U17305 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n21014) );
  INV_X1 U17306 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20988) );
  NOR3_X1 U17307 ( .A1(n14216), .A2(n21014), .A3(n20988), .ZN(n14206) );
  NAND3_X1 U17308 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n14205), .A3(n14206), 
        .ZN(n14192) );
  NOR4_X1 U17309 ( .A1(n15945), .A2(n14512), .A3(n21171), .A4(n14192), .ZN(
        n15930) );
  NAND2_X1 U17310 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n15930), .ZN(n15919) );
  NOR2_X1 U17311 ( .A1(n15920), .A2(n15919), .ZN(n14177) );
  NAND2_X1 U17312 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n14177), .ZN(n14168) );
  NOR2_X1 U17313 ( .A1(n21198), .A2(n14168), .ZN(n14155) );
  NAND2_X1 U17314 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n14155), .ZN(n14139) );
  NOR2_X1 U17315 ( .A1(n14473), .A2(n14139), .ZN(n14138) );
  NAND2_X1 U17316 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n14138), .ZN(n14112) );
  NOR2_X1 U17317 ( .A1(n21227), .A2(n14112), .ZN(n14100) );
  INV_X1 U17318 ( .A(n14100), .ZN(n14074) );
  AOI21_X1 U17319 ( .B1(n20069), .B2(n14074), .A(n20019), .ZN(n14115) );
  INV_X1 U17320 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n21183) );
  INV_X1 U17321 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21262) );
  OAI21_X1 U17322 ( .B1(n21183), .B2(n21262), .A(n20069), .ZN(n14075) );
  NAND2_X1 U17323 ( .A1(n14115), .A2(n14075), .ZN(n14089) );
  INV_X1 U17324 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n21233) );
  OAI22_X1 U17325 ( .A1(n20064), .A2(n21233), .B1(n14076), .B2(n20060), .ZN(
        n14078) );
  NAND3_X1 U17326 ( .A1(n20069), .A2(P1_REIP_REG_29__SCAN_IN), .A3(n14100), 
        .ZN(n14091) );
  NOR3_X1 U17327 ( .A1(n14091), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n21183), 
        .ZN(n14077) );
  AOI211_X1 U17328 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n14089), .A(n14078), 
        .B(n14077), .ZN(n14079) );
  OAI211_X1 U17329 ( .C1(n14594), .C2(n20073), .A(n14080), .B(n14079), .ZN(
        P1_U2809) );
  OAI22_X1 U17330 ( .A1(n14098), .A2(n14082), .B1(n9888), .B2(n14081), .ZN(
        n14083) );
  XOR2_X1 U17331 ( .A(n14084), .B(n14083), .Z(n14609) );
  NAND2_X1 U17332 ( .A1(n14442), .A2(n20031), .ZN(n14095) );
  INV_X1 U17333 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14088) );
  OAI22_X1 U17334 ( .A1(n14088), .A2(n20060), .B1(n20043), .B2(n14440), .ZN(
        n14093) );
  INV_X1 U17335 ( .A(n14089), .ZN(n14090) );
  AOI21_X1 U17336 ( .B1(n21183), .B2(n14091), .A(n14090), .ZN(n14092) );
  AOI211_X1 U17337 ( .C1(n20075), .C2(P1_EBX_REG_30__SCAN_IN), .A(n14093), .B(
        n14092), .ZN(n14094) );
  OAI211_X1 U17338 ( .C1(n20073), .C2(n14609), .A(n14095), .B(n14094), .ZN(
        P1_U2810) );
  OAI21_X1 U17339 ( .B1(n14096), .B2(n14097), .A(n14085), .ZN(n14451) );
  AOI21_X1 U17340 ( .B1(n14099), .B2(n9888), .A(n14098), .ZN(n14619) );
  NOR2_X1 U17341 ( .A1(n14115), .A2(n21262), .ZN(n14105) );
  AOI22_X1 U17342 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n20080), .B1(
        n20079), .B2(n14446), .ZN(n14102) );
  NAND3_X1 U17343 ( .A1(n20069), .A2(n14100), .A3(n21262), .ZN(n14101) );
  OAI211_X1 U17344 ( .C1(n20064), .C2(n14103), .A(n14102), .B(n14101), .ZN(
        n14104) );
  AOI211_X1 U17345 ( .C1(n14619), .C2(n20077), .A(n14105), .B(n14104), .ZN(
        n14106) );
  OAI21_X1 U17346 ( .B1(n14451), .B2(n15937), .A(n14106), .ZN(P1_U2811) );
  OR2_X1 U17347 ( .A1(n14124), .A2(n14107), .ZN(n14108) );
  NAND2_X1 U17348 ( .A1(n9888), .A2(n14108), .ZN(n14632) );
  AOI21_X1 U17349 ( .B1(n14110), .B2(n14109), .A(n14096), .ZN(n14460) );
  NAND2_X1 U17350 ( .A1(n14460), .A2(n20031), .ZN(n14119) );
  OAI22_X1 U17351 ( .A1(n14111), .A2(n20060), .B1(n20043), .B2(n14458), .ZN(
        n14117) );
  INV_X1 U17352 ( .A(n14112), .ZN(n14113) );
  AOI21_X1 U17353 ( .B1(n20069), .B2(n14113), .A(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n14114) );
  NOR2_X1 U17354 ( .A1(n14115), .A2(n14114), .ZN(n14116) );
  AOI211_X1 U17355 ( .C1(n20075), .C2(P1_EBX_REG_28__SCAN_IN), .A(n14117), .B(
        n14116), .ZN(n14118) );
  OAI211_X1 U17356 ( .C1(n20073), .C2(n14632), .A(n14119), .B(n14118), .ZN(
        P1_U2812) );
  OAI21_X1 U17357 ( .B1(n14120), .B2(n14121), .A(n14109), .ZN(n14469) );
  NOR2_X1 U17358 ( .A1(n14133), .A2(n14122), .ZN(n14123) );
  OR2_X1 U17359 ( .A1(n14124), .A2(n14123), .ZN(n14280) );
  INV_X1 U17360 ( .A(n14280), .ZN(n14641) );
  INV_X1 U17361 ( .A(n14138), .ZN(n14126) );
  AOI21_X1 U17362 ( .B1(n20069), .B2(n14126), .A(n20019), .ZN(n14137) );
  INV_X1 U17363 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21266) );
  INV_X1 U17364 ( .A(n14464), .ZN(n14125) );
  OAI22_X1 U17365 ( .A1(n14462), .A2(n20060), .B1(n20043), .B2(n14125), .ZN(
        n14128) );
  NOR3_X1 U17366 ( .A1(n20021), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14126), 
        .ZN(n14127) );
  AOI211_X1 U17367 ( .C1(P1_EBX_REG_27__SCAN_IN), .C2(n20075), .A(n14128), .B(
        n14127), .ZN(n14129) );
  OAI21_X1 U17368 ( .B1(n14137), .B2(n21266), .A(n14129), .ZN(n14130) );
  AOI21_X1 U17369 ( .B1(n14641), .B2(n20077), .A(n14130), .ZN(n14131) );
  OAI21_X1 U17370 ( .B1(n14469), .B2(n15937), .A(n14131), .ZN(P1_U2813) );
  AND2_X1 U17371 ( .A1(n14156), .A2(n14132), .ZN(n14134) );
  OR2_X1 U17372 ( .A1(n14134), .A2(n14133), .ZN(n14646) );
  AOI21_X1 U17373 ( .B1(n14136), .B2(n14149), .A(n14120), .ZN(n14477) );
  NAND2_X1 U17374 ( .A1(n14477), .A2(n20031), .ZN(n14148) );
  INV_X1 U17375 ( .A(n14137), .ZN(n14146) );
  NOR2_X1 U17376 ( .A1(n14139), .A2(n14138), .ZN(n14140) );
  NAND2_X1 U17377 ( .A1(n20069), .A2(n14140), .ZN(n14144) );
  NAND2_X1 U17378 ( .A1(n20075), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n14143) );
  INV_X1 U17379 ( .A(n14475), .ZN(n14141) );
  AOI22_X1 U17380 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n20080), .B1(
        n20079), .B2(n14141), .ZN(n14142) );
  NAND3_X1 U17381 ( .A1(n14144), .A2(n14143), .A3(n14142), .ZN(n14145) );
  AOI21_X1 U17382 ( .B1(n14146), .B2(P1_REIP_REG_26__SCAN_IN), .A(n14145), 
        .ZN(n14147) );
  OAI211_X1 U17383 ( .C1(n20073), .C2(n14646), .A(n14148), .B(n14147), .ZN(
        P1_U2814) );
  OAI21_X1 U17384 ( .B1(n14160), .B2(n14150), .A(n14149), .ZN(n14488) );
  NOR2_X1 U17385 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n20021), .ZN(n14154) );
  NAND2_X1 U17386 ( .A1(n20069), .A2(n14168), .ZN(n14151) );
  AND2_X1 U17387 ( .A1(n14151), .A2(n20059), .ZN(n14179) );
  NAND2_X1 U17388 ( .A1(n20069), .A2(n21198), .ZN(n14169) );
  INV_X1 U17389 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21212) );
  AOI21_X1 U17390 ( .B1(n14179), .B2(n14169), .A(n21212), .ZN(n14153) );
  OAI22_X1 U17391 ( .A1(n14485), .A2(n20060), .B1(n21193), .B2(n20064), .ZN(
        n14152) );
  AOI211_X1 U17392 ( .C1(n14155), .C2(n14154), .A(n14153), .B(n14152), .ZN(
        n14159) );
  AOI21_X1 U17393 ( .B1(n14157), .B2(n14164), .A(n14055), .ZN(n14661) );
  AOI22_X1 U17394 ( .A1(n14661), .A2(n20077), .B1(n14487), .B2(n20079), .ZN(
        n14158) );
  OAI211_X1 U17395 ( .C1(n14488), .C2(n15937), .A(n14159), .B(n14158), .ZN(
        P1_U2815) );
  AOI21_X1 U17396 ( .B1(n14161), .B2(n14174), .A(n14160), .ZN(n14162) );
  INV_X1 U17397 ( .A(n14162), .ZN(n14500) );
  OR2_X1 U17398 ( .A1(n14182), .A2(n14163), .ZN(n14165) );
  AND2_X1 U17399 ( .A1(n14165), .A2(n14164), .ZN(n14674) );
  NOR2_X1 U17400 ( .A1(n14179), .A2(n21198), .ZN(n14171) );
  AOI22_X1 U17401 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n20080), .B1(
        n20079), .B2(n14497), .ZN(n14167) );
  NAND2_X1 U17402 ( .A1(n20075), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n14166) );
  OAI211_X1 U17403 ( .C1(n14169), .C2(n14168), .A(n14167), .B(n14166), .ZN(
        n14170) );
  AOI211_X1 U17404 ( .C1(n14674), .C2(n20077), .A(n14171), .B(n14170), .ZN(
        n14172) );
  OAI21_X1 U17405 ( .B1(n14500), .B2(n15937), .A(n14172), .ZN(P1_U2816) );
  INV_X1 U17406 ( .A(n14174), .ZN(n14175) );
  AOI21_X1 U17407 ( .B1(n14176), .B2(n14173), .A(n14175), .ZN(n14507) );
  AOI21_X1 U17408 ( .B1(n20069), .B2(n14177), .A(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n14178) );
  OAI22_X1 U17409 ( .A1(n14179), .A2(n14178), .B1(n21168), .B2(n20064), .ZN(
        n14186) );
  INV_X1 U17410 ( .A(n15926), .ZN(n14181) );
  AOI21_X1 U17411 ( .B1(n14181), .B2(n15925), .A(n14180), .ZN(n14183) );
  OR2_X1 U17412 ( .A1(n14183), .A2(n14182), .ZN(n16057) );
  AOI22_X1 U17413 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n20080), .B1(
        n20079), .B2(n14503), .ZN(n14184) );
  OAI21_X1 U17414 ( .B1(n16057), .B2(n20073), .A(n14184), .ZN(n14185) );
  AOI211_X1 U17415 ( .C1(n14507), .C2(n20031), .A(n14186), .B(n14185), .ZN(
        n14187) );
  INV_X1 U17416 ( .A(n14187), .ZN(P1_U2817) );
  XNOR2_X1 U17417 ( .A(n14188), .B(n14288), .ZN(n14514) );
  OR2_X1 U17418 ( .A1(n14301), .A2(n14189), .ZN(n14190) );
  AND2_X1 U17419 ( .A1(n14291), .A2(n14190), .ZN(n16073) );
  INV_X1 U17420 ( .A(n14517), .ZN(n14191) );
  OAI22_X1 U17421 ( .A1(n20064), .A2(n21034), .B1(n14191), .B2(n20043), .ZN(
        n14196) );
  NOR2_X1 U17422 ( .A1(n20021), .A2(n14192), .ZN(n15946) );
  NAND2_X1 U17423 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n15946), .ZN(n15935) );
  AOI21_X1 U17424 ( .B1(n14192), .B2(n20069), .A(n20019), .ZN(n14207) );
  INV_X1 U17425 ( .A(n14207), .ZN(n15947) );
  AOI21_X1 U17426 ( .B1(n15946), .B2(n15945), .A(n15947), .ZN(n14194) );
  AOI21_X1 U17427 ( .B1(n20080), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n20048), .ZN(n14193) );
  OAI221_X1 U17428 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(n15935), .C1(n14512), 
        .C2(n14194), .A(n14193), .ZN(n14195) );
  AOI211_X1 U17429 ( .C1(n20077), .C2(n16073), .A(n14196), .B(n14195), .ZN(
        n14197) );
  OAI21_X1 U17430 ( .B1(n14514), .B2(n15937), .A(n14197), .ZN(P1_U2821) );
  OAI21_X1 U17431 ( .B1(n14198), .B2(n14200), .A(n14199), .ZN(n14534) );
  AND2_X1 U17432 ( .A1(n14311), .A2(n14201), .ZN(n14202) );
  NOR2_X1 U17433 ( .A1(n14299), .A2(n14202), .ZN(n16094) );
  INV_X1 U17434 ( .A(n14537), .ZN(n14204) );
  NAND2_X1 U17435 ( .A1(n20075), .A2(P1_EBX_REG_17__SCAN_IN), .ZN(n14203) );
  INV_X1 U17436 ( .A(n20048), .ZN(n14221) );
  OAI211_X1 U17437 ( .C1(n14204), .C2(n20043), .A(n14203), .B(n14221), .ZN(
        n14210) );
  NAND2_X1 U17438 ( .A1(n20069), .A2(n14205), .ZN(n14215) );
  INV_X1 U17439 ( .A(n14215), .ZN(n15969) );
  AOI21_X1 U17440 ( .B1(n14206), .B2(n15969), .A(P1_REIP_REG_17__SCAN_IN), 
        .ZN(n14208) );
  OAI22_X1 U17441 ( .A1(n14208), .A2(n14207), .B1(n14533), .B2(n20060), .ZN(
        n14209) );
  AOI211_X1 U17442 ( .C1(n16094), .C2(n20077), .A(n14210), .B(n14209), .ZN(
        n14211) );
  OAI21_X1 U17443 ( .B1(n14534), .B2(n15937), .A(n14211), .ZN(P1_U2823) );
  AOI21_X1 U17444 ( .B1(n14214), .B2(n14212), .A(n10303), .ZN(n14549) );
  INV_X1 U17445 ( .A(n14549), .ZN(n14394) );
  INV_X1 U17446 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n21016) );
  INV_X1 U17447 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20982) );
  NAND2_X1 U17448 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n14246) );
  OR3_X1 U17449 ( .A1(n20982), .A2(n14246), .A3(n14215), .ZN(n14233) );
  NOR2_X1 U17450 ( .A1(n21016), .A2(n14233), .ZN(n15956) );
  NAND2_X1 U17451 ( .A1(n20059), .A2(n20021), .ZN(n20074) );
  AOI21_X1 U17452 ( .B1(n14216), .B2(n20074), .A(n15974), .ZN(n15954) );
  AOI22_X1 U17453 ( .A1(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n20080), .B1(
        P1_EBX_REG_15__SCAN_IN), .B2(n20075), .ZN(n14217) );
  OAI21_X1 U17454 ( .B1(n15954), .B2(n20988), .A(n14217), .ZN(n14224) );
  INV_X1 U17455 ( .A(n14230), .ZN(n14219) );
  INV_X1 U17456 ( .A(n14309), .ZN(n14218) );
  AOI21_X1 U17457 ( .B1(n14220), .B2(n14219), .A(n14218), .ZN(n16101) );
  NAND2_X1 U17458 ( .A1(n16101), .A2(n20077), .ZN(n14222) );
  OAI211_X1 U17459 ( .C1(n14547), .C2(n20043), .A(n14222), .B(n14221), .ZN(
        n14223) );
  AOI211_X1 U17460 ( .C1(n15956), .C2(n20988), .A(n14224), .B(n14223), .ZN(
        n14225) );
  OAI21_X1 U17461 ( .B1(n14394), .B2(n15937), .A(n14225), .ZN(P1_U2825) );
  AOI21_X1 U17462 ( .B1(n14227), .B2(n14226), .A(n12003), .ZN(n16016) );
  INV_X1 U17463 ( .A(n16016), .ZN(n14397) );
  NOR2_X1 U17464 ( .A1(n14244), .A2(n14228), .ZN(n14229) );
  OR2_X1 U17465 ( .A1(n14230), .A2(n14229), .ZN(n16111) );
  OAI22_X1 U17466 ( .A1(n21236), .A2(n20064), .B1(n20073), .B2(n16111), .ZN(
        n14231) );
  AOI211_X1 U17467 ( .C1(n20080), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n20048), .B(n14231), .ZN(n14232) );
  INV_X1 U17468 ( .A(n14232), .ZN(n14235) );
  AOI21_X1 U17469 ( .B1(n21016), .B2(n14233), .A(n15954), .ZN(n14234) );
  AOI211_X1 U17470 ( .C1(n16015), .C2(n20079), .A(n14235), .B(n14234), .ZN(
        n14236) );
  OAI21_X1 U17471 ( .B1(n14397), .B2(n15937), .A(n14236), .ZN(P1_U2826) );
  OAI21_X1 U17472 ( .B1(n13560), .B2(n14238), .A(n14237), .ZN(n14404) );
  INV_X1 U17473 ( .A(n14403), .ZN(n14239) );
  OAI21_X1 U17474 ( .B1(n14404), .B2(n14239), .A(n14237), .ZN(n14325) );
  NAND2_X1 U17475 ( .A1(n14325), .A2(n14324), .ZN(n14323) );
  INV_X1 U17476 ( .A(n14240), .ZN(n14241) );
  AOI21_X1 U17477 ( .B1(n14323), .B2(n14241), .A(n11985), .ZN(n14561) );
  INV_X1 U17478 ( .A(n14561), .ZN(n14400) );
  AOI21_X1 U17479 ( .B1(n14246), .B2(n20074), .A(n15974), .ZN(n14242) );
  INV_X1 U17480 ( .A(n14242), .ZN(n15965) );
  AOI21_X1 U17481 ( .B1(n20080), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n20048), .ZN(n14243) );
  OAI21_X1 U17482 ( .B1(n20043), .B2(n14559), .A(n14243), .ZN(n14251) );
  AOI21_X1 U17483 ( .B1(n14245), .B2(n14322), .A(n14244), .ZN(n16124) );
  AOI22_X1 U17484 ( .A1(P1_EBX_REG_13__SCAN_IN), .A2(n20075), .B1(n20077), 
        .B2(n16124), .ZN(n14249) );
  INV_X1 U17485 ( .A(n14246), .ZN(n14247) );
  NAND3_X1 U17486 ( .A1(n14247), .A2(n20982), .A3(n15969), .ZN(n14248) );
  NAND2_X1 U17487 ( .A1(n14249), .A2(n14248), .ZN(n14250) );
  AOI211_X1 U17488 ( .C1(P1_REIP_REG_13__SCAN_IN), .C2(n15965), .A(n14251), 
        .B(n14250), .ZN(n14252) );
  OAI21_X1 U17489 ( .B1(n14400), .B2(n15937), .A(n14252), .ZN(P1_U2827) );
  INV_X1 U17490 ( .A(n14253), .ZN(n14257) );
  NAND2_X1 U17491 ( .A1(n14257), .A2(n11621), .ZN(n14254) );
  INV_X1 U17492 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n21230) );
  NAND4_X1 U17493 ( .A1(n20069), .A2(P1_REIP_REG_1__SCAN_IN), .A3(
        P1_REIP_REG_2__SCAN_IN), .A4(n21230), .ZN(n14265) );
  INV_X1 U17494 ( .A(n14255), .ZN(n14256) );
  NAND2_X1 U17495 ( .A1(n14257), .A2(n14256), .ZN(n20045) );
  INV_X1 U17496 ( .A(n20045), .ZN(n20078) );
  OAI221_X1 U17497 ( .B1(n20021), .B2(P1_REIP_REG_1__SCAN_IN), .C1(n20021), 
        .C2(P1_REIP_REG_2__SCAN_IN), .A(n20059), .ZN(n14258) );
  AOI22_X1 U17498 ( .A1(n20080), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n14258), .ZN(n14259) );
  OAI21_X1 U17499 ( .B1(n20043), .B2(n14260), .A(n14259), .ZN(n14261) );
  AOI21_X1 U17500 ( .B1(n20075), .B2(P1_EBX_REG_3__SCAN_IN), .A(n14261), .ZN(
        n14262) );
  OAI21_X1 U17501 ( .B1(n20073), .B2(n20178), .A(n14262), .ZN(n14263) );
  AOI21_X1 U17502 ( .B1(n20500), .B2(n20078), .A(n14263), .ZN(n14264) );
  OAI211_X1 U17503 ( .C1(n14266), .C2(n20087), .A(n14265), .B(n14264), .ZN(
        P1_U2837) );
  INV_X1 U17504 ( .A(n20087), .ZN(n20040) );
  NOR2_X1 U17505 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n20021), .ZN(n14267) );
  AOI22_X1 U17506 ( .A1(n20080), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        P1_REIP_REG_1__SCAN_IN), .B2(n14267), .ZN(n14268) );
  OAI21_X1 U17507 ( .B1(n20043), .B2(n14269), .A(n14268), .ZN(n14270) );
  AOI21_X1 U17508 ( .B1(n20075), .B2(P1_EBX_REG_2__SCAN_IN), .A(n14270), .ZN(
        n14271) );
  OAI21_X1 U17509 ( .B1(n20631), .B2(n20045), .A(n14271), .ZN(n14275) );
  INV_X1 U17510 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20889) );
  AOI21_X1 U17511 ( .B1(n20069), .B2(n20889), .A(n20019), .ZN(n14273) );
  INV_X1 U17512 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n21165) );
  OAI22_X1 U17513 ( .A1(n14273), .A2(n21165), .B1(n20073), .B2(n14272), .ZN(
        n14274) );
  AOI211_X1 U17514 ( .C1(n14276), .C2(n20040), .A(n14275), .B(n14274), .ZN(
        n14277) );
  INV_X1 U17515 ( .A(n14277), .ZN(P1_U2838) );
  OAI22_X1 U17516 ( .A1(n14594), .A2(n14316), .B1(n21233), .B2(n20101), .ZN(
        P1_U2841) );
  INV_X1 U17517 ( .A(n14442), .ZN(n14332) );
  INV_X1 U17518 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n21226) );
  OAI222_X1 U17519 ( .A1(n14326), .A2(n14332), .B1(n20101), .B2(n21226), .C1(
        n14609), .C2(n14316), .ZN(P1_U2842) );
  AOI22_X1 U17520 ( .A1(n14619), .A2(n20097), .B1(n14304), .B2(
        P1_EBX_REG_29__SCAN_IN), .ZN(n14278) );
  OAI21_X1 U17521 ( .B1(n14451), .B2(n14326), .A(n14278), .ZN(P1_U2843) );
  INV_X1 U17522 ( .A(n14460), .ZN(n14339) );
  OAI222_X1 U17523 ( .A1(n14279), .A2(n20101), .B1(n14316), .B2(n14632), .C1(
        n14339), .C2(n14326), .ZN(P1_U2844) );
  INV_X1 U17524 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14281) );
  OAI222_X1 U17525 ( .A1(n14281), .A2(n20101), .B1(n14316), .B2(n14280), .C1(
        n14469), .C2(n14326), .ZN(P1_U2845) );
  INV_X1 U17526 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n21259) );
  INV_X1 U17527 ( .A(n14477), .ZN(n14345) );
  OAI222_X1 U17528 ( .A1(n21259), .A2(n20101), .B1(n14316), .B2(n14646), .C1(
        n14345), .C2(n14326), .ZN(P1_U2846) );
  AOI22_X1 U17529 ( .A1(n14661), .A2(n20097), .B1(n14304), .B2(
        P1_EBX_REG_25__SCAN_IN), .ZN(n14282) );
  OAI21_X1 U17530 ( .B1(n14488), .B2(n14326), .A(n14282), .ZN(P1_U2847) );
  INV_X1 U17531 ( .A(n14674), .ZN(n14283) );
  OAI222_X1 U17532 ( .A1(n20999), .A2(n20101), .B1(n14316), .B2(n14283), .C1(
        n14500), .C2(n14326), .ZN(P1_U2848) );
  INV_X1 U17533 ( .A(n14507), .ZN(n14355) );
  OAI22_X1 U17534 ( .A1(n16057), .A2(n14316), .B1(n21168), .B2(n20101), .ZN(
        n14284) );
  INV_X1 U17535 ( .A(n14284), .ZN(n14285) );
  OAI21_X1 U17536 ( .B1(n14355), .B2(n14326), .A(n14285), .ZN(P1_U2849) );
  INV_X1 U17537 ( .A(n14286), .ZN(n14290) );
  OAI21_X1 U17538 ( .B1(n14188), .B2(n14288), .A(n14287), .ZN(n14289) );
  NAND2_X1 U17539 ( .A1(n14290), .A2(n14289), .ZN(n15998) );
  INV_X1 U17540 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14293) );
  OAI21_X1 U17541 ( .B1(n10278), .B2(n14292), .A(n9848), .ZN(n15936) );
  OAI222_X1 U17542 ( .A1(n15998), .A2(n14326), .B1(n20101), .B2(n14293), .C1(
        n15936), .C2(n14316), .ZN(P1_U2852) );
  NOR2_X1 U17543 ( .A1(n20101), .A2(n21034), .ZN(n14294) );
  AOI21_X1 U17544 ( .B1(n16073), .B2(n20097), .A(n14294), .ZN(n14295) );
  OAI21_X1 U17545 ( .B1(n14514), .B2(n14326), .A(n14295), .ZN(P1_U2853) );
  NAND2_X1 U17546 ( .A1(n14199), .A2(n14296), .ZN(n14297) );
  NOR2_X1 U17547 ( .A1(n14299), .A2(n14298), .ZN(n14300) );
  OR2_X1 U17548 ( .A1(n14301), .A2(n14300), .ZN(n16084) );
  OAI22_X1 U17549 ( .A1(n16084), .A2(n14316), .B1(n20959), .B2(n20101), .ZN(
        n14302) );
  AOI21_X1 U17550 ( .B1(n15950), .B2(n20098), .A(n14302), .ZN(n14303) );
  INV_X1 U17551 ( .A(n14303), .ZN(P1_U2854) );
  AOI22_X1 U17552 ( .A1(n16094), .A2(n20097), .B1(n14304), .B2(
        P1_EBX_REG_17__SCAN_IN), .ZN(n14305) );
  OAI21_X1 U17553 ( .B1(n14534), .B2(n14326), .A(n14305), .ZN(P1_U2855) );
  AOI21_X1 U17554 ( .B1(n14307), .B2(n14306), .A(n14198), .ZN(n16003) );
  NAND2_X1 U17555 ( .A1(n14309), .A2(n14308), .ZN(n14310) );
  NAND2_X1 U17556 ( .A1(n14311), .A2(n14310), .ZN(n15961) );
  OAI22_X1 U17557 ( .A1(n15961), .A2(n14316), .B1(n15953), .B2(n20101), .ZN(
        n14312) );
  AOI21_X1 U17558 ( .B1(n16003), .B2(n20098), .A(n14312), .ZN(n14313) );
  INV_X1 U17559 ( .A(n14313), .ZN(P1_U2856) );
  INV_X1 U17560 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14315) );
  INV_X1 U17561 ( .A(n16101), .ZN(n14314) );
  OAI222_X1 U17562 ( .A1(n14394), .A2(n14326), .B1(n20101), .B2(n14315), .C1(
        n14314), .C2(n14316), .ZN(P1_U2857) );
  OAI22_X1 U17563 ( .A1(n16111), .A2(n14316), .B1(n21236), .B2(n20101), .ZN(
        n14317) );
  AOI21_X1 U17564 ( .B1(n16016), .B2(n20098), .A(n14317), .ZN(n14318) );
  INV_X1 U17565 ( .A(n14318), .ZN(P1_U2858) );
  INV_X1 U17566 ( .A(n16124), .ZN(n14319) );
  OAI222_X1 U17567 ( .A1(n14400), .A2(n14326), .B1(n20101), .B2(n20998), .C1(
        n14316), .C2(n14319), .ZN(P1_U2859) );
  NAND2_X1 U17568 ( .A1(n15973), .A2(n14320), .ZN(n14321) );
  NAND2_X1 U17569 ( .A1(n14322), .A2(n14321), .ZN(n15962) );
  INV_X1 U17570 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n20972) );
  OAI21_X1 U17571 ( .B1(n14325), .B2(n14324), .A(n14323), .ZN(n15964) );
  OAI222_X1 U17572 ( .A1(n15962), .A2(n14316), .B1(n20101), .B2(n20972), .C1(
        n14326), .C2(n15964), .ZN(P1_U2860) );
  INV_X1 U17573 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20277) );
  OAI22_X1 U17574 ( .A1(n14362), .A2(n20277), .B1(n20975), .B2(n14391), .ZN(
        n14327) );
  INV_X1 U17575 ( .A(n14327), .ZN(n14331) );
  NOR3_X1 U17576 ( .A1(n14405), .A2(n20286), .A3(n14328), .ZN(n14329) );
  AOI22_X1 U17577 ( .A1(n14386), .A2(n14395), .B1(n14384), .B2(DATAI_30_), 
        .ZN(n14330) );
  OAI211_X1 U17578 ( .C1(n14332), .C2(n14409), .A(n14331), .B(n14330), .ZN(
        P1_U2874) );
  AOI22_X1 U17579 ( .A1(n14383), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n14405), .ZN(n14334) );
  AOI22_X1 U17580 ( .A1(n14386), .A2(n14398), .B1(n14384), .B2(DATAI_29_), 
        .ZN(n14333) );
  OAI211_X1 U17581 ( .C1(n14451), .C2(n14409), .A(n14334), .B(n14333), .ZN(
        P1_U2875) );
  INV_X1 U17582 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n14335) );
  OAI22_X1 U17583 ( .A1(n14362), .A2(n14335), .B1(n21275), .B2(n14391), .ZN(
        n14336) );
  INV_X1 U17584 ( .A(n14336), .ZN(n14338) );
  AOI22_X1 U17585 ( .A1(n14386), .A2(n14401), .B1(n14384), .B2(DATAI_28_), 
        .ZN(n14337) );
  OAI211_X1 U17586 ( .C1(n14339), .C2(n14409), .A(n14338), .B(n14337), .ZN(
        P1_U2876) );
  AOI22_X1 U17587 ( .A1(n14383), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n14405), .ZN(n14341) );
  AOI22_X1 U17588 ( .A1(n14386), .A2(n14406), .B1(n14384), .B2(DATAI_27_), 
        .ZN(n14340) );
  OAI211_X1 U17589 ( .C1(n14469), .C2(n14409), .A(n14341), .B(n14340), .ZN(
        P1_U2877) );
  AOI22_X1 U17590 ( .A1(n14383), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n14405), .ZN(n14344) );
  AOI22_X1 U17591 ( .A1(n14386), .A2(n14342), .B1(n14384), .B2(DATAI_26_), 
        .ZN(n14343) );
  OAI211_X1 U17592 ( .C1(n14345), .C2(n14409), .A(n14344), .B(n14343), .ZN(
        P1_U2878) );
  AOI22_X1 U17593 ( .A1(n14383), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n14405), .ZN(n14348) );
  AOI22_X1 U17594 ( .A1(n14386), .A2(n14346), .B1(n14384), .B2(DATAI_25_), 
        .ZN(n14347) );
  OAI211_X1 U17595 ( .C1(n14488), .C2(n14409), .A(n14348), .B(n14347), .ZN(
        P1_U2879) );
  AOI22_X1 U17596 ( .A1(n14383), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n14405), .ZN(n14351) );
  AOI22_X1 U17597 ( .A1(n14386), .A2(n14349), .B1(n14384), .B2(DATAI_24_), 
        .ZN(n14350) );
  OAI211_X1 U17598 ( .C1(n14500), .C2(n14409), .A(n14351), .B(n14350), .ZN(
        P1_U2880) );
  AOI22_X1 U17599 ( .A1(n14383), .A2(BUF1_REG_23__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n14405), .ZN(n14354) );
  AOI22_X1 U17600 ( .A1(n14386), .A2(n14352), .B1(n14384), .B2(DATAI_23_), 
        .ZN(n14353) );
  OAI211_X1 U17601 ( .C1(n14355), .C2(n14409), .A(n14354), .B(n14353), .ZN(
        P1_U2881) );
  OAI21_X1 U17602 ( .B1(n14357), .B2(n14356), .A(n14173), .ZN(n15924) );
  INV_X1 U17603 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20280) );
  OAI22_X1 U17604 ( .A1(n14362), .A2(n20280), .B1(n21244), .B2(n14391), .ZN(
        n14359) );
  INV_X1 U17605 ( .A(n14386), .ZN(n14365) );
  NOR2_X1 U17606 ( .A1(n14365), .A2(n20279), .ZN(n14358) );
  AOI211_X1 U17607 ( .C1(n14384), .C2(DATAI_22_), .A(n14359), .B(n14358), .ZN(
        n14360) );
  OAI21_X1 U17608 ( .B1(n15924), .B2(n14409), .A(n14360), .ZN(P1_U2882) );
  XOR2_X1 U17609 ( .A(n14361), .B(n14286), .Z(n15992) );
  INV_X1 U17610 ( .A(n15992), .ZN(n14369) );
  INV_X1 U17611 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20273) );
  NOR2_X1 U17612 ( .A1(n14362), .A2(n20273), .ZN(n14367) );
  INV_X1 U17613 ( .A(n14384), .ZN(n14364) );
  INV_X1 U17614 ( .A(DATAI_21_), .ZN(n14363) );
  OAI22_X1 U17615 ( .A1(n20272), .A2(n14365), .B1(n14364), .B2(n14363), .ZN(
        n14366) );
  AOI211_X1 U17616 ( .C1(n14405), .C2(P1_EAX_REG_21__SCAN_IN), .A(n14367), .B(
        n14366), .ZN(n14368) );
  OAI21_X1 U17617 ( .B1(n14369), .B2(n14409), .A(n14368), .ZN(P1_U2883) );
  AOI22_X1 U17618 ( .A1(n14383), .A2(BUF1_REG_20__SCAN_IN), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(n14405), .ZN(n14372) );
  AOI22_X1 U17619 ( .A1(n14386), .A2(n14370), .B1(n14384), .B2(DATAI_20_), 
        .ZN(n14371) );
  OAI211_X1 U17620 ( .C1(n15998), .C2(n14409), .A(n14372), .B(n14371), .ZN(
        P1_U2884) );
  AOI22_X1 U17621 ( .A1(n14383), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n14405), .ZN(n14375) );
  AOI22_X1 U17622 ( .A1(n14386), .A2(n14373), .B1(n14384), .B2(DATAI_19_), 
        .ZN(n14374) );
  OAI211_X1 U17623 ( .C1(n14514), .C2(n14409), .A(n14375), .B(n14374), .ZN(
        P1_U2885) );
  INV_X1 U17624 ( .A(n15950), .ZN(n14379) );
  AOI22_X1 U17625 ( .A1(n14383), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n14405), .ZN(n14378) );
  AOI22_X1 U17626 ( .A1(n14386), .A2(n14376), .B1(n14384), .B2(DATAI_18_), 
        .ZN(n14377) );
  OAI211_X1 U17627 ( .C1(n14379), .C2(n14409), .A(n14378), .B(n14377), .ZN(
        P1_U2886) );
  AOI22_X1 U17628 ( .A1(n14383), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n14405), .ZN(n14382) );
  AOI22_X1 U17629 ( .A1(n14386), .A2(n14380), .B1(n14384), .B2(DATAI_17_), 
        .ZN(n14381) );
  OAI211_X1 U17630 ( .C1(n14534), .C2(n14409), .A(n14382), .B(n14381), .ZN(
        P1_U2887) );
  INV_X1 U17631 ( .A(n16003), .ZN(n14389) );
  AOI22_X1 U17632 ( .A1(n14383), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n14405), .ZN(n14388) );
  AOI22_X1 U17633 ( .A1(n14386), .A2(n14385), .B1(n14384), .B2(DATAI_16_), 
        .ZN(n14387) );
  OAI211_X1 U17634 ( .C1(n14389), .C2(n14409), .A(n14388), .B(n14387), .ZN(
        P1_U2888) );
  OAI222_X1 U17635 ( .A1(n14394), .A2(n14409), .B1(n14393), .B2(n14392), .C1(
        n14391), .C2(n14390), .ZN(P1_U2889) );
  AOI22_X1 U17636 ( .A1(n14407), .A2(n14395), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n14405), .ZN(n14396) );
  OAI21_X1 U17637 ( .B1(n14397), .B2(n14409), .A(n14396), .ZN(P1_U2890) );
  AOI22_X1 U17638 ( .A1(n14407), .A2(n14398), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n14405), .ZN(n14399) );
  OAI21_X1 U17639 ( .B1(n14400), .B2(n14409), .A(n14399), .ZN(P1_U2891) );
  AOI22_X1 U17640 ( .A1(n14407), .A2(n14401), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n14405), .ZN(n14402) );
  OAI21_X1 U17641 ( .B1(n15964), .B2(n14409), .A(n14402), .ZN(P1_U2892) );
  XNOR2_X1 U17642 ( .A(n14404), .B(n14403), .ZN(n16029) );
  INV_X1 U17643 ( .A(n16029), .ZN(n14410) );
  AOI22_X1 U17644 ( .A1(n14407), .A2(n14406), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n14405), .ZN(n14408) );
  OAI21_X1 U17645 ( .B1(n14410), .B2(n14409), .A(n14408), .ZN(P1_U2893) );
  NAND2_X1 U17646 ( .A1(n13498), .A2(n16156), .ZN(n14412) );
  INV_X1 U17647 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16118) );
  NAND2_X1 U17648 ( .A1(n13498), .A2(n16118), .ZN(n14413) );
  NAND2_X1 U17649 ( .A1(n16008), .A2(n14413), .ZN(n14557) );
  INV_X1 U17650 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14713) );
  NAND2_X1 U17651 ( .A1(n13498), .A2(n14713), .ZN(n14555) );
  NAND2_X1 U17652 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14414) );
  NAND2_X1 U17653 ( .A1(n13498), .A2(n14414), .ZN(n14553) );
  NAND2_X1 U17654 ( .A1(n14555), .A2(n14553), .ZN(n14415) );
  NOR2_X1 U17655 ( .A1(n14557), .A2(n14415), .ZN(n16010) );
  NAND2_X1 U17656 ( .A1(n13498), .A2(n16110), .ZN(n14416) );
  NAND2_X1 U17657 ( .A1(n16010), .A2(n14416), .ZN(n14539) );
  OR2_X1 U17658 ( .A1(n13498), .A2(n16110), .ZN(n14417) );
  INV_X1 U17659 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14418) );
  OR2_X1 U17660 ( .A1(n13498), .A2(n14418), .ZN(n14543) );
  NAND2_X1 U17661 ( .A1(n13498), .A2(n14418), .ZN(n14691) );
  NAND2_X1 U17662 ( .A1(n14527), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14420) );
  NOR2_X1 U17663 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14551) );
  AND2_X1 U17664 ( .A1(n14551), .A2(n14713), .ZN(n14419) );
  NOR2_X1 U17665 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14421) );
  XNOR2_X1 U17666 ( .A(n16012), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14519) );
  INV_X1 U17667 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16078) );
  NAND2_X1 U17668 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14422) );
  NAND2_X1 U17669 ( .A1(n16078), .A2(n16089), .ZN(n14423) );
  INV_X1 U17670 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15892) );
  INV_X1 U17671 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15893) );
  NAND2_X1 U17672 ( .A1(n15892), .A2(n15893), .ZN(n14424) );
  NOR2_X1 U17673 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14479) );
  NAND2_X1 U17674 ( .A1(n14479), .A2(n14649), .ZN(n14425) );
  NAND2_X1 U17675 ( .A1(n14481), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14427) );
  AND2_X1 U17676 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14650) );
  NAND2_X1 U17677 ( .A1(n14650), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14653) );
  NAND2_X1 U17678 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14601) );
  XNOR2_X1 U17679 ( .A(n14429), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14608) );
  INV_X1 U17680 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21257) );
  NOR2_X1 U17681 ( .A1(n20207), .A2(n21257), .ZN(n14604) );
  AOI21_X1 U17682 ( .B1(n20151), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14604), .ZN(n14430) );
  OAI21_X1 U17683 ( .B1(n20164), .B2(n14431), .A(n14430), .ZN(n14432) );
  AOI21_X1 U17684 ( .B1(n14433), .B2(n20158), .A(n14432), .ZN(n14434) );
  OAI21_X1 U17685 ( .B1(n14608), .B2(n19988), .A(n14434), .ZN(P1_U2968) );
  NAND2_X1 U17686 ( .A1(n13498), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14436) );
  OAI21_X1 U17687 ( .B1(n14437), .B2(n14436), .A(n14435), .ZN(n14438) );
  XNOR2_X1 U17688 ( .A(n14438), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14616) );
  NOR2_X1 U17689 ( .A1(n20207), .A2(n21183), .ZN(n14613) );
  AOI21_X1 U17690 ( .B1(n20151), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14613), .ZN(n14439) );
  OAI21_X1 U17691 ( .B1(n20164), .B2(n14440), .A(n14439), .ZN(n14441) );
  AOI21_X1 U17692 ( .B1(n14442), .B2(n20158), .A(n14441), .ZN(n14443) );
  OAI21_X1 U17693 ( .B1(n14616), .B2(n19988), .A(n14443), .ZN(P1_U2969) );
  NAND2_X1 U17694 ( .A1(n20150), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14620) );
  OAI21_X1 U17695 ( .B1(n16041), .B2(n14444), .A(n14620), .ZN(n14445) );
  AOI21_X1 U17696 ( .B1(n14446), .B2(n16037), .A(n14445), .ZN(n14450) );
  XNOR2_X1 U17697 ( .A(n16012), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14447) );
  NAND2_X1 U17698 ( .A1(n14617), .A2(n20159), .ZN(n14449) );
  OAI211_X1 U17699 ( .C1(n14451), .C2(n15997), .A(n14450), .B(n14449), .ZN(
        P1_U2970) );
  NAND2_X1 U17700 ( .A1(n14452), .A2(n14652), .ZN(n14455) );
  NAND2_X1 U17701 ( .A1(n13498), .A2(n14653), .ZN(n14470) );
  NAND3_X1 U17702 ( .A1(n14502), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n14470), .ZN(n14454) );
  MUX2_X1 U17703 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n14652), .S(
        n13498), .Z(n14453) );
  AOI21_X1 U17704 ( .B1(n14455), .B2(n14454), .A(n14453), .ZN(n14456) );
  NOR2_X1 U17705 ( .A1(n20207), .A2(n21227), .ZN(n14628) );
  AOI21_X1 U17706 ( .B1(n20151), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14628), .ZN(n14457) );
  OAI21_X1 U17707 ( .B1(n20164), .B2(n14458), .A(n14457), .ZN(n14459) );
  AOI21_X1 U17708 ( .B1(n14460), .B2(n20158), .A(n14459), .ZN(n14461) );
  OAI21_X1 U17709 ( .B1(n19988), .B2(n14633), .A(n14461), .ZN(P1_U2971) );
  NOR2_X1 U17710 ( .A1(n20207), .A2(n21266), .ZN(n14637) );
  NOR2_X1 U17711 ( .A1(n16041), .A2(n14462), .ZN(n14463) );
  AOI211_X1 U17712 ( .C1(n16037), .C2(n14464), .A(n14637), .B(n14463), .ZN(
        n14468) );
  OAI211_X1 U17713 ( .C1(n14469), .C2(n15997), .A(n14468), .B(n14467), .ZN(
        P1_U2972) );
  INV_X1 U17714 ( .A(n14502), .ZN(n14480) );
  NOR2_X1 U17715 ( .A1(n14480), .A2(n16024), .ZN(n14471) );
  OAI21_X1 U17716 ( .B1(n14471), .B2(n14452), .A(n14470), .ZN(n14472) );
  XNOR2_X1 U17717 ( .A(n14472), .B(n14652), .ZN(n14658) );
  NOR2_X1 U17718 ( .A1(n20207), .A2(n14473), .ZN(n14647) );
  AOI21_X1 U17719 ( .B1(n20151), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n14647), .ZN(n14474) );
  OAI21_X1 U17720 ( .B1(n20164), .B2(n14475), .A(n14474), .ZN(n14476) );
  AOI21_X1 U17721 ( .B1(n14477), .B2(n20158), .A(n14476), .ZN(n14478) );
  OAI21_X1 U17722 ( .B1(n19988), .B2(n14658), .A(n14478), .ZN(P1_U2973) );
  NAND2_X1 U17723 ( .A1(n14480), .A2(n14479), .ZN(n14483) );
  AND2_X1 U17724 ( .A1(n14481), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14493) );
  NAND2_X1 U17725 ( .A1(n14493), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14482) );
  MUX2_X1 U17726 ( .A(n14483), .B(n14482), .S(n13498), .Z(n14484) );
  XNOR2_X1 U17727 ( .A(n14484), .B(n14649), .ZN(n14665) );
  NOR2_X1 U17728 ( .A1(n20207), .A2(n21212), .ZN(n14660) );
  NOR2_X1 U17729 ( .A1(n16041), .A2(n14485), .ZN(n14486) );
  AOI211_X1 U17730 ( .C1(n16037), .C2(n14487), .A(n14660), .B(n14486), .ZN(
        n14491) );
  INV_X1 U17731 ( .A(n14488), .ZN(n14489) );
  NAND2_X1 U17732 ( .A1(n14489), .A2(n20158), .ZN(n14490) );
  OAI211_X1 U17733 ( .C1(n14665), .C2(n19988), .A(n14491), .B(n14490), .ZN(
        P1_U2974) );
  NOR2_X1 U17734 ( .A1(n14493), .A2(n14502), .ZN(n14492) );
  MUX2_X1 U17735 ( .A(n14493), .B(n14492), .S(n16024), .Z(n14494) );
  XNOR2_X1 U17736 ( .A(n14494), .B(n14677), .ZN(n14670) );
  NAND2_X1 U17737 ( .A1(n14670), .A2(n20159), .ZN(n14499) );
  NOR2_X1 U17738 ( .A1(n20207), .A2(n21198), .ZN(n14673) );
  NOR2_X1 U17739 ( .A1(n16041), .A2(n14495), .ZN(n14496) );
  AOI211_X1 U17740 ( .C1(n16037), .C2(n14497), .A(n14673), .B(n14496), .ZN(
        n14498) );
  OAI211_X1 U17741 ( .C1(n14500), .C2(n15997), .A(n14499), .B(n14498), .ZN(
        P1_U2975) );
  XNOR2_X1 U17742 ( .A(n16012), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14501) );
  XNOR2_X1 U17743 ( .A(n14502), .B(n14501), .ZN(n16056) );
  INV_X1 U17744 ( .A(n14503), .ZN(n14505) );
  AOI22_X1 U17745 ( .A1(n20151), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(
        n20150), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n14504) );
  OAI21_X1 U17746 ( .B1(n20164), .B2(n14505), .A(n14504), .ZN(n14506) );
  AOI21_X1 U17747 ( .B1(n14507), .B2(n20158), .A(n14506), .ZN(n14508) );
  OAI21_X1 U17748 ( .B1(n16056), .B2(n19988), .A(n14508), .ZN(P1_U2976) );
  NAND2_X1 U17749 ( .A1(n14509), .A2(n16089), .ZN(n14510) );
  MUX2_X1 U17750 ( .A(n14510), .B(n14509), .S(n13498), .Z(n14511) );
  XNOR2_X1 U17751 ( .A(n14511), .B(n16078), .ZN(n16072) );
  INV_X1 U17752 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n14512) );
  OAI22_X1 U17753 ( .A1(n16041), .A2(n14513), .B1(n20207), .B2(n14512), .ZN(
        n14516) );
  NOR2_X1 U17754 ( .A1(n14514), .A2(n15997), .ZN(n14515) );
  AOI211_X1 U17755 ( .C1(n16037), .C2(n14517), .A(n14516), .B(n14515), .ZN(
        n14518) );
  OAI21_X1 U17756 ( .B1(n19988), .B2(n16072), .A(n14518), .ZN(P1_U2980) );
  OAI21_X1 U17757 ( .B1(n14520), .B2(n14519), .A(n14509), .ZN(n16085) );
  AOI22_X1 U17758 ( .A1(n20151), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n20150), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n14521) );
  OAI21_X1 U17759 ( .B1(n20164), .B2(n15948), .A(n14521), .ZN(n14522) );
  AOI21_X1 U17760 ( .B1(n15950), .B2(n20158), .A(n14522), .ZN(n14523) );
  OAI21_X1 U17761 ( .B1(n19988), .B2(n16085), .A(n14523), .ZN(P1_U2981) );
  NAND2_X1 U17762 ( .A1(n16024), .A2(n16090), .ZN(n14529) );
  NAND2_X1 U17763 ( .A1(n16025), .A2(n14525), .ZN(n16011) );
  INV_X1 U17764 ( .A(n14526), .ZN(n14692) );
  OAI21_X1 U17765 ( .B1(n16011), .B2(n14692), .A(n14527), .ZN(n14528) );
  MUX2_X1 U17766 ( .A(n16024), .B(n14529), .S(n14528), .Z(n14531) );
  INV_X1 U17767 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14530) );
  XNOR2_X1 U17768 ( .A(n14531), .B(n14530), .ZN(n16093) );
  INV_X1 U17769 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n14532) );
  OAI22_X1 U17770 ( .A1(n16041), .A2(n14533), .B1(n20207), .B2(n14532), .ZN(
        n14536) );
  NOR2_X1 U17771 ( .A1(n14534), .A2(n15997), .ZN(n14535) );
  AOI211_X1 U17772 ( .C1(n16037), .C2(n14537), .A(n14536), .B(n14535), .ZN(
        n14538) );
  OAI21_X1 U17773 ( .B1(n19988), .B2(n16093), .A(n14538), .ZN(P1_U2982) );
  INV_X1 U17774 ( .A(n16011), .ZN(n14540) );
  NOR2_X1 U17775 ( .A1(n14540), .A2(n14539), .ZN(n14693) );
  INV_X1 U17776 ( .A(n14541), .ZN(n14542) );
  NOR2_X1 U17777 ( .A1(n14693), .A2(n14542), .ZN(n14545) );
  NAND2_X1 U17778 ( .A1(n14543), .A2(n14691), .ZN(n14544) );
  XNOR2_X1 U17779 ( .A(n14545), .B(n14544), .ZN(n16100) );
  AOI22_X1 U17780 ( .A1(n20151), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20150), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n14546) );
  OAI21_X1 U17781 ( .B1(n20164), .B2(n14547), .A(n14546), .ZN(n14548) );
  AOI21_X1 U17782 ( .B1(n14549), .B2(n20158), .A(n14548), .ZN(n14550) );
  OAI21_X1 U17783 ( .B1(n16100), .B2(n19988), .A(n14550), .ZN(P1_U2984) );
  INV_X1 U17784 ( .A(n16025), .ZN(n14564) );
  INV_X1 U17785 ( .A(n14551), .ZN(n14552) );
  AOI22_X1 U17786 ( .A1(n14564), .A2(n14553), .B1(n16024), .B2(n14552), .ZN(
        n14711) );
  INV_X1 U17787 ( .A(n14555), .ZN(n14554) );
  AOI21_X1 U17788 ( .B1(n16024), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n14554), .ZN(n14710) );
  NAND2_X1 U17789 ( .A1(n14711), .A2(n14710), .ZN(n14709) );
  NAND2_X1 U17790 ( .A1(n14709), .A2(n14555), .ZN(n14556) );
  XOR2_X1 U17791 ( .A(n14557), .B(n14556), .Z(n16123) );
  INV_X1 U17792 ( .A(n16123), .ZN(n14563) );
  AOI22_X1 U17793 ( .A1(n20151), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n20150), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n14558) );
  OAI21_X1 U17794 ( .B1(n20164), .B2(n14559), .A(n14558), .ZN(n14560) );
  AOI21_X1 U17795 ( .B1(n14561), .B2(n20158), .A(n14560), .ZN(n14562) );
  OAI21_X1 U17796 ( .B1(n14563), .B2(n19988), .A(n14562), .ZN(P1_U2986) );
  NAND2_X1 U17797 ( .A1(n14567), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14566) );
  XNOR2_X1 U17798 ( .A(n14564), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14565) );
  MUX2_X1 U17799 ( .A(n14566), .B(n14565), .S(n13498), .Z(n14570) );
  INV_X1 U17800 ( .A(n14567), .ZN(n14569) );
  INV_X1 U17801 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14568) );
  NAND3_X1 U17802 ( .A1(n14569), .A2(n16024), .A3(n14568), .ZN(n16027) );
  NAND2_X1 U17803 ( .A1(n14570), .A2(n16027), .ZN(n16143) );
  INV_X1 U17804 ( .A(n16143), .ZN(n14576) );
  AOI22_X1 U17805 ( .A1(n20151), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n20150), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14571) );
  OAI21_X1 U17806 ( .B1(n20164), .B2(n14572), .A(n14571), .ZN(n14573) );
  AOI21_X1 U17807 ( .B1(n14574), .B2(n20158), .A(n14573), .ZN(n14575) );
  OAI21_X1 U17808 ( .B1(n14576), .B2(n19988), .A(n14575), .ZN(P1_U2989) );
  INV_X1 U17809 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14592) );
  INV_X1 U17810 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14591) );
  NAND2_X1 U17811 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16067) );
  NOR2_X1 U17812 ( .A1(n15892), .A2(n16078), .ZN(n14583) );
  NOR2_X1 U17813 ( .A1(n14578), .A2(n14577), .ZN(n16137) );
  NAND3_X1 U17814 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16140) );
  NAND2_X1 U17815 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16144) );
  NOR2_X1 U17816 ( .A1(n16140), .A2(n16144), .ZN(n14706) );
  NAND2_X1 U17817 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n14706), .ZN(
        n14716) );
  NOR2_X1 U17818 ( .A1(n14713), .A2(n14716), .ZN(n14580) );
  AND2_X1 U17819 ( .A1(n16137), .A2(n14580), .ZN(n16120) );
  NAND4_X1 U17820 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16082) );
  NOR2_X1 U17821 ( .A1(n16089), .A2(n16082), .ZN(n14597) );
  AND2_X1 U17822 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14597), .ZN(
        n14682) );
  NAND2_X1 U17823 ( .A1(n16120), .A2(n14682), .ZN(n14684) );
  NAND2_X1 U17824 ( .A1(n14580), .A2(n14579), .ZN(n14681) );
  NOR2_X1 U17825 ( .A1(n16118), .A2(n14681), .ZN(n16109) );
  AOI21_X1 U17826 ( .B1(n14597), .B2(n16109), .A(n20195), .ZN(n14581) );
  AOI211_X1 U17827 ( .C1(n14705), .C2(n14684), .A(n14581), .B(n14696), .ZN(
        n16075) );
  AOI22_X1 U17828 ( .A1(n14583), .A2(n16075), .B1(n14582), .B2(n20165), .ZN(
        n16064) );
  AOI21_X1 U17829 ( .B1(n20206), .B2(n16067), .A(n16064), .ZN(n16063) );
  NAND2_X1 U17830 ( .A1(n20193), .A2(n16062), .ZN(n14584) );
  AND2_X1 U17831 ( .A1(n16063), .A2(n14584), .ZN(n14667) );
  NAND2_X1 U17832 ( .A1(n20193), .A2(n14677), .ZN(n14587) );
  INV_X1 U17833 ( .A(n14653), .ZN(n14585) );
  OR2_X1 U17834 ( .A1(n16117), .A2(n14585), .ZN(n14586) );
  OAI211_X1 U17835 ( .C1(n14650), .C2(n14680), .A(n14587), .B(n14586), .ZN(
        n14588) );
  INV_X1 U17836 ( .A(n14588), .ZN(n14589) );
  NAND2_X1 U17837 ( .A1(n14667), .A2(n14589), .ZN(n14662) );
  OR2_X1 U17838 ( .A1(n14662), .A2(n20206), .ZN(n14590) );
  INV_X1 U17839 ( .A(n14590), .ZN(n14593) );
  OR2_X1 U17840 ( .A1(n14662), .A2(n14652), .ZN(n14655) );
  OAI21_X1 U17841 ( .B1(n14655), .B2(n14649), .A(n14590), .ZN(n14645) );
  OAI21_X1 U17842 ( .B1(n14428), .B2(n14593), .A(n14645), .ZN(n14624) );
  AOI211_X1 U17843 ( .C1(n14592), .C2(n20206), .A(n14591), .B(n14624), .ZN(
        n14611) );
  NOR3_X1 U17844 ( .A1(n14611), .A2(n14593), .A3(n14602), .ZN(n14606) );
  NOR2_X1 U17845 ( .A1(n14594), .A2(n20171), .ZN(n14605) );
  NAND2_X1 U17846 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n16120), .ZN(
        n14697) );
  NOR2_X1 U17847 ( .A1(n14708), .A2(n14697), .ZN(n14669) );
  AND2_X1 U17848 ( .A1(n20193), .A2(n16109), .ZN(n14595) );
  AND4_X1 U17849 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14596) );
  NAND2_X1 U17850 ( .A1(n14597), .A2(n14596), .ZN(n14666) );
  INV_X1 U17851 ( .A(n14666), .ZN(n14598) );
  NAND2_X1 U17852 ( .A1(n16091), .A2(n14598), .ZN(n14671) );
  INV_X1 U17853 ( .A(n14671), .ZN(n14600) );
  NOR2_X1 U17854 ( .A1(n14653), .A2(n14652), .ZN(n14599) );
  NAND2_X1 U17855 ( .A1(n14600), .A2(n14599), .ZN(n14639) );
  NOR2_X1 U17856 ( .A1(n14639), .A2(n14601), .ZN(n14618) );
  AND4_X1 U17857 ( .A1(n14618), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n14602), .ZN(n14603) );
  NOR4_X1 U17858 ( .A1(n14606), .A2(n14605), .A3(n14604), .A4(n14603), .ZN(
        n14607) );
  OAI21_X1 U17859 ( .B1(n14608), .B2(n20196), .A(n14607), .ZN(P1_U3000) );
  INV_X1 U17860 ( .A(n14609), .ZN(n14614) );
  AOI21_X1 U17861 ( .B1(n14618), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14610) );
  NOR2_X1 U17862 ( .A1(n14611), .A2(n14610), .ZN(n14612) );
  AOI211_X1 U17863 ( .C1(n20214), .C2(n14614), .A(n14613), .B(n14612), .ZN(
        n14615) );
  OAI21_X1 U17864 ( .B1(n14616), .B2(n20196), .A(n14615), .ZN(P1_U3001) );
  INV_X1 U17865 ( .A(n14617), .ZN(n14626) );
  INV_X1 U17866 ( .A(n14618), .ZN(n14622) );
  NAND2_X1 U17867 ( .A1(n14619), .A2(n20214), .ZN(n14621) );
  OAI211_X1 U17868 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n14622), .A(
        n14621), .B(n14620), .ZN(n14623) );
  AOI21_X1 U17869 ( .B1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n14624), .A(
        n14623), .ZN(n14625) );
  OAI21_X1 U17870 ( .B1(n14626), .B2(n20196), .A(n14625), .ZN(P1_U3002) );
  INV_X1 U17871 ( .A(n14645), .ZN(n14635) );
  INV_X1 U17872 ( .A(n14639), .ZN(n14630) );
  XNOR2_X1 U17873 ( .A(n14627), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14629) );
  AOI21_X1 U17874 ( .B1(n14630), .B2(n14629), .A(n14628), .ZN(n14631) );
  OAI21_X1 U17875 ( .B1(n14632), .B2(n20171), .A(n14631), .ZN(n14634) );
  INV_X1 U17876 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14644) );
  NAND2_X1 U17877 ( .A1(n14636), .A2(n20208), .ZN(n14643) );
  INV_X1 U17878 ( .A(n14637), .ZN(n14638) );
  OAI21_X1 U17879 ( .B1(n14639), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14638), .ZN(n14640) );
  AOI21_X1 U17880 ( .B1(n14641), .B2(n20214), .A(n14640), .ZN(n14642) );
  OAI211_X1 U17881 ( .C1(n14645), .C2(n14644), .A(n14643), .B(n14642), .ZN(
        P1_U3004) );
  INV_X1 U17882 ( .A(n14646), .ZN(n14648) );
  AOI21_X1 U17883 ( .B1(n14648), .B2(n20214), .A(n14647), .ZN(n14657) );
  NAND2_X1 U17884 ( .A1(n14650), .A2(n14649), .ZN(n14651) );
  NOR2_X1 U17885 ( .A1(n14671), .A2(n14651), .ZN(n14659) );
  OAI21_X1 U17886 ( .B1(n14671), .B2(n14653), .A(n14652), .ZN(n14654) );
  OAI21_X1 U17887 ( .B1(n14655), .B2(n14659), .A(n14654), .ZN(n14656) );
  OAI211_X1 U17888 ( .C1(n14658), .C2(n20196), .A(n14657), .B(n14656), .ZN(
        P1_U3005) );
  AOI211_X1 U17889 ( .C1(n14661), .C2(n20214), .A(n14660), .B(n14659), .ZN(
        n14664) );
  NAND2_X1 U17890 ( .A1(n14662), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14663) );
  OAI211_X1 U17891 ( .C1(n14665), .C2(n20196), .A(n14664), .B(n14663), .ZN(
        P1_U3006) );
  NOR2_X1 U17892 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n14666), .ZN(
        n16055) );
  INV_X1 U17893 ( .A(n14667), .ZN(n14668) );
  AOI21_X1 U17894 ( .B1(n14669), .B2(n16055), .A(n14668), .ZN(n14678) );
  NAND2_X1 U17895 ( .A1(n14670), .A2(n20208), .ZN(n14676) );
  NOR3_X1 U17896 ( .A1(n14671), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n16062), .ZN(n14672) );
  AOI211_X1 U17897 ( .C1(n14674), .C2(n20214), .A(n14673), .B(n14672), .ZN(
        n14675) );
  OAI211_X1 U17898 ( .C1(n14678), .C2(n14677), .A(n14676), .B(n14675), .ZN(
        P1_U3007) );
  NAND2_X1 U17899 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n16120), .ZN(
        n14679) );
  OAI22_X1 U17900 ( .A1(n20195), .A2(n14681), .B1(n14680), .B2(n14679), .ZN(
        n16121) );
  NAND2_X1 U17901 ( .A1(n14682), .A2(n16121), .ZN(n14683) );
  OAI221_X1 U17902 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n16117), 
        .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n14683), .A(n16075), .ZN(
        n14689) );
  NOR2_X1 U17903 ( .A1(n20207), .A2(n21171), .ZN(n16000) );
  OAI21_X1 U17904 ( .B1(n16117), .B2(n14684), .A(n14683), .ZN(n16079) );
  NAND2_X1 U17905 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n16079), .ZN(
        n15891) );
  NOR2_X1 U17906 ( .A1(n14685), .A2(n16024), .ZN(n15887) );
  NOR2_X1 U17907 ( .A1(n14686), .A2(n16012), .ZN(n15886) );
  NOR2_X1 U17908 ( .A1(n15887), .A2(n15886), .ZN(n14687) );
  XNOR2_X1 U17909 ( .A(n14687), .B(n15892), .ZN(n16002) );
  OAI22_X1 U17910 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15891), .B1(
        n16002), .B2(n20196), .ZN(n14688) );
  AOI211_X1 U17911 ( .C1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n14689), .A(
        n16000), .B(n14688), .ZN(n14690) );
  OAI21_X1 U17912 ( .B1(n20171), .B2(n15936), .A(n14690), .ZN(P1_U3011) );
  OAI21_X1 U17913 ( .B1(n14693), .B2(n14692), .A(n14691), .ZN(n14695) );
  XNOR2_X1 U17914 ( .A(n14695), .B(n14694), .ZN(n16004) );
  INV_X1 U17915 ( .A(n16004), .ZN(n14704) );
  INV_X1 U17916 ( .A(n16091), .ZN(n16083) );
  NOR3_X1 U17917 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n16083), .A3(
        n16110), .ZN(n16104) );
  AOI21_X1 U17918 ( .B1(n14705), .B2(n14697), .A(n14696), .ZN(n14698) );
  OAI21_X1 U17919 ( .B1(n16109), .B2(n20195), .A(n14698), .ZN(n16122) );
  AOI21_X1 U17920 ( .B1(n16110), .B2(n20206), .A(n16122), .ZN(n14699) );
  INV_X1 U17921 ( .A(n14699), .ZN(n16105) );
  OAI21_X1 U17922 ( .B1(n16104), .B2(n16105), .A(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14703) );
  NOR4_X1 U17923 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n16083), .A3(
        n16110), .A4(n14418), .ZN(n14701) );
  NOR2_X1 U17924 ( .A1(n15961), .A2(n20171), .ZN(n14700) );
  AOI211_X1 U17925 ( .C1(n20150), .C2(P1_REIP_REG_16__SCAN_IN), .A(n14701), 
        .B(n14700), .ZN(n14702) );
  OAI211_X1 U17926 ( .C1(n14704), .C2(n20196), .A(n14703), .B(n14702), .ZN(
        P1_U3015) );
  INV_X1 U17927 ( .A(n14705), .ZN(n20167) );
  AOI21_X1 U17928 ( .B1(n16137), .B2(n14706), .A(n20167), .ZN(n14707) );
  AOI211_X1 U17929 ( .C1(n20193), .C2(n14716), .A(n14707), .B(n16138), .ZN(
        n16136) );
  OAI21_X1 U17930 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n14708), .A(
        n16136), .ZN(n14718) );
  OAI21_X1 U17931 ( .B1(n14711), .B2(n14710), .A(n14709), .ZN(n14712) );
  INV_X1 U17932 ( .A(n14712), .ZN(n16023) );
  NAND2_X1 U17933 ( .A1(n14714), .A2(n14713), .ZN(n14715) );
  OAI22_X1 U17934 ( .A1(n16023), .A2(n20196), .B1(n14716), .B2(n14715), .ZN(
        n14717) );
  AOI21_X1 U17935 ( .B1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n14718), .A(
        n14717), .ZN(n14720) );
  NAND2_X1 U17936 ( .A1(n20150), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n14719) );
  OAI211_X1 U17937 ( .C1(n20171), .C2(n15962), .A(n14720), .B(n14719), .ZN(
        P1_U3019) );
  MUX2_X1 U17938 ( .A(n14721), .B(n20628), .S(n20766), .Z(n14722) );
  OAI21_X1 U17939 ( .B1(n14727), .B2(n20558), .A(n14722), .ZN(n14723) );
  MUX2_X1 U17940 ( .A(n14723), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        n14728), .Z(P1_U3477) );
  OR2_X1 U17941 ( .A1(n20766), .A2(n12580), .ZN(n14724) );
  AND2_X1 U17942 ( .A1(n14724), .A2(n20628), .ZN(n20472) );
  OAI21_X1 U17943 ( .B1(n14727), .B2(n20631), .A(n14726), .ZN(n14729) );
  MUX2_X1 U17944 ( .A(n14729), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        n14728), .Z(P1_U3476) );
  NOR3_X1 U17945 ( .A1(n14730), .A2(n14735), .A3(n11505), .ZN(n14733) );
  NOR2_X1 U17946 ( .A1(n20558), .A2(n14731), .ZN(n14732) );
  AOI211_X1 U17947 ( .C1(n14734), .C2(n11710), .A(n14733), .B(n14732), .ZN(
        n15854) );
  NOR3_X1 U17948 ( .A1(n11505), .A2(n14735), .A3(n15882), .ZN(n14736) );
  AOI21_X1 U17949 ( .B1(n14738), .B2(n14737), .A(n14736), .ZN(n14739) );
  OAI21_X1 U17950 ( .B1(n15854), .B2(n14744), .A(n14739), .ZN(n14740) );
  MUX2_X1 U17951 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14740), .S(
        n16185), .Z(P1_U3473) );
  INV_X1 U17952 ( .A(n14741), .ZN(n14745) );
  INV_X1 U17953 ( .A(n14742), .ZN(n14743) );
  OAI22_X1 U17954 ( .A1(n14745), .A2(n14744), .B1(n15882), .B2(n14743), .ZN(
        n14746) );
  MUX2_X1 U17955 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14746), .S(
        n16185), .Z(P1_U3469) );
  OAI21_X1 U17956 ( .B1(n19841), .B2(n19924), .A(n14747), .ZN(n14750) );
  NAND3_X1 U17957 ( .A1(n16347), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n19841), 
        .ZN(n14749) );
  MUX2_X1 U17958 ( .A(n14750), .B(n14749), .S(n14748), .Z(n14752) );
  OAI22_X1 U17959 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16364), .B1(n19851), 
        .B2(n19825), .ZN(n14751) );
  NAND2_X1 U17960 ( .A1(n14752), .A2(n14751), .ZN(n14755) );
  AOI21_X1 U17961 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n16363), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n14753) );
  AOI211_X1 U17962 ( .C1(n19835), .C2(n19218), .A(n14753), .B(n18911), .ZN(
        n14754) );
  MUX2_X1 U17963 ( .A(n14755), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n14754), 
        .Z(P2_U3610) );
  INV_X1 U17964 ( .A(n14825), .ZN(n14765) );
  NOR2_X1 U17965 ( .A1(n10145), .A2(n19831), .ZN(n18940) );
  NAND2_X1 U17966 ( .A1(n14756), .A2(n18940), .ZN(n14764) );
  INV_X1 U17967 ( .A(n14757), .ZN(n19123) );
  AOI22_X1 U17968 ( .A1(n19109), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19089), .ZN(n14758) );
  OAI21_X1 U17969 ( .B1(n19122), .B2(n14759), .A(n14758), .ZN(n14762) );
  NOR3_X1 U17970 ( .A1(n14760), .A2(P2_EBX_REG_30__SCAN_IN), .A3(n19106), .ZN(
        n14761) );
  AOI211_X1 U17971 ( .C1(n19036), .C2(n19123), .A(n14762), .B(n14761), .ZN(
        n14763) );
  OAI211_X1 U17972 ( .C1(n14765), .C2(n19115), .A(n14764), .B(n14763), .ZN(
        P2_U2824) );
  NAND2_X1 U17973 ( .A1(n14840), .A2(n14766), .ZN(n14767) );
  NAND2_X1 U17974 ( .A1(n14768), .A2(n14767), .ZN(n15239) );
  NAND2_X1 U17975 ( .A1(n9879), .A2(n14769), .ZN(n14770) );
  NAND2_X1 U17976 ( .A1(n14771), .A2(n14770), .ZN(n15236) );
  AOI22_X1 U17977 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n19080), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(n19109), .ZN(n14774) );
  INV_X1 U17978 ( .A(n19106), .ZN(n19081) );
  AOI22_X1 U17979 ( .A1(n14772), .A2(n19081), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19089), .ZN(n14773) );
  OAI211_X1 U17980 ( .C1(n15236), .C2(n19116), .A(n14774), .B(n14773), .ZN(
        n14777) );
  AOI211_X1 U17981 ( .C1(n15017), .C2(n9891), .A(n14775), .B(n19831), .ZN(
        n14776) );
  NOR2_X1 U17982 ( .A1(n14777), .A2(n14776), .ZN(n14778) );
  OAI21_X1 U17983 ( .B1(n15239), .B2(n19115), .A(n14778), .ZN(P2_U2826) );
  AOI211_X1 U17984 ( .C1(n15112), .C2(n14780), .A(n14779), .B(n19831), .ZN(
        n14782) );
  OAI22_X1 U17985 ( .A1(n15110), .A2(n19105), .B1(n10891), .B2(n19085), .ZN(
        n14781) );
  AOI211_X1 U17986 ( .C1(n19080), .C2(P2_REIP_REG_21__SCAN_IN), .A(n14782), 
        .B(n14781), .ZN(n14791) );
  NOR2_X1 U17987 ( .A1(n14784), .A2(n14783), .ZN(n14785) );
  OR2_X1 U17988 ( .A1(n12418), .A2(n14785), .ZN(n15331) );
  INV_X1 U17989 ( .A(n15331), .ZN(n14789) );
  NAND2_X1 U17990 ( .A1(n15339), .A2(n14786), .ZN(n14787) );
  AND2_X1 U17991 ( .A1(n14788), .A2(n14787), .ZN(n15328) );
  AOI22_X1 U17992 ( .A1(n14789), .A2(n11089), .B1(n15328), .B2(n19036), .ZN(
        n14790) );
  OAI211_X1 U17993 ( .C1(n14792), .C2(n19106), .A(n14791), .B(n14790), .ZN(
        P2_U2834) );
  XNOR2_X1 U17994 ( .A(n16296), .B(n14793), .ZN(n19154) );
  INV_X1 U17995 ( .A(n19154), .ZN(n15504) );
  NOR2_X1 U17996 ( .A1(n10145), .A2(n14794), .ZN(n14795) );
  XOR2_X1 U17997 ( .A(n14795), .B(n16263), .Z(n14796) );
  AOI22_X1 U17998 ( .A1(n15504), .A2(n19036), .B1(n19118), .B2(n14796), .ZN(
        n14802) );
  INV_X1 U17999 ( .A(n15499), .ZN(n16265) );
  INV_X1 U18000 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n14799) );
  OAI21_X1 U18001 ( .B1(n11008), .B2(n19085), .A(n19040), .ZN(n14797) );
  AOI21_X1 U18002 ( .B1(n19089), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n14797), .ZN(n14798) );
  OAI21_X1 U18003 ( .B1(n19122), .B2(n14799), .A(n14798), .ZN(n14800) );
  AOI21_X1 U18004 ( .B1(n16265), .B2(n11089), .A(n14800), .ZN(n14801) );
  OAI211_X1 U18005 ( .C1(n14803), .C2(n19106), .A(n14802), .B(n14801), .ZN(
        P2_U2846) );
  OAI211_X1 U18006 ( .C1(n14815), .C2(n14805), .A(n13535), .B(n14804), .ZN(
        n15537) );
  NOR2_X1 U18007 ( .A1(n13535), .A2(n19831), .ZN(n18934) );
  MUX2_X1 U18008 ( .A(n19089), .B(n18934), .S(n14806), .Z(n14809) );
  NOR2_X1 U18009 ( .A1(n19106), .A2(n14807), .ZN(n14808) );
  AOI211_X1 U18010 ( .C1(n19109), .C2(P2_EBX_REG_1__SCAN_IN), .A(n14809), .B(
        n14808), .ZN(n14811) );
  NAND2_X1 U18011 ( .A1(n19953), .A2(n19036), .ZN(n14810) );
  OAI211_X1 U18012 ( .C1(n19857), .C2(n19122), .A(n14811), .B(n14810), .ZN(
        n14813) );
  NOR2_X1 U18013 ( .A1(n19949), .A2(n14824), .ZN(n14812) );
  AOI211_X1 U18014 ( .C1(n11089), .C2(n13191), .A(n14813), .B(n14812), .ZN(
        n14814) );
  OAI21_X1 U18015 ( .B1(n15537), .B2(n19831), .A(n14814), .ZN(P2_U2854) );
  OAI21_X1 U18016 ( .B1(n19089), .B2(n18934), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14817) );
  INV_X1 U18017 ( .A(n14815), .ZN(n15526) );
  NAND2_X1 U18018 ( .A1(n15526), .A2(n18940), .ZN(n14816) );
  OAI211_X1 U18019 ( .C1(n19085), .C2(n12585), .A(n14817), .B(n14816), .ZN(
        n14819) );
  NOR2_X1 U18020 ( .A1(n19116), .A2(n16312), .ZN(n14818) );
  AOI211_X1 U18021 ( .C1(n19080), .C2(P2_REIP_REG_0__SCAN_IN), .A(n14819), .B(
        n14818), .ZN(n14820) );
  OAI21_X1 U18022 ( .B1(n19106), .B2(n14821), .A(n14820), .ZN(n14822) );
  AOI21_X1 U18023 ( .B1(n15525), .B2(n11089), .A(n14822), .ZN(n14823) );
  OAI21_X1 U18024 ( .B1(n19958), .B2(n14824), .A(n14823), .ZN(P2_U2855) );
  NAND2_X1 U18025 ( .A1(n14825), .A2(n14906), .ZN(n14826) );
  OAI21_X1 U18026 ( .B1(n14906), .B2(n14827), .A(n14826), .ZN(P2_U2856) );
  NAND2_X1 U18027 ( .A1(n14829), .A2(n14830), .ZN(n14922) );
  NAND3_X1 U18028 ( .A1(n14828), .A2(n14922), .A3(n14901), .ZN(n14832) );
  NAND2_X1 U18029 ( .A1(n14919), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14831) );
  OAI211_X1 U18030 ( .C1(n14919), .C2(n15239), .A(n14832), .B(n14831), .ZN(
        P2_U2858) );
  NAND2_X1 U18031 ( .A1(n14833), .A2(n14834), .ZN(n14836) );
  XNOR2_X1 U18032 ( .A(n14836), .B(n14835), .ZN(n14935) );
  OR2_X1 U18033 ( .A1(n14838), .A2(n14837), .ZN(n14839) );
  NAND2_X1 U18034 ( .A1(n14840), .A2(n14839), .ZN(n16201) );
  NOR2_X1 U18035 ( .A1(n16201), .A2(n14919), .ZN(n14841) );
  AOI21_X1 U18036 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n14919), .A(n14841), .ZN(
        n14842) );
  OAI21_X1 U18037 ( .B1(n14935), .B2(n14921), .A(n14842), .ZN(P2_U2859) );
  NAND2_X1 U18038 ( .A1(n14919), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14845) );
  OAI211_X1 U18039 ( .C1(n15260), .C2(n14919), .A(n14846), .B(n14845), .ZN(
        P2_U2860) );
  NOR2_X1 U18040 ( .A1(n14862), .A2(n14847), .ZN(n14848) );
  OR2_X1 U18041 ( .A1(n14849), .A2(n14848), .ZN(n16211) );
  AOI21_X1 U18042 ( .B1(n14850), .B2(n14852), .A(n14851), .ZN(n14942) );
  NAND2_X1 U18043 ( .A1(n14942), .A2(n14901), .ZN(n14854) );
  NAND2_X1 U18044 ( .A1(n14919), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n14853) );
  OAI211_X1 U18045 ( .C1(n16211), .C2(n14919), .A(n14854), .B(n14853), .ZN(
        P2_U2861) );
  OAI21_X1 U18046 ( .B1(n14856), .B2(n14858), .A(n14857), .ZN(n14958) );
  AND2_X1 U18047 ( .A1(n14860), .A2(n14859), .ZN(n14861) );
  NOR2_X1 U18048 ( .A1(n14862), .A2(n14861), .ZN(n16230) );
  NOR2_X1 U18049 ( .A1(n14906), .A2(n16222), .ZN(n14863) );
  AOI21_X1 U18050 ( .B1(n16230), .B2(n14906), .A(n14863), .ZN(n14864) );
  OAI21_X1 U18051 ( .B1(n14958), .B2(n14921), .A(n14864), .ZN(P2_U2862) );
  AOI21_X1 U18052 ( .B1(n14865), .B2(n14866), .A(n9854), .ZN(n14867) );
  XOR2_X1 U18053 ( .A(n14868), .B(n14867), .Z(n14964) );
  NOR2_X1 U18054 ( .A1(n15288), .A2(n14919), .ZN(n14869) );
  AOI21_X1 U18055 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n14919), .A(n14869), .ZN(
        n14870) );
  OAI21_X1 U18056 ( .B1(n14964), .B2(n14921), .A(n14870), .ZN(P2_U2863) );
  AOI21_X1 U18057 ( .B1(n14872), .B2(n14874), .A(n14873), .ZN(n14875) );
  INV_X1 U18058 ( .A(n14875), .ZN(n14972) );
  NAND2_X1 U18059 ( .A1(n14919), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n14877) );
  NAND2_X1 U18060 ( .A1(n15306), .A2(n14906), .ZN(n14876) );
  OAI211_X1 U18061 ( .C1(n14972), .C2(n14921), .A(n14877), .B(n14876), .ZN(
        P2_U2864) );
  AOI21_X1 U18062 ( .B1(n14879), .B2(n14878), .A(n11273), .ZN(n14880) );
  INV_X1 U18063 ( .A(n14880), .ZN(n14978) );
  MUX2_X1 U18064 ( .A(n14881), .B(n15319), .S(n14906), .Z(n14882) );
  OAI21_X1 U18065 ( .B1(n14978), .B2(n14921), .A(n14882), .ZN(P2_U2865) );
  OAI21_X1 U18066 ( .B1(n14883), .B2(n14884), .A(n14878), .ZN(n14984) );
  MUX2_X1 U18067 ( .A(n15331), .B(n10891), .S(n14919), .Z(n14885) );
  OAI21_X1 U18068 ( .B1(n14984), .B2(n14921), .A(n14885), .ZN(P2_U2866) );
  XNOR2_X1 U18069 ( .A(n14897), .B(n14886), .ZN(n18941) );
  AOI21_X1 U18070 ( .B1(n14889), .B2(n14888), .A(n14883), .ZN(n16235) );
  NAND2_X1 U18071 ( .A1(n16235), .A2(n14901), .ZN(n14891) );
  NAND2_X1 U18072 ( .A1(n14919), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n14890) );
  OAI211_X1 U18073 ( .C1(n18941), .C2(n14919), .A(n14891), .B(n14890), .ZN(
        P2_U2867) );
  OAI21_X1 U18074 ( .B1(n14893), .B2(n14894), .A(n14888), .ZN(n14996) );
  NAND2_X1 U18075 ( .A1(n14919), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n14899) );
  NAND2_X1 U18076 ( .A1(n14902), .A2(n14895), .ZN(n14896) );
  NAND2_X1 U18077 ( .A1(n14897), .A2(n14896), .ZN(n18954) );
  OR2_X1 U18078 ( .A1(n18954), .A2(n14919), .ZN(n14898) );
  OAI211_X1 U18079 ( .C1(n14996), .C2(n14921), .A(n14899), .B(n14898), .ZN(
        P2_U2868) );
  AOI21_X1 U18080 ( .B1(n14900), .B2(n13464), .A(n14893), .ZN(n16240) );
  NAND2_X1 U18081 ( .A1(n16240), .A2(n14901), .ZN(n14905) );
  OAI21_X1 U18082 ( .B1(n14909), .B2(n14903), .A(n14902), .ZN(n15141) );
  INV_X1 U18083 ( .A(n15141), .ZN(n18966) );
  NAND2_X1 U18084 ( .A1(n18966), .A2(n14906), .ZN(n14904) );
  OAI211_X1 U18085 ( .C1(n14906), .C2(n11040), .A(n14905), .B(n14904), .ZN(
        P2_U2869) );
  NOR2_X1 U18086 ( .A1(n9912), .A2(n14907), .ZN(n14908) );
  OR2_X1 U18087 ( .A1(n14909), .A2(n14908), .ZN(n18976) );
  NOR2_X1 U18088 ( .A1(n18976), .A2(n14919), .ZN(n14910) );
  AOI21_X1 U18089 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n14919), .A(n14910), .ZN(
        n14911) );
  OAI21_X1 U18090 ( .B1(n14912), .B2(n14921), .A(n14911), .ZN(P2_U2870) );
  AND2_X1 U18091 ( .A1(n14914), .A2(n14913), .ZN(n14915) );
  OR2_X1 U18092 ( .A1(n13465), .A2(n14915), .ZN(n19130) );
  AND2_X1 U18093 ( .A1(n14917), .A2(n14916), .ZN(n14918) );
  OR2_X1 U18094 ( .A1(n14918), .A2(n9912), .ZN(n18990) );
  MUX2_X1 U18095 ( .A(n18990), .B(n10888), .S(n14919), .Z(n14920) );
  OAI21_X1 U18096 ( .B1(n19130), .B2(n14921), .A(n14920), .ZN(P2_U2871) );
  NAND3_X1 U18097 ( .A1(n14828), .A2(n14922), .A3(n19137), .ZN(n14928) );
  INV_X1 U18098 ( .A(n15236), .ZN(n14925) );
  OAI22_X1 U18099 ( .A1(n14988), .A2(n19142), .B1(n19160), .B2(n14923), .ZN(
        n14924) );
  AOI21_X1 U18100 ( .B1(n14925), .B2(n19177), .A(n14924), .ZN(n14927) );
  AOI22_X1 U18101 ( .A1(n19128), .A2(BUF2_REG_29__SCAN_IN), .B1(n19129), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n14926) );
  NAND3_X1 U18102 ( .A1(n14928), .A2(n14927), .A3(n14926), .ZN(P2_U2890) );
  NAND2_X1 U18103 ( .A1(n12446), .A2(n14929), .ZN(n14930) );
  INV_X1 U18104 ( .A(n19145), .ZN(n14931) );
  OAI22_X1 U18105 ( .A1(n14988), .A2(n14931), .B1(n19160), .B2(n12723), .ZN(
        n14932) );
  AOI21_X1 U18106 ( .B1(n19177), .B2(n16204), .A(n14932), .ZN(n14934) );
  AOI22_X1 U18107 ( .A1(n19128), .A2(BUF2_REG_28__SCAN_IN), .B1(n19129), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n14933) );
  OAI211_X1 U18108 ( .C1(n14935), .C2(n19181), .A(n14934), .B(n14933), .ZN(
        P2_U2891) );
  INV_X1 U18109 ( .A(n14936), .ZN(n14941) );
  OAI22_X1 U18110 ( .A1(n14988), .A2(n19148), .B1(n19160), .B2(n14937), .ZN(
        n14938) );
  AOI21_X1 U18111 ( .B1(n19177), .B2(n15258), .A(n14938), .ZN(n14940) );
  AOI22_X1 U18112 ( .A1(n19128), .A2(BUF2_REG_27__SCAN_IN), .B1(n19129), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n14939) );
  OAI211_X1 U18113 ( .C1(n14941), .C2(n19181), .A(n14940), .B(n14939), .ZN(
        P2_U2892) );
  NAND2_X1 U18114 ( .A1(n14942), .A2(n19137), .ZN(n14949) );
  INV_X1 U18115 ( .A(n14988), .ZN(n19127) );
  AOI22_X1 U18116 ( .A1(n19127), .A2(n19150), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n19176), .ZN(n14948) );
  AOI22_X1 U18117 ( .A1(n19128), .A2(BUF2_REG_26__SCAN_IN), .B1(n19129), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n14947) );
  AND2_X1 U18118 ( .A1(n14952), .A2(n14943), .ZN(n14944) );
  NOR2_X1 U18119 ( .A1(n14945), .A2(n14944), .ZN(n16209) );
  NAND2_X1 U18120 ( .A1(n19177), .A2(n16209), .ZN(n14946) );
  NAND4_X1 U18121 ( .A1(n14949), .A2(n14948), .A3(n14947), .A4(n14946), .ZN(
        P2_U2893) );
  NAND2_X1 U18122 ( .A1(n9874), .A2(n14950), .ZN(n14951) );
  NAND2_X1 U18123 ( .A1(n14952), .A2(n14951), .ZN(n16232) );
  INV_X1 U18124 ( .A(n16232), .ZN(n14955) );
  OAI22_X1 U18125 ( .A1(n14988), .A2(n19153), .B1(n19160), .B2(n14953), .ZN(
        n14954) );
  AOI21_X1 U18126 ( .B1(n19177), .B2(n14955), .A(n14954), .ZN(n14957) );
  AOI22_X1 U18127 ( .A1(n19128), .A2(BUF2_REG_25__SCAN_IN), .B1(n19129), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n14956) );
  OAI211_X1 U18128 ( .C1(n14958), .C2(n19181), .A(n14957), .B(n14956), .ZN(
        P2_U2894) );
  INV_X1 U18129 ( .A(n15292), .ZN(n14961) );
  OAI22_X1 U18130 ( .A1(n14988), .A2(n19155), .B1(n19160), .B2(n14959), .ZN(
        n14960) );
  AOI21_X1 U18131 ( .B1(n19177), .B2(n14961), .A(n14960), .ZN(n14963) );
  AOI22_X1 U18132 ( .A1(n19128), .A2(BUF2_REG_24__SCAN_IN), .B1(n19129), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n14962) );
  OAI211_X1 U18133 ( .C1(n14964), .C2(n19181), .A(n14963), .B(n14962), .ZN(
        P2_U2895) );
  INV_X1 U18134 ( .A(n15304), .ZN(n14970) );
  OAI22_X1 U18135 ( .A1(n14988), .A2(n19157), .B1(n19160), .B2(n14965), .ZN(
        n14969) );
  INV_X1 U18136 ( .A(n19128), .ZN(n14991) );
  INV_X1 U18137 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n14967) );
  INV_X1 U18138 ( .A(n19129), .ZN(n14989) );
  INV_X1 U18139 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n14966) );
  OAI22_X1 U18140 ( .A1(n14991), .A2(n14967), .B1(n14989), .B2(n14966), .ZN(
        n14968) );
  AOI211_X1 U18141 ( .C1(n19177), .C2(n14970), .A(n14969), .B(n14968), .ZN(
        n14971) );
  OAI21_X1 U18142 ( .B1(n14972), .B2(n19181), .A(n14971), .ZN(P2_U2896) );
  OAI22_X1 U18143 ( .A1(n14988), .A2(n19159), .B1(n19160), .B2(n14973), .ZN(
        n14976) );
  INV_X1 U18144 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n14974) );
  OAI22_X1 U18145 ( .A1(n14991), .A2(n14974), .B1(n14989), .B2(n20280), .ZN(
        n14975) );
  AOI211_X1 U18146 ( .C1(n19177), .C2(n15315), .A(n14976), .B(n14975), .ZN(
        n14977) );
  OAI21_X1 U18147 ( .B1(n14978), .B2(n19181), .A(n14977), .ZN(P2_U2897) );
  INV_X1 U18148 ( .A(n19163), .ZN(n19268) );
  NAND2_X1 U18149 ( .A1(n19177), .A2(n15328), .ZN(n14980) );
  NAND2_X1 U18150 ( .A1(n19176), .A2(P2_EAX_REG_21__SCAN_IN), .ZN(n14979) );
  OAI211_X1 U18151 ( .C1(n19268), .C2(n14988), .A(n14980), .B(n14979), .ZN(
        n14981) );
  INV_X1 U18152 ( .A(n14981), .ZN(n14983) );
  AOI22_X1 U18153 ( .A1(n19128), .A2(BUF2_REG_21__SCAN_IN), .B1(n19129), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n14982) );
  OAI211_X1 U18154 ( .C1(n14984), .C2(n19181), .A(n14983), .B(n14982), .ZN(
        P2_U2898) );
  NOR2_X1 U18155 ( .A1(n14985), .A2(n15360), .ZN(n14986) );
  OR2_X1 U18156 ( .A1(n15341), .A2(n14986), .ZN(n18953) );
  INV_X1 U18157 ( .A(n18953), .ZN(n14994) );
  OAI22_X1 U18158 ( .A1(n14988), .A2(n19257), .B1(n19160), .B2(n14987), .ZN(
        n14993) );
  INV_X1 U18159 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n14990) );
  OAI22_X1 U18160 ( .A1(n14991), .A2(n14990), .B1(n14989), .B2(n20258), .ZN(
        n14992) );
  AOI211_X1 U18161 ( .C1(n19177), .C2(n14994), .A(n14993), .B(n14992), .ZN(
        n14995) );
  OAI21_X1 U18162 ( .B1(n14996), .B2(n19181), .A(n14995), .ZN(P2_U2900) );
  NAND2_X1 U18163 ( .A1(n14997), .A2(n15011), .ZN(n15002) );
  INV_X1 U18164 ( .A(n14998), .ZN(n14999) );
  NOR2_X1 U18165 ( .A1(n15000), .A2(n14999), .ZN(n15001) );
  XNOR2_X1 U18166 ( .A(n15002), .B(n15001), .ZN(n15227) );
  XOR2_X1 U18167 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n15014), .Z(
        n15225) );
  INV_X1 U18168 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15004) );
  OR2_X1 U18169 ( .A1(n19040), .A2(n15003), .ZN(n15216) );
  OAI21_X1 U18170 ( .B1(n19234), .B2(n15004), .A(n15216), .ZN(n15005) );
  AOI21_X1 U18171 ( .B1(n19222), .B2(n15006), .A(n15005), .ZN(n15007) );
  OAI21_X1 U18172 ( .B1(n15223), .B2(n13154), .A(n15007), .ZN(n15008) );
  AOI21_X1 U18173 ( .B1(n15225), .B2(n16283), .A(n15008), .ZN(n15009) );
  OAI21_X1 U18174 ( .B1(n15227), .B2(n19227), .A(n15009), .ZN(P2_U2984) );
  NAND2_X1 U18175 ( .A1(n15011), .A2(n15010), .ZN(n15013) );
  XOR2_X1 U18176 ( .A(n15013), .B(n15012), .Z(n15244) );
  AOI21_X1 U18177 ( .B1(n15234), .B2(n9830), .A(n15014), .ZN(n15242) );
  OAI21_X1 U18178 ( .B1(n19234), .B2(n15015), .A(n10364), .ZN(n15016) );
  AOI21_X1 U18179 ( .B1(n19222), .B2(n15017), .A(n15016), .ZN(n15018) );
  OAI21_X1 U18180 ( .B1(n15239), .B2(n13154), .A(n15018), .ZN(n15019) );
  AOI21_X1 U18181 ( .B1(n15242), .B2(n16283), .A(n15019), .ZN(n15020) );
  OAI21_X1 U18182 ( .B1(n15244), .B2(n19227), .A(n15020), .ZN(P2_U2985) );
  NAND2_X1 U18183 ( .A1(n15022), .A2(n9892), .ZN(n15024) );
  XNOR2_X1 U18184 ( .A(n15024), .B(n15023), .ZN(n15036) );
  INV_X1 U18185 ( .A(n15023), .ZN(n15025) );
  AOI22_X1 U18186 ( .A1(n15036), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n15025), .B2(n15024), .ZN(n15028) );
  XNOR2_X1 U18187 ( .A(n15026), .B(n10010), .ZN(n15027) );
  XNOR2_X1 U18188 ( .A(n15028), .B(n15027), .ZN(n15252) );
  INV_X1 U18189 ( .A(n9830), .ZN(n15030) );
  AOI21_X1 U18190 ( .B1(n10010), .B2(n15029), .A(n15030), .ZN(n15250) );
  INV_X1 U18191 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n16197) );
  NOR2_X1 U18192 ( .A1(n19083), .A2(n16197), .ZN(n15245) );
  NOR2_X1 U18193 ( .A1(n15211), .A2(n15031), .ZN(n15032) );
  AOI211_X1 U18194 ( .C1(n15162), .C2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15245), .B(n15032), .ZN(n15033) );
  OAI21_X1 U18195 ( .B1(n16201), .B2(n13154), .A(n15033), .ZN(n15034) );
  AOI21_X1 U18196 ( .B1(n15250), .B2(n16283), .A(n15034), .ZN(n15035) );
  OAI21_X1 U18197 ( .B1(n15252), .B2(n19227), .A(n15035), .ZN(P2_U2986) );
  XNOR2_X1 U18198 ( .A(n15036), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15265) );
  INV_X1 U18199 ( .A(n15228), .ZN(n15230) );
  NAND2_X1 U18200 ( .A1(n9815), .A2(n15230), .ZN(n15045) );
  INV_X1 U18201 ( .A(n15029), .ZN(n15038) );
  AOI21_X1 U18202 ( .B1(n15255), .B2(n15045), .A(n15038), .ZN(n15263) );
  OR2_X1 U18203 ( .A1(n19040), .A2(n19907), .ZN(n15256) );
  OAI21_X1 U18204 ( .B1(n19234), .B2(n15039), .A(n15256), .ZN(n15040) );
  AOI21_X1 U18205 ( .B1(n19222), .B2(n15041), .A(n15040), .ZN(n15042) );
  OAI21_X1 U18206 ( .B1(n15260), .B2(n13154), .A(n15042), .ZN(n15043) );
  AOI21_X1 U18207 ( .B1(n15263), .B2(n16283), .A(n15043), .ZN(n15044) );
  OAI21_X1 U18208 ( .B1(n15265), .B2(n19227), .A(n15044), .ZN(P2_U2987) );
  OAI21_X1 U18209 ( .B1(n15059), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15045), .ZN(n15277) );
  OAI21_X1 U18210 ( .B1(n15046), .B2(n15055), .A(n15056), .ZN(n15048) );
  XNOR2_X1 U18211 ( .A(n15048), .B(n15047), .ZN(n15275) );
  NOR2_X1 U18212 ( .A1(n19083), .A2(n15049), .ZN(n15267) );
  NOR2_X1 U18213 ( .A1(n15211), .A2(n15050), .ZN(n15051) );
  AOI211_X1 U18214 ( .C1(n15162), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15267), .B(n15051), .ZN(n15052) );
  OAI21_X1 U18215 ( .B1(n16211), .B2(n13154), .A(n15052), .ZN(n15053) );
  AOI21_X1 U18216 ( .B1(n15275), .B2(n16282), .A(n15053), .ZN(n15054) );
  OAI21_X1 U18217 ( .B1(n15277), .B2(n19225), .A(n15054), .ZN(P2_U2988) );
  INV_X1 U18218 ( .A(n15055), .ZN(n15057) );
  NAND2_X1 U18219 ( .A1(n15057), .A2(n15056), .ZN(n15058) );
  XNOR2_X1 U18220 ( .A(n15046), .B(n15058), .ZN(n15287) );
  AOI21_X1 U18221 ( .B1(n15060), .B2(n15066), .A(n15059), .ZN(n15278) );
  NAND2_X1 U18222 ( .A1(n15278), .A2(n16283), .ZN(n15065) );
  INV_X1 U18223 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19903) );
  NOR2_X1 U18224 ( .A1(n19083), .A2(n19903), .ZN(n15280) );
  AOI21_X1 U18225 ( .B1(n15162), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15280), .ZN(n15061) );
  OAI21_X1 U18226 ( .B1(n15211), .B2(n15062), .A(n15061), .ZN(n15063) );
  AOI21_X1 U18227 ( .B1(n16230), .B2(n19231), .A(n15063), .ZN(n15064) );
  OAI211_X1 U18228 ( .C1(n19227), .C2(n15287), .A(n15065), .B(n15064), .ZN(
        P2_U2989) );
  OAI21_X1 U18229 ( .B1(n9815), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15066), .ZN(n15301) );
  XNOR2_X1 U18230 ( .A(n15068), .B(n15289), .ZN(n15069) );
  XNOR2_X1 U18231 ( .A(n15067), .B(n15069), .ZN(n15299) );
  NAND2_X1 U18232 ( .A1(n19223), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n15291) );
  OAI21_X1 U18233 ( .B1(n19234), .B2(n15070), .A(n15291), .ZN(n15071) );
  AOI21_X1 U18234 ( .B1(n19222), .B2(n15072), .A(n15071), .ZN(n15073) );
  OAI21_X1 U18235 ( .B1(n15288), .B2(n13154), .A(n15073), .ZN(n15074) );
  AOI21_X1 U18236 ( .B1(n15299), .B2(n16282), .A(n15074), .ZN(n15075) );
  OAI21_X1 U18237 ( .B1(n15301), .B2(n19225), .A(n15075), .ZN(P2_U2990) );
  CLKBUF_X1 U18238 ( .A(n15076), .Z(n15077) );
  INV_X1 U18239 ( .A(n9815), .ZN(n15078) );
  OAI21_X1 U18240 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15077), .A(
        n15078), .ZN(n15312) );
  NAND2_X1 U18241 ( .A1(n19222), .A2(n15079), .ZN(n15080) );
  NAND2_X1 U18242 ( .A1(n19223), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n15302) );
  OAI211_X1 U18243 ( .C1(n19234), .C2(n10164), .A(n15080), .B(n15302), .ZN(
        n15081) );
  AOI21_X1 U18244 ( .B1(n15306), .B2(n19231), .A(n15081), .ZN(n15085) );
  XOR2_X1 U18245 ( .A(n15083), .B(n15082), .Z(n15310) );
  NAND2_X1 U18246 ( .A1(n15310), .A2(n16282), .ZN(n15084) );
  OAI211_X1 U18247 ( .C1(n15312), .C2(n19225), .A(n15085), .B(n15084), .ZN(
        P2_U2991) );
  OAI21_X1 U18249 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n15087), .A(
        n10042), .ZN(n15324) );
  NAND2_X1 U18250 ( .A1(n15089), .A2(n15088), .ZN(n15090) );
  XNOR2_X1 U18251 ( .A(n15091), .B(n15090), .ZN(n15322) );
  NOR2_X1 U18252 ( .A1(n19040), .A2(n19897), .ZN(n15314) );
  NOR2_X1 U18253 ( .A1(n15211), .A2(n15092), .ZN(n15093) );
  AOI211_X1 U18254 ( .C1(n15162), .C2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15314), .B(n15093), .ZN(n15094) );
  OAI21_X1 U18255 ( .B1(n15319), .B2(n13154), .A(n15094), .ZN(n15095) );
  AOI21_X1 U18256 ( .B1(n15322), .B2(n16282), .A(n15095), .ZN(n15096) );
  OAI21_X1 U18257 ( .B1(n15324), .B2(n19225), .A(n15096), .ZN(P2_U2992) );
  INV_X1 U18258 ( .A(n15434), .ZN(n15097) );
  INV_X1 U18259 ( .A(n15098), .ZN(n15160) );
  NAND2_X1 U18260 ( .A1(n15103), .A2(n15102), .ZN(n15117) );
  NAND2_X1 U18261 ( .A1(n15116), .A2(n15103), .ZN(n15107) );
  NAND2_X1 U18262 ( .A1(n15105), .A2(n15104), .ZN(n15106) );
  XNOR2_X1 U18263 ( .A(n15107), .B(n15106), .ZN(n15335) );
  AOI21_X1 U18264 ( .B1(n15109), .B2(n15108), .A(n15087), .ZN(n15333) );
  NOR2_X1 U18265 ( .A1(n19040), .A2(n19895), .ZN(n15327) );
  NOR2_X1 U18266 ( .A1(n19234), .A2(n15110), .ZN(n15111) );
  AOI211_X1 U18267 ( .C1(n19222), .C2(n15112), .A(n15327), .B(n15111), .ZN(
        n15113) );
  OAI21_X1 U18268 ( .B1(n15331), .B2(n13154), .A(n15113), .ZN(n15114) );
  AOI21_X1 U18269 ( .B1(n15333), .B2(n16283), .A(n15114), .ZN(n15115) );
  OAI21_X1 U18270 ( .B1(n15335), .B2(n19227), .A(n15115), .ZN(P2_U2993) );
  INV_X1 U18271 ( .A(n15108), .ZN(n15119) );
  AOI21_X1 U18272 ( .B1(n15338), .B2(n9877), .A(n15119), .ZN(n15347) );
  NOR2_X1 U18273 ( .A1(n19040), .A2(n19893), .ZN(n15343) );
  NOR2_X1 U18274 ( .A1(n15211), .A2(n15120), .ZN(n15121) );
  AOI211_X1 U18275 ( .C1(n15162), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15343), .B(n15121), .ZN(n15122) );
  OAI21_X1 U18276 ( .B1(n18941), .B2(n13154), .A(n15122), .ZN(n15123) );
  AOI21_X1 U18277 ( .B1(n15347), .B2(n16283), .A(n15123), .ZN(n15124) );
  INV_X1 U18278 ( .A(n15125), .ZN(n15126) );
  OAI21_X1 U18279 ( .B1(n15126), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n9877), .ZN(n15359) );
  INV_X1 U18280 ( .A(n15137), .ZN(n15127) );
  NAND2_X1 U18281 ( .A1(n15129), .A2(n15128), .ZN(n15130) );
  XNOR2_X1 U18282 ( .A(n15131), .B(n15130), .ZN(n15350) );
  NAND2_X1 U18283 ( .A1(n15350), .A2(n16282), .ZN(n15135) );
  NAND2_X1 U18284 ( .A1(n19223), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15352) );
  OAI21_X1 U18285 ( .B1(n19234), .B2(n18959), .A(n15352), .ZN(n15133) );
  NOR2_X1 U18286 ( .A1(n18954), .A2(n13154), .ZN(n15132) );
  AOI211_X1 U18287 ( .C1(n19222), .C2(n18952), .A(n15133), .B(n15132), .ZN(
        n15134) );
  OAI211_X1 U18288 ( .C1(n19225), .C2(n15359), .A(n15135), .B(n15134), .ZN(
        P2_U2995) );
  NAND2_X1 U18289 ( .A1(n15137), .A2(n15136), .ZN(n15138) );
  XNOR2_X1 U18290 ( .A(n15139), .B(n15138), .ZN(n15372) );
  INV_X1 U18291 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19889) );
  OAI22_X1 U18292 ( .A1(n19889), .A2(n19040), .B1(n15211), .B2(n15140), .ZN(
        n15143) );
  NOR2_X1 U18293 ( .A1(n15141), .A2(n13154), .ZN(n15142) );
  AOI211_X1 U18294 ( .C1(n15162), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15143), .B(n15142), .ZN(n15147) );
  INV_X1 U18295 ( .A(n15144), .ZN(n15145) );
  NAND2_X1 U18296 ( .A1(n15145), .A2(n15366), .ZN(n15369) );
  NAND3_X1 U18297 ( .A1(n15369), .A2(n16283), .A3(n15125), .ZN(n15146) );
  OAI211_X1 U18298 ( .C1(n15372), .C2(n19227), .A(n15147), .B(n15146), .ZN(
        P2_U2996) );
  NAND2_X1 U18299 ( .A1(n15149), .A2(n15148), .ZN(n15150) );
  XNOR2_X1 U18300 ( .A(n15151), .B(n15150), .ZN(n15373) );
  OAI21_X1 U18301 ( .B1(n15152), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n16283), .ZN(n15153) );
  NOR2_X1 U18302 ( .A1(n15153), .A2(n15144), .ZN(n15157) );
  OAI22_X1 U18303 ( .A1(n18982), .A2(n19234), .B1(n15211), .B2(n18975), .ZN(
        n15154) );
  NOR2_X1 U18304 ( .A1(n19040), .A2(n19887), .ZN(n15384) );
  NOR2_X1 U18305 ( .A1(n15154), .A2(n15384), .ZN(n15155) );
  OAI21_X1 U18306 ( .B1(n18976), .B2(n13154), .A(n15155), .ZN(n15156) );
  AOI211_X1 U18307 ( .C1(n15373), .C2(n16282), .A(n15157), .B(n15156), .ZN(
        n15158) );
  INV_X1 U18308 ( .A(n15158), .ZN(P2_U2997) );
  OAI21_X1 U18309 ( .B1(n15161), .B2(n15160), .A(n15159), .ZN(n15392) );
  INV_X1 U18310 ( .A(n18990), .ZN(n15397) );
  NOR2_X1 U18311 ( .A1(n19040), .A2(n19885), .ZN(n15396) );
  AOI21_X1 U18312 ( .B1(n15162), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n15396), .ZN(n15163) );
  OAI21_X1 U18313 ( .B1(n15211), .B2(n15164), .A(n15163), .ZN(n15167) );
  AOI211_X1 U18314 ( .C1(n15403), .C2(n15165), .A(n19225), .B(n15152), .ZN(
        n15166) );
  AOI211_X1 U18315 ( .C1(n19231), .C2(n15397), .A(n15167), .B(n15166), .ZN(
        n15168) );
  OAI21_X1 U18316 ( .B1(n19227), .B2(n15392), .A(n15168), .ZN(P2_U2998) );
  INV_X1 U18317 ( .A(n15170), .ZN(n15171) );
  NOR2_X1 U18318 ( .A1(n15174), .A2(n15171), .ZN(n15172) );
  OAI22_X1 U18319 ( .A1(n10245), .A2(n15174), .B1(n15173), .B2(n15172), .ZN(
        n15432) );
  NOR2_X1 U18320 ( .A1(n15477), .A2(n15441), .ZN(n15459) );
  AOI21_X1 U18321 ( .B1(n15459), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15177) );
  NOR2_X1 U18322 ( .A1(n15177), .A2(n15176), .ZN(n15430) );
  INV_X1 U18323 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n19881) );
  OAI22_X1 U18324 ( .A1(n19881), .A2(n19040), .B1(n15211), .B2(n15178), .ZN(
        n15180) );
  OAI22_X1 U18325 ( .A1(n15423), .A2(n13154), .B1(n10149), .B2(n19234), .ZN(
        n15179) );
  AOI211_X1 U18326 ( .C1(n15430), .C2(n16283), .A(n15180), .B(n15179), .ZN(
        n15181) );
  OAI21_X1 U18327 ( .B1(n15432), .B2(n19227), .A(n15181), .ZN(P2_U3000) );
  NAND2_X1 U18328 ( .A1(n15183), .A2(n15182), .ZN(n15184) );
  XNOR2_X1 U18329 ( .A(n15185), .B(n15184), .ZN(n15464) );
  INV_X1 U18330 ( .A(n15477), .ZN(n15186) );
  NOR2_X1 U18331 ( .A1(n15186), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15460) );
  NOR3_X1 U18332 ( .A1(n15460), .A2(n15459), .A3(n19225), .ZN(n15190) );
  INV_X1 U18333 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19877) );
  OAI22_X1 U18334 ( .A1(n19877), .A2(n19040), .B1(n15211), .B2(n15187), .ZN(
        n15189) );
  OAI22_X1 U18335 ( .A1(n15454), .A2(n13154), .B1(n10151), .B2(n19234), .ZN(
        n15188) );
  NOR3_X1 U18336 ( .A1(n15190), .A2(n15189), .A3(n15188), .ZN(n15191) );
  OAI21_X1 U18337 ( .B1(n19227), .B2(n15464), .A(n15191), .ZN(P2_U3002) );
  NAND2_X1 U18338 ( .A1(n15192), .A2(n15505), .ZN(n15197) );
  INV_X1 U18339 ( .A(n15193), .ZN(n15194) );
  NOR2_X1 U18340 ( .A1(n15195), .A2(n15194), .ZN(n15196) );
  XNOR2_X1 U18341 ( .A(n15197), .B(n15196), .ZN(n15496) );
  AOI21_X1 U18342 ( .B1(n15488), .B2(n15198), .A(n15199), .ZN(n15493) );
  INV_X1 U18343 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n19873) );
  OAI22_X1 U18344 ( .A1(n19873), .A2(n19040), .B1(n15211), .B2(n19060), .ZN(
        n15203) );
  INV_X1 U18345 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n15200) );
  OAI22_X1 U18346 ( .A1(n13154), .A2(n15201), .B1(n15200), .B2(n19234), .ZN(
        n15202) );
  AOI211_X1 U18347 ( .C1(n15493), .C2(n16283), .A(n15203), .B(n15202), .ZN(
        n15204) );
  OAI21_X1 U18348 ( .B1(n15496), .B2(n19227), .A(n15204), .ZN(P2_U3004) );
  XNOR2_X1 U18349 ( .A(n15206), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15207) );
  XNOR2_X1 U18350 ( .A(n9833), .B(n15207), .ZN(n15520) );
  INV_X1 U18351 ( .A(n16275), .ZN(n15209) );
  NAND2_X1 U18352 ( .A1(n15209), .A2(n16276), .ZN(n15210) );
  XNOR2_X1 U18353 ( .A(n15208), .B(n15210), .ZN(n15518) );
  OAI22_X1 U18354 ( .A1(n19867), .A2(n19040), .B1(n15211), .B2(n19079), .ZN(
        n15213) );
  OAI22_X1 U18355 ( .A1(n13154), .A2(n19086), .B1(n10168), .B2(n19234), .ZN(
        n15212) );
  AOI211_X1 U18356 ( .C1(n15518), .C2(n16282), .A(n15213), .B(n15212), .ZN(
        n15214) );
  OAI21_X1 U18357 ( .B1(n19225), .B2(n15520), .A(n15214), .ZN(P2_U3007) );
  INV_X1 U18358 ( .A(n15215), .ZN(n15217) );
  OAI21_X1 U18359 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15217), .A(
        n15216), .ZN(n15220) );
  NOR2_X1 U18360 ( .A1(n15218), .A2(n9832), .ZN(n15219) );
  AOI211_X1 U18361 ( .C1(n16299), .C2(n15221), .A(n15220), .B(n15219), .ZN(
        n15222) );
  OAI21_X1 U18362 ( .B1(n15223), .B2(n16314), .A(n15222), .ZN(n15224) );
  AOI21_X1 U18363 ( .B1(n15225), .B2(n16301), .A(n15224), .ZN(n15226) );
  OAI21_X1 U18364 ( .B1(n15227), .B2(n15495), .A(n15226), .ZN(P2_U3016) );
  INV_X1 U18365 ( .A(n15297), .ZN(n15269) );
  NOR2_X1 U18366 ( .A1(n15228), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15229) );
  NAND2_X1 U18367 ( .A1(n15269), .A2(n15229), .ZN(n15254) );
  NAND2_X1 U18368 ( .A1(n15290), .A2(n15230), .ZN(n15231) );
  NAND2_X1 U18369 ( .A1(n15231), .A2(n15316), .ZN(n15232) );
  NAND2_X1 U18370 ( .A1(n15233), .A2(n10010), .ZN(n15247) );
  AOI21_X1 U18371 ( .B1(n15253), .B2(n15247), .A(n15234), .ZN(n15241) );
  OAI211_X1 U18372 ( .C1(n16313), .C2(n15236), .A(n10364), .B(n10357), .ZN(
        n15237) );
  INV_X1 U18373 ( .A(n15237), .ZN(n15238) );
  OAI21_X1 U18374 ( .B1(n15239), .B2(n16314), .A(n15238), .ZN(n15240) );
  OAI21_X1 U18375 ( .B1(n15244), .B2(n15495), .A(n15243), .ZN(P2_U3017) );
  NOR2_X1 U18376 ( .A1(n15253), .A2(n10010), .ZN(n15249) );
  AOI21_X1 U18377 ( .B1(n16299), .B2(n16204), .A(n15245), .ZN(n15246) );
  OAI211_X1 U18378 ( .C1(n16201), .C2(n16314), .A(n15247), .B(n15246), .ZN(
        n15248) );
  AOI211_X1 U18379 ( .C1(n15250), .C2(n16301), .A(n15249), .B(n15248), .ZN(
        n15251) );
  OAI21_X1 U18380 ( .B1(n15252), .B2(n15495), .A(n15251), .ZN(P2_U3018) );
  AOI21_X1 U18381 ( .B1(n15255), .B2(n15254), .A(n15253), .ZN(n15262) );
  INV_X1 U18382 ( .A(n15256), .ZN(n15257) );
  AOI21_X1 U18383 ( .B1(n16299), .B2(n15258), .A(n15257), .ZN(n15259) );
  OAI21_X1 U18384 ( .B1(n15260), .B2(n16314), .A(n15259), .ZN(n15261) );
  AOI211_X1 U18385 ( .C1(n15263), .C2(n16301), .A(n15262), .B(n15261), .ZN(
        n15264) );
  OAI21_X1 U18386 ( .B1(n15265), .B2(n15495), .A(n15264), .ZN(P2_U3019) );
  NAND2_X1 U18387 ( .A1(n15290), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15279) );
  NOR3_X1 U18388 ( .A1(n15297), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n15289), .ZN(n15283) );
  AOI21_X1 U18389 ( .B1(n15316), .B2(n15279), .A(n15283), .ZN(n15273) );
  NOR2_X1 U18390 ( .A1(n16211), .A2(n16314), .ZN(n15266) );
  AOI211_X1 U18391 ( .C1(n16299), .C2(n16209), .A(n15267), .B(n15266), .ZN(
        n15271) );
  NAND3_X1 U18392 ( .A1(n15269), .A2(n15268), .A3(n15272), .ZN(n15270) );
  OAI211_X1 U18393 ( .C1(n15273), .C2(n15272), .A(n15271), .B(n15270), .ZN(
        n15274) );
  AOI21_X1 U18394 ( .B1(n15275), .B2(n16322), .A(n15274), .ZN(n15276) );
  OAI21_X1 U18395 ( .B1(n15277), .B2(n16326), .A(n15276), .ZN(P2_U3020) );
  NAND2_X1 U18396 ( .A1(n15278), .A2(n16301), .ZN(n15286) );
  NAND3_X1 U18397 ( .A1(n15279), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n15316), .ZN(n15282) );
  INV_X1 U18398 ( .A(n15280), .ZN(n15281) );
  OAI211_X1 U18399 ( .C1(n16313), .C2(n16232), .A(n15282), .B(n15281), .ZN(
        n15284) );
  AOI211_X1 U18400 ( .C1(n16304), .C2(n16230), .A(n15284), .B(n15283), .ZN(
        n15285) );
  OAI211_X1 U18401 ( .C1(n15287), .C2(n15495), .A(n15286), .B(n15285), .ZN(
        P2_U3021) );
  INV_X1 U18402 ( .A(n15288), .ZN(n15295) );
  NOR3_X1 U18403 ( .A1(n15290), .A2(n15473), .A3(n15289), .ZN(n15294) );
  OAI21_X1 U18404 ( .B1(n16313), .B2(n15292), .A(n15291), .ZN(n15293) );
  AOI211_X1 U18405 ( .C1(n15295), .C2(n16304), .A(n15294), .B(n15293), .ZN(
        n15296) );
  OAI21_X1 U18406 ( .B1(n15297), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15296), .ZN(n15298) );
  AOI21_X1 U18407 ( .B1(n15299), .B2(n16322), .A(n15298), .ZN(n15300) );
  OAI21_X1 U18408 ( .B1(n15301), .B2(n16326), .A(n15300), .ZN(P2_U3022) );
  XNOR2_X1 U18409 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15308) );
  NAND3_X1 U18410 ( .A1(n15325), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n15316), .ZN(n15303) );
  OAI211_X1 U18411 ( .C1(n16313), .C2(n15304), .A(n15303), .B(n15302), .ZN(
        n15305) );
  AOI21_X1 U18412 ( .B1(n15306), .B2(n16304), .A(n15305), .ZN(n15307) );
  OAI21_X1 U18413 ( .B1(n15313), .B2(n15308), .A(n15307), .ZN(n15309) );
  AOI21_X1 U18414 ( .B1(n15310), .B2(n16322), .A(n15309), .ZN(n15311) );
  OAI21_X1 U18415 ( .B1(n15312), .B2(n16326), .A(n15311), .ZN(P2_U3023) );
  NOR2_X1 U18416 ( .A1(n15313), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15321) );
  AOI21_X1 U18417 ( .B1(n16299), .B2(n15315), .A(n15314), .ZN(n15318) );
  NAND3_X1 U18418 ( .A1(n15325), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n15316), .ZN(n15317) );
  OAI211_X1 U18419 ( .C1(n15319), .C2(n16314), .A(n15318), .B(n15317), .ZN(
        n15320) );
  AOI211_X1 U18420 ( .C1(n15322), .C2(n16322), .A(n15321), .B(n15320), .ZN(
        n15323) );
  OAI21_X1 U18421 ( .B1(n15324), .B2(n16326), .A(n15323), .ZN(P2_U3024) );
  OAI21_X1 U18422 ( .B1(n15326), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15325), .ZN(n15330) );
  AOI21_X1 U18423 ( .B1(n16299), .B2(n15328), .A(n15327), .ZN(n15329) );
  OAI211_X1 U18424 ( .C1(n16314), .C2(n15331), .A(n15330), .B(n15329), .ZN(
        n15332) );
  AOI21_X1 U18425 ( .B1(n15333), .B2(n16301), .A(n15332), .ZN(n15334) );
  OAI21_X1 U18426 ( .B1(n15335), .B2(n15495), .A(n15334), .ZN(P2_U3025) );
  AOI211_X1 U18427 ( .C1(n15338), .C2(n15337), .A(n15336), .B(n15354), .ZN(
        n15346) );
  OAI21_X1 U18428 ( .B1(n15341), .B2(n15340), .A(n15339), .ZN(n16234) );
  NOR2_X1 U18429 ( .A1(n16313), .A2(n16234), .ZN(n15342) );
  AOI211_X1 U18430 ( .C1(n15362), .C2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15343), .B(n15342), .ZN(n15344) );
  OAI21_X1 U18431 ( .B1(n18941), .B2(n16314), .A(n15344), .ZN(n15345) );
  AOI211_X1 U18432 ( .C1(n15347), .C2(n16301), .A(n15346), .B(n15345), .ZN(
        n15348) );
  OAI21_X1 U18433 ( .B1(n15349), .B2(n15495), .A(n15348), .ZN(P2_U3026) );
  NAND2_X1 U18434 ( .A1(n15350), .A2(n16322), .ZN(n15358) );
  INV_X1 U18435 ( .A(n18954), .ZN(n15351) );
  NAND2_X1 U18436 ( .A1(n15351), .A2(n16304), .ZN(n15353) );
  OAI211_X1 U18437 ( .C1(n16313), .C2(n18953), .A(n15353), .B(n15352), .ZN(
        n15356) );
  NOR2_X1 U18438 ( .A1(n15354), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15355) );
  AOI211_X1 U18439 ( .C1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15362), .A(
        n15356), .B(n15355), .ZN(n15357) );
  OAI211_X1 U18440 ( .C1(n15359), .C2(n16326), .A(n15358), .B(n15357), .ZN(
        P2_U3027) );
  AOI21_X1 U18441 ( .B1(n9870), .B2(n15361), .A(n15360), .ZN(n18967) );
  INV_X1 U18442 ( .A(n15362), .ZN(n15367) );
  INV_X1 U18443 ( .A(n15458), .ZN(n15426) );
  NAND3_X1 U18444 ( .A1(n15426), .A2(n15363), .A3(n15366), .ZN(n15365) );
  AOI22_X1 U18445 ( .A1(n18966), .A2(n16304), .B1(n19223), .B2(
        P2_REIP_REG_18__SCAN_IN), .ZN(n15364) );
  OAI211_X1 U18446 ( .C1(n15367), .C2(n15366), .A(n15365), .B(n15364), .ZN(
        n15368) );
  AOI21_X1 U18447 ( .B1(n18967), .B2(n16299), .A(n15368), .ZN(n15371) );
  NAND3_X1 U18448 ( .A1(n15369), .A2(n16301), .A3(n15125), .ZN(n15370) );
  OAI211_X1 U18449 ( .C1(n15372), .C2(n15495), .A(n15371), .B(n15370), .ZN(
        P2_U3028) );
  INV_X1 U18450 ( .A(n15373), .ZN(n15391) );
  AND2_X1 U18451 ( .A1(n16326), .A2(n15374), .ZN(n15375) );
  OR2_X1 U18452 ( .A1(n15152), .A2(n15375), .ZN(n15380) );
  OR2_X1 U18453 ( .A1(n15381), .A2(n10041), .ZN(n15376) );
  NAND2_X1 U18454 ( .A1(n15445), .A2(n15376), .ZN(n15414) );
  NOR2_X1 U18455 ( .A1(n15377), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15378) );
  NOR2_X1 U18456 ( .A1(n15414), .A2(n15378), .ZN(n15379) );
  OAI21_X1 U18457 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15381), .A(
        n15404), .ZN(n15389) );
  NAND2_X1 U18458 ( .A1(n10041), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15382) );
  OAI22_X1 U18459 ( .A1(n15165), .A2(n16326), .B1(n15458), .B2(n15382), .ZN(
        n15400) );
  NAND3_X1 U18460 ( .A1(n15400), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n15383), .ZN(n15387) );
  INV_X1 U18461 ( .A(n18976), .ZN(n15385) );
  AOI21_X1 U18462 ( .B1(n15385), .B2(n16304), .A(n15384), .ZN(n15386) );
  OAI211_X1 U18463 ( .C1(n16313), .C2(n18977), .A(n15387), .B(n15386), .ZN(
        n15388) );
  AOI21_X1 U18464 ( .B1(n15389), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n15388), .ZN(n15390) );
  OAI21_X1 U18465 ( .B1(n15391), .B2(n15495), .A(n15390), .ZN(P2_U3029) );
  OR2_X1 U18466 ( .A1(n15392), .A2(n15495), .ZN(n15402) );
  AND2_X1 U18467 ( .A1(n9922), .A2(n15393), .ZN(n15395) );
  OR2_X1 U18468 ( .A1(n15395), .A2(n15394), .ZN(n19132) );
  AOI21_X1 U18469 ( .B1(n15397), .B2(n16304), .A(n15396), .ZN(n15398) );
  OAI21_X1 U18470 ( .B1(n19132), .B2(n16313), .A(n15398), .ZN(n15399) );
  AOI21_X1 U18471 ( .B1(n15400), .B2(n15403), .A(n15399), .ZN(n15401) );
  OAI211_X1 U18472 ( .C1(n15404), .C2(n15403), .A(n15402), .B(n15401), .ZN(
        P2_U3030) );
  NAND2_X1 U18473 ( .A1(n15406), .A2(n15405), .ZN(n15408) );
  XOR2_X1 U18474 ( .A(n15408), .B(n15407), .Z(n16246) );
  INV_X1 U18475 ( .A(n16246), .ZN(n15420) );
  INV_X1 U18476 ( .A(n15165), .ZN(n15409) );
  AOI21_X1 U18477 ( .B1(n15415), .B2(n15410), .A(n15409), .ZN(n16244) );
  OAI21_X1 U18478 ( .B1(n15421), .B2(n15411), .A(n9922), .ZN(n19139) );
  INV_X1 U18479 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19883) );
  NOR2_X1 U18480 ( .A1(n19883), .A2(n19040), .ZN(n15413) );
  NOR2_X1 U18481 ( .A1(n19001), .A2(n16314), .ZN(n15412) );
  AOI211_X1 U18482 ( .C1(n15414), .C2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15413), .B(n15412), .ZN(n15417) );
  NAND3_X1 U18483 ( .A1(n15426), .A2(n10041), .A3(n15415), .ZN(n15416) );
  OAI211_X1 U18484 ( .C1(n19139), .C2(n16313), .A(n15417), .B(n15416), .ZN(
        n15418) );
  AOI21_X1 U18485 ( .B1(n16244), .B2(n16301), .A(n15418), .ZN(n15419) );
  OAI21_X1 U18486 ( .B1(n15420), .B2(n15495), .A(n15419), .ZN(P2_U3031) );
  AOI21_X1 U18487 ( .B1(n15438), .B2(n15422), .A(n15421), .ZN(n19013) );
  INV_X1 U18488 ( .A(n19013), .ZN(n19141) );
  INV_X1 U18489 ( .A(n15445), .ZN(n15456) );
  OAI22_X1 U18490 ( .A1(n15423), .A2(n16314), .B1(n19881), .B2(n19083), .ZN(
        n15424) );
  AOI21_X1 U18491 ( .B1(n15456), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n15424), .ZN(n15428) );
  OAI211_X1 U18492 ( .C1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n15440), .A(
        n15426), .B(n15425), .ZN(n15427) );
  OAI211_X1 U18493 ( .C1(n19141), .C2(n16313), .A(n15428), .B(n15427), .ZN(
        n15429) );
  AOI21_X1 U18494 ( .B1(n15430), .B2(n16301), .A(n15429), .ZN(n15431) );
  OAI21_X1 U18495 ( .B1(n15432), .B2(n15495), .A(n15431), .ZN(P2_U3032) );
  AND2_X1 U18496 ( .A1(n15434), .A2(n15433), .ZN(n15435) );
  XNOR2_X1 U18497 ( .A(n15436), .B(n15435), .ZN(n16250) );
  INV_X1 U18498 ( .A(n16250), .ZN(n15449) );
  XNOR2_X1 U18499 ( .A(n15459), .B(n15437), .ZN(n16249) );
  OAI21_X1 U18500 ( .B1(n15451), .B2(n15439), .A(n15438), .ZN(n19143) );
  NOR2_X1 U18501 ( .A1(n19143), .A2(n16313), .ZN(n15447) );
  AOI211_X1 U18502 ( .C1(n15441), .C2(n15437), .A(n15440), .B(n15458), .ZN(
        n15443) );
  NOR2_X1 U18503 ( .A1(n19024), .A2(n16314), .ZN(n15442) );
  AOI211_X1 U18504 ( .C1(n19223), .C2(P2_REIP_REG_13__SCAN_IN), .A(n15443), 
        .B(n15442), .ZN(n15444) );
  OAI21_X1 U18505 ( .B1(n15445), .B2(n15437), .A(n15444), .ZN(n15446) );
  AOI211_X1 U18506 ( .C1(n16249), .C2(n16301), .A(n15447), .B(n15446), .ZN(
        n15448) );
  OAI21_X1 U18507 ( .B1(n15495), .B2(n15449), .A(n15448), .ZN(P2_U3033) );
  AOI21_X1 U18508 ( .B1(n15450), .B2(n15452), .A(n15451), .ZN(n19144) );
  NAND2_X1 U18509 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n19223), .ZN(n15453) );
  OAI21_X1 U18510 ( .B1(n16314), .B2(n15454), .A(n15453), .ZN(n15455) );
  AOI21_X1 U18511 ( .B1(n15456), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15455), .ZN(n15457) );
  OAI21_X1 U18512 ( .B1(n15458), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15457), .ZN(n15462) );
  NOR3_X1 U18513 ( .A1(n15460), .A2(n15459), .A3(n16326), .ZN(n15461) );
  AOI211_X1 U18514 ( .C1(n16299), .C2(n19144), .A(n15462), .B(n15461), .ZN(
        n15463) );
  OAI21_X1 U18515 ( .B1(n15495), .B2(n15464), .A(n15463), .ZN(P2_U3034) );
  OR2_X1 U18516 ( .A1(n15466), .A2(n10103), .ZN(n15467) );
  XNOR2_X1 U18517 ( .A(n15468), .B(n15467), .ZN(n16257) );
  INV_X1 U18518 ( .A(n16257), .ZN(n15482) );
  OAI21_X1 U18519 ( .B1(n15470), .B2(n15469), .A(n15450), .ZN(n19149) );
  INV_X1 U18520 ( .A(n19149), .ZN(n15480) );
  XNOR2_X1 U18521 ( .A(n15471), .B(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15472) );
  NAND2_X1 U18522 ( .A1(n15485), .A2(n15472), .ZN(n15475) );
  NOR2_X1 U18523 ( .A1(n15473), .A2(n15500), .ZN(n15486) );
  AOI22_X1 U18524 ( .A1(n19223), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15486), .ZN(n15474) );
  OAI211_X1 U18525 ( .C1(n19049), .C2(n16314), .A(n15475), .B(n15474), .ZN(
        n15479) );
  OR2_X1 U18526 ( .A1(n15199), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15476) );
  NAND2_X1 U18527 ( .A1(n15477), .A2(n15476), .ZN(n16256) );
  NOR2_X1 U18528 ( .A1(n16256), .A2(n16326), .ZN(n15478) );
  AOI211_X1 U18529 ( .C1(n16299), .C2(n15480), .A(n15479), .B(n15478), .ZN(
        n15481) );
  OAI21_X1 U18530 ( .B1(n15482), .B2(n15495), .A(n15481), .ZN(P2_U3035) );
  XNOR2_X1 U18531 ( .A(n15484), .B(n15483), .ZN(n19152) );
  NAND2_X1 U18532 ( .A1(n15485), .A2(n15488), .ZN(n15491) );
  INV_X1 U18533 ( .A(n15486), .ZN(n15487) );
  OAI22_X1 U18534 ( .A1(n19040), .A2(n19873), .B1(n15488), .B2(n15487), .ZN(
        n15489) );
  AOI21_X1 U18535 ( .B1(n16304), .B2(n19061), .A(n15489), .ZN(n15490) );
  OAI211_X1 U18536 ( .C1(n19152), .C2(n16313), .A(n15491), .B(n15490), .ZN(
        n15492) );
  AOI21_X1 U18537 ( .B1(n15493), .B2(n16301), .A(n15492), .ZN(n15494) );
  OAI21_X1 U18538 ( .B1(n15496), .B2(n15495), .A(n15494), .ZN(P2_U3036) );
  OR2_X1 U18539 ( .A1(n15497), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15498) );
  NAND2_X1 U18540 ( .A1(n15198), .A2(n15498), .ZN(n16268) );
  OAI22_X1 U18541 ( .A1(n16314), .A2(n15499), .B1(n14799), .B2(n19083), .ZN(
        n15503) );
  AOI21_X1 U18542 ( .B1(n13826), .B2(n15501), .A(n15500), .ZN(n15502) );
  AOI211_X1 U18543 ( .C1(n15504), .C2(n16299), .A(n15503), .B(n15502), .ZN(
        n15509) );
  NAND2_X1 U18544 ( .A1(n15506), .A2(n15505), .ZN(n15507) );
  XNOR2_X1 U18545 ( .A(n9901), .B(n15507), .ZN(n16264) );
  NAND2_X1 U18546 ( .A1(n16264), .A2(n16322), .ZN(n15508) );
  OAI211_X1 U18547 ( .C1(n16268), .C2(n16326), .A(n15509), .B(n15508), .ZN(
        P2_U3037) );
  NOR2_X1 U18548 ( .A1(n19867), .A2(n19040), .ZN(n15510) );
  AOI221_X1 U18549 ( .B1(n16307), .B2(n15511), .C1(n16300), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n15510), .ZN(n15512) );
  INV_X1 U18550 ( .A(n15512), .ZN(n15517) );
  OR2_X1 U18551 ( .A1(n15514), .A2(n15513), .ZN(n15515) );
  NAND2_X1 U18552 ( .A1(n15515), .A2(n16297), .ZN(n19158) );
  OAI22_X1 U18553 ( .A1(n19158), .A2(n16313), .B1(n16314), .B2(n19086), .ZN(
        n15516) );
  AOI211_X1 U18554 ( .C1(n15518), .C2(n16322), .A(n15517), .B(n15516), .ZN(
        n15519) );
  OAI21_X1 U18555 ( .B1(n16326), .B2(n15520), .A(n15519), .ZN(P2_U3039) );
  INV_X1 U18556 ( .A(n15521), .ZN(n15522) );
  NAND2_X1 U18557 ( .A1(n15523), .A2(n15522), .ZN(n15531) );
  MUX2_X1 U18558 ( .A(n15531), .B(n9821), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n15524) );
  AOI21_X1 U18559 ( .B1(n15525), .B2(n15550), .A(n15524), .ZN(n16331) );
  INV_X1 U18560 ( .A(n16331), .ZN(n15528) );
  AOI22_X1 U18561 ( .A1(n10145), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n15526), .B2(n13535), .ZN(n15539) );
  AOI222_X1 U18562 ( .A1(n15528), .A2(n15553), .B1(n15527), .B2(n16365), .C1(
        P2_STATE2_REG_1__SCAN_IN), .C2(n15539), .ZN(n15530) );
  NAND2_X1 U18563 ( .A1(n15557), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15529) );
  OAI21_X1 U18564 ( .B1(n15530), .B2(n15557), .A(n15529), .ZN(P2_U3601) );
  INV_X1 U18565 ( .A(n16365), .ZN(n15556) );
  OAI21_X1 U18566 ( .B1(n15532), .B2(n10478), .A(n15531), .ZN(n15535) );
  NAND2_X1 U18567 ( .A1(n9821), .A2(n15533), .ZN(n15534) );
  NAND2_X1 U18568 ( .A1(n15535), .A2(n15534), .ZN(n15536) );
  AOI21_X1 U18569 ( .B1(n13191), .B2(n15550), .A(n15536), .ZN(n16332) );
  INV_X1 U18570 ( .A(n15553), .ZN(n19925) );
  OAI21_X1 U18571 ( .B1(n13535), .B2(n15538), .A(n15537), .ZN(n15551) );
  NOR2_X1 U18572 ( .A1(n15539), .A2(n19832), .ZN(n15552) );
  INV_X1 U18573 ( .A(n15552), .ZN(n15540) );
  OAI222_X1 U18574 ( .A1(n15556), .A2(n19949), .B1(n16332), .B2(n19925), .C1(
        n15551), .C2(n15540), .ZN(n15541) );
  MUX2_X1 U18575 ( .A(n15541), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n15557), .Z(P2_U3600) );
  OAI21_X1 U18576 ( .B1(n12868), .B2(n15548), .A(n15542), .ZN(n15546) );
  OR2_X1 U18577 ( .A1(n15544), .A2(n15543), .ZN(n15545) );
  OAI211_X1 U18578 ( .C1(n15548), .C2(n15547), .A(n15546), .B(n15545), .ZN(
        n15549) );
  AOI21_X1 U18579 ( .B1(n13542), .B2(n15550), .A(n15549), .ZN(n16328) );
  INV_X1 U18580 ( .A(n16328), .ZN(n15554) );
  AOI22_X1 U18581 ( .A1(n15554), .A2(n15553), .B1(n15552), .B2(n15551), .ZN(
        n15555) );
  OAI21_X1 U18582 ( .B1(n19936), .B2(n15556), .A(n15555), .ZN(n15558) );
  INV_X1 U18583 ( .A(n15557), .ZN(n15664) );
  MUX2_X1 U18584 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n15558), .S(
        n15664), .Z(P2_U3599) );
  NOR2_X1 U18585 ( .A1(n17351), .A2(n17070), .ZN(n17058) );
  NAND2_X1 U18586 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17058), .ZN(n17000) );
  NOR2_X1 U18587 ( .A1(n17000), .A2(n15560), .ZN(n17005) );
  NAND2_X1 U18588 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17005), .ZN(n16994) );
  INV_X1 U18589 ( .A(n16994), .ZN(n16999) );
  NAND2_X1 U18590 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16999), .ZN(n15636) );
  AND3_X1 U18591 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(n16999), .ZN(n16988) );
  NOR2_X1 U18592 ( .A1(n17261), .A2(n16988), .ZN(n16989) );
  AOI22_X1 U18593 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15691), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15564) );
  AOI22_X1 U18594 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17019), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15563) );
  AOI22_X1 U18595 ( .A1(n9820), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17197), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15562) );
  AOI22_X1 U18596 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13703), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15561) );
  NAND4_X1 U18597 ( .A1(n15564), .A2(n15563), .A3(n15562), .A4(n15561), .ZN(
        n15570) );
  AOI22_X1 U18598 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n15699), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15568) );
  AOI22_X1 U18599 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15567) );
  AOI22_X1 U18600 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15566) );
  AOI22_X1 U18601 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15565) );
  NAND4_X1 U18602 ( .A1(n15568), .A2(n15567), .A3(n15566), .A4(n15565), .ZN(
        n15569) );
  NOR2_X1 U18603 ( .A1(n15570), .A2(n15569), .ZN(n15634) );
  AOI22_X1 U18604 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n16962), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15574) );
  AOI22_X1 U18605 ( .A1(n17197), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15573) );
  AOI22_X1 U18606 ( .A1(n9820), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17019), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15572) );
  AOI22_X1 U18607 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15571) );
  NAND4_X1 U18608 ( .A1(n15574), .A2(n15573), .A3(n15572), .A4(n15571), .ZN(
        n15580) );
  AOI22_X1 U18609 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15578) );
  AOI22_X1 U18610 ( .A1(n17208), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15577) );
  AOI22_X1 U18611 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n15699), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15576) );
  AOI22_X1 U18612 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n15691), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15575) );
  NAND4_X1 U18613 ( .A1(n15578), .A2(n15577), .A3(n15576), .A4(n15575), .ZN(
        n15579) );
  NOR2_X1 U18614 ( .A1(n15580), .A2(n15579), .ZN(n16996) );
  AOI22_X1 U18615 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15585) );
  AOI22_X1 U18616 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n15584) );
  AOI22_X1 U18617 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15583) );
  AOI22_X1 U18618 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17019), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15582) );
  NAND4_X1 U18619 ( .A1(n15585), .A2(n15584), .A3(n15583), .A4(n15582), .ZN(
        n15591) );
  AOI22_X1 U18620 ( .A1(n9820), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n15691), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15589) );
  AOI22_X1 U18621 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15588) );
  AOI22_X1 U18622 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n15587) );
  AOI22_X1 U18623 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n15699), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n15586) );
  NAND4_X1 U18624 ( .A1(n15589), .A2(n15588), .A3(n15587), .A4(n15586), .ZN(
        n15590) );
  NOR2_X1 U18625 ( .A1(n15591), .A2(n15590), .ZN(n17007) );
  AOI22_X1 U18626 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15601) );
  AOI22_X1 U18627 ( .A1(n9820), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15600) );
  AOI22_X1 U18628 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n15699), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15592) );
  OAI21_X1 U18629 ( .B1(n16970), .B2(n15746), .A(n15592), .ZN(n15598) );
  AOI22_X1 U18630 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17019), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15596) );
  AOI22_X1 U18631 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15595) );
  AOI22_X1 U18632 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15594) );
  AOI22_X1 U18633 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n15691), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15593) );
  NAND4_X1 U18634 ( .A1(n15596), .A2(n15595), .A3(n15594), .A4(n15593), .ZN(
        n15597) );
  AOI211_X1 U18635 ( .C1(n16962), .C2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n15598), .B(n15597), .ZN(n15599) );
  NAND3_X1 U18636 ( .A1(n15601), .A2(n15600), .A3(n15599), .ZN(n17013) );
  AOI22_X1 U18637 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n17179), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n17145), .ZN(n15613) );
  AOI22_X1 U18638 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n17188), .B1(
        n17019), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15612) );
  INV_X1 U18639 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17228) );
  AOI22_X1 U18640 ( .A1(n9820), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15602) );
  OAI21_X1 U18641 ( .B1(n17228), .B2(n17018), .A(n15602), .ZN(n15610) );
  AOI22_X1 U18642 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15608) );
  AOI22_X1 U18643 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n16962), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15607) );
  AOI22_X1 U18644 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n17143), .ZN(n15606) );
  AOI22_X1 U18645 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15605) );
  NAND4_X1 U18646 ( .A1(n15608), .A2(n15607), .A3(n15606), .A4(n15605), .ZN(
        n15609) );
  AOI211_X1 U18647 ( .C1(n17195), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n15610), .B(n15609), .ZN(n15611) );
  NAND3_X1 U18648 ( .A1(n15613), .A2(n15612), .A3(n15611), .ZN(n17014) );
  NAND2_X1 U18649 ( .A1(n17013), .A2(n17014), .ZN(n17012) );
  NOR2_X1 U18650 ( .A1(n17007), .A2(n17012), .ZN(n17006) );
  AOI22_X1 U18651 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15623) );
  AOI22_X1 U18652 ( .A1(n17208), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15622) );
  INV_X1 U18653 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17254) );
  AOI22_X1 U18654 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15691), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15614) );
  OAI21_X1 U18655 ( .B1(n16970), .B2(n17254), .A(n15614), .ZN(n15620) );
  AOI22_X1 U18656 ( .A1(n9820), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15618) );
  AOI22_X1 U18657 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n15699), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15617) );
  AOI22_X1 U18658 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13703), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15616) );
  AOI22_X1 U18659 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n16962), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15615) );
  NAND4_X1 U18660 ( .A1(n15618), .A2(n15617), .A3(n15616), .A4(n15615), .ZN(
        n15619) );
  AOI211_X1 U18661 ( .C1(n17195), .C2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n15620), .B(n15619), .ZN(n15621) );
  NAND3_X1 U18662 ( .A1(n15623), .A2(n15622), .A3(n15621), .ZN(n17003) );
  NAND2_X1 U18663 ( .A1(n17006), .A2(n17003), .ZN(n17002) );
  NOR2_X1 U18664 ( .A1(n16996), .A2(n17002), .ZN(n16995) );
  AOI22_X1 U18665 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17019), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15633) );
  AOI22_X1 U18666 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n15691), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15632) );
  INV_X1 U18667 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17242) );
  AOI22_X1 U18668 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15624) );
  OAI21_X1 U18669 ( .B1(n16970), .B2(n17242), .A(n15624), .ZN(n15630) );
  AOI22_X1 U18670 ( .A1(n9820), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15628) );
  AOI22_X1 U18671 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15627) );
  AOI22_X1 U18672 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13703), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15626) );
  AOI22_X1 U18673 ( .A1(n17208), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15699), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15625) );
  NAND4_X1 U18674 ( .A1(n15628), .A2(n15627), .A3(n15626), .A4(n15625), .ZN(
        n15629) );
  AOI211_X1 U18675 ( .C1(n17194), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n15630), .B(n15629), .ZN(n15631) );
  NAND3_X1 U18676 ( .A1(n15633), .A2(n15632), .A3(n15631), .ZN(n16992) );
  NAND2_X1 U18677 ( .A1(n16995), .A2(n16992), .ZN(n16991) );
  NOR2_X1 U18678 ( .A1(n15634), .A2(n16991), .ZN(n16986) );
  AOI21_X1 U18679 ( .B1(n15634), .B2(n16991), .A(n16986), .ZN(n17280) );
  AOI22_X1 U18680 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16989), .B1(n17280), 
        .B2(n17261), .ZN(n15635) );
  OAI21_X1 U18681 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n15636), .A(n15635), .ZN(
        P3_U2675) );
  AOI22_X1 U18682 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15691), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15647) );
  AOI22_X1 U18683 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15646) );
  INV_X1 U18684 ( .A(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15638) );
  AOI22_X1 U18685 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n16962), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15637) );
  OAI21_X1 U18686 ( .B1(n9871), .B2(n15638), .A(n15637), .ZN(n15644) );
  AOI22_X1 U18687 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17019), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15642) );
  AOI22_X1 U18688 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15641) );
  AOI22_X1 U18689 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13703), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15640) );
  AOI22_X1 U18690 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n15699), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15639) );
  NAND4_X1 U18691 ( .A1(n15642), .A2(n15641), .A3(n15640), .A4(n15639), .ZN(
        n15643) );
  AOI211_X1 U18692 ( .C1(n9820), .C2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A(
        n15644), .B(n15643), .ZN(n15645) );
  NAND3_X1 U18693 ( .A1(n15647), .A2(n15646), .A3(n15645), .ZN(n17357) );
  INV_X1 U18694 ( .A(n17357), .ZN(n15652) );
  INV_X1 U18695 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17172) );
  INV_X1 U18696 ( .A(n17244), .ZN(n17236) );
  NAND2_X1 U18697 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17226), .ZN(n17204) );
  NOR2_X1 U18698 ( .A1(n17172), .A2(n17204), .ZN(n17187) );
  NAND2_X1 U18699 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n17187), .ZN(n17169) );
  INV_X1 U18700 ( .A(n17169), .ZN(n17141) );
  AND2_X1 U18701 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17141), .ZN(n17158) );
  NAND2_X1 U18702 ( .A1(n15650), .A2(n17226), .ZN(n17102) );
  OAI21_X1 U18703 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17158), .A(n17102), .ZN(
        n15651) );
  AOI22_X1 U18704 ( .A1(n17261), .A2(n15652), .B1(n15651), .B2(n17246), .ZN(
        P3_U2690) );
  NAND2_X1 U18705 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18401) );
  AOI221_X1 U18706 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18401), .C1(n15654), 
        .C2(n18401), .A(n15653), .ZN(n18228) );
  NOR2_X1 U18707 ( .A1(n15655), .A2(n18699), .ZN(n15656) );
  OAI21_X1 U18708 ( .B1(n15656), .B2(n18520), .A(n18229), .ZN(n18226) );
  AOI22_X1 U18709 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18228), .B1(
        n18226), .B2(n18712), .ZN(P3_U2865) );
  INV_X1 U18710 ( .A(n15657), .ZN(n15660) );
  INV_X1 U18711 ( .A(n15658), .ZN(n16343) );
  NOR2_X1 U18712 ( .A1(n19925), .A2(n16343), .ZN(n15659) );
  NAND4_X1 U18713 ( .A1(n15661), .A2(n15664), .A3(n15660), .A4(n15659), .ZN(
        n15662) );
  OAI21_X1 U18714 ( .B1(n15664), .B2(n15663), .A(n15662), .ZN(P2_U3595) );
  INV_X1 U18715 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16407) );
  AOI22_X1 U18716 ( .A1(n17197), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n16962), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15675) );
  AOI22_X1 U18717 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15674) );
  AOI22_X1 U18718 ( .A1(n9820), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15666) );
  OAI21_X1 U18719 ( .B1(n9871), .B2(n17228), .A(n15666), .ZN(n15672) );
  AOI22_X1 U18720 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15670) );
  AOI22_X1 U18721 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13703), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15669) );
  AOI22_X1 U18722 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n15691), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15668) );
  AOI22_X1 U18723 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n15699), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15667) );
  NAND4_X1 U18724 ( .A1(n15670), .A2(n15669), .A3(n15668), .A4(n15667), .ZN(
        n15671) );
  AOI211_X1 U18725 ( .C1(n17196), .C2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n15672), .B(n15671), .ZN(n15673) );
  NAND3_X1 U18726 ( .A1(n15675), .A2(n15674), .A3(n15673), .ZN(n17382) );
  AOI22_X1 U18727 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15680) );
  AOI22_X1 U18728 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13697), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15679) );
  AOI22_X1 U18729 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15699), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15678) );
  AOI22_X1 U18730 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15677) );
  NAND4_X1 U18731 ( .A1(n15680), .A2(n15679), .A3(n15678), .A4(n15677), .ZN(
        n15686) );
  AOI22_X1 U18732 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15684) );
  AOI22_X1 U18733 ( .A1(n17197), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15683) );
  AOI22_X1 U18734 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15691), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15682) );
  AOI22_X1 U18735 ( .A1(n9820), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17019), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15681) );
  NAND4_X1 U18736 ( .A1(n15684), .A2(n15683), .A3(n15682), .A4(n15681), .ZN(
        n15685) );
  AOI22_X1 U18737 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15690) );
  AOI22_X1 U18738 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15689) );
  INV_X2 U18739 ( .A(n9883), .ZN(n17207) );
  AOI22_X1 U18740 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15688) );
  AOI22_X1 U18741 ( .A1(n9820), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15687) );
  NAND4_X1 U18742 ( .A1(n15690), .A2(n15689), .A3(n15688), .A4(n15687), .ZN(
        n15697) );
  AOI22_X1 U18743 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n15691), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15695) );
  AOI22_X1 U18744 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15699), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15694) );
  AOI22_X1 U18745 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15693) );
  AOI22_X1 U18746 ( .A1(n17197), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13703), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15692) );
  NAND4_X1 U18747 ( .A1(n15695), .A2(n15694), .A3(n15693), .A4(n15692), .ZN(
        n15696) );
  AOI22_X1 U18748 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15709) );
  AOI22_X1 U18749 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n15691), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15708) );
  INV_X1 U18750 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17256) );
  AOI22_X1 U18751 ( .A1(n15665), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n15581), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15698) );
  OAI21_X1 U18752 ( .B1(n9871), .B2(n17256), .A(n15698), .ZN(n15706) );
  AOI22_X1 U18753 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13698), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n15704) );
  AOI22_X1 U18754 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n15699), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15703) );
  AOI22_X1 U18755 ( .A1(n9820), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n15700), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n15702) );
  AOI22_X1 U18756 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15701) );
  NAND4_X1 U18757 ( .A1(n15704), .A2(n15703), .A3(n15702), .A4(n15701), .ZN(
        n15705) );
  AOI211_X1 U18758 ( .C1(n13697), .C2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n15706), .B(n15705), .ZN(n15707) );
  NAND3_X1 U18759 ( .A1(n15709), .A2(n15708), .A3(n15707), .ZN(n15819) );
  AOI22_X1 U18760 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15720) );
  AOI22_X1 U18761 ( .A1(n9820), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17146), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15719) );
  AOI22_X1 U18762 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n15711), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15712) );
  OAI21_X1 U18763 ( .B1(n9871), .B2(n17254), .A(n15712), .ZN(n15718) );
  AOI22_X1 U18764 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n15691), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15717) );
  AOI22_X1 U18765 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15716) );
  AOI22_X1 U18766 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17179), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15715) );
  AOI22_X1 U18767 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15714) );
  NAND2_X1 U18768 ( .A1(n15819), .A2(n17401), .ZN(n15818) );
  AOI22_X1 U18769 ( .A1(n9820), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15730) );
  AOI22_X1 U18770 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15729) );
  AOI22_X1 U18771 ( .A1(n17208), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15721) );
  OAI21_X1 U18772 ( .B1(n9871), .B2(n17242), .A(n15721), .ZN(n15727) );
  AOI22_X1 U18773 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13703), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15725) );
  AOI22_X1 U18774 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16962), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15724) );
  AOI22_X1 U18775 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n15691), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15723) );
  AOI22_X1 U18776 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17179), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15722) );
  NAND4_X1 U18777 ( .A1(n15725), .A2(n15724), .A3(n15723), .A4(n15722), .ZN(
        n15726) );
  AOI211_X1 U18778 ( .C1(n17197), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n15727), .B(n15726), .ZN(n15728) );
  NAND3_X1 U18779 ( .A1(n15730), .A2(n15729), .A3(n15728), .ZN(n15813) );
  NAND2_X1 U18780 ( .A1(n15743), .A2(n15813), .ZN(n15760) );
  AOI22_X1 U18781 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9820), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n15740) );
  AOI22_X1 U18782 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n15739) );
  INV_X1 U18783 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17232) );
  AOI22_X1 U18784 ( .A1(n13703), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n15731) );
  OAI21_X1 U18785 ( .B1(n9871), .B2(n17232), .A(n15731), .ZN(n15737) );
  AOI22_X1 U18786 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15735) );
  AOI22_X1 U18787 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n15734) );
  AOI22_X1 U18788 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n15733) );
  AOI22_X1 U18789 ( .A1(n17179), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15732) );
  NAND4_X1 U18790 ( .A1(n15735), .A2(n15734), .A3(n15733), .A4(n15732), .ZN(
        n15736) );
  AOI211_X1 U18791 ( .C1(n17174), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n15737), .B(n15736), .ZN(n15738) );
  NAND3_X1 U18792 ( .A1(n15740), .A2(n15739), .A3(n15738), .ZN(n17815) );
  NOR2_X4 U18793 ( .A1(n16392), .A2(n16440), .ZN(n17798) );
  INV_X1 U18794 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17528) );
  NAND2_X1 U18795 ( .A1(n17760), .A2(n17528), .ZN(n16438) );
  INV_X1 U18796 ( .A(n16438), .ZN(n15897) );
  INV_X1 U18797 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17929) );
  INV_X1 U18798 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18034) );
  INV_X1 U18799 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18146) );
  INV_X1 U18800 ( .A(n16440), .ZN(n15741) );
  OAI21_X1 U18801 ( .B1(n15741), .B2(n17382), .A(n17760), .ZN(n15765) );
  XOR2_X1 U18802 ( .A(n15742), .B(n17815), .Z(n15764) );
  INV_X1 U18803 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18171) );
  NOR2_X1 U18804 ( .A1(n18171), .A2(n15744), .ZN(n15759) );
  NOR2_X1 U18805 ( .A1(n15756), .A2(n15757), .ZN(n15758) );
  INV_X1 U18806 ( .A(n15819), .ZN(n17412) );
  INV_X1 U18807 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18845) );
  AOI22_X1 U18808 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15691), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15755) );
  AOI22_X1 U18809 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15754) );
  AOI22_X1 U18810 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15745) );
  OAI21_X1 U18811 ( .B1(n9871), .B2(n15746), .A(n15745), .ZN(n15752) );
  AOI22_X1 U18812 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n15711), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15750) );
  AOI22_X1 U18813 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15749) );
  AOI22_X1 U18814 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17179), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15748) );
  AOI22_X1 U18815 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15747) );
  NAND4_X1 U18816 ( .A1(n15750), .A2(n15749), .A3(n15748), .A4(n15747), .ZN(
        n15751) );
  AOI211_X1 U18817 ( .C1(n9820), .C2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A(
        n15752), .B(n15751), .ZN(n15753) );
  NAND3_X1 U18818 ( .A1(n15755), .A2(n15754), .A3(n15753), .ZN(n15917) );
  NAND2_X1 U18819 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15917), .ZN(
        n17893) );
  NOR2_X1 U18820 ( .A1(n17883), .A2(n17893), .ZN(n17882) );
  AOI21_X1 U18821 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n17412), .A(
        n17882), .ZN(n17874) );
  NOR2_X1 U18822 ( .A1(n17874), .A2(n17873), .ZN(n17872) );
  XNOR2_X1 U18823 ( .A(n15818), .B(n17397), .ZN(n17865) );
  XNOR2_X1 U18824 ( .A(n15760), .B(n17390), .ZN(n15762) );
  NOR2_X1 U18825 ( .A1(n15761), .A2(n15762), .ZN(n15763) );
  INV_X1 U18826 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17837) );
  XNOR2_X1 U18827 ( .A(n15762), .B(n15761), .ZN(n17836) );
  INV_X1 U18828 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18157) );
  XOR2_X1 U18829 ( .A(n18157), .B(n15764), .Z(n17824) );
  XNOR2_X1 U18830 ( .A(n15765), .B(n17679), .ZN(n17811) );
  NOR2_X1 U18831 ( .A1(n17679), .A2(n15765), .ZN(n15766) );
  INV_X1 U18832 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18135) );
  NAND2_X1 U18833 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18103) );
  NOR2_X1 U18834 ( .A1(n18103), .A2(n17758), .ZN(n18074) );
  NAND2_X1 U18835 ( .A1(n18074), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18055) );
  INV_X1 U18836 ( .A(n18055), .ZN(n18053) );
  NAND2_X1 U18837 ( .A1(n18053), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18058) );
  INV_X1 U18838 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17714) );
  NOR2_X1 U18839 ( .A1(n18058), .A2(n17714), .ZN(n18038) );
  NAND2_X1 U18840 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18038), .ZN(
        n16450) );
  NOR2_X1 U18841 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n10026), .ZN(
        n15769) );
  INV_X1 U18842 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18113) );
  INV_X1 U18843 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17764) );
  NAND2_X1 U18844 ( .A1(n18113), .A2(n17764), .ZN(n17763) );
  INV_X1 U18845 ( .A(n17763), .ZN(n17766) );
  NOR4_X1 U18846 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15768) );
  INV_X1 U18847 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18050) );
  NAND4_X1 U18848 ( .A1(n15769), .A2(n17766), .A3(n15768), .A4(n18050), .ZN(
        n15770) );
  NAND2_X1 U18849 ( .A1(n17760), .A2(n15770), .ZN(n15774) );
  OAI221_X1 U18850 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17760), 
        .C1(n18034), .C2(n15772), .A(n15774), .ZN(n17672) );
  INV_X1 U18851 ( .A(n15772), .ZN(n15773) );
  NAND2_X1 U18852 ( .A1(n15774), .A2(n15773), .ZN(n15778) );
  INV_X1 U18853 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18020) );
  NOR2_X1 U18854 ( .A1(n18034), .A2(n18020), .ZN(n17662) );
  INV_X1 U18855 ( .A(n17662), .ZN(n18013) );
  INV_X1 U18856 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17655) );
  INV_X1 U18857 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17968) );
  NAND2_X1 U18858 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17970) );
  NOR3_X1 U18859 ( .A1(n17655), .A2(n17968), .A3(n17970), .ZN(n17600) );
  NAND2_X1 U18860 ( .A1(n17600), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17901) );
  INV_X1 U18861 ( .A(n17901), .ZN(n17927) );
  NAND2_X1 U18862 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17927), .ZN(
        n17578) );
  NOR2_X1 U18863 ( .A1(n18013), .A2(n17578), .ZN(n15837) );
  NOR2_X1 U18864 ( .A1(n17798), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17663) );
  INV_X1 U18865 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17999) );
  NAND2_X1 U18866 ( .A1(n17663), .A2(n17999), .ZN(n15775) );
  NOR2_X1 U18867 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15775), .ZN(
        n17623) );
  NAND2_X1 U18868 ( .A1(n17623), .A2(n17968), .ZN(n17606) );
  NAND2_X1 U18869 ( .A1(n15776), .A2(n10360), .ZN(n15777) );
  OR2_X1 U18870 ( .A1(n17798), .A2(n17579), .ZN(n17565) );
  OAI221_X1 U18871 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17760), 
        .C1(n17929), .C2(n17566), .A(n17565), .ZN(n17553) );
  NOR2_X1 U18872 ( .A1(n17566), .A2(n17760), .ZN(n15780) );
  INV_X1 U18873 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17923) );
  NOR2_X1 U18874 ( .A1(n17929), .A2(n17923), .ZN(n15838) );
  INV_X1 U18875 ( .A(n15838), .ZN(n17906) );
  NAND2_X1 U18876 ( .A1(n17798), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16437) );
  AOI21_X1 U18877 ( .B1(n15897), .B2(n17540), .A(n15896), .ZN(n15783) );
  XNOR2_X1 U18878 ( .A(n16407), .B(n15783), .ZN(n16423) );
  NAND2_X1 U18879 ( .A1(n18244), .A2(n16578), .ZN(n15792) );
  NOR2_X1 U18880 ( .A1(n18263), .A2(n15792), .ZN(n15799) );
  INV_X1 U18881 ( .A(n15784), .ZN(n15785) );
  OAI21_X1 U18882 ( .B1(n15786), .B2(n15785), .A(n15795), .ZN(n18674) );
  INV_X1 U18883 ( .A(n18674), .ZN(n15790) );
  AOI21_X1 U18884 ( .B1(n18253), .B2(n15787), .A(n16376), .ZN(n15789) );
  AOI21_X1 U18885 ( .B1(n18889), .B2(n15791), .A(n18751), .ZN(n15793) );
  INV_X1 U18886 ( .A(n18890), .ZN(n18884) );
  AOI21_X1 U18887 ( .B1(n15793), .B2(n15792), .A(n18884), .ZN(n16556) );
  NAND3_X1 U18888 ( .A1(n15795), .A2(n16556), .A3(n15794), .ZN(n15796) );
  NAND2_X1 U18889 ( .A1(n15799), .A2(n15798), .ZN(n16441) );
  INV_X1 U18890 ( .A(n16441), .ZN(n18675) );
  NAND2_X1 U18891 ( .A1(n17382), .A2(n18675), .ZN(n17918) );
  NOR2_X2 U18892 ( .A1(n18207), .A2(n17918), .ZN(n18138) );
  OR3_X2 U18893 ( .A1(n18900), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18201) );
  INV_X2 U18894 ( .A(n18201), .ZN(n18218) );
  NOR2_X2 U18895 ( .A1(n15800), .A2(n15806), .ZN(n18696) );
  INV_X2 U18896 ( .A(n18696), .ZN(n18683) );
  XNOR2_X1 U18897 ( .A(n16578), .B(n17415), .ZN(n18902) );
  NOR2_X4 U18898 ( .A1(n18683), .A2(n18684), .ZN(n18112) );
  INV_X1 U18899 ( .A(n18112), .ZN(n17969) );
  NAND2_X1 U18900 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17925) );
  NOR2_X1 U18901 ( .A1(n17906), .A2(n17925), .ZN(n15807) );
  INV_X1 U18902 ( .A(n15807), .ZN(n17903) );
  NOR3_X1 U18903 ( .A1(n18171), .A2(n10170), .A3(n17837), .ZN(n18158) );
  NAND2_X1 U18904 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18158), .ZN(
        n18005) );
  NOR2_X1 U18905 ( .A1(n18146), .A2(n18005), .ZN(n18126) );
  NAND2_X1 U18906 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18126), .ZN(
        n15808) );
  NAND2_X1 U18907 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18129) );
  NOR2_X1 U18908 ( .A1(n15808), .A2(n18129), .ZN(n18027) );
  NAND2_X1 U18909 ( .A1(n10173), .A2(n18027), .ZN(n18009) );
  NOR2_X1 U18910 ( .A1(n18013), .A2(n18009), .ZN(n16451) );
  NAND2_X1 U18911 ( .A1(n17927), .A2(n16451), .ZN(n17904) );
  NOR2_X1 U18912 ( .A1(n17903), .A2(n17904), .ZN(n15844) );
  NOR3_X1 U18913 ( .A1(n15803), .A2(n15802), .A3(n18889), .ZN(n15805) );
  NOR2_X1 U18914 ( .A1(n15805), .A2(n15804), .ZN(n18686) );
  AND2_X1 U18915 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18027), .ZN(
        n18096) );
  NAND2_X1 U18916 ( .A1(n10173), .A2(n18096), .ZN(n18028) );
  NAND2_X1 U18917 ( .A1(n17662), .A2(n17600), .ZN(n17967) );
  NOR2_X1 U18918 ( .A1(n18028), .A2(n17967), .ZN(n17972) );
  NAND3_X1 U18919 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n15807), .A3(
        n17972), .ZN(n15845) );
  AOI21_X1 U18920 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18127) );
  NOR2_X1 U18921 ( .A1(n15808), .A2(n18127), .ZN(n18073) );
  INV_X1 U18922 ( .A(n18073), .ZN(n18054) );
  NOR3_X1 U18923 ( .A1(n18013), .A2(n16450), .A3(n18054), .ZN(n18011) );
  NAND2_X1 U18924 ( .A1(n17927), .A2(n18011), .ZN(n17947) );
  NOR2_X1 U18925 ( .A1(n17947), .A2(n17903), .ZN(n15843) );
  NOR2_X1 U18926 ( .A1(n15843), .A2(n18709), .ZN(n17905) );
  AOI221_X1 U18927 ( .B1(n15781), .B2(n18694), .C1(n15845), .C2(n18694), .A(
        n17905), .ZN(n15809) );
  OAI211_X1 U18928 ( .C1(n18696), .C2(n15844), .A(n15809), .B(n18194), .ZN(
        n15901) );
  AOI21_X1 U18929 ( .B1(n17969), .B2(n15781), .A(n15901), .ZN(n16448) );
  NAND2_X1 U18930 ( .A1(n18132), .A2(n17528), .ZN(n15840) );
  NAND2_X1 U18931 ( .A1(n18037), .A2(n18214), .ZN(n18212) );
  NOR2_X1 U18932 ( .A1(n15781), .A2(n17528), .ZN(n16418) );
  NAND2_X1 U18933 ( .A1(n16418), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16427) );
  INV_X1 U18934 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17581) );
  INV_X1 U18935 ( .A(n17815), .ZN(n17816) );
  INV_X1 U18936 ( .A(n15813), .ZN(n17393) );
  INV_X1 U18937 ( .A(n17397), .ZN(n15815) );
  INV_X1 U18938 ( .A(n15917), .ZN(n15820) );
  NOR2_X1 U18939 ( .A1(n17412), .A2(n15820), .ZN(n15821) );
  OR2_X1 U18940 ( .A1(n17401), .A2(n15821), .ZN(n15817) );
  NAND2_X1 U18941 ( .A1(n15815), .A2(n15817), .ZN(n15812) );
  INV_X1 U18942 ( .A(n17819), .ZN(n17817) );
  NAND2_X1 U18943 ( .A1(n15829), .A2(n17382), .ZN(n15830) );
  XOR2_X1 U18944 ( .A(n17815), .B(n17819), .Z(n15828) );
  XOR2_X1 U18945 ( .A(n17390), .B(n15810), .Z(n15811) );
  NAND2_X1 U18946 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15811), .ZN(
        n15827) );
  XOR2_X1 U18947 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n15811), .Z(
        n17834) );
  XNOR2_X1 U18948 ( .A(n15813), .B(n15812), .ZN(n15814) );
  NAND2_X1 U18949 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n15814), .ZN(
        n15826) );
  XOR2_X1 U18950 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n15814), .Z(
        n17849) );
  XOR2_X1 U18951 ( .A(n15815), .B(n15817), .Z(n15816) );
  NAND2_X1 U18952 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15816), .ZN(
        n15825) );
  XOR2_X1 U18953 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n15816), .Z(
        n17862) );
  OAI21_X1 U18954 ( .B1(n15820), .B2(n15818), .A(n15817), .ZN(n15823) );
  NAND2_X1 U18955 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n15823), .ZN(
        n15824) );
  NOR2_X1 U18956 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n15819), .ZN(
        n15822) );
  INV_X1 U18957 ( .A(n17883), .ZN(n17885) );
  INV_X1 U18958 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18846) );
  NAND2_X1 U18959 ( .A1(n15820), .A2(n18846), .ZN(n17892) );
  NOR2_X1 U18960 ( .A1(n17885), .A2(n17892), .ZN(n17884) );
  NOR3_X1 U18961 ( .A1(n15822), .A2(n15821), .A3(n17884), .ZN(n17877) );
  XNOR2_X1 U18962 ( .A(n15756), .B(n15823), .ZN(n17876) );
  NAND2_X1 U18963 ( .A1(n17877), .A2(n17876), .ZN(n17875) );
  NAND2_X1 U18964 ( .A1(n15824), .A2(n17875), .ZN(n17861) );
  NAND2_X1 U18965 ( .A1(n17862), .A2(n17861), .ZN(n17860) );
  NAND2_X1 U18966 ( .A1(n15825), .A2(n17860), .ZN(n17848) );
  NAND2_X1 U18967 ( .A1(n17849), .A2(n17848), .ZN(n17847) );
  NAND2_X1 U18968 ( .A1(n15826), .A2(n17847), .ZN(n17833) );
  NAND2_X1 U18969 ( .A1(n17834), .A2(n17833), .ZN(n17832) );
  NAND2_X1 U18970 ( .A1(n15827), .A2(n17832), .ZN(n17818) );
  AOI222_X1 U18971 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15828), .B1(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17818), .C1(n15828), .C2(
        n17818), .ZN(n17805) );
  XNOR2_X1 U18972 ( .A(n17382), .B(n15829), .ZN(n17806) );
  NAND2_X1 U18973 ( .A1(n17805), .A2(n17806), .ZN(n17804) );
  NAND2_X1 U18974 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17804), .ZN(
        n15833) );
  NOR2_X1 U18975 ( .A1(n15830), .A2(n15833), .ZN(n15835) );
  INV_X1 U18976 ( .A(n15830), .ZN(n15834) );
  NOR2_X1 U18977 ( .A1(n17805), .A2(n17806), .ZN(n15832) );
  NOR2_X1 U18978 ( .A1(n15834), .A2(n15833), .ZN(n15831) );
  AOI211_X1 U18979 ( .C1(n15834), .C2(n15833), .A(n15832), .B(n15831), .ZN(
        n17796) );
  NOR2_X1 U18980 ( .A1(n17796), .A2(n18135), .ZN(n17795) );
  INV_X1 U18981 ( .A(n17744), .ZN(n18094) );
  NAND2_X1 U18982 ( .A1(n18094), .A2(n10173), .ZN(n18036) );
  NAND2_X1 U18983 ( .A1(n15837), .A2(n17964), .ZN(n17944) );
  NOR2_X1 U18984 ( .A1(n17581), .A2(n17944), .ZN(n17563) );
  NAND2_X1 U18985 ( .A1(n15838), .A2(n17563), .ZN(n15842) );
  NOR2_X1 U18986 ( .A1(n16427), .A2(n15842), .ZN(n16419) );
  NAND2_X1 U18987 ( .A1(n16392), .A2(n18205), .ZN(n18142) );
  NAND2_X1 U18988 ( .A1(n15836), .A2(n17760), .ZN(n17699) );
  NAND2_X1 U18989 ( .A1(n17707), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17706) );
  NOR2_X1 U18990 ( .A1(n17706), .A2(n18050), .ZN(n17602) );
  NAND2_X1 U18991 ( .A1(n17602), .A2(n15837), .ZN(n17943) );
  NOR2_X1 U18992 ( .A1(n17943), .A2(n17581), .ZN(n17564) );
  NAND2_X1 U18993 ( .A1(n17564), .A2(n15838), .ZN(n17910) );
  NOR2_X1 U18994 ( .A1(n17910), .A2(n16427), .ZN(n16406) );
  OAI22_X1 U18995 ( .A1(n18212), .A2(n16419), .B1(n18142), .B2(n16406), .ZN(
        n15839) );
  INV_X1 U18996 ( .A(n15839), .ZN(n15902) );
  OAI221_X1 U18997 ( .B1(n18218), .B2(n16448), .C1(n18218), .C2(n15840), .A(
        n15902), .ZN(n15841) );
  AOI22_X1 U18998 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15841), .B1(
        n18218), .B2(P3_REIP_REG_29__SCAN_IN), .ZN(n15850) );
  INV_X1 U18999 ( .A(n17910), .ZN(n17527) );
  INV_X1 U19000 ( .A(n18142), .ZN(n17937) );
  INV_X1 U19001 ( .A(n15842), .ZN(n17908) );
  INV_X1 U19002 ( .A(n18212), .ZN(n18217) );
  AOI22_X1 U19003 ( .A1(n17527), .A2(n17937), .B1(n17908), .B2(n18217), .ZN(
        n15848) );
  AOI22_X1 U19004 ( .A1(n18683), .A2(n15844), .B1(n18684), .B2(n15843), .ZN(
        n15846) );
  AOI221_X1 U19005 ( .B1(n15846), .B2(n15845), .C1(n15846), .C2(n18104), .A(
        n18207), .ZN(n15847) );
  INV_X1 U19006 ( .A(n15847), .ZN(n16425) );
  NAND2_X1 U19007 ( .A1(n15848), .A2(n16425), .ZN(n15904) );
  NAND3_X1 U19008 ( .A1(n16418), .A2(n16407), .A3(n15904), .ZN(n15849) );
  OAI211_X1 U19009 ( .C1(n16423), .C2(n18124), .A(n15850), .B(n15849), .ZN(
        P3_U2833) );
  INV_X1 U19010 ( .A(n15859), .ZN(n15861) );
  NOR3_X1 U19011 ( .A1(n15852), .A2(n15851), .A3(n20686), .ZN(n15855) );
  OAI22_X1 U19012 ( .A1(n15854), .A2(n15853), .B1(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n15855), .ZN(n15857) );
  NAND2_X1 U19013 ( .A1(n15855), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n15856) );
  OAI211_X1 U19014 ( .C1(n15859), .C2(n15858), .A(n15857), .B(n15856), .ZN(
        n15860) );
  OAI21_X1 U19015 ( .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15861), .A(
        n15860), .ZN(n15863) );
  AOI222_X1 U19016 ( .A1(n15863), .A2(n20634), .B1(n15863), .B2(n15862), .C1(
        n20634), .C2(n15862), .ZN(n15871) );
  INV_X1 U19017 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n21301) );
  AOI21_X1 U19018 ( .B1(n21022), .B2(n21301), .A(n15864), .ZN(n15866) );
  NOR4_X1 U19019 ( .A1(n15868), .A2(n15867), .A3(n15866), .A4(n15865), .ZN(
        n15869) );
  OAI211_X1 U19020 ( .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n15871), .A(
        n15870), .B(n15869), .ZN(n15878) );
  NOR2_X1 U19021 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20898), .ZN(n15876) );
  NOR2_X1 U19022 ( .A1(n15872), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20899) );
  NAND4_X1 U19023 ( .A1(n15874), .A2(n15873), .A3(n20899), .A4(n20906), .ZN(
        n15875) );
  OAI221_X1 U19024 ( .B1(n15879), .B2(n15876), .C1(n15879), .C2(n20835), .A(
        n15875), .ZN(n16190) );
  AOI221_X1 U19025 ( .B1(n20902), .B2(n16192), .C1(n15878), .C2(n16192), .A(
        n16190), .ZN(n15880) );
  NOR2_X1 U19026 ( .A1(n15880), .A2(n20902), .ZN(n20828) );
  OAI211_X1 U19027 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20906), .A(n20828), 
        .B(n15877), .ZN(n16191) );
  AOI21_X1 U19028 ( .B1(n15879), .B2(n15878), .A(n16191), .ZN(n15885) );
  INV_X1 U19029 ( .A(n15880), .ZN(n15881) );
  OAI21_X1 U19030 ( .B1(n15882), .B2(n20901), .A(n15881), .ZN(n15883) );
  AOI22_X1 U19031 ( .A1(n15885), .A2(n15884), .B1(n20902), .B2(n15883), .ZN(
        P1_U3161) );
  AOI22_X1 U19032 ( .A1(n15887), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n15886), .B2(n15892), .ZN(n15888) );
  XNOR2_X1 U19033 ( .A(n15888), .B(n15893), .ZN(n15995) );
  AOI22_X1 U19034 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n16064), .B1(
        n20150), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15895) );
  NAND2_X1 U19035 ( .A1(n9848), .A2(n15889), .ZN(n15890) );
  AND2_X1 U19036 ( .A1(n15926), .A2(n15890), .ZN(n15981) );
  NOR2_X1 U19037 ( .A1(n15892), .A2(n15891), .ZN(n16068) );
  AOI22_X1 U19038 ( .A1(n15981), .A2(n20214), .B1(n16068), .B2(n15893), .ZN(
        n15894) );
  OAI211_X1 U19039 ( .C1(n15995), .C2(n20196), .A(n15895), .B(n15894), .ZN(
        P1_U3010) );
  NAND2_X1 U19040 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15896), .ZN(
        n16379) );
  INV_X1 U19041 ( .A(n16379), .ZN(n15899) );
  NAND2_X1 U19042 ( .A1(n17540), .A2(n15897), .ZN(n15898) );
  NOR2_X1 U19043 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15898), .ZN(
        n16377) );
  NOR2_X1 U19044 ( .A1(n15899), .A2(n16377), .ZN(n15900) );
  XOR2_X1 U19045 ( .A(n15900), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16405) );
  NOR2_X1 U19046 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16427), .ZN(
        n16401) );
  INV_X1 U19047 ( .A(n18132), .ZN(n18131) );
  NOR2_X1 U19048 ( .A1(n18207), .A2(n18131), .ZN(n18170) );
  AOI22_X1 U19049 ( .A1(n18170), .A2(n16427), .B1(n18201), .B2(n15901), .ZN(
        n16424) );
  INV_X1 U19050 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16380) );
  AOI21_X1 U19051 ( .B1(n16424), .B2(n15902), .A(n16380), .ZN(n15903) );
  AOI21_X1 U19052 ( .B1(n16401), .B2(n15904), .A(n15903), .ZN(n15905) );
  NAND2_X1 U19053 ( .A1(n18218), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16397) );
  OAI211_X1 U19054 ( .C1(n16405), .C2(n18124), .A(n15905), .B(n16397), .ZN(
        P3_U2832) );
  INV_X1 U19055 ( .A(HOLD), .ZN(n21232) );
  NOR2_X1 U19056 ( .A1(n20843), .A2(n21232), .ZN(n20831) );
  AOI22_X1 U19057 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n15907) );
  NAND2_X1 U19058 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20835), .ZN(n20836) );
  OAI211_X1 U19059 ( .C1(n20831), .C2(n15907), .A(n15906), .B(n20836), .ZN(
        P1_U3195) );
  AND2_X1 U19060 ( .A1(n15908), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR3_X1 U19061 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n15909) );
  NOR3_X1 U19062 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n18909), .A3(n19835), 
        .ZN(n19821) );
  NOR4_X1 U19063 ( .A1(n15909), .A2(n16364), .A3(n16373), .A4(n19821), .ZN(
        P2_U3178) );
  AOI221_X1 U19064 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16373), .C1(n19972), .C2(
        n16373), .A(n19758), .ZN(n19965) );
  INV_X1 U19065 ( .A(n19965), .ZN(n19962) );
  NOR2_X1 U19066 ( .A1(n16340), .A2(n19962), .ZN(P2_U3047) );
  INV_X1 U19067 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n21170) );
  OAI21_X1 U19068 ( .B1(n11621), .B2(n15910), .A(n20904), .ZN(n15911) );
  OAI211_X1 U19069 ( .C1(n20904), .C2(n21170), .A(n19985), .B(n15911), .ZN(
        P1_U3487) );
  NOR3_X1 U19070 ( .A1(n15912), .A2(n17415), .A3(n16578), .ZN(n15913) );
  NAND2_X1 U19071 ( .A1(n18268), .A2(n17264), .ZN(n17311) );
  AOI22_X1 U19072 ( .A1(n17409), .A2(BUF2_REG_0__SCAN_IN), .B1(n17383), .B2(
        n15917), .ZN(n15918) );
  OAI221_X1 U19073 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17311), .C1(n10049), 
        .C2(n17264), .A(n15918), .ZN(P3_U2735) );
  NOR3_X1 U19074 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n20021), .A3(n15919), 
        .ZN(n15923) );
  INV_X1 U19075 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20950) );
  OAI21_X1 U19076 ( .B1(n15930), .B2(n20021), .A(n20059), .ZN(n15940) );
  AOI21_X1 U19077 ( .B1(n20069), .B2(n20950), .A(n15940), .ZN(n15921) );
  INV_X1 U19078 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n21260) );
  OAI22_X1 U19079 ( .A1(n15921), .A2(n15920), .B1(n21260), .B2(n20064), .ZN(
        n15922) );
  AOI211_X1 U19080 ( .C1(n20080), .C2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15923), .B(n15922), .ZN(n15928) );
  INV_X1 U19081 ( .A(n15924), .ZN(n15987) );
  XNOR2_X1 U19082 ( .A(n15926), .B(n15925), .ZN(n16065) );
  AOI22_X1 U19083 ( .A1(n15987), .A2(n20031), .B1(n20077), .B2(n16065), .ZN(
        n15927) );
  OAI211_X1 U19084 ( .C1(n15990), .C2(n20043), .A(n15928), .B(n15927), .ZN(
        P1_U2818) );
  AOI22_X1 U19085 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n20080), .B1(
        P1_EBX_REG_21__SCAN_IN), .B2(n20075), .ZN(n15934) );
  NOR2_X1 U19086 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n20021), .ZN(n15929) );
  AOI22_X1 U19087 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n15940), .B1(n15930), 
        .B2(n15929), .ZN(n15933) );
  AOI22_X1 U19088 ( .A1(n15992), .A2(n20031), .B1(n20077), .B2(n15981), .ZN(
        n15932) );
  NAND2_X1 U19089 ( .A1(n15991), .A2(n20079), .ZN(n15931) );
  NAND4_X1 U19090 ( .A1(n15934), .A2(n15933), .A3(n15932), .A4(n15931), .ZN(
        P1_U2819) );
  AOI22_X1 U19091 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n20080), .B1(
        P1_EBX_REG_20__SCAN_IN), .B2(n20075), .ZN(n15942) );
  OAI21_X1 U19092 ( .B1(n14512), .B2(n15935), .A(n21171), .ZN(n15939) );
  OAI22_X1 U19093 ( .A1(n15998), .A2(n15937), .B1(n15936), .B2(n20073), .ZN(
        n15938) );
  AOI21_X1 U19094 ( .B1(n15940), .B2(n15939), .A(n15938), .ZN(n15941) );
  OAI211_X1 U19095 ( .C1(n15996), .C2(n20043), .A(n15942), .B(n15941), .ZN(
        P1_U2820) );
  AOI21_X1 U19096 ( .B1(n20080), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20048), .ZN(n15943) );
  OAI21_X1 U19097 ( .B1(n20959), .B2(n20064), .A(n15943), .ZN(n15944) );
  AOI221_X1 U19098 ( .B1(n15947), .B2(P1_REIP_REG_18__SCAN_IN), .C1(n15946), 
        .C2(n15945), .A(n15944), .ZN(n15952) );
  INV_X1 U19099 ( .A(n15948), .ZN(n15949) );
  AOI22_X1 U19100 ( .A1(n15950), .A2(n20031), .B1(n15949), .B2(n20079), .ZN(
        n15951) );
  OAI211_X1 U19101 ( .C1(n20073), .C2(n16084), .A(n15952), .B(n15951), .ZN(
        P1_U2822) );
  OAI22_X1 U19102 ( .A1(n15954), .A2(n21014), .B1(n15953), .B2(n20064), .ZN(
        n15955) );
  AOI211_X1 U19103 ( .C1(n20080), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n20048), .B(n15955), .ZN(n15958) );
  OAI221_X1 U19104 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(P1_REIP_REG_15__SCAN_IN), .C1(n21014), .C2(n20988), .A(n15956), .ZN(n15957) );
  OAI211_X1 U19105 ( .C1(n16007), .C2(n20043), .A(n15958), .B(n15957), .ZN(
        n15959) );
  AOI21_X1 U19106 ( .B1(n16003), .B2(n20031), .A(n15959), .ZN(n15960) );
  OAI21_X1 U19107 ( .B1(n20073), .B2(n15961), .A(n15960), .ZN(P1_U2824) );
  OAI22_X1 U19108 ( .A1(n20972), .A2(n20064), .B1(n20073), .B2(n15962), .ZN(
        n15963) );
  AOI211_X1 U19109 ( .C1(n20080), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n20048), .B(n15963), .ZN(n15968) );
  INV_X1 U19110 ( .A(n15964), .ZN(n16019) );
  AOI22_X1 U19111 ( .A1(n16020), .A2(n20079), .B1(n20031), .B2(n16019), .ZN(
        n15967) );
  OAI221_X1 U19112 ( .B1(P1_REIP_REG_12__SCAN_IN), .B2(P1_REIP_REG_11__SCAN_IN), .C1(P1_REIP_REG_12__SCAN_IN), .C2(n15969), .A(n15965), .ZN(n15966) );
  NAND3_X1 U19113 ( .A1(n15968), .A2(n15967), .A3(n15966), .ZN(P1_U2828) );
  INV_X1 U19114 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n21195) );
  AOI22_X1 U19115 ( .A1(P1_EBX_REG_11__SCAN_IN), .A2(n20075), .B1(n15969), 
        .B2(n21195), .ZN(n15979) );
  INV_X1 U19116 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15976) );
  NAND2_X1 U19117 ( .A1(n15971), .A2(n15970), .ZN(n15972) );
  AND2_X1 U19118 ( .A1(n15973), .A2(n15972), .ZN(n16129) );
  AOI22_X1 U19119 ( .A1(n20077), .A2(n16129), .B1(P1_REIP_REG_11__SCAN_IN), 
        .B2(n15974), .ZN(n15975) );
  OAI21_X1 U19120 ( .B1(n15976), .B2(n20060), .A(n15975), .ZN(n15977) );
  AOI211_X1 U19121 ( .C1(n16029), .C2(n20031), .A(n20048), .B(n15977), .ZN(
        n15978) );
  OAI211_X1 U19122 ( .C1(n16032), .C2(n20043), .A(n15979), .B(n15978), .ZN(
        P1_U2829) );
  AOI22_X1 U19123 ( .A1(n15987), .A2(n20098), .B1(n20097), .B2(n16065), .ZN(
        n15980) );
  OAI21_X1 U19124 ( .B1(n20101), .B2(n21260), .A(n15980), .ZN(P1_U2850) );
  AOI22_X1 U19125 ( .A1(n15992), .A2(n20098), .B1(n20097), .B2(n15981), .ZN(
        n15982) );
  OAI21_X1 U19126 ( .B1(n20101), .B2(n14039), .A(n15982), .ZN(P1_U2851) );
  INV_X1 U19127 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n21184) );
  AOI22_X1 U19128 ( .A1(n16029), .A2(n20098), .B1(n20097), .B2(n16129), .ZN(
        n15983) );
  OAI21_X1 U19129 ( .B1(n20101), .B2(n21184), .A(n15983), .ZN(P1_U2861) );
  AOI22_X1 U19130 ( .A1(n20151), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n20150), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n15989) );
  NAND2_X1 U19131 ( .A1(n15985), .A2(n15984), .ZN(n15986) );
  XNOR2_X1 U19132 ( .A(n15986), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16066) );
  AOI22_X1 U19133 ( .A1(n15987), .A2(n20158), .B1(n16066), .B2(n20159), .ZN(
        n15988) );
  OAI211_X1 U19134 ( .C1(n20164), .C2(n15990), .A(n15989), .B(n15988), .ZN(
        P1_U2977) );
  AOI22_X1 U19135 ( .A1(n20151), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n20150), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15994) );
  AOI22_X1 U19136 ( .A1(n15992), .A2(n20158), .B1(n16037), .B2(n15991), .ZN(
        n15993) );
  OAI211_X1 U19137 ( .C1(n15995), .C2(n19988), .A(n15994), .B(n15993), .ZN(
        P1_U2978) );
  OAI22_X1 U19138 ( .A1(n15998), .A2(n15997), .B1(n15996), .B2(n20164), .ZN(
        n15999) );
  AOI211_X1 U19139 ( .C1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n20151), .A(
        n16000), .B(n15999), .ZN(n16001) );
  OAI21_X1 U19140 ( .B1(n16002), .B2(n19988), .A(n16001), .ZN(P1_U2979) );
  AOI22_X1 U19141 ( .A1(n20151), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n20150), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n16006) );
  AOI22_X1 U19142 ( .A1(n16004), .A2(n20159), .B1(n20158), .B2(n16003), .ZN(
        n16005) );
  OAI211_X1 U19143 ( .C1(n20164), .C2(n16007), .A(n16006), .B(n16005), .ZN(
        P1_U2983) );
  INV_X1 U19144 ( .A(n16008), .ZN(n16009) );
  AOI21_X1 U19145 ( .B1(n16011), .B2(n16010), .A(n16009), .ZN(n16014) );
  XNOR2_X1 U19146 ( .A(n16012), .B(n16110), .ZN(n16013) );
  XNOR2_X1 U19147 ( .A(n16014), .B(n16013), .ZN(n16112) );
  AOI22_X1 U19148 ( .A1(n20151), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20150), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16018) );
  AOI22_X1 U19149 ( .A1(n16016), .A2(n20158), .B1(n16037), .B2(n16015), .ZN(
        n16017) );
  OAI211_X1 U19150 ( .C1(n16112), .C2(n19988), .A(n16018), .B(n16017), .ZN(
        P1_U2985) );
  AOI22_X1 U19151 ( .A1(n20151), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20150), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16022) );
  AOI22_X1 U19152 ( .A1(n16037), .A2(n16020), .B1(n20158), .B2(n16019), .ZN(
        n16021) );
  OAI211_X1 U19153 ( .C1(n16023), .C2(n19988), .A(n16022), .B(n16021), .ZN(
        P1_U2987) );
  AOI22_X1 U19154 ( .A1(n20151), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20150), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16031) );
  OR3_X1 U19155 ( .A1(n16025), .A2(n16024), .A3(n14568), .ZN(n16026) );
  NAND2_X1 U19156 ( .A1(n16027), .A2(n16026), .ZN(n16028) );
  XOR2_X1 U19157 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n16028), .Z(
        n16132) );
  AOI22_X1 U19158 ( .A1(n20159), .A2(n16132), .B1(n20158), .B2(n16029), .ZN(
        n16030) );
  OAI211_X1 U19159 ( .C1(n20164), .C2(n16032), .A(n16031), .B(n16030), .ZN(
        P1_U2988) );
  INV_X1 U19160 ( .A(n16033), .ZN(n16034) );
  AOI21_X1 U19161 ( .B1(n16036), .B2(n16035), .A(n16034), .ZN(n16164) );
  INV_X1 U19162 ( .A(n16164), .ZN(n16039) );
  INV_X1 U19163 ( .A(n20025), .ZN(n16038) );
  AOI222_X1 U19164 ( .A1(n16039), .A2(n20159), .B1(n16038), .B2(n16037), .C1(
        n20158), .C2(n20094), .ZN(n16040) );
  NAND2_X1 U19165 ( .A1(n20150), .A2(P1_REIP_REG_7__SCAN_IN), .ZN(n16162) );
  OAI211_X1 U19166 ( .C1(n16042), .C2(n16041), .A(n16040), .B(n16162), .ZN(
        P1_U2992) );
  AOI22_X1 U19167 ( .A1(n20151), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20150), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16047) );
  INV_X1 U19168 ( .A(n16043), .ZN(n16045) );
  INV_X1 U19169 ( .A(n16044), .ZN(n20030) );
  AOI22_X1 U19170 ( .A1(n16045), .A2(n20159), .B1(n20158), .B2(n20030), .ZN(
        n16046) );
  OAI211_X1 U19171 ( .C1(n20164), .C2(n20035), .A(n16047), .B(n16046), .ZN(
        P1_U2993) );
  AOI22_X1 U19172 ( .A1(n20151), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20150), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n16054) );
  OAI21_X1 U19173 ( .B1(n16050), .B2(n16049), .A(n16048), .ZN(n16051) );
  INV_X1 U19174 ( .A(n16051), .ZN(n16176) );
  INV_X1 U19175 ( .A(n16052), .ZN(n20099) );
  AOI22_X1 U19176 ( .A1(n16176), .A2(n20159), .B1(n20158), .B2(n20099), .ZN(
        n16053) );
  OAI211_X1 U19177 ( .C1(n20164), .C2(n20044), .A(n16054), .B(n16053), .ZN(
        P1_U2994) );
  AOI22_X1 U19178 ( .A1(n20150), .A2(P1_REIP_REG_23__SCAN_IN), .B1(n16055), 
        .B2(n16091), .ZN(n16061) );
  INV_X1 U19179 ( .A(n16056), .ZN(n16059) );
  INV_X1 U19180 ( .A(n16057), .ZN(n16058) );
  AOI22_X1 U19181 ( .A1(n16059), .A2(n20208), .B1(n20214), .B2(n16058), .ZN(
        n16060) );
  OAI211_X1 U19182 ( .C1(n16063), .C2(n16062), .A(n16061), .B(n16060), .ZN(
        P1_U3008) );
  AOI22_X1 U19183 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n16064), .B1(
        n20150), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n16071) );
  AOI22_X1 U19184 ( .A1(n16066), .A2(n20208), .B1(n20214), .B2(n16065), .ZN(
        n16070) );
  OAI211_X1 U19185 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16068), .B(n16067), .ZN(
        n16069) );
  NAND3_X1 U19186 ( .A1(n16071), .A2(n16070), .A3(n16069), .ZN(P1_U3009) );
  INV_X1 U19187 ( .A(n16072), .ZN(n16074) );
  AOI22_X1 U19188 ( .A1(n16074), .A2(n20208), .B1(n20214), .B2(n16073), .ZN(
        n16081) );
  INV_X1 U19189 ( .A(n16075), .ZN(n16077) );
  NOR2_X1 U19190 ( .A1(n20207), .A2(n14512), .ZN(n16076) );
  AOI221_X1 U19191 ( .B1(n16079), .B2(n16078), .C1(n16077), .C2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n16076), .ZN(n16080) );
  NAND2_X1 U19192 ( .A1(n16081), .A2(n16080), .ZN(P1_U3012) );
  AOI21_X1 U19193 ( .B1(n20206), .B2(n16082), .A(n16122), .ZN(n16099) );
  NOR3_X1 U19194 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16083), .A3(
        n16082), .ZN(n16087) );
  OAI22_X1 U19195 ( .A1(n16085), .A2(n20196), .B1(n20171), .B2(n16084), .ZN(
        n16086) );
  AOI211_X1 U19196 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n20150), .A(n16087), 
        .B(n16086), .ZN(n16088) );
  OAI21_X1 U19197 ( .B1(n16099), .B2(n16089), .A(n16088), .ZN(P1_U3013) );
  NOR3_X1 U19198 ( .A1(n14418), .A2(n16110), .A3(n16090), .ZN(n16092) );
  AOI21_X1 U19199 ( .B1(n16092), .B2(n16091), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16098) );
  INV_X1 U19200 ( .A(n16093), .ZN(n16095) );
  AOI22_X1 U19201 ( .A1(n16095), .A2(n20208), .B1(n20214), .B2(n16094), .ZN(
        n16097) );
  NAND2_X1 U19202 ( .A1(n20150), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n16096) );
  OAI211_X1 U19203 ( .C1(n16099), .C2(n16098), .A(n16097), .B(n16096), .ZN(
        P1_U3014) );
  INV_X1 U19204 ( .A(n16100), .ZN(n16102) );
  AOI22_X1 U19205 ( .A1(n16102), .A2(n20208), .B1(n20214), .B2(n16101), .ZN(
        n16107) );
  NOR2_X1 U19206 ( .A1(n20207), .A2(n20988), .ZN(n16103) );
  AOI211_X1 U19207 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16105), .A(
        n16104), .B(n16103), .ZN(n16106) );
  NAND2_X1 U19208 ( .A1(n16107), .A2(n16106), .ZN(P1_U3016) );
  NAND3_X1 U19209 ( .A1(n16110), .A2(n16109), .A3(n16108), .ZN(n16116) );
  NOR2_X1 U19210 ( .A1(n20207), .A2(n21016), .ZN(n16114) );
  OAI22_X1 U19211 ( .A1(n16112), .A2(n20196), .B1(n20171), .B2(n16111), .ZN(
        n16113) );
  AOI211_X1 U19212 ( .C1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n16122), .A(
        n16114), .B(n16113), .ZN(n16115) );
  NAND2_X1 U19213 ( .A1(n16116), .A2(n16115), .ZN(P1_U3017) );
  INV_X1 U19214 ( .A(n16117), .ZN(n16119) );
  OAI221_X1 U19215 ( .B1(n16121), .B2(n16120), .C1(n16121), .C2(n16119), .A(
        n16118), .ZN(n16128) );
  AOI22_X1 U19216 ( .A1(n16123), .A2(n20208), .B1(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16122), .ZN(n16127) );
  NAND2_X1 U19217 ( .A1(n20150), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n16126) );
  NAND2_X1 U19218 ( .A1(n16124), .A2(n20214), .ZN(n16125) );
  NAND4_X1 U19219 ( .A1(n16128), .A2(n16127), .A3(n16126), .A4(n16125), .ZN(
        P1_U3018) );
  INV_X1 U19220 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16135) );
  AOI22_X1 U19221 ( .A1(n16129), .A2(n20214), .B1(n20150), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n16134) );
  NOR2_X1 U19222 ( .A1(n16130), .A2(n16163), .ZN(n16152) );
  NOR2_X1 U19223 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16144), .ZN(
        n16131) );
  AOI22_X1 U19224 ( .A1(n20208), .A2(n16132), .B1(n16152), .B2(n16131), .ZN(
        n16133) );
  OAI211_X1 U19225 ( .C1(n16136), .C2(n16135), .A(n16134), .B(n16133), .ZN(
        P1_U3020) );
  NOR2_X1 U19226 ( .A1(n20167), .A2(n16137), .ZN(n16139) );
  AOI211_X1 U19227 ( .C1(n20206), .C2(n16140), .A(n16139), .B(n16138), .ZN(
        n16157) );
  OAI22_X1 U19228 ( .A1(n16141), .A2(n20171), .B1(n21026), .B2(n20207), .ZN(
        n16142) );
  AOI21_X1 U19229 ( .B1(n20208), .B2(n16143), .A(n16142), .ZN(n16146) );
  OAI211_X1 U19230 ( .C1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n16152), .B(n16144), .ZN(n16145) );
  OAI211_X1 U19231 ( .C1(n16157), .C2(n14568), .A(n16146), .B(n16145), .ZN(
        P1_U3021) );
  AND2_X1 U19232 ( .A1(n16148), .A2(n16147), .ZN(n16149) );
  OR2_X1 U19233 ( .A1(n16150), .A2(n16149), .ZN(n20088) );
  INV_X1 U19234 ( .A(n20088), .ZN(n20008) );
  AOI21_X1 U19235 ( .B1(n20008), .B2(n20214), .A(n16151), .ZN(n16155) );
  AOI22_X1 U19236 ( .A1(n16153), .A2(n20208), .B1(n16152), .B2(n16156), .ZN(
        n16154) );
  OAI211_X1 U19237 ( .C1(n16157), .C2(n16156), .A(n16155), .B(n16154), .ZN(
        P1_U3022) );
  INV_X1 U19238 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16168) );
  OR2_X1 U19239 ( .A1(n16159), .A2(n16158), .ZN(n16160) );
  AND2_X1 U19240 ( .A1(n16161), .A2(n16160), .ZN(n20093) );
  OAI21_X1 U19241 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16163), .A(
        n16162), .ZN(n16166) );
  NOR2_X1 U19242 ( .A1(n16164), .A2(n20196), .ZN(n16165) );
  AOI211_X1 U19243 ( .C1(n20214), .C2(n20093), .A(n16166), .B(n16165), .ZN(
        n16167) );
  OAI21_X1 U19244 ( .B1(n16169), .B2(n16168), .A(n16167), .ZN(P1_U3024) );
  AND2_X1 U19245 ( .A1(n16171), .A2(n16170), .ZN(n16172) );
  NOR2_X1 U19246 ( .A1(n16173), .A2(n16172), .ZN(n20096) );
  AOI22_X1 U19247 ( .A1(n20096), .A2(n20214), .B1(n20150), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n16178) );
  INV_X1 U19248 ( .A(n16174), .ZN(n16175) );
  AOI22_X1 U19249 ( .A1(n16176), .A2(n20208), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n16175), .ZN(n16177) );
  OAI211_X1 U19250 ( .C1(n20183), .C2(n16179), .A(n16178), .B(n16177), .ZN(
        P1_U3026) );
  NAND3_X1 U19251 ( .A1(n16182), .A2(n16181), .A3(n16180), .ZN(n16183) );
  OAI21_X1 U19252 ( .B1(n16185), .B2(n16184), .A(n16183), .ZN(P1_U3468) );
  NAND4_X1 U19253 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20898), .A4(n20906), .ZN(n16186) );
  AND2_X1 U19254 ( .A1(n16187), .A2(n16186), .ZN(n20827) );
  NAND2_X1 U19255 ( .A1(n16188), .A2(n20827), .ZN(n16189) );
  AOI22_X1 U19256 ( .A1(n16192), .A2(n16191), .B1(n16190), .B2(n16189), .ZN(
        P1_U3162) );
  OAI21_X1 U19257 ( .B1(n20828), .B2(n20641), .A(n16193), .ZN(P1_U3466) );
  AOI211_X1 U19258 ( .C1(n16195), .C2(n16194), .A(n9904), .B(n19831), .ZN(
        n16203) );
  AOI22_X1 U19259 ( .A1(n19109), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n19089), .ZN(n16196) );
  OAI21_X1 U19260 ( .B1(n19122), .B2(n16197), .A(n16196), .ZN(n16198) );
  AOI21_X1 U19261 ( .B1(n16199), .B2(n19081), .A(n16198), .ZN(n16200) );
  OAI21_X1 U19262 ( .B1(n16201), .B2(n19115), .A(n16200), .ZN(n16202) );
  AOI211_X1 U19263 ( .C1(n19036), .C2(n16204), .A(n16203), .B(n16202), .ZN(
        n16205) );
  INV_X1 U19264 ( .A(n16205), .ZN(P2_U2827) );
  AOI22_X1 U19265 ( .A1(P2_REIP_REG_26__SCAN_IN), .A2(n19080), .B1(
        P2_EBX_REG_26__SCAN_IN), .B2(n19109), .ZN(n16220) );
  OAI22_X1 U19266 ( .A1(n16207), .A2(n19106), .B1(n19105), .B2(n16206), .ZN(
        n16208) );
  INV_X1 U19267 ( .A(n16208), .ZN(n16219) );
  INV_X1 U19268 ( .A(n16209), .ZN(n16210) );
  OAI22_X1 U19269 ( .A1(n16211), .A2(n19115), .B1(n16210), .B2(n19116), .ZN(
        n16212) );
  INV_X1 U19270 ( .A(n16212), .ZN(n16218) );
  AOI21_X1 U19271 ( .B1(n16215), .B2(n16214), .A(n16213), .ZN(n16216) );
  NAND2_X1 U19272 ( .A1(n19118), .A2(n16216), .ZN(n16217) );
  NAND4_X1 U19273 ( .A1(n16220), .A2(n16219), .A3(n16218), .A4(n16217), .ZN(
        P2_U2829) );
  OAI211_X1 U19274 ( .C1(n9911), .C2(n16222), .A(n19081), .B(n16221), .ZN(
        n16224) );
  AOI22_X1 U19275 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19089), .B1(
        P2_EBX_REG_25__SCAN_IN), .B2(n19109), .ZN(n16223) );
  OAI211_X1 U19276 ( .C1(n19122), .C2(n19903), .A(n16224), .B(n16223), .ZN(
        n16229) );
  AOI211_X1 U19277 ( .C1(n16227), .C2(n16226), .A(n16225), .B(n19831), .ZN(
        n16228) );
  AOI211_X1 U19278 ( .C1(n11089), .C2(n16230), .A(n16229), .B(n16228), .ZN(
        n16231) );
  OAI21_X1 U19279 ( .B1(n16232), .B2(n19116), .A(n16231), .ZN(P2_U2830) );
  AOI22_X1 U19280 ( .A1(n19127), .A2(n16233), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n19176), .ZN(n16238) );
  AOI22_X1 U19281 ( .A1(n19129), .A2(BUF1_REG_20__SCAN_IN), .B1(n19128), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n16237) );
  INV_X1 U19282 ( .A(n16234), .ZN(n18942) );
  AOI22_X1 U19283 ( .A1(n16235), .A2(n19137), .B1(n19177), .B2(n18942), .ZN(
        n16236) );
  NAND3_X1 U19284 ( .A1(n16238), .A2(n16237), .A3(n16236), .ZN(P2_U2899) );
  AOI22_X1 U19285 ( .A1(n19127), .A2(n16239), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n19176), .ZN(n16243) );
  AOI22_X1 U19286 ( .A1(n19129), .A2(BUF1_REG_18__SCAN_IN), .B1(n19128), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n16242) );
  AOI22_X1 U19287 ( .A1(n16240), .A2(n19137), .B1(n19177), .B2(n18967), .ZN(
        n16241) );
  NAND3_X1 U19288 ( .A1(n16243), .A2(n16242), .A3(n16241), .ZN(P2_U2901) );
  AOI22_X1 U19289 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19223), .B1(n19222), 
        .B2(n19000), .ZN(n16248) );
  AOI222_X1 U19290 ( .A1(n16246), .A2(n16282), .B1(n19231), .B2(n16245), .C1(
        n16283), .C2(n16244), .ZN(n16247) );
  OAI211_X1 U19291 ( .C1(n18995), .C2(n19234), .A(n16248), .B(n16247), .ZN(
        P2_U2999) );
  AOI22_X1 U19292 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19223), .B1(n19222), 
        .B2(n19022), .ZN(n16255) );
  NAND2_X1 U19293 ( .A1(n16249), .A2(n16283), .ZN(n16252) );
  NAND2_X1 U19294 ( .A1(n16250), .A2(n16282), .ZN(n16251) );
  OAI211_X1 U19295 ( .C1(n13154), .C2(n19024), .A(n16252), .B(n16251), .ZN(
        n16253) );
  INV_X1 U19296 ( .A(n16253), .ZN(n16254) );
  OAI211_X1 U19297 ( .C1(n19017), .C2(n19234), .A(n16255), .B(n16254), .ZN(
        P2_U3001) );
  AOI22_X1 U19298 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19223), .B1(n19222), 
        .B2(n19047), .ZN(n16262) );
  OR2_X1 U19299 ( .A1(n16256), .A2(n19225), .ZN(n16259) );
  NAND2_X1 U19300 ( .A1(n16257), .A2(n16282), .ZN(n16258) );
  OAI211_X1 U19301 ( .C1(n13154), .C2(n19049), .A(n16259), .B(n16258), .ZN(
        n16260) );
  INV_X1 U19302 ( .A(n16260), .ZN(n16261) );
  OAI211_X1 U19303 ( .C1(n19042), .C2(n19234), .A(n16262), .B(n16261), .ZN(
        P2_U3003) );
  AOI22_X1 U19304 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19223), .B1(n19222), 
        .B2(n16263), .ZN(n16271) );
  NAND2_X1 U19305 ( .A1(n16264), .A2(n16282), .ZN(n16267) );
  NAND2_X1 U19306 ( .A1(n16265), .A2(n19231), .ZN(n16266) );
  OAI211_X1 U19307 ( .C1(n16268), .C2(n19225), .A(n16267), .B(n16266), .ZN(
        n16269) );
  INV_X1 U19308 ( .A(n16269), .ZN(n16270) );
  OAI211_X1 U19309 ( .C1(n16272), .C2(n19234), .A(n16271), .B(n16270), .ZN(
        P2_U3005) );
  AOI22_X1 U19310 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19223), .B1(n19222), 
        .B2(n19067), .ZN(n16287) );
  INV_X1 U19311 ( .A(n19072), .ZN(n16303) );
  XOR2_X1 U19312 ( .A(n16273), .B(n16274), .Z(n16302) );
  AOI21_X1 U19313 ( .B1(n15208), .B2(n16276), .A(n16275), .ZN(n16281) );
  INV_X1 U19314 ( .A(n16277), .ZN(n16278) );
  NOR2_X1 U19315 ( .A1(n16279), .A2(n16278), .ZN(n16280) );
  XNOR2_X1 U19316 ( .A(n16281), .B(n16280), .ZN(n16305) );
  AOI22_X1 U19317 ( .A1(n16302), .A2(n16283), .B1(n16282), .B2(n16305), .ZN(
        n16284) );
  INV_X1 U19318 ( .A(n16284), .ZN(n16285) );
  AOI21_X1 U19319 ( .B1(n19231), .B2(n16303), .A(n16285), .ZN(n16286) );
  OAI211_X1 U19320 ( .C1(n16288), .C2(n19234), .A(n16287), .B(n16286), .ZN(
        P2_U3006) );
  AOI22_X1 U19321 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n19223), .B1(n19222), 
        .B2(n19099), .ZN(n16294) );
  INV_X1 U19322 ( .A(n16289), .ZN(n16291) );
  OAI22_X1 U19323 ( .A1(n16291), .A2(n19227), .B1(n16290), .B2(n19225), .ZN(
        n16292) );
  AOI21_X1 U19324 ( .B1(n19231), .B2(n19100), .A(n16292), .ZN(n16293) );
  OAI211_X1 U19325 ( .C1(n16295), .C2(n19234), .A(n16294), .B(n16293), .ZN(
        P2_U3008) );
  AOI21_X1 U19326 ( .B1(n16298), .B2(n16297), .A(n16296), .ZN(n19071) );
  AOI22_X1 U19327 ( .A1(n16300), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n16299), .B2(n19071), .ZN(n16311) );
  AOI222_X1 U19328 ( .A1(n16305), .A2(n16322), .B1(n16304), .B2(n16303), .C1(
        n16302), .C2(n16301), .ZN(n16310) );
  NAND2_X1 U19329 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19223), .ZN(n16309) );
  OAI211_X1 U19330 ( .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n16307), .B(n16306), .ZN(n16308) );
  NAND4_X1 U19331 ( .A1(n16311), .A2(n16310), .A3(n16309), .A4(n16308), .ZN(
        P2_U3038) );
  OAI22_X1 U19332 ( .A1(n16315), .A2(n16314), .B1(n16313), .B2(n16312), .ZN(
        n16320) );
  INV_X1 U19333 ( .A(n16316), .ZN(n16317) );
  MUX2_X1 U19334 ( .A(n16318), .B(n16317), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n16319) );
  AOI211_X1 U19335 ( .C1(n16322), .C2(n16321), .A(n16320), .B(n16319), .ZN(
        n16324) );
  OAI211_X1 U19336 ( .C1(n16326), .C2(n16325), .A(n16324), .B(n16323), .ZN(
        P2_U3046) );
  MUX2_X1 U19337 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16327), .S(
        n16330), .Z(n16336) );
  INV_X1 U19338 ( .A(n16336), .ZN(n16360) );
  MUX2_X1 U19339 ( .A(n16329), .B(n16328), .S(n16330), .Z(n16359) );
  INV_X1 U19340 ( .A(n16330), .ZN(n16356) );
  INV_X1 U19341 ( .A(n16332), .ZN(n16334) );
  AOI22_X1 U19342 ( .A1(n16332), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n16331), .ZN(n16333) );
  AOI21_X1 U19343 ( .B1(n19955), .B2(n16334), .A(n16333), .ZN(n16335) );
  AOI211_X1 U19344 ( .C1(n16359), .C2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n16356), .B(n16335), .ZN(n16338) );
  NOR2_X1 U19345 ( .A1(n16359), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n16337) );
  OAI22_X1 U19346 ( .A1(n16338), .A2(n16337), .B1(n19935), .B2(n16336), .ZN(
        n16339) );
  OAI21_X1 U19347 ( .B1(n16360), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n16339), .ZN(n16341) );
  NAND2_X1 U19348 ( .A1(n16341), .A2(n16340), .ZN(n16358) );
  OAI21_X1 U19349 ( .B1(P2_MORE_REG_SCAN_IN), .B2(P2_FLUSH_REG_SCAN_IN), .A(
        n16342), .ZN(n16345) );
  OR3_X1 U19350 ( .A1(n15657), .A2(n16343), .A3(n11433), .ZN(n16344) );
  OAI211_X1 U19351 ( .C1(n16347), .C2(n16346), .A(n16345), .B(n16344), .ZN(
        n16355) );
  INV_X1 U19352 ( .A(n16348), .ZN(n16349) );
  AOI22_X1 U19353 ( .A1(n16354), .A2(n16351), .B1(n16350), .B2(n16349), .ZN(
        n16352) );
  OAI21_X1 U19354 ( .B1(n16354), .B2(n16353), .A(n16352), .ZN(n19973) );
  AOI211_X1 U19355 ( .C1(n16356), .C2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n16355), .B(n19973), .ZN(n16357) );
  OAI211_X1 U19356 ( .C1(n16360), .C2(n16359), .A(n16358), .B(n16357), .ZN(
        n16366) );
  AOI211_X1 U19357 ( .C1(n16362), .C2(n16366), .A(n16361), .B(n19821), .ZN(
        n16371) );
  AND3_X1 U19358 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n16363), .A3(n19851), 
        .ZN(n19823) );
  AOI21_X1 U19359 ( .B1(n16365), .B2(n16364), .A(n19823), .ZN(n16369) );
  OAI21_X1 U19360 ( .B1(n16366), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n19822) );
  NAND2_X1 U19361 ( .A1(n10914), .A2(n16367), .ZN(n16368) );
  NAND3_X1 U19362 ( .A1(n19822), .A2(n16368), .A3(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19828) );
  NAND2_X1 U19363 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19828), .ZN(n16374) );
  OAI21_X1 U19364 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16369), .A(n16374), 
        .ZN(n16370) );
  OAI211_X1 U19365 ( .C1(n19972), .C2(n16372), .A(n16371), .B(n16370), .ZN(
        P2_U3176) );
  AOI21_X1 U19366 ( .B1(n16374), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n16373), 
        .ZN(n16375) );
  INV_X1 U19367 ( .A(n16375), .ZN(P2_U3593) );
  OAI22_X2 U19368 ( .A1(n16376), .A2(n18677), .B1(n18674), .B2(n16441), .ZN(
        n18722) );
  NOR2_X1 U19369 ( .A1(n17798), .A2(n16377), .ZN(n16386) );
  OAI21_X1 U19370 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n17798), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16378) );
  OAI221_X1 U19371 ( .B1(n16380), .B2(n16379), .C1(n17798), .C2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A(n16378), .ZN(n16385) );
  INV_X1 U19372 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18844) );
  NAND2_X1 U19373 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18844), .ZN(
        n16426) );
  NAND2_X1 U19374 ( .A1(n16426), .A2(n16379), .ZN(n16383) );
  NAND2_X1 U19375 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17798), .ZN(
        n16381) );
  OAI22_X1 U19376 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17798), .B1(
        n16381), .B2(n16380), .ZN(n16382) );
  OAI21_X1 U19377 ( .B1(n16386), .B2(n16383), .A(n16382), .ZN(n16384) );
  OAI21_X1 U19378 ( .B1(n16386), .B2(n16385), .A(n16384), .ZN(n16435) );
  INV_X1 U19379 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16611) );
  NAND2_X1 U19380 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17845) );
  INV_X1 U19381 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17859) );
  NAND3_X1 U19382 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16812) );
  NAND2_X1 U19383 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17725) );
  NAND2_X1 U19384 ( .A1(n16779), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17685) );
  NAND2_X1 U19385 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17686) );
  NAND2_X1 U19386 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n17668), .ZN(
        n17645) );
  NAND2_X1 U19387 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17647) );
  NAND2_X1 U19388 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17612) );
  NAND2_X1 U19389 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17570) );
  NAND2_X1 U19390 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17535) );
  INV_X1 U19391 ( .A(n16388), .ZN(n16413) );
  INV_X1 U19392 ( .A(n16581), .ZN(n16409) );
  INV_X1 U19393 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18820) );
  NOR2_X1 U19394 ( .A1(n18820), .A2(n18201), .ZN(n16429) );
  NAND2_X1 U19395 ( .A1(n16388), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16389) );
  NAND2_X1 U19396 ( .A1(n18735), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17895) );
  OAI21_X1 U19397 ( .B1(n17890), .B2(n17633), .A(n18575), .ZN(n17684) );
  INV_X1 U19398 ( .A(n17684), .ZN(n17646) );
  OR2_X1 U19399 ( .A1(n16389), .A2(n17646), .ZN(n16399) );
  XNOR2_X1 U19400 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16390) );
  NOR2_X1 U19401 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17633), .ZN(
        n16410) );
  NAND2_X1 U19402 ( .A1(n18616), .A2(n16389), .ZN(n16414) );
  OAI211_X1 U19403 ( .C1(n16581), .C2(n17895), .A(n17894), .B(n16414), .ZN(
        n16417) );
  NOR2_X1 U19404 ( .A1(n16410), .A2(n16417), .ZN(n16398) );
  OAI22_X1 U19405 ( .A1(n16399), .A2(n16390), .B1(n16398), .B2(n10123), .ZN(
        n16391) );
  AOI211_X1 U19406 ( .C1(n17735), .C2(n16878), .A(n16429), .B(n16391), .ZN(
        n16396) );
  NAND2_X1 U19407 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16406), .ZN(
        n16393) );
  XOR2_X1 U19408 ( .A(n16393), .B(n18844), .Z(n16431) );
  NOR2_X1 U19409 ( .A1(n16578), .A2(n16558), .ZN(n17800) );
  NAND2_X1 U19410 ( .A1(n16419), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16394) );
  XOR2_X1 U19411 ( .A(n16394), .B(n18844), .Z(n16432) );
  AOI22_X1 U19412 ( .A1(n17745), .A2(n16431), .B1(n17800), .B2(n16432), .ZN(
        n16395) );
  OAI211_X1 U19413 ( .C1(n17773), .C2(n16435), .A(n16396), .B(n16395), .ZN(
        P3_U2799) );
  XNOR2_X1 U19414 ( .A(n10122), .B(n16408), .ZN(n16602) );
  OAI221_X1 U19415 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16399), .C1(
        n10122), .C2(n16398), .A(n16397), .ZN(n16400) );
  AOI21_X1 U19416 ( .B1(n17735), .B2(n16602), .A(n16400), .ZN(n16404) );
  OAI22_X1 U19417 ( .A1(n16406), .A2(n17803), .B1(n16419), .B2(n17899), .ZN(
        n16402) );
  OAI22_X1 U19418 ( .A1(n17744), .A2(n17899), .B1(n17803), .B2(n18099), .ZN(
        n17746) );
  NAND2_X1 U19419 ( .A1(n10173), .A2(n17746), .ZN(n17693) );
  NAND2_X1 U19420 ( .A1(n17927), .A2(n17610), .ZN(n17596) );
  NOR2_X1 U19421 ( .A1(n17903), .A2(n17596), .ZN(n17548) );
  AOI22_X1 U19422 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16402), .B1(
        n16401), .B2(n17548), .ZN(n16403) );
  OAI211_X1 U19423 ( .C1(n16405), .C2(n17773), .A(n16404), .B(n16403), .ZN(
        P3_U2800) );
  NAND2_X1 U19424 ( .A1(n17527), .A2(n16418), .ZN(n16444) );
  AOI211_X1 U19425 ( .C1(n16407), .C2(n16444), .A(n16406), .B(n17803), .ZN(
        n16416) );
  NAND2_X1 U19426 ( .A1(n18218), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16412) );
  AOI21_X1 U19427 ( .B1(n16611), .B2(n16409), .A(n16408), .ZN(n16610) );
  OAI21_X1 U19428 ( .B1(n16410), .B2(n17735), .A(n16610), .ZN(n16411) );
  OAI211_X1 U19429 ( .C1(n16414), .C2(n16413), .A(n16412), .B(n16411), .ZN(
        n16415) );
  AOI211_X1 U19430 ( .C1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n16417), .A(
        n16416), .B(n16415), .ZN(n16422) );
  AND2_X1 U19431 ( .A1(n16418), .A2(n17908), .ZN(n16442) );
  INV_X1 U19432 ( .A(n16419), .ZN(n16420) );
  OAI211_X1 U19433 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16442), .A(
        n17800), .B(n16420), .ZN(n16421) );
  OAI211_X1 U19434 ( .C1(n16423), .C2(n17773), .A(n16422), .B(n16421), .ZN(
        P3_U2801) );
  INV_X1 U19435 ( .A(n18170), .ZN(n18202) );
  OAI21_X1 U19436 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18202), .A(
        n16424), .ZN(n16430) );
  NOR3_X1 U19437 ( .A1(n16427), .A2(n16426), .A3(n16425), .ZN(n16428) );
  AOI211_X1 U19438 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n16430), .A(
        n16429), .B(n16428), .ZN(n16434) );
  AOI22_X1 U19439 ( .A1(n18217), .A2(n16432), .B1(n17937), .B2(n16431), .ZN(
        n16433) );
  OAI211_X1 U19440 ( .C1(n16435), .C2(n18124), .A(n16434), .B(n16433), .ZN(
        P3_U2831) );
  NAND4_X1 U19441 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17798), .A3(
        n16436), .A4(n17528), .ZN(n16460) );
  INV_X1 U19442 ( .A(n18205), .ZN(n18222) );
  NAND2_X1 U19443 ( .A1(n16438), .A2(n16437), .ZN(n17531) );
  INV_X1 U19444 ( .A(n17918), .ZN(n16439) );
  OAI21_X1 U19445 ( .B1(n16440), .B2(n17541), .A(n16439), .ZN(n16446) );
  NOR2_X1 U19446 ( .A1(n17382), .A2(n16441), .ZN(n18100) );
  NOR2_X1 U19447 ( .A1(n17990), .A2(n17528), .ZN(n16456) );
  NOR2_X1 U19448 ( .A1(n18013), .A2(n16450), .ZN(n17656) );
  INV_X1 U19449 ( .A(n18100), .ZN(n18076) );
  OAI22_X1 U19450 ( .A1(n17744), .A2(n18677), .B1(n18099), .B2(n18076), .ZN(
        n18008) );
  OAI21_X1 U19451 ( .B1(n18846), .B2(n18104), .A(n18696), .ZN(n18006) );
  AOI22_X1 U19452 ( .A1(n18684), .A2(n18011), .B1(n16451), .B2(n18006), .ZN(
        n16452) );
  INV_X1 U19453 ( .A(n16452), .ZN(n17926) );
  AOI21_X1 U19454 ( .B1(n17656), .B2(n18008), .A(n17926), .ZN(n17902) );
  NOR2_X1 U19455 ( .A1(n17902), .A2(n18207), .ZN(n17981) );
  NOR4_X1 U19456 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n15781), .A3(
        n17901), .A4(n17903), .ZN(n17533) );
  NAND2_X1 U19457 ( .A1(n18218), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17537) );
  INV_X1 U19458 ( .A(n17537), .ZN(n16453) );
  NAND3_X1 U19459 ( .A1(n18138), .A2(n17540), .A3(n17531), .ZN(n16458) );
  OAI211_X1 U19460 ( .C1(n16460), .C2(n18222), .A(n16459), .B(n16458), .ZN(
        P3_U2834) );
  NOR3_X1 U19461 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16462) );
  NOR4_X1 U19462 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16461) );
  INV_X2 U19463 ( .A(n16544), .ZN(U215) );
  NAND4_X1 U19464 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16462), .A3(n16461), .A4(
        U215), .ZN(U213) );
  INV_X1 U19465 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16546) );
  INV_X2 U19466 ( .A(U214), .ZN(n16507) );
  INV_X1 U19467 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16547) );
  OAI222_X1 U19468 ( .A1(U212), .A2(n16546), .B1(n16509), .B2(n20284), .C1(
        U214), .C2(n16547), .ZN(U216) );
  INV_X2 U19469 ( .A(U212), .ZN(n16506) );
  AOI22_X1 U19470 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16506), .ZN(n16464) );
  OAI21_X1 U19471 ( .B1(n20277), .B2(n16509), .A(n16464), .ZN(U217) );
  INV_X1 U19472 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20270) );
  AOI22_X1 U19473 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16506), .ZN(n16465) );
  OAI21_X1 U19474 ( .B1(n20270), .B2(n16509), .A(n16465), .ZN(U218) );
  AOI22_X1 U19475 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16506), .ZN(n16466) );
  OAI21_X1 U19476 ( .B1(n14335), .B2(n16509), .A(n16466), .ZN(U219) );
  INV_X1 U19477 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20255) );
  AOI22_X1 U19478 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16506), .ZN(n16467) );
  OAI21_X1 U19479 ( .B1(n20255), .B2(n16509), .A(n16467), .ZN(U220) );
  INV_X1 U19480 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20247) );
  AOI22_X1 U19481 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16506), .ZN(n16468) );
  OAI21_X1 U19482 ( .B1(n20247), .B2(n16509), .A(n16468), .ZN(U221) );
  INV_X1 U19483 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20240) );
  AOI22_X1 U19484 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16506), .ZN(n16469) );
  OAI21_X1 U19485 ( .B1(n20240), .B2(n16509), .A(n16469), .ZN(U222) );
  INV_X1 U19486 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20229) );
  AOI22_X1 U19487 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16506), .ZN(n16470) );
  OAI21_X1 U19488 ( .B1(n20229), .B2(n16509), .A(n16470), .ZN(U223) );
  AOI22_X1 U19489 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16506), .ZN(n16471) );
  OAI21_X1 U19490 ( .B1(n14966), .B2(n16509), .A(n16471), .ZN(U224) );
  AOI22_X1 U19491 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16506), .ZN(n16472) );
  OAI21_X1 U19492 ( .B1(n20280), .B2(n16509), .A(n16472), .ZN(U225) );
  AOI22_X1 U19493 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16506), .ZN(n16473) );
  OAI21_X1 U19494 ( .B1(n20273), .B2(n16509), .A(n16473), .ZN(U226) );
  INV_X1 U19495 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n20266) );
  AOI22_X1 U19496 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16506), .ZN(n16474) );
  OAI21_X1 U19497 ( .B1(n20266), .B2(n16509), .A(n16474), .ZN(U227) );
  INV_X1 U19498 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20258) );
  AOI22_X1 U19499 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16506), .ZN(n16475) );
  OAI21_X1 U19500 ( .B1(n20258), .B2(n16509), .A(n16475), .ZN(U228) );
  INV_X1 U19501 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20251) );
  AOI22_X1 U19502 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16506), .ZN(n16476) );
  OAI21_X1 U19503 ( .B1(n20251), .B2(n16509), .A(n16476), .ZN(U229) );
  INV_X1 U19504 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20243) );
  AOI22_X1 U19505 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16506), .ZN(n16477) );
  OAI21_X1 U19506 ( .B1(n20243), .B2(n16509), .A(n16477), .ZN(U230) );
  INV_X1 U19507 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20236) );
  AOI22_X1 U19508 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16506), .ZN(n16478) );
  OAI21_X1 U19509 ( .B1(n20236), .B2(n16509), .A(n16478), .ZN(U231) );
  INV_X1 U19510 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n16480) );
  AOI22_X1 U19511 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16506), .ZN(n16479) );
  OAI21_X1 U19512 ( .B1(n16480), .B2(n16509), .A(n16479), .ZN(U232) );
  INV_X1 U19513 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n16482) );
  AOI22_X1 U19514 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16506), .ZN(n16481) );
  OAI21_X1 U19515 ( .B1(n16482), .B2(n16509), .A(n16481), .ZN(U233) );
  AOI22_X1 U19516 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16506), .ZN(n16483) );
  OAI21_X1 U19517 ( .B1(n16484), .B2(n16509), .A(n16483), .ZN(U234) );
  INV_X1 U19518 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16486) );
  AOI22_X1 U19519 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16506), .ZN(n16485) );
  OAI21_X1 U19520 ( .B1(n16486), .B2(n16509), .A(n16485), .ZN(U235) );
  AOI22_X1 U19521 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16506), .ZN(n16487) );
  OAI21_X1 U19522 ( .B1(n12543), .B2(n16509), .A(n16487), .ZN(U236) );
  INV_X1 U19523 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16489) );
  AOI22_X1 U19524 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16506), .ZN(n16488) );
  OAI21_X1 U19525 ( .B1(n16489), .B2(n16509), .A(n16488), .ZN(U237) );
  AOI22_X1 U19526 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16506), .ZN(n16490) );
  OAI21_X1 U19527 ( .B1(n12517), .B2(n16509), .A(n16490), .ZN(U238) );
  INV_X1 U19528 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16492) );
  AOI22_X1 U19529 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16506), .ZN(n16491) );
  OAI21_X1 U19530 ( .B1(n16492), .B2(n16509), .A(n16491), .ZN(U239) );
  AOI22_X1 U19531 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16506), .ZN(n16493) );
  OAI21_X1 U19532 ( .B1(n12534), .B2(n16509), .A(n16493), .ZN(U240) );
  INV_X1 U19533 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16495) );
  AOI22_X1 U19534 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16506), .ZN(n16494) );
  OAI21_X1 U19535 ( .B1(n16495), .B2(n16509), .A(n16494), .ZN(U241) );
  AOI22_X1 U19536 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16506), .ZN(n16496) );
  OAI21_X1 U19537 ( .B1(n16497), .B2(n16509), .A(n16496), .ZN(U242) );
  INV_X1 U19538 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16499) );
  AOI22_X1 U19539 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16506), .ZN(n16498) );
  OAI21_X1 U19540 ( .B1(n16499), .B2(n16509), .A(n16498), .ZN(U243) );
  INV_X1 U19541 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16501) );
  AOI22_X1 U19542 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16506), .ZN(n16500) );
  OAI21_X1 U19543 ( .B1(n16501), .B2(n16509), .A(n16500), .ZN(U244) );
  INV_X1 U19544 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16503) );
  AOI22_X1 U19545 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16506), .ZN(n16502) );
  OAI21_X1 U19546 ( .B1(n16503), .B2(n16509), .A(n16502), .ZN(U245) );
  INV_X1 U19547 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16505) );
  AOI22_X1 U19548 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16506), .ZN(n16504) );
  OAI21_X1 U19549 ( .B1(n16505), .B2(n16509), .A(n16504), .ZN(U246) );
  INV_X1 U19550 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16510) );
  AOI22_X1 U19551 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16506), .ZN(n16508) );
  OAI21_X1 U19552 ( .B1(n16510), .B2(n16509), .A(n16508), .ZN(U247) );
  OAI22_X1 U19553 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16544), .ZN(n16511) );
  INV_X1 U19554 ( .A(n16511), .ZN(U251) );
  OAI22_X1 U19555 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16544), .ZN(n16512) );
  INV_X1 U19556 ( .A(n16512), .ZN(U252) );
  OAI22_X1 U19557 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16544), .ZN(n16513) );
  INV_X1 U19558 ( .A(n16513), .ZN(U253) );
  OAI22_X1 U19559 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16544), .ZN(n16514) );
  INV_X1 U19560 ( .A(n16514), .ZN(U254) );
  OAI22_X1 U19561 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16544), .ZN(n16515) );
  INV_X1 U19562 ( .A(n16515), .ZN(U255) );
  OAI22_X1 U19563 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16544), .ZN(n16516) );
  INV_X1 U19564 ( .A(n16516), .ZN(U256) );
  OAI22_X1 U19565 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16544), .ZN(n16517) );
  INV_X1 U19566 ( .A(n16517), .ZN(U257) );
  OAI22_X1 U19567 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16544), .ZN(n16518) );
  INV_X1 U19568 ( .A(n16518), .ZN(U258) );
  OAI22_X1 U19569 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16544), .ZN(n16519) );
  INV_X1 U19570 ( .A(n16519), .ZN(U259) );
  OAI22_X1 U19571 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16538), .ZN(n16520) );
  INV_X1 U19572 ( .A(n16520), .ZN(U260) );
  OAI22_X1 U19573 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16538), .ZN(n16521) );
  INV_X1 U19574 ( .A(n16521), .ZN(U261) );
  OAI22_X1 U19575 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16544), .ZN(n16522) );
  INV_X1 U19576 ( .A(n16522), .ZN(U262) );
  OAI22_X1 U19577 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16544), .ZN(n16523) );
  INV_X1 U19578 ( .A(n16523), .ZN(U263) );
  OAI22_X1 U19579 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16544), .ZN(n16524) );
  INV_X1 U19580 ( .A(n16524), .ZN(U264) );
  OAI22_X1 U19581 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16544), .ZN(n16525) );
  INV_X1 U19582 ( .A(n16525), .ZN(U265) );
  OAI22_X1 U19583 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16538), .ZN(n16526) );
  INV_X1 U19584 ( .A(n16526), .ZN(U266) );
  OAI22_X1 U19585 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16538), .ZN(n16527) );
  INV_X1 U19586 ( .A(n16527), .ZN(U267) );
  OAI22_X1 U19587 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16538), .ZN(n16528) );
  INV_X1 U19588 ( .A(n16528), .ZN(U268) );
  OAI22_X1 U19589 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16538), .ZN(n16529) );
  INV_X1 U19590 ( .A(n16529), .ZN(U269) );
  OAI22_X1 U19591 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16538), .ZN(n16530) );
  INV_X1 U19592 ( .A(n16530), .ZN(U270) );
  OAI22_X1 U19593 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16538), .ZN(n16531) );
  INV_X1 U19594 ( .A(n16531), .ZN(U271) );
  OAI22_X1 U19595 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16544), .ZN(n16532) );
  INV_X1 U19596 ( .A(n16532), .ZN(U272) );
  OAI22_X1 U19597 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16544), .ZN(n16533) );
  INV_X1 U19598 ( .A(n16533), .ZN(U273) );
  OAI22_X1 U19599 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16538), .ZN(n16534) );
  INV_X1 U19600 ( .A(n16534), .ZN(U274) );
  OAI22_X1 U19601 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16544), .ZN(n16535) );
  INV_X1 U19602 ( .A(n16535), .ZN(U275) );
  OAI22_X1 U19603 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16544), .ZN(n16536) );
  INV_X1 U19604 ( .A(n16536), .ZN(U276) );
  OAI22_X1 U19605 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16544), .ZN(n16537) );
  INV_X1 U19606 ( .A(n16537), .ZN(U277) );
  OAI22_X1 U19607 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16538), .ZN(n16539) );
  INV_X1 U19608 ( .A(n16539), .ZN(U278) );
  OAI22_X1 U19609 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16544), .ZN(n16540) );
  INV_X1 U19610 ( .A(n16540), .ZN(U279) );
  OAI22_X1 U19611 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16544), .ZN(n16541) );
  INV_X1 U19612 ( .A(n16541), .ZN(U280) );
  OAI22_X1 U19613 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16544), .ZN(n16543) );
  INV_X1 U19614 ( .A(n16543), .ZN(U281) );
  INV_X1 U19615 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n17270) );
  AOI22_X1 U19616 ( .A1(n16544), .A2(n16546), .B1(n17270), .B2(U215), .ZN(U282) );
  INV_X1 U19617 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16545) );
  AOI222_X1 U19618 ( .A1(n16547), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16546), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16545), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16548) );
  INV_X2 U19619 ( .A(n16550), .ZN(n16549) );
  INV_X1 U19620 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18780) );
  INV_X1 U19621 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19874) );
  AOI22_X1 U19622 ( .A1(n16549), .A2(n18780), .B1(n19874), .B2(n16550), .ZN(
        U347) );
  INV_X1 U19623 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18778) );
  INV_X1 U19624 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19872) );
  AOI22_X1 U19625 ( .A1(n16549), .A2(n18778), .B1(n19872), .B2(n16550), .ZN(
        U348) );
  INV_X1 U19626 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18775) );
  INV_X1 U19627 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19871) );
  AOI22_X1 U19628 ( .A1(n16549), .A2(n18775), .B1(n19871), .B2(n16550), .ZN(
        U349) );
  INV_X1 U19629 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18774) );
  INV_X1 U19630 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19869) );
  AOI22_X1 U19631 ( .A1(n16549), .A2(n18774), .B1(n19869), .B2(n16550), .ZN(
        U350) );
  INV_X1 U19632 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18772) );
  INV_X1 U19633 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19866) );
  AOI22_X1 U19634 ( .A1(n16549), .A2(n18772), .B1(n19866), .B2(n16550), .ZN(
        U351) );
  INV_X1 U19635 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18770) );
  INV_X1 U19636 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19864) );
  AOI22_X1 U19637 ( .A1(n16549), .A2(n18770), .B1(n19864), .B2(n16550), .ZN(
        U352) );
  INV_X1 U19638 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18768) );
  INV_X1 U19639 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19863) );
  AOI22_X1 U19640 ( .A1(n16549), .A2(n18768), .B1(n19863), .B2(n16550), .ZN(
        U353) );
  INV_X1 U19641 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18766) );
  AOI22_X1 U19642 ( .A1(n16549), .A2(n18766), .B1(n19861), .B2(n16550), .ZN(
        U354) );
  INV_X1 U19643 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18819) );
  INV_X1 U19644 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19910) );
  AOI22_X1 U19645 ( .A1(n16549), .A2(n18819), .B1(n19910), .B2(n16550), .ZN(
        U356) );
  INV_X1 U19646 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18816) );
  INV_X1 U19647 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19908) );
  AOI22_X1 U19648 ( .A1(n16549), .A2(n18816), .B1(n19908), .B2(n16550), .ZN(
        U357) );
  INV_X1 U19649 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18814) );
  INV_X1 U19650 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19906) );
  AOI22_X1 U19651 ( .A1(n16549), .A2(n18814), .B1(n19906), .B2(n16550), .ZN(
        U358) );
  INV_X1 U19652 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18812) );
  INV_X1 U19653 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19905) );
  AOI22_X1 U19654 ( .A1(n16549), .A2(n18812), .B1(n19905), .B2(n16550), .ZN(
        U359) );
  INV_X1 U19655 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18810) );
  INV_X1 U19656 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19904) );
  AOI22_X1 U19657 ( .A1(n16549), .A2(n18810), .B1(n19904), .B2(n16550), .ZN(
        U360) );
  INV_X1 U19658 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18808) );
  INV_X1 U19659 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19902) );
  AOI22_X1 U19660 ( .A1(n16549), .A2(n18808), .B1(n19902), .B2(n16550), .ZN(
        U361) );
  INV_X1 U19661 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18805) );
  INV_X1 U19662 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19900) );
  AOI22_X1 U19663 ( .A1(n16549), .A2(n18805), .B1(n19900), .B2(n16550), .ZN(
        U362) );
  INV_X1 U19664 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18804) );
  INV_X1 U19665 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19898) );
  AOI22_X1 U19666 ( .A1(n16549), .A2(n18804), .B1(n19898), .B2(n16550), .ZN(
        U363) );
  INV_X1 U19667 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18802) );
  INV_X1 U19668 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19896) );
  AOI22_X1 U19669 ( .A1(n16549), .A2(n18802), .B1(n19896), .B2(n16550), .ZN(
        U364) );
  INV_X1 U19670 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18764) );
  INV_X1 U19671 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19859) );
  AOI22_X1 U19672 ( .A1(n16549), .A2(n18764), .B1(n19859), .B2(n16550), .ZN(
        U365) );
  INV_X1 U19673 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18799) );
  INV_X1 U19674 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19894) );
  AOI22_X1 U19675 ( .A1(n16549), .A2(n18799), .B1(n19894), .B2(n16550), .ZN(
        U366) );
  INV_X1 U19676 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18798) );
  INV_X1 U19677 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19892) );
  AOI22_X1 U19678 ( .A1(n16549), .A2(n18798), .B1(n19892), .B2(n16550), .ZN(
        U367) );
  INV_X1 U19679 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18796) );
  INV_X1 U19680 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19890) );
  AOI22_X1 U19681 ( .A1(n16549), .A2(n18796), .B1(n19890), .B2(n16550), .ZN(
        U368) );
  INV_X1 U19682 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18794) );
  INV_X1 U19683 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19888) );
  AOI22_X1 U19684 ( .A1(n16549), .A2(n18794), .B1(n19888), .B2(n16550), .ZN(
        U369) );
  INV_X1 U19685 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18792) );
  INV_X1 U19686 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19886) );
  AOI22_X1 U19687 ( .A1(n16549), .A2(n18792), .B1(n19886), .B2(n16550), .ZN(
        U370) );
  INV_X1 U19688 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18789) );
  INV_X1 U19689 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19884) );
  AOI22_X1 U19690 ( .A1(n16549), .A2(n18789), .B1(n19884), .B2(n16550), .ZN(
        U371) );
  INV_X1 U19691 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18787) );
  INV_X1 U19692 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19882) );
  AOI22_X1 U19693 ( .A1(n16549), .A2(n18787), .B1(n19882), .B2(n16550), .ZN(
        U372) );
  INV_X1 U19694 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18786) );
  INV_X1 U19695 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19880) );
  AOI22_X1 U19696 ( .A1(n16549), .A2(n18786), .B1(n19880), .B2(n16550), .ZN(
        U373) );
  INV_X1 U19697 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18784) );
  INV_X1 U19698 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19878) );
  AOI22_X1 U19699 ( .A1(n16549), .A2(n18784), .B1(n19878), .B2(n16550), .ZN(
        U374) );
  INV_X1 U19700 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18782) );
  INV_X1 U19701 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19876) );
  AOI22_X1 U19702 ( .A1(n16549), .A2(n18782), .B1(n19876), .B2(n16550), .ZN(
        U375) );
  INV_X1 U19703 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18762) );
  INV_X1 U19704 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19858) );
  AOI22_X1 U19705 ( .A1(n16549), .A2(n18762), .B1(n19858), .B2(n16550), .ZN(
        U376) );
  NAND2_X1 U19706 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18761), .ZN(n16551) );
  AOI22_X1 U19707 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n16551), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18758), .ZN(n18833) );
  AOI21_X1 U19708 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18833), .ZN(n16552) );
  INV_X1 U19709 ( .A(n16552), .ZN(P3_U2633) );
  INV_X1 U19710 ( .A(n16574), .ZN(n18737) );
  OAI21_X1 U19711 ( .B1(n16557), .B2(n17414), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16553) );
  OAI21_X1 U19712 ( .B1(n16554), .B2(n18737), .A(n16553), .ZN(P3_U2634) );
  INV_X2 U19713 ( .A(n18898), .ZN(n18897) );
  AOI21_X1 U19714 ( .B1(n18758), .B2(n18761), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16555) );
  AOI22_X1 U19715 ( .A1(n18897), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16555), 
        .B2(n18898), .ZN(P3_U2635) );
  OAI21_X1 U19716 ( .B1(n18745), .B2(BS16), .A(n18833), .ZN(n18831) );
  OAI21_X1 U19717 ( .B1(n18833), .B2(n18888), .A(n18831), .ZN(P3_U2636) );
  NOR3_X1 U19718 ( .A1(n16557), .A2(n16556), .A3(n18673), .ZN(n18679) );
  NOR2_X1 U19719 ( .A1(n18679), .A2(n18732), .ZN(n18879) );
  OAI21_X1 U19720 ( .B1(n18879), .B2(n18224), .A(n16558), .ZN(P3_U2637) );
  NOR4_X1 U19721 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16562) );
  NOR4_X1 U19722 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16561) );
  NOR4_X1 U19723 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16560) );
  NOR4_X1 U19724 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16559) );
  NAND4_X1 U19725 ( .A1(n16562), .A2(n16561), .A3(n16560), .A4(n16559), .ZN(
        n16568) );
  NOR4_X1 U19726 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16566) );
  AOI211_X1 U19727 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16565) );
  NOR4_X1 U19728 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16564) );
  NOR4_X1 U19729 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16563) );
  NAND4_X1 U19730 ( .A1(n16566), .A2(n16565), .A3(n16564), .A4(n16563), .ZN(
        n16567) );
  NOR2_X1 U19731 ( .A1(n16568), .A2(n16567), .ZN(n18877) );
  INV_X1 U19732 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16570) );
  NOR3_X1 U19733 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16571) );
  OAI21_X1 U19734 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16571), .A(n18877), .ZN(
        n16569) );
  OAI21_X1 U19735 ( .B1(n18877), .B2(n16570), .A(n16569), .ZN(P3_U2638) );
  INV_X1 U19736 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18870) );
  INV_X1 U19737 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18832) );
  AOI21_X1 U19738 ( .B1(n18870), .B2(n18832), .A(n16571), .ZN(n16573) );
  INV_X1 U19739 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16572) );
  INV_X1 U19740 ( .A(n18877), .ZN(n18872) );
  AOI22_X1 U19741 ( .A1(n18877), .A2(n16573), .B1(n16572), .B2(n18872), .ZN(
        P3_U2639) );
  NOR3_X1 U19742 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .ZN(n18744) );
  NAND2_X1 U19743 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18744), .ZN(n16902) );
  NAND2_X1 U19744 ( .A1(n16574), .A2(n9814), .ZN(n18730) );
  INV_X1 U19745 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18806) );
  INV_X1 U19746 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18788) );
  INV_X1 U19747 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18785) );
  INV_X1 U19748 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18781) );
  INV_X1 U19749 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18771) );
  INV_X1 U19750 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18767) );
  NAND3_X1 U19751 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16910) );
  NOR2_X1 U19752 ( .A1(n18767), .A2(n16910), .ZN(n16885) );
  NAND2_X1 U19753 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16885), .ZN(n16862) );
  NOR2_X1 U19754 ( .A1(n18771), .A2(n16862), .ZN(n16863) );
  NAND3_X1 U19755 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(P3_REIP_REG_7__SCAN_IN), 
        .A3(n16863), .ZN(n16822) );
  INV_X1 U19756 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18779) );
  INV_X1 U19757 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18777) );
  NOR2_X1 U19758 ( .A1(n18779), .A2(n18777), .ZN(n16810) );
  INV_X1 U19759 ( .A(n16810), .ZN(n16833) );
  NOR3_X1 U19760 ( .A1(n18781), .A2(n16822), .A3(n16833), .ZN(n16789) );
  NAND2_X1 U19761 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16789), .ZN(n16786) );
  NOR3_X1 U19762 ( .A1(n18788), .A2(n18785), .A3(n16786), .ZN(n16684) );
  INV_X1 U19763 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18800) );
  INV_X1 U19764 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18790) );
  NAND2_X1 U19765 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .ZN(n16725) );
  NOR2_X1 U19766 ( .A1(n18790), .A2(n16725), .ZN(n16723) );
  NAND3_X1 U19767 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .A3(n16723), .ZN(n16706) );
  NOR2_X1 U19768 ( .A1(n18800), .A2(n16706), .ZN(n16685) );
  NAND4_X1 U19769 ( .A1(n16684), .A2(n16685), .A3(P3_REIP_REG_22__SCAN_IN), 
        .A4(P3_REIP_REG_21__SCAN_IN), .ZN(n16674) );
  NOR2_X1 U19770 ( .A1(n18806), .A2(n16674), .ZN(n16593) );
  NAND2_X1 U19771 ( .A1(n16593), .A2(n16955), .ZN(n16652) );
  NAND3_X1 U19772 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .A3(P3_REIP_REG_24__SCAN_IN), .ZN(n16594) );
  NOR2_X1 U19773 ( .A1(n16652), .A2(n16594), .ZN(n16629) );
  INV_X1 U19774 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18817) );
  INV_X1 U19775 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18818) );
  INV_X1 U19776 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18813) );
  NOR3_X1 U19777 ( .A1(n18817), .A2(n18818), .A3(n18813), .ZN(n16575) );
  OAI211_X1 U19778 ( .C1(n18751), .C2(n16578), .A(n18890), .B(n18888), .ZN(
        n18724) );
  NOR2_X1 U19779 ( .A1(n18901), .A2(n18237), .ZN(n16576) );
  NAND2_X1 U19780 ( .A1(n16955), .A2(n16915), .ZN(n16953) );
  AOI21_X1 U19781 ( .B1(n16629), .B2(n16575), .A(n16724), .ZN(n16614) );
  INV_X1 U19782 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n16577) );
  OAI211_X2 U19783 ( .C1(n16577), .C2(n18889), .A(n18724), .B(n16576), .ZN(
        n16952) );
  AOI22_X1 U19784 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n16614), .B1(
        P3_EBX_REG_31__SCAN_IN), .B2(n16940), .ZN(n16599) );
  NAND2_X1 U19785 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n16578), .ZN(n16579) );
  AOI211_X4 U19786 ( .C1(n18888), .C2(n18890), .A(n16580), .B(n16579), .ZN(
        n16926) );
  NOR3_X1 U19787 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16924) );
  NAND2_X1 U19788 ( .A1(n16924), .A2(n17241), .ZN(n16919) );
  NOR2_X1 U19789 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16919), .ZN(n16898) );
  NAND2_X1 U19790 ( .A1(n16898), .A2(n17235), .ZN(n16893) );
  INV_X1 U19791 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17224) );
  NAND2_X1 U19792 ( .A1(n16879), .A2(n17224), .ZN(n16868) );
  INV_X1 U19793 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16840) );
  NAND2_X1 U19794 ( .A1(n16852), .A2(n16840), .ZN(n16839) );
  INV_X1 U19795 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16819) );
  NAND2_X1 U19796 ( .A1(n16828), .A2(n16819), .ZN(n16818) );
  NAND2_X1 U19797 ( .A1(n16799), .A2(n16794), .ZN(n16793) );
  INV_X1 U19798 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16767) );
  NAND2_X1 U19799 ( .A1(n16775), .A2(n16767), .ZN(n16765) );
  INV_X1 U19800 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16748) );
  NAND2_X1 U19801 ( .A1(n16756), .A2(n16748), .ZN(n16747) );
  INV_X1 U19802 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16720) );
  NAND2_X1 U19803 ( .A1(n16730), .A2(n16720), .ZN(n16718) );
  INV_X1 U19804 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17044) );
  NAND2_X1 U19805 ( .A1(n16703), .A2(n17044), .ZN(n16696) );
  NAND2_X1 U19806 ( .A1(n16693), .A2(n16679), .ZN(n16678) );
  NAND2_X1 U19807 ( .A1(n16662), .A2(n16653), .ZN(n16642) );
  NOR2_X1 U19808 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16642), .ZN(n16641) );
  INV_X1 U19809 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16636) );
  NAND2_X1 U19810 ( .A1(n16641), .A2(n16636), .ZN(n16635) );
  NOR2_X1 U19811 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16635), .ZN(n16620) );
  INV_X1 U19812 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16987) );
  NAND2_X1 U19813 ( .A1(n16620), .A2(n16987), .ZN(n16600) );
  NOR2_X1 U19814 ( .A1(n16951), .A2(n16600), .ZN(n16605) );
  INV_X1 U19815 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16597) );
  INV_X1 U19816 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16582) );
  NOR2_X1 U19817 ( .A1(n17890), .A2(n17534), .ZN(n16584) );
  NAND2_X1 U19818 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16584), .ZN(
        n16583) );
  AOI21_X1 U19819 ( .B1(n16582), .B2(n16583), .A(n16581), .ZN(n17526) );
  OAI21_X1 U19820 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n16584), .A(
        n16583), .ZN(n17543) );
  INV_X1 U19821 ( .A(n17543), .ZN(n16632) );
  NAND2_X1 U19822 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9930), .ZN(
        n16585) );
  AOI21_X1 U19823 ( .B1(n10127), .B2(n16585), .A(n16584), .ZN(n17551) );
  NOR2_X1 U19824 ( .A1(n17890), .A2(n17569), .ZN(n16589) );
  AND2_X1 U19825 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16589), .ZN(
        n16586) );
  OAI21_X1 U19826 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16586), .A(
        n16585), .ZN(n16587) );
  INV_X1 U19827 ( .A(n16587), .ZN(n17562) );
  INV_X1 U19828 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17576) );
  XOR2_X1 U19829 ( .A(n17576), .B(n16589), .Z(n17585) );
  INV_X1 U19830 ( .A(n17585), .ZN(n16665) );
  NAND2_X1 U19831 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16588), .ZN(
        n17561) );
  AOI21_X1 U19832 ( .B1(n10126), .B2(n17561), .A(n16589), .ZN(n17588) );
  INV_X1 U19833 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16591) );
  INV_X1 U19834 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n16714) );
  NAND2_X1 U19835 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17632), .ZN(
        n16715) );
  NOR2_X1 U19836 ( .A1(n16714), .A2(n16715), .ZN(n16592) );
  NAND2_X1 U19837 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16592), .ZN(
        n16590) );
  AOI22_X1 U19838 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16588), .B1(
        n16591), .B2(n16590), .ZN(n17599) );
  INV_X1 U19839 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17620) );
  XNOR2_X1 U19840 ( .A(n17620), .B(n16592), .ZN(n17616) );
  AOI21_X1 U19841 ( .B1(n16714), .B2(n16715), .A(n16592), .ZN(n17634) );
  INV_X1 U19842 ( .A(n16715), .ZN(n17597) );
  NOR2_X1 U19843 ( .A1(n17890), .A2(n16778), .ZN(n16811) );
  INV_X1 U19844 ( .A(n16811), .ZN(n17721) );
  NOR2_X1 U19845 ( .A1(n17685), .A2(n17721), .ZN(n17683) );
  NAND2_X1 U19846 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17683), .ZN(
        n16764) );
  NOR2_X1 U19847 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16764), .ZN(
        n16733) );
  NOR2_X1 U19848 ( .A1(n17634), .A2(n16708), .ZN(n16707) );
  NOR2_X1 U19849 ( .A1(n16707), .A2(n16911), .ZN(n16695) );
  NOR2_X1 U19850 ( .A1(n17616), .A2(n16695), .ZN(n16694) );
  NOR2_X1 U19851 ( .A1(n16694), .A2(n16911), .ZN(n16687) );
  NOR2_X1 U19852 ( .A1(n17599), .A2(n16687), .ZN(n16686) );
  NOR2_X1 U19853 ( .A1(n16686), .A2(n16911), .ZN(n16673) );
  NOR2_X1 U19854 ( .A1(n17588), .A2(n16673), .ZN(n16672) );
  NOR2_X1 U19855 ( .A1(n16672), .A2(n16911), .ZN(n16664) );
  NOR2_X1 U19856 ( .A1(n16665), .A2(n16664), .ZN(n16663) );
  NOR2_X1 U19857 ( .A1(n16663), .A2(n16911), .ZN(n16656) );
  NOR2_X1 U19858 ( .A1(n17562), .A2(n16656), .ZN(n16655) );
  NOR2_X1 U19859 ( .A1(n16655), .A2(n16911), .ZN(n16644) );
  NOR2_X1 U19860 ( .A1(n17551), .A2(n16644), .ZN(n16643) );
  NOR2_X1 U19861 ( .A1(n16643), .A2(n16911), .ZN(n16631) );
  NOR2_X1 U19862 ( .A1(n16632), .A2(n16631), .ZN(n16630) );
  NOR2_X1 U19863 ( .A1(n16630), .A2(n16911), .ZN(n16622) );
  NOR2_X1 U19864 ( .A1(n17526), .A2(n16622), .ZN(n16621) );
  NOR2_X1 U19865 ( .A1(n16621), .A2(n16911), .ZN(n16609) );
  INV_X1 U19866 ( .A(n16902), .ZN(n18741) );
  NAND2_X1 U19867 ( .A1(n16878), .A2(n18741), .ZN(n16943) );
  NOR3_X1 U19868 ( .A1(n16602), .A2(n16601), .A3(n16943), .ZN(n16596) );
  INV_X1 U19869 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18822) );
  NAND2_X1 U19870 ( .A1(n16939), .A2(n16593), .ZN(n16671) );
  NOR2_X1 U19871 ( .A1(n16594), .A2(n16671), .ZN(n16619) );
  NAND4_X1 U19872 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16619), .ZN(n16603) );
  AOI221_X1 U19873 ( .B1(P3_REIP_REG_31__SCAN_IN), .B2(P3_REIP_REG_30__SCAN_IN), .C1(n18820), .C2(n18822), .A(n16603), .ZN(n16595) );
  AOI211_X1 U19874 ( .C1(n16605), .C2(n16597), .A(n16596), .B(n16595), .ZN(
        n16598) );
  OAI211_X1 U19875 ( .C1(n10123), .C2(n16942), .A(n16599), .B(n16598), .ZN(
        P3_U2640) );
  NAND2_X1 U19876 ( .A1(n16926), .A2(n16600), .ZN(n16617) );
  OAI22_X1 U19877 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16603), .B1(n10122), 
        .B2(n16942), .ZN(n16604) );
  OAI21_X1 U19878 ( .B1(n16940), .B2(n16605), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16606) );
  NOR2_X1 U19879 ( .A1(n16620), .A2(n16987), .ZN(n16618) );
  INV_X1 U19880 ( .A(n16607), .ZN(n16608) );
  AOI211_X1 U19881 ( .C1(n16610), .C2(n16609), .A(n16608), .B(n16902), .ZN(
        n16613) );
  OAI22_X1 U19882 ( .A1(n16611), .A2(n16942), .B1(n16952), .B2(n16987), .ZN(
        n16612) );
  AOI211_X1 U19883 ( .C1(n16614), .C2(P3_REIP_REG_29__SCAN_IN), .A(n16613), 
        .B(n16612), .ZN(n16616) );
  NAND4_X1 U19884 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16619), .A4(n18818), .ZN(n16615) );
  OAI211_X1 U19885 ( .C1(n16618), .C2(n16617), .A(n16616), .B(n16615), .ZN(
        P3_U2642) );
  NAND2_X1 U19886 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16619), .ZN(n16628) );
  AOI22_X1 U19887 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16873), .B1(
        n16940), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16627) );
  NAND2_X1 U19888 ( .A1(n16619), .A2(n18813), .ZN(n16638) );
  OAI21_X1 U19889 ( .B1(n16724), .B2(n16629), .A(n16638), .ZN(n16625) );
  AOI211_X1 U19890 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16635), .A(n16620), .B(
        n16951), .ZN(n16624) );
  AOI211_X1 U19891 ( .C1(n17526), .C2(n16622), .A(n16621), .B(n16902), .ZN(
        n16623) );
  AOI211_X1 U19892 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16625), .A(n16624), 
        .B(n16623), .ZN(n16626) );
  OAI211_X1 U19893 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16628), .A(n16627), 
        .B(n16626), .ZN(P3_U2643) );
  NOR2_X1 U19894 ( .A1(n16724), .A2(n16629), .ZN(n16640) );
  AOI211_X1 U19895 ( .C1(n16632), .C2(n16631), .A(n16630), .B(n16902), .ZN(
        n16634) );
  INV_X1 U19896 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17546) );
  OAI22_X1 U19897 ( .A1(n17546), .A2(n16942), .B1(n16952), .B2(n16636), .ZN(
        n16633) );
  AOI211_X1 U19898 ( .C1(n16640), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16634), 
        .B(n16633), .ZN(n16639) );
  OAI211_X1 U19899 ( .C1(n16641), .C2(n16636), .A(n16926), .B(n16635), .ZN(
        n16637) );
  NAND3_X1 U19900 ( .A1(n16639), .A2(n16638), .A3(n16637), .ZN(P3_U2644) );
  INV_X1 U19901 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18807) );
  NOR2_X1 U19902 ( .A1(n18807), .A2(n16671), .ZN(n16651) );
  AOI21_X1 U19903 ( .B1(P3_REIP_REG_25__SCAN_IN), .B2(n16651), .A(
        P3_REIP_REG_26__SCAN_IN), .ZN(n16650) );
  INV_X1 U19904 ( .A(n16640), .ZN(n16649) );
  AOI22_X1 U19905 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16873), .B1(
        n16940), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16648) );
  AOI211_X1 U19906 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16642), .A(n16641), .B(
        n16951), .ZN(n16646) );
  AOI211_X1 U19907 ( .C1(n17551), .C2(n16644), .A(n16643), .B(n16902), .ZN(
        n16645) );
  NOR2_X1 U19908 ( .A1(n16646), .A2(n16645), .ZN(n16647) );
  OAI211_X1 U19909 ( .C1(n16650), .C2(n16649), .A(n16648), .B(n16647), .ZN(
        P3_U2645) );
  INV_X1 U19910 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18809) );
  AOI22_X1 U19911 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n16873), .B1(
        n16651), .B2(n18809), .ZN(n16661) );
  NAND2_X1 U19912 ( .A1(n16953), .A2(n16652), .ZN(n16682) );
  OAI21_X1 U19913 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n16915), .A(n16682), 
        .ZN(n16659) );
  XOR2_X1 U19914 ( .A(P3_EBX_REG_25__SCAN_IN), .B(n16662), .Z(n16654) );
  OAI22_X1 U19915 ( .A1(n16951), .A2(n16654), .B1(n16653), .B2(n16952), .ZN(
        n16658) );
  AOI211_X1 U19916 ( .C1(n17562), .C2(n16656), .A(n16655), .B(n16902), .ZN(
        n16657) );
  AOI211_X1 U19917 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n16659), .A(n16658), 
        .B(n16657), .ZN(n16660) );
  NAND2_X1 U19918 ( .A1(n16661), .A2(n16660), .ZN(P3_U2646) );
  AOI22_X1 U19919 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16873), .B1(
        n16940), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n16670) );
  INV_X1 U19920 ( .A(n16682), .ZN(n16668) );
  AOI211_X1 U19921 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16678), .A(n16662), .B(
        n16951), .ZN(n16667) );
  AOI211_X1 U19922 ( .C1(n16665), .C2(n16664), .A(n16663), .B(n16902), .ZN(
        n16666) );
  AOI211_X1 U19923 ( .C1(n16668), .C2(P3_REIP_REG_24__SCAN_IN), .A(n16667), 
        .B(n16666), .ZN(n16669) );
  OAI211_X1 U19924 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16671), .A(n16670), 
        .B(n16669), .ZN(P3_U2647) );
  AOI211_X1 U19925 ( .C1(n17588), .C2(n16673), .A(n16672), .B(n16902), .ZN(
        n16677) );
  NOR3_X1 U19926 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16915), .A3(n16674), 
        .ZN(n16676) );
  OAI22_X1 U19927 ( .A1(n10126), .A2(n16942), .B1(n16952), .B2(n16679), .ZN(
        n16675) );
  NOR3_X1 U19928 ( .A1(n16677), .A2(n16676), .A3(n16675), .ZN(n16681) );
  OAI211_X1 U19929 ( .C1(n16693), .C2(n16679), .A(n16926), .B(n16678), .ZN(
        n16680) );
  OAI211_X1 U19930 ( .C1(n16682), .C2(n18806), .A(n16681), .B(n16680), .ZN(
        P3_U2648) );
  AOI21_X1 U19931 ( .B1(n16696), .B2(P3_EBX_REG_22__SCAN_IN), .A(n16951), .ZN(
        n16683) );
  AOI21_X1 U19932 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n16940), .A(n16683), .ZN(
        n16692) );
  OAI21_X1 U19933 ( .B1(n16915), .B2(n16684), .A(n16955), .ZN(n16783) );
  INV_X1 U19934 ( .A(n16783), .ZN(n16722) );
  OAI21_X1 U19935 ( .B1(n16724), .B2(n16685), .A(n16722), .ZN(n16710) );
  AOI22_X1 U19936 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n16873), .B1(
        P3_REIP_REG_22__SCAN_IN), .B2(n16710), .ZN(n16691) );
  INV_X1 U19937 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18803) );
  INV_X1 U19938 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18801) );
  NAND2_X1 U19939 ( .A1(n16685), .A2(n16763), .ZN(n16702) );
  AOI221_X1 U19940 ( .B1(P3_REIP_REG_22__SCAN_IN), .B2(P3_REIP_REG_21__SCAN_IN), .C1(n18803), .C2(n18801), .A(n16702), .ZN(n16689) );
  AOI211_X1 U19941 ( .C1(n17599), .C2(n16687), .A(n16686), .B(n16902), .ZN(
        n16688) );
  NOR2_X1 U19942 ( .A1(n16689), .A2(n16688), .ZN(n16690) );
  OAI211_X1 U19943 ( .C1(n16693), .C2(n16692), .A(n16691), .B(n16690), .ZN(
        P3_U2649) );
  INV_X1 U19944 ( .A(n16710), .ZN(n16701) );
  AOI211_X1 U19945 ( .C1(n17616), .C2(n16695), .A(n16694), .B(n16902), .ZN(
        n16699) );
  OAI211_X1 U19946 ( .C1(n16703), .C2(n17044), .A(n16926), .B(n16696), .ZN(
        n16697) );
  OAI21_X1 U19947 ( .B1(n17044), .B2(n16952), .A(n16697), .ZN(n16698) );
  AOI211_X1 U19948 ( .C1(n16873), .C2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n16699), .B(n16698), .ZN(n16700) );
  OAI221_X1 U19949 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n16702), .C1(n18801), 
        .C2(n16701), .A(n16700), .ZN(P3_U2650) );
  AOI211_X1 U19950 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16718), .A(n16703), .B(
        n16951), .ZN(n16704) );
  AOI21_X1 U19951 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16940), .A(n16704), .ZN(
        n16713) );
  INV_X1 U19952 ( .A(n16763), .ZN(n16705) );
  NOR2_X1 U19953 ( .A1(n16706), .A2(n16705), .ZN(n16711) );
  AOI211_X1 U19954 ( .C1(n17634), .C2(n16708), .A(n16707), .B(n16902), .ZN(
        n16709) );
  AOI221_X1 U19955 ( .B1(n16711), .B2(n18800), .C1(n16710), .C2(
        P3_REIP_REG_20__SCAN_IN), .A(n16709), .ZN(n16712) );
  OAI211_X1 U19956 ( .C1(n16714), .C2(n16942), .A(n16713), .B(n16712), .ZN(
        P3_U2651) );
  NOR2_X1 U19957 ( .A1(n17890), .A2(n17645), .ZN(n17644) );
  NAND2_X1 U19958 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17644), .ZN(
        n16732) );
  INV_X1 U19959 ( .A(n16732), .ZN(n16716) );
  AOI21_X1 U19960 ( .B1(n16733), .B2(n16716), .A(n16911), .ZN(n16717) );
  OAI21_X1 U19961 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16716), .A(
        n16715), .ZN(n17650) );
  XOR2_X1 U19962 ( .A(n16717), .B(n17650), .Z(n16729) );
  OAI211_X1 U19963 ( .C1(n16730), .C2(n16720), .A(n16926), .B(n16718), .ZN(
        n16719) );
  OAI211_X1 U19964 ( .C1(n16952), .C2(n16720), .A(n18201), .B(n16719), .ZN(
        n16721) );
  AOI21_X1 U19965 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16873), .A(
        n16721), .ZN(n16728) );
  OAI21_X1 U19966 ( .B1(n16724), .B2(n16723), .A(n16722), .ZN(n16746) );
  NAND2_X1 U19967 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n16763), .ZN(n16762) );
  NOR2_X1 U19968 ( .A1(n16725), .A2(n16762), .ZN(n16736) );
  INV_X1 U19969 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18797) );
  INV_X1 U19970 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18795) );
  XOR2_X1 U19971 ( .A(n18797), .B(n18795), .Z(n16726) );
  AOI22_X1 U19972 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n16746), .B1(n16736), 
        .B2(n16726), .ZN(n16727) );
  OAI211_X1 U19973 ( .C1(n16902), .C2(n16729), .A(n16728), .B(n16727), .ZN(
        P3_U2652) );
  INV_X1 U19974 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17660) );
  AOI211_X1 U19975 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16747), .A(n16730), .B(
        n16951), .ZN(n16731) );
  AOI211_X1 U19976 ( .C1(n16940), .C2(P3_EBX_REG_18__SCAN_IN), .A(n17990), .B(
        n16731), .ZN(n16738) );
  OAI21_X1 U19977 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17644), .A(
        n16732), .ZN(n17657) );
  INV_X1 U19978 ( .A(n16733), .ZN(n16753) );
  INV_X1 U19979 ( .A(n17644), .ZN(n16740) );
  OAI21_X1 U19980 ( .B1(n16753), .B2(n16740), .A(n16878), .ZN(n16742) );
  OAI21_X1 U19981 ( .B1(n17657), .B2(n16742), .A(n18741), .ZN(n16734) );
  AOI21_X1 U19982 ( .B1(n17657), .B2(n16742), .A(n16734), .ZN(n16735) );
  AOI221_X1 U19983 ( .B1(n16736), .B2(n18795), .C1(n16746), .C2(
        P3_REIP_REG_18__SCAN_IN), .A(n16735), .ZN(n16737) );
  OAI211_X1 U19984 ( .C1(n17660), .C2(n16942), .A(n16738), .B(n16737), .ZN(
        P3_U2653) );
  AOI22_X1 U19985 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16873), .B1(
        n16940), .B2(P3_EBX_REG_17__SCAN_IN), .ZN(n16751) );
  INV_X1 U19986 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18791) );
  NOR3_X1 U19987 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n18791), .A3(n16762), 
        .ZN(n16745) );
  INV_X1 U19988 ( .A(n17683), .ZN(n16739) );
  NOR2_X1 U19989 ( .A1(n17686), .A2(n16739), .ZN(n16752) );
  INV_X1 U19990 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16941) );
  OAI21_X1 U19991 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16752), .A(
        n16740), .ZN(n17669) );
  AOI21_X1 U19992 ( .B1(n16752), .B2(n16941), .A(n17669), .ZN(n16741) );
  OR2_X1 U19993 ( .A1(n16741), .A2(n16902), .ZN(n16743) );
  NOR2_X1 U19994 ( .A1(n16902), .A2(n16878), .ZN(n16897) );
  INV_X1 U19995 ( .A(n16897), .ZN(n16938) );
  AOI22_X1 U19996 ( .A1(n16743), .A2(n16938), .B1(n17669), .B2(n16742), .ZN(
        n16744) );
  AOI211_X1 U19997 ( .C1(P3_REIP_REG_17__SCAN_IN), .C2(n16746), .A(n16745), 
        .B(n16744), .ZN(n16750) );
  OAI211_X1 U19998 ( .C1(n16756), .C2(n16748), .A(n16926), .B(n16747), .ZN(
        n16749) );
  NAND4_X1 U19999 ( .A1(n16751), .A2(n16750), .A3(n18201), .A4(n16749), .ZN(
        P3_U2654) );
  AOI21_X1 U20000 ( .B1(n16953), .B2(n18790), .A(n16783), .ZN(n16774) );
  INV_X1 U20001 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16757) );
  AOI21_X1 U20002 ( .B1(n16757), .B2(n16764), .A(n16752), .ZN(n16755) );
  NAND2_X1 U20003 ( .A1(n16753), .A2(n16878), .ZN(n16754) );
  INV_X1 U20004 ( .A(n16754), .ZN(n16770) );
  INV_X1 U20005 ( .A(n16755), .ZN(n17689) );
  AOI221_X1 U20006 ( .B1(n16755), .B2(n16770), .C1(n17689), .C2(n16754), .A(
        n16902), .ZN(n16760) );
  AOI211_X1 U20007 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16765), .A(n16756), .B(
        n16951), .ZN(n16759) );
  INV_X1 U20008 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17113) );
  OAI22_X1 U20009 ( .A1(n16757), .A2(n16942), .B1(n16952), .B2(n17113), .ZN(
        n16758) );
  NOR4_X1 U20010 ( .A1(n18218), .A2(n16760), .A3(n16759), .A4(n16758), .ZN(
        n16761) );
  OAI221_X1 U20011 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(n16762), .C1(n18791), 
        .C2(n16774), .A(n16761), .ZN(P3_U2655) );
  NOR2_X1 U20012 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n16763), .ZN(n16773) );
  OAI21_X1 U20013 ( .B1(n16911), .B2(n16941), .A(n18741), .ZN(n16950) );
  OAI21_X1 U20014 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17683), .A(
        n16764), .ZN(n17694) );
  AOI211_X1 U20015 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n16938), .A(
        n16950), .B(n17694), .ZN(n16769) );
  OAI211_X1 U20016 ( .C1(n16775), .C2(n16767), .A(n16926), .B(n16765), .ZN(
        n16766) );
  OAI211_X1 U20017 ( .C1(n16952), .C2(n16767), .A(n18201), .B(n16766), .ZN(
        n16768) );
  AOI211_X1 U20018 ( .C1(n16873), .C2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16769), .B(n16768), .ZN(n16772) );
  NAND3_X1 U20019 ( .A1(n18741), .A2(n16770), .A3(n17694), .ZN(n16771) );
  OAI211_X1 U20020 ( .C1(n16774), .C2(n16773), .A(n16772), .B(n16771), .ZN(
        P3_U2656) );
  INV_X1 U20021 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17709) );
  AOI211_X1 U20022 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16793), .A(n16775), .B(
        n16951), .ZN(n16776) );
  AOI211_X1 U20023 ( .C1(n16940), .C2(P3_EBX_REG_14__SCAN_IN), .A(n17990), .B(
        n16776), .ZN(n16785) );
  NOR3_X1 U20024 ( .A1(n16915), .A2(n18785), .A3(n16786), .ZN(n16782) );
  NAND2_X1 U20025 ( .A1(n16779), .A2(n16811), .ZN(n16777) );
  AOI21_X1 U20026 ( .B1(n17709), .B2(n16777), .A(n17683), .ZN(n17711) );
  NAND2_X1 U20027 ( .A1(n16941), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16886) );
  OAI21_X1 U20028 ( .B1(n16778), .B2(n16886), .A(n16878), .ZN(n16802) );
  OAI21_X1 U20029 ( .B1(n16779), .B2(n16911), .A(n16802), .ZN(n16788) );
  OAI21_X1 U20030 ( .B1(n17711), .B2(n16788), .A(n18741), .ZN(n16780) );
  AOI21_X1 U20031 ( .B1(n17711), .B2(n16788), .A(n16780), .ZN(n16781) );
  AOI221_X1 U20032 ( .B1(P3_REIP_REG_14__SCAN_IN), .B2(n16783), .C1(n16782), 
        .C2(n16783), .A(n16781), .ZN(n16784) );
  OAI211_X1 U20033 ( .C1(n17709), .C2(n16942), .A(n16785), .B(n16784), .ZN(
        P3_U2657) );
  AOI21_X1 U20034 ( .B1(n16940), .B2(P3_EBX_REG_13__SCAN_IN), .A(n17990), .ZN(
        n16798) );
  NOR2_X1 U20035 ( .A1(n16915), .A2(n16786), .ZN(n16787) );
  AOI22_X1 U20036 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n16873), .B1(
        n16787), .B2(n18785), .ZN(n16797) );
  AND2_X1 U20037 ( .A1(n16788), .A2(n18741), .ZN(n16792) );
  INV_X1 U20038 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16805) );
  NOR2_X1 U20039 ( .A1(n16805), .A2(n17721), .ZN(n16801) );
  OAI22_X1 U20040 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n16801), .B1(
        n17721), .B2(n17725), .ZN(n17727) );
  INV_X1 U20041 ( .A(n16789), .ZN(n16804) );
  AOI21_X1 U20042 ( .B1(n16939), .B2(n16804), .A(n16947), .ZN(n16815) );
  INV_X1 U20043 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18783) );
  NAND2_X1 U20044 ( .A1(n16939), .A2(n18783), .ZN(n16803) );
  AOI21_X1 U20045 ( .B1(n16815), .B2(n16803), .A(n18785), .ZN(n16791) );
  AOI211_X1 U20046 ( .C1(n16878), .C2(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n16950), .B(n17727), .ZN(n16790) );
  AOI211_X1 U20047 ( .C1(n16792), .C2(n17727), .A(n16791), .B(n16790), .ZN(
        n16796) );
  OAI211_X1 U20048 ( .C1(n16799), .C2(n16794), .A(n16926), .B(n16793), .ZN(
        n16795) );
  NAND4_X1 U20049 ( .A1(n16798), .A2(n16797), .A3(n16796), .A4(n16795), .ZN(
        P3_U2658) );
  AOI211_X1 U20050 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16818), .A(n16799), .B(
        n16951), .ZN(n16800) );
  AOI21_X1 U20051 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n16940), .A(n16800), .ZN(
        n16809) );
  AOI21_X1 U20052 ( .B1(n16805), .B2(n17721), .A(n16801), .ZN(n17734) );
  XNOR2_X1 U20053 ( .A(n17734), .B(n16802), .ZN(n16807) );
  OAI22_X1 U20054 ( .A1(n16805), .A2(n16942), .B1(n16804), .B2(n16803), .ZN(
        n16806) );
  AOI211_X1 U20055 ( .C1(n18741), .C2(n16807), .A(n17990), .B(n16806), .ZN(
        n16808) );
  OAI211_X1 U20056 ( .C1(n16815), .C2(n18783), .A(n16809), .B(n16808), .ZN(
        P3_U2659) );
  INV_X1 U20057 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18776) );
  NAND3_X1 U20058 ( .A1(n16939), .A2(P3_REIP_REG_7__SCAN_IN), .A3(n16863), 
        .ZN(n16851) );
  NOR2_X1 U20059 ( .A1(n18776), .A2(n16851), .ZN(n16845) );
  AOI21_X1 U20060 ( .B1(n16810), .B2(n16845), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16816) );
  INV_X1 U20061 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17790) );
  NOR3_X1 U20062 ( .A1(n17890), .A2(n17787), .A3(n17790), .ZN(n16836) );
  NAND3_X1 U20063 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A3(n16836), .ZN(n16823) );
  AOI21_X1 U20064 ( .B1(n17750), .B2(n16823), .A(n16811), .ZN(n17753) );
  OR2_X1 U20065 ( .A1(n17787), .A2(n16886), .ZN(n16849) );
  OAI21_X1 U20066 ( .B1(n16812), .B2(n16849), .A(n16878), .ZN(n16813) );
  XOR2_X1 U20067 ( .A(n17753), .B(n16813), .Z(n16814) );
  OAI22_X1 U20068 ( .A1(n16816), .A2(n16815), .B1(n16902), .B2(n16814), .ZN(
        n16817) );
  AOI211_X1 U20069 ( .C1(n16940), .C2(P3_EBX_REG_11__SCAN_IN), .A(n17990), .B(
        n16817), .ZN(n16821) );
  OAI211_X1 U20070 ( .C1(n16828), .C2(n16819), .A(n16926), .B(n16818), .ZN(
        n16820) );
  OAI211_X1 U20071 ( .C1(n16942), .C2(n17750), .A(n16821), .B(n16820), .ZN(
        P3_U2660) );
  AOI21_X1 U20072 ( .B1(n16939), .B2(n16822), .A(n16947), .ZN(n16850) );
  INV_X1 U20073 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17778) );
  INV_X1 U20074 ( .A(n16836), .ZN(n16848) );
  NOR2_X1 U20075 ( .A1(n17778), .A2(n16848), .ZN(n16824) );
  OAI21_X1 U20076 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16824), .A(
        n16823), .ZN(n17769) );
  INV_X1 U20077 ( .A(n17769), .ZN(n16827) );
  NOR3_X1 U20078 ( .A1(n17790), .A2(n17778), .A3(n16849), .ZN(n16825) );
  NOR2_X1 U20079 ( .A1(n16825), .A2(n16911), .ZN(n16838) );
  INV_X1 U20080 ( .A(n16838), .ZN(n16826) );
  AOI221_X1 U20081 ( .B1(n16827), .B2(n16838), .C1(n17769), .C2(n16826), .A(
        n16902), .ZN(n16832) );
  AOI211_X1 U20082 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16839), .A(n16828), .B(
        n16951), .ZN(n16831) );
  AOI22_X1 U20083 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16873), .B1(
        n16940), .B2(P3_EBX_REG_10__SCAN_IN), .ZN(n16829) );
  INV_X1 U20084 ( .A(n16829), .ZN(n16830) );
  NOR4_X1 U20085 ( .A1(n18218), .A2(n16832), .A3(n16831), .A4(n16830), .ZN(
        n16835) );
  OAI211_X1 U20086 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(P3_REIP_REG_9__SCAN_IN), 
        .A(n16845), .B(n16833), .ZN(n16834) );
  OAI211_X1 U20087 ( .C1(n16850), .C2(n18779), .A(n16835), .B(n16834), .ZN(
        P3_U2661) );
  AOI22_X1 U20088 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16848), .B1(
        n16836), .B2(n17778), .ZN(n17780) );
  NOR2_X1 U20089 ( .A1(n17790), .A2(n16849), .ZN(n16837) );
  AOI22_X1 U20090 ( .A1(n16838), .A2(n17780), .B1(n16837), .B2(n17778), .ZN(
        n16847) );
  OAI22_X1 U20091 ( .A1(n18777), .A2(n16850), .B1(n17780), .B2(n16938), .ZN(
        n16844) );
  AOI22_X1 U20092 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16873), .B1(
        n16940), .B2(P3_EBX_REG_9__SCAN_IN), .ZN(n16842) );
  OAI211_X1 U20093 ( .C1(n16852), .C2(n16840), .A(n16926), .B(n16839), .ZN(
        n16841) );
  NAND3_X1 U20094 ( .A1(n16842), .A2(n18201), .A3(n16841), .ZN(n16843) );
  AOI211_X1 U20095 ( .C1(n16845), .C2(n18777), .A(n16844), .B(n16843), .ZN(
        n16846) );
  OAI21_X1 U20096 ( .B1(n16847), .B2(n16902), .A(n16846), .ZN(P3_U2662) );
  NOR2_X1 U20097 ( .A1(n17890), .A2(n17787), .ZN(n16858) );
  OAI21_X1 U20098 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16858), .A(
        n16848), .ZN(n17792) );
  NAND2_X1 U20099 ( .A1(n16878), .A2(n16849), .ZN(n16860) );
  XNOR2_X1 U20100 ( .A(n17792), .B(n16860), .ZN(n16857) );
  AOI21_X1 U20101 ( .B1(n16940), .B2(P3_EBX_REG_8__SCAN_IN), .A(n17990), .ZN(
        n16856) );
  AOI21_X1 U20102 ( .B1(n18776), .B2(n16851), .A(n16850), .ZN(n16854) );
  AOI211_X1 U20103 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16868), .A(n16852), .B(
        n16951), .ZN(n16853) );
  AOI211_X1 U20104 ( .C1(n16873), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16854), .B(n16853), .ZN(n16855) );
  OAI211_X1 U20105 ( .C1(n16902), .C2(n16857), .A(n16856), .B(n16855), .ZN(
        P3_U2663) );
  NOR2_X1 U20106 ( .A1(n17890), .A2(n17826), .ZN(n16887) );
  NAND2_X1 U20107 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16887), .ZN(
        n16872) );
  AOI21_X1 U20108 ( .B1(n10129), .B2(n16872), .A(n16858), .ZN(n17812) );
  INV_X1 U20109 ( .A(n17812), .ZN(n16861) );
  NOR2_X1 U20110 ( .A1(n10134), .A2(n16886), .ZN(n16871) );
  OAI21_X1 U20111 ( .B1(n16871), .B2(n16861), .A(n18741), .ZN(n16859) );
  AOI22_X1 U20112 ( .A1(n16861), .A2(n16860), .B1(n16938), .B2(n16859), .ZN(
        n16867) );
  AOI21_X1 U20113 ( .B1(n16939), .B2(n16862), .A(n16947), .ZN(n16891) );
  NAND4_X1 U20114 ( .A1(n16939), .A2(P3_REIP_REG_5__SCAN_IN), .A3(n16885), 
        .A4(n18771), .ZN(n16877) );
  INV_X1 U20115 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18773) );
  AOI21_X1 U20116 ( .B1(n16891), .B2(n16877), .A(n18773), .ZN(n16866) );
  NAND2_X1 U20117 ( .A1(n16939), .A2(n16863), .ZN(n16864) );
  OAI22_X1 U20118 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n16864), .B1(n16952), 
        .B2(n17224), .ZN(n16865) );
  NOR4_X1 U20119 ( .A1(n17990), .A2(n16867), .A3(n16866), .A4(n16865), .ZN(
        n16870) );
  OAI211_X1 U20120 ( .C1(n16879), .C2(n17224), .A(n16926), .B(n16868), .ZN(
        n16869) );
  OAI211_X1 U20121 ( .C1(n16942), .C2(n10129), .A(n16870), .B(n16869), .ZN(
        P3_U2664) );
  NOR2_X1 U20122 ( .A1(n16871), .A2(n16943), .ZN(n16876) );
  OAI21_X1 U20123 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16887), .A(
        n16872), .ZN(n17828) );
  AOI22_X1 U20124 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16873), .B1(
        n16940), .B2(P3_EBX_REG_6__SCAN_IN), .ZN(n16874) );
  INV_X1 U20125 ( .A(n16874), .ZN(n16875) );
  AOI21_X1 U20126 ( .B1(n16876), .B2(n17828), .A(n16875), .ZN(n16884) );
  INV_X1 U20127 ( .A(n16877), .ZN(n16882) );
  AOI211_X1 U20128 ( .C1(n16878), .C2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16950), .B(n17828), .ZN(n16881) );
  AOI211_X1 U20129 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16893), .A(n16879), .B(
        n16951), .ZN(n16880) );
  NOR4_X1 U20130 ( .A1(n18218), .A2(n16882), .A3(n16881), .A4(n16880), .ZN(
        n16883) );
  OAI211_X1 U20131 ( .C1(n16891), .C2(n18771), .A(n16884), .B(n16883), .ZN(
        P3_U2665) );
  AOI21_X1 U20132 ( .B1(n16939), .B2(n16885), .A(P3_REIP_REG_5__SCAN_IN), .ZN(
        n16890) );
  INV_X1 U20133 ( .A(n16886), .ZN(n16935) );
  AOI21_X1 U20134 ( .B1(n17838), .B2(n16935), .A(n16911), .ZN(n16901) );
  AND2_X1 U20135 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17838), .ZN(
        n16896) );
  INV_X1 U20136 ( .A(n16887), .ZN(n16888) );
  OAI21_X1 U20137 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n16896), .A(
        n16888), .ZN(n17841) );
  XOR2_X1 U20138 ( .A(n16901), .B(n17841), .Z(n16889) );
  OAI22_X1 U20139 ( .A1(n16891), .A2(n16890), .B1(n16902), .B2(n16889), .ZN(
        n16892) );
  AOI211_X1 U20140 ( .C1(n16940), .C2(P3_EBX_REG_5__SCAN_IN), .A(n17990), .B(
        n16892), .ZN(n16895) );
  OAI211_X1 U20141 ( .C1(n16898), .C2(n17235), .A(n16926), .B(n16893), .ZN(
        n16894) );
  OAI211_X1 U20142 ( .C1(n16942), .C2(n10133), .A(n16895), .B(n16894), .ZN(
        P3_U2666) );
  NAND2_X1 U20143 ( .A1(n16939), .A2(n18767), .ZN(n16909) );
  OR2_X1 U20144 ( .A1(n17890), .A2(n17845), .ZN(n16912) );
  AOI21_X1 U20145 ( .B1(n17859), .B2(n16912), .A(n16896), .ZN(n17856) );
  AOI22_X1 U20146 ( .A1(n16940), .A2(P3_EBX_REG_4__SCAN_IN), .B1(n17856), .B2(
        n16897), .ZN(n16908) );
  AOI211_X1 U20147 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16919), .A(n16898), .B(
        n16951), .ZN(n16906) );
  NAND2_X1 U20148 ( .A1(n18237), .A2(n18886), .ZN(n18904) );
  INV_X1 U20149 ( .A(n18904), .ZN(n16933) );
  OAI21_X1 U20150 ( .B1(n17195), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n16933), .ZN(n16899) );
  OAI211_X1 U20151 ( .C1(n17859), .C2(n16942), .A(n18201), .B(n16899), .ZN(
        n16905) );
  NOR2_X1 U20152 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17845), .ZN(
        n17851) );
  INV_X1 U20153 ( .A(n17856), .ZN(n16900) );
  AOI22_X1 U20154 ( .A1(n16935), .A2(n17851), .B1(n16901), .B2(n16900), .ZN(
        n16903) );
  AOI21_X1 U20155 ( .B1(n16939), .B2(n16910), .A(n16947), .ZN(n16914) );
  OAI22_X1 U20156 ( .A1(n16903), .A2(n16902), .B1(n18767), .B2(n16914), .ZN(
        n16904) );
  NOR3_X1 U20157 ( .A1(n16906), .A2(n16905), .A3(n16904), .ZN(n16907) );
  OAI211_X1 U20158 ( .C1(n16910), .C2(n16909), .A(n16908), .B(n16907), .ZN(
        P3_U2667) );
  INV_X1 U20159 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16922) );
  AOI21_X1 U20160 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n16935), .A(
        n16911), .ZN(n16934) );
  INV_X1 U20161 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17881) );
  NOR2_X1 U20162 ( .A1(n17890), .A2(n17881), .ZN(n16913) );
  OAI21_X1 U20163 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n16913), .A(
        n16912), .ZN(n17869) );
  XNOR2_X1 U20164 ( .A(n16934), .B(n17869), .ZN(n16918) );
  INV_X1 U20165 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18765) );
  NAND2_X1 U20166 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16928) );
  AOI221_X1 U20167 ( .B1(n16915), .B2(n18765), .C1(n16928), .C2(n18765), .A(
        n16914), .ZN(n16917) );
  INV_X1 U20168 ( .A(n18690), .ZN(n18706) );
  NOR2_X1 U20169 ( .A1(n18869), .A2(n18706), .ZN(n16923) );
  INV_X1 U20170 ( .A(n16923), .ZN(n18692) );
  AOI21_X1 U20171 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18692), .A(
        n17143), .ZN(n18836) );
  OAI22_X1 U20172 ( .A1(n18836), .A2(n18904), .B1(n16952), .B2(n17241), .ZN(
        n16916) );
  AOI211_X1 U20173 ( .C1(n18741), .C2(n16918), .A(n16917), .B(n16916), .ZN(
        n16921) );
  OAI211_X1 U20174 ( .C1(n16924), .C2(n17241), .A(n16926), .B(n16919), .ZN(
        n16920) );
  OAI211_X1 U20175 ( .C1(n16942), .C2(n16922), .A(n16921), .B(n16920), .ZN(
        P3_U2668) );
  AOI22_X1 U20176 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17881), .B1(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17890), .ZN(n17878) );
  AOI21_X1 U20177 ( .B1(n18851), .B2(n18704), .A(n16923), .ZN(n18848) );
  OAI22_X1 U20178 ( .A1(n17881), .A2(n16942), .B1(n16952), .B2(n17250), .ZN(
        n16932) );
  INV_X1 U20179 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18763) );
  NOR2_X1 U20180 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n16927) );
  INV_X1 U20181 ( .A(n16924), .ZN(n16925) );
  OAI211_X1 U20182 ( .C1(n16927), .C2(n17250), .A(n16926), .B(n16925), .ZN(
        n16930) );
  OAI211_X1 U20183 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n16939), .B(n16928), .ZN(n16929) );
  OAI211_X1 U20184 ( .C1(n18763), .C2(n16955), .A(n16930), .B(n16929), .ZN(
        n16931) );
  AOI211_X1 U20185 ( .C1(n18848), .C2(n16933), .A(n16932), .B(n16931), .ZN(
        n16937) );
  OAI211_X1 U20186 ( .C1(n16935), .C2(n17878), .A(n18741), .B(n16934), .ZN(
        n16936) );
  OAI211_X1 U20187 ( .C1(n16938), .C2(n17878), .A(n16937), .B(n16936), .ZN(
        P3_U2669) );
  AOI22_X1 U20188 ( .A1(n16940), .A2(P3_EBX_REG_1__SCAN_IN), .B1(n16939), .B2(
        n18870), .ZN(n16949) );
  AOI221_X1 U20189 ( .B1(n16943), .B2(n16942), .C1(n16941), .C2(n16942), .A(
        n17890), .ZN(n16946) );
  OAI21_X1 U20190 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n17251), .ZN(n17259) );
  NAND2_X1 U20191 ( .A1(n18704), .A2(n16944), .ZN(n18853) );
  OAI22_X1 U20192 ( .A1(n16951), .A2(n17259), .B1(n18853), .B2(n18904), .ZN(
        n16945) );
  AOI211_X1 U20193 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(n16947), .A(n16946), .B(
        n16945), .ZN(n16948) );
  OAI211_X1 U20194 ( .C1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n16950), .A(
        n16949), .B(n16948), .ZN(P3_U2670) );
  NAND2_X1 U20195 ( .A1(n16952), .A2(n16951), .ZN(n16954) );
  AOI22_X1 U20196 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n16954), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n16953), .ZN(n16957) );
  NAND3_X1 U20197 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18900), .A3(
        n16955), .ZN(n16956) );
  OAI211_X1 U20198 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n18904), .A(
        n16957), .B(n16956), .ZN(P3_U2671) );
  AOI22_X1 U20199 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n9817), .B1(
        P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n17188), .ZN(n16961) );
  AOI22_X1 U20200 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16960) );
  AOI22_X1 U20201 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n17195), .ZN(n16959) );
  AOI22_X1 U20202 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17213), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16958) );
  NAND4_X1 U20203 ( .A1(n16961), .A2(n16960), .A3(n16959), .A4(n16958), .ZN(
        n16968) );
  AOI22_X1 U20204 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n17019), .B1(
        n13703), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16966) );
  AOI22_X1 U20205 ( .A1(n9820), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16965) );
  AOI22_X1 U20206 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17179), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16964) );
  AOI22_X1 U20207 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n16962), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16963) );
  NAND4_X1 U20208 ( .A1(n16966), .A2(n16965), .A3(n16964), .A4(n16963), .ZN(
        n16967) );
  NOR2_X1 U20209 ( .A1(n16968), .A2(n16967), .ZN(n16980) );
  AOI22_X1 U20210 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16979) );
  AOI22_X1 U20211 ( .A1(n9820), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16978) );
  AOI22_X1 U20212 ( .A1(n17179), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n15691), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16969) );
  OAI21_X1 U20213 ( .B1(n16970), .B2(n17232), .A(n16969), .ZN(n16976) );
  AOI22_X1 U20214 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16974) );
  AOI22_X1 U20215 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13697), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16973) );
  AOI22_X1 U20216 ( .A1(n17197), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n16962), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16972) );
  AOI22_X1 U20217 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13703), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16971) );
  NAND4_X1 U20218 ( .A1(n16974), .A2(n16973), .A3(n16972), .A4(n16971), .ZN(
        n16975) );
  AOI211_X1 U20219 ( .C1(n9817), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n16976), .B(n16975), .ZN(n16977) );
  NAND3_X1 U20220 ( .A1(n16979), .A2(n16978), .A3(n16977), .ZN(n16985) );
  NAND2_X1 U20221 ( .A1(n16986), .A2(n16985), .ZN(n16984) );
  XNOR2_X1 U20222 ( .A(n16980), .B(n16984), .ZN(n17272) );
  NOR2_X1 U20223 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16981), .ZN(n16983) );
  OAI22_X1 U20224 ( .A1(n17272), .A2(n17246), .B1(n16983), .B2(n16982), .ZN(
        P3_U2673) );
  OAI21_X1 U20225 ( .B1(n16986), .B2(n16985), .A(n16984), .ZN(n17279) );
  AOI22_X1 U20226 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16989), .B1(n16988), 
        .B2(n16987), .ZN(n16990) );
  OAI21_X1 U20227 ( .B1(n17279), .B2(n17246), .A(n16990), .ZN(P3_U2674) );
  OAI21_X1 U20228 ( .B1(n16995), .B2(n16992), .A(n16991), .ZN(n17288) );
  NAND3_X1 U20229 ( .A1(n16994), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n17246), 
        .ZN(n16993) );
  OAI221_X1 U20230 ( .B1(n16994), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n17246), 
        .C2(n17288), .A(n16993), .ZN(P3_U2676) );
  AOI21_X1 U20231 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17246), .A(n17005), .ZN(
        n16998) );
  AOI21_X1 U20232 ( .B1(n16996), .B2(n17002), .A(n16995), .ZN(n17289) );
  INV_X1 U20233 ( .A(n17289), .ZN(n16997) );
  OAI22_X1 U20234 ( .A1(n16999), .A2(n16998), .B1(n16997), .B2(n17246), .ZN(
        P3_U2677) );
  INV_X1 U20235 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n17001) );
  INV_X1 U20236 ( .A(n17000), .ZN(n17045) );
  NAND2_X1 U20237 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17045), .ZN(n17031) );
  NOR2_X1 U20238 ( .A1(n17001), .A2(n17031), .ZN(n17011) );
  AND2_X1 U20239 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n17011), .ZN(n17016) );
  AND2_X1 U20240 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17016), .ZN(n17010) );
  AOI21_X1 U20241 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17246), .A(n17010), .ZN(
        n17004) );
  OAI21_X1 U20242 ( .B1(n17006), .B2(n17003), .A(n17002), .ZN(n17298) );
  OAI22_X1 U20243 ( .A1(n17005), .A2(n17004), .B1(n17298), .B2(n17246), .ZN(
        P3_U2678) );
  AOI21_X1 U20244 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17246), .A(n17016), .ZN(
        n17009) );
  AOI21_X1 U20245 ( .B1(n17007), .B2(n17012), .A(n17006), .ZN(n17299) );
  INV_X1 U20246 ( .A(n17299), .ZN(n17008) );
  OAI22_X1 U20247 ( .A1(n17010), .A2(n17009), .B1(n17008), .B2(n17246), .ZN(
        P3_U2679) );
  AOI21_X1 U20248 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17246), .A(n17011), .ZN(
        n17015) );
  OAI21_X1 U20249 ( .B1(n17014), .B2(n17013), .A(n17012), .ZN(n17309) );
  OAI22_X1 U20250 ( .A1(n17016), .A2(n17015), .B1(n17309), .B2(n17246), .ZN(
        P3_U2680) );
  AOI22_X1 U20251 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n15699), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17028) );
  AOI22_X1 U20252 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17027) );
  AOI22_X1 U20253 ( .A1(n17197), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17017) );
  OAI21_X1 U20254 ( .B1(n17018), .B2(n17232), .A(n17017), .ZN(n17025) );
  AOI22_X1 U20255 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17023) );
  AOI22_X1 U20256 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17022) );
  AOI22_X1 U20257 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17019), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17021) );
  AOI22_X1 U20258 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17020) );
  NAND4_X1 U20259 ( .A1(n17023), .A2(n17022), .A3(n17021), .A4(n17020), .ZN(
        n17024) );
  AOI211_X1 U20260 ( .C1(n9820), .C2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n17025), .B(n17024), .ZN(n17026) );
  NAND3_X1 U20261 ( .A1(n17028), .A2(n17027), .A3(n17026), .ZN(n17310) );
  INV_X1 U20262 ( .A(n17310), .ZN(n17030) );
  NAND3_X1 U20263 ( .A1(n17031), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17246), 
        .ZN(n17029) );
  OAI221_X1 U20264 ( .B1(n17031), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17246), 
        .C2(n17030), .A(n17029), .ZN(P3_U2681) );
  AOI22_X1 U20265 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9820), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17035) );
  AOI22_X1 U20266 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17034) );
  AOI22_X1 U20267 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n15691), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17033) );
  AOI22_X1 U20268 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17032) );
  NAND4_X1 U20269 ( .A1(n17035), .A2(n17034), .A3(n17033), .A4(n17032), .ZN(
        n17041) );
  AOI22_X1 U20270 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13703), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17039) );
  AOI22_X1 U20271 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17179), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17038) );
  AOI22_X1 U20272 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17037) );
  AOI22_X1 U20273 ( .A1(n17197), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17036) );
  NAND4_X1 U20274 ( .A1(n17039), .A2(n17038), .A3(n17037), .A4(n17036), .ZN(
        n17040) );
  NOR2_X1 U20275 ( .A1(n17041), .A2(n17040), .ZN(n17317) );
  NOR2_X1 U20276 ( .A1(n17042), .A2(n17070), .ZN(n17043) );
  NOR2_X1 U20277 ( .A1(n17261), .A2(n17043), .ZN(n17057) );
  AOI22_X1 U20278 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17057), .B1(n17045), 
        .B2(n17044), .ZN(n17046) );
  OAI21_X1 U20279 ( .B1(n17317), .B2(n17246), .A(n17046), .ZN(P3_U2682) );
  AOI22_X1 U20280 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17050) );
  AOI22_X1 U20281 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17049) );
  AOI22_X1 U20282 ( .A1(n15710), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n15700), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17048) );
  AOI22_X1 U20283 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n15713), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17047) );
  NAND4_X1 U20284 ( .A1(n17050), .A2(n17049), .A3(n17048), .A4(n17047), .ZN(
        n17056) );
  AOI22_X1 U20285 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17054) );
  AOI22_X1 U20286 ( .A1(n17197), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n16962), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17053) );
  AOI22_X1 U20287 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17052) );
  AOI22_X1 U20288 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17051) );
  NAND4_X1 U20289 ( .A1(n17054), .A2(n17053), .A3(n17052), .A4(n17051), .ZN(
        n17055) );
  NOR2_X1 U20290 ( .A1(n17056), .A2(n17055), .ZN(n17324) );
  OAI21_X1 U20291 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17058), .A(n17057), .ZN(
        n17059) );
  OAI21_X1 U20292 ( .B1(n17324), .B2(n17246), .A(n17059), .ZN(P3_U2683) );
  AOI22_X1 U20293 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17063) );
  AOI22_X1 U20294 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17062) );
  AOI22_X1 U20295 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17061) );
  AOI22_X1 U20296 ( .A1(n15700), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17060) );
  NAND4_X1 U20297 ( .A1(n17063), .A2(n17062), .A3(n17061), .A4(n17060), .ZN(
        n17069) );
  AOI22_X1 U20298 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n15711), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17067) );
  AOI22_X1 U20299 ( .A1(n9820), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n16962), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17066) );
  AOI22_X1 U20300 ( .A1(n17208), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17065) );
  AOI22_X1 U20301 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15713), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17064) );
  NAND4_X1 U20302 ( .A1(n17067), .A2(n17066), .A3(n17065), .A4(n17064), .ZN(
        n17068) );
  NOR2_X1 U20303 ( .A1(n17069), .A2(n17068), .ZN(n17329) );
  OAI21_X1 U20304 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17071), .A(n17070), .ZN(
        n17072) );
  AOI22_X1 U20305 ( .A1(n17261), .A2(n17329), .B1(n17072), .B2(n17246), .ZN(
        P3_U2684) );
  NAND2_X1 U20306 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17073), .ZN(n17086) );
  AOI22_X1 U20307 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15713), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17077) );
  AOI22_X1 U20308 ( .A1(n17197), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15711), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17076) );
  AOI22_X1 U20309 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17075) );
  AOI22_X1 U20310 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17074) );
  NAND4_X1 U20311 ( .A1(n17077), .A2(n17076), .A3(n17075), .A4(n17074), .ZN(
        n17083) );
  AOI22_X1 U20312 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17081) );
  AOI22_X1 U20313 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17080) );
  AOI22_X1 U20314 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9820), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17079) );
  AOI22_X1 U20315 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17078) );
  NAND4_X1 U20316 ( .A1(n17081), .A2(n17080), .A3(n17079), .A4(n17078), .ZN(
        n17082) );
  NOR2_X1 U20317 ( .A1(n17083), .A2(n17082), .ZN(n17334) );
  NAND2_X1 U20318 ( .A1(n18268), .A2(n17257), .ZN(n17263) );
  INV_X1 U20319 ( .A(n17263), .ZN(n17239) );
  NAND4_X1 U20320 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17097), .A3(n17239), 
        .A4(n17084), .ZN(n17085) );
  OAI221_X1 U20321 ( .B1(n17261), .B2(n17086), .C1(n17246), .C2(n17334), .A(
        n17085), .ZN(P3_U2685) );
  AOI22_X1 U20322 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17090) );
  AOI22_X1 U20323 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17089) );
  AOI22_X1 U20324 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n16962), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17088) );
  AOI22_X1 U20325 ( .A1(n15700), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17087) );
  NAND4_X1 U20326 ( .A1(n17090), .A2(n17089), .A3(n17088), .A4(n17087), .ZN(
        n17096) );
  AOI22_X1 U20327 ( .A1(n17197), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17094) );
  AOI22_X1 U20328 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17093) );
  AOI22_X1 U20329 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9820), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17092) );
  AOI22_X1 U20330 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n15699), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17091) );
  NAND4_X1 U20331 ( .A1(n17094), .A2(n17093), .A3(n17092), .A4(n17091), .ZN(
        n17095) );
  NOR2_X1 U20332 ( .A1(n17096), .A2(n17095), .ZN(n17339) );
  AND2_X1 U20333 ( .A1(n17097), .A2(n17239), .ZN(n17099) );
  NOR2_X1 U20334 ( .A1(n17351), .A2(n17097), .ZN(n17101) );
  NAND2_X1 U20335 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17257), .ZN(n17098) );
  OAI22_X1 U20336 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17099), .B1(n17101), 
        .B2(n17098), .ZN(n17100) );
  OAI21_X1 U20337 ( .B1(n17339), .B2(n17246), .A(n17100), .ZN(P3_U2686) );
  INV_X1 U20338 ( .A(n17101), .ZN(n17115) );
  INV_X1 U20339 ( .A(n17102), .ZN(n17138) );
  NAND2_X1 U20340 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17140), .ZN(n17114) );
  AOI22_X1 U20341 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17106) );
  AOI22_X1 U20342 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n15711), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17105) );
  AOI22_X1 U20343 ( .A1(n9820), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17197), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17104) );
  AOI22_X1 U20344 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n15700), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17103) );
  NAND4_X1 U20345 ( .A1(n17106), .A2(n17105), .A3(n17104), .A4(n17103), .ZN(
        n17112) );
  AOI22_X1 U20346 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17110) );
  AOI22_X1 U20347 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17109) );
  AOI22_X1 U20348 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17179), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17108) );
  AOI22_X1 U20349 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17019), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17107) );
  NAND4_X1 U20350 ( .A1(n17110), .A2(n17109), .A3(n17108), .A4(n17107), .ZN(
        n17111) );
  NOR2_X1 U20351 ( .A1(n17112), .A2(n17111), .ZN(n17345) );
  NAND2_X1 U20352 ( .A1(n17246), .A2(n17114), .ZN(n17126) );
  OAI222_X1 U20353 ( .A1(n17115), .A2(n17114), .B1(n17246), .B2(n17345), .C1(
        n17113), .C2(n17126), .ZN(P3_U2687) );
  AOI22_X1 U20354 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n9817), .B1(
        P3_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n17179), .ZN(n17119) );
  AOI22_X1 U20355 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17118) );
  AOI22_X1 U20356 ( .A1(n15700), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n16962), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17117) );
  AOI22_X1 U20357 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n17188), .B1(
        n15711), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17116) );
  NAND4_X1 U20358 ( .A1(n17119), .A2(n17118), .A3(n17117), .A4(n17116), .ZN(
        n17125) );
  AOI22_X1 U20359 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n17213), .ZN(n17123) );
  AOI22_X1 U20360 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n17197), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n17145), .ZN(n17122) );
  AOI22_X1 U20361 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n17143), .ZN(n17121) );
  AOI22_X1 U20362 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17019), .B1(
        n9820), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17120) );
  NAND4_X1 U20363 ( .A1(n17123), .A2(n17122), .A3(n17121), .A4(n17120), .ZN(
        n17124) );
  NOR2_X1 U20364 ( .A1(n17125), .A2(n17124), .ZN(n17349) );
  NOR2_X1 U20365 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17140), .ZN(n17127) );
  OAI22_X1 U20366 ( .A1(n17349), .A2(n17246), .B1(n17127), .B2(n17126), .ZN(
        P3_U2688) );
  AOI22_X1 U20367 ( .A1(n17197), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17131) );
  AOI22_X1 U20368 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17019), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17130) );
  AOI22_X1 U20369 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17129) );
  AOI22_X1 U20370 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17128) );
  NAND4_X1 U20371 ( .A1(n17131), .A2(n17130), .A3(n17129), .A4(n17128), .ZN(
        n17137) );
  AOI22_X1 U20372 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n15711), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17135) );
  AOI22_X1 U20373 ( .A1(n17208), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17179), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17134) );
  AOI22_X1 U20374 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17133) );
  AOI22_X1 U20375 ( .A1(n9820), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17132) );
  NAND4_X1 U20376 ( .A1(n17135), .A2(n17134), .A3(n17133), .A4(n17132), .ZN(
        n17136) );
  NOR2_X1 U20377 ( .A1(n17137), .A2(n17136), .ZN(n17353) );
  OAI21_X1 U20378 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17138), .A(n17246), .ZN(
        n17139) );
  OAI22_X1 U20379 ( .A1(n17353), .A2(n17246), .B1(n17140), .B2(n17139), .ZN(
        P3_U2689) );
  OAI21_X1 U20380 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17141), .A(n17246), .ZN(
        n17157) );
  AOI22_X1 U20381 ( .A1(n17179), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17155) );
  AOI22_X1 U20382 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16962), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17154) );
  AOI22_X1 U20383 ( .A1(n9820), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17197), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17142) );
  OAI21_X1 U20384 ( .B1(n9883), .B2(n17242), .A(n17142), .ZN(n17152) );
  AOI22_X1 U20385 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17150) );
  AOI22_X1 U20386 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17149) );
  AOI22_X1 U20387 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17148) );
  AOI22_X1 U20388 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17147) );
  NAND4_X1 U20389 ( .A1(n17150), .A2(n17149), .A3(n17148), .A4(n17147), .ZN(
        n17151) );
  AOI211_X1 U20390 ( .C1(n17196), .C2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A(
        n17152), .B(n17151), .ZN(n17153) );
  NAND3_X1 U20391 ( .A1(n17155), .A2(n17154), .A3(n17153), .ZN(n17361) );
  INV_X1 U20392 ( .A(n17361), .ZN(n17156) );
  OAI22_X1 U20393 ( .A1(n17158), .A2(n17157), .B1(n17156), .B2(n17246), .ZN(
        P3_U2691) );
  AOI22_X1 U20394 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17168) );
  AOI22_X1 U20395 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17167) );
  INV_X1 U20396 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17247) );
  AOI22_X1 U20397 ( .A1(n17208), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17159) );
  OAI21_X1 U20398 ( .B1(n9883), .B2(n17247), .A(n17159), .ZN(n17165) );
  AOI22_X1 U20399 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17163) );
  AOI22_X1 U20400 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17179), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17162) );
  AOI22_X1 U20401 ( .A1(n9820), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17161) );
  AOI22_X1 U20402 ( .A1(n17197), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16962), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17160) );
  NAND4_X1 U20403 ( .A1(n17163), .A2(n17162), .A3(n17161), .A4(n17160), .ZN(
        n17164) );
  AOI211_X1 U20404 ( .C1(n17214), .C2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A(
        n17165), .B(n17164), .ZN(n17166) );
  NAND3_X1 U20405 ( .A1(n17168), .A2(n17167), .A3(n17166), .ZN(n17365) );
  INV_X1 U20406 ( .A(n17365), .ZN(n17171) );
  OAI21_X1 U20407 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17187), .A(n17169), .ZN(
        n17170) );
  AOI22_X1 U20408 ( .A1(n17261), .A2(n17171), .B1(n17170), .B2(n17246), .ZN(
        P3_U2692) );
  AOI21_X1 U20409 ( .B1(n17172), .B2(n17204), .A(n17261), .ZN(n17173) );
  INV_X1 U20410 ( .A(n17173), .ZN(n17186) );
  AOI22_X1 U20411 ( .A1(n17208), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17178) );
  AOI22_X1 U20412 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n16962), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17177) );
  AOI22_X1 U20413 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17197), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17176) );
  AOI22_X1 U20414 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17175) );
  NAND4_X1 U20415 ( .A1(n17178), .A2(n17177), .A3(n17176), .A4(n17175), .ZN(
        n17185) );
  AOI22_X1 U20416 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17019), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17183) );
  AOI22_X1 U20417 ( .A1(n15700), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17179), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17182) );
  AOI22_X1 U20418 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17181) );
  AOI22_X1 U20419 ( .A1(n9820), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13703), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17180) );
  NAND4_X1 U20420 ( .A1(n17183), .A2(n17182), .A3(n17181), .A4(n17180), .ZN(
        n17184) );
  NOR2_X1 U20421 ( .A1(n17185), .A2(n17184), .ZN(n17368) );
  OAI22_X1 U20422 ( .A1(n17187), .A2(n17186), .B1(n17368), .B2(n17246), .ZN(
        P3_U2693) );
  AOI22_X1 U20423 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17193) );
  AOI22_X1 U20424 ( .A1(n17208), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17019), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17192) );
  AOI22_X1 U20425 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n15711), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17191) );
  AOI22_X1 U20426 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17179), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17190) );
  NAND4_X1 U20427 ( .A1(n17193), .A2(n17192), .A3(n17191), .A4(n17190), .ZN(
        n17203) );
  AOI22_X1 U20428 ( .A1(n15700), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17201) );
  AOI22_X1 U20429 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9820), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17200) );
  AOI22_X1 U20430 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17199) );
  AOI22_X1 U20431 ( .A1(n17197), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n16962), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17198) );
  NAND4_X1 U20432 ( .A1(n17201), .A2(n17200), .A3(n17199), .A4(n17198), .ZN(
        n17202) );
  NOR2_X1 U20433 ( .A1(n17203), .A2(n17202), .ZN(n17373) );
  OAI21_X1 U20434 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17226), .A(n17204), .ZN(
        n17205) );
  AOI22_X1 U20435 ( .A1(n17261), .A2(n17373), .B1(n17205), .B2(n17246), .ZN(
        P3_U2694) );
  AOI22_X1 U20436 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17212) );
  AOI22_X1 U20437 ( .A1(n15710), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17211) );
  AOI22_X1 U20438 ( .A1(n17208), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17210) );
  AOI22_X1 U20439 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15691), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17209) );
  NAND4_X1 U20440 ( .A1(n17212), .A2(n17211), .A3(n17210), .A4(n17209), .ZN(
        n17223) );
  AOI22_X1 U20441 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17221) );
  AOI22_X1 U20442 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n15711), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17220) );
  AOI22_X1 U20443 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15713), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17219) );
  AOI22_X1 U20444 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17218) );
  NAND4_X1 U20445 ( .A1(n17221), .A2(n17220), .A3(n17219), .A4(n17218), .ZN(
        n17222) );
  NOR2_X1 U20446 ( .A1(n17223), .A2(n17222), .ZN(n17380) );
  NOR3_X1 U20447 ( .A1(n17351), .A2(n17235), .A3(n17236), .ZN(n17231) );
  NAND2_X1 U20448 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17231), .ZN(n17227) );
  NOR2_X1 U20449 ( .A1(n17224), .A2(n17227), .ZN(n17230) );
  AOI21_X1 U20450 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17246), .A(n17230), .ZN(
        n17225) );
  OAI22_X1 U20451 ( .A1(n17380), .A2(n17246), .B1(n17226), .B2(n17225), .ZN(
        P3_U2695) );
  INV_X1 U20452 ( .A(n17227), .ZN(n17234) );
  AOI21_X1 U20453 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17246), .A(n17234), .ZN(
        n17229) );
  OAI22_X1 U20454 ( .A1(n17230), .A2(n17229), .B1(n17228), .B2(n17246), .ZN(
        P3_U2696) );
  AOI21_X1 U20455 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17246), .A(n17231), .ZN(
        n17233) );
  OAI22_X1 U20456 ( .A1(n17234), .A2(n17233), .B1(n17232), .B2(n17246), .ZN(
        P3_U2697) );
  INV_X1 U20457 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17238) );
  AOI22_X1 U20458 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17236), .B1(n17244), .B2(
        n17235), .ZN(n17237) );
  AOI22_X1 U20459 ( .A1(n17261), .A2(n17238), .B1(n17237), .B2(n17246), .ZN(
        P3_U2698) );
  NAND2_X1 U20460 ( .A1(n17240), .A2(n17239), .ZN(n17245) );
  NOR2_X1 U20461 ( .A1(n17241), .A2(n17245), .ZN(n17249) );
  AOI21_X1 U20462 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17246), .A(n17249), .ZN(
        n17243) );
  OAI22_X1 U20463 ( .A1(n17244), .A2(n17243), .B1(n17242), .B2(n17246), .ZN(
        P3_U2699) );
  INV_X1 U20464 ( .A(n17245), .ZN(n17253) );
  AOI21_X1 U20465 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17246), .A(n17253), .ZN(
        n17248) );
  OAI22_X1 U20466 ( .A1(n17249), .A2(n17248), .B1(n17247), .B2(n17246), .ZN(
        P3_U2700) );
  OAI21_X1 U20467 ( .B1(n17260), .B2(n17251), .A(n17250), .ZN(n17252) );
  INV_X1 U20468 ( .A(n17252), .ZN(n17255) );
  AOI221_X1 U20469 ( .B1(n17255), .B2(n17246), .C1(n17254), .C2(n17261), .A(
        n17253), .ZN(P3_U2701) );
  INV_X1 U20470 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17258) );
  OAI222_X1 U20471 ( .A1(n17263), .A2(n17259), .B1(n17258), .B2(n17257), .C1(
        n17256), .C2(n17246), .ZN(P3_U2702) );
  AOI22_X1 U20472 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17261), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17260), .ZN(n17262) );
  OAI21_X1 U20473 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17263), .A(n17262), .ZN(
        P3_U2703) );
  INV_X1 U20474 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17489) );
  INV_X1 U20475 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17424) );
  INV_X1 U20476 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17485) );
  INV_X1 U20477 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17483) );
  INV_X1 U20478 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17445) );
  INV_X1 U20479 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17504) );
  INV_X1 U20480 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17496) );
  INV_X1 U20481 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17461) );
  NAND4_X1 U20482 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(P3_EAX_REG_2__SCAN_IN), 
        .A3(P3_EAX_REG_6__SCAN_IN), .A4(P3_EAX_REG_5__SCAN_IN), .ZN(n17265) );
  NOR2_X1 U20483 ( .A1(n17461), .A2(n17265), .ZN(n17381) );
  INV_X1 U20484 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17510) );
  INV_X1 U20485 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17451) );
  NOR2_X1 U20486 ( .A1(n17510), .A2(n17451), .ZN(n17360) );
  AND2_X1 U20487 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17360), .ZN(n17356) );
  NAND4_X1 U20488 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .A3(n17376), .A4(n17356), .ZN(n17350) );
  NAND4_X1 U20489 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n17266)
         );
  NAND2_X1 U20490 ( .A1(n18268), .A2(n17305), .ZN(n17300) );
  NOR2_X1 U20491 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n9872), .ZN(n17268) );
  NAND2_X1 U20492 ( .A1(n17400), .A2(n9872), .ZN(n17275) );
  OAI21_X1 U20493 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17311), .A(n17275), .ZN(
        n17267) );
  AOI22_X1 U20494 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17268), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17267), .ZN(n17269) );
  OAI21_X1 U20495 ( .B1(n17270), .B2(n17316), .A(n17269), .ZN(P3_U2704) );
  INV_X1 U20496 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17417) );
  NOR2_X2 U20497 ( .A1(n17271), .A2(n17400), .ZN(n17341) );
  INV_X1 U20498 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n18261) );
  OAI22_X1 U20499 ( .A1(n17272), .A2(n17411), .B1(n18261), .B2(n17316), .ZN(
        n17273) );
  AOI21_X1 U20500 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17341), .A(n17273), .ZN(
        n17274) );
  OAI221_X1 U20501 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n9872), .C1(n17417), 
        .C2(n17275), .A(n17274), .ZN(P3_U2705) );
  AOI22_X1 U20502 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17341), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17340), .ZN(n17278) );
  OAI211_X1 U20503 ( .C1(n17276), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17400), .B(
        n9872), .ZN(n17277) );
  OAI211_X1 U20504 ( .C1(n17279), .C2(n17411), .A(n17278), .B(n17277), .ZN(
        P3_U2706) );
  INV_X1 U20505 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n18251) );
  AOI22_X1 U20506 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17341), .B1(n17383), .B2(
        n17280), .ZN(n17283) );
  OAI211_X1 U20507 ( .C1(n17284), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17400), .B(
        n17281), .ZN(n17282) );
  OAI211_X1 U20508 ( .C1(n17316), .C2(n18251), .A(n17283), .B(n17282), .ZN(
        P3_U2707) );
  AOI22_X1 U20509 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17341), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17340), .ZN(n17287) );
  AOI211_X1 U20510 ( .C1(n17489), .C2(n17290), .A(n17284), .B(n17406), .ZN(
        n17285) );
  INV_X1 U20511 ( .A(n17285), .ZN(n17286) );
  OAI211_X1 U20512 ( .C1(n17288), .C2(n17411), .A(n17287), .B(n17286), .ZN(
        P3_U2708) );
  INV_X1 U20513 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n17293) );
  AOI22_X1 U20514 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17341), .B1(n17383), .B2(
        n17289), .ZN(n17292) );
  OAI211_X1 U20515 ( .C1(n17294), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17400), .B(
        n17290), .ZN(n17291) );
  OAI211_X1 U20516 ( .C1(n17316), .C2(n17293), .A(n17292), .B(n17291), .ZN(
        P3_U2709) );
  AOI22_X1 U20517 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17341), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17340), .ZN(n17297) );
  AOI211_X1 U20518 ( .C1(n17424), .C2(n17301), .A(n17294), .B(n17406), .ZN(
        n17295) );
  INV_X1 U20519 ( .A(n17295), .ZN(n17296) );
  OAI211_X1 U20520 ( .C1(n17298), .C2(n17411), .A(n17297), .B(n17296), .ZN(
        P3_U2710) );
  INV_X1 U20521 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n18230) );
  AOI22_X1 U20522 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17341), .B1(n17383), .B2(
        n17299), .ZN(n17304) );
  OAI21_X1 U20523 ( .B1(n17485), .B2(n17406), .A(n17300), .ZN(n17302) );
  NAND2_X1 U20524 ( .A1(n17302), .A2(n17301), .ZN(n17303) );
  OAI211_X1 U20525 ( .C1(n17316), .C2(n18230), .A(n17304), .B(n17303), .ZN(
        P3_U2711) );
  AOI211_X1 U20526 ( .C1(n17483), .C2(n9890), .A(n17406), .B(n17305), .ZN(
        n17306) );
  AOI21_X1 U20527 ( .B1(n17340), .B2(BUF2_REG_23__SCAN_IN), .A(n17306), .ZN(
        n17308) );
  NAND2_X1 U20528 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17341), .ZN(n17307) );
  OAI211_X1 U20529 ( .C1(n17309), .C2(n17411), .A(n17308), .B(n17307), .ZN(
        P3_U2712) );
  INV_X1 U20530 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17430) );
  INV_X1 U20531 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17434) );
  INV_X1 U20532 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17441) );
  NAND2_X1 U20533 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17336), .ZN(n17335) );
  NAND2_X1 U20534 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17325), .ZN(n17321) );
  OR2_X1 U20535 ( .A1(n17430), .A2(n17321), .ZN(n17315) );
  AOI22_X1 U20536 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17340), .B1(n17383), .B2(
        n17310), .ZN(n17314) );
  NAND2_X1 U20537 ( .A1(n17400), .A2(n17321), .ZN(n17320) );
  OAI21_X1 U20538 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17311), .A(n17320), .ZN(
        n17312) );
  AOI22_X1 U20539 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17341), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17312), .ZN(n17313) );
  OAI211_X1 U20540 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n17315), .A(n17314), .B(
        n17313), .ZN(P3_U2713) );
  INV_X1 U20541 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n19264) );
  OAI22_X1 U20542 ( .A1(n17317), .A2(n17411), .B1(n19264), .B2(n17316), .ZN(
        n17318) );
  AOI21_X1 U20543 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17341), .A(n17318), .ZN(
        n17319) );
  OAI221_X1 U20544 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17321), .C1(n17430), 
        .C2(n17320), .A(n17319), .ZN(P3_U2714) );
  AOI22_X1 U20545 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17341), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17340), .ZN(n17323) );
  OAI211_X1 U20546 ( .C1(n17325), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17400), .B(
        n17321), .ZN(n17322) );
  OAI211_X1 U20547 ( .C1(n17324), .C2(n17411), .A(n17323), .B(n17322), .ZN(
        P3_U2715) );
  AOI22_X1 U20548 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17341), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17340), .ZN(n17328) );
  AOI211_X1 U20549 ( .C1(n17434), .C2(n17330), .A(n17325), .B(n17406), .ZN(
        n17326) );
  INV_X1 U20550 ( .A(n17326), .ZN(n17327) );
  OAI211_X1 U20551 ( .C1(n17329), .C2(n17411), .A(n17328), .B(n17327), .ZN(
        P3_U2716) );
  AOI22_X1 U20552 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17341), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17340), .ZN(n17333) );
  OAI211_X1 U20553 ( .C1(n17331), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17400), .B(
        n17330), .ZN(n17332) );
  OAI211_X1 U20554 ( .C1(n17334), .C2(n17411), .A(n17333), .B(n17332), .ZN(
        P3_U2717) );
  AOI22_X1 U20555 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17341), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17340), .ZN(n17338) );
  OAI211_X1 U20556 ( .C1(n17336), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17400), .B(
        n17335), .ZN(n17337) );
  OAI211_X1 U20557 ( .C1(n17339), .C2(n17411), .A(n17338), .B(n17337), .ZN(
        P3_U2718) );
  AOI22_X1 U20558 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17341), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17340), .ZN(n17344) );
  INV_X1 U20559 ( .A(n17346), .ZN(n17342) );
  OAI221_X1 U20560 ( .B1(n17342), .B2(P3_EAX_REG_16__SCAN_IN), .C1(n17346), 
        .C2(n17441), .A(n17400), .ZN(n17343) );
  OAI211_X1 U20561 ( .C1(n17345), .C2(n17411), .A(n17344), .B(n17343), .ZN(
        P3_U2719) );
  OAI211_X1 U20562 ( .C1(P3_EAX_REG_15__SCAN_IN), .C2(n17355), .A(n17400), .B(
        n17346), .ZN(n17348) );
  NAND2_X1 U20563 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17409), .ZN(n17347) );
  OAI211_X1 U20564 ( .C1(n17349), .C2(n17411), .A(n17348), .B(n17347), .ZN(
        P3_U2720) );
  INV_X1 U20565 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n17519) );
  OAI22_X1 U20566 ( .A1(n17351), .A2(n17350), .B1(n17445), .B2(n17406), .ZN(
        n17352) );
  INV_X1 U20567 ( .A(n17352), .ZN(n17354) );
  OAI222_X1 U20568 ( .A1(n17405), .A2(n17519), .B1(n17355), .B2(n17354), .C1(
        n17411), .C2(n17353), .ZN(P3_U2721) );
  INV_X1 U20569 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17453) );
  NAND2_X1 U20570 ( .A1(n18268), .A2(n17376), .ZN(n17371) );
  NAND2_X1 U20571 ( .A1(n17356), .A2(n17375), .ZN(n17359) );
  INV_X1 U20572 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17514) );
  NAND2_X1 U20573 ( .A1(n17400), .A2(n17359), .ZN(n17363) );
  AOI22_X1 U20574 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17409), .B1(n17383), .B2(
        n17357), .ZN(n17358) );
  OAI221_X1 U20575 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17359), .C1(n17514), 
        .C2(n17363), .A(n17358), .ZN(P3_U2722) );
  NAND2_X1 U20576 ( .A1(n17360), .A2(n17375), .ZN(n17364) );
  INV_X1 U20577 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17448) );
  AOI22_X1 U20578 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17409), .B1(n17383), .B2(
        n17361), .ZN(n17362) );
  OAI221_X1 U20579 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17364), .C1(n17448), 
        .C2(n17363), .A(n17362), .ZN(P3_U2723) );
  NAND2_X1 U20580 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17375), .ZN(n17367) );
  NAND2_X1 U20581 ( .A1(n17400), .A2(n17367), .ZN(n17370) );
  AOI22_X1 U20582 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17409), .B1(n17383), .B2(
        n17365), .ZN(n17366) );
  OAI221_X1 U20583 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17367), .C1(n17510), 
        .C2(n17370), .A(n17366), .ZN(P3_U2724) );
  INV_X1 U20584 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17508) );
  NOR2_X1 U20585 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17375), .ZN(n17369) );
  OAI222_X1 U20586 ( .A1(n17405), .A2(n17508), .B1(n17370), .B2(n17369), .C1(
        n17411), .C2(n17368), .ZN(P3_U2725) );
  INV_X1 U20587 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17506) );
  OAI21_X1 U20588 ( .B1(n17453), .B2(n17406), .A(n17371), .ZN(n17372) );
  INV_X1 U20589 ( .A(n17372), .ZN(n17374) );
  OAI222_X1 U20590 ( .A1(n17405), .A2(n17506), .B1(n17375), .B2(n17374), .C1(
        n17411), .C2(n17373), .ZN(P3_U2726) );
  AOI211_X1 U20591 ( .C1(n17504), .C2(n17377), .A(n17406), .B(n17376), .ZN(
        n17378) );
  AOI21_X1 U20592 ( .B1(n17409), .B2(BUF2_REG_8__SCAN_IN), .A(n17378), .ZN(
        n17379) );
  OAI21_X1 U20593 ( .B1(n17380), .B2(n17411), .A(n17379), .ZN(P3_U2727) );
  NAND3_X1 U20594 ( .A1(n18268), .A2(n9929), .A3(n17381), .ZN(n17386) );
  NAND2_X1 U20595 ( .A1(n17386), .A2(P3_EAX_REG_7__SCAN_IN), .ZN(n17385) );
  AOI22_X1 U20596 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17409), .B1(n17383), .B2(
        n17382), .ZN(n17384) );
  OAI221_X1 U20597 ( .B1(n17386), .B2(P3_EAX_REG_7__SCAN_IN), .C1(n17385), 
        .C2(n17406), .A(n17384), .ZN(P3_U2728) );
  INV_X1 U20598 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18262) );
  INV_X1 U20599 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17459) );
  INV_X1 U20600 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17463) );
  NAND3_X1 U20601 ( .A1(n18268), .A2(n9929), .A3(P3_EAX_REG_2__SCAN_IN), .ZN(
        n17396) );
  NOR2_X1 U20602 ( .A1(n17463), .A2(n17396), .ZN(n17398) );
  NAND2_X1 U20603 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17398), .ZN(n17389) );
  NOR2_X1 U20604 ( .A1(n17459), .A2(n17389), .ZN(n17391) );
  AOI21_X1 U20605 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17400), .A(n17391), .ZN(
        n17388) );
  INV_X1 U20606 ( .A(n17386), .ZN(n17387) );
  OAI222_X1 U20607 ( .A1(n17405), .A2(n18262), .B1(n17388), .B2(n17387), .C1(
        n17411), .C2(n17816), .ZN(P3_U2729) );
  INV_X1 U20608 ( .A(n17389), .ZN(n17394) );
  AOI21_X1 U20609 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17400), .A(n17394), .ZN(
        n17392) );
  OAI222_X1 U20610 ( .A1(n17405), .A2(n18257), .B1(n17392), .B2(n17391), .C1(
        n17411), .C2(n17390), .ZN(P3_U2730) );
  INV_X1 U20611 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18252) );
  AOI21_X1 U20612 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17400), .A(n17398), .ZN(
        n17395) );
  OAI222_X1 U20613 ( .A1(n17405), .A2(n18252), .B1(n17395), .B2(n17394), .C1(
        n17411), .C2(n17393), .ZN(P3_U2731) );
  INV_X1 U20614 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18247) );
  INV_X1 U20615 ( .A(n17396), .ZN(n17403) );
  AOI21_X1 U20616 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17400), .A(n17403), .ZN(
        n17399) );
  OAI222_X1 U20617 ( .A1(n17405), .A2(n18247), .B1(n17399), .B2(n17398), .C1(
        n17411), .C2(n17397), .ZN(P3_U2732) );
  INV_X1 U20618 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18243) );
  AOI22_X1 U20619 ( .A1(n18268), .A2(n9929), .B1(P3_EAX_REG_2__SCAN_IN), .B2(
        n17400), .ZN(n17404) );
  INV_X1 U20620 ( .A(n17401), .ZN(n17402) );
  OAI222_X1 U20621 ( .A1(n17405), .A2(n18243), .B1(n17404), .B2(n17403), .C1(
        n17411), .C2(n17402), .ZN(P3_U2733) );
  AOI211_X1 U20622 ( .C1(n17496), .C2(n17407), .A(n17406), .B(n9929), .ZN(
        n17408) );
  AOI21_X1 U20623 ( .B1(n17409), .B2(BUF2_REG_1__SCAN_IN), .A(n17408), .ZN(
        n17410) );
  OAI21_X1 U20624 ( .B1(n17412), .B2(n17411), .A(n17410), .ZN(P3_U2734) );
  NAND2_X1 U20625 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17722), .ZN(n18883) );
  INV_X2 U20626 ( .A(n18883), .ZN(n17468) );
  AND2_X1 U20627 ( .A1(n17438), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U20628 ( .A1(n17442), .A2(n17415), .ZN(n17440) );
  AOI22_X1 U20629 ( .A1(n17468), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(n17467), .ZN(n17416) );
  OAI21_X1 U20630 ( .B1(n17417), .B2(n17440), .A(n17416), .ZN(P3_U2737) );
  INV_X1 U20631 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17492) );
  AOI22_X1 U20632 ( .A1(n17468), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17467), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17418) );
  OAI21_X1 U20633 ( .B1(n17492), .B2(n17440), .A(n17418), .ZN(P3_U2738) );
  AOI22_X1 U20634 ( .A1(n17468), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17467), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17419) );
  OAI21_X1 U20635 ( .B1(n10045), .B2(n17440), .A(n17419), .ZN(P3_U2739) );
  AOI22_X1 U20636 ( .A1(n17468), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17438), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17420) );
  OAI21_X1 U20637 ( .B1(n17489), .B2(n17440), .A(n17420), .ZN(P3_U2740) );
  INV_X1 U20638 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17422) );
  AOI22_X1 U20639 ( .A1(n17468), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17438), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17421) );
  OAI21_X1 U20640 ( .B1(n17422), .B2(n17440), .A(n17421), .ZN(P3_U2741) );
  AOI22_X1 U20641 ( .A1(n17468), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17467), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17423) );
  OAI21_X1 U20642 ( .B1(n17424), .B2(n17440), .A(n17423), .ZN(P3_U2742) );
  AOI22_X1 U20643 ( .A1(n17468), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17438), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17425) );
  OAI21_X1 U20644 ( .B1(n17485), .B2(n17440), .A(n17425), .ZN(P3_U2743) );
  AOI22_X1 U20645 ( .A1(n17468), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17467), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17426) );
  OAI21_X1 U20646 ( .B1(n17483), .B2(n17440), .A(n17426), .ZN(P3_U2744) );
  INV_X1 U20647 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17428) );
  AOI22_X1 U20648 ( .A1(n17468), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17438), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17427) );
  OAI21_X1 U20649 ( .B1(n17428), .B2(n17440), .A(n17427), .ZN(P3_U2745) );
  AOI22_X1 U20650 ( .A1(n17468), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17438), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17429) );
  OAI21_X1 U20651 ( .B1(n17430), .B2(n17440), .A(n17429), .ZN(P3_U2746) );
  INV_X1 U20652 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17432) );
  AOI22_X1 U20653 ( .A1(n17468), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17438), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17431) );
  OAI21_X1 U20654 ( .B1(n17432), .B2(n17440), .A(n17431), .ZN(P3_U2747) );
  AOI22_X1 U20655 ( .A1(n17468), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17438), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17433) );
  OAI21_X1 U20656 ( .B1(n17434), .B2(n17440), .A(n17433), .ZN(P3_U2748) );
  INV_X1 U20657 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17436) );
  AOI22_X1 U20658 ( .A1(n17468), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17438), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17435) );
  OAI21_X1 U20659 ( .B1(n17436), .B2(n17440), .A(n17435), .ZN(P3_U2749) );
  INV_X1 U20660 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17476) );
  AOI22_X1 U20661 ( .A1(n17468), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17438), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17437) );
  OAI21_X1 U20662 ( .B1(n17476), .B2(n17440), .A(n17437), .ZN(P3_U2750) );
  AOI22_X1 U20663 ( .A1(n17468), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17438), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17439) );
  OAI21_X1 U20664 ( .B1(n17441), .B2(n17440), .A(n17439), .ZN(P3_U2751) );
  INV_X1 U20665 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17524) );
  AOI22_X1 U20666 ( .A1(n17468), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17467), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17443) );
  OAI21_X1 U20667 ( .B1(n17524), .B2(n17470), .A(n17443), .ZN(P3_U2752) );
  AOI22_X1 U20668 ( .A1(n17468), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17467), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17444) );
  OAI21_X1 U20669 ( .B1(n17445), .B2(n17470), .A(n17444), .ZN(P3_U2753) );
  AOI22_X1 U20670 ( .A1(n17468), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17467), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17446) );
  OAI21_X1 U20671 ( .B1(n17514), .B2(n17470), .A(n17446), .ZN(P3_U2754) );
  AOI22_X1 U20672 ( .A1(n17468), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17467), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17447) );
  OAI21_X1 U20673 ( .B1(n17448), .B2(n17470), .A(n17447), .ZN(P3_U2755) );
  AOI22_X1 U20674 ( .A1(n17468), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17467), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17449) );
  OAI21_X1 U20675 ( .B1(n17510), .B2(n17470), .A(n17449), .ZN(P3_U2756) );
  AOI22_X1 U20676 ( .A1(n17468), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17467), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17450) );
  OAI21_X1 U20677 ( .B1(n17451), .B2(n17470), .A(n17450), .ZN(P3_U2757) );
  AOI22_X1 U20678 ( .A1(n17468), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17467), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17452) );
  OAI21_X1 U20679 ( .B1(n17453), .B2(n17470), .A(n17452), .ZN(P3_U2758) );
  AOI22_X1 U20680 ( .A1(n17468), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17467), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17454) );
  OAI21_X1 U20681 ( .B1(n17504), .B2(n17470), .A(n17454), .ZN(P3_U2759) );
  AOI22_X1 U20682 ( .A1(n17468), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17467), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17455) );
  OAI21_X1 U20683 ( .B1(n10051), .B2(n17470), .A(n17455), .ZN(P3_U2760) );
  INV_X1 U20684 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17457) );
  AOI22_X1 U20685 ( .A1(n17468), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17467), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17456) );
  OAI21_X1 U20686 ( .B1(n17457), .B2(n17470), .A(n17456), .ZN(P3_U2761) );
  AOI22_X1 U20687 ( .A1(n17468), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17467), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17458) );
  OAI21_X1 U20688 ( .B1(n17459), .B2(n17470), .A(n17458), .ZN(P3_U2762) );
  AOI22_X1 U20689 ( .A1(n17468), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17467), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17460) );
  OAI21_X1 U20690 ( .B1(n17461), .B2(n17470), .A(n17460), .ZN(P3_U2763) );
  AOI22_X1 U20691 ( .A1(n17468), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17467), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17462) );
  OAI21_X1 U20692 ( .B1(n17463), .B2(n17470), .A(n17462), .ZN(P3_U2764) );
  INV_X1 U20693 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17465) );
  AOI22_X1 U20694 ( .A1(n17468), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17467), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17464) );
  OAI21_X1 U20695 ( .B1(n17465), .B2(n17470), .A(n17464), .ZN(P3_U2765) );
  AOI22_X1 U20696 ( .A1(n17468), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17467), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17466) );
  OAI21_X1 U20697 ( .B1(n17496), .B2(n17470), .A(n17466), .ZN(P3_U2766) );
  AOI22_X1 U20698 ( .A1(n17468), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17467), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17469) );
  OAI21_X1 U20699 ( .B1(n10049), .B2(n17470), .A(n17469), .ZN(P3_U2767) );
  INV_X1 U20700 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18231) );
  OAI211_X1 U20701 ( .C1(n18890), .C2(n18889), .A(n17471), .B(n17473), .ZN(
        n17520) );
  NAND2_X1 U20702 ( .A1(n17473), .A2(n17472), .ZN(n17523) );
  AOI22_X1 U20703 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17516), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17515), .ZN(n17474) );
  OAI21_X1 U20704 ( .B1(n18231), .B2(n17518), .A(n17474), .ZN(P3_U2768) );
  AOI22_X1 U20705 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17521), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17515), .ZN(n17475) );
  OAI21_X1 U20706 ( .B1(n17476), .B2(n17523), .A(n17475), .ZN(P3_U2769) );
  AOI22_X1 U20707 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17516), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17515), .ZN(n17477) );
  OAI21_X1 U20708 ( .B1(n18243), .B2(n17518), .A(n17477), .ZN(P3_U2770) );
  AOI22_X1 U20709 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17516), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17515), .ZN(n17478) );
  OAI21_X1 U20710 ( .B1(n18247), .B2(n17518), .A(n17478), .ZN(P3_U2771) );
  AOI22_X1 U20711 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17516), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17515), .ZN(n17479) );
  OAI21_X1 U20712 ( .B1(n18252), .B2(n17518), .A(n17479), .ZN(P3_U2772) );
  AOI22_X1 U20713 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17516), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17515), .ZN(n17480) );
  OAI21_X1 U20714 ( .B1(n18257), .B2(n17518), .A(n17480), .ZN(P3_U2773) );
  AOI22_X1 U20715 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17516), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17515), .ZN(n17481) );
  OAI21_X1 U20716 ( .B1(n18262), .B2(n17518), .A(n17481), .ZN(P3_U2774) );
  AOI22_X1 U20717 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17521), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17515), .ZN(n17482) );
  OAI21_X1 U20718 ( .B1(n17483), .B2(n17523), .A(n17482), .ZN(P3_U2775) );
  AOI22_X1 U20719 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17521), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17515), .ZN(n17484) );
  OAI21_X1 U20720 ( .B1(n17485), .B2(n17523), .A(n17484), .ZN(P3_U2776) );
  AOI22_X1 U20721 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17516), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17515), .ZN(n17486) );
  OAI21_X1 U20722 ( .B1(n17506), .B2(n17518), .A(n17486), .ZN(P3_U2777) );
  AOI22_X1 U20723 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17516), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17515), .ZN(n17487) );
  OAI21_X1 U20724 ( .B1(n17508), .B2(n17518), .A(n17487), .ZN(P3_U2778) );
  AOI22_X1 U20725 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17521), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17515), .ZN(n17488) );
  OAI21_X1 U20726 ( .B1(n17489), .B2(n17523), .A(n17488), .ZN(P3_U2779) );
  INV_X1 U20727 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17512) );
  AOI22_X1 U20728 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17516), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17515), .ZN(n17490) );
  OAI21_X1 U20729 ( .B1(n17512), .B2(n17518), .A(n17490), .ZN(P3_U2780) );
  AOI22_X1 U20730 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17521), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17515), .ZN(n17491) );
  OAI21_X1 U20731 ( .B1(n17492), .B2(n17523), .A(n17491), .ZN(P3_U2781) );
  AOI22_X1 U20732 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17516), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17515), .ZN(n17493) );
  OAI21_X1 U20733 ( .B1(n17519), .B2(n17518), .A(n17493), .ZN(P3_U2782) );
  AOI22_X1 U20734 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17516), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17515), .ZN(n17494) );
  OAI21_X1 U20735 ( .B1(n18231), .B2(n17518), .A(n17494), .ZN(P3_U2783) );
  AOI22_X1 U20736 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17521), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17515), .ZN(n17495) );
  OAI21_X1 U20737 ( .B1(n17496), .B2(n17523), .A(n17495), .ZN(P3_U2784) );
  AOI22_X1 U20738 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17516), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17515), .ZN(n17497) );
  OAI21_X1 U20739 ( .B1(n18243), .B2(n17518), .A(n17497), .ZN(P3_U2785) );
  AOI22_X1 U20740 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17516), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17520), .ZN(n17498) );
  OAI21_X1 U20741 ( .B1(n18247), .B2(n17518), .A(n17498), .ZN(P3_U2786) );
  AOI22_X1 U20742 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17516), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17520), .ZN(n17499) );
  OAI21_X1 U20743 ( .B1(n18252), .B2(n17518), .A(n17499), .ZN(P3_U2787) );
  AOI22_X1 U20744 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17516), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17520), .ZN(n17500) );
  OAI21_X1 U20745 ( .B1(n18257), .B2(n17518), .A(n17500), .ZN(P3_U2788) );
  AOI22_X1 U20746 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17516), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17520), .ZN(n17501) );
  OAI21_X1 U20747 ( .B1(n18262), .B2(n17518), .A(n17501), .ZN(P3_U2789) );
  AOI22_X1 U20748 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17521), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17520), .ZN(n17502) );
  OAI21_X1 U20749 ( .B1(n10051), .B2(n17523), .A(n17502), .ZN(P3_U2790) );
  AOI22_X1 U20750 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17521), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17520), .ZN(n17503) );
  OAI21_X1 U20751 ( .B1(n17504), .B2(n17523), .A(n17503), .ZN(P3_U2791) );
  AOI22_X1 U20752 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17516), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17520), .ZN(n17505) );
  OAI21_X1 U20753 ( .B1(n17506), .B2(n17518), .A(n17505), .ZN(P3_U2792) );
  AOI22_X1 U20754 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17516), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17515), .ZN(n17507) );
  OAI21_X1 U20755 ( .B1(n17508), .B2(n17518), .A(n17507), .ZN(P3_U2793) );
  AOI22_X1 U20756 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17521), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17520), .ZN(n17509) );
  OAI21_X1 U20757 ( .B1(n17510), .B2(n17523), .A(n17509), .ZN(P3_U2794) );
  AOI22_X1 U20758 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17516), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17515), .ZN(n17511) );
  OAI21_X1 U20759 ( .B1(n17512), .B2(n17518), .A(n17511), .ZN(P3_U2795) );
  AOI22_X1 U20760 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17521), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17520), .ZN(n17513) );
  OAI21_X1 U20761 ( .B1(n17514), .B2(n17523), .A(n17513), .ZN(P3_U2796) );
  AOI22_X1 U20762 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17516), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17515), .ZN(n17517) );
  OAI21_X1 U20763 ( .B1(n17519), .B2(n17518), .A(n17517), .ZN(P3_U2797) );
  AOI22_X1 U20764 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17521), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17520), .ZN(n17522) );
  OAI21_X1 U20765 ( .B1(n17524), .B2(n17523), .A(n17522), .ZN(P3_U2798) );
  AOI21_X1 U20766 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n9930), .A(
        n17895), .ZN(n17525) );
  AOI211_X1 U20767 ( .C1(n17846), .C2(n17534), .A(n17844), .B(n17525), .ZN(
        n17559) );
  OAI21_X1 U20768 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17633), .A(
        n17559), .ZN(n17545) );
  AOI22_X1 U20769 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17545), .B1(
        n17735), .B2(n17526), .ZN(n17539) );
  NAND2_X1 U20770 ( .A1(n17803), .A2(n17899), .ZN(n17604) );
  INV_X1 U20771 ( .A(n17604), .ZN(n17631) );
  OAI22_X1 U20772 ( .A1(n17527), .A2(n17803), .B1(n17908), .B2(n17899), .ZN(
        n17555) );
  NOR2_X1 U20773 ( .A1(n15781), .A2(n17555), .ZN(n17529) );
  NOR3_X1 U20774 ( .A1(n17631), .A2(n17529), .A3(n17528), .ZN(n17532) );
  NOR2_X1 U20775 ( .A1(n17646), .A2(n17534), .ZN(n17547) );
  OAI211_X1 U20776 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17547), .B(n17535), .ZN(n17536) );
  NAND4_X1 U20777 ( .A1(n17539), .A2(n17538), .A3(n17537), .A4(n17536), .ZN(
        P3_U2802) );
  NAND2_X1 U20778 ( .A1(n10181), .A2(n17541), .ZN(n17542) );
  XOR2_X1 U20779 ( .A(n17760), .B(n17542), .Z(n17916) );
  OAI22_X1 U20780 ( .A1(n18201), .A2(n18813), .B1(n17728), .B2(n17543), .ZN(
        n17544) );
  AOI221_X1 U20781 ( .B1(n17547), .B2(n17546), .C1(n17545), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n17544), .ZN(n17550) );
  AOI22_X1 U20782 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17555), .B1(
        n17548), .B2(n15781), .ZN(n17549) );
  OAI211_X1 U20783 ( .C1(n17916), .C2(n17773), .A(n17550), .B(n17549), .ZN(
        P3_U2803) );
  AOI21_X1 U20784 ( .B1(n9930), .B2(n18616), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17558) );
  NAND2_X1 U20785 ( .A1(n17728), .A2(n17633), .ZN(n17855) );
  AOI22_X1 U20786 ( .A1(n18218), .A2(P3_REIP_REG_26__SCAN_IN), .B1(n17551), 
        .B2(n17855), .ZN(n17557) );
  AOI21_X1 U20787 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17553), .A(
        n17552), .ZN(n17917) );
  INV_X1 U20788 ( .A(n17925), .ZN(n17928) );
  NAND3_X1 U20789 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17928), .A3(
        n17923), .ZN(n17920) );
  OAI22_X1 U20790 ( .A1(n17917), .A2(n17773), .B1(n17596), .B2(n17920), .ZN(
        n17554) );
  AOI21_X1 U20791 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17555), .A(
        n17554), .ZN(n17556) );
  OAI211_X1 U20792 ( .C1(n17559), .C2(n17558), .A(n17557), .B(n17556), .ZN(
        P3_U2804) );
  AND2_X1 U20793 ( .A1(n17569), .A2(n18616), .ZN(n17560) );
  AOI211_X1 U20794 ( .C1(n17722), .C2(n17561), .A(n17844), .B(n17560), .ZN(
        n17592) );
  OAI21_X1 U20795 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17633), .A(
        n17592), .ZN(n17575) );
  AOI22_X1 U20796 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17575), .B1(
        n17735), .B2(n17562), .ZN(n17574) );
  XOR2_X1 U20797 ( .A(n17563), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17935) );
  XOR2_X1 U20798 ( .A(n17564), .B(n17929), .Z(n17934) );
  OAI21_X1 U20799 ( .B1(n17760), .B2(n17566), .A(n17565), .ZN(n17567) );
  XOR2_X1 U20800 ( .A(n17567), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17940) );
  OAI22_X1 U20801 ( .A1(n17803), .A2(n17934), .B1(n17773), .B2(n17940), .ZN(
        n17568) );
  AOI21_X1 U20802 ( .B1(n17800), .B2(n17935), .A(n17568), .ZN(n17573) );
  NOR2_X1 U20803 ( .A1(n18201), .A2(n18809), .ZN(n17933) );
  INV_X1 U20804 ( .A(n17933), .ZN(n17572) );
  NOR2_X1 U20805 ( .A1(n17646), .A2(n17569), .ZN(n17577) );
  OAI211_X1 U20806 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17577), .B(n17570), .ZN(n17571) );
  NAND4_X1 U20807 ( .A1(n17574), .A2(n17573), .A3(n17572), .A4(n17571), .ZN(
        P3_U2805) );
  NOR2_X1 U20808 ( .A1(n18201), .A2(n18807), .ZN(n17941) );
  AOI221_X1 U20809 ( .B1(n17577), .B2(n17576), .C1(n17575), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17941), .ZN(n17584) );
  NOR2_X1 U20810 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17578), .ZN(
        n17942) );
  AOI22_X1 U20811 ( .A1(n17745), .A2(n17943), .B1(n17800), .B2(n17944), .ZN(
        n17595) );
  AOI21_X1 U20812 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17580), .A(
        n17579), .ZN(n17952) );
  OAI22_X1 U20813 ( .A1(n17595), .A2(n17581), .B1(n17952), .B2(n17773), .ZN(
        n17582) );
  AOI21_X1 U20814 ( .B1(n17610), .B2(n17942), .A(n17582), .ZN(n17583) );
  OAI211_X1 U20815 ( .C1(n17728), .C2(n17585), .A(n17584), .B(n17583), .ZN(
        P3_U2806) );
  INV_X1 U20816 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17953) );
  INV_X1 U20817 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17608) );
  OAI21_X1 U20818 ( .B1(n17665), .B2(n17901), .A(n17606), .ZN(n17586) );
  OAI211_X1 U20819 ( .C1(n17798), .C2(n17608), .A(n17586), .B(n17628), .ZN(
        n17587) );
  XOR2_X1 U20820 ( .A(n17953), .B(n17587), .Z(n17957) );
  AOI21_X1 U20821 ( .B1(n16588), .B2(n18616), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17591) );
  INV_X1 U20822 ( .A(n17633), .ZN(n17589) );
  OAI21_X1 U20823 ( .B1(n17735), .B2(n17589), .A(n17588), .ZN(n17590) );
  NAND2_X1 U20824 ( .A1(n18218), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17958) );
  OAI211_X1 U20825 ( .C1(n17592), .C2(n17591), .A(n17590), .B(n17958), .ZN(
        n17593) );
  AOI21_X1 U20826 ( .B1(n17799), .B2(n17957), .A(n17593), .ZN(n17594) );
  OAI221_X1 U20827 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17596), 
        .C1(n17953), .C2(n17595), .A(n17594), .ZN(P3_U2807) );
  OAI21_X1 U20828 ( .B1(n17597), .B2(n17895), .A(n17894), .ZN(n17598) );
  AOI21_X1 U20829 ( .B1(n17846), .B2(n17611), .A(n17598), .ZN(n17637) );
  OAI21_X1 U20830 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17633), .A(
        n17637), .ZN(n17619) );
  AOI22_X1 U20831 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17619), .B1(
        n17735), .B2(n17599), .ZN(n17615) );
  INV_X1 U20832 ( .A(n17600), .ZN(n17601) );
  NOR2_X1 U20833 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17601), .ZN(
        n17961) );
  INV_X1 U20834 ( .A(n17602), .ZN(n17963) );
  AOI22_X1 U20835 ( .A1(n17963), .A2(n17745), .B1(n18036), .B2(n17800), .ZN(
        n17692) );
  INV_X1 U20836 ( .A(n17692), .ZN(n17603) );
  AOI21_X1 U20837 ( .B1(n17967), .B2(n17604), .A(n17603), .ZN(n17627) );
  AOI221_X1 U20838 ( .B1(n17680), .B2(n17606), .C1(n17967), .C2(n17606), .A(
        n17605), .ZN(n17607) );
  XOR2_X1 U20839 ( .A(n17608), .B(n17607), .Z(n17960) );
  OAI22_X1 U20840 ( .A1(n17627), .A2(n17608), .B1(n17773), .B2(n17960), .ZN(
        n17609) );
  AOI21_X1 U20841 ( .B1(n17610), .B2(n17961), .A(n17609), .ZN(n17614) );
  NAND2_X1 U20842 ( .A1(n18218), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17975) );
  NOR2_X1 U20843 ( .A1(n17646), .A2(n17611), .ZN(n17621) );
  OAI211_X1 U20844 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17621), .B(n17612), .ZN(n17613) );
  NAND4_X1 U20845 ( .A1(n17615), .A2(n17614), .A3(n17975), .A4(n17613), .ZN(
        P3_U2808) );
  INV_X1 U20846 ( .A(n17616), .ZN(n17617) );
  OAI22_X1 U20847 ( .A1(n18201), .A2(n18801), .B1(n17728), .B2(n17617), .ZN(
        n17618) );
  AOI221_X1 U20848 ( .B1(n17621), .B2(n17620), .C1(n17619), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17618), .ZN(n17626) );
  INV_X1 U20849 ( .A(n17970), .ZN(n17979) );
  AND3_X1 U20850 ( .A1(n17798), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17622), .ZN(n17642) );
  AOI22_X1 U20851 ( .A1(n17979), .A2(n17642), .B1(n17665), .B2(n17623), .ZN(
        n17624) );
  XOR2_X1 U20852 ( .A(n17968), .B(n17624), .Z(n17983) );
  NOR2_X1 U20853 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17970), .ZN(
        n17982) );
  NAND2_X1 U20854 ( .A1(n17662), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17977) );
  NOR2_X1 U20855 ( .A1(n17693), .A2(n17977), .ZN(n17653) );
  AOI22_X1 U20856 ( .A1(n17799), .A2(n17983), .B1(n17982), .B2(n17653), .ZN(
        n17625) );
  OAI211_X1 U20857 ( .C1(n17627), .C2(n17968), .A(n17626), .B(n17625), .ZN(
        P3_U2809) );
  OAI221_X1 U20858 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17663), 
        .C1(n17999), .C2(n17642), .A(n17628), .ZN(n17629) );
  XOR2_X1 U20859 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17629), .Z(
        n17998) );
  NOR2_X1 U20860 ( .A1(n17999), .A2(n17977), .ZN(n17630) );
  INV_X1 U20861 ( .A(n17630), .ZN(n17989) );
  NOR2_X1 U20862 ( .A1(n17693), .A2(n17989), .ZN(n17640) );
  INV_X1 U20863 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17639) );
  OAI21_X1 U20864 ( .B1(n17631), .B2(n17630), .A(n17692), .ZN(n17652) );
  AOI21_X1 U20865 ( .B1(n17632), .B2(n18616), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17636) );
  OAI21_X1 U20866 ( .B1(n17735), .B2(n17589), .A(n17634), .ZN(n17635) );
  NAND2_X1 U20867 ( .A1(n18218), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n17996) );
  OAI211_X1 U20868 ( .C1(n17637), .C2(n17636), .A(n17635), .B(n17996), .ZN(
        n17638) );
  AOI221_X1 U20869 ( .B1(n17640), .B2(n17639), .C1(n17652), .C2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A(n17638), .ZN(n17641) );
  OAI21_X1 U20870 ( .B1(n17773), .B2(n17998), .A(n17641), .ZN(P3_U2810) );
  AOI21_X1 U20871 ( .B1(n17665), .B2(n17663), .A(n17642), .ZN(n17643) );
  XOR2_X1 U20872 ( .A(n17643), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Z(
        n18004) );
  AOI21_X1 U20873 ( .B1(n17846), .B2(n17645), .A(n17844), .ZN(n17677) );
  OAI21_X1 U20874 ( .B1(n17644), .B2(n17895), .A(n17677), .ZN(n17659) );
  AOI22_X1 U20875 ( .A1(n18218), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17659), .ZN(n17649) );
  NOR2_X1 U20876 ( .A1(n17646), .A2(n17645), .ZN(n17661) );
  OAI211_X1 U20877 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17661), .B(n17647), .ZN(n17648) );
  OAI211_X1 U20878 ( .C1(n17728), .C2(n17650), .A(n17649), .B(n17648), .ZN(
        n17651) );
  AOI221_X1 U20879 ( .B1(n17653), .B2(n17999), .C1(n17652), .C2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n17651), .ZN(n17654) );
  OAI21_X1 U20880 ( .B1(n18004), .B2(n17773), .A(n17654), .ZN(P3_U2811) );
  INV_X1 U20881 ( .A(n17746), .ZN(n17786) );
  NAND2_X1 U20882 ( .A1(n17656), .A2(n17655), .ZN(n18018) );
  OAI22_X1 U20883 ( .A1(n18201), .A2(n18795), .B1(n17728), .B2(n17657), .ZN(
        n17658) );
  AOI221_X1 U20884 ( .B1(n17661), .B2(n17660), .C1(n17659), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17658), .ZN(n17667) );
  OAI21_X1 U20885 ( .B1(n17662), .B2(n17693), .A(n17692), .ZN(n17674) );
  AOI21_X1 U20886 ( .B1(n17798), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17663), .ZN(n17664) );
  XOR2_X1 U20887 ( .A(n17665), .B(n17664), .Z(n18014) );
  AOI22_X1 U20888 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17674), .B1(
        n17799), .B2(n18014), .ZN(n17666) );
  OAI211_X1 U20889 ( .C1(n17786), .C2(n18018), .A(n17667), .B(n17666), .ZN(
        P3_U2812) );
  AOI21_X1 U20890 ( .B1(n18616), .B2(n17668), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17678) );
  INV_X1 U20891 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18793) );
  OAI22_X1 U20892 ( .A1(n18201), .A2(n18793), .B1(n17669), .B2(n17891), .ZN(
        n17670) );
  INV_X1 U20893 ( .A(n17670), .ZN(n17676) );
  AOI21_X1 U20894 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17672), .A(
        n17671), .ZN(n18019) );
  NAND2_X1 U20895 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18020), .ZN(
        n18026) );
  OAI22_X1 U20896 ( .A1(n18019), .A2(n17773), .B1(n17693), .B2(n18026), .ZN(
        n17673) );
  AOI21_X1 U20897 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17674), .A(
        n17673), .ZN(n17675) );
  OAI211_X1 U20898 ( .C1(n17678), .C2(n17677), .A(n17676), .B(n17675), .ZN(
        P3_U2813) );
  AOI22_X1 U20899 ( .A1(n17774), .A2(n10173), .B1(n17680), .B2(n17760), .ZN(
        n17681) );
  XOR2_X1 U20900 ( .A(n18034), .B(n17681), .Z(n18031) );
  AOI21_X1 U20901 ( .B1(n17846), .B2(n17682), .A(n17844), .ZN(n17708) );
  OAI21_X1 U20902 ( .B1(n17683), .B2(n17895), .A(n17708), .ZN(n17696) );
  AOI22_X1 U20903 ( .A1(n18218), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17696), .ZN(n17688) );
  NAND2_X1 U20904 ( .A1(n17724), .A2(n17684), .ZN(n17738) );
  NOR2_X1 U20905 ( .A1(n17685), .A2(n17738), .ZN(n17698) );
  OAI211_X1 U20906 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17698), .B(n17686), .ZN(n17687) );
  OAI211_X1 U20907 ( .C1(n17728), .C2(n17689), .A(n17688), .B(n17687), .ZN(
        n17690) );
  AOI21_X1 U20908 ( .B1(n17799), .B2(n18031), .A(n17690), .ZN(n17691) );
  OAI221_X1 U20909 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17693), 
        .C1(n18034), .C2(n17692), .A(n17691), .ZN(P3_U2814) );
  AND2_X1 U20910 ( .A1(n17706), .A2(n18050), .ZN(n18042) );
  NAND2_X1 U20911 ( .A1(n17745), .A2(n17963), .ZN(n17705) );
  INV_X1 U20912 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17697) );
  NAND2_X1 U20913 ( .A1(n18218), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18048) );
  OAI21_X1 U20914 ( .B1(n17728), .B2(n17694), .A(n18048), .ZN(n17695) );
  AOI221_X1 U20915 ( .B1(n17698), .B2(n17697), .C1(n17696), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17695), .ZN(n17704) );
  NAND3_X1 U20916 ( .A1(n18074), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        n17774), .ZN(n17719) );
  NOR2_X1 U20917 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17699), .ZN(
        n17775) );
  NAND2_X1 U20918 ( .A1(n17766), .A2(n17775), .ZN(n17747) );
  OR3_X1 U20919 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n17747), .ZN(n17715) );
  INV_X1 U20920 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18092) );
  NOR2_X1 U20921 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18092), .ZN(
        n18072) );
  AOI221_X1 U20922 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17719), 
        .C1(n17714), .C2(n17715), .A(n18072), .ZN(n17700) );
  XOR2_X1 U20923 ( .A(n17700), .B(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .Z(
        n18046) );
  NOR2_X1 U20924 ( .A1(n17964), .A2(n17899), .ZN(n17702) );
  NOR3_X1 U20925 ( .A1(n17744), .A2(n17714), .A3(n18058), .ZN(n17712) );
  NOR2_X1 U20926 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17712), .ZN(
        n18044) );
  INV_X1 U20927 ( .A(n18044), .ZN(n17701) );
  AOI22_X1 U20928 ( .A1(n17799), .A2(n18046), .B1(n17702), .B2(n17701), .ZN(
        n17703) );
  OAI211_X1 U20929 ( .C1(n18042), .C2(n17705), .A(n17704), .B(n17703), .ZN(
        P3_U2815) );
  OAI21_X1 U20930 ( .B1(n17707), .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n17706), .ZN(n18069) );
  NAND2_X1 U20931 ( .A1(n18616), .A2(n17724), .ZN(n17752) );
  AOI221_X1 U20932 ( .B1(n17725), .B2(n17709), .C1(n17752), .C2(n17709), .A(
        n17708), .ZN(n17710) );
  NOR2_X1 U20933 ( .A1(n18201), .A2(n18788), .ZN(n18064) );
  AOI211_X1 U20934 ( .C1(n17711), .C2(n17855), .A(n17710), .B(n18064), .ZN(
        n17718) );
  INV_X1 U20935 ( .A(n18058), .ZN(n18060) );
  NAND2_X1 U20936 ( .A1(n18060), .A2(n18094), .ZN(n17713) );
  AOI21_X1 U20937 ( .B1(n17714), .B2(n17713), .A(n17712), .ZN(n18066) );
  AOI21_X1 U20938 ( .B1(n17715), .B2(n17719), .A(n18072), .ZN(n17716) );
  XOR2_X1 U20939 ( .A(n17716), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(
        n18065) );
  AOI22_X1 U20940 ( .A1(n17800), .A2(n18066), .B1(n17799), .B2(n18065), .ZN(
        n17717) );
  OAI211_X1 U20941 ( .C1(n17803), .C2(n18069), .A(n17718), .B(n17717), .ZN(
        P3_U2816) );
  INV_X1 U20942 ( .A(n17774), .ZN(n17759) );
  INV_X1 U20943 ( .A(n18074), .ZN(n18070) );
  OAI22_X1 U20944 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17747), .B1(
        n17759), .B2(n18070), .ZN(n17733) );
  NAND2_X1 U20945 ( .A1(n18092), .A2(n17733), .ZN(n17732) );
  OAI21_X1 U20946 ( .B1(n17747), .B2(n17732), .A(n17719), .ZN(n17720) );
  XNOR2_X1 U20947 ( .A(n17720), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18084) );
  INV_X1 U20948 ( .A(n17846), .ZN(n17789) );
  AOI21_X1 U20949 ( .B1(n17722), .B2(n17721), .A(n17844), .ZN(n17723) );
  OAI21_X1 U20950 ( .B1(n17724), .B2(n17789), .A(n17723), .ZN(n17736) );
  NOR2_X1 U20951 ( .A1(n18201), .A2(n18785), .ZN(n18071) );
  OAI21_X1 U20952 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17725), .ZN(n17726) );
  OAI22_X1 U20953 ( .A1(n17728), .A2(n17727), .B1(n17738), .B2(n17726), .ZN(
        n17729) );
  AOI211_X1 U20954 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17736), .A(
        n18071), .B(n17729), .ZN(n17731) );
  NOR2_X1 U20955 ( .A1(n18099), .A2(n18055), .ZN(n18077) );
  NOR2_X1 U20956 ( .A1(n17744), .A2(n18055), .ZN(n18075) );
  OAI22_X1 U20957 ( .A1(n18077), .A2(n17803), .B1(n18075), .B2(n17899), .ZN(
        n17740) );
  NOR2_X1 U20958 ( .A1(n17786), .A2(n18070), .ZN(n17741) );
  AOI22_X1 U20959 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17740), .B1(
        n18072), .B2(n17741), .ZN(n17730) );
  OAI211_X1 U20960 ( .C1(n18084), .C2(n17773), .A(n17731), .B(n17730), .ZN(
        P3_U2817) );
  OAI21_X1 U20961 ( .B1(n17733), .B2(n18092), .A(n17732), .ZN(n18089) );
  INV_X1 U20962 ( .A(n18089), .ZN(n17743) );
  AOI22_X1 U20963 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17736), .B1(
        n17735), .B2(n17734), .ZN(n17737) );
  NAND2_X1 U20964 ( .A1(n18218), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18090) );
  OAI211_X1 U20965 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n17738), .A(
        n17737), .B(n18090), .ZN(n17739) );
  AOI221_X1 U20966 ( .B1(n17741), .B2(n18092), .C1(n17740), .C2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17739), .ZN(n17742) );
  OAI21_X1 U20967 ( .B1(n17743), .B2(n17773), .A(n17742), .ZN(P3_U2818) );
  AOI22_X1 U20968 ( .A1(n17745), .A2(n18099), .B1(n17800), .B2(n17744), .ZN(
        n17785) );
  NAND2_X1 U20969 ( .A1(n18103), .A2(n17746), .ZN(n17765) );
  OAI21_X1 U20970 ( .B1(n17759), .B2(n18103), .A(n17747), .ZN(n17748) );
  XNOR2_X1 U20971 ( .A(n17758), .B(n17748), .ZN(n18093) );
  INV_X1 U20972 ( .A(n18103), .ZN(n17749) );
  NAND2_X1 U20973 ( .A1(n17749), .A2(n17758), .ZN(n18110) );
  NAND4_X1 U20974 ( .A1(n18616), .A2(n17788), .A3(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17779) );
  NOR2_X1 U20975 ( .A1(n17778), .A2(n17779), .ZN(n17777) );
  NAND2_X1 U20976 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17777), .ZN(
        n17767) );
  OAI21_X1 U20977 ( .B1(n17889), .B2(n17750), .A(n17767), .ZN(n17751) );
  AOI22_X1 U20978 ( .A1(n17753), .A2(n17855), .B1(n17752), .B2(n17751), .ZN(
        n17755) );
  NAND2_X1 U20979 ( .A1(n18218), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n17754) );
  OAI211_X1 U20980 ( .C1(n17786), .C2(n18110), .A(n17755), .B(n17754), .ZN(
        n17756) );
  AOI21_X1 U20981 ( .B1(n17799), .B2(n18093), .A(n17756), .ZN(n17757) );
  OAI221_X1 U20982 ( .B1(n17758), .B2(n17785), .C1(n17758), .C2(n17765), .A(
        n17757), .ZN(P3_U2819) );
  OAI221_X1 U20983 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n17759), 
        .C1(n17764), .C2(n17774), .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17762) );
  NAND4_X1 U20984 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n9921), .A3(
        n17760), .A4(n18113), .ZN(n17761) );
  OAI211_X1 U20985 ( .C1(n17775), .C2(n17763), .A(n17762), .B(n17761), .ZN(
        n18118) );
  OAI22_X1 U20986 ( .A1(n17766), .A2(n17765), .B1(n17785), .B2(n17764), .ZN(
        n17771) );
  INV_X1 U20987 ( .A(n17889), .ZN(n17825) );
  OAI211_X1 U20988 ( .C1(n17777), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n17825), .B(n17767), .ZN(n17768) );
  NAND2_X1 U20989 ( .A1(n18218), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n18116) );
  OAI211_X1 U20990 ( .C1(n17891), .C2(n17769), .A(n17768), .B(n18116), .ZN(
        n17770) );
  NOR2_X1 U20991 ( .A1(n17771), .A2(n17770), .ZN(n17772) );
  OAI21_X1 U20992 ( .B1(n18118), .B2(n17773), .A(n17772), .ZN(P3_U2820) );
  NOR2_X1 U20993 ( .A1(n17775), .A2(n17774), .ZN(n17776) );
  XOR2_X1 U20994 ( .A(n17776), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n18125) );
  INV_X1 U20995 ( .A(n18125), .ZN(n17783) );
  AOI211_X1 U20996 ( .C1(n17779), .C2(n17778), .A(n17889), .B(n17777), .ZN(
        n17782) );
  NAND2_X1 U20997 ( .A1(n18218), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n18122) );
  OAI21_X1 U20998 ( .B1(n17891), .B2(n17780), .A(n18122), .ZN(n17781) );
  AOI211_X1 U20999 ( .C1(n17799), .C2(n17783), .A(n17782), .B(n17781), .ZN(
        n17784) );
  OAI221_X1 U21000 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17786), .C1(
        n18113), .C2(n17785), .A(n17784), .ZN(P3_U2821) );
  AOI221_X1 U21001 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C1(n17787), .C2(n17790), .A(n18575), .ZN(n17794) );
  OAI21_X1 U21002 ( .B1(n17789), .B2(n17788), .A(n17894), .ZN(n17808) );
  INV_X1 U21003 ( .A(n17808), .ZN(n17791) );
  OAI22_X1 U21004 ( .A1(n17891), .A2(n17792), .B1(n17791), .B2(n17790), .ZN(
        n17793) );
  AOI211_X1 U21005 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n18218), .A(n17794), .B(
        n17793), .ZN(n17802) );
  AOI21_X1 U21006 ( .B1(n17796), .B2(n18135), .A(n17795), .ZN(n18139) );
  AOI21_X1 U21007 ( .B1(n17798), .B2(n18143), .A(n17797), .ZN(n18137) );
  AOI22_X1 U21008 ( .A1(n17800), .A2(n18139), .B1(n17799), .B2(n18137), .ZN(
        n17801) );
  OAI211_X1 U21009 ( .C1(n17803), .C2(n18143), .A(n17802), .B(n17801), .ZN(
        P3_U2822) );
  OAI21_X1 U21010 ( .B1(n17806), .B2(n17805), .A(n17804), .ZN(n17807) );
  XOR2_X1 U21011 ( .A(n17807), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18152) );
  NOR2_X1 U21012 ( .A1(n18575), .A2(n10134), .ZN(n17809) );
  NOR2_X1 U21013 ( .A1(n18201), .A2(n18773), .ZN(n18148) );
  AOI221_X1 U21014 ( .B1(n17809), .B2(n10129), .C1(n17808), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18148), .ZN(n17814) );
  AOI21_X1 U21015 ( .B1(n18146), .B2(n17811), .A(n17810), .ZN(n18149) );
  AOI22_X1 U21016 ( .A1(n9816), .A2(n18149), .B1(n17812), .B2(n17855), .ZN(
        n17813) );
  OAI211_X1 U21017 ( .C1(n17899), .C2(n18152), .A(n17814), .B(n17813), .ZN(
        P3_U2823) );
  AOI22_X1 U21018 ( .A1(n17816), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n18157), .B2(n17815), .ZN(n17821) );
  AOI22_X1 U21019 ( .A1(n17819), .A2(n17832), .B1(n17818), .B2(n17817), .ZN(
        n17820) );
  XNOR2_X1 U21020 ( .A(n17821), .B(n17820), .ZN(n18154) );
  NOR2_X1 U21021 ( .A1(n18575), .A2(n17826), .ZN(n17822) );
  AOI22_X1 U21022 ( .A1(n18218), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n17822), 
        .B2(n17827), .ZN(n17831) );
  AOI21_X1 U21023 ( .B1(n9943), .B2(n17824), .A(n17823), .ZN(n18156) );
  OAI21_X1 U21024 ( .B1(n17826), .B2(n18575), .A(n17825), .ZN(n17839) );
  OAI22_X1 U21025 ( .A1(n17891), .A2(n17828), .B1(n17827), .B2(n17839), .ZN(
        n17829) );
  AOI21_X1 U21026 ( .B1(n9816), .B2(n18156), .A(n17829), .ZN(n17830) );
  OAI211_X1 U21027 ( .C1(n18154), .C2(n17899), .A(n17831), .B(n17830), .ZN(
        P3_U2824) );
  OAI21_X1 U21028 ( .B1(n17834), .B2(n17833), .A(n17832), .ZN(n18168) );
  AOI21_X1 U21029 ( .B1(n17837), .B2(n17836), .A(n17835), .ZN(n18165) );
  AOI21_X1 U21030 ( .B1(n17838), .B2(n17894), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17840) );
  OAI22_X1 U21031 ( .A1(n17891), .A2(n17841), .B1(n17840), .B2(n17839), .ZN(
        n17842) );
  AOI21_X1 U21032 ( .B1(n9816), .B2(n18165), .A(n17842), .ZN(n17843) );
  NAND2_X1 U21033 ( .A1(n18218), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18166) );
  OAI211_X1 U21034 ( .C1(n17899), .C2(n18168), .A(n17843), .B(n18166), .ZN(
        P3_U2825) );
  AOI21_X1 U21035 ( .B1(n17846), .B2(n17845), .A(n17844), .ZN(n17867) );
  OAI21_X1 U21036 ( .B1(n17849), .B2(n17848), .A(n17847), .ZN(n18178) );
  OAI22_X1 U21037 ( .A1(n17899), .A2(n18178), .B1(n18201), .B2(n18767), .ZN(
        n17850) );
  AOI21_X1 U21038 ( .B1(n18616), .B2(n17851), .A(n17850), .ZN(n17858) );
  AOI21_X1 U21039 ( .B1(n17854), .B2(n17853), .A(n17852), .ZN(n18176) );
  AOI22_X1 U21040 ( .A1(n9816), .A2(n18176), .B1(n17856), .B2(n17855), .ZN(
        n17857) );
  OAI211_X1 U21041 ( .C1(n17859), .C2(n17867), .A(n17858), .B(n17857), .ZN(
        P3_U2826) );
  OAI21_X1 U21042 ( .B1(n17862), .B2(n17861), .A(n17860), .ZN(n18186) );
  OAI21_X1 U21043 ( .B1(n17865), .B2(n17864), .A(n17863), .ZN(n17866) );
  XOR2_X1 U21044 ( .A(n17866), .B(n10170), .Z(n18184) );
  AOI21_X1 U21045 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17894), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17868) );
  OAI22_X1 U21046 ( .A1(n17891), .A2(n17869), .B1(n17868), .B2(n17867), .ZN(
        n17870) );
  AOI21_X1 U21047 ( .B1(n9816), .B2(n18184), .A(n17870), .ZN(n17871) );
  NAND2_X1 U21048 ( .A1(n18218), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18182) );
  OAI211_X1 U21049 ( .C1(n17899), .C2(n18186), .A(n17871), .B(n18182), .ZN(
        P3_U2827) );
  AOI21_X1 U21050 ( .B1(n17874), .B2(n17873), .A(n17872), .ZN(n18198) );
  NOR2_X1 U21051 ( .A1(n18201), .A2(n18763), .ZN(n18197) );
  OAI21_X1 U21052 ( .B1(n17877), .B2(n17876), .A(n17875), .ZN(n18200) );
  OAI22_X1 U21053 ( .A1(n17891), .A2(n17878), .B1(n17899), .B2(n18200), .ZN(
        n17879) );
  AOI211_X1 U21054 ( .C1(n9816), .C2(n18198), .A(n18197), .B(n17879), .ZN(
        n17880) );
  OAI221_X1 U21055 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18575), .C1(
        n17881), .C2(n17894), .A(n17880), .ZN(P3_U2828) );
  AOI21_X1 U21056 ( .B1(n17883), .B2(n17893), .A(n17882), .ZN(n18206) );
  AOI21_X1 U21057 ( .B1(n17885), .B2(n17892), .A(n17884), .ZN(n18213) );
  OAI22_X1 U21058 ( .A1(n18213), .A2(n17899), .B1(n18201), .B2(n18870), .ZN(
        n17886) );
  AOI21_X1 U21059 ( .B1(n9816), .B2(n18206), .A(n17886), .ZN(n17888) );
  OAI221_X1 U21060 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17891), .C1(
        n17890), .C2(n17889), .A(n17888), .ZN(P3_U2829) );
  NAND2_X1 U21061 ( .A1(n17893), .A2(n17892), .ZN(n18221) );
  INV_X1 U21062 ( .A(n18221), .ZN(n17900) );
  NAND3_X1 U21063 ( .A1(n18847), .A2(n17895), .A3(n17894), .ZN(n17896) );
  AOI22_X1 U21064 ( .A1(n18218), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17896), .ZN(n17897) );
  OAI221_X1 U21065 ( .B1(n17900), .B2(n17899), .C1(n18221), .C2(n17898), .A(
        n17897), .ZN(P3_U2830) );
  OR2_X1 U21066 ( .A1(n17902), .A2(n17901), .ZN(n17954) );
  NOR2_X1 U21067 ( .A1(n17903), .A2(n17954), .ZN(n17912) );
  NOR2_X1 U21068 ( .A1(n18683), .A2(n18694), .ZN(n18187) );
  INV_X1 U21069 ( .A(n18187), .ZN(n18130) );
  NAND2_X1 U21070 ( .A1(n18694), .A2(n18846), .ZN(n18188) );
  INV_X1 U21071 ( .A(n18188), .ZN(n18128) );
  AOI21_X1 U21072 ( .B1(n17904), .B2(n18130), .A(n18128), .ZN(n17946) );
  OAI21_X1 U21073 ( .B1(n17928), .B2(n18187), .A(n17946), .ZN(n17924) );
  AOI211_X1 U21074 ( .C1(n17906), .C2(n18130), .A(n17905), .B(n17924), .ZN(
        n17907) );
  OAI21_X1 U21075 ( .B1(n17908), .B2(n18677), .A(n17907), .ZN(n17909) );
  AOI21_X1 U21076 ( .B1(n18100), .B2(n17910), .A(n17909), .ZN(n17919) );
  INV_X1 U21077 ( .A(n17919), .ZN(n17911) );
  MUX2_X1 U21078 ( .A(n17912), .B(n17911), .S(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(n17913) );
  AOI22_X1 U21079 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18209), .B1(
        n18214), .B2(n17913), .ZN(n17915) );
  NAND2_X1 U21080 ( .A1(n18218), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17914) );
  OAI211_X1 U21081 ( .C1(n17916), .C2(n18124), .A(n17915), .B(n17914), .ZN(
        P3_U2835) );
  OAI222_X1 U21082 ( .A1(n17920), .A2(n17954), .B1(n17923), .B2(n17919), .C1(
        n17918), .C2(n17917), .ZN(n17921) );
  AOI22_X1 U21083 ( .A1(n18218), .A2(P3_REIP_REG_26__SCAN_IN), .B1(n18214), 
        .B2(n17921), .ZN(n17922) );
  OAI21_X1 U21084 ( .B1(n17923), .B2(n18194), .A(n17922), .ZN(P3_U2836) );
  AOI221_X1 U21085 ( .B1(n17947), .B2(n18684), .C1(n17925), .C2(n18684), .A(
        n17924), .ZN(n17931) );
  NAND3_X1 U21086 ( .A1(n17928), .A2(n17927), .A3(n17926), .ZN(n17930) );
  AOI221_X1 U21087 ( .B1(n17931), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), 
        .C1(n17930), .C2(n17929), .A(n18207), .ZN(n17932) );
  AOI211_X1 U21088 ( .C1(n18209), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17933), .B(n17932), .ZN(n17939) );
  INV_X1 U21089 ( .A(n17934), .ZN(n17936) );
  AOI22_X1 U21090 ( .A1(n17937), .A2(n17936), .B1(n18217), .B2(n17935), .ZN(
        n17938) );
  OAI211_X1 U21091 ( .C1(n18124), .C2(n17940), .A(n17939), .B(n17938), .ZN(
        P3_U2837) );
  AOI21_X1 U21092 ( .B1(n17942), .B2(n17981), .A(n17941), .ZN(n17951) );
  AOI22_X1 U21093 ( .A1(n18037), .A2(n17944), .B1(n18100), .B2(n17943), .ZN(
        n17945) );
  NAND3_X1 U21094 ( .A1(n17946), .A2(n17945), .A3(n18194), .ZN(n17949) );
  AOI211_X1 U21095 ( .C1(n18684), .C2(n17947), .A(n17953), .B(n17949), .ZN(
        n17948) );
  NOR2_X1 U21096 ( .A1(n17990), .A2(n17948), .ZN(n17956) );
  OAI211_X1 U21097 ( .C1(n18132), .C2(n17949), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17956), .ZN(n17950) );
  OAI211_X1 U21098 ( .C1(n17952), .C2(n18124), .A(n17951), .B(n17950), .ZN(
        P3_U2838) );
  OAI21_X1 U21099 ( .B1(n18209), .B2(n17954), .A(n17953), .ZN(n17955) );
  AOI22_X1 U21100 ( .A1(n18138), .A2(n17957), .B1(n17956), .B2(n17955), .ZN(
        n17959) );
  NAND2_X1 U21101 ( .A1(n17959), .A2(n17958), .ZN(P3_U2839) );
  INV_X1 U21102 ( .A(n17960), .ZN(n17962) );
  AOI22_X1 U21103 ( .A1(n18138), .A2(n17962), .B1(n17981), .B2(n17961), .ZN(
        n17976) );
  NAND2_X1 U21104 ( .A1(n18100), .A2(n17963), .ZN(n18043) );
  OAI211_X1 U21105 ( .C1(n17964), .C2(n18677), .A(n18214), .B(n18043), .ZN(
        n18030) );
  NAND2_X1 U21106 ( .A1(n18677), .A2(n18076), .ZN(n18102) );
  AOI21_X1 U21107 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n18011), .A(
        n18709), .ZN(n17965) );
  AOI221_X1 U21108 ( .B1(n18009), .B2(n18683), .C1(n17989), .C2(n18683), .A(
        n17965), .ZN(n17987) );
  OAI21_X1 U21109 ( .B1(n18696), .B2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n17987), .ZN(n17966) );
  AOI21_X1 U21110 ( .B1(n17967), .B2(n18102), .A(n17966), .ZN(n17978) );
  AOI22_X1 U21111 ( .A1(n18684), .A2(n17970), .B1(n17969), .B2(n17968), .ZN(
        n17971) );
  OAI211_X1 U21112 ( .C1(n18104), .C2(n17972), .A(n17978), .B(n17971), .ZN(
        n17973) );
  OAI211_X1 U21113 ( .C1(n18030), .C2(n17973), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n18201), .ZN(n17974) );
  NAND3_X1 U21114 ( .A1(n17976), .A2(n17975), .A3(n17974), .ZN(P3_U2840) );
  NOR2_X1 U21115 ( .A1(n18684), .A2(n18694), .ZN(n18208) );
  AOI221_X1 U21116 ( .B1(n18028), .B2(n18694), .C1(n17977), .C2(n18694), .A(
        n18030), .ZN(n17992) );
  OAI211_X1 U21117 ( .C1(n17979), .C2(n18208), .A(n17992), .B(n17978), .ZN(
        n17980) );
  NAND2_X1 U21118 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17980), .ZN(
        n17985) );
  NAND2_X1 U21119 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17981), .ZN(
        n17986) );
  INV_X1 U21120 ( .A(n17986), .ZN(n18000) );
  AOI22_X1 U21121 ( .A1(n18138), .A2(n17983), .B1(n17982), .B2(n18000), .ZN(
        n17984) );
  OAI221_X1 U21122 ( .B1(n18218), .B2(n17985), .C1(n18201), .C2(n18801), .A(
        n17984), .ZN(P3_U2841) );
  OR2_X1 U21123 ( .A1(n17999), .A2(n17986), .ZN(n17995) );
  INV_X1 U21124 ( .A(n17987), .ZN(n17988) );
  AOI21_X1 U21125 ( .B1(n17989), .B2(n18102), .A(n17988), .ZN(n17991) );
  AOI21_X1 U21126 ( .B1(n17992), .B2(n17991), .A(n17990), .ZN(n18001) );
  NOR3_X1 U21127 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18208), .A3(
        n18726), .ZN(n17993) );
  NOR2_X1 U21128 ( .A1(n18001), .A2(n17993), .ZN(n17994) );
  MUX2_X1 U21129 ( .A(n17995), .B(n17994), .S(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .Z(n17997) );
  OAI211_X1 U21130 ( .C1(n17998), .C2(n18124), .A(n17997), .B(n17996), .ZN(
        P3_U2842) );
  AOI22_X1 U21131 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18001), .B1(
        n18000), .B2(n17999), .ZN(n18003) );
  NAND2_X1 U21132 ( .A1(n18218), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18002) );
  OAI211_X1 U21133 ( .C1(n18004), .C2(n18124), .A(n18003), .B(n18002), .ZN(
        P3_U2843) );
  INV_X1 U21134 ( .A(n18005), .ZN(n18007) );
  INV_X1 U21135 ( .A(n18006), .ZN(n18189) );
  OAI22_X1 U21136 ( .A1(n18127), .A2(n18709), .B1(n18129), .B2(n18189), .ZN(
        n18180) );
  NAND2_X1 U21137 ( .A1(n18007), .A2(n18180), .ZN(n18145) );
  NOR3_X1 U21138 ( .A1(n18135), .A2(n18146), .A3(n18145), .ZN(n18059) );
  OAI21_X1 U21139 ( .B1(n18059), .B2(n18008), .A(n18214), .ZN(n18109) );
  OAI21_X1 U21140 ( .B1(n18009), .B2(n18034), .A(n18130), .ZN(n18010) );
  OAI211_X1 U21141 ( .C1(n18011), .C2(n18709), .A(n18188), .B(n18010), .ZN(
        n18012) );
  AOI211_X1 U21142 ( .C1(n18013), .C2(n18102), .A(n18030), .B(n18012), .ZN(
        n18021) );
  AOI221_X1 U21143 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18021), 
        .C1(n18187), .C2(n18021), .A(n18218), .ZN(n18015) );
  AOI22_X1 U21144 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18015), .B1(
        n18138), .B2(n18014), .ZN(n18017) );
  NAND2_X1 U21145 ( .A1(n18218), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18016) );
  OAI211_X1 U21146 ( .C1(n18018), .C2(n18109), .A(n18017), .B(n18016), .ZN(
        P3_U2844) );
  INV_X1 U21147 ( .A(n18109), .ZN(n18121) );
  NAND2_X1 U21148 ( .A1(n10173), .A2(n18121), .ZN(n18035) );
  INV_X1 U21149 ( .A(n18019), .ZN(n18023) );
  NOR3_X1 U21150 ( .A1(n18218), .A2(n18021), .A3(n18020), .ZN(n18022) );
  AOI21_X1 U21151 ( .B1(n18138), .B2(n18023), .A(n18022), .ZN(n18025) );
  NAND2_X1 U21152 ( .A1(n18218), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n18024) );
  OAI211_X1 U21153 ( .C1(n18026), .C2(n18035), .A(n18025), .B(n18024), .ZN(
        P3_U2845) );
  NOR2_X1 U21154 ( .A1(n18696), .A2(n18027), .ZN(n18051) );
  AOI21_X1 U21155 ( .B1(n18684), .B2(n18054), .A(n18051), .ZN(n18095) );
  OAI21_X1 U21156 ( .B1(n18050), .B2(n18694), .A(n18028), .ZN(n18029) );
  OAI211_X1 U21157 ( .C1(n18112), .C2(n18038), .A(n18095), .B(n18029), .ZN(
        n18039) );
  OAI221_X1 U21158 ( .B1(n18030), .B2(n18132), .C1(n18030), .C2(n18039), .A(
        n18201), .ZN(n18033) );
  AOI22_X1 U21159 ( .A1(n18218), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n18138), 
        .B2(n18031), .ZN(n18032) );
  OAI221_X1 U21160 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18035), 
        .C1(n18034), .C2(n18033), .A(n18032), .ZN(P3_U2846) );
  NAND2_X1 U21161 ( .A1(n18037), .A2(n18036), .ZN(n18045) );
  AOI21_X1 U21162 ( .B1(n18038), .B2(n18059), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18041) );
  INV_X1 U21163 ( .A(n18039), .ZN(n18040) );
  OAI222_X1 U21164 ( .A1(n18045), .A2(n18044), .B1(n18043), .B2(n18042), .C1(
        n18041), .C2(n18040), .ZN(n18047) );
  AOI22_X1 U21165 ( .A1(n18214), .A2(n18047), .B1(n18138), .B2(n18046), .ZN(
        n18049) );
  OAI211_X1 U21166 ( .C1(n18194), .C2(n18050), .A(n18049), .B(n18048), .ZN(
        P3_U2847) );
  INV_X1 U21167 ( .A(n18051), .ZN(n18052) );
  OAI221_X1 U21168 ( .B1(n18104), .B2(n18053), .C1(n18104), .C2(n18096), .A(
        n18052), .ZN(n18079) );
  OAI21_X1 U21169 ( .B1(n18055), .B2(n18054), .A(n18684), .ZN(n18056) );
  OAI211_X1 U21170 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n18208), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n18056), .ZN(n18057) );
  AOI211_X1 U21171 ( .C1(n18683), .C2(n18058), .A(n18079), .B(n18057), .ZN(
        n18062) );
  AOI21_X1 U21172 ( .B1(n18060), .B2(n18059), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18061) );
  NOR3_X1 U21173 ( .A1(n18062), .A2(n18061), .A3(n18207), .ZN(n18063) );
  AOI211_X1 U21174 ( .C1(n18209), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n18064), .B(n18063), .ZN(n18068) );
  AOI22_X1 U21175 ( .A1(n18217), .A2(n18066), .B1(n18138), .B2(n18065), .ZN(
        n18067) );
  OAI211_X1 U21176 ( .C1(n18142), .C2(n18069), .A(n18068), .B(n18067), .ZN(
        P3_U2848) );
  NOR2_X1 U21177 ( .A1(n18070), .A2(n18109), .ZN(n18085) );
  AOI21_X1 U21178 ( .B1(n18072), .B2(n18085), .A(n18071), .ZN(n18083) );
  NOR2_X1 U21179 ( .A1(n18073), .A2(n18709), .ZN(n18080) );
  NOR2_X1 U21180 ( .A1(n18112), .A2(n18074), .ZN(n18106) );
  OAI22_X1 U21181 ( .A1(n18077), .A2(n18076), .B1(n18075), .B2(n18677), .ZN(
        n18078) );
  NOR4_X1 U21182 ( .A1(n18080), .A2(n18106), .A3(n18079), .A4(n18078), .ZN(
        n18087) );
  OAI211_X1 U21183 ( .C1(n18112), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18214), .B(n18087), .ZN(n18081) );
  NAND3_X1 U21184 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18201), .A3(
        n18081), .ZN(n18082) );
  OAI211_X1 U21185 ( .C1(n18084), .C2(n18124), .A(n18083), .B(n18082), .ZN(
        P3_U2849) );
  AOI21_X1 U21186 ( .B1(n18214), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18085), .ZN(n18086) );
  AOI21_X1 U21187 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18087), .A(
        n18086), .ZN(n18088) );
  AOI21_X1 U21188 ( .B1(n18138), .B2(n18089), .A(n18088), .ZN(n18091) );
  OAI211_X1 U21189 ( .C1(n18194), .C2(n18092), .A(n18091), .B(n18090), .ZN(
        P3_U2850) );
  AOI22_X1 U21190 ( .A1(n18218), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18138), 
        .B2(n18093), .ZN(n18108) );
  NOR2_X1 U21191 ( .A1(n18677), .A2(n18094), .ZN(n18098) );
  OAI211_X1 U21192 ( .C1(n18104), .C2(n18096), .A(n18214), .B(n18095), .ZN(
        n18097) );
  AOI211_X1 U21193 ( .C1(n18100), .C2(n18099), .A(n18098), .B(n18097), .ZN(
        n18119) );
  OAI21_X1 U21194 ( .B1(n18104), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n18119), .ZN(n18101) );
  AOI21_X1 U21195 ( .B1(n18103), .B2(n18102), .A(n18101), .ZN(n18111) );
  OAI21_X1 U21196 ( .B1(n18104), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18111), .ZN(n18105) );
  OAI211_X1 U21197 ( .C1(n18106), .C2(n18105), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18201), .ZN(n18107) );
  OAI211_X1 U21198 ( .C1(n18110), .C2(n18109), .A(n18108), .B(n18107), .ZN(
        P3_U2851) );
  AOI221_X1 U21199 ( .B1(n18112), .B2(n18111), .C1(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18111), .A(n18218), .ZN(
        n18115) );
  NOR2_X1 U21200 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18113), .ZN(
        n18114) );
  AOI22_X1 U21201 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18115), .B1(
        n18121), .B2(n18114), .ZN(n18117) );
  OAI211_X1 U21202 ( .C1(n18124), .C2(n18118), .A(n18117), .B(n18116), .ZN(
        P3_U2852) );
  OAI21_X1 U21203 ( .B1(n18218), .B2(n18119), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18120) );
  OAI21_X1 U21204 ( .B1(n18121), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n18120), .ZN(n18123) );
  OAI211_X1 U21205 ( .C1(n18125), .C2(n18124), .A(n18123), .B(n18122), .ZN(
        P3_U2853) );
  AND3_X1 U21206 ( .A1(n18126), .A2(n18214), .A3(n18180), .ZN(n18136) );
  AND2_X1 U21207 ( .A1(n18684), .A2(n18127), .ZN(n18193) );
  AOI211_X1 U21208 ( .C1(n18130), .C2(n18129), .A(n18128), .B(n18193), .ZN(
        n18169) );
  OAI21_X1 U21209 ( .B1(n18131), .B2(n18158), .A(n18169), .ZN(n18153) );
  AOI211_X1 U21210 ( .C1(n18132), .C2(n18157), .A(n18146), .B(n18153), .ZN(
        n18144) );
  OAI21_X1 U21211 ( .B1(n18144), .B2(n18202), .A(n18194), .ZN(n18134) );
  NOR2_X1 U21212 ( .A1(n18201), .A2(n18776), .ZN(n18133) );
  AOI221_X1 U21213 ( .B1(n18136), .B2(n18135), .C1(n18134), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18133), .ZN(n18141) );
  AOI22_X1 U21214 ( .A1(n18217), .A2(n18139), .B1(n18138), .B2(n18137), .ZN(
        n18140) );
  OAI211_X1 U21215 ( .C1(n18143), .C2(n18142), .A(n18141), .B(n18140), .ZN(
        P3_U2854) );
  AOI211_X1 U21216 ( .C1(n18146), .C2(n18145), .A(n18144), .B(n18207), .ZN(
        n18147) );
  AOI211_X1 U21217 ( .C1(n18209), .C2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18148), .B(n18147), .ZN(n18151) );
  NAND2_X1 U21218 ( .A1(n18205), .A2(n18149), .ZN(n18150) );
  OAI211_X1 U21219 ( .C1(n18152), .C2(n18212), .A(n18151), .B(n18150), .ZN(
        P3_U2855) );
  AOI21_X1 U21220 ( .B1(n18214), .B2(n18153), .A(n18209), .ZN(n18161) );
  OAI22_X1 U21221 ( .A1(n18154), .A2(n18212), .B1(n18161), .B2(n18157), .ZN(
        n18155) );
  AOI21_X1 U21222 ( .B1(n18205), .B2(n18156), .A(n18155), .ZN(n18160) );
  NAND4_X1 U21223 ( .A1(n18214), .A2(n18158), .A3(n18157), .A4(n18180), .ZN(
        n18159) );
  OAI211_X1 U21224 ( .C1(n18771), .C2(n18201), .A(n18160), .B(n18159), .ZN(
        P3_U2856) );
  NAND3_X1 U21225 ( .A1(n18214), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18180), .ZN(n18172) );
  NOR2_X1 U21226 ( .A1(n18171), .A2(n18172), .ZN(n18163) );
  INV_X1 U21227 ( .A(n18161), .ZN(n18162) );
  MUX2_X1 U21228 ( .A(n18163), .B(n18162), .S(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(n18164) );
  AOI21_X1 U21229 ( .B1(n18205), .B2(n18165), .A(n18164), .ZN(n18167) );
  OAI211_X1 U21230 ( .C1(n18212), .C2(n18168), .A(n18167), .B(n18166), .ZN(
        P3_U2857) );
  NOR2_X1 U21231 ( .A1(n18201), .A2(n18767), .ZN(n18175) );
  NAND2_X1 U21232 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18169), .ZN(
        n18179) );
  AOI21_X1 U21233 ( .B1(n18170), .B2(n18179), .A(n18209), .ZN(n18173) );
  AOI22_X1 U21234 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18173), .B1(
        n18172), .B2(n18171), .ZN(n18174) );
  AOI211_X1 U21235 ( .C1(n18176), .C2(n18205), .A(n18175), .B(n18174), .ZN(
        n18177) );
  OAI21_X1 U21236 ( .B1(n18212), .B2(n18178), .A(n18177), .ZN(P3_U2858) );
  OAI211_X1 U21237 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n18180), .A(
        n18214), .B(n18179), .ZN(n18181) );
  OAI211_X1 U21238 ( .C1(n18194), .C2(n10170), .A(n18182), .B(n18181), .ZN(
        n18183) );
  AOI21_X1 U21239 ( .B1(n18205), .B2(n18184), .A(n18183), .ZN(n18185) );
  OAI21_X1 U21240 ( .B1(n18212), .B2(n18186), .A(n18185), .ZN(P3_U2859) );
  AOI211_X1 U21241 ( .C1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n18188), .A(
        n18187), .B(n15756), .ZN(n18192) );
  NAND2_X1 U21242 ( .A1(n18684), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18190) );
  AOI221_X1 U21243 ( .B1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n18190), .C1(
        n15756), .C2(n18189), .A(n18845), .ZN(n18191) );
  NOR3_X1 U21244 ( .A1(n18193), .A2(n18192), .A3(n18191), .ZN(n18195) );
  OAI22_X1 U21245 ( .A1(n18195), .A2(n18207), .B1(n15756), .B2(n18194), .ZN(
        n18196) );
  AOI211_X1 U21246 ( .C1(n18205), .C2(n18198), .A(n18197), .B(n18196), .ZN(
        n18199) );
  OAI21_X1 U21247 ( .B1(n18212), .B2(n18200), .A(n18199), .ZN(P3_U2860) );
  NOR2_X1 U21248 ( .A1(n18201), .A2(n18870), .ZN(n18204) );
  AOI211_X1 U21249 ( .C1(n18696), .C2(n18846), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18202), .ZN(n18203) );
  AOI211_X1 U21250 ( .C1(n18206), .C2(n18205), .A(n18204), .B(n18203), .ZN(
        n18211) );
  NOR3_X1 U21251 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18208), .A3(
        n18207), .ZN(n18216) );
  OAI21_X1 U21252 ( .B1(n18209), .B2(n18216), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18210) );
  OAI211_X1 U21253 ( .C1(n18213), .C2(n18212), .A(n18211), .B(n18210), .ZN(
        P3_U2861) );
  AOI211_X1 U21254 ( .C1(n18696), .C2(n18214), .A(n18218), .B(n18846), .ZN(
        n18215) );
  AOI211_X1 U21255 ( .C1(n18217), .C2(n18221), .A(n18216), .B(n18215), .ZN(
        n18220) );
  NAND2_X1 U21256 ( .A1(n18218), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n18219) );
  OAI211_X1 U21257 ( .C1(n18222), .C2(n18221), .A(n18220), .B(n18219), .ZN(
        P3_U2862) );
  AOI211_X1 U21258 ( .C1(n18224), .C2(n18223), .A(n18726), .B(n18847), .ZN(
        n18727) );
  OAI21_X1 U21259 ( .B1(n18727), .B2(n18273), .A(n18229), .ZN(n18225) );
  OAI221_X1 U21260 ( .B1(n18518), .B2(n18881), .C1(n18518), .C2(n18229), .A(
        n18225), .ZN(P3_U2863) );
  INV_X1 U21261 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18715) );
  NOR2_X1 U21262 ( .A1(n18715), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18519) );
  NAND2_X1 U21263 ( .A1(n18715), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18356) );
  INV_X1 U21264 ( .A(n18356), .ZN(n18404) );
  NOR2_X1 U21265 ( .A1(n18519), .A2(n18404), .ZN(n18227) );
  OAI22_X1 U21266 ( .A1(n18228), .A2(n18715), .B1(n18227), .B2(n18226), .ZN(
        P3_U2866) );
  NOR2_X1 U21267 ( .A1(n18716), .A2(n18229), .ZN(P3_U2867) );
  NOR2_X1 U21268 ( .A1(n18712), .A2(n18715), .ZN(n18233) );
  NAND2_X1 U21269 ( .A1(n18699), .A2(n18233), .ZN(n18545) );
  NOR2_X2 U21270 ( .A1(n18518), .A2(n18545), .ZN(n18662) );
  INV_X1 U21271 ( .A(n18662), .ZN(n18646) );
  NOR2_X1 U21272 ( .A1(n18230), .A2(n18575), .ZN(n18612) );
  INV_X1 U21273 ( .A(n18612), .ZN(n18581) );
  NOR2_X2 U21274 ( .A1(n18426), .A2(n18231), .ZN(n18611) );
  NOR2_X1 U21275 ( .A1(n18715), .A2(n18401), .ZN(n18614) );
  NAND2_X1 U21276 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18614), .ZN(
        n18312) );
  INV_X1 U21277 ( .A(n18312), .ZN(n18664) );
  NOR2_X1 U21278 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18425) );
  NOR2_X1 U21279 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18313) );
  NAND2_X1 U21280 ( .A1(n18425), .A2(n18313), .ZN(n18333) );
  NOR2_X1 U21281 ( .A1(n18664), .A2(n18326), .ZN(n18292) );
  NOR2_X1 U21282 ( .A1(n9814), .A2(n18292), .ZN(n18266) );
  NAND2_X1 U21283 ( .A1(n18616), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18620) );
  INV_X1 U21284 ( .A(n18620), .ZN(n18574) );
  NOR2_X1 U21285 ( .A1(n18699), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18472) );
  NAND2_X1 U21286 ( .A1(n18233), .A2(n18472), .ZN(n18598) );
  INV_X1 U21287 ( .A(n18598), .ZN(n18605) );
  AOI22_X1 U21288 ( .A1(n18611), .A2(n18266), .B1(n18574), .B2(n18605), .ZN(
        n18239) );
  INV_X1 U21289 ( .A(n18426), .ZN(n18524) );
  AOI21_X1 U21290 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18292), .ZN(n18234) );
  NOR2_X1 U21291 ( .A1(n18518), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18452) );
  NOR2_X1 U21292 ( .A1(n18472), .A2(n18452), .ZN(n18522) );
  INV_X1 U21293 ( .A(n18522), .ZN(n18232) );
  NAND2_X1 U21294 ( .A1(n18233), .A2(n18232), .ZN(n18573) );
  NOR2_X1 U21295 ( .A1(n18426), .A2(n18573), .ZN(n18578) );
  AOI22_X1 U21296 ( .A1(n18524), .A2(n18234), .B1(n18520), .B2(n18578), .ZN(
        n18269) );
  NAND2_X1 U21297 ( .A1(n18236), .A2(n18235), .ZN(n18267) );
  NOR2_X2 U21298 ( .A1(n18237), .A2(n18267), .ZN(n18617) );
  AOI22_X1 U21299 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18269), .B1(
        n18326), .B2(n18617), .ZN(n18238) );
  OAI211_X1 U21300 ( .C1(n18646), .C2(n18581), .A(n18239), .B(n18238), .ZN(
        P3_U2868) );
  INV_X1 U21301 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n18240) );
  NOR2_X1 U21302 ( .A1(n18240), .A2(n18575), .ZN(n18582) );
  INV_X1 U21303 ( .A(n18582), .ZN(n18626) );
  AND2_X1 U21304 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18524), .ZN(n18621) );
  AND2_X1 U21305 ( .A1(BUF2_REG_17__SCAN_IN), .A2(n18616), .ZN(n18622) );
  AOI22_X1 U21306 ( .A1(n18266), .A2(n18621), .B1(n18605), .B2(n18622), .ZN(
        n18242) );
  NOR2_X1 U21307 ( .A1(n18889), .A2(n18267), .ZN(n18623) );
  AOI22_X1 U21308 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18269), .B1(
        n18326), .B2(n18623), .ZN(n18241) );
  OAI211_X1 U21309 ( .C1(n18646), .C2(n18626), .A(n18242), .B(n18241), .ZN(
        P3_U2869) );
  NAND2_X1 U21310 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n18616), .ZN(n18554) );
  NAND2_X1 U21311 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18616), .ZN(n18632) );
  INV_X1 U21312 ( .A(n18632), .ZN(n18551) );
  NOR2_X2 U21313 ( .A1(n18243), .A2(n18426), .ZN(n18627) );
  AOI22_X1 U21314 ( .A1(n18662), .A2(n18551), .B1(n18266), .B2(n18627), .ZN(
        n18246) );
  NOR2_X2 U21315 ( .A1(n18244), .A2(n18267), .ZN(n18629) );
  AOI22_X1 U21316 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18269), .B1(
        n18326), .B2(n18629), .ZN(n18245) );
  OAI211_X1 U21317 ( .C1(n18598), .C2(n18554), .A(n18246), .B(n18245), .ZN(
        P3_U2870) );
  NAND2_X1 U21318 ( .A1(BUF2_REG_19__SCAN_IN), .A2(n18616), .ZN(n18638) );
  NAND2_X1 U21319 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18616), .ZN(n18591) );
  INV_X1 U21320 ( .A(n18591), .ZN(n18634) );
  NOR2_X2 U21321 ( .A1(n18247), .A2(n18426), .ZN(n18633) );
  AOI22_X1 U21322 ( .A1(n18662), .A2(n18634), .B1(n18266), .B2(n18633), .ZN(
        n18250) );
  NOR2_X2 U21323 ( .A1(n18248), .A2(n18267), .ZN(n18635) );
  AOI22_X1 U21324 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18269), .B1(
        n18326), .B2(n18635), .ZN(n18249) );
  OAI211_X1 U21325 ( .C1(n18598), .C2(n18638), .A(n18250), .B(n18249), .ZN(
        P3_U2871) );
  NOR2_X1 U21326 ( .A1(n18251), .A2(n18575), .ZN(n18641) );
  INV_X1 U21327 ( .A(n18641), .ZN(n18561) );
  NOR2_X2 U21328 ( .A1(n18252), .A2(n18426), .ZN(n18639) );
  NAND2_X1 U21329 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n18616), .ZN(n18645) );
  INV_X1 U21330 ( .A(n18645), .ZN(n18557) );
  AOI22_X1 U21331 ( .A1(n18266), .A2(n18639), .B1(n18605), .B2(n18557), .ZN(
        n18255) );
  NOR2_X2 U21332 ( .A1(n18253), .A2(n18267), .ZN(n18642) );
  AOI22_X1 U21333 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18269), .B1(
        n18326), .B2(n18642), .ZN(n18254) );
  OAI211_X1 U21334 ( .C1(n18646), .C2(n18561), .A(n18255), .B(n18254), .ZN(
        P3_U2872) );
  INV_X1 U21335 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18256) );
  INV_X1 U21336 ( .A(n18594), .ZN(n18652) );
  NOR2_X2 U21337 ( .A1(n18257), .A2(n18426), .ZN(n18647) );
  NOR2_X2 U21338 ( .A1(n19264), .A2(n18575), .ZN(n18648) );
  AOI22_X1 U21339 ( .A1(n18266), .A2(n18647), .B1(n18605), .B2(n18648), .ZN(
        n18260) );
  NOR2_X1 U21340 ( .A1(n18258), .A2(n18267), .ZN(n18649) );
  AOI22_X1 U21341 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18269), .B1(
        n18326), .B2(n18649), .ZN(n18259) );
  OAI211_X1 U21342 ( .C1(n18646), .C2(n18652), .A(n18260), .B(n18259), .ZN(
        P3_U2873) );
  NOR2_X1 U21343 ( .A1(n18261), .A2(n18575), .ZN(n18564) );
  INV_X1 U21344 ( .A(n18564), .ZN(n18658) );
  NOR2_X2 U21345 ( .A1(n18262), .A2(n18426), .ZN(n18653) );
  NAND2_X1 U21346 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18616), .ZN(n18567) );
  INV_X1 U21347 ( .A(n18567), .ZN(n18654) );
  AOI22_X1 U21348 ( .A1(n18266), .A2(n18653), .B1(n18605), .B2(n18654), .ZN(
        n18265) );
  NOR2_X2 U21349 ( .A1(n18263), .A2(n18267), .ZN(n18655) );
  AOI22_X1 U21350 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18269), .B1(
        n18326), .B2(n18655), .ZN(n18264) );
  OAI211_X1 U21351 ( .C1(n18646), .C2(n18658), .A(n18265), .B(n18264), .ZN(
        P3_U2874) );
  NAND2_X1 U21352 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18616), .ZN(n18609) );
  NAND2_X1 U21353 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n18616), .ZN(n18669) );
  INV_X1 U21354 ( .A(n18669), .ZN(n18604) );
  AND2_X1 U21355 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18524), .ZN(n18660) );
  AOI22_X1 U21356 ( .A1(n18662), .A2(n18604), .B1(n18266), .B2(n18660), .ZN(
        n18271) );
  NOR2_X2 U21357 ( .A1(n18268), .A2(n18267), .ZN(n18663) );
  AOI22_X1 U21358 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18269), .B1(
        n18326), .B2(n18663), .ZN(n18270) );
  OAI211_X1 U21359 ( .C1(n18598), .C2(n18609), .A(n18271), .B(n18270), .ZN(
        P3_U2875) );
  INV_X1 U21360 ( .A(n18313), .ZN(n18272) );
  AOI22_X1 U21361 ( .A1(n18664), .A2(n18574), .B1(n18611), .B2(n18288), .ZN(
        n18275) );
  NOR2_X1 U21362 ( .A1(n18426), .A2(n18273), .ZN(n18613) );
  AND2_X1 U21363 ( .A1(n18699), .A2(n18613), .ZN(n18450) );
  AOI22_X1 U21364 ( .A1(n18616), .A2(n18614), .B1(n18313), .B2(n18450), .ZN(
        n18289) );
  NAND2_X1 U21365 ( .A1(n18452), .A2(n18313), .ZN(n18355) );
  AOI22_X1 U21366 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18289), .B1(
        n18617), .B2(n18346), .ZN(n18274) );
  OAI211_X1 U21367 ( .C1(n18581), .C2(n18598), .A(n18275), .B(n18274), .ZN(
        P3_U2876) );
  AOI22_X1 U21368 ( .A1(n18664), .A2(n18622), .B1(n18621), .B2(n18288), .ZN(
        n18277) );
  AOI22_X1 U21369 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18289), .B1(
        n18623), .B2(n18346), .ZN(n18276) );
  OAI211_X1 U21370 ( .C1(n18598), .C2(n18626), .A(n18277), .B(n18276), .ZN(
        P3_U2877) );
  INV_X1 U21371 ( .A(n18554), .ZN(n18628) );
  AOI22_X1 U21372 ( .A1(n18664), .A2(n18628), .B1(n18627), .B2(n18288), .ZN(
        n18279) );
  AOI22_X1 U21373 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18289), .B1(
        n18629), .B2(n18346), .ZN(n18278) );
  OAI211_X1 U21374 ( .C1(n18598), .C2(n18632), .A(n18279), .B(n18278), .ZN(
        P3_U2878) );
  AOI22_X1 U21375 ( .A1(n18605), .A2(n18634), .B1(n18633), .B2(n18288), .ZN(
        n18281) );
  AOI22_X1 U21376 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18289), .B1(
        n18635), .B2(n18346), .ZN(n18280) );
  OAI211_X1 U21377 ( .C1(n18312), .C2(n18638), .A(n18281), .B(n18280), .ZN(
        P3_U2879) );
  AOI22_X1 U21378 ( .A1(n18664), .A2(n18557), .B1(n18639), .B2(n18288), .ZN(
        n18283) );
  AOI22_X1 U21379 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18289), .B1(
        n18642), .B2(n18346), .ZN(n18282) );
  OAI211_X1 U21380 ( .C1(n18598), .C2(n18561), .A(n18283), .B(n18282), .ZN(
        P3_U2880) );
  AOI22_X1 U21381 ( .A1(n18664), .A2(n18648), .B1(n18647), .B2(n18288), .ZN(
        n18285) );
  AOI22_X1 U21382 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18289), .B1(
        n18649), .B2(n18346), .ZN(n18284) );
  OAI211_X1 U21383 ( .C1(n18598), .C2(n18652), .A(n18285), .B(n18284), .ZN(
        P3_U2881) );
  AOI22_X1 U21384 ( .A1(n18605), .A2(n18564), .B1(n18653), .B2(n18288), .ZN(
        n18287) );
  AOI22_X1 U21385 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18289), .B1(
        n18655), .B2(n18346), .ZN(n18286) );
  OAI211_X1 U21386 ( .C1(n18312), .C2(n18567), .A(n18287), .B(n18286), .ZN(
        P3_U2882) );
  AOI22_X1 U21387 ( .A1(n18605), .A2(n18604), .B1(n18660), .B2(n18288), .ZN(
        n18291) );
  AOI22_X1 U21388 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18289), .B1(
        n18663), .B2(n18346), .ZN(n18290) );
  OAI211_X1 U21389 ( .C1(n18312), .C2(n18609), .A(n18291), .B(n18290), .ZN(
        P3_U2883) );
  NAND2_X1 U21390 ( .A1(n18472), .A2(n18313), .ZN(n18378) );
  NOR2_X1 U21391 ( .A1(n18346), .A2(n18371), .ZN(n18334) );
  NOR2_X1 U21392 ( .A1(n9814), .A2(n18334), .ZN(n18308) );
  AOI22_X1 U21393 ( .A1(n18326), .A2(n18574), .B1(n18611), .B2(n18308), .ZN(
        n18295) );
  OAI21_X1 U21394 ( .B1(n18292), .B2(n18473), .A(n18334), .ZN(n18293) );
  OAI211_X1 U21395 ( .C1(n18371), .C2(n18863), .A(n18524), .B(n18293), .ZN(
        n18309) );
  AOI22_X1 U21396 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18309), .B1(
        n18617), .B2(n18371), .ZN(n18294) );
  OAI211_X1 U21397 ( .C1(n18581), .C2(n18312), .A(n18295), .B(n18294), .ZN(
        P3_U2884) );
  INV_X1 U21398 ( .A(n18623), .ZN(n18585) );
  AOI22_X1 U21399 ( .A1(n18664), .A2(n18582), .B1(n18621), .B2(n18308), .ZN(
        n18297) );
  AOI22_X1 U21400 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18309), .B1(
        n18326), .B2(n18622), .ZN(n18296) );
  OAI211_X1 U21401 ( .C1(n18585), .C2(n18378), .A(n18297), .B(n18296), .ZN(
        P3_U2885) );
  AOI22_X1 U21402 ( .A1(n18326), .A2(n18628), .B1(n18627), .B2(n18308), .ZN(
        n18299) );
  AOI22_X1 U21403 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18309), .B1(
        n18629), .B2(n18371), .ZN(n18298) );
  OAI211_X1 U21404 ( .C1(n18312), .C2(n18632), .A(n18299), .B(n18298), .ZN(
        P3_U2886) );
  AOI22_X1 U21405 ( .A1(n18664), .A2(n18634), .B1(n18633), .B2(n18308), .ZN(
        n18301) );
  AOI22_X1 U21406 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18309), .B1(
        n18635), .B2(n18371), .ZN(n18300) );
  OAI211_X1 U21407 ( .C1(n18333), .C2(n18638), .A(n18301), .B(n18300), .ZN(
        P3_U2887) );
  AOI22_X1 U21408 ( .A1(n18326), .A2(n18557), .B1(n18639), .B2(n18308), .ZN(
        n18303) );
  AOI22_X1 U21409 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18309), .B1(
        n18642), .B2(n18371), .ZN(n18302) );
  OAI211_X1 U21410 ( .C1(n18312), .C2(n18561), .A(n18303), .B(n18302), .ZN(
        P3_U2888) );
  AOI22_X1 U21411 ( .A1(n18664), .A2(n18594), .B1(n18647), .B2(n18308), .ZN(
        n18305) );
  AOI22_X1 U21412 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18309), .B1(
        n18326), .B2(n18648), .ZN(n18304) );
  OAI211_X1 U21413 ( .C1(n18597), .C2(n18378), .A(n18305), .B(n18304), .ZN(
        P3_U2889) );
  AOI22_X1 U21414 ( .A1(n18326), .A2(n18654), .B1(n18653), .B2(n18308), .ZN(
        n18307) );
  AOI22_X1 U21415 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18309), .B1(
        n18655), .B2(n18371), .ZN(n18306) );
  OAI211_X1 U21416 ( .C1(n18312), .C2(n18658), .A(n18307), .B(n18306), .ZN(
        P3_U2890) );
  INV_X1 U21417 ( .A(n18609), .ZN(n18661) );
  AOI22_X1 U21418 ( .A1(n18326), .A2(n18661), .B1(n18660), .B2(n18308), .ZN(
        n18311) );
  AOI22_X1 U21419 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18309), .B1(
        n18663), .B2(n18371), .ZN(n18310) );
  OAI211_X1 U21420 ( .C1(n18312), .C2(n18669), .A(n18311), .B(n18310), .ZN(
        P3_U2891) );
  NAND2_X1 U21421 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18313), .ZN(
        n18357) );
  NOR2_X1 U21422 ( .A1(n9814), .A2(n18357), .ZN(n18329) );
  AOI22_X1 U21423 ( .A1(n18612), .A2(n18326), .B1(n18611), .B2(n18329), .ZN(
        n18315) );
  NOR2_X2 U21424 ( .A1(n18518), .A2(n18357), .ZN(n18393) );
  AOI21_X1 U21425 ( .B1(n18699), .B2(n18473), .A(n18426), .ZN(n18403) );
  OAI211_X1 U21426 ( .C1(n18393), .C2(n18863), .A(n18313), .B(n18403), .ZN(
        n18330) );
  AOI22_X1 U21427 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18330), .B1(
        n18617), .B2(n18393), .ZN(n18314) );
  OAI211_X1 U21428 ( .C1(n18620), .C2(n18355), .A(n18315), .B(n18314), .ZN(
        P3_U2892) );
  AOI22_X1 U21429 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18330), .B1(
        n18621), .B2(n18329), .ZN(n18317) );
  AOI22_X1 U21430 ( .A1(n18623), .A2(n18393), .B1(n18622), .B2(n18346), .ZN(
        n18316) );
  OAI211_X1 U21431 ( .C1(n18333), .C2(n18626), .A(n18317), .B(n18316), .ZN(
        P3_U2893) );
  AOI22_X1 U21432 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18330), .B1(
        n18627), .B2(n18329), .ZN(n18319) );
  AOI22_X1 U21433 ( .A1(n18628), .A2(n18346), .B1(n18629), .B2(n18393), .ZN(
        n18318) );
  OAI211_X1 U21434 ( .C1(n18333), .C2(n18632), .A(n18319), .B(n18318), .ZN(
        P3_U2894) );
  AOI22_X1 U21435 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18330), .B1(
        n18633), .B2(n18329), .ZN(n18321) );
  INV_X1 U21436 ( .A(n18638), .ZN(n18588) );
  AOI22_X1 U21437 ( .A1(n18588), .A2(n18346), .B1(n18635), .B2(n18393), .ZN(
        n18320) );
  OAI211_X1 U21438 ( .C1(n18333), .C2(n18591), .A(n18321), .B(n18320), .ZN(
        P3_U2895) );
  AOI22_X1 U21439 ( .A1(n18557), .A2(n18346), .B1(n18639), .B2(n18329), .ZN(
        n18323) );
  AOI22_X1 U21440 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18330), .B1(
        n18642), .B2(n18393), .ZN(n18322) );
  OAI211_X1 U21441 ( .C1(n18333), .C2(n18561), .A(n18323), .B(n18322), .ZN(
        P3_U2896) );
  AOI22_X1 U21442 ( .A1(n18326), .A2(n18594), .B1(n18647), .B2(n18329), .ZN(
        n18325) );
  AOI22_X1 U21443 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18330), .B1(
        n18648), .B2(n18346), .ZN(n18324) );
  OAI211_X1 U21444 ( .C1(n18597), .C2(n18400), .A(n18325), .B(n18324), .ZN(
        P3_U2897) );
  AOI22_X1 U21445 ( .A1(n18326), .A2(n18564), .B1(n18653), .B2(n18329), .ZN(
        n18328) );
  AOI22_X1 U21446 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18330), .B1(
        n18655), .B2(n18393), .ZN(n18327) );
  OAI211_X1 U21447 ( .C1(n18567), .C2(n18355), .A(n18328), .B(n18327), .ZN(
        P3_U2898) );
  AOI22_X1 U21448 ( .A1(n18661), .A2(n18346), .B1(n18660), .B2(n18329), .ZN(
        n18332) );
  AOI22_X1 U21449 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18330), .B1(
        n18663), .B2(n18393), .ZN(n18331) );
  OAI211_X1 U21450 ( .C1(n18333), .C2(n18669), .A(n18332), .B(n18331), .ZN(
        P3_U2899) );
  INV_X1 U21451 ( .A(n18425), .ZN(n18701) );
  INV_X1 U21452 ( .A(n18409), .ZN(n18424) );
  AOI21_X1 U21453 ( .B1(n18424), .B2(n18400), .A(n9814), .ZN(n18351) );
  AOI22_X1 U21454 ( .A1(n18611), .A2(n18351), .B1(n18574), .B2(n18371), .ZN(
        n18337) );
  AOI221_X1 U21455 ( .B1(n18334), .B2(n18400), .C1(n18473), .C2(n18400), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18335) );
  OAI21_X1 U21456 ( .B1(n18409), .B2(n18335), .A(n18524), .ZN(n18352) );
  AOI22_X1 U21457 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18352), .B1(
        n18617), .B2(n18409), .ZN(n18336) );
  OAI211_X1 U21458 ( .C1(n18581), .C2(n18355), .A(n18337), .B(n18336), .ZN(
        P3_U2900) );
  AOI22_X1 U21459 ( .A1(n18622), .A2(n18371), .B1(n18621), .B2(n18351), .ZN(
        n18339) );
  AOI22_X1 U21460 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18352), .B1(
        n18623), .B2(n18409), .ZN(n18338) );
  OAI211_X1 U21461 ( .C1(n18626), .C2(n18355), .A(n18339), .B(n18338), .ZN(
        P3_U2901) );
  AOI22_X1 U21462 ( .A1(n18628), .A2(n18371), .B1(n18627), .B2(n18351), .ZN(
        n18341) );
  AOI22_X1 U21463 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18352), .B1(
        n18629), .B2(n18409), .ZN(n18340) );
  OAI211_X1 U21464 ( .C1(n18632), .C2(n18355), .A(n18341), .B(n18340), .ZN(
        P3_U2902) );
  AOI22_X1 U21465 ( .A1(n18588), .A2(n18371), .B1(n18633), .B2(n18351), .ZN(
        n18343) );
  AOI22_X1 U21466 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18352), .B1(
        n18635), .B2(n18409), .ZN(n18342) );
  OAI211_X1 U21467 ( .C1(n18591), .C2(n18355), .A(n18343), .B(n18342), .ZN(
        P3_U2903) );
  AOI22_X1 U21468 ( .A1(n18641), .A2(n18346), .B1(n18639), .B2(n18351), .ZN(
        n18345) );
  AOI22_X1 U21469 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18352), .B1(
        n18642), .B2(n18409), .ZN(n18344) );
  OAI211_X1 U21470 ( .C1(n18645), .C2(n18378), .A(n18345), .B(n18344), .ZN(
        P3_U2904) );
  AOI22_X1 U21471 ( .A1(n18594), .A2(n18346), .B1(n18647), .B2(n18351), .ZN(
        n18348) );
  AOI22_X1 U21472 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18352), .B1(
        n18648), .B2(n18371), .ZN(n18347) );
  OAI211_X1 U21473 ( .C1(n18597), .C2(n18424), .A(n18348), .B(n18347), .ZN(
        P3_U2905) );
  AOI22_X1 U21474 ( .A1(n18654), .A2(n18371), .B1(n18653), .B2(n18351), .ZN(
        n18350) );
  AOI22_X1 U21475 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18352), .B1(
        n18655), .B2(n18409), .ZN(n18349) );
  OAI211_X1 U21476 ( .C1(n18658), .C2(n18355), .A(n18350), .B(n18349), .ZN(
        P3_U2906) );
  AOI22_X1 U21477 ( .A1(n18661), .A2(n18371), .B1(n18660), .B2(n18351), .ZN(
        n18354) );
  AOI22_X1 U21478 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18352), .B1(
        n18663), .B2(n18409), .ZN(n18353) );
  OAI211_X1 U21479 ( .C1(n18669), .C2(n18355), .A(n18354), .B(n18353), .ZN(
        P3_U2907) );
  AOI22_X1 U21480 ( .A1(n18612), .A2(n18371), .B1(n18611), .B2(n18374), .ZN(
        n18360) );
  INV_X1 U21481 ( .A(n18357), .ZN(n18358) );
  AOI22_X1 U21482 ( .A1(n18616), .A2(n18358), .B1(n18450), .B2(n18404), .ZN(
        n18375) );
  NAND2_X1 U21483 ( .A1(n18452), .A2(n18404), .ZN(n18449) );
  AOI22_X1 U21484 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18375), .B1(
        n18617), .B2(n18441), .ZN(n18359) );
  OAI211_X1 U21485 ( .C1(n18620), .C2(n18400), .A(n18360), .B(n18359), .ZN(
        P3_U2908) );
  AOI22_X1 U21486 ( .A1(n18622), .A2(n18393), .B1(n18621), .B2(n18374), .ZN(
        n18362) );
  AOI22_X1 U21487 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18375), .B1(
        n18623), .B2(n18441), .ZN(n18361) );
  OAI211_X1 U21488 ( .C1(n18626), .C2(n18378), .A(n18362), .B(n18361), .ZN(
        P3_U2909) );
  AOI22_X1 U21489 ( .A1(n18627), .A2(n18374), .B1(n18551), .B2(n18371), .ZN(
        n18364) );
  AOI22_X1 U21490 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18375), .B1(
        n18629), .B2(n18441), .ZN(n18363) );
  OAI211_X1 U21491 ( .C1(n18554), .C2(n18400), .A(n18364), .B(n18363), .ZN(
        P3_U2910) );
  AOI22_X1 U21492 ( .A1(n18634), .A2(n18371), .B1(n18633), .B2(n18374), .ZN(
        n18366) );
  AOI22_X1 U21493 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18375), .B1(
        n18635), .B2(n18441), .ZN(n18365) );
  OAI211_X1 U21494 ( .C1(n18638), .C2(n18400), .A(n18366), .B(n18365), .ZN(
        P3_U2911) );
  AOI22_X1 U21495 ( .A1(n18641), .A2(n18371), .B1(n18639), .B2(n18374), .ZN(
        n18368) );
  AOI22_X1 U21496 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18375), .B1(
        n18642), .B2(n18441), .ZN(n18367) );
  OAI211_X1 U21497 ( .C1(n18645), .C2(n18400), .A(n18368), .B(n18367), .ZN(
        P3_U2912) );
  AOI22_X1 U21498 ( .A1(n18648), .A2(n18393), .B1(n18647), .B2(n18374), .ZN(
        n18370) );
  AOI22_X1 U21499 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18375), .B1(
        n18649), .B2(n18441), .ZN(n18369) );
  OAI211_X1 U21500 ( .C1(n18652), .C2(n18378), .A(n18370), .B(n18369), .ZN(
        P3_U2913) );
  AOI22_X1 U21501 ( .A1(n18564), .A2(n18371), .B1(n18653), .B2(n18374), .ZN(
        n18373) );
  AOI22_X1 U21502 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18375), .B1(
        n18655), .B2(n18441), .ZN(n18372) );
  OAI211_X1 U21503 ( .C1(n18567), .C2(n18400), .A(n18373), .B(n18372), .ZN(
        P3_U2914) );
  AOI22_X1 U21504 ( .A1(n18661), .A2(n18393), .B1(n18660), .B2(n18374), .ZN(
        n18377) );
  AOI22_X1 U21505 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18375), .B1(
        n18663), .B2(n18441), .ZN(n18376) );
  OAI211_X1 U21506 ( .C1(n18669), .C2(n18378), .A(n18377), .B(n18376), .ZN(
        P3_U2915) );
  NAND2_X1 U21507 ( .A1(n18472), .A2(n18404), .ZN(n18444) );
  NOR2_X1 U21508 ( .A1(n18441), .A2(n18468), .ZN(n18427) );
  NOR2_X1 U21509 ( .A1(n9814), .A2(n18427), .ZN(n18396) );
  AOI22_X1 U21510 ( .A1(n18612), .A2(n18393), .B1(n18611), .B2(n18396), .ZN(
        n18382) );
  NOR2_X1 U21511 ( .A1(n18409), .A2(n18393), .ZN(n18379) );
  OAI21_X1 U21512 ( .B1(n18379), .B2(n18473), .A(n18427), .ZN(n18380) );
  OAI211_X1 U21513 ( .C1(n18468), .C2(n18863), .A(n18524), .B(n18380), .ZN(
        n18397) );
  AOI22_X1 U21514 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18397), .B1(
        n18617), .B2(n18468), .ZN(n18381) );
  OAI211_X1 U21515 ( .C1(n18620), .C2(n18424), .A(n18382), .B(n18381), .ZN(
        P3_U2916) );
  AOI22_X1 U21516 ( .A1(n18582), .A2(n18393), .B1(n18621), .B2(n18396), .ZN(
        n18384) );
  AOI22_X1 U21517 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18397), .B1(
        n18622), .B2(n18409), .ZN(n18383) );
  OAI211_X1 U21518 ( .C1(n18585), .C2(n18444), .A(n18384), .B(n18383), .ZN(
        P3_U2917) );
  AOI22_X1 U21519 ( .A1(n18627), .A2(n18396), .B1(n18551), .B2(n18393), .ZN(
        n18386) );
  AOI22_X1 U21520 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18397), .B1(
        n18629), .B2(n18468), .ZN(n18385) );
  OAI211_X1 U21521 ( .C1(n18554), .C2(n18424), .A(n18386), .B(n18385), .ZN(
        P3_U2918) );
  AOI22_X1 U21522 ( .A1(n18634), .A2(n18393), .B1(n18633), .B2(n18396), .ZN(
        n18388) );
  AOI22_X1 U21523 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18397), .B1(
        n18635), .B2(n18468), .ZN(n18387) );
  OAI211_X1 U21524 ( .C1(n18638), .C2(n18424), .A(n18388), .B(n18387), .ZN(
        P3_U2919) );
  AOI22_X1 U21525 ( .A1(n18557), .A2(n18409), .B1(n18639), .B2(n18396), .ZN(
        n18390) );
  AOI22_X1 U21526 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18397), .B1(
        n18642), .B2(n18468), .ZN(n18389) );
  OAI211_X1 U21527 ( .C1(n18561), .C2(n18400), .A(n18390), .B(n18389), .ZN(
        P3_U2920) );
  AOI22_X1 U21528 ( .A1(n18594), .A2(n18393), .B1(n18647), .B2(n18396), .ZN(
        n18392) );
  AOI22_X1 U21529 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18397), .B1(
        n18648), .B2(n18409), .ZN(n18391) );
  OAI211_X1 U21530 ( .C1(n18597), .C2(n18444), .A(n18392), .B(n18391), .ZN(
        P3_U2921) );
  AOI22_X1 U21531 ( .A1(n18564), .A2(n18393), .B1(n18653), .B2(n18396), .ZN(
        n18395) );
  AOI22_X1 U21532 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18397), .B1(
        n18655), .B2(n18468), .ZN(n18394) );
  OAI211_X1 U21533 ( .C1(n18567), .C2(n18424), .A(n18395), .B(n18394), .ZN(
        P3_U2922) );
  AOI22_X1 U21534 ( .A1(n18661), .A2(n18409), .B1(n18660), .B2(n18396), .ZN(
        n18399) );
  AOI22_X1 U21535 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18397), .B1(
        n18663), .B2(n18468), .ZN(n18398) );
  OAI211_X1 U21536 ( .C1(n18669), .C2(n18400), .A(n18399), .B(n18398), .ZN(
        P3_U2923) );
  NOR2_X1 U21537 ( .A1(n18401), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18451) );
  INV_X1 U21538 ( .A(n18451), .ZN(n18402) );
  NOR2_X1 U21539 ( .A1(n9814), .A2(n18402), .ZN(n18420) );
  AOI22_X1 U21540 ( .A1(n18612), .A2(n18409), .B1(n18611), .B2(n18420), .ZN(
        n18406) );
  NAND2_X1 U21541 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18451), .ZN(
        n18490) );
  INV_X1 U21542 ( .A(n18490), .ZN(n18492) );
  OAI211_X1 U21543 ( .C1(n18492), .C2(n18863), .A(n18404), .B(n18403), .ZN(
        n18421) );
  AOI22_X1 U21544 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18421), .B1(
        n18617), .B2(n18492), .ZN(n18405) );
  OAI211_X1 U21545 ( .C1(n18620), .C2(n18449), .A(n18406), .B(n18405), .ZN(
        P3_U2924) );
  AOI22_X1 U21546 ( .A1(n18582), .A2(n18409), .B1(n18621), .B2(n18420), .ZN(
        n18408) );
  AOI22_X1 U21547 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18421), .B1(
        n18622), .B2(n18441), .ZN(n18407) );
  OAI211_X1 U21548 ( .C1(n18585), .C2(n18490), .A(n18408), .B(n18407), .ZN(
        P3_U2925) );
  AOI22_X1 U21549 ( .A1(n18627), .A2(n18420), .B1(n18551), .B2(n18409), .ZN(
        n18411) );
  AOI22_X1 U21550 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18421), .B1(
        n18629), .B2(n18492), .ZN(n18410) );
  OAI211_X1 U21551 ( .C1(n18554), .C2(n18449), .A(n18411), .B(n18410), .ZN(
        P3_U2926) );
  AOI22_X1 U21552 ( .A1(n18634), .A2(n18409), .B1(n18633), .B2(n18420), .ZN(
        n18413) );
  AOI22_X1 U21553 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18421), .B1(
        n18635), .B2(n18492), .ZN(n18412) );
  OAI211_X1 U21554 ( .C1(n18638), .C2(n18449), .A(n18413), .B(n18412), .ZN(
        P3_U2927) );
  AOI22_X1 U21555 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18421), .B1(
        n18639), .B2(n18420), .ZN(n18415) );
  AOI22_X1 U21556 ( .A1(n18641), .A2(n18409), .B1(n18642), .B2(n18492), .ZN(
        n18414) );
  OAI211_X1 U21557 ( .C1(n18645), .C2(n18449), .A(n18415), .B(n18414), .ZN(
        P3_U2928) );
  AOI22_X1 U21558 ( .A1(n18594), .A2(n18409), .B1(n18647), .B2(n18420), .ZN(
        n18417) );
  AOI22_X1 U21559 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18421), .B1(
        n18648), .B2(n18441), .ZN(n18416) );
  OAI211_X1 U21560 ( .C1(n18597), .C2(n18490), .A(n18417), .B(n18416), .ZN(
        P3_U2929) );
  AOI22_X1 U21561 ( .A1(n18564), .A2(n18409), .B1(n18653), .B2(n18420), .ZN(
        n18419) );
  AOI22_X1 U21562 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18421), .B1(
        n18655), .B2(n18492), .ZN(n18418) );
  OAI211_X1 U21563 ( .C1(n18567), .C2(n18449), .A(n18419), .B(n18418), .ZN(
        P3_U2930) );
  AOI22_X1 U21564 ( .A1(n18661), .A2(n18441), .B1(n18660), .B2(n18420), .ZN(
        n18423) );
  AOI22_X1 U21565 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18421), .B1(
        n18663), .B2(n18492), .ZN(n18422) );
  OAI211_X1 U21566 ( .C1(n18669), .C2(n18424), .A(n18423), .B(n18422), .ZN(
        P3_U2931) );
  NAND2_X1 U21567 ( .A1(n18425), .A2(n18519), .ZN(n18517) );
  NOR2_X1 U21568 ( .A1(n18510), .A2(n18492), .ZN(n18474) );
  NOR2_X1 U21569 ( .A1(n9814), .A2(n18474), .ZN(n18445) );
  AOI22_X1 U21570 ( .A1(n18612), .A2(n18441), .B1(n18611), .B2(n18445), .ZN(
        n18430) );
  OAI22_X1 U21571 ( .A1(n18427), .A2(n18575), .B1(n18474), .B2(n18426), .ZN(
        n18428) );
  OAI21_X1 U21572 ( .B1(n18510), .B2(n18863), .A(n18428), .ZN(n18446) );
  AOI22_X1 U21573 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18446), .B1(
        n18617), .B2(n18510), .ZN(n18429) );
  OAI211_X1 U21574 ( .C1(n18620), .C2(n18444), .A(n18430), .B(n18429), .ZN(
        P3_U2932) );
  AOI22_X1 U21575 ( .A1(n18582), .A2(n18441), .B1(n18621), .B2(n18445), .ZN(
        n18432) );
  AOI22_X1 U21576 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18446), .B1(
        n18622), .B2(n18468), .ZN(n18431) );
  OAI211_X1 U21577 ( .C1(n18585), .C2(n18517), .A(n18432), .B(n18431), .ZN(
        P3_U2933) );
  AOI22_X1 U21578 ( .A1(n18628), .A2(n18468), .B1(n18627), .B2(n18445), .ZN(
        n18434) );
  AOI22_X1 U21579 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18446), .B1(
        n18629), .B2(n18510), .ZN(n18433) );
  OAI211_X1 U21580 ( .C1(n18632), .C2(n18449), .A(n18434), .B(n18433), .ZN(
        P3_U2934) );
  AOI22_X1 U21581 ( .A1(n18634), .A2(n18441), .B1(n18633), .B2(n18445), .ZN(
        n18436) );
  AOI22_X1 U21582 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18446), .B1(
        n18635), .B2(n18510), .ZN(n18435) );
  OAI211_X1 U21583 ( .C1(n18638), .C2(n18444), .A(n18436), .B(n18435), .ZN(
        P3_U2935) );
  AOI22_X1 U21584 ( .A1(n18641), .A2(n18441), .B1(n18639), .B2(n18445), .ZN(
        n18438) );
  AOI22_X1 U21585 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18446), .B1(
        n18642), .B2(n18510), .ZN(n18437) );
  OAI211_X1 U21586 ( .C1(n18645), .C2(n18444), .A(n18438), .B(n18437), .ZN(
        P3_U2936) );
  AOI22_X1 U21587 ( .A1(n18594), .A2(n18441), .B1(n18647), .B2(n18445), .ZN(
        n18440) );
  AOI22_X1 U21588 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18446), .B1(
        n18648), .B2(n18468), .ZN(n18439) );
  OAI211_X1 U21589 ( .C1(n18597), .C2(n18517), .A(n18440), .B(n18439), .ZN(
        P3_U2937) );
  AOI22_X1 U21590 ( .A1(n18564), .A2(n18441), .B1(n18653), .B2(n18445), .ZN(
        n18443) );
  AOI22_X1 U21591 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18446), .B1(
        n18655), .B2(n18510), .ZN(n18442) );
  OAI211_X1 U21592 ( .C1(n18567), .C2(n18444), .A(n18443), .B(n18442), .ZN(
        P3_U2938) );
  AOI22_X1 U21593 ( .A1(n18661), .A2(n18468), .B1(n18660), .B2(n18445), .ZN(
        n18448) );
  AOI22_X1 U21594 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18446), .B1(
        n18663), .B2(n18510), .ZN(n18447) );
  OAI211_X1 U21595 ( .C1(n18669), .C2(n18449), .A(n18448), .B(n18447), .ZN(
        P3_U2939) );
  INV_X1 U21596 ( .A(n18519), .ZN(n18496) );
  AOI22_X1 U21597 ( .A1(n18612), .A2(n18468), .B1(n18611), .B2(n18467), .ZN(
        n18454) );
  AOI22_X1 U21598 ( .A1(n18616), .A2(n18451), .B1(n18450), .B2(n18519), .ZN(
        n18469) );
  NAND2_X1 U21599 ( .A1(n18452), .A2(n18519), .ZN(n18544) );
  INV_X1 U21600 ( .A(n18544), .ZN(n18537) );
  AOI22_X1 U21601 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18469), .B1(
        n18617), .B2(n18537), .ZN(n18453) );
  OAI211_X1 U21602 ( .C1(n18620), .C2(n18490), .A(n18454), .B(n18453), .ZN(
        P3_U2940) );
  AOI22_X1 U21603 ( .A1(n18582), .A2(n18468), .B1(n18621), .B2(n18467), .ZN(
        n18456) );
  AOI22_X1 U21604 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18469), .B1(
        n18622), .B2(n18492), .ZN(n18455) );
  OAI211_X1 U21605 ( .C1(n18585), .C2(n18544), .A(n18456), .B(n18455), .ZN(
        P3_U2941) );
  AOI22_X1 U21606 ( .A1(n18627), .A2(n18467), .B1(n18551), .B2(n18468), .ZN(
        n18458) );
  AOI22_X1 U21607 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18469), .B1(
        n18629), .B2(n18537), .ZN(n18457) );
  OAI211_X1 U21608 ( .C1(n18554), .C2(n18490), .A(n18458), .B(n18457), .ZN(
        P3_U2942) );
  AOI22_X1 U21609 ( .A1(n18634), .A2(n18468), .B1(n18633), .B2(n18467), .ZN(
        n18460) );
  AOI22_X1 U21610 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18469), .B1(
        n18635), .B2(n18537), .ZN(n18459) );
  OAI211_X1 U21611 ( .C1(n18638), .C2(n18490), .A(n18460), .B(n18459), .ZN(
        P3_U2943) );
  AOI22_X1 U21612 ( .A1(n18641), .A2(n18468), .B1(n18639), .B2(n18467), .ZN(
        n18462) );
  AOI22_X1 U21613 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18469), .B1(
        n18642), .B2(n18537), .ZN(n18461) );
  OAI211_X1 U21614 ( .C1(n18645), .C2(n18490), .A(n18462), .B(n18461), .ZN(
        P3_U2944) );
  AOI22_X1 U21615 ( .A1(n18594), .A2(n18468), .B1(n18647), .B2(n18467), .ZN(
        n18464) );
  AOI22_X1 U21616 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18469), .B1(
        n18648), .B2(n18492), .ZN(n18463) );
  OAI211_X1 U21617 ( .C1(n18597), .C2(n18544), .A(n18464), .B(n18463), .ZN(
        P3_U2945) );
  AOI22_X1 U21618 ( .A1(n18564), .A2(n18468), .B1(n18653), .B2(n18467), .ZN(
        n18466) );
  AOI22_X1 U21619 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18469), .B1(
        n18655), .B2(n18537), .ZN(n18465) );
  OAI211_X1 U21620 ( .C1(n18567), .C2(n18490), .A(n18466), .B(n18465), .ZN(
        P3_U2946) );
  AOI22_X1 U21621 ( .A1(n18604), .A2(n18468), .B1(n18660), .B2(n18467), .ZN(
        n18471) );
  AOI22_X1 U21622 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18469), .B1(
        n18663), .B2(n18537), .ZN(n18470) );
  OAI211_X1 U21623 ( .C1(n18609), .C2(n18490), .A(n18471), .B(n18470), .ZN(
        P3_U2947) );
  AOI22_X1 U21624 ( .A1(n18611), .A2(n18491), .B1(n18574), .B2(n18510), .ZN(
        n18477) );
  NAND2_X1 U21625 ( .A1(n18472), .A2(n18519), .ZN(n18560) );
  AOI221_X1 U21626 ( .B1(n18474), .B2(n18544), .C1(n18473), .C2(n18544), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18475) );
  OAI21_X1 U21627 ( .B1(n18569), .B2(n18475), .A(n18524), .ZN(n18493) );
  AOI22_X1 U21628 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18493), .B1(
        n18617), .B2(n18569), .ZN(n18476) );
  OAI211_X1 U21629 ( .C1(n18581), .C2(n18490), .A(n18477), .B(n18476), .ZN(
        P3_U2948) );
  AOI22_X1 U21630 ( .A1(n18622), .A2(n18510), .B1(n18621), .B2(n18491), .ZN(
        n18479) );
  AOI22_X1 U21631 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18493), .B1(
        n18623), .B2(n18569), .ZN(n18478) );
  OAI211_X1 U21632 ( .C1(n18626), .C2(n18490), .A(n18479), .B(n18478), .ZN(
        P3_U2949) );
  AOI22_X1 U21633 ( .A1(n18627), .A2(n18491), .B1(n18551), .B2(n18492), .ZN(
        n18481) );
  AOI22_X1 U21634 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18493), .B1(
        n18629), .B2(n18569), .ZN(n18480) );
  OAI211_X1 U21635 ( .C1(n18554), .C2(n18517), .A(n18481), .B(n18480), .ZN(
        P3_U2950) );
  AOI22_X1 U21636 ( .A1(n18634), .A2(n18492), .B1(n18633), .B2(n18491), .ZN(
        n18483) );
  AOI22_X1 U21637 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18493), .B1(
        n18635), .B2(n18569), .ZN(n18482) );
  OAI211_X1 U21638 ( .C1(n18638), .C2(n18517), .A(n18483), .B(n18482), .ZN(
        P3_U2951) );
  AOI22_X1 U21639 ( .A1(n18557), .A2(n18510), .B1(n18639), .B2(n18491), .ZN(
        n18485) );
  AOI22_X1 U21640 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18493), .B1(
        n18642), .B2(n18569), .ZN(n18484) );
  OAI211_X1 U21641 ( .C1(n18561), .C2(n18490), .A(n18485), .B(n18484), .ZN(
        P3_U2952) );
  AOI22_X1 U21642 ( .A1(n18594), .A2(n18492), .B1(n18647), .B2(n18491), .ZN(
        n18487) );
  AOI22_X1 U21643 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18493), .B1(
        n18648), .B2(n18510), .ZN(n18486) );
  OAI211_X1 U21644 ( .C1(n18597), .C2(n18560), .A(n18487), .B(n18486), .ZN(
        P3_U2953) );
  AOI22_X1 U21645 ( .A1(n18654), .A2(n18510), .B1(n18653), .B2(n18491), .ZN(
        n18489) );
  AOI22_X1 U21646 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18493), .B1(
        n18655), .B2(n18569), .ZN(n18488) );
  OAI211_X1 U21647 ( .C1(n18658), .C2(n18490), .A(n18489), .B(n18488), .ZN(
        P3_U2954) );
  AOI22_X1 U21648 ( .A1(n18604), .A2(n18492), .B1(n18660), .B2(n18491), .ZN(
        n18495) );
  AOI22_X1 U21649 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18493), .B1(
        n18663), .B2(n18569), .ZN(n18494) );
  OAI211_X1 U21650 ( .C1(n18609), .C2(n18517), .A(n18495), .B(n18494), .ZN(
        P3_U2955) );
  NOR2_X1 U21651 ( .A1(n18699), .A2(n18496), .ZN(n18546) );
  INV_X1 U21652 ( .A(n18546), .ZN(n18497) );
  NOR2_X1 U21653 ( .A1(n9814), .A2(n18497), .ZN(n18513) );
  AOI22_X1 U21654 ( .A1(n18611), .A2(n18513), .B1(n18574), .B2(n18537), .ZN(
        n18499) );
  OAI211_X1 U21655 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18616), .A(
        n18613), .B(n18519), .ZN(n18514) );
  NAND2_X1 U21656 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18546), .ZN(
        n18601) );
  AOI22_X1 U21657 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18514), .B1(
        n18617), .B2(n18603), .ZN(n18498) );
  OAI211_X1 U21658 ( .C1(n18581), .C2(n18517), .A(n18499), .B(n18498), .ZN(
        P3_U2956) );
  AOI22_X1 U21659 ( .A1(n18622), .A2(n18537), .B1(n18621), .B2(n18513), .ZN(
        n18501) );
  AOI22_X1 U21660 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18514), .B1(
        n18623), .B2(n18603), .ZN(n18500) );
  OAI211_X1 U21661 ( .C1(n18626), .C2(n18517), .A(n18501), .B(n18500), .ZN(
        P3_U2957) );
  AOI22_X1 U21662 ( .A1(n18627), .A2(n18513), .B1(n18551), .B2(n18510), .ZN(
        n18503) );
  AOI22_X1 U21663 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18514), .B1(
        n18629), .B2(n18603), .ZN(n18502) );
  OAI211_X1 U21664 ( .C1(n18554), .C2(n18544), .A(n18503), .B(n18502), .ZN(
        P3_U2958) );
  AOI22_X1 U21665 ( .A1(n18588), .A2(n18537), .B1(n18633), .B2(n18513), .ZN(
        n18505) );
  AOI22_X1 U21666 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18514), .B1(
        n18635), .B2(n18603), .ZN(n18504) );
  OAI211_X1 U21667 ( .C1(n18591), .C2(n18517), .A(n18505), .B(n18504), .ZN(
        P3_U2959) );
  AOI22_X1 U21668 ( .A1(n18641), .A2(n18510), .B1(n18639), .B2(n18513), .ZN(
        n18507) );
  AOI22_X1 U21669 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18514), .B1(
        n18642), .B2(n18603), .ZN(n18506) );
  OAI211_X1 U21670 ( .C1(n18645), .C2(n18544), .A(n18507), .B(n18506), .ZN(
        P3_U2960) );
  AOI22_X1 U21671 ( .A1(n18594), .A2(n18510), .B1(n18647), .B2(n18513), .ZN(
        n18509) );
  AOI22_X1 U21672 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18514), .B1(
        n18648), .B2(n18537), .ZN(n18508) );
  OAI211_X1 U21673 ( .C1(n18597), .C2(n18601), .A(n18509), .B(n18508), .ZN(
        P3_U2961) );
  AOI22_X1 U21674 ( .A1(n18564), .A2(n18510), .B1(n18653), .B2(n18513), .ZN(
        n18512) );
  AOI22_X1 U21675 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18514), .B1(
        n18655), .B2(n18603), .ZN(n18511) );
  OAI211_X1 U21676 ( .C1(n18567), .C2(n18544), .A(n18512), .B(n18511), .ZN(
        P3_U2962) );
  AOI22_X1 U21677 ( .A1(n18661), .A2(n18537), .B1(n18660), .B2(n18513), .ZN(
        n18516) );
  AOI22_X1 U21678 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18514), .B1(
        n18663), .B2(n18603), .ZN(n18515) );
  OAI211_X1 U21679 ( .C1(n18669), .C2(n18517), .A(n18516), .B(n18515), .ZN(
        P3_U2963) );
  INV_X1 U21680 ( .A(n18545), .ZN(n18615) );
  NAND2_X1 U21681 ( .A1(n18518), .A2(n18615), .ZN(n18668) );
  INV_X1 U21682 ( .A(n18668), .ZN(n18640) );
  NOR2_X1 U21683 ( .A1(n18603), .A2(n18640), .ZN(n18576) );
  NOR2_X1 U21684 ( .A1(n9814), .A2(n18576), .ZN(n18540) );
  AOI22_X1 U21685 ( .A1(n18611), .A2(n18540), .B1(n18574), .B2(n18569), .ZN(
        n18526) );
  NAND2_X1 U21686 ( .A1(n18520), .A2(n18519), .ZN(n18521) );
  OAI21_X1 U21687 ( .B1(n18522), .B2(n18521), .A(n18576), .ZN(n18523) );
  OAI211_X1 U21688 ( .C1(n18640), .C2(n18863), .A(n18524), .B(n18523), .ZN(
        n18541) );
  AOI22_X1 U21689 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18541), .B1(
        n18617), .B2(n18640), .ZN(n18525) );
  OAI211_X1 U21690 ( .C1(n18581), .C2(n18544), .A(n18526), .B(n18525), .ZN(
        P3_U2964) );
  AOI22_X1 U21691 ( .A1(n18582), .A2(n18537), .B1(n18621), .B2(n18540), .ZN(
        n18528) );
  AOI22_X1 U21692 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18541), .B1(
        n18622), .B2(n18569), .ZN(n18527) );
  OAI211_X1 U21693 ( .C1(n18585), .C2(n18668), .A(n18528), .B(n18527), .ZN(
        P3_U2965) );
  AOI22_X1 U21694 ( .A1(n18628), .A2(n18569), .B1(n18627), .B2(n18540), .ZN(
        n18530) );
  AOI22_X1 U21695 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18541), .B1(
        n18629), .B2(n18640), .ZN(n18529) );
  OAI211_X1 U21696 ( .C1(n18632), .C2(n18544), .A(n18530), .B(n18529), .ZN(
        P3_U2966) );
  AOI22_X1 U21697 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18541), .B1(
        n18633), .B2(n18540), .ZN(n18532) );
  AOI22_X1 U21698 ( .A1(n18635), .A2(n18640), .B1(n18634), .B2(n18537), .ZN(
        n18531) );
  OAI211_X1 U21699 ( .C1(n18638), .C2(n18560), .A(n18532), .B(n18531), .ZN(
        P3_U2967) );
  AOI22_X1 U21700 ( .A1(n18641), .A2(n18537), .B1(n18639), .B2(n18540), .ZN(
        n18534) );
  AOI22_X1 U21701 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18541), .B1(
        n18642), .B2(n18640), .ZN(n18533) );
  OAI211_X1 U21702 ( .C1(n18645), .C2(n18560), .A(n18534), .B(n18533), .ZN(
        P3_U2968) );
  AOI22_X1 U21703 ( .A1(n18648), .A2(n18569), .B1(n18647), .B2(n18540), .ZN(
        n18536) );
  AOI22_X1 U21704 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18541), .B1(
        n18649), .B2(n18640), .ZN(n18535) );
  OAI211_X1 U21705 ( .C1(n18652), .C2(n18544), .A(n18536), .B(n18535), .ZN(
        P3_U2969) );
  AOI22_X1 U21706 ( .A1(n18564), .A2(n18537), .B1(n18653), .B2(n18540), .ZN(
        n18539) );
  AOI22_X1 U21707 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18541), .B1(
        n18655), .B2(n18640), .ZN(n18538) );
  OAI211_X1 U21708 ( .C1(n18567), .C2(n18560), .A(n18539), .B(n18538), .ZN(
        P3_U2970) );
  AOI22_X1 U21709 ( .A1(n18661), .A2(n18569), .B1(n18660), .B2(n18540), .ZN(
        n18543) );
  AOI22_X1 U21710 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18541), .B1(
        n18663), .B2(n18640), .ZN(n18542) );
  OAI211_X1 U21711 ( .C1(n18669), .C2(n18544), .A(n18543), .B(n18542), .ZN(
        P3_U2971) );
  NOR2_X1 U21712 ( .A1(n9814), .A2(n18545), .ZN(n18568) );
  AOI22_X1 U21713 ( .A1(n18611), .A2(n18568), .B1(n18574), .B2(n18603), .ZN(
        n18548) );
  AOI22_X1 U21714 ( .A1(n18616), .A2(n18546), .B1(n18615), .B2(n18613), .ZN(
        n18570) );
  AOI22_X1 U21715 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18570), .B1(
        n18662), .B2(n18617), .ZN(n18547) );
  OAI211_X1 U21716 ( .C1(n18581), .C2(n18560), .A(n18548), .B(n18547), .ZN(
        P3_U2972) );
  AOI22_X1 U21717 ( .A1(n18582), .A2(n18569), .B1(n18621), .B2(n18568), .ZN(
        n18550) );
  AOI22_X1 U21718 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18570), .B1(
        n18622), .B2(n18603), .ZN(n18549) );
  OAI211_X1 U21719 ( .C1(n18646), .C2(n18585), .A(n18550), .B(n18549), .ZN(
        P3_U2973) );
  AOI22_X1 U21720 ( .A1(n18627), .A2(n18568), .B1(n18551), .B2(n18569), .ZN(
        n18553) );
  AOI22_X1 U21721 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18570), .B1(
        n18662), .B2(n18629), .ZN(n18552) );
  OAI211_X1 U21722 ( .C1(n18554), .C2(n18601), .A(n18553), .B(n18552), .ZN(
        P3_U2974) );
  AOI22_X1 U21723 ( .A1(n18634), .A2(n18569), .B1(n18633), .B2(n18568), .ZN(
        n18556) );
  AOI22_X1 U21724 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18570), .B1(
        n18662), .B2(n18635), .ZN(n18555) );
  OAI211_X1 U21725 ( .C1(n18638), .C2(n18601), .A(n18556), .B(n18555), .ZN(
        P3_U2975) );
  AOI22_X1 U21726 ( .A1(n18557), .A2(n18603), .B1(n18639), .B2(n18568), .ZN(
        n18559) );
  AOI22_X1 U21727 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18570), .B1(
        n18662), .B2(n18642), .ZN(n18558) );
  OAI211_X1 U21728 ( .C1(n18561), .C2(n18560), .A(n18559), .B(n18558), .ZN(
        P3_U2976) );
  AOI22_X1 U21729 ( .A1(n18594), .A2(n18569), .B1(n18647), .B2(n18568), .ZN(
        n18563) );
  AOI22_X1 U21730 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18570), .B1(
        n18648), .B2(n18603), .ZN(n18562) );
  OAI211_X1 U21731 ( .C1(n18646), .C2(n18597), .A(n18563), .B(n18562), .ZN(
        P3_U2977) );
  AOI22_X1 U21732 ( .A1(n18564), .A2(n18569), .B1(n18653), .B2(n18568), .ZN(
        n18566) );
  AOI22_X1 U21733 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18570), .B1(
        n18662), .B2(n18655), .ZN(n18565) );
  OAI211_X1 U21734 ( .C1(n18567), .C2(n18601), .A(n18566), .B(n18565), .ZN(
        P3_U2978) );
  AOI22_X1 U21735 ( .A1(n18604), .A2(n18569), .B1(n18660), .B2(n18568), .ZN(
        n18572) );
  AOI22_X1 U21736 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18570), .B1(
        n18662), .B2(n18663), .ZN(n18571) );
  OAI211_X1 U21737 ( .C1(n18609), .C2(n18601), .A(n18572), .B(n18571), .ZN(
        P3_U2979) );
  NOR2_X1 U21738 ( .A1(n9814), .A2(n18573), .ZN(n18602) );
  AOI22_X1 U21739 ( .A1(n18611), .A2(n18602), .B1(n18574), .B2(n18640), .ZN(
        n18580) );
  NOR2_X1 U21740 ( .A1(n18576), .A2(n18575), .ZN(n18577) );
  OAI22_X1 U21741 ( .A1(n18578), .A2(n18577), .B1(n18605), .B2(n18863), .ZN(
        n18606) );
  AOI22_X1 U21742 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18606), .B1(
        n18617), .B2(n18605), .ZN(n18579) );
  OAI211_X1 U21743 ( .C1(n18581), .C2(n18601), .A(n18580), .B(n18579), .ZN(
        P3_U2980) );
  AOI22_X1 U21744 ( .A1(n18582), .A2(n18603), .B1(n18621), .B2(n18602), .ZN(
        n18584) );
  AOI22_X1 U21745 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18606), .B1(
        n18622), .B2(n18640), .ZN(n18583) );
  OAI211_X1 U21746 ( .C1(n18598), .C2(n18585), .A(n18584), .B(n18583), .ZN(
        P3_U2981) );
  AOI22_X1 U21747 ( .A1(n18628), .A2(n18640), .B1(n18627), .B2(n18602), .ZN(
        n18587) );
  AOI22_X1 U21748 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18606), .B1(
        n18605), .B2(n18629), .ZN(n18586) );
  OAI211_X1 U21749 ( .C1(n18632), .C2(n18601), .A(n18587), .B(n18586), .ZN(
        P3_U2982) );
  AOI22_X1 U21750 ( .A1(n18588), .A2(n18640), .B1(n18633), .B2(n18602), .ZN(
        n18590) );
  AOI22_X1 U21751 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18606), .B1(
        n18605), .B2(n18635), .ZN(n18589) );
  OAI211_X1 U21752 ( .C1(n18591), .C2(n18601), .A(n18590), .B(n18589), .ZN(
        P3_U2983) );
  AOI22_X1 U21753 ( .A1(n18641), .A2(n18603), .B1(n18639), .B2(n18602), .ZN(
        n18593) );
  AOI22_X1 U21754 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18606), .B1(
        n18605), .B2(n18642), .ZN(n18592) );
  OAI211_X1 U21755 ( .C1(n18645), .C2(n18668), .A(n18593), .B(n18592), .ZN(
        P3_U2984) );
  AOI22_X1 U21756 ( .A1(n18594), .A2(n18603), .B1(n18647), .B2(n18602), .ZN(
        n18596) );
  AOI22_X1 U21757 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18606), .B1(
        n18648), .B2(n18640), .ZN(n18595) );
  OAI211_X1 U21758 ( .C1(n18598), .C2(n18597), .A(n18596), .B(n18595), .ZN(
        P3_U2985) );
  AOI22_X1 U21759 ( .A1(n18654), .A2(n18640), .B1(n18653), .B2(n18602), .ZN(
        n18600) );
  AOI22_X1 U21760 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18606), .B1(
        n18605), .B2(n18655), .ZN(n18599) );
  OAI211_X1 U21761 ( .C1(n18658), .C2(n18601), .A(n18600), .B(n18599), .ZN(
        P3_U2986) );
  AOI22_X1 U21762 ( .A1(n18604), .A2(n18603), .B1(n18660), .B2(n18602), .ZN(
        n18608) );
  AOI22_X1 U21763 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18606), .B1(
        n18605), .B2(n18663), .ZN(n18607) );
  OAI211_X1 U21764 ( .C1(n18609), .C2(n18668), .A(n18608), .B(n18607), .ZN(
        P3_U2987) );
  INV_X1 U21765 ( .A(n18614), .ZN(n18610) );
  NOR2_X1 U21766 ( .A1(n9814), .A2(n18610), .ZN(n18659) );
  AOI22_X1 U21767 ( .A1(n18612), .A2(n18640), .B1(n18611), .B2(n18659), .ZN(
        n18619) );
  AOI22_X1 U21768 ( .A1(n18616), .A2(n18615), .B1(n18614), .B2(n18613), .ZN(
        n18665) );
  AOI22_X1 U21769 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18665), .B1(
        n18664), .B2(n18617), .ZN(n18618) );
  OAI211_X1 U21770 ( .C1(n18646), .C2(n18620), .A(n18619), .B(n18618), .ZN(
        P3_U2988) );
  AOI22_X1 U21771 ( .A1(n18662), .A2(n18622), .B1(n18621), .B2(n18659), .ZN(
        n18625) );
  AOI22_X1 U21772 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18665), .B1(
        n18664), .B2(n18623), .ZN(n18624) );
  OAI211_X1 U21773 ( .C1(n18626), .C2(n18668), .A(n18625), .B(n18624), .ZN(
        P3_U2989) );
  AOI22_X1 U21774 ( .A1(n18662), .A2(n18628), .B1(n18627), .B2(n18659), .ZN(
        n18631) );
  AOI22_X1 U21775 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18665), .B1(
        n18664), .B2(n18629), .ZN(n18630) );
  OAI211_X1 U21776 ( .C1(n18632), .C2(n18668), .A(n18631), .B(n18630), .ZN(
        P3_U2990) );
  AOI22_X1 U21777 ( .A1(n18634), .A2(n18640), .B1(n18633), .B2(n18659), .ZN(
        n18637) );
  AOI22_X1 U21778 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18665), .B1(
        n18664), .B2(n18635), .ZN(n18636) );
  OAI211_X1 U21779 ( .C1(n18646), .C2(n18638), .A(n18637), .B(n18636), .ZN(
        P3_U2991) );
  AOI22_X1 U21780 ( .A1(n18641), .A2(n18640), .B1(n18639), .B2(n18659), .ZN(
        n18644) );
  AOI22_X1 U21781 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18665), .B1(
        n18664), .B2(n18642), .ZN(n18643) );
  OAI211_X1 U21782 ( .C1(n18646), .C2(n18645), .A(n18644), .B(n18643), .ZN(
        P3_U2992) );
  AOI22_X1 U21783 ( .A1(n18662), .A2(n18648), .B1(n18647), .B2(n18659), .ZN(
        n18651) );
  AOI22_X1 U21784 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18665), .B1(
        n18664), .B2(n18649), .ZN(n18650) );
  OAI211_X1 U21785 ( .C1(n18652), .C2(n18668), .A(n18651), .B(n18650), .ZN(
        P3_U2993) );
  AOI22_X1 U21786 ( .A1(n18662), .A2(n18654), .B1(n18653), .B2(n18659), .ZN(
        n18657) );
  AOI22_X1 U21787 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18665), .B1(
        n18664), .B2(n18655), .ZN(n18656) );
  OAI211_X1 U21788 ( .C1(n18658), .C2(n18668), .A(n18657), .B(n18656), .ZN(
        P3_U2994) );
  AOI22_X1 U21789 ( .A1(n18662), .A2(n18661), .B1(n18660), .B2(n18659), .ZN(
        n18667) );
  AOI22_X1 U21790 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18665), .B1(
        n18664), .B2(n18663), .ZN(n18666) );
  OAI211_X1 U21791 ( .C1(n18669), .C2(n18668), .A(n18667), .B(n18666), .ZN(
        P3_U2995) );
  NAND2_X1 U21792 ( .A1(n18671), .A2(n18670), .ZN(n18672) );
  AOI22_X1 U21793 ( .A1(n18675), .A2(n18674), .B1(n18673), .B2(n18672), .ZN(
        n18676) );
  OAI221_X1 U21794 ( .B1(n18678), .B2(n18709), .C1(n18678), .C2(n18677), .A(
        n18676), .ZN(n18880) );
  OAI21_X1 U21795 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18679), .ZN(n18680) );
  OAI211_X1 U21796 ( .C1(n18710), .C2(n18682), .A(n18681), .B(n18680), .ZN(
        n18721) );
  NAND2_X1 U21797 ( .A1(n18851), .A2(n18704), .ZN(n18689) );
  AOI21_X1 U21798 ( .B1(n18694), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n18683), .ZN(n18697) );
  INV_X1 U21799 ( .A(n18697), .ZN(n18705) );
  AOI22_X1 U21800 ( .A1(n18684), .A2(n18689), .B1(n18690), .B2(n18705), .ZN(
        n18685) );
  NOR2_X1 U21801 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18685), .ZN(
        n18838) );
  OAI21_X1 U21802 ( .B1(n18688), .B2(n18687), .A(n18686), .ZN(n18703) );
  OAI21_X1 U21803 ( .B1(n18696), .B2(n18690), .A(n18689), .ZN(n18691) );
  AOI21_X1 U21804 ( .B1(n18703), .B2(n18692), .A(n18691), .ZN(n18839) );
  NAND2_X1 U21805 ( .A1(n18710), .A2(n18839), .ZN(n18693) );
  AOI22_X1 U21806 ( .A1(n18710), .A2(n18838), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18693), .ZN(n18719) );
  NOR2_X1 U21807 ( .A1(n18695), .A2(n18694), .ZN(n18698) );
  AOI22_X1 U21808 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18696), .B1(
        n18698), .B2(n18869), .ZN(n18864) );
  NOR2_X1 U21809 ( .A1(n18864), .A2(n18699), .ZN(n18702) );
  OAI22_X1 U21810 ( .A1(n18698), .A2(n18853), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18697), .ZN(n18857) );
  OAI221_X1 U21811 ( .B1(n18857), .B2(n18864), .C1(n18857), .C2(n18699), .A(
        n18710), .ZN(n18700) );
  AOI22_X1 U21812 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18702), .B1(
        n18701), .B2(n18700), .ZN(n18713) );
  NAND3_X1 U21813 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18704), .A3(
        n18703), .ZN(n18708) );
  OAI211_X1 U21814 ( .C1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n18706), .B(n18705), .ZN(
        n18707) );
  OAI211_X1 U21815 ( .C1(n18848), .C2(n18709), .A(n18708), .B(n18707), .ZN(
        n18849) );
  MUX2_X1 U21816 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n18849), .S(
        n18710), .Z(n18714) );
  AND2_X1 U21817 ( .A1(n18713), .A2(n18714), .ZN(n18711) );
  OAI221_X1 U21818 ( .B1(n18713), .B2(n18714), .C1(n18712), .C2(n18711), .A(
        n18716), .ZN(n18718) );
  AOI21_X1 U21819 ( .B1(n18716), .B2(n18715), .A(n18714), .ZN(n18717) );
  AOI222_X1 U21820 ( .A1(n18719), .A2(n18718), .B1(n18719), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18718), .C2(n18717), .ZN(
        n18720) );
  NOR4_X1 U21821 ( .A1(n18722), .A2(n18880), .A3(n18721), .A4(n18720), .ZN(
        n18733) );
  INV_X1 U21822 ( .A(n18854), .ZN(n18865) );
  NOR2_X1 U21823 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18892) );
  AOI22_X1 U21824 ( .A1(n18865), .A2(n18892), .B1(n18884), .B2(n17468), .ZN(
        n18723) );
  INV_X1 U21825 ( .A(n18723), .ZN(n18729) );
  OAI211_X1 U21826 ( .C1(n18725), .C2(n18724), .A(n18882), .B(n18733), .ZN(
        n18835) );
  NAND2_X1 U21827 ( .A1(n18884), .A2(n18726), .ZN(n18734) );
  NAND2_X1 U21828 ( .A1(n18835), .A2(n18734), .ZN(n18736) );
  NOR2_X1 U21829 ( .A1(n18727), .A2(n18736), .ZN(n18728) );
  MUX2_X1 U21830 ( .A(n18729), .B(n18728), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18731) );
  OAI211_X1 U21831 ( .C1(n18733), .C2(n18732), .A(n18731), .B(n18730), .ZN(
        P3_U2996) );
  NOR2_X1 U21832 ( .A1(n18890), .A2(n18883), .ZN(n18740) );
  NOR3_X1 U21833 ( .A1(n18847), .A2(n18735), .A3(n18734), .ZN(n18743) );
  NOR3_X1 U21834 ( .A1(n9814), .A2(n18737), .A3(n18736), .ZN(n18739) );
  OR4_X1 U21835 ( .A1(n18741), .A2(n18740), .A3(n18743), .A4(n18739), .ZN(
        P3_U2997) );
  NOR4_X1 U21836 ( .A1(n18892), .A2(n18744), .A3(n18743), .A4(n18742), .ZN(
        P3_U2998) );
  AND2_X1 U21837 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18830), .ZN(
        P3_U2999) );
  AND2_X1 U21838 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18830), .ZN(
        P3_U3000) );
  AND2_X1 U21839 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18830), .ZN(
        P3_U3001) );
  AND2_X1 U21840 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18830), .ZN(
        P3_U3002) );
  AND2_X1 U21841 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18830), .ZN(
        P3_U3003) );
  AND2_X1 U21842 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18830), .ZN(
        P3_U3004) );
  AND2_X1 U21843 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18830), .ZN(
        P3_U3005) );
  AND2_X1 U21844 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18830), .ZN(
        P3_U3006) );
  AND2_X1 U21845 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18830), .ZN(
        P3_U3007) );
  AND2_X1 U21846 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18830), .ZN(
        P3_U3008) );
  AND2_X1 U21847 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18830), .ZN(
        P3_U3009) );
  AND2_X1 U21848 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18830), .ZN(
        P3_U3010) );
  AND2_X1 U21849 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18830), .ZN(
        P3_U3011) );
  AND2_X1 U21850 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18830), .ZN(
        P3_U3012) );
  AND2_X1 U21851 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18830), .ZN(
        P3_U3013) );
  AND2_X1 U21852 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18830), .ZN(
        P3_U3014) );
  AND2_X1 U21853 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18830), .ZN(
        P3_U3015) );
  AND2_X1 U21854 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18830), .ZN(
        P3_U3016) );
  AND2_X1 U21855 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18830), .ZN(
        P3_U3017) );
  AND2_X1 U21856 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18830), .ZN(
        P3_U3018) );
  AND2_X1 U21857 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18830), .ZN(
        P3_U3019) );
  AND2_X1 U21858 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18830), .ZN(
        P3_U3020) );
  AND2_X1 U21859 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18830), .ZN(P3_U3021) );
  AND2_X1 U21860 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18830), .ZN(P3_U3022) );
  AND2_X1 U21861 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18830), .ZN(P3_U3023) );
  AND2_X1 U21862 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18830), .ZN(P3_U3024) );
  AND2_X1 U21863 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18830), .ZN(P3_U3025) );
  AND2_X1 U21864 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18830), .ZN(P3_U3026) );
  AND2_X1 U21865 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18830), .ZN(P3_U3027) );
  AND2_X1 U21866 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18830), .ZN(P3_U3028) );
  NAND2_X1 U21867 ( .A1(n18884), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18754) );
  OAI21_X1 U21868 ( .B1(n18745), .B2(n21232), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18747) );
  INV_X1 U21869 ( .A(NA), .ZN(n21180) );
  NOR3_X1 U21870 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .A3(n21180), .ZN(n18746) );
  AOI21_X1 U21871 ( .B1(n18898), .B2(n18747), .A(n18746), .ZN(n18748) );
  OAI221_X1 U21872 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(P3_STATE_REG_0__SCAN_IN), .C1(P3_STATE_REG_2__SCAN_IN), .C2(n18754), .A(n18748), .ZN(P3_U3029) );
  AOI21_X1 U21873 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(HOLD), .A(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18749) );
  AOI21_X1 U21874 ( .B1(HOLD), .B2(P3_STATE_REG_2__SCAN_IN), .A(n18749), .ZN(
        n18750) );
  AOI22_X1 U21875 ( .A1(n18884), .A2(P3_STATE_REG_1__SCAN_IN), .B1(
        P3_STATE_REG_0__SCAN_IN), .B2(n18750), .ZN(n18752) );
  INV_X1 U21876 ( .A(n18751), .ZN(n18887) );
  NAND2_X1 U21877 ( .A1(n18752), .A2(n18887), .ZN(P3_U3030) );
  INV_X1 U21878 ( .A(n18754), .ZN(n18753) );
  AOI221_X1 U21879 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n18758), .C1(n21180), 
        .C2(n18758), .A(n18753), .ZN(n18759) );
  NOR2_X1 U21880 ( .A1(n18761), .A2(n21232), .ZN(n18756) );
  OAI22_X1 U21881 ( .A1(NA), .A2(n18754), .B1(P3_STATE_REG_1__SCAN_IN), .B2(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18755) );
  OAI22_X1 U21882 ( .A1(n18756), .A2(n18755), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18757) );
  OAI22_X1 U21883 ( .A1(n18759), .A2(n18761), .B1(n18758), .B2(n18757), .ZN(
        P3_U3031) );
  OAI222_X1 U21884 ( .A1(n18870), .A2(n18823), .B1(n18762), .B2(n18897), .C1(
        n18763), .C2(n18815), .ZN(P3_U3032) );
  OAI222_X1 U21885 ( .A1(n18815), .A2(n18765), .B1(n18764), .B2(n18897), .C1(
        n18763), .C2(n18823), .ZN(P3_U3033) );
  OAI222_X1 U21886 ( .A1(n18815), .A2(n18767), .B1(n18766), .B2(n18897), .C1(
        n18765), .C2(n18823), .ZN(P3_U3034) );
  INV_X1 U21887 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18769) );
  OAI222_X1 U21888 ( .A1(n18815), .A2(n18769), .B1(n18768), .B2(n18897), .C1(
        n18767), .C2(n18823), .ZN(P3_U3035) );
  OAI222_X1 U21889 ( .A1(n18815), .A2(n18771), .B1(n18770), .B2(n18897), .C1(
        n18769), .C2(n18823), .ZN(P3_U3036) );
  OAI222_X1 U21890 ( .A1(n18815), .A2(n18773), .B1(n18772), .B2(n18897), .C1(
        n18771), .C2(n18823), .ZN(P3_U3037) );
  OAI222_X1 U21891 ( .A1(n18815), .A2(n18776), .B1(n18774), .B2(n18897), .C1(
        n18773), .C2(n18823), .ZN(P3_U3038) );
  OAI222_X1 U21892 ( .A1(n18776), .A2(n18823), .B1(n18775), .B2(n18897), .C1(
        n18777), .C2(n18815), .ZN(P3_U3039) );
  OAI222_X1 U21893 ( .A1(n18815), .A2(n18779), .B1(n18778), .B2(n18897), .C1(
        n18777), .C2(n18823), .ZN(P3_U3040) );
  OAI222_X1 U21894 ( .A1(n18815), .A2(n18781), .B1(n18780), .B2(n18897), .C1(
        n18779), .C2(n18823), .ZN(P3_U3041) );
  OAI222_X1 U21895 ( .A1(n18815), .A2(n18783), .B1(n18782), .B2(n18897), .C1(
        n18781), .C2(n18823), .ZN(P3_U3042) );
  OAI222_X1 U21896 ( .A1(n18815), .A2(n18785), .B1(n18784), .B2(n18897), .C1(
        n18783), .C2(n18823), .ZN(P3_U3043) );
  OAI222_X1 U21897 ( .A1(n18815), .A2(n18788), .B1(n18786), .B2(n18897), .C1(
        n18785), .C2(n18823), .ZN(P3_U3044) );
  OAI222_X1 U21898 ( .A1(n18788), .A2(n18823), .B1(n18787), .B2(n18897), .C1(
        n18790), .C2(n18815), .ZN(P3_U3045) );
  OAI222_X1 U21899 ( .A1(n18790), .A2(n18823), .B1(n18789), .B2(n18897), .C1(
        n18791), .C2(n18815), .ZN(P3_U3046) );
  OAI222_X1 U21900 ( .A1(n18815), .A2(n18793), .B1(n18792), .B2(n18897), .C1(
        n18791), .C2(n18823), .ZN(P3_U3047) );
  OAI222_X1 U21901 ( .A1(n18815), .A2(n18795), .B1(n18794), .B2(n18897), .C1(
        n18793), .C2(n18823), .ZN(P3_U3048) );
  OAI222_X1 U21902 ( .A1(n18815), .A2(n18797), .B1(n18796), .B2(n18897), .C1(
        n18795), .C2(n18823), .ZN(P3_U3049) );
  OAI222_X1 U21903 ( .A1(n18815), .A2(n18800), .B1(n18798), .B2(n18897), .C1(
        n18797), .C2(n18823), .ZN(P3_U3050) );
  OAI222_X1 U21904 ( .A1(n18800), .A2(n18823), .B1(n18799), .B2(n18897), .C1(
        n18801), .C2(n18815), .ZN(P3_U3051) );
  OAI222_X1 U21905 ( .A1(n18815), .A2(n18803), .B1(n18802), .B2(n18897), .C1(
        n18801), .C2(n18823), .ZN(P3_U3052) );
  OAI222_X1 U21906 ( .A1(n18815), .A2(n18806), .B1(n18804), .B2(n18897), .C1(
        n18803), .C2(n18823), .ZN(P3_U3053) );
  OAI222_X1 U21907 ( .A1(n18806), .A2(n18823), .B1(n18805), .B2(n18897), .C1(
        n18807), .C2(n18815), .ZN(P3_U3054) );
  OAI222_X1 U21908 ( .A1(n18815), .A2(n18809), .B1(n18808), .B2(n18897), .C1(
        n18807), .C2(n18823), .ZN(P3_U3055) );
  INV_X1 U21909 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18811) );
  OAI222_X1 U21910 ( .A1(n18815), .A2(n18811), .B1(n18810), .B2(n18897), .C1(
        n18809), .C2(n18823), .ZN(P3_U3056) );
  OAI222_X1 U21911 ( .A1(n18815), .A2(n18813), .B1(n18812), .B2(n18897), .C1(
        n18811), .C2(n18823), .ZN(P3_U3057) );
  OAI222_X1 U21912 ( .A1(n18815), .A2(n18817), .B1(n18814), .B2(n18897), .C1(
        n18813), .C2(n18823), .ZN(P3_U3058) );
  OAI222_X1 U21913 ( .A1(n18817), .A2(n18823), .B1(n18816), .B2(n18897), .C1(
        n18818), .C2(n18815), .ZN(P3_U3059) );
  OAI222_X1 U21914 ( .A1(n18815), .A2(n18822), .B1(n18819), .B2(n18897), .C1(
        n18818), .C2(n18823), .ZN(P3_U3060) );
  INV_X1 U21915 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18821) );
  OAI222_X1 U21916 ( .A1(n18823), .A2(n18822), .B1(n18821), .B2(n18897), .C1(
        n18820), .C2(n18815), .ZN(P3_U3061) );
  OAI22_X1 U21917 ( .A1(n18898), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18897), .ZN(n18824) );
  INV_X1 U21918 ( .A(n18824), .ZN(P3_U3274) );
  OAI22_X1 U21919 ( .A1(n18898), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18897), .ZN(n18825) );
  INV_X1 U21920 ( .A(n18825), .ZN(P3_U3275) );
  OAI22_X1 U21921 ( .A1(n18898), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18897), .ZN(n18826) );
  INV_X1 U21922 ( .A(n18826), .ZN(P3_U3276) );
  OAI22_X1 U21923 ( .A1(n18898), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18897), .ZN(n18827) );
  INV_X1 U21924 ( .A(n18827), .ZN(P3_U3277) );
  INV_X1 U21925 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18829) );
  INV_X1 U21926 ( .A(n18831), .ZN(n18828) );
  AOI21_X1 U21927 ( .B1(n18830), .B2(n18829), .A(n18828), .ZN(P3_U3280) );
  OAI21_X1 U21928 ( .B1(n18833), .B2(n18832), .A(n18831), .ZN(P3_U3281) );
  OAI221_X1 U21929 ( .B1(n18863), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18863), 
        .C2(n18835), .A(n18834), .ZN(P3_U3282) );
  INV_X1 U21930 ( .A(n18900), .ZN(n18858) );
  INV_X1 U21931 ( .A(n18836), .ZN(n18837) );
  AOI22_X1 U21932 ( .A1(n18858), .A2(n18838), .B1(n18865), .B2(n18837), .ZN(
        n18843) );
  INV_X1 U21933 ( .A(n18868), .ZN(n18859) );
  OAI21_X1 U21934 ( .B1(n18900), .B2(n18839), .A(n18859), .ZN(n18840) );
  INV_X1 U21935 ( .A(n18840), .ZN(n18842) );
  OAI22_X1 U21936 ( .A1(n18868), .A2(n18843), .B1(n18842), .B2(n18841), .ZN(
        P3_U3285) );
  AOI22_X1 U21937 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n18845), .B2(n18844), .ZN(
        n18855) );
  NOR2_X1 U21938 ( .A1(n18847), .A2(n18846), .ZN(n18852) );
  AOI222_X1 U21939 ( .A1(n18849), .A2(n18858), .B1(n18855), .B2(n18852), .C1(
        n18865), .C2(n18848), .ZN(n18850) );
  AOI22_X1 U21940 ( .A1(n18868), .A2(n18851), .B1(n18850), .B2(n18859), .ZN(
        P3_U3288) );
  INV_X1 U21941 ( .A(n18852), .ZN(n18862) );
  OAI22_X1 U21942 ( .A1(n18855), .A2(n18862), .B1(n18854), .B2(n18853), .ZN(
        n18856) );
  AOI21_X1 U21943 ( .B1(n18858), .B2(n18857), .A(n18856), .ZN(n18860) );
  AOI22_X1 U21944 ( .A1(n18868), .A2(n18861), .B1(n18860), .B2(n18859), .ZN(
        P3_U3289) );
  OAI221_X1 U21945 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(n18864), .C1(
        P3_STATE2_REG_1__SCAN_IN), .C2(n18863), .A(n18862), .ZN(n18867) );
  AOI21_X1 U21946 ( .B1(n18869), .B2(n18865), .A(n18868), .ZN(n18866) );
  AOI22_X1 U21947 ( .A1(n18869), .A2(n18868), .B1(n18867), .B2(n18866), .ZN(
        P3_U3290) );
  AOI21_X1 U21948 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18871) );
  AOI22_X1 U21949 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18871), .B2(n18870), .ZN(n18874) );
  INV_X1 U21950 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18873) );
  AOI22_X1 U21951 ( .A1(n18877), .A2(n18874), .B1(n18873), .B2(n18872), .ZN(
        P3_U3292) );
  INV_X1 U21952 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18876) );
  OAI21_X1 U21953 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18877), .ZN(n18875) );
  OAI21_X1 U21954 ( .B1(n18877), .B2(n18876), .A(n18875), .ZN(P3_U3293) );
  INV_X1 U21955 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18878) );
  AOI22_X1 U21956 ( .A1(n18897), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18878), 
        .B2(n18898), .ZN(P3_U3294) );
  MUX2_X1 U21957 ( .A(P3_MORE_REG_SCAN_IN), .B(n18880), .S(n18879), .Z(
        P3_U3295) );
  OAI22_X1 U21958 ( .A1(n18884), .A2(n18883), .B1(n18882), .B2(n18881), .ZN(
        n18885) );
  NOR2_X1 U21959 ( .A1(n18886), .A2(n18885), .ZN(n18896) );
  AOI21_X1 U21960 ( .B1(n18889), .B2(n18888), .A(n18887), .ZN(n18891) );
  OAI211_X1 U21961 ( .C1(n18891), .C2(n18902), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18890), .ZN(n18893) );
  AOI21_X1 U21962 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18893), .A(n18892), 
        .ZN(n18895) );
  NAND2_X1 U21963 ( .A1(n18896), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18894) );
  OAI21_X1 U21964 ( .B1(n18896), .B2(n18895), .A(n18894), .ZN(P3_U3296) );
  OAI22_X1 U21965 ( .A1(n18898), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18897), .ZN(n18899) );
  INV_X1 U21966 ( .A(n18899), .ZN(P3_U3297) );
  OAI21_X1 U21967 ( .B1(n18900), .B2(P3_STATE2_REG_2__SCAN_IN), .A(n18901), 
        .ZN(n18905) );
  OAI22_X1 U21968 ( .A1(n18902), .A2(n18901), .B1(n18905), .B2(
        P3_READREQUEST_REG_SCAN_IN), .ZN(n18903) );
  INV_X1 U21969 ( .A(n18903), .ZN(P3_U3298) );
  OAI21_X1 U21970 ( .B1(n18905), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n18904), 
        .ZN(n18906) );
  INV_X1 U21971 ( .A(n18906), .ZN(P3_U3299) );
  NAND2_X1 U21972 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19856), .ZN(n19843) );
  AOI22_X1 U21973 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19843), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n19837), .ZN(n19921) );
  AOI21_X1 U21974 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19921), .ZN(n18907) );
  INV_X1 U21975 ( .A(n18907), .ZN(P2_U2815) );
  INV_X1 U21976 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18910) );
  OAI22_X1 U21977 ( .A1(n18911), .A2(n18910), .B1(n18909), .B2(n18908), .ZN(
        P2_U2816) );
  NOR2_X2 U21978 ( .A1(n19848), .A2(P2_STATE_REG_0__SCAN_IN), .ZN(n19912) );
  AOI21_X1 U21979 ( .B1(n19837), .B2(n19856), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18912) );
  AOI22_X1 U21980 ( .A1(n19868), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n18912), 
        .B2(n19978), .ZN(P2_U2817) );
  INV_X1 U21981 ( .A(n19836), .ZN(n19846) );
  OAI21_X1 U21982 ( .B1(n19846), .B2(BS16), .A(n19921), .ZN(n19919) );
  OAI21_X1 U21983 ( .B1(n19921), .B2(n19924), .A(n19919), .ZN(P2_U2818) );
  NOR4_X1 U21984 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18916) );
  NOR4_X1 U21985 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n18915) );
  NOR4_X1 U21986 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18914) );
  NOR4_X1 U21987 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18913) );
  NAND4_X1 U21988 ( .A1(n18916), .A2(n18915), .A3(n18914), .A4(n18913), .ZN(
        n18922) );
  NOR4_X1 U21989 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n18920) );
  AOI211_X1 U21990 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n18919) );
  NOR4_X1 U21991 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n18918) );
  NOR4_X1 U21992 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n18917) );
  NAND4_X1 U21993 ( .A1(n18920), .A2(n18919), .A3(n18918), .A4(n18917), .ZN(
        n18921) );
  NOR2_X1 U21994 ( .A1(n18922), .A2(n18921), .ZN(n18933) );
  INV_X1 U21995 ( .A(n18933), .ZN(n18931) );
  NOR2_X1 U21996 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18931), .ZN(n18925) );
  INV_X1 U21997 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18923) );
  AOI22_X1 U21998 ( .A1(n18925), .A2(n18926), .B1(n18931), .B2(n18923), .ZN(
        P2_U2820) );
  OR3_X1 U21999 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18930) );
  INV_X1 U22000 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18924) );
  AOI22_X1 U22001 ( .A1(n18925), .A2(n18930), .B1(n18931), .B2(n18924), .ZN(
        P2_U2821) );
  INV_X1 U22002 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19920) );
  NAND2_X1 U22003 ( .A1(n18925), .A2(n19920), .ZN(n18929) );
  OAI21_X1 U22004 ( .B1(n18926), .B2(n19857), .A(n18933), .ZN(n18927) );
  OAI21_X1 U22005 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18933), .A(n18927), 
        .ZN(n18928) );
  OAI221_X1 U22006 ( .B1(n18929), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18929), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18928), .ZN(P2_U2822) );
  INV_X1 U22007 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18932) );
  OAI221_X1 U22008 ( .B1(n18933), .B2(n18932), .C1(n18931), .C2(n18930), .A(
        n18929), .ZN(P2_U2823) );
  AOI22_X1 U22009 ( .A1(n18935), .A2(n19081), .B1(n18938), .B2(n18934), .ZN(
        n18947) );
  AOI22_X1 U22010 ( .A1(P2_REIP_REG_20__SCAN_IN), .A2(n19080), .B1(
        P2_EBX_REG_20__SCAN_IN), .B2(n19109), .ZN(n18946) );
  AOI21_X1 U22011 ( .B1(n18938), .B2(n18937), .A(n18936), .ZN(n18939) );
  AOI22_X1 U22012 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19089), .B1(
        n18940), .B2(n18939), .ZN(n18945) );
  INV_X1 U22013 ( .A(n18941), .ZN(n18943) );
  AOI22_X1 U22014 ( .A1(n18943), .A2(n11089), .B1(n19036), .B2(n18942), .ZN(
        n18944) );
  NAND4_X1 U22015 ( .A1(n18947), .A2(n18946), .A3(n18945), .A4(n18944), .ZN(
        P2_U2835) );
  OAI22_X1 U22016 ( .A1(n18948), .A2(n19106), .B1(n19891), .B2(n19122), .ZN(
        n18949) );
  AOI211_X1 U22017 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n19109), .A(n19223), .B(
        n18949), .ZN(n18958) );
  NOR2_X1 U22018 ( .A1(n10145), .A2(n18950), .ZN(n18951) );
  XOR2_X1 U22019 ( .A(n18952), .B(n18951), .Z(n18956) );
  OAI22_X1 U22020 ( .A1(n18954), .A2(n19115), .B1(n18953), .B2(n19116), .ZN(
        n18955) );
  AOI21_X1 U22021 ( .B1(n18956), .B2(n19118), .A(n18955), .ZN(n18957) );
  OAI211_X1 U22022 ( .C1(n18959), .C2(n19105), .A(n18958), .B(n18957), .ZN(
        P2_U2836) );
  NAND2_X1 U22023 ( .A1(n13535), .A2(n18960), .ZN(n18961) );
  XOR2_X1 U22024 ( .A(n18962), .B(n18961), .Z(n18970) );
  OAI21_X1 U22025 ( .B1(n11040), .B2(n19085), .A(n19040), .ZN(n18965) );
  OAI22_X1 U22026 ( .A1(n18963), .A2(n19106), .B1(n19889), .B2(n19122), .ZN(
        n18964) );
  AOI211_X1 U22027 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n19089), .A(
        n18965), .B(n18964), .ZN(n18969) );
  AOI22_X1 U22028 ( .A1(n18967), .A2(n19036), .B1(n18966), .B2(n11089), .ZN(
        n18968) );
  OAI211_X1 U22029 ( .C1(n19831), .C2(n18970), .A(n18969), .B(n18968), .ZN(
        P2_U2837) );
  OAI22_X1 U22030 ( .A1(n18971), .A2(n19106), .B1(n19887), .B2(n19122), .ZN(
        n18972) );
  AOI211_X1 U22031 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n19109), .A(n19223), .B(
        n18972), .ZN(n18981) );
  NOR2_X1 U22032 ( .A1(n10145), .A2(n18973), .ZN(n18974) );
  XNOR2_X1 U22033 ( .A(n18975), .B(n18974), .ZN(n18979) );
  OAI22_X1 U22034 ( .A1(n18977), .A2(n19116), .B1(n19115), .B2(n18976), .ZN(
        n18978) );
  AOI21_X1 U22035 ( .B1(n18979), .B2(n19118), .A(n18978), .ZN(n18980) );
  OAI211_X1 U22036 ( .C1(n18982), .C2(n19105), .A(n18981), .B(n18980), .ZN(
        P2_U2838) );
  NAND2_X1 U22037 ( .A1(n13535), .A2(n18983), .ZN(n18984) );
  XOR2_X1 U22038 ( .A(n18985), .B(n18984), .Z(n18994) );
  OAI21_X1 U22039 ( .B1(n10888), .B2(n19085), .A(n19040), .ZN(n18989) );
  INV_X1 U22040 ( .A(n18986), .ZN(n18987) );
  OAI22_X1 U22041 ( .A1(n18987), .A2(n19106), .B1(n19885), .B2(n19122), .ZN(
        n18988) );
  AOI211_X1 U22042 ( .C1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n19089), .A(
        n18989), .B(n18988), .ZN(n18993) );
  OAI22_X1 U22043 ( .A1(n19132), .A2(n19116), .B1(n19115), .B2(n18990), .ZN(
        n18991) );
  INV_X1 U22044 ( .A(n18991), .ZN(n18992) );
  OAI211_X1 U22045 ( .C1(n19831), .C2(n18994), .A(n18993), .B(n18992), .ZN(
        P2_U2839) );
  OAI22_X1 U22046 ( .A1(n18996), .A2(n19106), .B1(n19105), .B2(n18995), .ZN(
        n18997) );
  AOI211_X1 U22047 ( .C1(P2_EBX_REG_15__SCAN_IN), .C2(n19109), .A(n19223), .B(
        n18997), .ZN(n19005) );
  NOR2_X1 U22048 ( .A1(n10145), .A2(n18998), .ZN(n18999) );
  XOR2_X1 U22049 ( .A(n19000), .B(n18999), .Z(n19003) );
  OAI22_X1 U22050 ( .A1(n19139), .A2(n19116), .B1(n19115), .B2(n19001), .ZN(
        n19002) );
  AOI21_X1 U22051 ( .B1(n19003), .B2(n19118), .A(n19002), .ZN(n19004) );
  OAI211_X1 U22052 ( .C1(n19883), .C2(n19122), .A(n19005), .B(n19004), .ZN(
        P2_U2840) );
  NAND2_X1 U22053 ( .A1(n13535), .A2(n19006), .ZN(n19007) );
  XOR2_X1 U22054 ( .A(n19008), .B(n19007), .Z(n19016) );
  AOI22_X1 U22055 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n19080), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19089), .ZN(n19009) );
  OAI21_X1 U22056 ( .B1(n19010), .B2(n19106), .A(n19009), .ZN(n19011) );
  AOI211_X1 U22057 ( .C1(P2_EBX_REG_14__SCAN_IN), .C2(n19109), .A(n19223), .B(
        n19011), .ZN(n19015) );
  AOI22_X1 U22058 ( .A1(n19013), .A2(n19036), .B1(n11089), .B2(n19012), .ZN(
        n19014) );
  OAI211_X1 U22059 ( .C1(n19831), .C2(n19016), .A(n19015), .B(n19014), .ZN(
        P2_U2841) );
  OAI21_X1 U22060 ( .B1(n11022), .B2(n19085), .A(n19040), .ZN(n19020) );
  OAI22_X1 U22061 ( .A1(n19018), .A2(n19106), .B1(n19105), .B2(n19017), .ZN(
        n19019) );
  AOI211_X1 U22062 ( .C1(P2_REIP_REG_13__SCAN_IN), .C2(n19080), .A(n19020), 
        .B(n19019), .ZN(n19028) );
  NOR2_X1 U22063 ( .A1(n10145), .A2(n19021), .ZN(n19023) );
  XOR2_X1 U22064 ( .A(n19023), .B(n19022), .Z(n19026) );
  INV_X1 U22065 ( .A(n19024), .ZN(n19025) );
  AOI22_X1 U22066 ( .A1(n19026), .A2(n19118), .B1(n11089), .B2(n19025), .ZN(
        n19027) );
  OAI211_X1 U22067 ( .C1(n19143), .C2(n19116), .A(n19028), .B(n19027), .ZN(
        P2_U2842) );
  NAND2_X1 U22068 ( .A1(n13535), .A2(n19029), .ZN(n19030) );
  XOR2_X1 U22069 ( .A(n19031), .B(n19030), .Z(n19039) );
  AOI22_X1 U22070 ( .A1(n19032), .A2(n19081), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19089), .ZN(n19033) );
  OAI211_X1 U22071 ( .C1(n11019), .C2(n19085), .A(n19033), .B(n19083), .ZN(
        n19034) );
  AOI21_X1 U22072 ( .B1(P2_REIP_REG_12__SCAN_IN), .B2(n19080), .A(n19034), 
        .ZN(n19038) );
  AOI22_X1 U22073 ( .A1(n19144), .A2(n19036), .B1(n11089), .B2(n19035), .ZN(
        n19037) );
  OAI211_X1 U22074 ( .C1(n19831), .C2(n19039), .A(n19038), .B(n19037), .ZN(
        P2_U2843) );
  OAI21_X1 U22075 ( .B1(n19041), .B2(n19085), .A(n19040), .ZN(n19045) );
  OAI22_X1 U22076 ( .A1(n19043), .A2(n19106), .B1(n19105), .B2(n19042), .ZN(
        n19044) );
  AOI211_X1 U22077 ( .C1(P2_REIP_REG_11__SCAN_IN), .C2(n19080), .A(n19045), 
        .B(n19044), .ZN(n19053) );
  NOR2_X1 U22078 ( .A1(n10145), .A2(n19046), .ZN(n19048) );
  XOR2_X1 U22079 ( .A(n19048), .B(n19047), .Z(n19051) );
  INV_X1 U22080 ( .A(n19049), .ZN(n19050) );
  AOI22_X1 U22081 ( .A1(n19051), .A2(n19118), .B1(n11089), .B2(n19050), .ZN(
        n19052) );
  OAI211_X1 U22082 ( .C1(n19149), .C2(n19116), .A(n19053), .B(n19052), .ZN(
        P2_U2844) );
  AOI22_X1 U22083 ( .A1(n19054), .A2(n19081), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19089), .ZN(n19055) );
  OAI211_X1 U22084 ( .C1(n19056), .C2(n19085), .A(n19055), .B(n19083), .ZN(
        n19057) );
  AOI21_X1 U22085 ( .B1(P2_REIP_REG_10__SCAN_IN), .B2(n19080), .A(n19057), 
        .ZN(n19064) );
  NAND2_X1 U22086 ( .A1(n13535), .A2(n19058), .ZN(n19059) );
  XOR2_X1 U22087 ( .A(n19060), .B(n19059), .Z(n19062) );
  AOI22_X1 U22088 ( .A1(n19062), .A2(n19118), .B1(n11089), .B2(n19061), .ZN(
        n19063) );
  OAI211_X1 U22089 ( .C1(n19152), .C2(n19116), .A(n19064), .B(n19063), .ZN(
        P2_U2845) );
  NAND2_X1 U22090 ( .A1(n13535), .A2(n19065), .ZN(n19066) );
  XOR2_X1 U22091 ( .A(n19067), .B(n19066), .Z(n19076) );
  AOI22_X1 U22092 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19080), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19089), .ZN(n19068) );
  OAI21_X1 U22093 ( .B1(n19069), .B2(n19106), .A(n19068), .ZN(n19070) );
  AOI211_X1 U22094 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n19109), .A(n19223), .B(
        n19070), .ZN(n19075) );
  INV_X1 U22095 ( .A(n19071), .ZN(n19156) );
  OAI22_X1 U22096 ( .A1(n19072), .A2(n19115), .B1(n19116), .B2(n19156), .ZN(
        n19073) );
  INV_X1 U22097 ( .A(n19073), .ZN(n19074) );
  OAI211_X1 U22098 ( .C1(n19831), .C2(n19076), .A(n19075), .B(n19074), .ZN(
        P2_U2847) );
  NOR2_X1 U22099 ( .A1(n10145), .A2(n19077), .ZN(n19078) );
  XOR2_X1 U22100 ( .A(n19079), .B(n19078), .Z(n19091) );
  AOI22_X1 U22101 ( .A1(n19082), .A2(n19081), .B1(P2_REIP_REG_7__SCAN_IN), 
        .B2(n19080), .ZN(n19084) );
  OAI211_X1 U22102 ( .C1(n10997), .C2(n19085), .A(n19084), .B(n19083), .ZN(
        n19088) );
  OAI22_X1 U22103 ( .A1(n19158), .A2(n19116), .B1(n19115), .B2(n19086), .ZN(
        n19087) );
  AOI211_X1 U22104 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19089), .A(
        n19088), .B(n19087), .ZN(n19090) );
  OAI21_X1 U22105 ( .B1(n19831), .B2(n19091), .A(n19090), .ZN(P2_U2848) );
  AOI21_X1 U22106 ( .B1(P2_EBX_REG_6__SCAN_IN), .B2(n19109), .A(n19223), .ZN(
        n19095) );
  OAI22_X1 U22107 ( .A1(n19092), .A2(n19106), .B1(n19105), .B2(n16295), .ZN(
        n19093) );
  INV_X1 U22108 ( .A(n19093), .ZN(n19094) );
  OAI211_X1 U22109 ( .C1(n19865), .C2(n19122), .A(n19095), .B(n19094), .ZN(
        n19096) );
  INV_X1 U22110 ( .A(n19096), .ZN(n19103) );
  NAND2_X1 U22111 ( .A1(n13535), .A2(n19097), .ZN(n19098) );
  XNOR2_X1 U22112 ( .A(n19099), .B(n19098), .ZN(n19101) );
  AOI22_X1 U22113 ( .A1(n19101), .A2(n19118), .B1(n11089), .B2(n19100), .ZN(
        n19102) );
  OAI211_X1 U22114 ( .C1(n19116), .C2(n19161), .A(n19103), .B(n19102), .ZN(
        P2_U2849) );
  OAI22_X1 U22115 ( .A1(n19107), .A2(n19106), .B1(n19105), .B2(n19104), .ZN(
        n19108) );
  AOI211_X1 U22116 ( .C1(P2_EBX_REG_5__SCAN_IN), .C2(n19109), .A(n19223), .B(
        n19108), .ZN(n19121) );
  NOR2_X1 U22117 ( .A1(n10145), .A2(n19110), .ZN(n19112) );
  XNOR2_X1 U22118 ( .A(n19113), .B(n19112), .ZN(n19119) );
  OAI22_X1 U22119 ( .A1(n19168), .A2(n19116), .B1(n19115), .B2(n19114), .ZN(
        n19117) );
  AOI21_X1 U22120 ( .B1(n19119), .B2(n19118), .A(n19117), .ZN(n19120) );
  OAI211_X1 U22121 ( .C1(n13404), .C2(n19122), .A(n19121), .B(n19120), .ZN(
        P2_U2850) );
  AOI22_X1 U22122 ( .A1(n19123), .A2(n19177), .B1(n19129), .B2(
        BUF1_REG_31__SCAN_IN), .ZN(n19125) );
  AOI22_X1 U22123 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19176), .B1(n19128), 
        .B2(BUF2_REG_31__SCAN_IN), .ZN(n19124) );
  NAND2_X1 U22124 ( .A1(n19125), .A2(n19124), .ZN(P2_U2888) );
  INV_X1 U22125 ( .A(n19239), .ZN(n19126) );
  AOI22_X1 U22126 ( .A1(n19127), .A2(n19126), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n19176), .ZN(n19136) );
  AOI22_X1 U22127 ( .A1(n19129), .A2(BUF1_REG_16__SCAN_IN), .B1(n19128), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n19135) );
  OAI22_X1 U22128 ( .A1(n19132), .A2(n19131), .B1(n19181), .B2(n19130), .ZN(
        n19133) );
  INV_X1 U22129 ( .A(n19133), .ZN(n19134) );
  NAND3_X1 U22130 ( .A1(n19136), .A2(n19135), .A3(n19134), .ZN(P2_U2903) );
  OAI222_X1 U22131 ( .A1(n19139), .A2(n19169), .B1(n12509), .B2(n19160), .C1(
        n19138), .C2(n19185), .ZN(P2_U2904) );
  INV_X1 U22132 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19189) );
  OAI222_X1 U22133 ( .A1(n19141), .A2(n19169), .B1(n19189), .B2(n19160), .C1(
        n19185), .C2(n19140), .ZN(P2_U2905) );
  INV_X1 U22134 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19191) );
  OAI222_X1 U22135 ( .A1(n19143), .A2(n19169), .B1(n19191), .B2(n19160), .C1(
        n19185), .C2(n19142), .ZN(P2_U2906) );
  INV_X1 U22136 ( .A(n19144), .ZN(n19147) );
  AOI22_X1 U22137 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19176), .B1(n19145), 
        .B2(n19162), .ZN(n19146) );
  OAI21_X1 U22138 ( .B1(n19169), .B2(n19147), .A(n19146), .ZN(P2_U2907) );
  INV_X1 U22139 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19195) );
  OAI222_X1 U22140 ( .A1(n19149), .A2(n19169), .B1(n19195), .B2(n19160), .C1(
        n19185), .C2(n19148), .ZN(P2_U2908) );
  AOI22_X1 U22141 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19176), .B1(n19150), 
        .B2(n19162), .ZN(n19151) );
  OAI21_X1 U22142 ( .B1(n19169), .B2(n19152), .A(n19151), .ZN(P2_U2909) );
  INV_X1 U22143 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19199) );
  OAI222_X1 U22144 ( .A1(n19154), .A2(n19169), .B1(n19199), .B2(n19160), .C1(
        n19185), .C2(n19153), .ZN(P2_U2910) );
  INV_X1 U22145 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19201) );
  OAI222_X1 U22146 ( .A1(n19156), .A2(n19169), .B1(n19201), .B2(n19160), .C1(
        n19185), .C2(n19155), .ZN(P2_U2911) );
  INV_X1 U22147 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19203) );
  OAI222_X1 U22148 ( .A1(n19158), .A2(n19169), .B1(n19203), .B2(n19160), .C1(
        n19185), .C2(n19157), .ZN(P2_U2912) );
  INV_X1 U22149 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19206) );
  OAI222_X1 U22150 ( .A1(n19161), .A2(n19169), .B1(n19206), .B2(n19160), .C1(
        n19185), .C2(n19159), .ZN(P2_U2913) );
  AOI22_X1 U22151 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19176), .B1(n19163), .B2(
        n19162), .ZN(n19167) );
  OR3_X1 U22152 ( .A1(n19165), .A2(n19164), .A3(n19181), .ZN(n19166) );
  OAI211_X1 U22153 ( .C1(n19169), .C2(n19168), .A(n19167), .B(n19166), .ZN(
        P2_U2914) );
  AOI22_X1 U22154 ( .A1(n19927), .A2(n19177), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19176), .ZN(n19175) );
  AOI21_X1 U22155 ( .B1(n19172), .B2(n19171), .A(n19170), .ZN(n19173) );
  OR2_X1 U22156 ( .A1(n19173), .A2(n19181), .ZN(n19174) );
  OAI211_X1 U22157 ( .C1(n19257), .C2(n19185), .A(n19175), .B(n19174), .ZN(
        P2_U2916) );
  AOI22_X1 U22158 ( .A1(n19177), .A2(n19953), .B1(n19176), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19184) );
  AOI21_X1 U22159 ( .B1(n19180), .B2(n19179), .A(n19178), .ZN(n19182) );
  OR2_X1 U22160 ( .A1(n19182), .A2(n19181), .ZN(n19183) );
  OAI211_X1 U22161 ( .C1(n19248), .C2(n19185), .A(n19184), .B(n19183), .ZN(
        P2_U2918) );
  AND2_X1 U22162 ( .A1(n19204), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  AOI22_X1 U22163 ( .A1(n19218), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19217), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19187) );
  OAI21_X1 U22164 ( .B1(n12509), .B2(n19220), .A(n19187), .ZN(P2_U2936) );
  AOI22_X1 U22165 ( .A1(n19218), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19217), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19188) );
  OAI21_X1 U22166 ( .B1(n19189), .B2(n19220), .A(n19188), .ZN(P2_U2937) );
  AOI22_X1 U22167 ( .A1(n19218), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19217), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19190) );
  OAI21_X1 U22168 ( .B1(n19191), .B2(n19220), .A(n19190), .ZN(P2_U2938) );
  AOI22_X1 U22169 ( .A1(n19218), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19217), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19192) );
  OAI21_X1 U22170 ( .B1(n19193), .B2(n19220), .A(n19192), .ZN(P2_U2939) );
  AOI22_X1 U22171 ( .A1(n19218), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19204), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19194) );
  OAI21_X1 U22172 ( .B1(n19195), .B2(n19220), .A(n19194), .ZN(P2_U2940) );
  AOI22_X1 U22173 ( .A1(n19218), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19204), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19196) );
  OAI21_X1 U22174 ( .B1(n19197), .B2(n19220), .A(n19196), .ZN(P2_U2941) );
  AOI22_X1 U22175 ( .A1(n19218), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19204), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19198) );
  OAI21_X1 U22176 ( .B1(n19199), .B2(n19220), .A(n19198), .ZN(P2_U2942) );
  AOI22_X1 U22177 ( .A1(n19218), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19204), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19200) );
  OAI21_X1 U22178 ( .B1(n19201), .B2(n19220), .A(n19200), .ZN(P2_U2943) );
  AOI22_X1 U22179 ( .A1(n19218), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19204), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19202) );
  OAI21_X1 U22180 ( .B1(n19203), .B2(n19220), .A(n19202), .ZN(P2_U2944) );
  AOI22_X1 U22181 ( .A1(n19218), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19204), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19205) );
  OAI21_X1 U22182 ( .B1(n19206), .B2(n19220), .A(n19205), .ZN(P2_U2945) );
  INV_X1 U22183 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19208) );
  AOI22_X1 U22184 ( .A1(n19218), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19217), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19207) );
  OAI21_X1 U22185 ( .B1(n19208), .B2(n19220), .A(n19207), .ZN(P2_U2946) );
  INV_X1 U22186 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19210) );
  AOI22_X1 U22187 ( .A1(n19218), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19217), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19209) );
  OAI21_X1 U22188 ( .B1(n19210), .B2(n19220), .A(n19209), .ZN(P2_U2947) );
  INV_X1 U22189 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19212) );
  AOI22_X1 U22190 ( .A1(n19218), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19217), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19211) );
  OAI21_X1 U22191 ( .B1(n19212), .B2(n19220), .A(n19211), .ZN(P2_U2948) );
  INV_X1 U22192 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19214) );
  AOI22_X1 U22193 ( .A1(n19218), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19217), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19213) );
  OAI21_X1 U22194 ( .B1(n19214), .B2(n19220), .A(n19213), .ZN(P2_U2949) );
  INV_X1 U22195 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19216) );
  AOI22_X1 U22196 ( .A1(n19218), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19217), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19215) );
  OAI21_X1 U22197 ( .B1(n19216), .B2(n19220), .A(n19215), .ZN(P2_U2950) );
  AOI22_X1 U22198 ( .A1(n19218), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19217), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19219) );
  OAI21_X1 U22199 ( .B1(n12512), .B2(n19220), .A(n19219), .ZN(P2_U2951) );
  AOI22_X1 U22200 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19223), .B1(n19222), 
        .B2(n19221), .ZN(n19233) );
  INV_X1 U22201 ( .A(n19224), .ZN(n19228) );
  OAI22_X1 U22202 ( .A1(n19228), .A2(n19227), .B1(n19226), .B2(n19225), .ZN(
        n19229) );
  AOI21_X1 U22203 ( .B1(n19231), .B2(n19230), .A(n19229), .ZN(n19232) );
  OAI211_X1 U22204 ( .C1(n19235), .C2(n19234), .A(n19233), .B(n19232), .ZN(
        P2_U3010) );
  AOI22_X1 U22205 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19274), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19273), .ZN(n19764) );
  NAND2_X1 U22206 ( .A1(n19670), .A2(n19753), .ZN(n19800) );
  AOI22_X1 U22207 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19273), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n19274), .ZN(n19706) );
  INV_X1 U22208 ( .A(n19266), .ZN(n19275) );
  NAND2_X1 U22209 ( .A1(n19935), .A2(n19946), .ZN(n19345) );
  OR2_X1 U22210 ( .A1(n19345), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19288) );
  NOR2_X1 U22211 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19288), .ZN(
        n19276) );
  AOI22_X1 U22212 ( .A1(n19815), .A2(n19761), .B1(n19692), .B2(n19276), .ZN(
        n19246) );
  AOI21_X1 U22213 ( .B1(n19800), .B2(n19319), .A(n19924), .ZN(n19236) );
  NOR2_X1 U22214 ( .A1(n19236), .A2(n19931), .ZN(n19241) );
  INV_X1 U22215 ( .A(n19760), .ZN(n19810) );
  AOI21_X1 U22216 ( .B1(n19242), .B2(n19938), .A(n19923), .ZN(n19237) );
  AOI21_X1 U22217 ( .B1(n19241), .B2(n19810), .A(n19237), .ZN(n19238) );
  OAI21_X1 U22218 ( .B1(n19238), .B2(n19276), .A(n19758), .ZN(n19279) );
  OAI21_X1 U22219 ( .B1(n19760), .B2(n19276), .A(n19241), .ZN(n19244) );
  OAI21_X1 U22220 ( .B1(n19242), .B2(n19276), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19243) );
  NAND2_X1 U22221 ( .A1(n19244), .A2(n19243), .ZN(n19278) );
  AOI22_X1 U22222 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19279), .B1(
        n19240), .B2(n19278), .ZN(n19245) );
  OAI211_X1 U22223 ( .C1(n19764), .C2(n19319), .A(n19246), .B(n19245), .ZN(
        P2_U3048) );
  AOI22_X1 U22224 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19274), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19273), .ZN(n19640) );
  AOI22_X1 U22225 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19274), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19273), .ZN(n19771) );
  NOR2_X2 U22226 ( .A1(n19247), .A2(n19266), .ZN(n19707) );
  AOI22_X1 U22227 ( .A1(n19815), .A2(n19637), .B1(n19707), .B2(n19276), .ZN(
        n19251) );
  AOI22_X1 U22228 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19279), .B1(
        n19249), .B2(n19278), .ZN(n19250) );
  OAI211_X1 U22229 ( .C1(n19640), .C2(n19319), .A(n19251), .B(n19250), .ZN(
        P2_U3049) );
  AOI22_X1 U22230 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19274), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19273), .ZN(n19644) );
  AOI22_X1 U22231 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19274), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19273), .ZN(n19778) );
  NOR2_X2 U22232 ( .A1(n19252), .A2(n19266), .ZN(n19710) );
  AOI22_X1 U22233 ( .A1(n19815), .A2(n19641), .B1(n19710), .B2(n19276), .ZN(
        n19256) );
  AOI22_X1 U22234 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19279), .B1(
        n19254), .B2(n19278), .ZN(n19255) );
  OAI211_X1 U22235 ( .C1(n19644), .C2(n19319), .A(n19256), .B(n19255), .ZN(
        P2_U3050) );
  AOI22_X1 U22236 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19274), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19273), .ZN(n19785) );
  AOI22_X1 U22237 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19274), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19273), .ZN(n19718) );
  AOI22_X1 U22238 ( .A1(n19815), .A2(n19782), .B1(n19713), .B2(n19276), .ZN(
        n19259) );
  NOR2_X2 U22239 ( .A1(n19257), .A2(n19665), .ZN(n19715) );
  AOI22_X1 U22240 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19279), .B1(
        n19715), .B2(n19278), .ZN(n19258) );
  OAI211_X1 U22241 ( .C1(n19785), .C2(n19319), .A(n19259), .B(n19258), .ZN(
        P2_U3051) );
  AOI22_X1 U22242 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19274), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19273), .ZN(n19724) );
  AOI22_X1 U22243 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19274), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19273), .ZN(n19792) );
  NOR2_X2 U22244 ( .A1(n10905), .A2(n19266), .ZN(n19719) );
  AOI22_X1 U22245 ( .A1(n19815), .A2(n19720), .B1(n19719), .B2(n19276), .ZN(
        n19262) );
  NOR2_X2 U22246 ( .A1(n19260), .A2(n19665), .ZN(n19721) );
  AOI22_X1 U22247 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19279), .B1(
        n19721), .B2(n19278), .ZN(n19261) );
  OAI211_X1 U22248 ( .C1(n19724), .C2(n19319), .A(n19262), .B(n19261), .ZN(
        P2_U3052) );
  INV_X1 U22249 ( .A(n19274), .ZN(n19265) );
  INV_X1 U22250 ( .A(n19273), .ZN(n19263) );
  AOI22_X1 U22251 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19274), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19273), .ZN(n19730) );
  NOR2_X2 U22252 ( .A1(n19267), .A2(n19266), .ZN(n19725) );
  AOI22_X1 U22253 ( .A1(n19815), .A2(n19796), .B1(n19725), .B2(n19276), .ZN(
        n19270) );
  NOR2_X2 U22254 ( .A1(n19268), .A2(n19665), .ZN(n19727) );
  AOI22_X1 U22255 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19279), .B1(
        n19727), .B2(n19278), .ZN(n19269) );
  OAI211_X1 U22256 ( .C1(n19801), .C2(n19319), .A(n19270), .B(n19269), .ZN(
        P2_U3053) );
  AOI22_X1 U22257 ( .A1(n19815), .A2(n19651), .B1(n19731), .B2(n19276), .ZN(
        n19272) );
  AOI22_X1 U22258 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19279), .B1(
        n19732), .B2(n19278), .ZN(n19271) );
  OAI211_X1 U22259 ( .C1(n19654), .C2(n19319), .A(n19272), .B(n19271), .ZN(
        P2_U3054) );
  AOI22_X1 U22260 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19274), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19273), .ZN(n19745) );
  AOI22_X1 U22261 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19274), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19273), .ZN(n19820) );
  AOI22_X1 U22262 ( .A1(n19815), .A2(n19738), .B1(n19737), .B2(n19276), .ZN(
        n19281) );
  AOI22_X1 U22263 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19279), .B1(
        n19741), .B2(n19278), .ZN(n19280) );
  OAI211_X1 U22264 ( .C1(n19745), .C2(n19319), .A(n19281), .B(n19280), .ZN(
        P2_U3055) );
  NOR2_X1 U22265 ( .A1(n19525), .A2(n19345), .ZN(n19291) );
  INV_X1 U22266 ( .A(n19291), .ZN(n19313) );
  NAND2_X1 U22267 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19313), .ZN(n19282) );
  NOR2_X1 U22268 ( .A1(n13368), .A2(n19282), .ZN(n19287) );
  NOR2_X1 U22269 ( .A1(n19938), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19824) );
  INV_X1 U22270 ( .A(n19288), .ZN(n19283) );
  NOR2_X1 U22271 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19283), .ZN(n19284) );
  OR3_X1 U22272 ( .A1(n19287), .A2(n19824), .A3(n19284), .ZN(n19314) );
  INV_X1 U22273 ( .A(n19240), .ZN(n19751) );
  INV_X1 U22274 ( .A(n19692), .ZN(n19750) );
  OAI22_X1 U22275 ( .A1(n19314), .A2(n19751), .B1(n19750), .B2(n19313), .ZN(
        n19285) );
  INV_X1 U22276 ( .A(n19285), .ZN(n19294) );
  NAND2_X1 U22277 ( .A1(n19286), .A2(n19530), .ZN(n19289) );
  AOI21_X1 U22278 ( .B1(n19289), .B2(n19288), .A(n19287), .ZN(n19290) );
  OAI211_X1 U22279 ( .C1(n19291), .C2(n19938), .A(n19290), .B(n19758), .ZN(
        n19316) );
  INV_X1 U22280 ( .A(n19530), .ZN(n19292) );
  INV_X1 U22281 ( .A(n19764), .ZN(n19693) );
  AOI22_X1 U22282 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19316), .B1(
        n19341), .B2(n19693), .ZN(n19293) );
  OAI211_X1 U22283 ( .C1(n19706), .C2(n19319), .A(n19294), .B(n19293), .ZN(
        P2_U3056) );
  INV_X1 U22284 ( .A(n19249), .ZN(n19766) );
  INV_X1 U22285 ( .A(n19707), .ZN(n19765) );
  OAI22_X1 U22286 ( .A1(n19314), .A2(n19766), .B1(n19765), .B2(n19313), .ZN(
        n19295) );
  INV_X1 U22287 ( .A(n19295), .ZN(n19297) );
  INV_X1 U22288 ( .A(n19640), .ZN(n19768) );
  AOI22_X1 U22289 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19316), .B1(
        n19341), .B2(n19768), .ZN(n19296) );
  OAI211_X1 U22290 ( .C1(n19771), .C2(n19319), .A(n19297), .B(n19296), .ZN(
        P2_U3057) );
  INV_X1 U22291 ( .A(n19254), .ZN(n19773) );
  INV_X1 U22292 ( .A(n19710), .ZN(n19772) );
  OAI22_X1 U22293 ( .A1(n19314), .A2(n19773), .B1(n19772), .B2(n19313), .ZN(
        n19298) );
  INV_X1 U22294 ( .A(n19298), .ZN(n19300) );
  INV_X1 U22295 ( .A(n19644), .ZN(n19775) );
  AOI22_X1 U22296 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19316), .B1(
        n19341), .B2(n19775), .ZN(n19299) );
  OAI211_X1 U22297 ( .C1(n19778), .C2(n19319), .A(n19300), .B(n19299), .ZN(
        P2_U3058) );
  INV_X1 U22298 ( .A(n19715), .ZN(n19780) );
  INV_X1 U22299 ( .A(n19713), .ZN(n19779) );
  OAI22_X1 U22300 ( .A1(n19314), .A2(n19780), .B1(n19779), .B2(n19313), .ZN(
        n19301) );
  INV_X1 U22301 ( .A(n19301), .ZN(n19303) );
  INV_X1 U22302 ( .A(n19785), .ZN(n19714) );
  AOI22_X1 U22303 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19316), .B1(
        n19341), .B2(n19714), .ZN(n19302) );
  OAI211_X1 U22304 ( .C1(n19718), .C2(n19319), .A(n19303), .B(n19302), .ZN(
        P2_U3059) );
  INV_X1 U22305 ( .A(n19721), .ZN(n19787) );
  INV_X1 U22306 ( .A(n19719), .ZN(n19786) );
  OAI22_X1 U22307 ( .A1(n19314), .A2(n19787), .B1(n19786), .B2(n19313), .ZN(
        n19304) );
  INV_X1 U22308 ( .A(n19304), .ZN(n19306) );
  INV_X1 U22309 ( .A(n19724), .ZN(n19789) );
  AOI22_X1 U22310 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19316), .B1(
        n19341), .B2(n19789), .ZN(n19305) );
  OAI211_X1 U22311 ( .C1(n19792), .C2(n19319), .A(n19306), .B(n19305), .ZN(
        P2_U3060) );
  INV_X1 U22312 ( .A(n19727), .ZN(n19794) );
  INV_X1 U22313 ( .A(n19725), .ZN(n19793) );
  OAI22_X1 U22314 ( .A1(n19314), .A2(n19794), .B1(n19793), .B2(n19313), .ZN(
        n19307) );
  INV_X1 U22315 ( .A(n19307), .ZN(n19309) );
  AOI22_X1 U22316 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19316), .B1(
        n19341), .B2(n19726), .ZN(n19308) );
  OAI211_X1 U22317 ( .C1(n19730), .C2(n19319), .A(n19309), .B(n19308), .ZN(
        P2_U3061) );
  INV_X1 U22318 ( .A(n19732), .ZN(n19803) );
  OAI22_X1 U22319 ( .A1(n19314), .A2(n19803), .B1(n19802), .B2(n19313), .ZN(
        n19310) );
  INV_X1 U22320 ( .A(n19310), .ZN(n19312) );
  AOI22_X1 U22321 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19316), .B1(
        n19341), .B2(n19805), .ZN(n19311) );
  OAI211_X1 U22322 ( .C1(n19808), .C2(n19319), .A(n19312), .B(n19311), .ZN(
        P2_U3062) );
  INV_X1 U22323 ( .A(n19741), .ZN(n19811) );
  INV_X1 U22324 ( .A(n19737), .ZN(n19809) );
  OAI22_X1 U22325 ( .A1(n19314), .A2(n19811), .B1(n19809), .B2(n19313), .ZN(
        n19315) );
  INV_X1 U22326 ( .A(n19315), .ZN(n19318) );
  INV_X1 U22327 ( .A(n19745), .ZN(n19814) );
  AOI22_X1 U22328 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19316), .B1(
        n19341), .B2(n19814), .ZN(n19317) );
  OAI211_X1 U22329 ( .C1(n19820), .C2(n19319), .A(n19318), .B(n19317), .ZN(
        P2_U3063) );
  NOR2_X1 U22330 ( .A1(n19563), .A2(n19345), .ZN(n19339) );
  OAI21_X1 U22331 ( .B1(n13369), .B2(n19339), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19320) );
  OR2_X1 U22332 ( .A1(n19568), .A2(n19345), .ZN(n19321) );
  NAND2_X1 U22333 ( .A1(n19320), .A2(n19321), .ZN(n19340) );
  AOI22_X1 U22334 ( .A1(n19340), .A2(n19240), .B1(n19692), .B2(n19339), .ZN(
        n19326) );
  AOI21_X1 U22335 ( .B1(n13588), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19324) );
  OAI21_X1 U22336 ( .B1(n19365), .B2(n19341), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19322) );
  NAND3_X1 U22337 ( .A1(n19322), .A2(n19923), .A3(n19321), .ZN(n19323) );
  OAI211_X1 U22338 ( .C1(n19339), .C2(n19324), .A(n19323), .B(n19758), .ZN(
        n19342) );
  AOI22_X1 U22339 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19342), .B1(
        n19341), .B2(n19761), .ZN(n19325) );
  OAI211_X1 U22340 ( .C1(n19764), .C2(n19374), .A(n19326), .B(n19325), .ZN(
        P2_U3064) );
  AOI22_X1 U22341 ( .A1(n19340), .A2(n19249), .B1(n19707), .B2(n19339), .ZN(
        n19328) );
  AOI22_X1 U22342 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19342), .B1(
        n19341), .B2(n19637), .ZN(n19327) );
  OAI211_X1 U22343 ( .C1(n19640), .C2(n19374), .A(n19328), .B(n19327), .ZN(
        P2_U3065) );
  AOI22_X1 U22344 ( .A1(n19340), .A2(n19254), .B1(n19710), .B2(n19339), .ZN(
        n19330) );
  AOI22_X1 U22345 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19342), .B1(
        n19341), .B2(n19641), .ZN(n19329) );
  OAI211_X1 U22346 ( .C1(n19644), .C2(n19374), .A(n19330), .B(n19329), .ZN(
        P2_U3066) );
  AOI22_X1 U22347 ( .A1(n19340), .A2(n19715), .B1(n19713), .B2(n19339), .ZN(
        n19332) );
  AOI22_X1 U22348 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19342), .B1(
        n19341), .B2(n19782), .ZN(n19331) );
  OAI211_X1 U22349 ( .C1(n19785), .C2(n19374), .A(n19332), .B(n19331), .ZN(
        P2_U3067) );
  AOI22_X1 U22350 ( .A1(n19340), .A2(n19721), .B1(n19719), .B2(n19339), .ZN(
        n19334) );
  AOI22_X1 U22351 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19342), .B1(
        n19341), .B2(n19720), .ZN(n19333) );
  OAI211_X1 U22352 ( .C1(n19724), .C2(n19374), .A(n19334), .B(n19333), .ZN(
        P2_U3068) );
  AOI22_X1 U22353 ( .A1(n19340), .A2(n19727), .B1(n19725), .B2(n19339), .ZN(
        n19336) );
  AOI22_X1 U22354 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19342), .B1(
        n19341), .B2(n19796), .ZN(n19335) );
  OAI211_X1 U22355 ( .C1(n19801), .C2(n19374), .A(n19336), .B(n19335), .ZN(
        P2_U3069) );
  AOI22_X1 U22356 ( .A1(n19340), .A2(n19732), .B1(n19731), .B2(n19339), .ZN(
        n19338) );
  AOI22_X1 U22357 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19342), .B1(
        n19341), .B2(n19651), .ZN(n19337) );
  OAI211_X1 U22358 ( .C1(n19654), .C2(n19374), .A(n19338), .B(n19337), .ZN(
        P2_U3070) );
  AOI22_X1 U22359 ( .A1(n19340), .A2(n19741), .B1(n19737), .B2(n19339), .ZN(
        n19344) );
  AOI22_X1 U22360 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19342), .B1(
        n19341), .B2(n19738), .ZN(n19343) );
  OAI211_X1 U22361 ( .C1(n19745), .C2(n19374), .A(n19344), .B(n19343), .ZN(
        P2_U3071) );
  NOR2_X2 U22362 ( .A1(n19415), .A2(n19598), .ZN(n19401) );
  INV_X1 U22363 ( .A(n19401), .ZN(n19368) );
  NOR2_X1 U22364 ( .A1(n19592), .A2(n19345), .ZN(n19369) );
  AOI22_X1 U22365 ( .A1(n19365), .A2(n19761), .B1(n19369), .B2(n19692), .ZN(
        n19354) );
  OAI21_X1 U22366 ( .B1(n19405), .B2(n19598), .A(n19923), .ZN(n19352) );
  NOR2_X1 U22367 ( .A1(n19955), .A2(n19345), .ZN(n19349) );
  INV_X1 U22368 ( .A(n13367), .ZN(n19347) );
  INV_X1 U22369 ( .A(n19369), .ZN(n19346) );
  OAI211_X1 U22370 ( .C1(n19347), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19346), 
        .B(n19931), .ZN(n19348) );
  OAI211_X1 U22371 ( .C1(n19352), .C2(n19349), .A(n19758), .B(n19348), .ZN(
        n19371) );
  INV_X1 U22372 ( .A(n19349), .ZN(n19351) );
  OAI21_X1 U22373 ( .B1(n13367), .B2(n19369), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19350) );
  OAI21_X1 U22374 ( .B1(n19352), .B2(n19351), .A(n19350), .ZN(n19370) );
  AOI22_X1 U22375 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19371), .B1(
        n19240), .B2(n19370), .ZN(n19353) );
  OAI211_X1 U22376 ( .C1(n19764), .C2(n19368), .A(n19354), .B(n19353), .ZN(
        P2_U3072) );
  AOI22_X1 U22377 ( .A1(n19637), .A2(n19365), .B1(n19369), .B2(n19707), .ZN(
        n19356) );
  AOI22_X1 U22378 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19371), .B1(
        n19249), .B2(n19370), .ZN(n19355) );
  OAI211_X1 U22379 ( .C1(n19640), .C2(n19368), .A(n19356), .B(n19355), .ZN(
        P2_U3073) );
  AOI22_X1 U22380 ( .A1(n19775), .A2(n19401), .B1(n19369), .B2(n19710), .ZN(
        n19358) );
  AOI22_X1 U22381 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19371), .B1(
        n19254), .B2(n19370), .ZN(n19357) );
  OAI211_X1 U22382 ( .C1(n19778), .C2(n19374), .A(n19358), .B(n19357), .ZN(
        P2_U3074) );
  AOI22_X1 U22383 ( .A1(n19782), .A2(n19365), .B1(n19369), .B2(n19713), .ZN(
        n19360) );
  AOI22_X1 U22384 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19371), .B1(
        n19715), .B2(n19370), .ZN(n19359) );
  OAI211_X1 U22385 ( .C1(n19785), .C2(n19368), .A(n19360), .B(n19359), .ZN(
        P2_U3075) );
  AOI22_X1 U22386 ( .A1(n19789), .A2(n19401), .B1(n19369), .B2(n19719), .ZN(
        n19362) );
  AOI22_X1 U22387 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19371), .B1(
        n19721), .B2(n19370), .ZN(n19361) );
  OAI211_X1 U22388 ( .C1(n19792), .C2(n19374), .A(n19362), .B(n19361), .ZN(
        P2_U3076) );
  AOI22_X1 U22389 ( .A1(n19726), .A2(n19401), .B1(n19369), .B2(n19725), .ZN(
        n19364) );
  AOI22_X1 U22390 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19371), .B1(
        n19727), .B2(n19370), .ZN(n19363) );
  OAI211_X1 U22391 ( .C1(n19730), .C2(n19374), .A(n19364), .B(n19363), .ZN(
        P2_U3077) );
  AOI22_X1 U22392 ( .A1(n19651), .A2(n19365), .B1(n19731), .B2(n19369), .ZN(
        n19367) );
  AOI22_X1 U22393 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19371), .B1(
        n19732), .B2(n19370), .ZN(n19366) );
  OAI211_X1 U22394 ( .C1(n19654), .C2(n19368), .A(n19367), .B(n19366), .ZN(
        P2_U3078) );
  AOI22_X1 U22395 ( .A1(n19814), .A2(n19401), .B1(n19369), .B2(n19737), .ZN(
        n19373) );
  AOI22_X1 U22396 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19371), .B1(
        n19741), .B2(n19370), .ZN(n19372) );
  OAI211_X1 U22397 ( .C1(n19820), .C2(n19374), .A(n19373), .B(n19372), .ZN(
        P2_U3079) );
  NOR2_X1 U22398 ( .A1(n19378), .A2(n19377), .ZN(n19633) );
  NAND2_X1 U22399 ( .A1(n19633), .A2(n19935), .ZN(n19383) );
  NAND3_X1 U22400 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19935), .A3(
        n19955), .ZN(n19412) );
  NOR2_X1 U22401 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19412), .ZN(
        n19399) );
  OAI21_X1 U22402 ( .B1(n19380), .B2(n19399), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19379) );
  OAI21_X1 U22403 ( .B1(n19383), .B2(n19931), .A(n19379), .ZN(n19400) );
  AOI22_X1 U22404 ( .A1(n19400), .A2(n19240), .B1(n19692), .B2(n19399), .ZN(
        n19386) );
  OAI21_X1 U22405 ( .B1(n19401), .B2(n19429), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19382) );
  AOI211_X1 U22406 ( .C1(n19380), .C2(n19938), .A(n19399), .B(n19923), .ZN(
        n19381) );
  AOI211_X1 U22407 ( .C1(n19383), .C2(n19382), .A(n19665), .B(n19381), .ZN(
        n19384) );
  AOI22_X1 U22408 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19402), .B1(
        n19401), .B2(n19761), .ZN(n19385) );
  OAI211_X1 U22409 ( .C1(n19764), .C2(n19439), .A(n19386), .B(n19385), .ZN(
        P2_U3080) );
  AOI22_X1 U22410 ( .A1(n19400), .A2(n19249), .B1(n19707), .B2(n19399), .ZN(
        n19388) );
  AOI22_X1 U22411 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19402), .B1(
        n19401), .B2(n19637), .ZN(n19387) );
  OAI211_X1 U22412 ( .C1(n19640), .C2(n19439), .A(n19388), .B(n19387), .ZN(
        P2_U3081) );
  AOI22_X1 U22413 ( .A1(n19400), .A2(n19254), .B1(n19710), .B2(n19399), .ZN(
        n19390) );
  AOI22_X1 U22414 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19402), .B1(
        n19401), .B2(n19641), .ZN(n19389) );
  OAI211_X1 U22415 ( .C1(n19644), .C2(n19439), .A(n19390), .B(n19389), .ZN(
        P2_U3082) );
  AOI22_X1 U22416 ( .A1(n19400), .A2(n19715), .B1(n19713), .B2(n19399), .ZN(
        n19392) );
  AOI22_X1 U22417 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19402), .B1(
        n19401), .B2(n19782), .ZN(n19391) );
  OAI211_X1 U22418 ( .C1(n19785), .C2(n19439), .A(n19392), .B(n19391), .ZN(
        P2_U3083) );
  AOI22_X1 U22419 ( .A1(n19400), .A2(n19721), .B1(n19719), .B2(n19399), .ZN(
        n19394) );
  AOI22_X1 U22420 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19402), .B1(
        n19401), .B2(n19720), .ZN(n19393) );
  OAI211_X1 U22421 ( .C1(n19724), .C2(n19439), .A(n19394), .B(n19393), .ZN(
        P2_U3084) );
  AOI22_X1 U22422 ( .A1(n19400), .A2(n19727), .B1(n19725), .B2(n19399), .ZN(
        n19396) );
  AOI22_X1 U22423 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19402), .B1(
        n19401), .B2(n19796), .ZN(n19395) );
  OAI211_X1 U22424 ( .C1(n19801), .C2(n19439), .A(n19396), .B(n19395), .ZN(
        P2_U3085) );
  AOI22_X1 U22425 ( .A1(n19400), .A2(n19732), .B1(n19731), .B2(n19399), .ZN(
        n19398) );
  AOI22_X1 U22426 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19402), .B1(
        n19401), .B2(n19651), .ZN(n19397) );
  OAI211_X1 U22427 ( .C1(n19654), .C2(n19439), .A(n19398), .B(n19397), .ZN(
        P2_U3086) );
  AOI22_X1 U22428 ( .A1(n19400), .A2(n19741), .B1(n19737), .B2(n19399), .ZN(
        n19404) );
  AOI22_X1 U22429 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19402), .B1(
        n19401), .B2(n19738), .ZN(n19403) );
  OAI211_X1 U22430 ( .C1(n19745), .C2(n19439), .A(n19404), .B(n19403), .ZN(
        P2_U3087) );
  OAI21_X1 U22431 ( .B1(n19405), .B2(n19414), .A(n19923), .ZN(n19413) );
  INV_X1 U22432 ( .A(n19412), .ZN(n19406) );
  OR2_X1 U22433 ( .A1(n19413), .A2(n19406), .ZN(n19410) );
  NAND2_X1 U22434 ( .A1(n13356), .A2(n19938), .ZN(n19408) );
  NOR2_X1 U22435 ( .A1(n19964), .A2(n19412), .ZN(n19441) );
  NOR2_X1 U22436 ( .A1(n19923), .A2(n19441), .ZN(n19407) );
  AOI21_X1 U22437 ( .B1(n19408), .B2(n19407), .A(n19665), .ZN(n19409) );
  INV_X1 U22438 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n19418) );
  AOI22_X1 U22439 ( .A1(n19761), .A2(n19429), .B1(n19441), .B2(n19692), .ZN(
        n19417) );
  OAI21_X1 U22440 ( .B1(n13356), .B2(n19441), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19411) );
  OAI21_X1 U22441 ( .B1(n19413), .B2(n19412), .A(n19411), .ZN(n19435) );
  NOR2_X2 U22442 ( .A1(n19415), .A2(n19414), .ZN(n19464) );
  AOI22_X1 U22443 ( .A1(n19240), .A2(n19435), .B1(n19464), .B2(n19693), .ZN(
        n19416) );
  OAI211_X1 U22444 ( .C1(n19422), .C2(n19418), .A(n19417), .B(n19416), .ZN(
        P2_U3088) );
  INV_X1 U22445 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n19421) );
  AOI22_X1 U22446 ( .A1(n19637), .A2(n19429), .B1(n19441), .B2(n19707), .ZN(
        n19420) );
  AOI22_X1 U22447 ( .A1(n19249), .A2(n19435), .B1(n19464), .B2(n19768), .ZN(
        n19419) );
  OAI211_X1 U22448 ( .C1(n19422), .C2(n19421), .A(n19420), .B(n19419), .ZN(
        P2_U3089) );
  AOI22_X1 U22449 ( .A1(n19775), .A2(n19464), .B1(n19710), .B2(n19441), .ZN(
        n19424) );
  AOI22_X1 U22450 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19436), .B1(
        n19254), .B2(n19435), .ZN(n19423) );
  OAI211_X1 U22451 ( .C1(n19778), .C2(n19439), .A(n19424), .B(n19423), .ZN(
        P2_U3090) );
  INV_X1 U22452 ( .A(n19464), .ZN(n19432) );
  AOI22_X1 U22453 ( .A1(n19782), .A2(n19429), .B1(n19441), .B2(n19713), .ZN(
        n19426) );
  AOI22_X1 U22454 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19436), .B1(
        n19715), .B2(n19435), .ZN(n19425) );
  OAI211_X1 U22455 ( .C1(n19785), .C2(n19432), .A(n19426), .B(n19425), .ZN(
        P2_U3091) );
  AOI22_X1 U22456 ( .A1(n19720), .A2(n19429), .B1(n19441), .B2(n19719), .ZN(
        n19428) );
  AOI22_X1 U22457 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19436), .B1(
        n19721), .B2(n19435), .ZN(n19427) );
  OAI211_X1 U22458 ( .C1(n19724), .C2(n19432), .A(n19428), .B(n19427), .ZN(
        P2_U3092) );
  AOI22_X1 U22459 ( .A1(n19796), .A2(n19429), .B1(n19441), .B2(n19725), .ZN(
        n19431) );
  AOI22_X1 U22460 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19436), .B1(
        n19727), .B2(n19435), .ZN(n19430) );
  OAI211_X1 U22461 ( .C1(n19801), .C2(n19432), .A(n19431), .B(n19430), .ZN(
        P2_U3093) );
  AOI22_X1 U22462 ( .A1(n19805), .A2(n19464), .B1(n19731), .B2(n19441), .ZN(
        n19434) );
  AOI22_X1 U22463 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19436), .B1(
        n19732), .B2(n19435), .ZN(n19433) );
  OAI211_X1 U22464 ( .C1(n19808), .C2(n19439), .A(n19434), .B(n19433), .ZN(
        P2_U3094) );
  AOI22_X1 U22465 ( .A1(n19814), .A2(n19464), .B1(n19441), .B2(n19737), .ZN(
        n19438) );
  AOI22_X1 U22466 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19436), .B1(
        n19741), .B2(n19435), .ZN(n19437) );
  OAI211_X1 U22467 ( .C1(n19820), .C2(n19439), .A(n19438), .B(n19437), .ZN(
        P2_U3095) );
  NOR2_X1 U22468 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19440), .ZN(
        n19462) );
  NOR2_X1 U22469 ( .A1(n19441), .A2(n19462), .ZN(n19446) );
  OAI21_X1 U22470 ( .B1(n19443), .B2(n19462), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19442) );
  OAI21_X1 U22471 ( .B1(n19446), .B2(n19931), .A(n19442), .ZN(n19463) );
  AOI22_X1 U22472 ( .A1(n19463), .A2(n19240), .B1(n19692), .B2(n19462), .ZN(
        n19449) );
  OAI21_X1 U22473 ( .B1(n19464), .B2(n19473), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19445) );
  AOI211_X1 U22474 ( .C1(n19443), .C2(n19938), .A(n19462), .B(n19923), .ZN(
        n19444) );
  AOI211_X1 U22475 ( .C1(n19446), .C2(n19445), .A(n19665), .B(n19444), .ZN(
        n19447) );
  AOI22_X1 U22476 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19465), .B1(
        n19464), .B2(n19761), .ZN(n19448) );
  OAI211_X1 U22477 ( .C1(n19764), .C2(n19487), .A(n19449), .B(n19448), .ZN(
        P2_U3096) );
  AOI22_X1 U22478 ( .A1(n19463), .A2(n19249), .B1(n19707), .B2(n19462), .ZN(
        n19451) );
  AOI22_X1 U22479 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19465), .B1(
        n19464), .B2(n19637), .ZN(n19450) );
  OAI211_X1 U22480 ( .C1(n19640), .C2(n19487), .A(n19451), .B(n19450), .ZN(
        P2_U3097) );
  AOI22_X1 U22481 ( .A1(n19463), .A2(n19254), .B1(n19710), .B2(n19462), .ZN(
        n19453) );
  AOI22_X1 U22482 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19465), .B1(
        n19464), .B2(n19641), .ZN(n19452) );
  OAI211_X1 U22483 ( .C1(n19644), .C2(n19487), .A(n19453), .B(n19452), .ZN(
        P2_U3098) );
  AOI22_X1 U22484 ( .A1(n19463), .A2(n19715), .B1(n19713), .B2(n19462), .ZN(
        n19455) );
  AOI22_X1 U22485 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19465), .B1(
        n19464), .B2(n19782), .ZN(n19454) );
  OAI211_X1 U22486 ( .C1(n19785), .C2(n19487), .A(n19455), .B(n19454), .ZN(
        P2_U3099) );
  AOI22_X1 U22487 ( .A1(n19463), .A2(n19721), .B1(n19719), .B2(n19462), .ZN(
        n19457) );
  AOI22_X1 U22488 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19465), .B1(
        n19464), .B2(n19720), .ZN(n19456) );
  OAI211_X1 U22489 ( .C1(n19724), .C2(n19487), .A(n19457), .B(n19456), .ZN(
        P2_U3100) );
  AOI22_X1 U22490 ( .A1(n19463), .A2(n19727), .B1(n19725), .B2(n19462), .ZN(
        n19459) );
  AOI22_X1 U22491 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19465), .B1(
        n19464), .B2(n19796), .ZN(n19458) );
  OAI211_X1 U22492 ( .C1(n19801), .C2(n19487), .A(n19459), .B(n19458), .ZN(
        P2_U3101) );
  AOI22_X1 U22493 ( .A1(n19463), .A2(n19732), .B1(n19731), .B2(n19462), .ZN(
        n19461) );
  AOI22_X1 U22494 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19465), .B1(
        n19464), .B2(n19651), .ZN(n19460) );
  OAI211_X1 U22495 ( .C1(n19654), .C2(n19487), .A(n19461), .B(n19460), .ZN(
        P2_U3102) );
  AOI22_X1 U22496 ( .A1(n19463), .A2(n19741), .B1(n19737), .B2(n19462), .ZN(
        n19467) );
  AOI22_X1 U22497 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19465), .B1(
        n19464), .B2(n19738), .ZN(n19466) );
  OAI211_X1 U22498 ( .C1(n19745), .C2(n19487), .A(n19467), .B(n19466), .ZN(
        P2_U3103) );
  INV_X1 U22499 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n19470) );
  AOI22_X1 U22500 ( .A1(n19483), .A2(n19240), .B1(n19692), .B2(n19491), .ZN(
        n19469) );
  AOI22_X1 U22501 ( .A1(n19473), .A2(n19761), .B1(n19516), .B2(n19693), .ZN(
        n19468) );
  OAI211_X1 U22502 ( .C1(n19476), .C2(n19470), .A(n19469), .B(n19468), .ZN(
        P2_U3104) );
  AOI22_X1 U22503 ( .A1(n19483), .A2(n19249), .B1(n19707), .B2(n19491), .ZN(
        n19472) );
  AOI22_X1 U22504 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19484), .B1(
        n19516), .B2(n19768), .ZN(n19471) );
  OAI211_X1 U22505 ( .C1(n19771), .C2(n19487), .A(n19472), .B(n19471), .ZN(
        P2_U3105) );
  AOI22_X1 U22506 ( .A1(n19483), .A2(n19254), .B1(n19710), .B2(n19491), .ZN(
        n19475) );
  AOI22_X1 U22507 ( .A1(n19473), .A2(n19641), .B1(n19516), .B2(n19775), .ZN(
        n19474) );
  OAI211_X1 U22508 ( .C1(n19476), .C2(n11169), .A(n19475), .B(n19474), .ZN(
        P2_U3106) );
  AOI22_X1 U22509 ( .A1(n19483), .A2(n19715), .B1(n19713), .B2(n19491), .ZN(
        n19478) );
  AOI22_X1 U22510 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19484), .B1(
        n19516), .B2(n19714), .ZN(n19477) );
  OAI211_X1 U22511 ( .C1(n19718), .C2(n19487), .A(n19478), .B(n19477), .ZN(
        P2_U3107) );
  AOI22_X1 U22512 ( .A1(n19483), .A2(n19721), .B1(n19719), .B2(n19491), .ZN(
        n19480) );
  AOI22_X1 U22513 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19484), .B1(
        n19516), .B2(n19789), .ZN(n19479) );
  OAI211_X1 U22514 ( .C1(n19792), .C2(n19487), .A(n19480), .B(n19479), .ZN(
        P2_U3108) );
  AOI22_X1 U22515 ( .A1(n19483), .A2(n19727), .B1(n19725), .B2(n19491), .ZN(
        n19482) );
  AOI22_X1 U22516 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19484), .B1(
        n19516), .B2(n19726), .ZN(n19481) );
  OAI211_X1 U22517 ( .C1(n19730), .C2(n19487), .A(n19482), .B(n19481), .ZN(
        P2_U3109) );
  AOI22_X1 U22518 ( .A1(n19483), .A2(n19741), .B1(n19737), .B2(n19491), .ZN(
        n19486) );
  AOI22_X1 U22519 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19484), .B1(
        n19516), .B2(n19814), .ZN(n19485) );
  OAI211_X1 U22520 ( .C1(n19820), .C2(n19487), .A(n19486), .B(n19485), .ZN(
        P2_U3111) );
  NAND2_X1 U22521 ( .A1(n19690), .A2(n19530), .ZN(n19548) );
  INV_X1 U22522 ( .A(n19516), .ZN(n19489) );
  AOI21_X1 U22523 ( .B1(n19548), .B2(n19489), .A(n19924), .ZN(n19490) );
  NOR2_X1 U22524 ( .A1(n19490), .A2(n19931), .ZN(n19493) );
  NAND2_X1 U22525 ( .A1(n19946), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19597) );
  INV_X1 U22526 ( .A(n19597), .ZN(n19591) );
  NAND2_X1 U22527 ( .A1(n19591), .A2(n19955), .ZN(n19532) );
  NOR2_X1 U22528 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19532), .ZN(
        n19515) );
  NOR2_X1 U22529 ( .A1(n19515), .A2(n19491), .ZN(n19494) );
  AOI211_X1 U22530 ( .C1(n13365), .C2(n19938), .A(n19515), .B(n19923), .ZN(
        n19492) );
  INV_X1 U22531 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n19499) );
  AOI22_X1 U22532 ( .A1(n19551), .A2(n19693), .B1(n19692), .B2(n19515), .ZN(
        n19498) );
  INV_X1 U22533 ( .A(n19493), .ZN(n19496) );
  OAI21_X1 U22534 ( .B1(n13365), .B2(n19515), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19495) );
  AOI22_X1 U22535 ( .A1(n19240), .A2(n19517), .B1(n19516), .B2(n19761), .ZN(
        n19497) );
  OAI211_X1 U22536 ( .C1(n19521), .C2(n19499), .A(n19498), .B(n19497), .ZN(
        P2_U3112) );
  INV_X1 U22537 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n19502) );
  AOI22_X1 U22538 ( .A1(n19551), .A2(n19768), .B1(n19707), .B2(n19515), .ZN(
        n19501) );
  AOI22_X1 U22539 ( .A1(n19249), .A2(n19517), .B1(n19516), .B2(n19637), .ZN(
        n19500) );
  OAI211_X1 U22540 ( .C1(n19521), .C2(n19502), .A(n19501), .B(n19500), .ZN(
        P2_U3113) );
  AOI22_X1 U22541 ( .A1(n19551), .A2(n19775), .B1(n19710), .B2(n19515), .ZN(
        n19504) );
  AOI22_X1 U22542 ( .A1(n19254), .A2(n19517), .B1(n19516), .B2(n19641), .ZN(
        n19503) );
  OAI211_X1 U22543 ( .C1(n19521), .C2(n11170), .A(n19504), .B(n19503), .ZN(
        P2_U3114) );
  INV_X1 U22544 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n19507) );
  AOI22_X1 U22545 ( .A1(n19551), .A2(n19714), .B1(n19713), .B2(n19515), .ZN(
        n19506) );
  AOI22_X1 U22546 ( .A1(n19715), .A2(n19517), .B1(n19516), .B2(n19782), .ZN(
        n19505) );
  OAI211_X1 U22547 ( .C1(n19521), .C2(n19507), .A(n19506), .B(n19505), .ZN(
        P2_U3115) );
  INV_X1 U22548 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n19510) );
  AOI22_X1 U22549 ( .A1(n19551), .A2(n19789), .B1(n19719), .B2(n19515), .ZN(
        n19509) );
  AOI22_X1 U22550 ( .A1(n19721), .A2(n19517), .B1(n19516), .B2(n19720), .ZN(
        n19508) );
  OAI211_X1 U22551 ( .C1(n19521), .C2(n19510), .A(n19509), .B(n19508), .ZN(
        P2_U3116) );
  AOI22_X1 U22552 ( .A1(n19726), .A2(n19551), .B1(n19725), .B2(n19515), .ZN(
        n19512) );
  AOI22_X1 U22553 ( .A1(n19727), .A2(n19517), .B1(n19516), .B2(n19796), .ZN(
        n19511) );
  OAI211_X1 U22554 ( .C1(n19521), .C2(n11212), .A(n19512), .B(n19511), .ZN(
        P2_U3117) );
  AOI22_X1 U22555 ( .A1(n19551), .A2(n19805), .B1(n19731), .B2(n19515), .ZN(
        n19514) );
  AOI22_X1 U22556 ( .A1(n19732), .A2(n19517), .B1(n19516), .B2(n19651), .ZN(
        n19513) );
  OAI211_X1 U22557 ( .C1(n19521), .C2(n13582), .A(n19514), .B(n19513), .ZN(
        P2_U3118) );
  INV_X1 U22558 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n19520) );
  AOI22_X1 U22559 ( .A1(n19551), .A2(n19814), .B1(n19737), .B2(n19515), .ZN(
        n19519) );
  AOI22_X1 U22560 ( .A1(n19741), .A2(n19517), .B1(n19516), .B2(n19738), .ZN(
        n19518) );
  OAI211_X1 U22561 ( .C1(n19521), .C2(n19520), .A(n19519), .B(n19518), .ZN(
        P2_U3119) );
  NOR2_X1 U22562 ( .A1(n19522), .A2(n19924), .ZN(n19754) );
  NAND2_X1 U22563 ( .A1(n19754), .A2(n19530), .ZN(n19523) );
  NAND2_X1 U22564 ( .A1(n19523), .A2(n19923), .ZN(n19533) );
  INV_X1 U22565 ( .A(n19532), .ZN(n19524) );
  OR2_X1 U22566 ( .A1(n19533), .A2(n19524), .ZN(n19529) );
  NOR2_X1 U22567 ( .A1(n19525), .A2(n19597), .ZN(n19559) );
  INV_X1 U22568 ( .A(n19559), .ZN(n19526) );
  OAI211_X1 U22569 ( .C1(n13357), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19526), 
        .B(n19931), .ZN(n19527) );
  AND2_X1 U22570 ( .A1(n19527), .A2(n19758), .ZN(n19528) );
  AND2_X1 U22571 ( .A1(n19529), .A2(n19528), .ZN(n19537) );
  INV_X1 U22572 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n19536) );
  AOI22_X1 U22573 ( .A1(n19693), .A2(n19587), .B1(n19692), .B2(n19559), .ZN(
        n19535) );
  OAI21_X1 U22574 ( .B1(n13190), .B2(n19559), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19531) );
  OAI21_X1 U22575 ( .B1(n19533), .B2(n19532), .A(n19531), .ZN(n19552) );
  AOI22_X1 U22576 ( .A1(n19240), .A2(n19552), .B1(n19551), .B2(n19761), .ZN(
        n19534) );
  OAI211_X1 U22577 ( .C1(n19537), .C2(n19536), .A(n19535), .B(n19534), .ZN(
        P2_U3120) );
  AOI22_X1 U22578 ( .A1(n19551), .A2(n19637), .B1(n19707), .B2(n19559), .ZN(
        n19539) );
  INV_X1 U22579 ( .A(n19537), .ZN(n19553) );
  AOI22_X1 U22580 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19553), .B1(
        n19249), .B2(n19552), .ZN(n19538) );
  OAI211_X1 U22581 ( .C1(n19640), .C2(n19557), .A(n19539), .B(n19538), .ZN(
        P2_U3121) );
  AOI22_X1 U22582 ( .A1(n19551), .A2(n19641), .B1(n19710), .B2(n19559), .ZN(
        n19541) );
  AOI22_X1 U22583 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19553), .B1(
        n19254), .B2(n19552), .ZN(n19540) );
  OAI211_X1 U22584 ( .C1(n19644), .C2(n19557), .A(n19541), .B(n19540), .ZN(
        P2_U3122) );
  AOI22_X1 U22585 ( .A1(n19714), .A2(n19587), .B1(n19713), .B2(n19559), .ZN(
        n19543) );
  AOI22_X1 U22586 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19553), .B1(
        n19715), .B2(n19552), .ZN(n19542) );
  OAI211_X1 U22587 ( .C1(n19718), .C2(n19548), .A(n19543), .B(n19542), .ZN(
        P2_U3123) );
  AOI22_X1 U22588 ( .A1(n19789), .A2(n19587), .B1(n19719), .B2(n19559), .ZN(
        n19545) );
  AOI22_X1 U22589 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19553), .B1(
        n19721), .B2(n19552), .ZN(n19544) );
  OAI211_X1 U22590 ( .C1(n19792), .C2(n19548), .A(n19545), .B(n19544), .ZN(
        P2_U3124) );
  AOI22_X1 U22591 ( .A1(n19726), .A2(n19587), .B1(n19725), .B2(n19559), .ZN(
        n19547) );
  AOI22_X1 U22592 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19553), .B1(
        n19727), .B2(n19552), .ZN(n19546) );
  OAI211_X1 U22593 ( .C1(n19730), .C2(n19548), .A(n19547), .B(n19546), .ZN(
        P2_U3125) );
  AOI22_X1 U22594 ( .A1(n19551), .A2(n19651), .B1(n19731), .B2(n19559), .ZN(
        n19550) );
  AOI22_X1 U22595 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19553), .B1(
        n19732), .B2(n19552), .ZN(n19549) );
  OAI211_X1 U22596 ( .C1(n19654), .C2(n19557), .A(n19550), .B(n19549), .ZN(
        P2_U3126) );
  AOI22_X1 U22597 ( .A1(n19551), .A2(n19738), .B1(n19737), .B2(n19559), .ZN(
        n19555) );
  AOI22_X1 U22598 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19553), .B1(
        n19741), .B2(n19552), .ZN(n19554) );
  OAI211_X1 U22599 ( .C1(n19745), .C2(n19557), .A(n19555), .B(n19554), .ZN(
        P2_U3127) );
  NAND2_X1 U22600 ( .A1(n13366), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19562) );
  INV_X1 U22601 ( .A(n19690), .ZN(n19556) );
  AOI21_X1 U22602 ( .B1(n19614), .B2(n19557), .A(n19924), .ZN(n19558) );
  NOR2_X1 U22603 ( .A1(n19559), .A2(n19558), .ZN(n19560) );
  NOR2_X1 U22604 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19560), .ZN(n19561) );
  NAND2_X1 U22605 ( .A1(n19562), .A2(n19561), .ZN(n19565) );
  NOR2_X1 U22606 ( .A1(n19563), .A2(n19597), .ZN(n19585) );
  INV_X1 U22607 ( .A(n19585), .ZN(n19564) );
  AOI21_X1 U22608 ( .B1(n19565), .B2(n19564), .A(n19665), .ZN(n19574) );
  OAI21_X1 U22609 ( .B1(n19566), .B2(n19585), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19567) );
  OAI21_X1 U22610 ( .B1(n19597), .B2(n19568), .A(n19567), .ZN(n19586) );
  AOI22_X1 U22611 ( .A1(n19586), .A2(n19240), .B1(n19692), .B2(n19585), .ZN(
        n19570) );
  AOI22_X1 U22612 ( .A1(n19587), .A2(n19761), .B1(n19619), .B2(n19693), .ZN(
        n19569) );
  OAI211_X1 U22613 ( .C1(n19574), .C2(n11245), .A(n19570), .B(n19569), .ZN(
        P2_U3128) );
  AOI22_X1 U22614 ( .A1(n19586), .A2(n19249), .B1(n19707), .B2(n19585), .ZN(
        n19572) );
  AOI22_X1 U22615 ( .A1(n19587), .A2(n19637), .B1(n19619), .B2(n19768), .ZN(
        n19571) );
  OAI211_X1 U22616 ( .C1(n19574), .C2(n19573), .A(n19572), .B(n19571), .ZN(
        P2_U3129) );
  AOI22_X1 U22617 ( .A1(n19586), .A2(n19254), .B1(n19710), .B2(n19585), .ZN(
        n19576) );
  AOI22_X1 U22618 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19588), .B1(
        n19587), .B2(n19641), .ZN(n19575) );
  OAI211_X1 U22619 ( .C1(n19644), .C2(n19614), .A(n19576), .B(n19575), .ZN(
        P2_U3130) );
  AOI22_X1 U22620 ( .A1(n19586), .A2(n19715), .B1(n19713), .B2(n19585), .ZN(
        n19578) );
  AOI22_X1 U22621 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19588), .B1(
        n19587), .B2(n19782), .ZN(n19577) );
  OAI211_X1 U22622 ( .C1(n19785), .C2(n19614), .A(n19578), .B(n19577), .ZN(
        P2_U3131) );
  AOI22_X1 U22623 ( .A1(n19586), .A2(n19721), .B1(n19719), .B2(n19585), .ZN(
        n19580) );
  AOI22_X1 U22624 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19588), .B1(
        n19587), .B2(n19720), .ZN(n19579) );
  OAI211_X1 U22625 ( .C1(n19724), .C2(n19614), .A(n19580), .B(n19579), .ZN(
        P2_U3132) );
  AOI22_X1 U22626 ( .A1(n19586), .A2(n19727), .B1(n19725), .B2(n19585), .ZN(
        n19582) );
  AOI22_X1 U22627 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19588), .B1(
        n19587), .B2(n19796), .ZN(n19581) );
  OAI211_X1 U22628 ( .C1(n19801), .C2(n19614), .A(n19582), .B(n19581), .ZN(
        P2_U3133) );
  AOI22_X1 U22629 ( .A1(n19586), .A2(n19732), .B1(n19731), .B2(n19585), .ZN(
        n19584) );
  AOI22_X1 U22630 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19588), .B1(
        n19587), .B2(n19651), .ZN(n19583) );
  OAI211_X1 U22631 ( .C1(n19654), .C2(n19614), .A(n19584), .B(n19583), .ZN(
        P2_U3134) );
  AOI22_X1 U22632 ( .A1(n19586), .A2(n19741), .B1(n19737), .B2(n19585), .ZN(
        n19590) );
  AOI22_X1 U22633 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19588), .B1(
        n19587), .B2(n19738), .ZN(n19589) );
  OAI211_X1 U22634 ( .C1(n19745), .C2(n19614), .A(n19590), .B(n19589), .ZN(
        P2_U3135) );
  NAND2_X1 U22635 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19591), .ZN(
        n19595) );
  NOR2_X1 U22636 ( .A1(n19592), .A2(n19597), .ZN(n19617) );
  OAI21_X1 U22637 ( .B1(n19593), .B2(n19617), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19594) );
  OAI21_X1 U22638 ( .B1(n19595), .B2(n19931), .A(n19594), .ZN(n19618) );
  AOI22_X1 U22639 ( .A1(n19618), .A2(n19240), .B1(n19692), .B2(n19617), .ZN(
        n19603) );
  AOI21_X1 U22640 ( .B1(n19596), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19601) );
  INV_X1 U22641 ( .A(n19754), .ZN(n19599) );
  OAI22_X1 U22642 ( .A1(n19599), .A2(n19598), .B1(n19597), .B2(n19955), .ZN(
        n19600) );
  OAI211_X1 U22643 ( .C1(n19617), .C2(n19601), .A(n19600), .B(n19758), .ZN(
        n19620) );
  NAND2_X1 U22644 ( .A1(n19670), .A2(n19922), .ZN(n19628) );
  AOI22_X1 U22645 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19620), .B1(
        n19657), .B2(n19693), .ZN(n19602) );
  OAI211_X1 U22646 ( .C1(n19706), .C2(n19614), .A(n19603), .B(n19602), .ZN(
        P2_U3136) );
  AOI22_X1 U22647 ( .A1(n19618), .A2(n19249), .B1(n19707), .B2(n19617), .ZN(
        n19605) );
  AOI22_X1 U22648 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19620), .B1(
        n19657), .B2(n19768), .ZN(n19604) );
  OAI211_X1 U22649 ( .C1(n19771), .C2(n19614), .A(n19605), .B(n19604), .ZN(
        P2_U3137) );
  AOI22_X1 U22650 ( .A1(n19618), .A2(n19254), .B1(n19710), .B2(n19617), .ZN(
        n19607) );
  AOI22_X1 U22651 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19620), .B1(
        n19619), .B2(n19641), .ZN(n19606) );
  OAI211_X1 U22652 ( .C1(n19644), .C2(n19628), .A(n19607), .B(n19606), .ZN(
        P2_U3138) );
  AOI22_X1 U22653 ( .A1(n19618), .A2(n19715), .B1(n19713), .B2(n19617), .ZN(
        n19609) );
  AOI22_X1 U22654 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19620), .B1(
        n19657), .B2(n19714), .ZN(n19608) );
  OAI211_X1 U22655 ( .C1(n19718), .C2(n19614), .A(n19609), .B(n19608), .ZN(
        P2_U3139) );
  AOI22_X1 U22656 ( .A1(n19618), .A2(n19721), .B1(n19719), .B2(n19617), .ZN(
        n19611) );
  AOI22_X1 U22657 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19620), .B1(
        n19619), .B2(n19720), .ZN(n19610) );
  OAI211_X1 U22658 ( .C1(n19724), .C2(n19628), .A(n19611), .B(n19610), .ZN(
        P2_U3140) );
  AOI22_X1 U22659 ( .A1(n19618), .A2(n19727), .B1(n19725), .B2(n19617), .ZN(
        n19613) );
  AOI22_X1 U22660 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19620), .B1(
        n19657), .B2(n19726), .ZN(n19612) );
  OAI211_X1 U22661 ( .C1(n19730), .C2(n19614), .A(n19613), .B(n19612), .ZN(
        P2_U3141) );
  AOI22_X1 U22662 ( .A1(n19618), .A2(n19732), .B1(n19731), .B2(n19617), .ZN(
        n19616) );
  AOI22_X1 U22663 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19620), .B1(
        n19619), .B2(n19651), .ZN(n19615) );
  OAI211_X1 U22664 ( .C1(n19654), .C2(n19628), .A(n19616), .B(n19615), .ZN(
        P2_U3142) );
  AOI22_X1 U22665 ( .A1(n19618), .A2(n19741), .B1(n19737), .B2(n19617), .ZN(
        n19622) );
  AOI22_X1 U22666 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19620), .B1(
        n19619), .B2(n19738), .ZN(n19621) );
  OAI211_X1 U22667 ( .C1(n19745), .C2(n19628), .A(n19622), .B(n19621), .ZN(
        P2_U3143) );
  INV_X1 U22668 ( .A(n19623), .ZN(n19627) );
  INV_X1 U22669 ( .A(n19633), .ZN(n19626) );
  NAND3_X1 U22670 ( .A1(n19955), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19661) );
  INV_X1 U22671 ( .A(n19661), .ZN(n19668) );
  NAND2_X1 U22672 ( .A1(n19964), .A2(n19668), .ZN(n19629) );
  INV_X1 U22673 ( .A(n19629), .ZN(n19655) );
  OAI21_X1 U22674 ( .B1(n19624), .B2(n19655), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19625) );
  OAI21_X1 U22675 ( .B1(n19627), .B2(n19626), .A(n19625), .ZN(n19656) );
  AOI22_X1 U22676 ( .A1(n19656), .A2(n19240), .B1(n19692), .B2(n19655), .ZN(
        n19636) );
  AOI21_X1 U22677 ( .B1(n19689), .B2(n19628), .A(n19924), .ZN(n19634) );
  OAI211_X1 U22678 ( .C1(n19630), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19629), 
        .B(n19931), .ZN(n19631) );
  AND2_X1 U22679 ( .A1(n19631), .A2(n19758), .ZN(n19632) );
  OAI211_X1 U22680 ( .C1(n19634), .C2(n19633), .A(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n19632), .ZN(n19658) );
  AOI22_X1 U22681 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19658), .B1(
        n19657), .B2(n19761), .ZN(n19635) );
  OAI211_X1 U22682 ( .C1(n19764), .C2(n19689), .A(n19636), .B(n19635), .ZN(
        P2_U3144) );
  AOI22_X1 U22683 ( .A1(n19656), .A2(n19249), .B1(n19707), .B2(n19655), .ZN(
        n19639) );
  AOI22_X1 U22684 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19658), .B1(
        n19657), .B2(n19637), .ZN(n19638) );
  OAI211_X1 U22685 ( .C1(n19640), .C2(n19689), .A(n19639), .B(n19638), .ZN(
        P2_U3145) );
  AOI22_X1 U22686 ( .A1(n19656), .A2(n19254), .B1(n19710), .B2(n19655), .ZN(
        n19643) );
  AOI22_X1 U22687 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19658), .B1(
        n19657), .B2(n19641), .ZN(n19642) );
  OAI211_X1 U22688 ( .C1(n19644), .C2(n19689), .A(n19643), .B(n19642), .ZN(
        P2_U3146) );
  AOI22_X1 U22689 ( .A1(n19656), .A2(n19715), .B1(n19713), .B2(n19655), .ZN(
        n19646) );
  AOI22_X1 U22690 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19658), .B1(
        n19657), .B2(n19782), .ZN(n19645) );
  OAI211_X1 U22691 ( .C1(n19785), .C2(n19689), .A(n19646), .B(n19645), .ZN(
        P2_U3147) );
  AOI22_X1 U22692 ( .A1(n19656), .A2(n19721), .B1(n19719), .B2(n19655), .ZN(
        n19648) );
  AOI22_X1 U22693 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19658), .B1(
        n19657), .B2(n19720), .ZN(n19647) );
  OAI211_X1 U22694 ( .C1(n19724), .C2(n19689), .A(n19648), .B(n19647), .ZN(
        P2_U3148) );
  AOI22_X1 U22695 ( .A1(n19656), .A2(n19727), .B1(n19725), .B2(n19655), .ZN(
        n19650) );
  AOI22_X1 U22696 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19658), .B1(
        n19657), .B2(n19796), .ZN(n19649) );
  OAI211_X1 U22697 ( .C1(n19801), .C2(n19689), .A(n19650), .B(n19649), .ZN(
        P2_U3149) );
  AOI22_X1 U22698 ( .A1(n19656), .A2(n19732), .B1(n19731), .B2(n19655), .ZN(
        n19653) );
  AOI22_X1 U22699 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19658), .B1(
        n19657), .B2(n19651), .ZN(n19652) );
  OAI211_X1 U22700 ( .C1(n19654), .C2(n19689), .A(n19653), .B(n19652), .ZN(
        P2_U3150) );
  AOI22_X1 U22701 ( .A1(n19656), .A2(n19741), .B1(n19737), .B2(n19655), .ZN(
        n19660) );
  AOI22_X1 U22702 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19658), .B1(
        n19657), .B2(n19738), .ZN(n19659) );
  OAI211_X1 U22703 ( .C1(n19745), .C2(n19689), .A(n19660), .B(n19659), .ZN(
        P2_U3151) );
  NOR2_X1 U22704 ( .A1(n19964), .A2(n19661), .ZN(n19695) );
  NOR3_X1 U22705 ( .A1(n19662), .A2(n19695), .A3(n19825), .ZN(n19664) );
  AOI21_X1 U22706 ( .B1(n19938), .B2(n19668), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19663) );
  AOI22_X1 U22707 ( .A1(n19685), .A2(n19240), .B1(n19692), .B2(n19695), .ZN(
        n19672) );
  INV_X1 U22708 ( .A(n19695), .ZN(n19666) );
  AOI211_X1 U22709 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19666), .A(n19665), 
        .B(n19664), .ZN(n19667) );
  OAI221_X1 U22710 ( .B1(n19668), .B2(n19669), .C1(n19668), .C2(n19754), .A(
        n19667), .ZN(n19686) );
  AOI22_X1 U22711 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19686), .B1(
        n19739), .B2(n19693), .ZN(n19671) );
  OAI211_X1 U22712 ( .C1(n19706), .C2(n19689), .A(n19672), .B(n19671), .ZN(
        P2_U3152) );
  AOI22_X1 U22713 ( .A1(n19685), .A2(n19249), .B1(n19707), .B2(n19695), .ZN(
        n19674) );
  AOI22_X1 U22714 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19686), .B1(
        n19739), .B2(n19768), .ZN(n19673) );
  OAI211_X1 U22715 ( .C1(n19771), .C2(n19689), .A(n19674), .B(n19673), .ZN(
        P2_U3153) );
  AOI22_X1 U22716 ( .A1(n19685), .A2(n19254), .B1(n19710), .B2(n19695), .ZN(
        n19676) );
  AOI22_X1 U22717 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19686), .B1(
        n19739), .B2(n19775), .ZN(n19675) );
  OAI211_X1 U22718 ( .C1(n19778), .C2(n19689), .A(n19676), .B(n19675), .ZN(
        P2_U3154) );
  AOI22_X1 U22719 ( .A1(n19685), .A2(n19715), .B1(n19713), .B2(n19695), .ZN(
        n19678) );
  AOI22_X1 U22720 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19686), .B1(
        n19739), .B2(n19714), .ZN(n19677) );
  OAI211_X1 U22721 ( .C1(n19718), .C2(n19689), .A(n19678), .B(n19677), .ZN(
        P2_U3155) );
  AOI22_X1 U22722 ( .A1(n19685), .A2(n19721), .B1(n19719), .B2(n19695), .ZN(
        n19680) );
  AOI22_X1 U22723 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19686), .B1(
        n19739), .B2(n19789), .ZN(n19679) );
  OAI211_X1 U22724 ( .C1(n19792), .C2(n19689), .A(n19680), .B(n19679), .ZN(
        P2_U3156) );
  AOI22_X1 U22725 ( .A1(n19685), .A2(n19727), .B1(n19725), .B2(n19695), .ZN(
        n19682) );
  AOI22_X1 U22726 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19686), .B1(
        n19739), .B2(n19726), .ZN(n19681) );
  OAI211_X1 U22727 ( .C1(n19730), .C2(n19689), .A(n19682), .B(n19681), .ZN(
        P2_U3157) );
  AOI22_X1 U22728 ( .A1(n19685), .A2(n19732), .B1(n19731), .B2(n19695), .ZN(
        n19684) );
  AOI22_X1 U22729 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19686), .B1(
        n19739), .B2(n19805), .ZN(n19683) );
  OAI211_X1 U22730 ( .C1(n19808), .C2(n19689), .A(n19684), .B(n19683), .ZN(
        P2_U3158) );
  AOI22_X1 U22731 ( .A1(n19685), .A2(n19741), .B1(n19737), .B2(n19695), .ZN(
        n19688) );
  AOI22_X1 U22732 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19686), .B1(
        n19739), .B2(n19814), .ZN(n19687) );
  OAI211_X1 U22733 ( .C1(n19820), .C2(n19689), .A(n19688), .B(n19687), .ZN(
        P2_U3159) );
  NAND2_X1 U22734 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19691), .ZN(
        n19756) );
  NOR2_X1 U22735 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19756), .ZN(
        n19736) );
  AOI22_X1 U22736 ( .A1(n19797), .A2(n19693), .B1(n19692), .B2(n19736), .ZN(
        n19705) );
  OAI21_X1 U22737 ( .B1(n19797), .B2(n19739), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19694) );
  NAND2_X1 U22738 ( .A1(n19694), .A2(n19923), .ZN(n19703) );
  NOR2_X1 U22739 ( .A1(n19736), .A2(n19695), .ZN(n19702) );
  INV_X1 U22740 ( .A(n19702), .ZN(n19699) );
  INV_X1 U22741 ( .A(n19700), .ZN(n19697) );
  INV_X1 U22742 ( .A(n19736), .ZN(n19696) );
  OAI211_X1 U22743 ( .C1(n19697), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19696), 
        .B(n19931), .ZN(n19698) );
  OAI211_X1 U22744 ( .C1(n19703), .C2(n19699), .A(n19758), .B(n19698), .ZN(
        n19742) );
  OAI21_X1 U22745 ( .B1(n19700), .B2(n19736), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19701) );
  AOI22_X1 U22746 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19742), .B1(
        n19240), .B2(n19740), .ZN(n19704) );
  OAI211_X1 U22747 ( .C1(n19706), .C2(n19735), .A(n19705), .B(n19704), .ZN(
        P2_U3160) );
  AOI22_X1 U22748 ( .A1(n19797), .A2(n19768), .B1(n19707), .B2(n19736), .ZN(
        n19709) );
  AOI22_X1 U22749 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19742), .B1(
        n19249), .B2(n19740), .ZN(n19708) );
  OAI211_X1 U22750 ( .C1(n19771), .C2(n19735), .A(n19709), .B(n19708), .ZN(
        P2_U3161) );
  AOI22_X1 U22751 ( .A1(n19797), .A2(n19775), .B1(n19710), .B2(n19736), .ZN(
        n19712) );
  AOI22_X1 U22752 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19742), .B1(
        n19254), .B2(n19740), .ZN(n19711) );
  OAI211_X1 U22753 ( .C1(n19778), .C2(n19735), .A(n19712), .B(n19711), .ZN(
        P2_U3162) );
  AOI22_X1 U22754 ( .A1(n19797), .A2(n19714), .B1(n19713), .B2(n19736), .ZN(
        n19717) );
  AOI22_X1 U22755 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19742), .B1(
        n19715), .B2(n19740), .ZN(n19716) );
  OAI211_X1 U22756 ( .C1(n19718), .C2(n19735), .A(n19717), .B(n19716), .ZN(
        P2_U3163) );
  AOI22_X1 U22757 ( .A1(n19739), .A2(n19720), .B1(n19719), .B2(n19736), .ZN(
        n19723) );
  AOI22_X1 U22758 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19742), .B1(
        n19721), .B2(n19740), .ZN(n19722) );
  OAI211_X1 U22759 ( .C1(n19724), .C2(n19819), .A(n19723), .B(n19722), .ZN(
        P2_U3164) );
  AOI22_X1 U22760 ( .A1(n19726), .A2(n19797), .B1(n19725), .B2(n19736), .ZN(
        n19729) );
  AOI22_X1 U22761 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19742), .B1(
        n19727), .B2(n19740), .ZN(n19728) );
  OAI211_X1 U22762 ( .C1(n19730), .C2(n19735), .A(n19729), .B(n19728), .ZN(
        P2_U3165) );
  AOI22_X1 U22763 ( .A1(n19797), .A2(n19805), .B1(n19731), .B2(n19736), .ZN(
        n19734) );
  AOI22_X1 U22764 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19742), .B1(
        n19732), .B2(n19740), .ZN(n19733) );
  OAI211_X1 U22765 ( .C1(n19808), .C2(n19735), .A(n19734), .B(n19733), .ZN(
        P2_U3166) );
  AOI22_X1 U22766 ( .A1(n19739), .A2(n19738), .B1(n19737), .B2(n19736), .ZN(
        n19744) );
  AOI22_X1 U22767 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19742), .B1(
        n19741), .B2(n19740), .ZN(n19743) );
  OAI211_X1 U22768 ( .C1(n19745), .C2(n19819), .A(n19744), .B(n19743), .ZN(
        P2_U3167) );
  NAND2_X1 U22769 ( .A1(n19810), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19746) );
  NOR2_X1 U22770 ( .A1(n19747), .A2(n19746), .ZN(n19755) );
  INV_X1 U22771 ( .A(n19756), .ZN(n19748) );
  AOI21_X1 U22772 ( .B1(n19938), .B2(n19748), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19749) );
  OR2_X1 U22773 ( .A1(n19755), .A2(n19749), .ZN(n19812) );
  OAI22_X1 U22774 ( .A1(n19812), .A2(n19751), .B1(n19810), .B2(n19750), .ZN(
        n19752) );
  INV_X1 U22775 ( .A(n19752), .ZN(n19763) );
  NAND2_X1 U22776 ( .A1(n19754), .A2(n19753), .ZN(n19757) );
  AOI21_X1 U22777 ( .B1(n19757), .B2(n19756), .A(n19755), .ZN(n19759) );
  OAI211_X1 U22778 ( .C1(n19760), .C2(n19938), .A(n19759), .B(n19758), .ZN(
        n19816) );
  AOI22_X1 U22779 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19816), .B1(
        n19797), .B2(n19761), .ZN(n19762) );
  OAI211_X1 U22780 ( .C1(n19764), .C2(n19800), .A(n19763), .B(n19762), .ZN(
        P2_U3168) );
  OAI22_X1 U22781 ( .A1(n19812), .A2(n19766), .B1(n19810), .B2(n19765), .ZN(
        n19767) );
  INV_X1 U22782 ( .A(n19767), .ZN(n19770) );
  AOI22_X1 U22783 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19816), .B1(
        n19815), .B2(n19768), .ZN(n19769) );
  OAI211_X1 U22784 ( .C1(n19771), .C2(n19819), .A(n19770), .B(n19769), .ZN(
        P2_U3169) );
  OAI22_X1 U22785 ( .A1(n19812), .A2(n19773), .B1(n19810), .B2(n19772), .ZN(
        n19774) );
  INV_X1 U22786 ( .A(n19774), .ZN(n19777) );
  AOI22_X1 U22787 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19816), .B1(
        n19815), .B2(n19775), .ZN(n19776) );
  OAI211_X1 U22788 ( .C1(n19778), .C2(n19819), .A(n19777), .B(n19776), .ZN(
        P2_U3170) );
  OAI22_X1 U22789 ( .A1(n19812), .A2(n19780), .B1(n19810), .B2(n19779), .ZN(
        n19781) );
  INV_X1 U22790 ( .A(n19781), .ZN(n19784) );
  AOI22_X1 U22791 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19816), .B1(
        n19797), .B2(n19782), .ZN(n19783) );
  OAI211_X1 U22792 ( .C1(n19785), .C2(n19800), .A(n19784), .B(n19783), .ZN(
        P2_U3171) );
  OAI22_X1 U22793 ( .A1(n19812), .A2(n19787), .B1(n19810), .B2(n19786), .ZN(
        n19788) );
  INV_X1 U22794 ( .A(n19788), .ZN(n19791) );
  AOI22_X1 U22795 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19816), .B1(
        n19815), .B2(n19789), .ZN(n19790) );
  OAI211_X1 U22796 ( .C1(n19792), .C2(n19819), .A(n19791), .B(n19790), .ZN(
        P2_U3172) );
  OAI22_X1 U22797 ( .A1(n19812), .A2(n19794), .B1(n19810), .B2(n19793), .ZN(
        n19795) );
  INV_X1 U22798 ( .A(n19795), .ZN(n19799) );
  AOI22_X1 U22799 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19816), .B1(
        n19797), .B2(n19796), .ZN(n19798) );
  OAI211_X1 U22800 ( .C1(n19801), .C2(n19800), .A(n19799), .B(n19798), .ZN(
        P2_U3173) );
  OAI22_X1 U22801 ( .A1(n19812), .A2(n19803), .B1(n19810), .B2(n19802), .ZN(
        n19804) );
  INV_X1 U22802 ( .A(n19804), .ZN(n19807) );
  AOI22_X1 U22803 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19816), .B1(
        n19815), .B2(n19805), .ZN(n19806) );
  OAI211_X1 U22804 ( .C1(n19808), .C2(n19819), .A(n19807), .B(n19806), .ZN(
        P2_U3174) );
  OAI22_X1 U22805 ( .A1(n19812), .A2(n19811), .B1(n19810), .B2(n19809), .ZN(
        n19813) );
  INV_X1 U22806 ( .A(n19813), .ZN(n19818) );
  AOI22_X1 U22807 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19816), .B1(
        n19815), .B2(n19814), .ZN(n19817) );
  OAI211_X1 U22808 ( .C1(n19820), .C2(n19819), .A(n19818), .B(n19817), .ZN(
        P2_U3175) );
  AOI21_X1 U22809 ( .B1(n19823), .B2(n19822), .A(n19821), .ZN(n19833) );
  INV_X1 U22810 ( .A(n19824), .ZN(n19827) );
  NAND2_X1 U22811 ( .A1(n19851), .A2(n19825), .ZN(n19826) );
  NAND4_X1 U22812 ( .A1(n19829), .A2(n19828), .A3(n19827), .A4(n19826), .ZN(
        n19830) );
  OAI211_X1 U22813 ( .C1(n19833), .C2(n19832), .A(n19831), .B(n19830), .ZN(
        P2_U3177) );
  AND2_X1 U22814 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19834), .ZN(
        P2_U3179) );
  AND2_X1 U22815 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19834), .ZN(
        P2_U3180) );
  AND2_X1 U22816 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19834), .ZN(
        P2_U3181) );
  AND2_X1 U22817 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19834), .ZN(
        P2_U3182) );
  AND2_X1 U22818 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19834), .ZN(
        P2_U3183) );
  AND2_X1 U22819 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19834), .ZN(
        P2_U3184) );
  AND2_X1 U22820 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19834), .ZN(
        P2_U3185) );
  AND2_X1 U22821 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19834), .ZN(
        P2_U3186) );
  AND2_X1 U22822 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19834), .ZN(
        P2_U3187) );
  AND2_X1 U22823 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19834), .ZN(
        P2_U3188) );
  AND2_X1 U22824 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19834), .ZN(
        P2_U3189) );
  AND2_X1 U22825 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19834), .ZN(
        P2_U3190) );
  AND2_X1 U22826 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19834), .ZN(
        P2_U3191) );
  AND2_X1 U22827 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19834), .ZN(
        P2_U3192) );
  AND2_X1 U22828 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19834), .ZN(
        P2_U3193) );
  AND2_X1 U22829 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19834), .ZN(
        P2_U3194) );
  AND2_X1 U22830 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19834), .ZN(
        P2_U3195) );
  AND2_X1 U22831 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19834), .ZN(
        P2_U3196) );
  AND2_X1 U22832 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19834), .ZN(
        P2_U3197) );
  AND2_X1 U22833 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19834), .ZN(
        P2_U3198) );
  AND2_X1 U22834 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19834), .ZN(
        P2_U3199) );
  AND2_X1 U22835 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19834), .ZN(
        P2_U3200) );
  AND2_X1 U22836 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19834), .ZN(P2_U3201) );
  AND2_X1 U22837 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19834), .ZN(P2_U3202) );
  AND2_X1 U22838 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19834), .ZN(P2_U3203) );
  AND2_X1 U22839 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19834), .ZN(P2_U3204) );
  AND2_X1 U22840 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19834), .ZN(P2_U3205) );
  AND2_X1 U22841 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19834), .ZN(P2_U3206) );
  AND2_X1 U22842 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19834), .ZN(P2_U3207) );
  AND2_X1 U22843 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19834), .ZN(P2_U3208) );
  NOR2_X1 U22844 ( .A1(n19848), .A2(n19835), .ZN(n19844) );
  INV_X1 U22845 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19845) );
  NOR3_X1 U22846 ( .A1(n19844), .A2(n19845), .A3(n19837), .ZN(n19839) );
  OAI211_X1 U22847 ( .C1(HOLD), .C2(n19845), .A(n19836), .B(n19978), .ZN(
        n19838) );
  NAND3_X1 U22848 ( .A1(n19837), .A2(n19848), .A3(NA), .ZN(n19847) );
  OAI211_X1 U22849 ( .C1(P2_STATE_REG_2__SCAN_IN), .C2(n19839), .A(n19838), 
        .B(n19847), .ZN(P2_U3209) );
  AOI21_X1 U22850 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21232), .A(n19856), 
        .ZN(n19849) );
  NOR3_X1 U22851 ( .A1(n19849), .A2(n19845), .A3(n19837), .ZN(n19840) );
  NOR2_X1 U22852 ( .A1(n19840), .A2(n19844), .ZN(n19842) );
  OAI211_X1 U22853 ( .C1(n21232), .C2(n19843), .A(n19842), .B(n19841), .ZN(
        P2_U3210) );
  AOI22_X1 U22854 ( .A1(n19846), .A2(n19845), .B1(n19844), .B2(n21180), .ZN(
        n19855) );
  OAI21_X1 U22855 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .ZN(n19854) );
  INV_X1 U22856 ( .A(n19847), .ZN(n19853) );
  NOR2_X1 U22857 ( .A1(n19848), .A2(n19856), .ZN(n19850) );
  AOI21_X1 U22858 ( .B1(n19851), .B2(n19850), .A(n19849), .ZN(n19852) );
  OAI22_X1 U22859 ( .A1(n19855), .A2(n19854), .B1(n19853), .B2(n19852), .ZN(
        P2_U3211) );
  OAI222_X1 U22860 ( .A1(n19914), .A2(n19860), .B1(n19858), .B2(n19912), .C1(
        n19857), .C2(n19911), .ZN(P2_U3212) );
  OAI222_X1 U22861 ( .A1(n19911), .A2(n19860), .B1(n19859), .B2(n19912), .C1(
        n13272), .C2(n19914), .ZN(P2_U3213) );
  OAI222_X1 U22862 ( .A1(n19911), .A2(n13272), .B1(n19861), .B2(n19912), .C1(
        n19862), .C2(n19914), .ZN(P2_U3214) );
  OAI222_X1 U22863 ( .A1(n19914), .A2(n13404), .B1(n19863), .B2(n19912), .C1(
        n19862), .C2(n19911), .ZN(P2_U3215) );
  OAI222_X1 U22864 ( .A1(n19914), .A2(n19865), .B1(n19864), .B2(n19912), .C1(
        n13404), .C2(n19911), .ZN(P2_U3216) );
  OAI222_X1 U22865 ( .A1(n19914), .A2(n19867), .B1(n19866), .B2(n19912), .C1(
        n19865), .C2(n19911), .ZN(P2_U3217) );
  INV_X1 U22866 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n19870) );
  OAI222_X1 U22867 ( .A1(n19914), .A2(n19870), .B1(n19869), .B2(n19868), .C1(
        n19867), .C2(n19911), .ZN(P2_U3218) );
  OAI222_X1 U22868 ( .A1(n19914), .A2(n14799), .B1(n19871), .B2(n19912), .C1(
        n19870), .C2(n19911), .ZN(P2_U3219) );
  OAI222_X1 U22869 ( .A1(n19914), .A2(n19873), .B1(n19872), .B2(n19868), .C1(
        n14799), .C2(n19911), .ZN(P2_U3220) );
  INV_X1 U22870 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n19875) );
  OAI222_X1 U22871 ( .A1(n19914), .A2(n19875), .B1(n19874), .B2(n19868), .C1(
        n19873), .C2(n19911), .ZN(P2_U3221) );
  OAI222_X1 U22872 ( .A1(n19914), .A2(n19877), .B1(n19876), .B2(n19868), .C1(
        n19875), .C2(n19911), .ZN(P2_U3222) );
  INV_X1 U22873 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n19879) );
  OAI222_X1 U22874 ( .A1(n19914), .A2(n19879), .B1(n19878), .B2(n19868), .C1(
        n19877), .C2(n19911), .ZN(P2_U3223) );
  OAI222_X1 U22875 ( .A1(n19914), .A2(n19881), .B1(n19880), .B2(n19868), .C1(
        n19879), .C2(n19911), .ZN(P2_U3224) );
  OAI222_X1 U22876 ( .A1(n19914), .A2(n19883), .B1(n19882), .B2(n19868), .C1(
        n19881), .C2(n19911), .ZN(P2_U3225) );
  OAI222_X1 U22877 ( .A1(n19914), .A2(n19885), .B1(n19884), .B2(n19868), .C1(
        n19883), .C2(n19911), .ZN(P2_U3226) );
  OAI222_X1 U22878 ( .A1(n19914), .A2(n19887), .B1(n19886), .B2(n19868), .C1(
        n19885), .C2(n19911), .ZN(P2_U3227) );
  OAI222_X1 U22879 ( .A1(n19914), .A2(n19889), .B1(n19888), .B2(n19868), .C1(
        n19887), .C2(n19911), .ZN(P2_U3228) );
  OAI222_X1 U22880 ( .A1(n19914), .A2(n19891), .B1(n19890), .B2(n19868), .C1(
        n19889), .C2(n19911), .ZN(P2_U3229) );
  OAI222_X1 U22881 ( .A1(n19914), .A2(n19893), .B1(n19892), .B2(n19868), .C1(
        n19891), .C2(n19911), .ZN(P2_U3230) );
  OAI222_X1 U22882 ( .A1(n19914), .A2(n19895), .B1(n19894), .B2(n19868), .C1(
        n19893), .C2(n19911), .ZN(P2_U3231) );
  OAI222_X1 U22883 ( .A1(n19914), .A2(n19897), .B1(n19896), .B2(n19868), .C1(
        n19895), .C2(n19911), .ZN(P2_U3232) );
  OAI222_X1 U22884 ( .A1(n19914), .A2(n19899), .B1(n19898), .B2(n19868), .C1(
        n19897), .C2(n19911), .ZN(P2_U3233) );
  OAI222_X1 U22885 ( .A1(n19914), .A2(n19901), .B1(n19900), .B2(n19912), .C1(
        n19899), .C2(n19911), .ZN(P2_U3234) );
  OAI222_X1 U22886 ( .A1(n19914), .A2(n19903), .B1(n19902), .B2(n19912), .C1(
        n19901), .C2(n19911), .ZN(P2_U3235) );
  OAI222_X1 U22887 ( .A1(n19914), .A2(n15049), .B1(n19904), .B2(n19912), .C1(
        n19903), .C2(n19911), .ZN(P2_U3236) );
  OAI222_X1 U22888 ( .A1(n19914), .A2(n19907), .B1(n19905), .B2(n19912), .C1(
        n15049), .C2(n19911), .ZN(P2_U3237) );
  OAI222_X1 U22889 ( .A1(n19911), .A2(n19907), .B1(n19906), .B2(n19912), .C1(
        n16197), .C2(n19914), .ZN(P2_U3238) );
  OAI222_X1 U22890 ( .A1(n19914), .A2(n19909), .B1(n19908), .B2(n19912), .C1(
        n16197), .C2(n19911), .ZN(P2_U3239) );
  OAI222_X1 U22891 ( .A1(n19914), .A2(n15003), .B1(n19910), .B2(n19912), .C1(
        n19909), .C2(n19911), .ZN(P2_U3240) );
  INV_X1 U22892 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19913) );
  OAI222_X1 U22893 ( .A1(n19914), .A2(n14759), .B1(n19913), .B2(n19912), .C1(
        n15003), .C2(n19911), .ZN(P2_U3241) );
  OAI22_X1 U22894 ( .A1(n19978), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n19912), .ZN(n19915) );
  INV_X1 U22895 ( .A(n19915), .ZN(P2_U3585) );
  MUX2_X1 U22896 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n19978), .Z(P2_U3586) );
  OAI22_X1 U22897 ( .A1(n19978), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n19912), .ZN(n19916) );
  INV_X1 U22898 ( .A(n19916), .ZN(P2_U3587) );
  OAI22_X1 U22899 ( .A1(n19978), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n19912), .ZN(n19917) );
  INV_X1 U22900 ( .A(n19917), .ZN(P2_U3588) );
  OAI21_X1 U22901 ( .B1(n19921), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19919), 
        .ZN(n19918) );
  INV_X1 U22902 ( .A(n19918), .ZN(P2_U3591) );
  OAI21_X1 U22903 ( .B1(n19921), .B2(n19920), .A(n19919), .ZN(P2_U3592) );
  AND2_X1 U22904 ( .A1(n19923), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19950) );
  NAND2_X1 U22905 ( .A1(n19922), .A2(n19950), .ZN(n19940) );
  OAI21_X1 U22906 ( .B1(n19949), .B2(n19924), .A(n19923), .ZN(n19926) );
  AND2_X1 U22907 ( .A1(n19926), .A2(n19925), .ZN(n19937) );
  NAND2_X1 U22908 ( .A1(n19940), .A2(n19937), .ZN(n19929) );
  AOI22_X1 U22909 ( .A1(n19929), .A2(n19928), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n19927), .ZN(n19930) );
  OAI21_X1 U22910 ( .B1(n19932), .B2(n19931), .A(n19930), .ZN(n19933) );
  INV_X1 U22911 ( .A(n19933), .ZN(n19934) );
  AOI22_X1 U22912 ( .A1(n19965), .A2(n19935), .B1(n19934), .B2(n19962), .ZN(
        P2_U3602) );
  INV_X1 U22913 ( .A(n19936), .ZN(n19944) );
  INV_X1 U22914 ( .A(n19937), .ZN(n19943) );
  NOR2_X1 U22915 ( .A1(n19939), .A2(n19938), .ZN(n19942) );
  INV_X1 U22916 ( .A(n19940), .ZN(n19941) );
  AOI211_X1 U22917 ( .C1(n19944), .C2(n19943), .A(n19942), .B(n19941), .ZN(
        n19945) );
  AOI22_X1 U22918 ( .A1(n19965), .A2(n19946), .B1(n19945), .B2(n19962), .ZN(
        P2_U3603) );
  INV_X1 U22919 ( .A(n19947), .ZN(n19957) );
  AND2_X1 U22920 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19948) );
  NOR2_X1 U22921 ( .A1(n19957), .A2(n19948), .ZN(n19951) );
  MUX2_X1 U22922 ( .A(n19951), .B(n19950), .S(n19949), .Z(n19952) );
  AOI21_X1 U22923 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19953), .A(n19952), 
        .ZN(n19954) );
  AOI22_X1 U22924 ( .A1(n19965), .A2(n19955), .B1(n19954), .B2(n19962), .ZN(
        P2_U3604) );
  OAI21_X1 U22925 ( .B1(n19958), .B2(n19957), .A(n19956), .ZN(n19959) );
  AOI21_X1 U22926 ( .B1(n19961), .B2(n19960), .A(n19959), .ZN(n19963) );
  AOI22_X1 U22927 ( .A1(n19965), .A2(n19964), .B1(n19963), .B2(n19962), .ZN(
        P2_U3605) );
  INV_X1 U22928 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19966) );
  AOI22_X1 U22929 ( .A1(n19868), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19966), 
        .B2(n19978), .ZN(P2_U3608) );
  INV_X1 U22930 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n19977) );
  INV_X1 U22931 ( .A(n19967), .ZN(n19971) );
  INV_X1 U22932 ( .A(n19968), .ZN(n19970) );
  AOI22_X1 U22933 ( .A1(n19972), .A2(n19971), .B1(n19970), .B2(n19969), .ZN(
        n19975) );
  NOR2_X1 U22934 ( .A1(n19973), .A2(n19976), .ZN(n19974) );
  AOI22_X1 U22935 ( .A1(n19977), .A2(n19976), .B1(n19975), .B2(n19974), .ZN(
        P2_U3609) );
  OAI22_X1 U22936 ( .A1(n19978), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n19912), .ZN(n19979) );
  INV_X1 U22937 ( .A(n19979), .ZN(P2_U3611) );
  NOR2_X2 U22938 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20834), .ZN(n20909) );
  INV_X1 U22939 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n21199) );
  NAND2_X1 U22940 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20843), .ZN(n19980) );
  AOI21_X1 U22941 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n19980), .A(n20909), 
        .ZN(n20888) );
  OAI21_X1 U22942 ( .B1(n20909), .B2(n21199), .A(n20829), .ZN(P1_U2802) );
  INV_X1 U22943 ( .A(n19981), .ZN(n19983) );
  OAI21_X1 U22944 ( .B1(n19983), .B2(n19982), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19984) );
  OAI21_X1 U22945 ( .B1(n19985), .B2(n20902), .A(n19984), .ZN(P1_U2803) );
  INV_X1 U22946 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n20986) );
  NOR2_X1 U22947 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19987) );
  NOR2_X1 U22948 ( .A1(n20909), .A2(n19987), .ZN(n19986) );
  AOI22_X1 U22949 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(n20909), .B1(n20986), 
        .B2(n19986), .ZN(P1_U2804) );
  OAI21_X1 U22950 ( .B1(BS16), .B2(n19987), .A(n20888), .ZN(n20886) );
  OAI21_X1 U22951 ( .B1(n20888), .B2(n21280), .A(n20886), .ZN(P1_U2805) );
  OAI21_X1 U22952 ( .B1(n19989), .B2(n21022), .A(n19988), .ZN(P1_U2806) );
  NOR4_X1 U22953 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19993) );
  NOR4_X1 U22954 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19992) );
  NOR4_X1 U22955 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19991) );
  NOR4_X1 U22956 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19990) );
  NAND4_X1 U22957 ( .A1(n19993), .A2(n19992), .A3(n19991), .A4(n19990), .ZN(
        n19999) );
  NOR4_X1 U22958 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19997) );
  AOI211_X1 U22959 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19996) );
  NOR4_X1 U22960 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19995) );
  NOR4_X1 U22961 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19994) );
  NAND4_X1 U22962 ( .A1(n19997), .A2(n19996), .A3(n19995), .A4(n19994), .ZN(
        n19998) );
  NOR2_X1 U22963 ( .A1(n19999), .A2(n19998), .ZN(n20893) );
  INV_X1 U22964 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20962) );
  NOR3_X1 U22965 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20001) );
  OAI21_X1 U22966 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20001), .A(n20893), .ZN(
        n20000) );
  OAI21_X1 U22967 ( .B1(n20893), .B2(n20962), .A(n20000), .ZN(P1_U2807) );
  INV_X1 U22968 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20887) );
  AOI21_X1 U22969 ( .B1(n20889), .B2(n20887), .A(n20001), .ZN(n20002) );
  INV_X1 U22970 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21242) );
  INV_X1 U22971 ( .A(n20893), .ZN(n20895) );
  AOI22_X1 U22972 ( .A1(n20893), .A2(n20002), .B1(n21242), .B2(n20895), .ZN(
        P1_U2808) );
  NOR4_X1 U22973 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n21208), .A3(n20003), .A4(
        n20038), .ZN(n20004) );
  AOI21_X1 U22974 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(n20005), .A(n20004), .ZN(
        n20013) );
  INV_X1 U22975 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n20092) );
  OAI22_X1 U22976 ( .A1(n20006), .A2(n20060), .B1(n20092), .B2(n20064), .ZN(
        n20007) );
  AOI211_X1 U22977 ( .C1(n20077), .C2(n20008), .A(n20048), .B(n20007), .ZN(
        n20012) );
  INV_X1 U22978 ( .A(n20089), .ZN(n20010) );
  AOI22_X1 U22979 ( .A1(n20010), .A2(n20031), .B1(n20079), .B2(n20009), .ZN(
        n20011) );
  NAND3_X1 U22980 ( .A1(n20013), .A2(n20012), .A3(n20011), .ZN(P1_U2831) );
  AOI22_X1 U22981 ( .A1(P1_EBX_REG_7__SCAN_IN), .A2(n20075), .B1(n20077), .B2(
        n20093), .ZN(n20017) );
  INV_X1 U22982 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21272) );
  NOR2_X1 U22983 ( .A1(n21235), .A2(n21272), .ZN(n20022) );
  INV_X1 U22984 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20015) );
  INV_X1 U22985 ( .A(n20038), .ZN(n20014) );
  NAND3_X1 U22986 ( .A1(n20022), .A2(n20015), .A3(n20014), .ZN(n20016) );
  NAND2_X1 U22987 ( .A1(n20017), .A2(n20016), .ZN(n20018) );
  AOI211_X1 U22988 ( .C1(n20080), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n20048), .B(n20018), .ZN(n20024) );
  AOI21_X1 U22989 ( .B1(n20069), .B2(n20020), .A(n20019), .ZN(n20054) );
  OAI21_X1 U22990 ( .B1(n20022), .B2(n20021), .A(n20054), .ZN(n20032) );
  AOI22_X1 U22991 ( .A1(n20032), .A2(P1_REIP_REG_7__SCAN_IN), .B1(n20094), 
        .B2(n20031), .ZN(n20023) );
  OAI211_X1 U22992 ( .C1(n20025), .C2(n20043), .A(n20024), .B(n20023), .ZN(
        P1_U2833) );
  NOR2_X1 U22993 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20038), .ZN(n20026) );
  AOI22_X1 U22994 ( .A1(P1_EBX_REG_6__SCAN_IN), .A2(n20075), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n20026), .ZN(n20027) );
  OAI21_X1 U22995 ( .B1(n20073), .B2(n20028), .A(n20027), .ZN(n20029) );
  AOI211_X1 U22996 ( .C1(n20080), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n20048), .B(n20029), .ZN(n20034) );
  AOI22_X1 U22997 ( .A1(n20032), .A2(P1_REIP_REG_6__SCAN_IN), .B1(n20031), 
        .B2(n20030), .ZN(n20033) );
  OAI211_X1 U22998 ( .C1(n20035), .C2(n20043), .A(n20034), .B(n20033), .ZN(
        P1_U2834) );
  OAI22_X1 U22999 ( .A1(n20054), .A2(n21272), .B1(n20036), .B2(n20060), .ZN(
        n20037) );
  AOI211_X1 U23000 ( .C1(n20077), .C2(n20096), .A(n20048), .B(n20037), .ZN(
        n20042) );
  INV_X1 U23001 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n21265) );
  OAI22_X1 U23002 ( .A1(n20038), .A2(P1_REIP_REG_5__SCAN_IN), .B1(n21265), 
        .B2(n20064), .ZN(n20039) );
  AOI21_X1 U23003 ( .B1(n20099), .B2(n20040), .A(n20039), .ZN(n20041) );
  OAI211_X1 U23004 ( .C1(n20044), .C2(n20043), .A(n20042), .B(n20041), .ZN(
        P1_U2835) );
  OAI22_X1 U23005 ( .A1(n20073), .A2(n20172), .B1(n20046), .B2(n20045), .ZN(
        n20047) );
  AOI211_X1 U23006 ( .C1(n20080), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20048), .B(n20047), .ZN(n20057) );
  NOR3_X1 U23007 ( .A1(n21230), .A2(n20889), .A3(n21165), .ZN(n20049) );
  AOI21_X1 U23008 ( .B1(n20069), .B2(n20049), .A(P1_REIP_REG_4__SCAN_IN), .ZN(
        n20053) );
  INV_X1 U23009 ( .A(n20163), .ZN(n20050) );
  NAND2_X1 U23010 ( .A1(n20079), .A2(n20050), .ZN(n20052) );
  OR2_X1 U23011 ( .A1(n20156), .A2(n20087), .ZN(n20051) );
  OAI211_X1 U23012 ( .C1(n20054), .C2(n20053), .A(n20052), .B(n20051), .ZN(
        n20055) );
  INV_X1 U23013 ( .A(n20055), .ZN(n20056) );
  OAI211_X1 U23014 ( .C1(n20058), .C2(n20064), .A(n20057), .B(n20056), .ZN(
        P1_U2836) );
  OAI22_X1 U23015 ( .A1(n20060), .A2(n20062), .B1(n20889), .B2(n20059), .ZN(
        n20061) );
  AOI21_X1 U23016 ( .B1(n20079), .B2(n20062), .A(n20061), .ZN(n20063) );
  OAI21_X1 U23017 ( .B1(n20065), .B2(n20064), .A(n20063), .ZN(n20068) );
  NOR2_X1 U23018 ( .A1(n20066), .A2(n20087), .ZN(n20067) );
  AOI211_X1 U23019 ( .C1(n20078), .C2(n20726), .A(n20068), .B(n20067), .ZN(
        n20071) );
  NAND2_X1 U23020 ( .A1(n20069), .A2(n20889), .ZN(n20070) );
  OAI211_X1 U23021 ( .C1(n20073), .C2(n20072), .A(n20071), .B(n20070), .ZN(
        P1_U2839) );
  AOI22_X1 U23022 ( .A1(P1_EBX_REG_0__SCAN_IN), .A2(n20075), .B1(
        P1_REIP_REG_0__SCAN_IN), .B2(n20074), .ZN(n20085) );
  NAND2_X1 U23023 ( .A1(n20077), .A2(n20076), .ZN(n20083) );
  NAND2_X1 U23024 ( .A1(n20078), .A2(n11839), .ZN(n20082) );
  OAI21_X1 U23025 ( .B1(n20080), .B2(n20079), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n20081) );
  AND3_X1 U23026 ( .A1(n20083), .A2(n20082), .A3(n20081), .ZN(n20084) );
  OAI211_X1 U23027 ( .C1(n20087), .C2(n20086), .A(n20085), .B(n20084), .ZN(
        P1_U2840) );
  OAI22_X1 U23028 ( .A1(n20089), .A2(n14326), .B1(n14316), .B2(n20088), .ZN(
        n20090) );
  INV_X1 U23029 ( .A(n20090), .ZN(n20091) );
  OAI21_X1 U23030 ( .B1(n20101), .B2(n20092), .A(n20091), .ZN(P1_U2863) );
  AOI22_X1 U23031 ( .A1(n20094), .A2(n20098), .B1(n20097), .B2(n20093), .ZN(
        n20095) );
  OAI21_X1 U23032 ( .B1(n20101), .B2(n21201), .A(n20095), .ZN(P1_U2865) );
  AOI22_X1 U23033 ( .A1(n20099), .A2(n20098), .B1(n20097), .B2(n20096), .ZN(
        n20100) );
  OAI21_X1 U23034 ( .B1(n20101), .B2(n21265), .A(n20100), .ZN(P1_U2867) );
  AOI22_X1 U23035 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20105), .B1(n15908), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20102) );
  OAI21_X1 U23036 ( .B1(n20104), .B2(n20103), .A(n20102), .ZN(P1_U2921) );
  INV_X1 U23037 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20107) );
  AOI22_X1 U23038 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20106) );
  OAI21_X1 U23039 ( .B1(n20107), .B2(n20134), .A(n20106), .ZN(P1_U2922) );
  INV_X1 U23040 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20109) );
  AOI22_X1 U23041 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20108) );
  OAI21_X1 U23042 ( .B1(n20109), .B2(n20134), .A(n20108), .ZN(P1_U2923) );
  INV_X1 U23043 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20111) );
  AOI22_X1 U23044 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20110) );
  OAI21_X1 U23045 ( .B1(n20111), .B2(n20134), .A(n20110), .ZN(P1_U2924) );
  INV_X1 U23046 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20113) );
  AOI22_X1 U23047 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20112) );
  OAI21_X1 U23048 ( .B1(n20113), .B2(n20134), .A(n20112), .ZN(P1_U2925) );
  INV_X1 U23049 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20115) );
  AOI22_X1 U23050 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20114) );
  OAI21_X1 U23051 ( .B1(n20115), .B2(n20134), .A(n20114), .ZN(P1_U2926) );
  INV_X1 U23052 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20117) );
  AOI22_X1 U23053 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20116) );
  OAI21_X1 U23054 ( .B1(n20117), .B2(n20134), .A(n20116), .ZN(P1_U2927) );
  AOI22_X1 U23055 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20118) );
  OAI21_X1 U23056 ( .B1(n20119), .B2(n20134), .A(n20118), .ZN(P1_U2928) );
  AOI22_X1 U23057 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20120) );
  OAI21_X1 U23058 ( .B1(n13292), .B2(n20134), .A(n20120), .ZN(P1_U2929) );
  AOI22_X1 U23059 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20121) );
  OAI21_X1 U23060 ( .B1(n20122), .B2(n20134), .A(n20121), .ZN(P1_U2930) );
  AOI22_X1 U23061 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20123) );
  OAI21_X1 U23062 ( .B1(n13137), .B2(n20134), .A(n20123), .ZN(P1_U2931) );
  AOI22_X1 U23063 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20124) );
  OAI21_X1 U23064 ( .B1(n20125), .B2(n20134), .A(n20124), .ZN(P1_U2932) );
  AOI22_X1 U23065 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20126) );
  OAI21_X1 U23066 ( .B1(n20127), .B2(n20134), .A(n20126), .ZN(P1_U2933) );
  AOI22_X1 U23067 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20128) );
  OAI21_X1 U23068 ( .B1(n20129), .B2(n20134), .A(n20128), .ZN(P1_U2934) );
  AOI22_X1 U23069 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20130) );
  OAI21_X1 U23070 ( .B1(n20131), .B2(n20134), .A(n20130), .ZN(P1_U2935) );
  AOI22_X1 U23071 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20132), .B1(n15908), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20133) );
  OAI21_X1 U23072 ( .B1(n20135), .B2(n20134), .A(n20133), .ZN(P1_U2936) );
  AOI22_X1 U23073 ( .A1(n20147), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20146), .ZN(n20137) );
  NAND2_X1 U23074 ( .A1(n20137), .A2(n20136), .ZN(P1_U2961) );
  AOI22_X1 U23075 ( .A1(n20147), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n20146), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n20139) );
  NAND2_X1 U23076 ( .A1(n20139), .A2(n20138), .ZN(P1_U2962) );
  AOI22_X1 U23077 ( .A1(n20147), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20146), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n20141) );
  NAND2_X1 U23078 ( .A1(n20141), .A2(n20140), .ZN(P1_U2963) );
  AOI22_X1 U23079 ( .A1(n20147), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n20146), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20143) );
  NAND2_X1 U23080 ( .A1(n20143), .A2(n20142), .ZN(P1_U2964) );
  AOI22_X1 U23081 ( .A1(n20147), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20146), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20145) );
  NAND2_X1 U23082 ( .A1(n20145), .A2(n20144), .ZN(P1_U2965) );
  AOI22_X1 U23083 ( .A1(n20147), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n20146), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20149) );
  NAND2_X1 U23084 ( .A1(n20149), .A2(n20148), .ZN(P1_U2966) );
  AOI22_X1 U23085 ( .A1(n20151), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20150), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20162) );
  OR2_X1 U23086 ( .A1(n20153), .A2(n20152), .ZN(n20154) );
  NAND2_X1 U23087 ( .A1(n20155), .A2(n20154), .ZN(n20170) );
  INV_X1 U23088 ( .A(n20170), .ZN(n20160) );
  INV_X1 U23089 ( .A(n20156), .ZN(n20157) );
  AOI22_X1 U23090 ( .A1(n20160), .A2(n20159), .B1(n20158), .B2(n20157), .ZN(
        n20161) );
  OAI211_X1 U23091 ( .C1(n20164), .C2(n20163), .A(n20162), .B(n20161), .ZN(
        P1_U2995) );
  NOR2_X1 U23092 ( .A1(n20203), .A2(n20217), .ZN(n20166) );
  OAI21_X1 U23093 ( .B1(n20167), .B2(n20166), .A(n20165), .ZN(n20191) );
  AOI21_X1 U23094 ( .B1(n20193), .B2(n20168), .A(n20191), .ZN(n20188) );
  AOI211_X1 U23095 ( .C1(n20177), .C2(n20187), .A(n20169), .B(n20183), .ZN(
        n20175) );
  NOR2_X1 U23096 ( .A1(n20170), .A2(n20196), .ZN(n20174) );
  INV_X1 U23097 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20846) );
  OAI22_X1 U23098 ( .A1(n20172), .A2(n20171), .B1(n20846), .B2(n20207), .ZN(
        n20173) );
  NOR3_X1 U23099 ( .A1(n20175), .A2(n20174), .A3(n20173), .ZN(n20176) );
  OAI21_X1 U23100 ( .B1(n20188), .B2(n20177), .A(n20176), .ZN(P1_U3027) );
  INV_X1 U23101 ( .A(n20178), .ZN(n20181) );
  INV_X1 U23102 ( .A(n20179), .ZN(n20180) );
  AOI21_X1 U23103 ( .B1(n20181), .B2(n20214), .A(n20180), .ZN(n20186) );
  OAI22_X1 U23104 ( .A1(n20183), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        n20182), .B2(n20196), .ZN(n20184) );
  INV_X1 U23105 ( .A(n20184), .ZN(n20185) );
  OAI211_X1 U23106 ( .C1(n20188), .C2(n20187), .A(n20186), .B(n20185), .ZN(
        P1_U3028) );
  INV_X1 U23107 ( .A(n20189), .ZN(n20204) );
  NOR2_X1 U23108 ( .A1(n20190), .A2(n20217), .ZN(n20192) );
  AOI21_X1 U23109 ( .B1(n20193), .B2(n20192), .A(n20191), .ZN(n20202) );
  OAI22_X1 U23110 ( .A1(n20195), .A2(n20194), .B1(n21165), .B2(n20207), .ZN(
        n20199) );
  NOR2_X1 U23111 ( .A1(n20197), .A2(n20196), .ZN(n20198) );
  AOI211_X1 U23112 ( .C1(n20214), .C2(n20200), .A(n20199), .B(n20198), .ZN(
        n20201) );
  OAI221_X1 U23113 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20204), .C1(
        n20203), .C2(n20202), .A(n20201), .ZN(P1_U3029) );
  NAND2_X1 U23114 ( .A1(n20206), .A2(n20205), .ZN(n20218) );
  NOR2_X1 U23115 ( .A1(n20207), .A2(n20889), .ZN(n20212) );
  AND3_X1 U23116 ( .A1(n20210), .A2(n20209), .A3(n20208), .ZN(n20211) );
  AOI211_X1 U23117 ( .C1(n20214), .C2(n20213), .A(n20212), .B(n20211), .ZN(
        n20215) );
  OAI221_X1 U23118 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20218), .C1(
        n20217), .C2(n20216), .A(n20215), .ZN(P1_U3030) );
  NOR2_X1 U23119 ( .A1(n12321), .A2(n20219), .ZN(P1_U3032) );
  NAND2_X1 U23120 ( .A1(n20559), .A2(n20501), .ZN(n20391) );
  INV_X1 U23121 ( .A(n20233), .ZN(n20220) );
  NOR2_X1 U23122 ( .A1(n20220), .A2(n20898), .ZN(n20633) );
  INV_X1 U23123 ( .A(n20563), .ZN(n20327) );
  NOR3_X1 U23124 ( .A1(n20319), .A2(n20820), .A3(n12580), .ZN(n20223) );
  INV_X1 U23125 ( .A(n20628), .ZN(n20222) );
  NOR2_X1 U23126 ( .A1(n20223), .A2(n20222), .ZN(n20235) );
  INV_X1 U23127 ( .A(n20631), .ZN(n20224) );
  OR2_X1 U23128 ( .A1(n20500), .A2(n20224), .ZN(n20359) );
  OR2_X1 U23129 ( .A1(n20359), .A2(n20726), .ZN(n20234) );
  INV_X1 U23130 ( .A(n20234), .ZN(n20225) );
  NOR3_X1 U23131 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20302) );
  INV_X1 U23132 ( .A(n20302), .ZN(n20299) );
  NOR2_X1 U23133 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20299), .ZN(
        n20288) );
  OAI22_X1 U23134 ( .A1(n20235), .A2(n20225), .B1(n20288), .B2(n20641), .ZN(
        n20226) );
  INV_X1 U23135 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20239) );
  INV_X1 U23136 ( .A(DATAI_24_), .ZN(n21210) );
  OAI22_X2 U23137 ( .A1(n20229), .A2(n20291), .B1(n21210), .B2(n20290), .ZN(
        n20773) );
  NOR2_X2 U23138 ( .A1(n20287), .A2(n20231), .ZN(n20764) );
  AOI22_X1 U23139 ( .A1(n20820), .A2(n20773), .B1(n20764), .B2(n20288), .ZN(
        n20238) );
  NOR2_X1 U23140 ( .A1(n20233), .A2(n20898), .ZN(n20561) );
  INV_X1 U23141 ( .A(n20561), .ZN(n20503) );
  OAI22_X1 U23142 ( .A1(n20235), .A2(n20234), .B1(n20503), .B2(n20391), .ZN(
        n20292) );
  INV_X1 U23143 ( .A(DATAI_16_), .ZN(n21001) );
  OAI22_X1 U23144 ( .A1(n20236), .A2(n20291), .B1(n21001), .B2(n20290), .ZN(
        n20693) );
  AOI22_X1 U23145 ( .A1(n20765), .A2(n20292), .B1(n20319), .B2(n20693), .ZN(
        n20237) );
  OAI211_X1 U23146 ( .C1(n20296), .C2(n20239), .A(n20238), .B(n20237), .ZN(
        P1_U3033) );
  INV_X1 U23147 ( .A(DATAI_25_), .ZN(n21186) );
  OAI22_X2 U23148 ( .A1(n20240), .A2(n20291), .B1(n21186), .B2(n20290), .ZN(
        n20779) );
  NOR2_X2 U23149 ( .A1(n20287), .A2(n20241), .ZN(n20777) );
  AOI22_X1 U23150 ( .A1(n20820), .A2(n20779), .B1(n20777), .B2(n20288), .ZN(
        n20245) );
  INV_X1 U23151 ( .A(DATAI_17_), .ZN(n20945) );
  OAI22_X1 U23152 ( .A1(n20243), .A2(n20291), .B1(n20945), .B2(n20290), .ZN(
        n20697) );
  AOI22_X1 U23153 ( .A1(n20778), .A2(n20292), .B1(n20319), .B2(n20697), .ZN(
        n20244) );
  OAI211_X1 U23154 ( .C1(n20296), .C2(n20246), .A(n20245), .B(n20244), .ZN(
        P1_U3034) );
  INV_X1 U23155 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n20254) );
  INV_X1 U23156 ( .A(DATAI_26_), .ZN(n21167) );
  OAI22_X2 U23157 ( .A1(n20247), .A2(n20291), .B1(n21167), .B2(n20290), .ZN(
        n20735) );
  NOR2_X2 U23158 ( .A1(n20287), .A2(n20248), .ZN(n20783) );
  AOI22_X1 U23159 ( .A1(n20820), .A2(n20735), .B1(n20783), .B2(n20288), .ZN(
        n20253) );
  INV_X1 U23160 ( .A(DATAI_18_), .ZN(n20250) );
  OAI22_X1 U23161 ( .A1(n20251), .A2(n20291), .B1(n20250), .B2(n20290), .ZN(
        n20785) );
  AOI22_X1 U23162 ( .A1(n20784), .A2(n20292), .B1(n20319), .B2(n20785), .ZN(
        n20252) );
  OAI211_X1 U23163 ( .C1(n20296), .C2(n20254), .A(n20253), .B(n20252), .ZN(
        P1_U3035) );
  INV_X1 U23164 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n20262) );
  INV_X1 U23165 ( .A(DATAI_27_), .ZN(n21104) );
  NOR2_X2 U23166 ( .A1(n20287), .A2(n20256), .ZN(n20789) );
  AOI22_X1 U23167 ( .A1(n20820), .A2(n20739), .B1(n20789), .B2(n20288), .ZN(
        n20261) );
  INV_X1 U23168 ( .A(DATAI_19_), .ZN(n20259) );
  OAI22_X1 U23169 ( .A1(n20259), .A2(n20290), .B1(n20258), .B2(n20291), .ZN(
        n20791) );
  AOI22_X1 U23170 ( .A1(n20790), .A2(n20292), .B1(n20319), .B2(n20791), .ZN(
        n20260) );
  OAI211_X1 U23171 ( .C1(n20296), .C2(n20262), .A(n20261), .B(n20260), .ZN(
        P1_U3036) );
  INV_X1 U23172 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n20269) );
  INV_X1 U23173 ( .A(DATAI_28_), .ZN(n21274) );
  NOR2_X2 U23174 ( .A1(n20287), .A2(n20263), .ZN(n20795) );
  AOI22_X1 U23175 ( .A1(n20820), .A2(n20743), .B1(n20795), .B2(n20288), .ZN(
        n20268) );
  INV_X1 U23176 ( .A(DATAI_20_), .ZN(n20265) );
  OAI22_X1 U23177 ( .A1(n20266), .A2(n20291), .B1(n20265), .B2(n20290), .ZN(
        n20797) );
  AOI22_X1 U23178 ( .A1(n20796), .A2(n20292), .B1(n20319), .B2(n20797), .ZN(
        n20267) );
  OAI211_X1 U23179 ( .C1(n20296), .C2(n20269), .A(n20268), .B(n20267), .ZN(
        P1_U3037) );
  INV_X1 U23180 ( .A(DATAI_29_), .ZN(n21196) );
  OAI22_X2 U23181 ( .A1(n20270), .A2(n20291), .B1(n21196), .B2(n20290), .ZN(
        n20803) );
  NOR2_X2 U23182 ( .A1(n20287), .A2(n20271), .ZN(n20801) );
  AOI22_X1 U23183 ( .A1(n20820), .A2(n20803), .B1(n20801), .B2(n20288), .ZN(
        n20275) );
  OAI22_X1 U23184 ( .A1(n20273), .A2(n20291), .B1(n14363), .B2(n20290), .ZN(
        n20707) );
  AOI22_X1 U23185 ( .A1(n20802), .A2(n20292), .B1(n20319), .B2(n20707), .ZN(
        n20274) );
  OAI211_X1 U23186 ( .C1(n20296), .C2(n20276), .A(n20275), .B(n20274), .ZN(
        P1_U3038) );
  INV_X1 U23187 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n20283) );
  INV_X1 U23188 ( .A(DATAI_30_), .ZN(n21251) );
  NOR2_X2 U23189 ( .A1(n20287), .A2(n20278), .ZN(n20809) );
  AOI22_X1 U23190 ( .A1(n20820), .A2(n20749), .B1(n20809), .B2(n20288), .ZN(
        n20282) );
  INV_X1 U23191 ( .A(DATAI_22_), .ZN(n21207) );
  OAI22_X1 U23192 ( .A1(n20280), .A2(n20291), .B1(n21207), .B2(n20290), .ZN(
        n20811) );
  AOI22_X1 U23193 ( .A1(n20810), .A2(n20292), .B1(n20319), .B2(n20811), .ZN(
        n20281) );
  OAI211_X1 U23194 ( .C1(n20296), .C2(n20283), .A(n20282), .B(n20281), .ZN(
        P1_U3039) );
  INV_X1 U23195 ( .A(DATAI_31_), .ZN(n20285) );
  NOR2_X2 U23196 ( .A1(n20287), .A2(n20286), .ZN(n20816) );
  AOI22_X1 U23197 ( .A1(n20820), .A2(n20755), .B1(n20816), .B2(n20288), .ZN(
        n20294) );
  INV_X1 U23198 ( .A(DATAI_23_), .ZN(n21003) );
  OAI22_X1 U23199 ( .A1(n14966), .A2(n20291), .B1(n21003), .B2(n20290), .ZN(
        n20819) );
  AOI22_X1 U23200 ( .A1(n20818), .A2(n20292), .B1(n20319), .B2(n20819), .ZN(
        n20293) );
  OAI211_X1 U23201 ( .C1(n20296), .C2(n20295), .A(n20294), .B(n20293), .ZN(
        P1_U3040) );
  INV_X1 U23202 ( .A(n20693), .ZN(n20776) );
  INV_X1 U23203 ( .A(n20359), .ZN(n20298) );
  INV_X1 U23204 ( .A(n20297), .ZN(n20687) );
  NOR2_X1 U23205 ( .A1(n20686), .A2(n20299), .ZN(n20317) );
  AOI21_X1 U23206 ( .B1(n20298), .B2(n20687), .A(n20317), .ZN(n20300) );
  OAI22_X1 U23207 ( .A1(n20300), .A2(n12580), .B1(n20299), .B2(n20898), .ZN(
        n20318) );
  AOI22_X1 U23208 ( .A1(n20765), .A2(n20318), .B1(n20764), .B2(n20317), .ZN(
        n20304) );
  OAI211_X1 U23209 ( .C1(n20368), .C2(n21280), .A(n20598), .B(n20300), .ZN(
        n20301) );
  OAI211_X1 U23210 ( .C1(n20598), .C2(n20302), .A(n20770), .B(n20301), .ZN(
        n20320) );
  AOI22_X1 U23211 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20320), .B1(
        n20319), .B2(n20773), .ZN(n20303) );
  OAI211_X1 U23212 ( .C1(n20776), .C2(n20351), .A(n20304), .B(n20303), .ZN(
        P1_U3041) );
  INV_X1 U23213 ( .A(n20697), .ZN(n20782) );
  AOI22_X1 U23214 ( .A1(n20778), .A2(n20318), .B1(n20777), .B2(n20317), .ZN(
        n20306) );
  AOI22_X1 U23215 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20320), .B1(
        n20319), .B2(n20779), .ZN(n20305) );
  OAI211_X1 U23216 ( .C1(n20782), .C2(n20351), .A(n20306), .B(n20305), .ZN(
        P1_U3042) );
  INV_X1 U23217 ( .A(n20785), .ZN(n20738) );
  AOI22_X1 U23218 ( .A1(n20784), .A2(n20318), .B1(n20783), .B2(n20317), .ZN(
        n20308) );
  AOI22_X1 U23219 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20320), .B1(
        n20319), .B2(n20735), .ZN(n20307) );
  OAI211_X1 U23220 ( .C1(n20738), .C2(n20351), .A(n20308), .B(n20307), .ZN(
        P1_U3043) );
  INV_X1 U23221 ( .A(n20791), .ZN(n20742) );
  AOI22_X1 U23222 ( .A1(n20790), .A2(n20318), .B1(n20789), .B2(n20317), .ZN(
        n20310) );
  AOI22_X1 U23223 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20320), .B1(
        n20319), .B2(n20739), .ZN(n20309) );
  OAI211_X1 U23224 ( .C1(n20742), .C2(n20351), .A(n20310), .B(n20309), .ZN(
        P1_U3044) );
  INV_X1 U23225 ( .A(n20797), .ZN(n20746) );
  AOI22_X1 U23226 ( .A1(n20796), .A2(n20318), .B1(n20795), .B2(n20317), .ZN(
        n20312) );
  AOI22_X1 U23227 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20320), .B1(
        n20319), .B2(n20743), .ZN(n20311) );
  OAI211_X1 U23228 ( .C1(n20746), .C2(n20351), .A(n20312), .B(n20311), .ZN(
        P1_U3045) );
  INV_X1 U23229 ( .A(n20707), .ZN(n20808) );
  AOI22_X1 U23230 ( .A1(n20802), .A2(n20318), .B1(n20801), .B2(n20317), .ZN(
        n20314) );
  AOI22_X1 U23231 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20320), .B1(
        n20319), .B2(n20803), .ZN(n20313) );
  OAI211_X1 U23232 ( .C1(n20808), .C2(n20351), .A(n20314), .B(n20313), .ZN(
        P1_U3046) );
  INV_X1 U23233 ( .A(n20811), .ZN(n20752) );
  AOI22_X1 U23234 ( .A1(n20810), .A2(n20318), .B1(n20809), .B2(n20317), .ZN(
        n20316) );
  AOI22_X1 U23235 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20320), .B1(
        n20319), .B2(n20749), .ZN(n20315) );
  OAI211_X1 U23236 ( .C1(n20752), .C2(n20351), .A(n20316), .B(n20315), .ZN(
        P1_U3047) );
  INV_X1 U23237 ( .A(n20819), .ZN(n20760) );
  AOI22_X1 U23238 ( .A1(n20818), .A2(n20318), .B1(n20816), .B2(n20317), .ZN(
        n20322) );
  AOI22_X1 U23239 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20320), .B1(
        n20319), .B2(n20755), .ZN(n20321) );
  OAI211_X1 U23240 ( .C1(n20760), .C2(n20351), .A(n20322), .B(n20321), .ZN(
        P1_U3048) );
  NAND2_X1 U23241 ( .A1(n20351), .A2(n20598), .ZN(n20324) );
  OAI21_X1 U23242 ( .B1(n20384), .B2(n20324), .A(n20628), .ZN(n20326) );
  NOR2_X1 U23243 ( .A1(n20359), .A2(n20558), .ZN(n20329) );
  INV_X1 U23244 ( .A(n20765), .ZN(n20645) );
  NOR3_X1 U23245 ( .A1(n20325), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20357) );
  NAND2_X1 U23246 ( .A1(n20686), .A2(n20357), .ZN(n20350) );
  INV_X1 U23247 ( .A(n20350), .ZN(n20343) );
  AOI22_X1 U23248 ( .A1(n20384), .A2(n20693), .B1(n20764), .B2(n20343), .ZN(
        n20332) );
  INV_X1 U23249 ( .A(n20326), .ZN(n20330) );
  NOR2_X1 U23250 ( .A1(n10355), .A2(n20898), .ZN(n20444) );
  AOI211_X1 U23251 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n20350), .A(n20444), 
        .B(n20327), .ZN(n20328) );
  INV_X1 U23252 ( .A(n20351), .ZN(n20344) );
  AOI22_X1 U23253 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20353), .B1(
        n20344), .B2(n20773), .ZN(n20331) );
  OAI211_X1 U23254 ( .C1(n20356), .C2(n20645), .A(n20332), .B(n20331), .ZN(
        P1_U3049) );
  INV_X1 U23255 ( .A(n20778), .ZN(n20651) );
  AOI22_X1 U23256 ( .A1(n20384), .A2(n20697), .B1(n20777), .B2(n20343), .ZN(
        n20334) );
  AOI22_X1 U23257 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20353), .B1(
        n20344), .B2(n20779), .ZN(n20333) );
  OAI211_X1 U23258 ( .C1(n20356), .C2(n20651), .A(n20334), .B(n20333), .ZN(
        P1_U3050) );
  INV_X1 U23259 ( .A(n20784), .ZN(n20656) );
  AOI22_X1 U23260 ( .A1(n20384), .A2(n20785), .B1(n20783), .B2(n20343), .ZN(
        n20336) );
  AOI22_X1 U23261 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20353), .B1(
        n20344), .B2(n20735), .ZN(n20335) );
  OAI211_X1 U23262 ( .C1(n20356), .C2(n20656), .A(n20336), .B(n20335), .ZN(
        P1_U3051) );
  INV_X1 U23263 ( .A(n20790), .ZN(n20661) );
  INV_X1 U23264 ( .A(n20739), .ZN(n20794) );
  INV_X1 U23265 ( .A(n20789), .ZN(n20657) );
  OAI22_X1 U23266 ( .A1(n20351), .A2(n20794), .B1(n20657), .B2(n20350), .ZN(
        n20337) );
  INV_X1 U23267 ( .A(n20337), .ZN(n20339) );
  AOI22_X1 U23268 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20353), .B1(
        n20384), .B2(n20791), .ZN(n20338) );
  OAI211_X1 U23269 ( .C1(n20356), .C2(n20661), .A(n20339), .B(n20338), .ZN(
        P1_U3052) );
  INV_X1 U23270 ( .A(n20796), .ZN(n20666) );
  INV_X1 U23271 ( .A(n20743), .ZN(n20800) );
  INV_X1 U23272 ( .A(n20795), .ZN(n20662) );
  OAI22_X1 U23273 ( .A1(n20351), .A2(n20800), .B1(n20662), .B2(n20350), .ZN(
        n20340) );
  INV_X1 U23274 ( .A(n20340), .ZN(n20342) );
  AOI22_X1 U23275 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20353), .B1(
        n20384), .B2(n20797), .ZN(n20341) );
  OAI211_X1 U23276 ( .C1(n20356), .C2(n20666), .A(n20342), .B(n20341), .ZN(
        P1_U3053) );
  INV_X1 U23277 ( .A(n20802), .ZN(n20671) );
  AOI22_X1 U23278 ( .A1(n20384), .A2(n20707), .B1(n20801), .B2(n20343), .ZN(
        n20346) );
  AOI22_X1 U23279 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20353), .B1(
        n20344), .B2(n20803), .ZN(n20345) );
  OAI211_X1 U23280 ( .C1(n20356), .C2(n20671), .A(n20346), .B(n20345), .ZN(
        P1_U3054) );
  INV_X1 U23281 ( .A(n20810), .ZN(n20676) );
  INV_X1 U23282 ( .A(n20749), .ZN(n20814) );
  INV_X1 U23283 ( .A(n20809), .ZN(n20672) );
  OAI22_X1 U23284 ( .A1(n20351), .A2(n20814), .B1(n20672), .B2(n20350), .ZN(
        n20347) );
  INV_X1 U23285 ( .A(n20347), .ZN(n20349) );
  AOI22_X1 U23286 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20353), .B1(
        n20384), .B2(n20811), .ZN(n20348) );
  OAI211_X1 U23287 ( .C1(n20356), .C2(n20676), .A(n20349), .B(n20348), .ZN(
        P1_U3055) );
  INV_X1 U23288 ( .A(n20818), .ZN(n20684) );
  INV_X1 U23289 ( .A(n20755), .ZN(n20825) );
  INV_X1 U23290 ( .A(n20816), .ZN(n20678) );
  OAI22_X1 U23291 ( .A1(n20351), .A2(n20825), .B1(n20678), .B2(n20350), .ZN(
        n20352) );
  INV_X1 U23292 ( .A(n20352), .ZN(n20355) );
  AOI22_X1 U23293 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20353), .B1(
        n20384), .B2(n20819), .ZN(n20354) );
  OAI211_X1 U23294 ( .C1(n20356), .C2(n20684), .A(n20355), .B(n20354), .ZN(
        P1_U3056) );
  INV_X1 U23295 ( .A(n20357), .ZN(n20364) );
  INV_X1 U23296 ( .A(n20472), .ZN(n20597) );
  AOI21_X1 U23297 ( .B1(n20368), .B2(n20598), .A(n20597), .ZN(n20367) );
  NAND2_X1 U23298 ( .A1(n11839), .A2(n20358), .ZN(n20593) );
  OR2_X1 U23299 ( .A1(n20359), .A2(n20593), .ZN(n20361) );
  NOR2_X1 U23300 ( .A1(n20591), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20383) );
  INV_X1 U23301 ( .A(n20383), .ZN(n20360) );
  OAI22_X1 U23302 ( .A1(n20898), .A2(n20364), .B1(n20367), .B2(n20363), .ZN(
        n20362) );
  AOI22_X1 U23303 ( .A1(n20384), .A2(n20773), .B1(n20764), .B2(n20383), .ZN(
        n20370) );
  INV_X1 U23304 ( .A(n20363), .ZN(n20366) );
  INV_X1 U23305 ( .A(n20770), .ZN(n20600) );
  AOI21_X1 U23306 ( .B1(n12580), .B2(n20364), .A(n20600), .ZN(n20365) );
  OAI21_X1 U23307 ( .B1(n20367), .B2(n20366), .A(n20365), .ZN(n20385) );
  AOI22_X1 U23308 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20385), .B1(
        n20413), .B2(n20693), .ZN(n20369) );
  OAI211_X1 U23309 ( .C1(n20388), .C2(n20645), .A(n20370), .B(n20369), .ZN(
        P1_U3057) );
  AOI22_X1 U23310 ( .A1(n20384), .A2(n20779), .B1(n20777), .B2(n20383), .ZN(
        n20372) );
  AOI22_X1 U23311 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20385), .B1(
        n20413), .B2(n20697), .ZN(n20371) );
  OAI211_X1 U23312 ( .C1(n20388), .C2(n20651), .A(n20372), .B(n20371), .ZN(
        P1_U3058) );
  AOI22_X1 U23313 ( .A1(n20413), .A2(n20785), .B1(n20783), .B2(n20383), .ZN(
        n20374) );
  AOI22_X1 U23314 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20385), .B1(
        n20384), .B2(n20735), .ZN(n20373) );
  OAI211_X1 U23315 ( .C1(n20388), .C2(n20656), .A(n20374), .B(n20373), .ZN(
        P1_U3059) );
  AOI22_X1 U23316 ( .A1(n20384), .A2(n20739), .B1(n20789), .B2(n20383), .ZN(
        n20376) );
  AOI22_X1 U23317 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20385), .B1(
        n20413), .B2(n20791), .ZN(n20375) );
  OAI211_X1 U23318 ( .C1(n20388), .C2(n20661), .A(n20376), .B(n20375), .ZN(
        P1_U3060) );
  AOI22_X1 U23319 ( .A1(n20413), .A2(n20797), .B1(n20795), .B2(n20383), .ZN(
        n20378) );
  AOI22_X1 U23320 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20385), .B1(
        n20384), .B2(n20743), .ZN(n20377) );
  OAI211_X1 U23321 ( .C1(n20388), .C2(n20666), .A(n20378), .B(n20377), .ZN(
        P1_U3061) );
  AOI22_X1 U23322 ( .A1(n20413), .A2(n20707), .B1(n20801), .B2(n20383), .ZN(
        n20380) );
  AOI22_X1 U23323 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20385), .B1(
        n20384), .B2(n20803), .ZN(n20379) );
  OAI211_X1 U23324 ( .C1(n20388), .C2(n20671), .A(n20380), .B(n20379), .ZN(
        P1_U3062) );
  AOI22_X1 U23325 ( .A1(n20384), .A2(n20749), .B1(n20809), .B2(n20383), .ZN(
        n20382) );
  AOI22_X1 U23326 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20385), .B1(
        n20413), .B2(n20811), .ZN(n20381) );
  OAI211_X1 U23327 ( .C1(n20388), .C2(n20676), .A(n20382), .B(n20381), .ZN(
        P1_U3063) );
  AOI22_X1 U23328 ( .A1(n20384), .A2(n20755), .B1(n20816), .B2(n20383), .ZN(
        n20387) );
  AOI22_X1 U23329 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20385), .B1(
        n20413), .B2(n20819), .ZN(n20386) );
  OAI211_X1 U23330 ( .C1(n20388), .C2(n20684), .A(n20387), .B(n20386), .ZN(
        P1_U3064) );
  INV_X1 U23331 ( .A(n20633), .ZN(n20721) );
  NOR2_X1 U23332 ( .A1(n20631), .A2(n20389), .ZN(n20469) );
  NAND3_X1 U23333 ( .A1(n20469), .A2(n20627), .A3(n20558), .ZN(n20390) );
  OAI21_X1 U23334 ( .B1(n20391), .B2(n20721), .A(n20390), .ZN(n20412) );
  NOR3_X1 U23335 ( .A1(n15858), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20420) );
  INV_X1 U23336 ( .A(n20420), .ZN(n20417) );
  NOR2_X1 U23337 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20417), .ZN(
        n20411) );
  AOI22_X1 U23338 ( .A1(n20765), .A2(n20412), .B1(n20764), .B2(n20411), .ZN(
        n20398) );
  INV_X1 U23339 ( .A(n20413), .ZN(n20392) );
  AOI21_X1 U23340 ( .B1(n20392), .B2(n20440), .A(n21280), .ZN(n20393) );
  AOI21_X1 U23341 ( .B1(n20469), .B2(n20558), .A(n20393), .ZN(n20394) );
  NOR2_X1 U23342 ( .A1(n20394), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20396) );
  AOI22_X1 U23343 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20414), .B1(
        n20413), .B2(n20773), .ZN(n20397) );
  OAI211_X1 U23344 ( .C1(n20776), .C2(n20440), .A(n20398), .B(n20397), .ZN(
        P1_U3065) );
  AOI22_X1 U23345 ( .A1(n20778), .A2(n20412), .B1(n20777), .B2(n20411), .ZN(
        n20400) );
  AOI22_X1 U23346 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20414), .B1(
        n20413), .B2(n20779), .ZN(n20399) );
  OAI211_X1 U23347 ( .C1(n20782), .C2(n20440), .A(n20400), .B(n20399), .ZN(
        P1_U3066) );
  AOI22_X1 U23348 ( .A1(n20784), .A2(n20412), .B1(n20783), .B2(n20411), .ZN(
        n20402) );
  AOI22_X1 U23349 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20414), .B1(
        n20413), .B2(n20735), .ZN(n20401) );
  OAI211_X1 U23350 ( .C1(n20738), .C2(n20440), .A(n20402), .B(n20401), .ZN(
        P1_U3067) );
  AOI22_X1 U23351 ( .A1(n20790), .A2(n20412), .B1(n20789), .B2(n20411), .ZN(
        n20404) );
  AOI22_X1 U23352 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20414), .B1(
        n20413), .B2(n20739), .ZN(n20403) );
  OAI211_X1 U23353 ( .C1(n20742), .C2(n20440), .A(n20404), .B(n20403), .ZN(
        P1_U3068) );
  AOI22_X1 U23354 ( .A1(n20796), .A2(n20412), .B1(n20795), .B2(n20411), .ZN(
        n20406) );
  AOI22_X1 U23355 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20414), .B1(
        n20413), .B2(n20743), .ZN(n20405) );
  OAI211_X1 U23356 ( .C1(n20746), .C2(n20440), .A(n20406), .B(n20405), .ZN(
        P1_U3069) );
  AOI22_X1 U23357 ( .A1(n20802), .A2(n20412), .B1(n20801), .B2(n20411), .ZN(
        n20408) );
  AOI22_X1 U23358 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20414), .B1(
        n20413), .B2(n20803), .ZN(n20407) );
  OAI211_X1 U23359 ( .C1(n20808), .C2(n20440), .A(n20408), .B(n20407), .ZN(
        P1_U3070) );
  AOI22_X1 U23360 ( .A1(n20810), .A2(n20412), .B1(n20809), .B2(n20411), .ZN(
        n20410) );
  AOI22_X1 U23361 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20414), .B1(
        n20413), .B2(n20749), .ZN(n20409) );
  OAI211_X1 U23362 ( .C1(n20752), .C2(n20440), .A(n20410), .B(n20409), .ZN(
        P1_U3071) );
  AOI22_X1 U23363 ( .A1(n20818), .A2(n20412), .B1(n20816), .B2(n20411), .ZN(
        n20416) );
  AOI22_X1 U23364 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20414), .B1(
        n20413), .B2(n20755), .ZN(n20415) );
  OAI211_X1 U23365 ( .C1(n20760), .C2(n20440), .A(n20416), .B(n20415), .ZN(
        P1_U3072) );
  INV_X1 U23366 ( .A(n20773), .ZN(n20696) );
  NOR2_X1 U23367 ( .A1(n20686), .A2(n20417), .ZN(n20435) );
  AOI21_X1 U23368 ( .B1(n20469), .B2(n20687), .A(n20435), .ZN(n20418) );
  OAI22_X1 U23369 ( .A1(n20418), .A2(n12580), .B1(n20417), .B2(n20898), .ZN(
        n20436) );
  AOI22_X1 U23370 ( .A1(n20765), .A2(n20436), .B1(n20764), .B2(n20435), .ZN(
        n20422) );
  OAI211_X1 U23371 ( .C1(n20471), .C2(n21280), .A(n20598), .B(n20418), .ZN(
        n20419) );
  OAI211_X1 U23372 ( .C1(n20598), .C2(n20420), .A(n20770), .B(n20419), .ZN(
        n20437) );
  AOI22_X1 U23373 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20437), .B1(
        n20464), .B2(n20693), .ZN(n20421) );
  OAI211_X1 U23374 ( .C1(n20696), .C2(n20440), .A(n20422), .B(n20421), .ZN(
        P1_U3073) );
  INV_X1 U23375 ( .A(n20779), .ZN(n20700) );
  AOI22_X1 U23376 ( .A1(n20778), .A2(n20436), .B1(n20777), .B2(n20435), .ZN(
        n20424) );
  AOI22_X1 U23377 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20437), .B1(
        n20464), .B2(n20697), .ZN(n20423) );
  OAI211_X1 U23378 ( .C1(n20700), .C2(n20440), .A(n20424), .B(n20423), .ZN(
        P1_U3074) );
  INV_X1 U23379 ( .A(n20735), .ZN(n20788) );
  AOI22_X1 U23380 ( .A1(n20784), .A2(n20436), .B1(n20783), .B2(n20435), .ZN(
        n20426) );
  AOI22_X1 U23381 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20437), .B1(
        n20464), .B2(n20785), .ZN(n20425) );
  OAI211_X1 U23382 ( .C1(n20788), .C2(n20440), .A(n20426), .B(n20425), .ZN(
        P1_U3075) );
  AOI22_X1 U23383 ( .A1(n20790), .A2(n20436), .B1(n20789), .B2(n20435), .ZN(
        n20428) );
  AOI22_X1 U23384 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20437), .B1(
        n20464), .B2(n20791), .ZN(n20427) );
  OAI211_X1 U23385 ( .C1(n20794), .C2(n20440), .A(n20428), .B(n20427), .ZN(
        P1_U3076) );
  AOI22_X1 U23386 ( .A1(n20796), .A2(n20436), .B1(n20795), .B2(n20435), .ZN(
        n20430) );
  AOI22_X1 U23387 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20437), .B1(
        n20464), .B2(n20797), .ZN(n20429) );
  OAI211_X1 U23388 ( .C1(n20800), .C2(n20440), .A(n20430), .B(n20429), .ZN(
        P1_U3077) );
  INV_X1 U23389 ( .A(n20803), .ZN(n20710) );
  AOI22_X1 U23390 ( .A1(n20802), .A2(n20436), .B1(n20801), .B2(n20435), .ZN(
        n20432) );
  AOI22_X1 U23391 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20437), .B1(
        n20464), .B2(n20707), .ZN(n20431) );
  OAI211_X1 U23392 ( .C1(n20710), .C2(n20440), .A(n20432), .B(n20431), .ZN(
        P1_U3078) );
  AOI22_X1 U23393 ( .A1(n20810), .A2(n20436), .B1(n20809), .B2(n20435), .ZN(
        n20434) );
  AOI22_X1 U23394 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20437), .B1(
        n20464), .B2(n20811), .ZN(n20433) );
  OAI211_X1 U23395 ( .C1(n20814), .C2(n20440), .A(n20434), .B(n20433), .ZN(
        P1_U3079) );
  AOI22_X1 U23396 ( .A1(n20818), .A2(n20436), .B1(n20816), .B2(n20435), .ZN(
        n20439) );
  AOI22_X1 U23397 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20437), .B1(
        n20464), .B2(n20819), .ZN(n20438) );
  OAI211_X1 U23398 ( .C1(n20825), .C2(n20440), .A(n20439), .B(n20438), .ZN(
        P1_U3080) );
  NAND3_X1 U23399 ( .A1(n20448), .A2(n20441), .A3(n20598), .ZN(n20442) );
  NAND2_X1 U23400 ( .A1(n20442), .A2(n20628), .ZN(n20446) );
  AND2_X1 U23401 ( .A1(n20469), .A2(n20726), .ZN(n20443) );
  NOR2_X1 U23402 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20470), .ZN(
        n20463) );
  AOI22_X1 U23403 ( .A1(n20464), .A2(n20773), .B1(n20764), .B2(n20463), .ZN(
        n20450) );
  INV_X1 U23404 ( .A(n20443), .ZN(n20445) );
  AOI21_X1 U23405 ( .B1(n20446), .B2(n20445), .A(n20444), .ZN(n20447) );
  OAI211_X1 U23406 ( .C1(n20463), .C2(n20641), .A(n20729), .B(n20447), .ZN(
        n20465) );
  AOI22_X1 U23407 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20465), .B1(
        n20494), .B2(n20693), .ZN(n20449) );
  OAI211_X1 U23408 ( .C1(n20468), .C2(n20645), .A(n20450), .B(n20449), .ZN(
        P1_U3081) );
  AOI22_X1 U23409 ( .A1(n20494), .A2(n20697), .B1(n20777), .B2(n20463), .ZN(
        n20452) );
  AOI22_X1 U23410 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20465), .B1(
        n20464), .B2(n20779), .ZN(n20451) );
  OAI211_X1 U23411 ( .C1(n20468), .C2(n20651), .A(n20452), .B(n20451), .ZN(
        P1_U3082) );
  AOI22_X1 U23412 ( .A1(n20464), .A2(n20735), .B1(n20783), .B2(n20463), .ZN(
        n20454) );
  AOI22_X1 U23413 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20465), .B1(
        n20494), .B2(n20785), .ZN(n20453) );
  OAI211_X1 U23414 ( .C1(n20468), .C2(n20656), .A(n20454), .B(n20453), .ZN(
        P1_U3083) );
  AOI22_X1 U23415 ( .A1(n20464), .A2(n20739), .B1(n20789), .B2(n20463), .ZN(
        n20456) );
  AOI22_X1 U23416 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20465), .B1(
        n20494), .B2(n20791), .ZN(n20455) );
  OAI211_X1 U23417 ( .C1(n20468), .C2(n20661), .A(n20456), .B(n20455), .ZN(
        P1_U3084) );
  AOI22_X1 U23418 ( .A1(n20494), .A2(n20797), .B1(n20795), .B2(n20463), .ZN(
        n20458) );
  AOI22_X1 U23419 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20465), .B1(
        n20464), .B2(n20743), .ZN(n20457) );
  OAI211_X1 U23420 ( .C1(n20468), .C2(n20666), .A(n20458), .B(n20457), .ZN(
        P1_U3085) );
  AOI22_X1 U23421 ( .A1(n20464), .A2(n20803), .B1(n20801), .B2(n20463), .ZN(
        n20460) );
  AOI22_X1 U23422 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20465), .B1(
        n20494), .B2(n20707), .ZN(n20459) );
  OAI211_X1 U23423 ( .C1(n20468), .C2(n20671), .A(n20460), .B(n20459), .ZN(
        P1_U3086) );
  AOI22_X1 U23424 ( .A1(n20464), .A2(n20749), .B1(n20809), .B2(n20463), .ZN(
        n20462) );
  AOI22_X1 U23425 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20465), .B1(
        n20494), .B2(n20811), .ZN(n20461) );
  OAI211_X1 U23426 ( .C1(n20468), .C2(n20676), .A(n20462), .B(n20461), .ZN(
        P1_U3087) );
  AOI22_X1 U23427 ( .A1(n20464), .A2(n20755), .B1(n20816), .B2(n20463), .ZN(
        n20467) );
  AOI22_X1 U23428 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20465), .B1(
        n20494), .B2(n20819), .ZN(n20466) );
  OAI211_X1 U23429 ( .C1(n20468), .C2(n20684), .A(n20467), .B(n20466), .ZN(
        P1_U3088) );
  INV_X1 U23430 ( .A(n20593), .ZN(n20761) );
  AOI21_X1 U23431 ( .B1(n20469), .B2(n20761), .A(n20492), .ZN(n20474) );
  OAI22_X1 U23432 ( .A1(n20474), .A2(n12580), .B1(n20470), .B2(n20898), .ZN(
        n20493) );
  AOI22_X1 U23433 ( .A1(n20765), .A2(n20493), .B1(n20764), .B2(n20492), .ZN(
        n20479) );
  INV_X1 U23434 ( .A(n20470), .ZN(n20477) );
  INV_X1 U23435 ( .A(n20471), .ZN(n20473) );
  OAI21_X1 U23436 ( .B1(n20473), .B2(n12580), .A(n20472), .ZN(n20475) );
  NAND2_X1 U23437 ( .A1(n20475), .A2(n20474), .ZN(n20476) );
  OAI211_X1 U23438 ( .C1(n20477), .C2(n20598), .A(n20770), .B(n20476), .ZN(
        n20495) );
  AOI22_X1 U23439 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20495), .B1(
        n20494), .B2(n20773), .ZN(n20478) );
  OAI211_X1 U23440 ( .C1(n20776), .C2(n20504), .A(n20479), .B(n20478), .ZN(
        P1_U3089) );
  AOI22_X1 U23441 ( .A1(n20778), .A2(n20493), .B1(n20777), .B2(n20492), .ZN(
        n20481) );
  AOI22_X1 U23442 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20495), .B1(
        n20494), .B2(n20779), .ZN(n20480) );
  OAI211_X1 U23443 ( .C1(n20782), .C2(n20504), .A(n20481), .B(n20480), .ZN(
        P1_U3090) );
  AOI22_X1 U23444 ( .A1(n20784), .A2(n20493), .B1(n20783), .B2(n20492), .ZN(
        n20483) );
  AOI22_X1 U23445 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20495), .B1(
        n20494), .B2(n20735), .ZN(n20482) );
  OAI211_X1 U23446 ( .C1(n20738), .C2(n20504), .A(n20483), .B(n20482), .ZN(
        P1_U3091) );
  AOI22_X1 U23447 ( .A1(n20790), .A2(n20493), .B1(n20789), .B2(n20492), .ZN(
        n20485) );
  AOI22_X1 U23448 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20495), .B1(
        n20494), .B2(n20739), .ZN(n20484) );
  OAI211_X1 U23449 ( .C1(n20742), .C2(n20504), .A(n20485), .B(n20484), .ZN(
        P1_U3092) );
  AOI22_X1 U23450 ( .A1(n20796), .A2(n20493), .B1(n20795), .B2(n20492), .ZN(
        n20487) );
  AOI22_X1 U23451 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20495), .B1(
        n20494), .B2(n20743), .ZN(n20486) );
  OAI211_X1 U23452 ( .C1(n20746), .C2(n20504), .A(n20487), .B(n20486), .ZN(
        P1_U3093) );
  AOI22_X1 U23453 ( .A1(n20802), .A2(n20493), .B1(n20801), .B2(n20492), .ZN(
        n20489) );
  AOI22_X1 U23454 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20495), .B1(
        n20494), .B2(n20803), .ZN(n20488) );
  OAI211_X1 U23455 ( .C1(n20808), .C2(n20504), .A(n20489), .B(n20488), .ZN(
        P1_U3094) );
  AOI22_X1 U23456 ( .A1(n20810), .A2(n20493), .B1(n20809), .B2(n20492), .ZN(
        n20491) );
  AOI22_X1 U23457 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20495), .B1(
        n20494), .B2(n20749), .ZN(n20490) );
  OAI211_X1 U23458 ( .C1(n20752), .C2(n20504), .A(n20491), .B(n20490), .ZN(
        P1_U3095) );
  AOI22_X1 U23459 ( .A1(n20818), .A2(n20493), .B1(n20816), .B2(n20492), .ZN(
        n20497) );
  AOI22_X1 U23460 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20495), .B1(
        n20494), .B2(n20755), .ZN(n20496) );
  OAI211_X1 U23461 ( .C1(n20760), .C2(n20504), .A(n20497), .B(n20496), .ZN(
        P1_U3096) );
  INV_X1 U23462 ( .A(n20498), .ZN(n20499) );
  NAND2_X1 U23463 ( .A1(n20500), .A2(n20631), .ZN(n20594) );
  INV_X1 U23464 ( .A(n20594), .ZN(n20529) );
  NOR3_X1 U23465 ( .A1(n20634), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20533) );
  INV_X1 U23466 ( .A(n20533), .ZN(n20530) );
  NOR2_X1 U23467 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20530), .ZN(
        n20523) );
  AOI21_X1 U23468 ( .B1(n20529), .B2(n20558), .A(n20523), .ZN(n20506) );
  INV_X1 U23469 ( .A(n20559), .ZN(n20502) );
  NOR2_X1 U23470 ( .A1(n20502), .A2(n20501), .ZN(n20632) );
  INV_X1 U23471 ( .A(n20632), .ZN(n20637) );
  OAI22_X1 U23472 ( .A1(n20506), .A2(n12580), .B1(n20637), .B2(n20503), .ZN(
        n20524) );
  AOI22_X1 U23473 ( .A1(n20765), .A2(n20524), .B1(n20764), .B2(n20523), .ZN(
        n20510) );
  INV_X1 U23474 ( .A(n20554), .ZN(n20505) );
  OAI21_X1 U23475 ( .B1(n20505), .B2(n20525), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20507) );
  NAND2_X1 U23476 ( .A1(n20507), .A2(n20506), .ZN(n20508) );
  AOI22_X1 U23477 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20526), .B1(
        n20525), .B2(n20773), .ZN(n20509) );
  OAI211_X1 U23478 ( .C1(n20776), .C2(n20554), .A(n20510), .B(n20509), .ZN(
        P1_U3097) );
  AOI22_X1 U23479 ( .A1(n20778), .A2(n20524), .B1(n20777), .B2(n20523), .ZN(
        n20512) );
  AOI22_X1 U23480 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20526), .B1(
        n20525), .B2(n20779), .ZN(n20511) );
  OAI211_X1 U23481 ( .C1(n20782), .C2(n20554), .A(n20512), .B(n20511), .ZN(
        P1_U3098) );
  AOI22_X1 U23482 ( .A1(n20784), .A2(n20524), .B1(n20783), .B2(n20523), .ZN(
        n20514) );
  AOI22_X1 U23483 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20526), .B1(
        n20525), .B2(n20735), .ZN(n20513) );
  OAI211_X1 U23484 ( .C1(n20738), .C2(n20554), .A(n20514), .B(n20513), .ZN(
        P1_U3099) );
  AOI22_X1 U23485 ( .A1(n20790), .A2(n20524), .B1(n20789), .B2(n20523), .ZN(
        n20516) );
  AOI22_X1 U23486 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20526), .B1(
        n20525), .B2(n20739), .ZN(n20515) );
  OAI211_X1 U23487 ( .C1(n20742), .C2(n20554), .A(n20516), .B(n20515), .ZN(
        P1_U3100) );
  AOI22_X1 U23488 ( .A1(n20796), .A2(n20524), .B1(n20795), .B2(n20523), .ZN(
        n20518) );
  AOI22_X1 U23489 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20526), .B1(
        n20525), .B2(n20743), .ZN(n20517) );
  OAI211_X1 U23490 ( .C1(n20746), .C2(n20554), .A(n20518), .B(n20517), .ZN(
        P1_U3101) );
  AOI22_X1 U23491 ( .A1(n20802), .A2(n20524), .B1(n20801), .B2(n20523), .ZN(
        n20520) );
  AOI22_X1 U23492 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20526), .B1(
        n20525), .B2(n20803), .ZN(n20519) );
  OAI211_X1 U23493 ( .C1(n20808), .C2(n20554), .A(n20520), .B(n20519), .ZN(
        P1_U3102) );
  AOI22_X1 U23494 ( .A1(n20810), .A2(n20524), .B1(n20809), .B2(n20523), .ZN(
        n20522) );
  AOI22_X1 U23495 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20526), .B1(
        n20525), .B2(n20749), .ZN(n20521) );
  OAI211_X1 U23496 ( .C1(n20752), .C2(n20554), .A(n20522), .B(n20521), .ZN(
        P1_U3103) );
  AOI22_X1 U23497 ( .A1(n20818), .A2(n20524), .B1(n20816), .B2(n20523), .ZN(
        n20528) );
  AOI22_X1 U23498 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20526), .B1(
        n20525), .B2(n20755), .ZN(n20527) );
  OAI211_X1 U23499 ( .C1(n20760), .C2(n20554), .A(n20528), .B(n20527), .ZN(
        P1_U3104) );
  NOR2_X1 U23500 ( .A1(n20686), .A2(n20530), .ZN(n20549) );
  AOI21_X1 U23501 ( .B1(n20529), .B2(n20687), .A(n20549), .ZN(n20531) );
  OAI22_X1 U23502 ( .A1(n20531), .A2(n12580), .B1(n20530), .B2(n20898), .ZN(
        n20550) );
  AOI22_X1 U23503 ( .A1(n20765), .A2(n20550), .B1(n20764), .B2(n20549), .ZN(
        n20536) );
  INV_X1 U23504 ( .A(n20590), .ZN(n20599) );
  OAI211_X1 U23505 ( .C1(n20599), .C2(n21280), .A(n20598), .B(n20531), .ZN(
        n20532) );
  OAI211_X1 U23506 ( .C1(n20598), .C2(n20533), .A(n20770), .B(n20532), .ZN(
        n20551) );
  AOI22_X1 U23507 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20551), .B1(
        n20583), .B2(n20693), .ZN(n20535) );
  OAI211_X1 U23508 ( .C1(n20696), .C2(n20554), .A(n20536), .B(n20535), .ZN(
        P1_U3105) );
  AOI22_X1 U23509 ( .A1(n20778), .A2(n20550), .B1(n20777), .B2(n20549), .ZN(
        n20538) );
  AOI22_X1 U23510 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20551), .B1(
        n20583), .B2(n20697), .ZN(n20537) );
  OAI211_X1 U23511 ( .C1(n20700), .C2(n20554), .A(n20538), .B(n20537), .ZN(
        P1_U3106) );
  AOI22_X1 U23512 ( .A1(n20784), .A2(n20550), .B1(n20783), .B2(n20549), .ZN(
        n20540) );
  AOI22_X1 U23513 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20551), .B1(
        n20583), .B2(n20785), .ZN(n20539) );
  OAI211_X1 U23514 ( .C1(n20788), .C2(n20554), .A(n20540), .B(n20539), .ZN(
        P1_U3107) );
  AOI22_X1 U23515 ( .A1(n20790), .A2(n20550), .B1(n20789), .B2(n20549), .ZN(
        n20542) );
  AOI22_X1 U23516 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20551), .B1(
        n20583), .B2(n20791), .ZN(n20541) );
  OAI211_X1 U23517 ( .C1(n20794), .C2(n20554), .A(n20542), .B(n20541), .ZN(
        P1_U3108) );
  AOI22_X1 U23518 ( .A1(n20796), .A2(n20550), .B1(n20795), .B2(n20549), .ZN(
        n20544) );
  AOI22_X1 U23519 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20551), .B1(
        n20583), .B2(n20797), .ZN(n20543) );
  OAI211_X1 U23520 ( .C1(n20800), .C2(n20554), .A(n20544), .B(n20543), .ZN(
        P1_U3109) );
  AOI22_X1 U23521 ( .A1(n20802), .A2(n20550), .B1(n20801), .B2(n20549), .ZN(
        n20546) );
  AOI22_X1 U23522 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20551), .B1(
        n20583), .B2(n20707), .ZN(n20545) );
  OAI211_X1 U23523 ( .C1(n20710), .C2(n20554), .A(n20546), .B(n20545), .ZN(
        P1_U3110) );
  AOI22_X1 U23524 ( .A1(n20810), .A2(n20550), .B1(n20809), .B2(n20549), .ZN(
        n20548) );
  AOI22_X1 U23525 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20551), .B1(
        n20583), .B2(n20811), .ZN(n20547) );
  OAI211_X1 U23526 ( .C1(n20814), .C2(n20554), .A(n20548), .B(n20547), .ZN(
        P1_U3111) );
  AOI22_X1 U23527 ( .A1(n20818), .A2(n20550), .B1(n20816), .B2(n20549), .ZN(
        n20553) );
  AOI22_X1 U23528 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20551), .B1(
        n20583), .B2(n20819), .ZN(n20552) );
  OAI211_X1 U23529 ( .C1(n20825), .C2(n20554), .A(n20553), .B(n20552), .ZN(
        P1_U3112) );
  INV_X1 U23530 ( .A(n20583), .ZN(n20555) );
  NAND2_X1 U23531 ( .A1(n20555), .A2(n20598), .ZN(n20557) );
  OAI21_X1 U23532 ( .B1(n20557), .B2(n20621), .A(n20628), .ZN(n20566) );
  NOR2_X1 U23533 ( .A1(n20594), .A2(n20558), .ZN(n20562) );
  OR2_X1 U23534 ( .A1(n20559), .A2(n20634), .ZN(n20720) );
  INV_X1 U23535 ( .A(n20720), .ZN(n20560) );
  NAND3_X1 U23536 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n15858), .ZN(n20601) );
  NOR2_X1 U23537 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20601), .ZN(
        n20582) );
  AOI22_X1 U23538 ( .A1(n20583), .A2(n20773), .B1(n20764), .B2(n20582), .ZN(
        n20569) );
  INV_X1 U23539 ( .A(n20562), .ZN(n20565) );
  NAND2_X1 U23540 ( .A1(n20720), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20728) );
  OAI211_X1 U23541 ( .C1(n20641), .C2(n20582), .A(n20728), .B(n20563), .ZN(
        n20564) );
  AOI21_X1 U23542 ( .B1(n20566), .B2(n20565), .A(n20564), .ZN(n20567) );
  AOI22_X1 U23543 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20584), .B1(
        n20621), .B2(n20693), .ZN(n20568) );
  OAI211_X1 U23544 ( .C1(n20587), .C2(n20645), .A(n20569), .B(n20568), .ZN(
        P1_U3113) );
  AOI22_X1 U23545 ( .A1(n20621), .A2(n20697), .B1(n20777), .B2(n20582), .ZN(
        n20571) );
  AOI22_X1 U23546 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20584), .B1(
        n20583), .B2(n20779), .ZN(n20570) );
  OAI211_X1 U23547 ( .C1(n20587), .C2(n20651), .A(n20571), .B(n20570), .ZN(
        P1_U3114) );
  AOI22_X1 U23548 ( .A1(n20621), .A2(n20785), .B1(n20783), .B2(n20582), .ZN(
        n20573) );
  AOI22_X1 U23549 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20584), .B1(
        n20583), .B2(n20735), .ZN(n20572) );
  OAI211_X1 U23550 ( .C1(n20587), .C2(n20656), .A(n20573), .B(n20572), .ZN(
        P1_U3115) );
  AOI22_X1 U23551 ( .A1(n20621), .A2(n20791), .B1(n20789), .B2(n20582), .ZN(
        n20575) );
  AOI22_X1 U23552 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20584), .B1(
        n20583), .B2(n20739), .ZN(n20574) );
  OAI211_X1 U23553 ( .C1(n20587), .C2(n20661), .A(n20575), .B(n20574), .ZN(
        P1_U3116) );
  AOI22_X1 U23554 ( .A1(n20583), .A2(n20743), .B1(n20795), .B2(n20582), .ZN(
        n20577) );
  AOI22_X1 U23555 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20584), .B1(
        n20621), .B2(n20797), .ZN(n20576) );
  OAI211_X1 U23556 ( .C1(n20587), .C2(n20666), .A(n20577), .B(n20576), .ZN(
        P1_U3117) );
  AOI22_X1 U23557 ( .A1(n20583), .A2(n20803), .B1(n20801), .B2(n20582), .ZN(
        n20579) );
  AOI22_X1 U23558 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20584), .B1(
        n20621), .B2(n20707), .ZN(n20578) );
  OAI211_X1 U23559 ( .C1(n20587), .C2(n20671), .A(n20579), .B(n20578), .ZN(
        P1_U3118) );
  AOI22_X1 U23560 ( .A1(n20583), .A2(n20749), .B1(n20809), .B2(n20582), .ZN(
        n20581) );
  AOI22_X1 U23561 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20584), .B1(
        n20621), .B2(n20811), .ZN(n20580) );
  OAI211_X1 U23562 ( .C1(n20587), .C2(n20676), .A(n20581), .B(n20580), .ZN(
        P1_U3119) );
  AOI22_X1 U23563 ( .A1(n20621), .A2(n20819), .B1(n20816), .B2(n20582), .ZN(
        n20586) );
  AOI22_X1 U23564 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20584), .B1(
        n20583), .B2(n20755), .ZN(n20585) );
  OAI211_X1 U23565 ( .C1(n20587), .C2(n20684), .A(n20586), .B(n20585), .ZN(
        P1_U3120) );
  INV_X1 U23566 ( .A(n20588), .ZN(n20589) );
  INV_X1 U23567 ( .A(n20591), .ZN(n20592) );
  NAND2_X1 U23568 ( .A1(n20592), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20596) );
  OAI21_X1 U23569 ( .B1(n20594), .B2(n20593), .A(n20596), .ZN(n20603) );
  INV_X1 U23570 ( .A(n20603), .ZN(n20595) );
  OAI22_X1 U23571 ( .A1(n20595), .A2(n12580), .B1(n20601), .B2(n20898), .ZN(
        n20620) );
  INV_X1 U23572 ( .A(n20596), .ZN(n20619) );
  AOI22_X1 U23573 ( .A1(n20765), .A2(n20620), .B1(n20764), .B2(n20619), .ZN(
        n20606) );
  AOI21_X1 U23574 ( .B1(n20599), .B2(n20598), .A(n20597), .ZN(n20604) );
  AOI21_X1 U23575 ( .B1(n20601), .B2(n12580), .A(n20600), .ZN(n20602) );
  AOI22_X1 U23576 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20773), .ZN(n20605) );
  OAI211_X1 U23577 ( .C1(n20776), .C2(n20642), .A(n20606), .B(n20605), .ZN(
        P1_U3121) );
  AOI22_X1 U23578 ( .A1(n20778), .A2(n20620), .B1(n20777), .B2(n20619), .ZN(
        n20608) );
  AOI22_X1 U23579 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20779), .ZN(n20607) );
  OAI211_X1 U23580 ( .C1(n20782), .C2(n20642), .A(n20608), .B(n20607), .ZN(
        P1_U3122) );
  AOI22_X1 U23581 ( .A1(n20784), .A2(n20620), .B1(n20783), .B2(n20619), .ZN(
        n20610) );
  AOI22_X1 U23582 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20735), .ZN(n20609) );
  OAI211_X1 U23583 ( .C1(n20738), .C2(n20642), .A(n20610), .B(n20609), .ZN(
        P1_U3123) );
  AOI22_X1 U23584 ( .A1(n20790), .A2(n20620), .B1(n20789), .B2(n20619), .ZN(
        n20612) );
  AOI22_X1 U23585 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20739), .ZN(n20611) );
  OAI211_X1 U23586 ( .C1(n20742), .C2(n20642), .A(n20612), .B(n20611), .ZN(
        P1_U3124) );
  AOI22_X1 U23587 ( .A1(n20796), .A2(n20620), .B1(n20795), .B2(n20619), .ZN(
        n20614) );
  AOI22_X1 U23588 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20743), .ZN(n20613) );
  OAI211_X1 U23589 ( .C1(n20746), .C2(n20642), .A(n20614), .B(n20613), .ZN(
        P1_U3125) );
  AOI22_X1 U23590 ( .A1(n20802), .A2(n20620), .B1(n20801), .B2(n20619), .ZN(
        n20616) );
  AOI22_X1 U23591 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20803), .ZN(n20615) );
  OAI211_X1 U23592 ( .C1(n20808), .C2(n20642), .A(n20616), .B(n20615), .ZN(
        P1_U3126) );
  AOI22_X1 U23593 ( .A1(n20810), .A2(n20620), .B1(n20809), .B2(n20619), .ZN(
        n20618) );
  AOI22_X1 U23594 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20749), .ZN(n20617) );
  OAI211_X1 U23595 ( .C1(n20752), .C2(n20642), .A(n20618), .B(n20617), .ZN(
        P1_U3127) );
  AOI22_X1 U23596 ( .A1(n20818), .A2(n20620), .B1(n20816), .B2(n20619), .ZN(
        n20624) );
  AOI22_X1 U23597 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20755), .ZN(n20623) );
  OAI211_X1 U23598 ( .C1(n20760), .C2(n20642), .A(n20624), .B(n20623), .ZN(
        P1_U3128) );
  NAND3_X1 U23599 ( .A1(n20642), .A2(n20627), .A3(n20718), .ZN(n20629) );
  NAND2_X1 U23600 ( .A1(n20629), .A2(n20628), .ZN(n20639) );
  OR2_X1 U23601 ( .A1(n20631), .A2(n20630), .ZN(n20723) );
  NOR2_X1 U23602 ( .A1(n20723), .A2(n20726), .ZN(n20636) );
  INV_X1 U23603 ( .A(n20718), .ZN(n20635) );
  NOR3_X1 U23604 ( .A1(n15858), .A2(n20634), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20691) );
  INV_X1 U23605 ( .A(n20691), .ZN(n20688) );
  NOR2_X1 U23606 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20688), .ZN(
        n20646) );
  AOI22_X1 U23607 ( .A1(n20635), .A2(n20693), .B1(n20764), .B2(n20646), .ZN(
        n20644) );
  INV_X1 U23608 ( .A(n20636), .ZN(n20638) );
  AOI22_X1 U23609 ( .A1(n20639), .A2(n20638), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20637), .ZN(n20640) );
  AOI22_X1 U23610 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20681), .B1(
        n20680), .B2(n20773), .ZN(n20643) );
  OAI211_X1 U23611 ( .C1(n20685), .C2(n20645), .A(n20644), .B(n20643), .ZN(
        P1_U3129) );
  INV_X1 U23612 ( .A(n20777), .ZN(n20647) );
  INV_X1 U23613 ( .A(n20646), .ZN(n20677) );
  OAI22_X1 U23614 ( .A1(n20718), .A2(n20782), .B1(n20647), .B2(n20677), .ZN(
        n20648) );
  INV_X1 U23615 ( .A(n20648), .ZN(n20650) );
  AOI22_X1 U23616 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20681), .B1(
        n20680), .B2(n20779), .ZN(n20649) );
  OAI211_X1 U23617 ( .C1(n20685), .C2(n20651), .A(n20650), .B(n20649), .ZN(
        P1_U3130) );
  INV_X1 U23618 ( .A(n20783), .ZN(n20652) );
  OAI22_X1 U23619 ( .A1(n20718), .A2(n20738), .B1(n20652), .B2(n20677), .ZN(
        n20653) );
  INV_X1 U23620 ( .A(n20653), .ZN(n20655) );
  AOI22_X1 U23621 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20681), .B1(
        n20680), .B2(n20735), .ZN(n20654) );
  OAI211_X1 U23622 ( .C1(n20685), .C2(n20656), .A(n20655), .B(n20654), .ZN(
        P1_U3131) );
  OAI22_X1 U23623 ( .A1(n20718), .A2(n20742), .B1(n20657), .B2(n20677), .ZN(
        n20658) );
  INV_X1 U23624 ( .A(n20658), .ZN(n20660) );
  AOI22_X1 U23625 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20681), .B1(
        n20680), .B2(n20739), .ZN(n20659) );
  OAI211_X1 U23626 ( .C1(n20685), .C2(n20661), .A(n20660), .B(n20659), .ZN(
        P1_U3132) );
  OAI22_X1 U23627 ( .A1(n20718), .A2(n20746), .B1(n20662), .B2(n20677), .ZN(
        n20663) );
  INV_X1 U23628 ( .A(n20663), .ZN(n20665) );
  AOI22_X1 U23629 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20681), .B1(
        n20680), .B2(n20743), .ZN(n20664) );
  OAI211_X1 U23630 ( .C1(n20685), .C2(n20666), .A(n20665), .B(n20664), .ZN(
        P1_U3133) );
  INV_X1 U23631 ( .A(n20801), .ZN(n20667) );
  OAI22_X1 U23632 ( .A1(n20718), .A2(n20808), .B1(n20667), .B2(n20677), .ZN(
        n20668) );
  INV_X1 U23633 ( .A(n20668), .ZN(n20670) );
  AOI22_X1 U23634 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20681), .B1(
        n20680), .B2(n20803), .ZN(n20669) );
  OAI211_X1 U23635 ( .C1(n20685), .C2(n20671), .A(n20670), .B(n20669), .ZN(
        P1_U3134) );
  OAI22_X1 U23636 ( .A1(n20718), .A2(n20752), .B1(n20672), .B2(n20677), .ZN(
        n20673) );
  INV_X1 U23637 ( .A(n20673), .ZN(n20675) );
  AOI22_X1 U23638 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20681), .B1(
        n20680), .B2(n20749), .ZN(n20674) );
  OAI211_X1 U23639 ( .C1(n20685), .C2(n20676), .A(n20675), .B(n20674), .ZN(
        P1_U3135) );
  OAI22_X1 U23640 ( .A1(n20718), .A2(n20760), .B1(n20678), .B2(n20677), .ZN(
        n20679) );
  INV_X1 U23641 ( .A(n20679), .ZN(n20683) );
  AOI22_X1 U23642 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20681), .B1(
        n20680), .B2(n20755), .ZN(n20682) );
  OAI211_X1 U23643 ( .C1(n20685), .C2(n20684), .A(n20683), .B(n20682), .ZN(
        P1_U3136) );
  INV_X1 U23644 ( .A(n20723), .ZN(n20762) );
  NOR2_X1 U23645 ( .A1(n20686), .A2(n20688), .ZN(n20713) );
  AOI21_X1 U23646 ( .B1(n20762), .B2(n20687), .A(n20713), .ZN(n20689) );
  OAI22_X1 U23647 ( .A1(n20689), .A2(n12580), .B1(n20688), .B2(n20898), .ZN(
        n20714) );
  AOI22_X1 U23648 ( .A1(n20765), .A2(n20714), .B1(n20764), .B2(n20713), .ZN(
        n20695) );
  OAI21_X1 U23649 ( .B1(n20691), .B2(n20690), .A(n20770), .ZN(n20715) );
  OR2_X1 U23650 ( .A1(n20769), .A2(n20692), .ZN(n20724) );
  AOI22_X1 U23651 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20715), .B1(
        n20756), .B2(n20693), .ZN(n20694) );
  OAI211_X1 U23652 ( .C1(n20696), .C2(n20718), .A(n20695), .B(n20694), .ZN(
        P1_U3137) );
  AOI22_X1 U23653 ( .A1(n20778), .A2(n20714), .B1(n20777), .B2(n20713), .ZN(
        n20699) );
  AOI22_X1 U23654 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20715), .B1(
        n20756), .B2(n20697), .ZN(n20698) );
  OAI211_X1 U23655 ( .C1(n20700), .C2(n20718), .A(n20699), .B(n20698), .ZN(
        P1_U3138) );
  AOI22_X1 U23656 ( .A1(n20784), .A2(n20714), .B1(n20783), .B2(n20713), .ZN(
        n20702) );
  AOI22_X1 U23657 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20715), .B1(
        n20756), .B2(n20785), .ZN(n20701) );
  OAI211_X1 U23658 ( .C1(n20788), .C2(n20718), .A(n20702), .B(n20701), .ZN(
        P1_U3139) );
  AOI22_X1 U23659 ( .A1(n20790), .A2(n20714), .B1(n20789), .B2(n20713), .ZN(
        n20704) );
  AOI22_X1 U23660 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20715), .B1(
        n20756), .B2(n20791), .ZN(n20703) );
  OAI211_X1 U23661 ( .C1(n20794), .C2(n20718), .A(n20704), .B(n20703), .ZN(
        P1_U3140) );
  AOI22_X1 U23662 ( .A1(n20796), .A2(n20714), .B1(n20795), .B2(n20713), .ZN(
        n20706) );
  AOI22_X1 U23663 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20715), .B1(
        n20756), .B2(n20797), .ZN(n20705) );
  OAI211_X1 U23664 ( .C1(n20800), .C2(n20718), .A(n20706), .B(n20705), .ZN(
        P1_U3141) );
  AOI22_X1 U23665 ( .A1(n20802), .A2(n20714), .B1(n20801), .B2(n20713), .ZN(
        n20709) );
  AOI22_X1 U23666 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20715), .B1(
        n20756), .B2(n20707), .ZN(n20708) );
  OAI211_X1 U23667 ( .C1(n20710), .C2(n20718), .A(n20709), .B(n20708), .ZN(
        P1_U3142) );
  AOI22_X1 U23668 ( .A1(n20810), .A2(n20714), .B1(n20809), .B2(n20713), .ZN(
        n20712) );
  AOI22_X1 U23669 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20715), .B1(
        n20756), .B2(n20811), .ZN(n20711) );
  OAI211_X1 U23670 ( .C1(n20814), .C2(n20718), .A(n20712), .B(n20711), .ZN(
        P1_U3143) );
  AOI22_X1 U23671 ( .A1(n20818), .A2(n20714), .B1(n20816), .B2(n20713), .ZN(
        n20717) );
  AOI22_X1 U23672 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20715), .B1(
        n20756), .B2(n20819), .ZN(n20716) );
  OAI211_X1 U23673 ( .C1(n20825), .C2(n20718), .A(n20717), .B(n20716), .ZN(
        P1_U3144) );
  NAND2_X1 U23674 ( .A1(n20726), .A2(n20598), .ZN(n20722) );
  OAI22_X1 U23675 ( .A1(n20723), .A2(n20722), .B1(n20721), .B2(n20720), .ZN(
        n20754) );
  NOR2_X1 U23676 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20763), .ZN(
        n20753) );
  AOI22_X1 U23677 ( .A1(n20765), .A2(n20754), .B1(n20764), .B2(n20753), .ZN(
        n20732) );
  AOI21_X1 U23678 ( .B1(n20824), .B2(n20724), .A(n21280), .ZN(n20725) );
  AOI21_X1 U23679 ( .B1(n20762), .B2(n20726), .A(n20725), .ZN(n20727) );
  NOR2_X1 U23680 ( .A1(n20727), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20730) );
  AOI22_X1 U23681 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20757), .B1(
        n20756), .B2(n20773), .ZN(n20731) );
  OAI211_X1 U23682 ( .C1(n20776), .C2(n20824), .A(n20732), .B(n20731), .ZN(
        P1_U3145) );
  AOI22_X1 U23683 ( .A1(n20778), .A2(n20754), .B1(n20777), .B2(n20753), .ZN(
        n20734) );
  AOI22_X1 U23684 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20757), .B1(
        n20756), .B2(n20779), .ZN(n20733) );
  OAI211_X1 U23685 ( .C1(n20782), .C2(n20824), .A(n20734), .B(n20733), .ZN(
        P1_U3146) );
  AOI22_X1 U23686 ( .A1(n20784), .A2(n20754), .B1(n20783), .B2(n20753), .ZN(
        n20737) );
  AOI22_X1 U23687 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20757), .B1(
        n20756), .B2(n20735), .ZN(n20736) );
  OAI211_X1 U23688 ( .C1(n20738), .C2(n20824), .A(n20737), .B(n20736), .ZN(
        P1_U3147) );
  AOI22_X1 U23689 ( .A1(n20790), .A2(n20754), .B1(n20789), .B2(n20753), .ZN(
        n20741) );
  AOI22_X1 U23690 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20757), .B1(
        n20756), .B2(n20739), .ZN(n20740) );
  OAI211_X1 U23691 ( .C1(n20742), .C2(n20824), .A(n20741), .B(n20740), .ZN(
        P1_U3148) );
  AOI22_X1 U23692 ( .A1(n20796), .A2(n20754), .B1(n20795), .B2(n20753), .ZN(
        n20745) );
  AOI22_X1 U23693 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20757), .B1(
        n20756), .B2(n20743), .ZN(n20744) );
  OAI211_X1 U23694 ( .C1(n20746), .C2(n20824), .A(n20745), .B(n20744), .ZN(
        P1_U3149) );
  AOI22_X1 U23695 ( .A1(n20802), .A2(n20754), .B1(n20801), .B2(n20753), .ZN(
        n20748) );
  AOI22_X1 U23696 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20757), .B1(
        n20756), .B2(n20803), .ZN(n20747) );
  OAI211_X1 U23697 ( .C1(n20808), .C2(n20824), .A(n20748), .B(n20747), .ZN(
        P1_U3150) );
  AOI22_X1 U23698 ( .A1(n20810), .A2(n20754), .B1(n20809), .B2(n20753), .ZN(
        n20751) );
  AOI22_X1 U23699 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20757), .B1(
        n20756), .B2(n20749), .ZN(n20750) );
  OAI211_X1 U23700 ( .C1(n20752), .C2(n20824), .A(n20751), .B(n20750), .ZN(
        P1_U3151) );
  AOI22_X1 U23701 ( .A1(n20818), .A2(n20754), .B1(n20816), .B2(n20753), .ZN(
        n20759) );
  AOI22_X1 U23702 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20757), .B1(
        n20756), .B2(n20755), .ZN(n20758) );
  OAI211_X1 U23703 ( .C1(n20760), .C2(n20824), .A(n20759), .B(n20758), .ZN(
        P1_U3152) );
  AOI21_X1 U23704 ( .B1(n20762), .B2(n20761), .A(n20815), .ZN(n20767) );
  OAI22_X1 U23705 ( .A1(n20767), .A2(n12580), .B1(n20763), .B2(n20898), .ZN(
        n20817) );
  AOI22_X1 U23706 ( .A1(n20765), .A2(n20817), .B1(n20764), .B2(n20815), .ZN(
        n20775) );
  NAND2_X1 U23707 ( .A1(n20766), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20768) );
  OAI21_X1 U23708 ( .B1(n20769), .B2(n20768), .A(n20767), .ZN(n20771) );
  OAI221_X1 U23709 ( .B1(n20598), .B2(n20772), .C1(n12580), .C2(n20771), .A(
        n20770), .ZN(n20821) );
  INV_X1 U23710 ( .A(n20824), .ZN(n20804) );
  AOI22_X1 U23711 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20821), .B1(
        n20804), .B2(n20773), .ZN(n20774) );
  OAI211_X1 U23712 ( .C1(n20776), .C2(n20807), .A(n20775), .B(n20774), .ZN(
        P1_U3153) );
  AOI22_X1 U23713 ( .A1(n20778), .A2(n20817), .B1(n20777), .B2(n20815), .ZN(
        n20781) );
  AOI22_X1 U23714 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20821), .B1(
        n20804), .B2(n20779), .ZN(n20780) );
  OAI211_X1 U23715 ( .C1(n20782), .C2(n20807), .A(n20781), .B(n20780), .ZN(
        P1_U3154) );
  AOI22_X1 U23716 ( .A1(n20784), .A2(n20817), .B1(n20783), .B2(n20815), .ZN(
        n20787) );
  AOI22_X1 U23717 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20821), .B1(
        n20820), .B2(n20785), .ZN(n20786) );
  OAI211_X1 U23718 ( .C1(n20788), .C2(n20824), .A(n20787), .B(n20786), .ZN(
        P1_U3155) );
  AOI22_X1 U23719 ( .A1(n20790), .A2(n20817), .B1(n20789), .B2(n20815), .ZN(
        n20793) );
  AOI22_X1 U23720 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20821), .B1(
        n20820), .B2(n20791), .ZN(n20792) );
  OAI211_X1 U23721 ( .C1(n20794), .C2(n20824), .A(n20793), .B(n20792), .ZN(
        P1_U3156) );
  AOI22_X1 U23722 ( .A1(n20796), .A2(n20817), .B1(n20795), .B2(n20815), .ZN(
        n20799) );
  AOI22_X1 U23723 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20821), .B1(
        n20820), .B2(n20797), .ZN(n20798) );
  OAI211_X1 U23724 ( .C1(n20800), .C2(n20824), .A(n20799), .B(n20798), .ZN(
        P1_U3157) );
  AOI22_X1 U23725 ( .A1(n20802), .A2(n20817), .B1(n20801), .B2(n20815), .ZN(
        n20806) );
  AOI22_X1 U23726 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20821), .B1(
        n20804), .B2(n20803), .ZN(n20805) );
  OAI211_X1 U23727 ( .C1(n20808), .C2(n20807), .A(n20806), .B(n20805), .ZN(
        P1_U3158) );
  AOI22_X1 U23728 ( .A1(n20810), .A2(n20817), .B1(n20809), .B2(n20815), .ZN(
        n20813) );
  AOI22_X1 U23729 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20821), .B1(
        n20820), .B2(n20811), .ZN(n20812) );
  OAI211_X1 U23730 ( .C1(n20814), .C2(n20824), .A(n20813), .B(n20812), .ZN(
        P1_U3159) );
  AOI22_X1 U23731 ( .A1(n20818), .A2(n20817), .B1(n20816), .B2(n20815), .ZN(
        n20823) );
  AOI22_X1 U23732 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20821), .B1(
        n20820), .B2(n20819), .ZN(n20822) );
  OAI211_X1 U23733 ( .C1(n20825), .C2(n20824), .A(n20823), .B(n20822), .ZN(
        P1_U3160) );
  OAI211_X1 U23734 ( .C1(n20828), .C2(n20898), .A(n20827), .B(n20826), .ZN(
        P1_U3163) );
  AND2_X1 U23735 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20829), .ZN(
        P1_U3164) );
  AND2_X1 U23736 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20829), .ZN(
        P1_U3165) );
  AND2_X1 U23737 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20829), .ZN(
        P1_U3166) );
  AND2_X1 U23738 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20829), .ZN(
        P1_U3167) );
  AND2_X1 U23739 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20829), .ZN(
        P1_U3168) );
  AND2_X1 U23740 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20829), .ZN(
        P1_U3169) );
  AND2_X1 U23741 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20829), .ZN(
        P1_U3170) );
  AND2_X1 U23742 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20829), .ZN(
        P1_U3171) );
  AND2_X1 U23743 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20829), .ZN(
        P1_U3172) );
  AND2_X1 U23744 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20829), .ZN(
        P1_U3173) );
  AND2_X1 U23745 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20829), .ZN(
        P1_U3174) );
  AND2_X1 U23746 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20829), .ZN(
        P1_U3175) );
  AND2_X1 U23747 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20829), .ZN(
        P1_U3176) );
  AND2_X1 U23748 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20829), .ZN(
        P1_U3177) );
  AND2_X1 U23749 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20829), .ZN(
        P1_U3178) );
  AND2_X1 U23750 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20829), .ZN(
        P1_U3179) );
  AND2_X1 U23751 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20829), .ZN(
        P1_U3180) );
  AND2_X1 U23752 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20829), .ZN(
        P1_U3181) );
  AND2_X1 U23753 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20829), .ZN(
        P1_U3182) );
  AND2_X1 U23754 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20829), .ZN(
        P1_U3183) );
  AND2_X1 U23755 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20829), .ZN(
        P1_U3184) );
  AND2_X1 U23756 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20829), .ZN(
        P1_U3185) );
  AND2_X1 U23757 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20829), .ZN(P1_U3186) );
  AND2_X1 U23758 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20829), .ZN(P1_U3187) );
  AND2_X1 U23759 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20829), .ZN(P1_U3188) );
  AND2_X1 U23760 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20829), .ZN(P1_U3189) );
  AND2_X1 U23761 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20829), .ZN(P1_U3190) );
  AND2_X1 U23762 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20829), .ZN(P1_U3191) );
  AND2_X1 U23763 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20829), .ZN(P1_U3192) );
  AND2_X1 U23764 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20829), .ZN(P1_U3193) );
  NAND2_X1 U23765 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20836), .ZN(n20839) );
  INV_X1 U23766 ( .A(n20839), .ZN(n20833) );
  INV_X1 U23767 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21216) );
  OAI22_X1 U23768 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21180), .B1(n20834), 
        .B2(n21232), .ZN(n20830) );
  NOR3_X1 U23769 ( .A1(n20831), .A2(n21216), .A3(n20830), .ZN(n20832) );
  OAI22_X1 U23770 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20833), .B1(n20909), 
        .B2(n20832), .ZN(P1_U3194) );
  AOI211_X1 U23771 ( .C1(n20835), .C2(n21180), .A(P1_STATE_REG_2__SCAN_IN), 
        .B(n20834), .ZN(n20842) );
  AOI21_X1 U23772 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(n20843), .A(n21232), .ZN(n20838) );
  INV_X1 U23773 ( .A(n20836), .ZN(n20837) );
  OAI221_X1 U23774 ( .B1(n20838), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .C1(
        n20838), .C2(n20837), .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20841) );
  OAI211_X1 U23775 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n21180), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n20839), .ZN(n20840) );
  OAI21_X1 U23776 ( .B1(n20842), .B2(n20841), .A(n20840), .ZN(P1_U3196) );
  OR2_X1 U23777 ( .A1(n20876), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20853) );
  INV_X2 U23778 ( .A(n20853), .ZN(n20877) );
  NOR2_X1 U23779 ( .A1(n20843), .A2(n20876), .ZN(n20872) );
  INV_X1 U23780 ( .A(n20872), .ZN(n20851) );
  INV_X1 U23781 ( .A(n20851), .ZN(n20879) );
  AOI222_X1 U23782 ( .A1(n20877), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n20876), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n20879), .ZN(n20844) );
  INV_X1 U23783 ( .A(n20844), .ZN(P1_U3197) );
  AOI222_X1 U23784 ( .A1(n20879), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20876), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20877), .ZN(n20845) );
  INV_X1 U23785 ( .A(n20845), .ZN(P1_U3198) );
  OAI222_X1 U23786 ( .A1(n20851), .A2(n21230), .B1(n20847), .B2(n20909), .C1(
        n20846), .C2(n20853), .ZN(P1_U3199) );
  AOI222_X1 U23787 ( .A1(n20877), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20876), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20872), .ZN(n20848) );
  INV_X1 U23788 ( .A(n20848), .ZN(P1_U3200) );
  AOI222_X1 U23789 ( .A1(n20879), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20876), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20877), .ZN(n20849) );
  INV_X1 U23790 ( .A(n20849), .ZN(P1_U3201) );
  AOI22_X1 U23791 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n20876), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20877), .ZN(n20850) );
  OAI21_X1 U23792 ( .B1(n21235), .B2(n20851), .A(n20850), .ZN(P1_U3202) );
  AOI22_X1 U23793 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n20876), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20872), .ZN(n20852) );
  OAI21_X1 U23794 ( .B1(n21208), .B2(n20853), .A(n20852), .ZN(P1_U3203) );
  AOI222_X1 U23795 ( .A1(n20879), .A2(P1_REIP_REG_8__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20876), .C1(P1_REIP_REG_9__SCAN_IN), 
        .C2(n20877), .ZN(n20854) );
  INV_X1 U23796 ( .A(n20854), .ZN(P1_U3204) );
  AOI222_X1 U23797 ( .A1(n20879), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20876), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20877), .ZN(n20855) );
  INV_X1 U23798 ( .A(n20855), .ZN(P1_U3205) );
  AOI222_X1 U23799 ( .A1(n20877), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20876), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20879), .ZN(n20856) );
  INV_X1 U23800 ( .A(n20856), .ZN(P1_U3206) );
  AOI222_X1 U23801 ( .A1(n20879), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20876), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20877), .ZN(n20857) );
  INV_X1 U23802 ( .A(n20857), .ZN(P1_U3207) );
  AOI222_X1 U23803 ( .A1(n20879), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20876), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n20877), .ZN(n20858) );
  INV_X1 U23804 ( .A(n20858), .ZN(P1_U3208) );
  AOI222_X1 U23805 ( .A1(n20879), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n20876), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20877), .ZN(n20859) );
  INV_X1 U23806 ( .A(n20859), .ZN(P1_U3209) );
  AOI222_X1 U23807 ( .A1(n20877), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20876), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20879), .ZN(n20860) );
  INV_X1 U23808 ( .A(n20860), .ZN(P1_U3210) );
  AOI222_X1 U23809 ( .A1(n20879), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20876), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20877), .ZN(n20861) );
  INV_X1 U23810 ( .A(n20861), .ZN(P1_U3211) );
  AOI222_X1 U23811 ( .A1(n20872), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n20876), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n20877), .ZN(n20862) );
  INV_X1 U23812 ( .A(n20862), .ZN(P1_U3212) );
  AOI222_X1 U23813 ( .A1(n20872), .A2(P1_REIP_REG_17__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n20876), .C1(P1_REIP_REG_18__SCAN_IN), 
        .C2(n20877), .ZN(n20863) );
  INV_X1 U23814 ( .A(n20863), .ZN(P1_U3213) );
  AOI222_X1 U23815 ( .A1(n20877), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20876), .C1(P1_REIP_REG_18__SCAN_IN), 
        .C2(n20879), .ZN(n20864) );
  INV_X1 U23816 ( .A(n20864), .ZN(P1_U3214) );
  AOI222_X1 U23817 ( .A1(n20877), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n20876), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20879), .ZN(n20865) );
  INV_X1 U23818 ( .A(n20865), .ZN(P1_U3215) );
  AOI222_X1 U23819 ( .A1(n20872), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n20876), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20877), .ZN(n20866) );
  INV_X1 U23820 ( .A(n20866), .ZN(P1_U3216) );
  AOI222_X1 U23821 ( .A1(n20872), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20876), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n20877), .ZN(n20867) );
  INV_X1 U23822 ( .A(n20867), .ZN(P1_U3217) );
  AOI222_X1 U23823 ( .A1(n20872), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n20876), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20877), .ZN(n20868) );
  INV_X1 U23824 ( .A(n20868), .ZN(P1_U3218) );
  AOI222_X1 U23825 ( .A1(n20879), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20876), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n20877), .ZN(n20869) );
  INV_X1 U23826 ( .A(n20869), .ZN(P1_U3219) );
  AOI222_X1 U23827 ( .A1(n20872), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20876), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20877), .ZN(n20870) );
  INV_X1 U23828 ( .A(n20870), .ZN(P1_U3220) );
  AOI222_X1 U23829 ( .A1(n20879), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20876), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20877), .ZN(n20871) );
  INV_X1 U23830 ( .A(n20871), .ZN(P1_U3221) );
  AOI222_X1 U23831 ( .A1(n20872), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20876), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20877), .ZN(n20873) );
  INV_X1 U23832 ( .A(n20873), .ZN(P1_U3222) );
  AOI222_X1 U23833 ( .A1(n20879), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20876), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20877), .ZN(n20874) );
  INV_X1 U23834 ( .A(n20874), .ZN(P1_U3223) );
  AOI222_X1 U23835 ( .A1(n20879), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20876), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20877), .ZN(n20875) );
  INV_X1 U23836 ( .A(n20875), .ZN(P1_U3224) );
  AOI222_X1 U23837 ( .A1(n20877), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20876), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20879), .ZN(n20878) );
  INV_X1 U23838 ( .A(n20878), .ZN(P1_U3225) );
  AOI222_X1 U23839 ( .A1(n20879), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20876), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20877), .ZN(n20880) );
  INV_X1 U23840 ( .A(n20880), .ZN(P1_U3226) );
  OAI22_X1 U23841 ( .A1(n20876), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20909), .ZN(n20881) );
  INV_X1 U23842 ( .A(n20881), .ZN(P1_U3458) );
  OAI22_X1 U23843 ( .A1(n20876), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20909), .ZN(n20882) );
  INV_X1 U23844 ( .A(n20882), .ZN(P1_U3459) );
  OAI22_X1 U23845 ( .A1(n20876), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20909), .ZN(n20883) );
  INV_X1 U23846 ( .A(n20883), .ZN(P1_U3460) );
  OAI22_X1 U23847 ( .A1(n20876), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20909), .ZN(n20884) );
  INV_X1 U23848 ( .A(n20884), .ZN(P1_U3461) );
  OAI21_X1 U23849 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20888), .A(n20886), 
        .ZN(n20885) );
  INV_X1 U23850 ( .A(n20885), .ZN(P1_U3464) );
  OAI21_X1 U23851 ( .B1(n20888), .B2(n20887), .A(n20886), .ZN(P1_U3465) );
  AOI21_X1 U23852 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20890) );
  AOI22_X1 U23853 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20890), .B2(n20889), .ZN(n20892) );
  INV_X1 U23854 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20891) );
  AOI22_X1 U23855 ( .A1(n20893), .A2(n20892), .B1(n20891), .B2(n20895), .ZN(
        P1_U3481) );
  INV_X1 U23856 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20896) );
  INV_X1 U23857 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n21162) );
  NOR2_X1 U23858 ( .A1(n20895), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20894) );
  AOI22_X1 U23859 ( .A1(n20896), .A2(n20895), .B1(n21162), .B2(n20894), .ZN(
        P1_U3482) );
  OAI22_X1 U23860 ( .A1(n20876), .A2(n21170), .B1(P1_W_R_N_REG_SCAN_IN), .B2(
        n20909), .ZN(n20897) );
  INV_X1 U23861 ( .A(n20897), .ZN(P1_U3483) );
  NOR3_X1 U23862 ( .A1(n20900), .A2(n20899), .A3(n20898), .ZN(n20903) );
  OAI21_X1 U23863 ( .B1(n20903), .B2(n20902), .A(n20901), .ZN(n20908) );
  AOI211_X1 U23864 ( .C1(n20132), .C2(n20906), .A(n20905), .B(n20904), .ZN(
        n20907) );
  MUX2_X1 U23865 ( .A(n20908), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n20907), 
        .Z(P1_U3485) );
  AOI22_X1 U23866 ( .A1(n20909), .A2(n21181), .B1(n21241), .B2(n20876), .ZN(
        P1_U3486) );
  AOI22_X1 U23867 ( .A1(n16548), .A2(P3_ADDRESS_REG_29__SCAN_IN), .B1(
        P2_ADDRESS_REG_29__SCAN_IN), .B2(n16550), .ZN(n21303) );
  OAI22_X1 U23868 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(keyinput_g56), .B1(
        keyinput_g7), .B2(DATAI_25_), .ZN(n20910) );
  AOI221_X1 U23869 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(keyinput_g56), .C1(
        DATAI_25_), .C2(keyinput_g7), .A(n20910), .ZN(n20917) );
  OAI22_X1 U23870 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(keyinput_g110), .B1(
        P1_REIP_REG_25__SCAN_IN), .B2(keyinput_g58), .ZN(n20911) );
  AOI221_X1 U23871 ( .B1(P1_EBX_REG_5__SCAN_IN), .B2(keyinput_g110), .C1(
        keyinput_g58), .C2(P1_REIP_REG_25__SCAN_IN), .A(n20911), .ZN(n20916)
         );
  OAI22_X1 U23872 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(keyinput_g83), .B1(BS16), 
        .B2(keyinput_g35), .ZN(n20912) );
  AOI221_X1 U23873 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(keyinput_g83), .C1(
        keyinput_g35), .C2(BS16), .A(n20912), .ZN(n20915) );
  OAI22_X1 U23874 ( .A1(P1_EBX_REG_29__SCAN_IN), .A2(keyinput_g86), .B1(
        keyinput_g88), .B2(P1_EBX_REG_27__SCAN_IN), .ZN(n20913) );
  AOI221_X1 U23875 ( .B1(P1_EBX_REG_29__SCAN_IN), .B2(keyinput_g86), .C1(
        P1_EBX_REG_27__SCAN_IN), .C2(keyinput_g88), .A(n20913), .ZN(n20914) );
  NAND4_X1 U23876 ( .A1(n20917), .A2(n20916), .A3(n20915), .A4(n20914), .ZN(
        n21051) );
  OAI22_X1 U23877 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(keyinput_g65), .B1(
        keyinput_g11), .B2(DATAI_21_), .ZN(n20918) );
  AOI221_X1 U23878 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(keyinput_g65), .C1(
        DATAI_21_), .C2(keyinput_g11), .A(n20918), .ZN(n20943) );
  OAI22_X1 U23879 ( .A1(P1_EBX_REG_15__SCAN_IN), .A2(keyinput_g100), .B1(
        keyinput_g3), .B2(DATAI_29_), .ZN(n20919) );
  AOI221_X1 U23880 ( .B1(P1_EBX_REG_15__SCAN_IN), .B2(keyinput_g100), .C1(
        DATAI_29_), .C2(keyinput_g3), .A(n20919), .ZN(n20922) );
  OAI22_X1 U23881 ( .A1(P1_EBX_REG_1__SCAN_IN), .A2(keyinput_g114), .B1(
        P1_EBX_REG_11__SCAN_IN), .B2(keyinput_g104), .ZN(n20920) );
  AOI221_X1 U23882 ( .B1(P1_EBX_REG_1__SCAN_IN), .B2(keyinput_g114), .C1(
        keyinput_g104), .C2(P1_EBX_REG_11__SCAN_IN), .A(n20920), .ZN(n20921)
         );
  OAI211_X1 U23883 ( .C1(n21216), .C2(keyinput_g43), .A(n20922), .B(n20921), 
        .ZN(n20923) );
  AOI21_X1 U23884 ( .B1(n21216), .B2(keyinput_g43), .A(n20923), .ZN(n20942) );
  AOI22_X1 U23885 ( .A1(P1_W_R_N_REG_SCAN_IN), .A2(keyinput_g47), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(keyinput_g75), .ZN(n20924) );
  OAI221_X1 U23886 ( .B1(P1_W_R_N_REG_SCAN_IN), .B2(keyinput_g47), .C1(
        P1_REIP_REG_8__SCAN_IN), .C2(keyinput_g75), .A(n20924), .ZN(n20931) );
  AOI22_X1 U23887 ( .A1(DATAI_2_), .A2(keyinput_g30), .B1(DATAI_24_), .B2(
        keyinput_g8), .ZN(n20925) );
  OAI221_X1 U23888 ( .B1(DATAI_2_), .B2(keyinput_g30), .C1(DATAI_24_), .C2(
        keyinput_g8), .A(n20925), .ZN(n20930) );
  AOI22_X1 U23889 ( .A1(DATAI_15_), .A2(keyinput_g17), .B1(
        P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_g44), .ZN(n20926) );
  OAI221_X1 U23890 ( .B1(DATAI_15_), .B2(keyinput_g17), .C1(
        P1_STATEBS16_REG_SCAN_IN), .C2(keyinput_g44), .A(n20926), .ZN(n20929)
         );
  AOI22_X1 U23891 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(keyinput_g76), .B1(
        P1_EBX_REG_26__SCAN_IN), .B2(keyinput_g89), .ZN(n20927) );
  OAI221_X1 U23892 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(keyinput_g76), .C1(
        P1_EBX_REG_26__SCAN_IN), .C2(keyinput_g89), .A(n20927), .ZN(n20928) );
  NOR4_X1 U23893 ( .A1(n20931), .A2(n20930), .A3(n20929), .A4(n20928), .ZN(
        n20941) );
  AOI22_X1 U23894 ( .A1(DATAI_4_), .A2(keyinput_g28), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(keyinput_g85), .ZN(n20932) );
  OAI221_X1 U23895 ( .B1(DATAI_4_), .B2(keyinput_g28), .C1(
        P1_EBX_REG_30__SCAN_IN), .C2(keyinput_g85), .A(n20932), .ZN(n20939) );
  AOI22_X1 U23896 ( .A1(DATAI_19_), .A2(keyinput_g13), .B1(
        P1_EBX_REG_31__SCAN_IN), .B2(keyinput_g84), .ZN(n20933) );
  OAI221_X1 U23897 ( .B1(DATAI_19_), .B2(keyinput_g13), .C1(
        P1_EBX_REG_31__SCAN_IN), .C2(keyinput_g84), .A(n20933), .ZN(n20938) );
  AOI22_X1 U23898 ( .A1(P1_BYTEENABLE_REG_0__SCAN_IN), .A2(keyinput_g48), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(keyinput_g120), .ZN(n20934) );
  OAI221_X1 U23899 ( .B1(P1_BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_g48), 
        .C1(P1_EAX_REG_27__SCAN_IN), .C2(keyinput_g120), .A(n20934), .ZN(
        n20937) );
  AOI22_X1 U23900 ( .A1(P1_EBX_REG_10__SCAN_IN), .A2(keyinput_g105), .B1(
        P1_EBX_REG_9__SCAN_IN), .B2(keyinput_g106), .ZN(n20935) );
  OAI221_X1 U23901 ( .B1(P1_EBX_REG_10__SCAN_IN), .B2(keyinput_g105), .C1(
        P1_EBX_REG_9__SCAN_IN), .C2(keyinput_g106), .A(n20935), .ZN(n20936) );
  NOR4_X1 U23902 ( .A1(n20939), .A2(n20938), .A3(n20937), .A4(n20936), .ZN(
        n20940) );
  NAND4_X1 U23903 ( .A1(n20943), .A2(n20942), .A3(n20941), .A4(n20940), .ZN(
        n21050) );
  INV_X1 U23904 ( .A(DATAI_0_), .ZN(n20946) );
  AOI22_X1 U23905 ( .A1(n20946), .A2(keyinput_g32), .B1(n20945), .B2(
        keyinput_g15), .ZN(n20944) );
  OAI221_X1 U23906 ( .B1(n20946), .B2(keyinput_g32), .C1(n20945), .C2(
        keyinput_g15), .A(n20944), .ZN(n20957) );
  AOI22_X1 U23907 ( .A1(n21256), .A2(keyinput_g127), .B1(keyinput_g109), .B2(
        n20948), .ZN(n20947) );
  OAI221_X1 U23908 ( .B1(n21256), .B2(keyinput_g127), .C1(n20948), .C2(
        keyinput_g109), .A(n20947), .ZN(n20956) );
  INV_X1 U23909 ( .A(DATAI_14_), .ZN(n20951) );
  AOI22_X1 U23910 ( .A1(n20951), .A2(keyinput_g18), .B1(n20950), .B2(
        keyinput_g62), .ZN(n20949) );
  OAI221_X1 U23911 ( .B1(n20951), .B2(keyinput_g18), .C1(n20950), .C2(
        keyinput_g62), .A(n20949), .ZN(n20955) );
  AOI22_X1 U23912 ( .A1(n20953), .A2(keyinput_g118), .B1(keyinput_g74), .B2(
        n13635), .ZN(n20952) );
  OAI221_X1 U23913 ( .B1(n20953), .B2(keyinput_g118), .C1(n13635), .C2(
        keyinput_g74), .A(n20952), .ZN(n20954) );
  NOR4_X1 U23914 ( .A1(n20957), .A2(n20956), .A3(n20955), .A4(n20954), .ZN(
        n20996) );
  AOI22_X1 U23915 ( .A1(n21170), .A2(keyinput_g38), .B1(n20959), .B2(
        keyinput_g97), .ZN(n20958) );
  OAI221_X1 U23916 ( .B1(n21170), .B2(keyinput_g38), .C1(n20959), .C2(
        keyinput_g97), .A(n20958), .ZN(n20970) );
  INV_X1 U23917 ( .A(DATAI_9_), .ZN(n20961) );
  AOI22_X1 U23918 ( .A1(n20962), .A2(keyinput_g49), .B1(n20961), .B2(
        keyinput_g23), .ZN(n20960) );
  OAI221_X1 U23919 ( .B1(n20962), .B2(keyinput_g49), .C1(n20961), .C2(
        keyinput_g23), .A(n20960), .ZN(n20969) );
  INV_X1 U23920 ( .A(DATAI_3_), .ZN(n21245) );
  INV_X1 U23921 ( .A(DATAI_10_), .ZN(n20964) );
  AOI22_X1 U23922 ( .A1(n21245), .A2(keyinput_g29), .B1(n20964), .B2(
        keyinput_g22), .ZN(n20963) );
  OAI221_X1 U23923 ( .B1(n21245), .B2(keyinput_g29), .C1(n20964), .C2(
        keyinput_g22), .A(n20963), .ZN(n20968) );
  INV_X1 U23924 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n20966) );
  AOI22_X1 U23925 ( .A1(n20966), .A2(keyinput_g71), .B1(n21187), .B2(
        keyinput_g123), .ZN(n20965) );
  OAI221_X1 U23926 ( .B1(n20966), .B2(keyinput_g71), .C1(n21187), .C2(
        keyinput_g123), .A(n20965), .ZN(n20967) );
  NOR4_X1 U23927 ( .A1(n20970), .A2(n20969), .A3(n20968), .A4(n20967), .ZN(
        n20995) );
  AOI22_X1 U23928 ( .A1(n20972), .A2(keyinput_g103), .B1(keyinput_g10), .B2(
        n21207), .ZN(n20971) );
  OAI221_X1 U23929 ( .B1(n20972), .B2(keyinput_g103), .C1(n21207), .C2(
        keyinput_g10), .A(n20971), .ZN(n20980) );
  AOI22_X1 U23930 ( .A1(n21183), .A2(keyinput_g53), .B1(keyinput_g59), .B2(
        n21198), .ZN(n20973) );
  OAI221_X1 U23931 ( .B1(n21183), .B2(keyinput_g53), .C1(n21198), .C2(
        keyinput_g59), .A(n20973), .ZN(n20979) );
  AOI22_X1 U23932 ( .A1(n12796), .A2(keyinput_g115), .B1(n20975), .B2(
        keyinput_g117), .ZN(n20974) );
  OAI221_X1 U23933 ( .B1(n12796), .B2(keyinput_g115), .C1(n20975), .C2(
        keyinput_g117), .A(n20974), .ZN(n20978) );
  INV_X1 U23934 ( .A(DATAI_1_), .ZN(n21229) );
  AOI22_X1 U23935 ( .A1(n21171), .A2(keyinput_g63), .B1(keyinput_g31), .B2(
        n21229), .ZN(n20976) );
  OAI221_X1 U23936 ( .B1(n21171), .B2(keyinput_g63), .C1(n21229), .C2(
        keyinput_g31), .A(n20976), .ZN(n20977) );
  NOR4_X1 U23937 ( .A1(n20980), .A2(n20979), .A3(n20978), .A4(n20977), .ZN(
        n20994) );
  AOI22_X1 U23938 ( .A1(n20982), .A2(keyinput_g70), .B1(keyinput_g34), .B2(
        n21180), .ZN(n20981) );
  OAI221_X1 U23939 ( .B1(n20982), .B2(keyinput_g70), .C1(n21180), .C2(
        keyinput_g34), .A(n20981), .ZN(n20992) );
  AOI22_X1 U23940 ( .A1(n20984), .A2(keyinput_g126), .B1(keyinput_g121), .B2(
        n21215), .ZN(n20983) );
  OAI221_X1 U23941 ( .B1(n20984), .B2(keyinput_g126), .C1(n21215), .C2(
        keyinput_g121), .A(n20983), .ZN(n20991) );
  AOI22_X1 U23942 ( .A1(n20986), .A2(keyinput_g42), .B1(n21279), .B2(
        keyinput_g122), .ZN(n20985) );
  OAI221_X1 U23943 ( .B1(n20986), .B2(keyinput_g42), .C1(n21279), .C2(
        keyinput_g122), .A(n20985), .ZN(n20990) );
  AOI22_X1 U23944 ( .A1(n20988), .A2(keyinput_g68), .B1(n21195), .B2(
        keyinput_g72), .ZN(n20987) );
  OAI221_X1 U23945 ( .B1(n20988), .B2(keyinput_g68), .C1(n21195), .C2(
        keyinput_g72), .A(n20987), .ZN(n20989) );
  NOR4_X1 U23946 ( .A1(n20992), .A2(n20991), .A3(n20990), .A4(n20989), .ZN(
        n20993) );
  NAND4_X1 U23947 ( .A1(n20996), .A2(n20995), .A3(n20994), .A4(n20993), .ZN(
        n21049) );
  INV_X1 U23948 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n20998) );
  AOI22_X1 U23949 ( .A1(n20999), .A2(keyinput_g91), .B1(keyinput_g102), .B2(
        n20998), .ZN(n20997) );
  OAI221_X1 U23950 ( .B1(n20999), .B2(keyinput_g91), .C1(n20998), .C2(
        keyinput_g102), .A(n20997), .ZN(n21008) );
  AOI22_X1 U23951 ( .A1(n21001), .A2(keyinput_g16), .B1(keyinput_g39), .B2(
        n21199), .ZN(n21000) );
  OAI221_X1 U23952 ( .B1(n21001), .B2(keyinput_g16), .C1(n21199), .C2(
        keyinput_g39), .A(n21000), .ZN(n21007) );
  AOI22_X1 U23953 ( .A1(n21003), .A2(keyinput_g9), .B1(n21201), .B2(
        keyinput_g108), .ZN(n21002) );
  OAI221_X1 U23954 ( .B1(n21003), .B2(keyinput_g9), .C1(n21201), .C2(
        keyinput_g108), .A(n21002), .ZN(n21006) );
  AOI22_X1 U23955 ( .A1(n21235), .A2(keyinput_g77), .B1(n21227), .B2(
        keyinput_g55), .ZN(n21004) );
  OAI221_X1 U23956 ( .B1(n21235), .B2(keyinput_g77), .C1(n21227), .C2(
        keyinput_g55), .A(n21004), .ZN(n21005) );
  NOR4_X1 U23957 ( .A1(n21008), .A2(n21007), .A3(n21006), .A4(n21005), .ZN(
        n21047) );
  INV_X1 U23958 ( .A(P1_EAX_REG_31__SCAN_IN), .ZN(n21010) );
  AOI22_X1 U23959 ( .A1(n21010), .A2(keyinput_g116), .B1(keyinput_g2), .B2(
        n21251), .ZN(n21009) );
  OAI221_X1 U23960 ( .B1(n21010), .B2(keyinput_g116), .C1(n21251), .C2(
        keyinput_g2), .A(n21009), .ZN(n21020) );
  INV_X1 U23961 ( .A(READY2), .ZN(n21012) );
  AOI22_X1 U23962 ( .A1(n21012), .A2(keyinput_g37), .B1(keyinput_g0), .B2(
        n21181), .ZN(n21011) );
  OAI221_X1 U23963 ( .B1(n21012), .B2(keyinput_g37), .C1(n21181), .C2(
        keyinput_g0), .A(n21011), .ZN(n21019) );
  AOI22_X1 U23964 ( .A1(n21167), .A2(keyinput_g6), .B1(n21014), .B2(
        keyinput_g67), .ZN(n21013) );
  OAI221_X1 U23965 ( .B1(n21167), .B2(keyinput_g6), .C1(n21014), .C2(
        keyinput_g67), .A(n21013), .ZN(n21018) );
  AOI22_X1 U23966 ( .A1(n21016), .A2(keyinput_g69), .B1(n14512), .B2(
        keyinput_g64), .ZN(n21015) );
  OAI221_X1 U23967 ( .B1(n21016), .B2(keyinput_g69), .C1(n14512), .C2(
        keyinput_g64), .A(n21015), .ZN(n21017) );
  NOR4_X1 U23968 ( .A1(n21020), .A2(n21019), .A3(n21018), .A4(n21017), .ZN(
        n21046) );
  AOI22_X1 U23969 ( .A1(n21274), .A2(keyinput_g4), .B1(keyinput_g46), .B2(
        n21022), .ZN(n21021) );
  OAI221_X1 U23970 ( .B1(n21274), .B2(keyinput_g4), .C1(n21022), .C2(
        keyinput_g46), .A(n21021), .ZN(n21031) );
  INV_X1 U23971 ( .A(DATAI_12_), .ZN(n21024) );
  AOI22_X1 U23972 ( .A1(n21024), .A2(keyinput_g20), .B1(n21244), .B2(
        keyinput_g125), .ZN(n21023) );
  OAI221_X1 U23973 ( .B1(n21024), .B2(keyinput_g20), .C1(n21244), .C2(
        keyinput_g125), .A(n21023), .ZN(n21030) );
  AOI22_X1 U23974 ( .A1(n21026), .A2(keyinput_g73), .B1(n21236), .B2(
        keyinput_g101), .ZN(n21025) );
  OAI221_X1 U23975 ( .B1(n21026), .B2(keyinput_g73), .C1(n21236), .C2(
        keyinput_g101), .A(n21025), .ZN(n21029) );
  AOI22_X1 U23976 ( .A1(n21165), .A2(keyinput_g81), .B1(n21230), .B2(
        keyinput_g80), .ZN(n21027) );
  OAI221_X1 U23977 ( .B1(n21165), .B2(keyinput_g81), .C1(n21230), .C2(
        keyinput_g80), .A(n21027), .ZN(n21028) );
  NOR4_X1 U23978 ( .A1(n21031), .A2(n21030), .A3(n21029), .A4(n21028), .ZN(
        n21045) );
  INV_X1 U23979 ( .A(DATAI_13_), .ZN(n21263) );
  AOI22_X1 U23980 ( .A1(n21241), .A2(keyinput_g41), .B1(n21263), .B2(
        keyinput_g19), .ZN(n21032) );
  OAI221_X1 U23981 ( .B1(n21241), .B2(keyinput_g41), .C1(n21263), .C2(
        keyinput_g19), .A(n21032), .ZN(n21043) );
  INV_X1 U23982 ( .A(READY1), .ZN(n21035) );
  AOI22_X1 U23983 ( .A1(n21035), .A2(keyinput_g36), .B1(keyinput_g96), .B2(
        n21034), .ZN(n21033) );
  OAI221_X1 U23984 ( .B1(n21035), .B2(keyinput_g36), .C1(n21034), .C2(
        keyinput_g96), .A(n21033), .ZN(n21042) );
  INV_X1 U23985 ( .A(DATAI_5_), .ZN(n21177) );
  AOI22_X1 U23986 ( .A1(n21168), .A2(keyinput_g92), .B1(keyinput_g27), .B2(
        n21177), .ZN(n21036) );
  OAI221_X1 U23987 ( .B1(n21168), .B2(keyinput_g92), .C1(n21177), .C2(
        keyinput_g27), .A(n21036), .ZN(n21041) );
  INV_X1 U23988 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n21039) );
  INV_X1 U23989 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n21038) );
  AOI22_X1 U23990 ( .A1(n21039), .A2(keyinput_g98), .B1(keyinput_g60), .B2(
        n21038), .ZN(n21037) );
  OAI221_X1 U23991 ( .B1(n21039), .B2(keyinput_g98), .C1(n21038), .C2(
        keyinput_g60), .A(n21037), .ZN(n21040) );
  NOR4_X1 U23992 ( .A1(n21043), .A2(n21042), .A3(n21041), .A4(n21040), .ZN(
        n21044) );
  NAND4_X1 U23993 ( .A1(n21047), .A2(n21046), .A3(n21045), .A4(n21044), .ZN(
        n21048) );
  NOR4_X1 U23994 ( .A1(n21051), .A2(n21050), .A3(n21049), .A4(n21048), .ZN(
        n21089) );
  OAI22_X1 U23995 ( .A1(P1_EBX_REG_22__SCAN_IN), .A2(keyinput_g93), .B1(
        P1_BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_g51), .ZN(n21052) );
  AOI221_X1 U23996 ( .B1(P1_EBX_REG_22__SCAN_IN), .B2(keyinput_g93), .C1(
        keyinput_g51), .C2(P1_BYTEENABLE_REG_3__SCAN_IN), .A(n21052), .ZN(
        n21059) );
  OAI22_X1 U23997 ( .A1(P1_EBX_REG_25__SCAN_IN), .A2(keyinput_g90), .B1(
        DATAI_31_), .B2(keyinput_g1), .ZN(n21053) );
  AOI221_X1 U23998 ( .B1(P1_EBX_REG_25__SCAN_IN), .B2(keyinput_g90), .C1(
        keyinput_g1), .C2(DATAI_31_), .A(n21053), .ZN(n21058) );
  OAI22_X1 U23999 ( .A1(DATAI_8_), .A2(keyinput_g24), .B1(DATAI_6_), .B2(
        keyinput_g26), .ZN(n21054) );
  AOI221_X1 U24000 ( .B1(DATAI_8_), .B2(keyinput_g24), .C1(keyinput_g26), .C2(
        DATAI_6_), .A(n21054), .ZN(n21057) );
  OAI22_X1 U24001 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(keyinput_g79), .B1(
        keyinput_g12), .B2(DATAI_20_), .ZN(n21055) );
  AOI221_X1 U24002 ( .B1(P1_REIP_REG_4__SCAN_IN), .B2(keyinput_g79), .C1(
        DATAI_20_), .C2(keyinput_g12), .A(n21055), .ZN(n21056) );
  NAND4_X1 U24003 ( .A1(n21059), .A2(n21058), .A3(n21057), .A4(n21056), .ZN(
        n21087) );
  OAI22_X1 U24004 ( .A1(DATAI_11_), .A2(keyinput_g21), .B1(keyinput_g33), .B2(
        HOLD), .ZN(n21060) );
  AOI221_X1 U24005 ( .B1(DATAI_11_), .B2(keyinput_g21), .C1(HOLD), .C2(
        keyinput_g33), .A(n21060), .ZN(n21067) );
  OAI22_X1 U24006 ( .A1(P1_EBX_REG_2__SCAN_IN), .A2(keyinput_g113), .B1(
        P1_REIP_REG_26__SCAN_IN), .B2(keyinput_g57), .ZN(n21061) );
  AOI221_X1 U24007 ( .B1(P1_EBX_REG_2__SCAN_IN), .B2(keyinput_g113), .C1(
        keyinput_g57), .C2(P1_REIP_REG_26__SCAN_IN), .A(n21061), .ZN(n21066)
         );
  OAI22_X1 U24008 ( .A1(P1_EAX_REG_28__SCAN_IN), .A2(keyinput_g119), .B1(
        DATAI_7_), .B2(keyinput_g25), .ZN(n21062) );
  AOI221_X1 U24009 ( .B1(P1_EAX_REG_28__SCAN_IN), .B2(keyinput_g119), .C1(
        keyinput_g25), .C2(DATAI_7_), .A(n21062), .ZN(n21065) );
  OAI22_X1 U24010 ( .A1(P1_EAX_REG_23__SCAN_IN), .A2(keyinput_g124), .B1(
        keyinput_g94), .B2(P1_EBX_REG_21__SCAN_IN), .ZN(n21063) );
  AOI221_X1 U24011 ( .B1(P1_EAX_REG_23__SCAN_IN), .B2(keyinput_g124), .C1(
        P1_EBX_REG_21__SCAN_IN), .C2(keyinput_g94), .A(n21063), .ZN(n21064) );
  NAND4_X1 U24012 ( .A1(n21067), .A2(n21066), .A3(n21065), .A4(n21064), .ZN(
        n21086) );
  OAI22_X1 U24013 ( .A1(P1_REIP_REG_31__SCAN_IN), .A2(keyinput_g52), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(keyinput_g61), .ZN(n21068) );
  AOI221_X1 U24014 ( .B1(P1_REIP_REG_31__SCAN_IN), .B2(keyinput_g52), .C1(
        keyinput_g61), .C2(P1_REIP_REG_22__SCAN_IN), .A(n21068), .ZN(n21075)
         );
  OAI22_X1 U24015 ( .A1(P1_EBX_REG_28__SCAN_IN), .A2(keyinput_g87), .B1(
        keyinput_g54), .B2(P1_REIP_REG_29__SCAN_IN), .ZN(n21069) );
  AOI221_X1 U24016 ( .B1(P1_EBX_REG_28__SCAN_IN), .B2(keyinput_g87), .C1(
        P1_REIP_REG_29__SCAN_IN), .C2(keyinput_g54), .A(n21069), .ZN(n21074)
         );
  OAI22_X1 U24017 ( .A1(P1_EBX_REG_20__SCAN_IN), .A2(keyinput_g95), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(keyinput_g78), .ZN(n21070) );
  AOI221_X1 U24018 ( .B1(P1_EBX_REG_20__SCAN_IN), .B2(keyinput_g95), .C1(
        keyinput_g78), .C2(P1_REIP_REG_5__SCAN_IN), .A(n21070), .ZN(n21073) );
  OAI22_X1 U24019 ( .A1(P1_EBX_REG_3__SCAN_IN), .A2(keyinput_g112), .B1(
        keyinput_g82), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n21071) );
  AOI221_X1 U24020 ( .B1(P1_EBX_REG_3__SCAN_IN), .B2(keyinput_g112), .C1(
        P1_REIP_REG_1__SCAN_IN), .C2(keyinput_g82), .A(n21071), .ZN(n21072) );
  NAND4_X1 U24021 ( .A1(n21075), .A2(n21074), .A3(n21073), .A4(n21072), .ZN(
        n21085) );
  OAI22_X1 U24022 ( .A1(P1_EBX_REG_16__SCAN_IN), .A2(keyinput_g99), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(keyinput_g66), .ZN(n21076) );
  AOI221_X1 U24023 ( .B1(P1_EBX_REG_16__SCAN_IN), .B2(keyinput_g99), .C1(
        keyinput_g66), .C2(P1_REIP_REG_17__SCAN_IN), .A(n21076), .ZN(n21083)
         );
  OAI22_X1 U24024 ( .A1(P1_EBX_REG_8__SCAN_IN), .A2(keyinput_g107), .B1(
        keyinput_g50), .B2(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21077) );
  AOI221_X1 U24025 ( .B1(P1_EBX_REG_8__SCAN_IN), .B2(keyinput_g107), .C1(
        P1_BYTEENABLE_REG_2__SCAN_IN), .C2(keyinput_g50), .A(n21077), .ZN(
        n21082) );
  OAI22_X1 U24026 ( .A1(P1_EBX_REG_4__SCAN_IN), .A2(keyinput_g111), .B1(
        P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_g40), .ZN(n21078) );
  AOI221_X1 U24027 ( .B1(P1_EBX_REG_4__SCAN_IN), .B2(keyinput_g111), .C1(
        keyinput_g40), .C2(P1_CODEFETCH_REG_SCAN_IN), .A(n21078), .ZN(n21081)
         );
  OAI22_X1 U24028 ( .A1(n21104), .A2(keyinput_g5), .B1(keyinput_g14), .B2(
        DATAI_18_), .ZN(n21079) );
  AOI221_X1 U24029 ( .B1(n21104), .B2(keyinput_g5), .C1(DATAI_18_), .C2(
        keyinput_g14), .A(n21079), .ZN(n21080) );
  NAND4_X1 U24030 ( .A1(n21083), .A2(n21082), .A3(n21081), .A4(n21080), .ZN(
        n21084) );
  NOR4_X1 U24031 ( .A1(n21087), .A2(n21086), .A3(n21085), .A4(n21084), .ZN(
        n21088) );
  AOI22_X1 U24032 ( .A1(n21089), .A2(n21088), .B1(keyinput_g45), .B2(n21301), 
        .ZN(n21300) );
  INV_X1 U24033 ( .A(keyinput_f45), .ZN(n21298) );
  AOI22_X1 U24034 ( .A1(READY2), .A2(keyinput_f37), .B1(DATAI_12_), .B2(
        keyinput_f20), .ZN(n21090) );
  OAI221_X1 U24035 ( .B1(READY2), .B2(keyinput_f37), .C1(DATAI_12_), .C2(
        keyinput_f20), .A(n21090), .ZN(n21097) );
  AOI22_X1 U24036 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(keyinput_f82), .B1(
        P1_EBX_REG_6__SCAN_IN), .B2(keyinput_f109), .ZN(n21091) );
  OAI221_X1 U24037 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(keyinput_f82), .C1(
        P1_EBX_REG_6__SCAN_IN), .C2(keyinput_f109), .A(n21091), .ZN(n21096) );
  AOI22_X1 U24038 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(keyinput_f62), .B1(
        P1_EBX_REG_18__SCAN_IN), .B2(keyinput_f97), .ZN(n21092) );
  OAI221_X1 U24039 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(keyinput_f62), .C1(
        P1_EBX_REG_18__SCAN_IN), .C2(keyinput_f97), .A(n21092), .ZN(n21095) );
  AOI22_X1 U24040 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(keyinput_f69), .B1(
        P1_EBX_REG_17__SCAN_IN), .B2(keyinput_f98), .ZN(n21093) );
  OAI221_X1 U24041 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(keyinput_f69), .C1(
        P1_EBX_REG_17__SCAN_IN), .C2(keyinput_f98), .A(n21093), .ZN(n21094) );
  NOR4_X1 U24042 ( .A1(n21097), .A2(n21096), .A3(n21095), .A4(n21094), .ZN(
        n21296) );
  AOI22_X1 U24043 ( .A1(P1_EBX_REG_1__SCAN_IN), .A2(keyinput_f114), .B1(
        P1_EBX_REG_21__SCAN_IN), .B2(keyinput_f94), .ZN(n21098) );
  OAI221_X1 U24044 ( .B1(P1_EBX_REG_1__SCAN_IN), .B2(keyinput_f114), .C1(
        P1_EBX_REG_21__SCAN_IN), .C2(keyinput_f94), .A(n21098), .ZN(n21124) );
  OAI22_X1 U24045 ( .A1(DATAI_21_), .A2(keyinput_f11), .B1(DATAI_19_), .B2(
        keyinput_f13), .ZN(n21099) );
  AOI221_X1 U24046 ( .B1(DATAI_21_), .B2(keyinput_f11), .C1(keyinput_f13), 
        .C2(DATAI_19_), .A(n21099), .ZN(n21103) );
  AOI22_X1 U24047 ( .A1(keyinput_f47), .A2(P1_W_R_N_REG_SCAN_IN), .B1(
        P1_EBX_REG_2__SCAN_IN), .B2(keyinput_f113), .ZN(n21100) );
  OAI221_X1 U24048 ( .B1(keyinput_f47), .B2(P1_W_R_N_REG_SCAN_IN), .C1(
        P1_EBX_REG_2__SCAN_IN), .C2(keyinput_f113), .A(n21100), .ZN(n21101) );
  AOI21_X1 U24049 ( .B1(keyinput_f5), .B2(n21104), .A(n21101), .ZN(n21102) );
  OAI211_X1 U24050 ( .C1(keyinput_f5), .C2(n21104), .A(n21103), .B(n21102), 
        .ZN(n21123) );
  OAI22_X1 U24051 ( .A1(P1_EAX_REG_21__SCAN_IN), .A2(keyinput_f126), .B1(
        P1_REIP_REG_4__SCAN_IN), .B2(keyinput_f79), .ZN(n21105) );
  AOI221_X1 U24052 ( .B1(P1_EAX_REG_21__SCAN_IN), .B2(keyinput_f126), .C1(
        keyinput_f79), .C2(P1_REIP_REG_4__SCAN_IN), .A(n21105), .ZN(n21112) );
  OAI22_X1 U24053 ( .A1(P1_EBX_REG_8__SCAN_IN), .A2(keyinput_f107), .B1(
        DATAI_10_), .B2(keyinput_f22), .ZN(n21106) );
  AOI221_X1 U24054 ( .B1(P1_EBX_REG_8__SCAN_IN), .B2(keyinput_f107), .C1(
        keyinput_f22), .C2(DATAI_10_), .A(n21106), .ZN(n21111) );
  OAI22_X1 U24055 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(keyinput_f65), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(keyinput_f67), .ZN(n21107) );
  AOI221_X1 U24056 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(keyinput_f65), .C1(
        keyinput_f67), .C2(P1_REIP_REG_16__SCAN_IN), .A(n21107), .ZN(n21110)
         );
  OAI22_X1 U24057 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(keyinput_f68), .B1(
        P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_f40), .ZN(n21108) );
  AOI221_X1 U24058 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(keyinput_f68), .C1(
        keyinput_f40), .C2(P1_CODEFETCH_REG_SCAN_IN), .A(n21108), .ZN(n21109)
         );
  NAND4_X1 U24059 ( .A1(n21112), .A2(n21111), .A3(n21110), .A4(n21109), .ZN(
        n21122) );
  OAI22_X1 U24060 ( .A1(P1_EBX_REG_20__SCAN_IN), .A2(keyinput_f95), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(keyinput_f76), .ZN(n21113) );
  AOI221_X1 U24061 ( .B1(P1_EBX_REG_20__SCAN_IN), .B2(keyinput_f95), .C1(
        keyinput_f76), .C2(P1_REIP_REG_7__SCAN_IN), .A(n21113), .ZN(n21120) );
  OAI22_X1 U24062 ( .A1(READY1), .A2(keyinput_f36), .B1(DATAI_11_), .B2(
        keyinput_f21), .ZN(n21114) );
  AOI221_X1 U24063 ( .B1(READY1), .B2(keyinput_f36), .C1(keyinput_f21), .C2(
        DATAI_11_), .A(n21114), .ZN(n21119) );
  OAI22_X1 U24064 ( .A1(DATAI_8_), .A2(keyinput_f24), .B1(DATAI_20_), .B2(
        keyinput_f12), .ZN(n21115) );
  AOI221_X1 U24065 ( .B1(DATAI_8_), .B2(keyinput_f24), .C1(keyinput_f12), .C2(
        DATAI_20_), .A(n21115), .ZN(n21118) );
  OAI22_X1 U24066 ( .A1(P1_EBX_REG_19__SCAN_IN), .A2(keyinput_f96), .B1(
        keyinput_f60), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n21116) );
  AOI221_X1 U24067 ( .B1(P1_EBX_REG_19__SCAN_IN), .B2(keyinput_f96), .C1(
        P1_REIP_REG_23__SCAN_IN), .C2(keyinput_f60), .A(n21116), .ZN(n21117)
         );
  NAND4_X1 U24068 ( .A1(n21120), .A2(n21119), .A3(n21118), .A4(n21117), .ZN(
        n21121) );
  NOR4_X1 U24069 ( .A1(n21124), .A2(n21123), .A3(n21122), .A4(n21121), .ZN(
        n21295) );
  OAI22_X1 U24070 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(keyinput_f57), .B1(
        keyinput_f71), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n21125) );
  AOI221_X1 U24071 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(keyinput_f57), .C1(
        P1_REIP_REG_12__SCAN_IN), .C2(keyinput_f71), .A(n21125), .ZN(n21132)
         );
  OAI22_X1 U24072 ( .A1(P1_EBX_REG_28__SCAN_IN), .A2(keyinput_f87), .B1(
        keyinput_f48), .B2(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21126) );
  AOI221_X1 U24073 ( .B1(P1_EBX_REG_28__SCAN_IN), .B2(keyinput_f87), .C1(
        P1_BYTEENABLE_REG_0__SCAN_IN), .C2(keyinput_f48), .A(n21126), .ZN(
        n21131) );
  OAI22_X1 U24074 ( .A1(P1_EBX_REG_9__SCAN_IN), .A2(keyinput_f106), .B1(
        DATAI_23_), .B2(keyinput_f9), .ZN(n21127) );
  AOI221_X1 U24075 ( .B1(P1_EBX_REG_9__SCAN_IN), .B2(keyinput_f106), .C1(
        keyinput_f9), .C2(DATAI_23_), .A(n21127), .ZN(n21130) );
  OAI22_X1 U24076 ( .A1(P1_EBX_REG_16__SCAN_IN), .A2(keyinput_f99), .B1(
        DATAI_16_), .B2(keyinput_f16), .ZN(n21128) );
  AOI221_X1 U24077 ( .B1(P1_EBX_REG_16__SCAN_IN), .B2(keyinput_f99), .C1(
        keyinput_f16), .C2(DATAI_16_), .A(n21128), .ZN(n21129) );
  NAND4_X1 U24078 ( .A1(n21132), .A2(n21131), .A3(n21130), .A4(n21129), .ZN(
        n21160) );
  OAI22_X1 U24079 ( .A1(DATAI_31_), .A2(keyinput_f1), .B1(keyinput_f64), .B2(
        P1_REIP_REG_19__SCAN_IN), .ZN(n21133) );
  AOI221_X1 U24080 ( .B1(DATAI_31_), .B2(keyinput_f1), .C1(
        P1_REIP_REG_19__SCAN_IN), .C2(keyinput_f64), .A(n21133), .ZN(n21140)
         );
  OAI22_X1 U24081 ( .A1(DATAI_7_), .A2(keyinput_f25), .B1(keyinput_f49), .B2(
        P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21134) );
  AOI221_X1 U24082 ( .B1(DATAI_7_), .B2(keyinput_f25), .C1(
        P1_BYTEENABLE_REG_1__SCAN_IN), .C2(keyinput_f49), .A(n21134), .ZN(
        n21139) );
  OAI22_X1 U24083 ( .A1(P1_EBX_REG_4__SCAN_IN), .A2(keyinput_f111), .B1(
        keyinput_f15), .B2(DATAI_17_), .ZN(n21135) );
  AOI221_X1 U24084 ( .B1(P1_EBX_REG_4__SCAN_IN), .B2(keyinput_f111), .C1(
        DATAI_17_), .C2(keyinput_f15), .A(n21135), .ZN(n21138) );
  OAI22_X1 U24085 ( .A1(P1_EBX_REG_29__SCAN_IN), .A2(keyinput_f86), .B1(
        keyinput_f88), .B2(P1_EBX_REG_27__SCAN_IN), .ZN(n21136) );
  AOI221_X1 U24086 ( .B1(P1_EBX_REG_29__SCAN_IN), .B2(keyinput_f86), .C1(
        P1_EBX_REG_27__SCAN_IN), .C2(keyinput_f88), .A(n21136), .ZN(n21137) );
  NAND4_X1 U24087 ( .A1(n21140), .A2(n21139), .A3(n21138), .A4(n21137), .ZN(
        n21159) );
  OAI22_X1 U24088 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(keyinput_f73), .B1(
        keyinput_f23), .B2(DATAI_9_), .ZN(n21141) );
  AOI221_X1 U24089 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(keyinput_f73), .C1(
        DATAI_9_), .C2(keyinput_f23), .A(n21141), .ZN(n21148) );
  OAI22_X1 U24090 ( .A1(P1_EBX_REG_13__SCAN_IN), .A2(keyinput_f102), .B1(
        keyinput_f42), .B2(P1_D_C_N_REG_SCAN_IN), .ZN(n21142) );
  AOI221_X1 U24091 ( .B1(P1_EBX_REG_13__SCAN_IN), .B2(keyinput_f102), .C1(
        P1_D_C_N_REG_SCAN_IN), .C2(keyinput_f42), .A(n21142), .ZN(n21147) );
  OAI22_X1 U24092 ( .A1(P1_EBX_REG_24__SCAN_IN), .A2(keyinput_f91), .B1(
        keyinput_f70), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n21143) );
  AOI221_X1 U24093 ( .B1(P1_EBX_REG_24__SCAN_IN), .B2(keyinput_f91), .C1(
        P1_REIP_REG_13__SCAN_IN), .C2(keyinput_f70), .A(n21143), .ZN(n21146)
         );
  OAI22_X1 U24094 ( .A1(P1_EAX_REG_30__SCAN_IN), .A2(keyinput_f117), .B1(
        keyinput_f32), .B2(DATAI_0_), .ZN(n21144) );
  AOI221_X1 U24095 ( .B1(P1_EAX_REG_30__SCAN_IN), .B2(keyinput_f117), .C1(
        DATAI_0_), .C2(keyinput_f32), .A(n21144), .ZN(n21145) );
  NAND4_X1 U24096 ( .A1(n21148), .A2(n21147), .A3(n21146), .A4(n21145), .ZN(
        n21158) );
  OAI22_X1 U24097 ( .A1(P1_EAX_REG_31__SCAN_IN), .A2(keyinput_f116), .B1(
        keyinput_f14), .B2(DATAI_18_), .ZN(n21149) );
  AOI221_X1 U24098 ( .B1(P1_EAX_REG_31__SCAN_IN), .B2(keyinput_f116), .C1(
        DATAI_18_), .C2(keyinput_f14), .A(n21149), .ZN(n21156) );
  OAI22_X1 U24099 ( .A1(P1_EBX_REG_12__SCAN_IN), .A2(keyinput_f103), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(keyinput_f61), .ZN(n21150) );
  AOI221_X1 U24100 ( .B1(P1_EBX_REG_12__SCAN_IN), .B2(keyinput_f103), .C1(
        keyinput_f61), .C2(P1_REIP_REG_22__SCAN_IN), .A(n21150), .ZN(n21155)
         );
  OAI22_X1 U24101 ( .A1(DATAI_14_), .A2(keyinput_f18), .B1(
        P1_FLUSH_REG_SCAN_IN), .B2(keyinput_f46), .ZN(n21151) );
  AOI221_X1 U24102 ( .B1(DATAI_14_), .B2(keyinput_f18), .C1(keyinput_f46), 
        .C2(P1_FLUSH_REG_SCAN_IN), .A(n21151), .ZN(n21154) );
  OAI22_X1 U24103 ( .A1(P1_EAX_REG_27__SCAN_IN), .A2(keyinput_f120), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(keyinput_f118), .ZN(n21152) );
  AOI221_X1 U24104 ( .B1(P1_EAX_REG_27__SCAN_IN), .B2(keyinput_f120), .C1(
        keyinput_f118), .C2(P1_EAX_REG_29__SCAN_IN), .A(n21152), .ZN(n21153)
         );
  NAND4_X1 U24105 ( .A1(n21156), .A2(n21155), .A3(n21154), .A4(n21153), .ZN(
        n21157) );
  NOR4_X1 U24106 ( .A1(n21160), .A2(n21159), .A3(n21158), .A4(n21157), .ZN(
        n21294) );
  AOI22_X1 U24107 ( .A1(DATAI_15_), .A2(keyinput_f17), .B1(n21162), .B2(
        keyinput_f83), .ZN(n21161) );
  OAI221_X1 U24108 ( .B1(DATAI_15_), .B2(keyinput_f17), .C1(n21162), .C2(
        keyinput_f83), .A(n21161), .ZN(n21175) );
  INV_X1 U24109 ( .A(keyinput_f50), .ZN(n21164) );
  AOI22_X1 U24110 ( .A1(n21165), .A2(keyinput_f81), .B1(
        P1_BYTEENABLE_REG_2__SCAN_IN), .B2(n21164), .ZN(n21163) );
  OAI221_X1 U24111 ( .B1(n21165), .B2(keyinput_f81), .C1(n21164), .C2(
        P1_BYTEENABLE_REG_2__SCAN_IN), .A(n21163), .ZN(n21174) );
  AOI22_X1 U24112 ( .A1(n21168), .A2(keyinput_f92), .B1(keyinput_f6), .B2(
        n21167), .ZN(n21166) );
  OAI221_X1 U24113 ( .B1(n21168), .B2(keyinput_f92), .C1(n21167), .C2(
        keyinput_f6), .A(n21166), .ZN(n21173) );
  AOI22_X1 U24114 ( .A1(n21171), .A2(keyinput_f63), .B1(keyinput_f38), .B2(
        n21170), .ZN(n21169) );
  OAI221_X1 U24115 ( .B1(n21171), .B2(keyinput_f63), .C1(n21170), .C2(
        keyinput_f38), .A(n21169), .ZN(n21172) );
  NOR4_X1 U24116 ( .A1(n21175), .A2(n21174), .A3(n21173), .A4(n21172), .ZN(
        n21224) );
  INV_X1 U24117 ( .A(DATAI_2_), .ZN(n21178) );
  AOI22_X1 U24118 ( .A1(n21178), .A2(keyinput_f30), .B1(n21177), .B2(
        keyinput_f27), .ZN(n21176) );
  OAI221_X1 U24119 ( .B1(n21178), .B2(keyinput_f30), .C1(n21177), .C2(
        keyinput_f27), .A(n21176), .ZN(n21191) );
  AOI22_X1 U24120 ( .A1(n21181), .A2(keyinput_f0), .B1(keyinput_f34), .B2(
        n21180), .ZN(n21179) );
  OAI221_X1 U24121 ( .B1(n21181), .B2(keyinput_f0), .C1(n21180), .C2(
        keyinput_f34), .A(n21179), .ZN(n21190) );
  AOI22_X1 U24122 ( .A1(n21184), .A2(keyinput_f104), .B1(keyinput_f53), .B2(
        n21183), .ZN(n21182) );
  OAI221_X1 U24123 ( .B1(n21184), .B2(keyinput_f104), .C1(n21183), .C2(
        keyinput_f53), .A(n21182), .ZN(n21189) );
  AOI22_X1 U24124 ( .A1(n21187), .A2(keyinput_f123), .B1(keyinput_f7), .B2(
        n21186), .ZN(n21185) );
  OAI221_X1 U24125 ( .B1(n21187), .B2(keyinput_f123), .C1(n21186), .C2(
        keyinput_f7), .A(n21185), .ZN(n21188) );
  NOR4_X1 U24126 ( .A1(n21191), .A2(n21190), .A3(n21189), .A4(n21188), .ZN(
        n21223) );
  AOI22_X1 U24127 ( .A1(n14532), .A2(keyinput_f66), .B1(n21193), .B2(
        keyinput_f90), .ZN(n21192) );
  OAI221_X1 U24128 ( .B1(n14532), .B2(keyinput_f66), .C1(n21193), .C2(
        keyinput_f90), .A(n21192), .ZN(n21205) );
  AOI22_X1 U24129 ( .A1(n21196), .A2(keyinput_f3), .B1(n21195), .B2(
        keyinput_f72), .ZN(n21194) );
  OAI221_X1 U24130 ( .B1(n21196), .B2(keyinput_f3), .C1(n21195), .C2(
        keyinput_f72), .A(n21194), .ZN(n21204) );
  AOI22_X1 U24131 ( .A1(n21199), .A2(keyinput_f39), .B1(n21198), .B2(
        keyinput_f59), .ZN(n21197) );
  OAI221_X1 U24132 ( .B1(n21199), .B2(keyinput_f39), .C1(n21198), .C2(
        keyinput_f59), .A(n21197), .ZN(n21203) );
  AOI22_X1 U24133 ( .A1(n13564), .A2(keyinput_f105), .B1(n21201), .B2(
        keyinput_f108), .ZN(n21200) );
  OAI221_X1 U24134 ( .B1(n13564), .B2(keyinput_f105), .C1(n21201), .C2(
        keyinput_f108), .A(n21200), .ZN(n21202) );
  NOR4_X1 U24135 ( .A1(n21205), .A2(n21204), .A3(n21203), .A4(n21202), .ZN(
        n21222) );
  AOI22_X1 U24136 ( .A1(n21208), .A2(keyinput_f75), .B1(keyinput_f10), .B2(
        n21207), .ZN(n21206) );
  OAI221_X1 U24137 ( .B1(n21208), .B2(keyinput_f75), .C1(n21207), .C2(
        keyinput_f10), .A(n21206), .ZN(n21220) );
  AOI22_X1 U24138 ( .A1(n21210), .A2(keyinput_f8), .B1(n13635), .B2(
        keyinput_f74), .ZN(n21209) );
  OAI221_X1 U24139 ( .B1(n21210), .B2(keyinput_f8), .C1(n13635), .C2(
        keyinput_f74), .A(n21209), .ZN(n21219) );
  INV_X1 U24140 ( .A(DATAI_4_), .ZN(n21213) );
  AOI22_X1 U24141 ( .A1(n21213), .A2(keyinput_f28), .B1(n21212), .B2(
        keyinput_f58), .ZN(n21211) );
  OAI221_X1 U24142 ( .B1(n21213), .B2(keyinput_f28), .C1(n21212), .C2(
        keyinput_f58), .A(n21211), .ZN(n21218) );
  AOI22_X1 U24143 ( .A1(n21216), .A2(keyinput_f43), .B1(n21215), .B2(
        keyinput_f121), .ZN(n21214) );
  OAI221_X1 U24144 ( .B1(n21216), .B2(keyinput_f43), .C1(n21215), .C2(
        keyinput_f121), .A(n21214), .ZN(n21217) );
  NOR4_X1 U24145 ( .A1(n21220), .A2(n21219), .A3(n21218), .A4(n21217), .ZN(
        n21221) );
  NAND4_X1 U24146 ( .A1(n21224), .A2(n21223), .A3(n21222), .A4(n21221), .ZN(
        n21292) );
  AOI22_X1 U24147 ( .A1(n21227), .A2(keyinput_f55), .B1(n21226), .B2(
        keyinput_f85), .ZN(n21225) );
  OAI221_X1 U24148 ( .B1(n21227), .B2(keyinput_f55), .C1(n21226), .C2(
        keyinput_f85), .A(n21225), .ZN(n21291) );
  OAI22_X1 U24149 ( .A1(n21230), .A2(keyinput_f80), .B1(n21229), .B2(
        keyinput_f31), .ZN(n21228) );
  AOI221_X1 U24150 ( .B1(n21230), .B2(keyinput_f80), .C1(keyinput_f31), .C2(
        n21229), .A(n21228), .ZN(n21239) );
  OAI22_X1 U24151 ( .A1(n21233), .A2(keyinput_f84), .B1(n21232), .B2(
        keyinput_f33), .ZN(n21231) );
  AOI221_X1 U24152 ( .B1(n21233), .B2(keyinput_f84), .C1(keyinput_f33), .C2(
        n21232), .A(n21231), .ZN(n21238) );
  OAI22_X1 U24153 ( .A1(n21236), .A2(keyinput_f101), .B1(n21235), .B2(
        keyinput_f77), .ZN(n21234) );
  AOI221_X1 U24154 ( .B1(n21236), .B2(keyinput_f101), .C1(keyinput_f77), .C2(
        n21235), .A(n21234), .ZN(n21237) );
  NAND3_X1 U24155 ( .A1(n21239), .A2(n21238), .A3(n21237), .ZN(n21290) );
  OAI22_X1 U24156 ( .A1(keyinput_f51), .A2(n21242), .B1(n21241), .B2(
        keyinput_f41), .ZN(n21240) );
  AOI221_X1 U24157 ( .B1(n21242), .B2(keyinput_f51), .C1(n21241), .C2(
        keyinput_f41), .A(n21240), .ZN(n21288) );
  AOI22_X1 U24158 ( .A1(n21245), .A2(keyinput_f29), .B1(n21244), .B2(
        keyinput_f125), .ZN(n21243) );
  OAI221_X1 U24159 ( .B1(n21245), .B2(keyinput_f29), .C1(n21244), .C2(
        keyinput_f125), .A(n21243), .ZN(n21254) );
  AOI22_X1 U24160 ( .A1(n21248), .A2(keyinput_f112), .B1(n21247), .B2(
        keyinput_f124), .ZN(n21246) );
  OAI221_X1 U24161 ( .B1(n21248), .B2(keyinput_f112), .C1(n21247), .C2(
        keyinput_f124), .A(n21246), .ZN(n21253) );
  INV_X1 U24162 ( .A(BS16), .ZN(n21250) );
  AOI22_X1 U24163 ( .A1(n21251), .A2(keyinput_f2), .B1(keyinput_f35), .B2(
        n21250), .ZN(n21249) );
  OAI221_X1 U24164 ( .B1(n21251), .B2(keyinput_f2), .C1(n21250), .C2(
        keyinput_f35), .A(n21249), .ZN(n21252) );
  NOR3_X1 U24165 ( .A1(n21254), .A2(n21253), .A3(n21252), .ZN(n21287) );
  AOI22_X1 U24166 ( .A1(n21257), .A2(keyinput_f52), .B1(n21256), .B2(
        keyinput_f127), .ZN(n21255) );
  OAI221_X1 U24167 ( .B1(n21257), .B2(keyinput_f52), .C1(n21256), .C2(
        keyinput_f127), .A(n21255), .ZN(n21270) );
  AOI22_X1 U24168 ( .A1(n21260), .A2(keyinput_f93), .B1(n21259), .B2(
        keyinput_f89), .ZN(n21258) );
  OAI221_X1 U24169 ( .B1(n21260), .B2(keyinput_f93), .C1(n21259), .C2(
        keyinput_f89), .A(n21258), .ZN(n21269) );
  AOI22_X1 U24170 ( .A1(n21263), .A2(keyinput_f19), .B1(n21262), .B2(
        keyinput_f54), .ZN(n21261) );
  OAI221_X1 U24171 ( .B1(n21263), .B2(keyinput_f19), .C1(n21262), .C2(
        keyinput_f54), .A(n21261), .ZN(n21268) );
  AOI22_X1 U24172 ( .A1(n21266), .A2(keyinput_f56), .B1(n21265), .B2(
        keyinput_f110), .ZN(n21264) );
  OAI221_X1 U24173 ( .B1(n21266), .B2(keyinput_f56), .C1(n21265), .C2(
        keyinput_f110), .A(n21264), .ZN(n21267) );
  NOR4_X1 U24174 ( .A1(n21270), .A2(n21269), .A3(n21268), .A4(n21267), .ZN(
        n21286) );
  AOI22_X1 U24175 ( .A1(n21272), .A2(keyinput_f78), .B1(n12796), .B2(
        keyinput_f115), .ZN(n21271) );
  OAI221_X1 U24176 ( .B1(n21272), .B2(keyinput_f78), .C1(n12796), .C2(
        keyinput_f115), .A(n21271), .ZN(n21284) );
  AOI22_X1 U24177 ( .A1(n21275), .A2(keyinput_f119), .B1(keyinput_f4), .B2(
        n21274), .ZN(n21273) );
  OAI221_X1 U24178 ( .B1(n21275), .B2(keyinput_f119), .C1(n21274), .C2(
        keyinput_f4), .A(n21273), .ZN(n21283) );
  INV_X1 U24179 ( .A(DATAI_6_), .ZN(n21277) );
  AOI22_X1 U24180 ( .A1(n14315), .A2(keyinput_f100), .B1(keyinput_f26), .B2(
        n21277), .ZN(n21276) );
  OAI221_X1 U24181 ( .B1(n14315), .B2(keyinput_f100), .C1(n21277), .C2(
        keyinput_f26), .A(n21276), .ZN(n21282) );
  AOI22_X1 U24182 ( .A1(n21280), .A2(keyinput_f44), .B1(keyinput_f122), .B2(
        n21279), .ZN(n21278) );
  OAI221_X1 U24183 ( .B1(n21280), .B2(keyinput_f44), .C1(n21279), .C2(
        keyinput_f122), .A(n21278), .ZN(n21281) );
  NOR4_X1 U24184 ( .A1(n21284), .A2(n21283), .A3(n21282), .A4(n21281), .ZN(
        n21285) );
  NAND4_X1 U24185 ( .A1(n21288), .A2(n21287), .A3(n21286), .A4(n21285), .ZN(
        n21289) );
  NOR4_X1 U24186 ( .A1(n21292), .A2(n21291), .A3(n21290), .A4(n21289), .ZN(
        n21293) );
  NAND4_X1 U24187 ( .A1(n21296), .A2(n21295), .A3(n21294), .A4(n21293), .ZN(
        n21297) );
  OAI221_X1 U24188 ( .B1(P1_MORE_REG_SCAN_IN), .B2(keyinput_f45), .C1(n21301), 
        .C2(n21298), .A(n21297), .ZN(n21299) );
  OAI211_X1 U24189 ( .C1(keyinput_g45), .C2(n21301), .A(n21300), .B(n21299), 
        .ZN(n21302) );
  XOR2_X1 U24190 ( .A(n21303), .B(n21302), .Z(U355) );
  AND2_X1 U11596 ( .A1(n10320), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10478) );
  AND2_X1 U16366 ( .A1(n21304), .A2(n13198), .ZN(n19593) );
  INV_X1 U11262 ( .A(n14067), .ZN(n14070) );
  NAND3_X1 U11266 ( .A1(n10320), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10433) );
  CLKBUF_X1 U11316 ( .A(n11714), .Z(n11745) );
  AND2_X1 U11319 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n10472), .ZN(
        n10558) );
  CLKBUF_X1 U11336 ( .A(n10855), .Z(n9818) );
  INV_X1 U11348 ( .A(n10748), .ZN(n10768) );
  CLKBUF_X1 U11368 ( .A(n15175), .Z(n15477) );
  CLKBUF_X1 U11529 ( .A(n11121), .Z(n11122) );
  INV_X1 U11550 ( .A(n13366), .ZN(n19566) );
  CLKBUF_X1 U11573 ( .A(n15665), .Z(n17206) );
  CLKBUF_X1 U11590 ( .A(n19204), .Z(n19217) );
  CLKBUF_X2 U11672 ( .A(n15037), .Z(n9815) );
  CLKBUF_X1 U12439 ( .A(n15086), .Z(n15087) );
  CLKBUF_X1 U12584 ( .A(n17887), .Z(n9816) );
  AND2_X2 U12982 ( .A1(n13188), .A2(n13192), .ZN(n21304) );
endmodule

