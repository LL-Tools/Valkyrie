

module b22_C_gen_AntiSAT_k_128_3 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0,
         keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5,
         keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10,
         keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15,
         keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20,
         keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25,
         keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30,
         keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35,
         keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40,
         keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45,
         keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50,
         keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55,
         keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60,
         keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410;

  XNOR2_X1 U7218 ( .A(n8072), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14216) );
  CLKBUF_X2 U7219 ( .A(n8632), .Z(n6474) );
  NAND2_X1 U7220 ( .A1(n8908), .A2(n8912), .ZN(n8921) );
  NAND2_X1 U7221 ( .A1(n6830), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6829) );
  MUX2_X1 U7222 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8906), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8908) );
  INV_X1 U7223 ( .A(n8248), .ZN(n7693) );
  NAND4_X1 U7224 ( .A1(n6715), .A2(n7608), .A3(n7501), .A4(n7500), .ZN(n7503)
         );
  INV_X1 U7225 ( .A(n12773), .ZN(n12644) );
  INV_X2 U7226 ( .A(n12454), .ZN(n12441) );
  INV_X1 U7227 ( .A(n7552), .ZN(n7750) );
  NOR2_X2 U7228 ( .A1(n7503), .A2(n7588), .ZN(n7744) );
  OR2_X1 U7229 ( .A1(n12538), .A2(n8840), .ZN(n12201) );
  INV_X1 U7230 ( .A(n6725), .ZN(n13134) );
  AND2_X1 U7231 ( .A1(n10453), .A2(n10002), .ZN(n6519) );
  CLKBUF_X2 U7232 ( .A(n8632), .Z(n6475) );
  OAI21_X1 U7233 ( .B1(n8462), .B2(P3_IR_REG_18__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8453) );
  OR2_X1 U7234 ( .A1(n14439), .A2(n14438), .ZN(n14441) );
  NAND2_X1 U7235 ( .A1(n13638), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8973) );
  CLKBUF_X2 U7237 ( .A(n7644), .Z(n6492) );
  OAI21_X1 U7238 ( .B1(n9929), .B2(n7371), .A(n7370), .ZN(n13955) );
  INV_X1 U7239 ( .A(n14724), .ZN(n11494) );
  NAND2_X1 U7240 ( .A1(n7045), .A2(n7042), .ZN(n12121) );
  NAND2_X1 U7241 ( .A1(n9093), .A2(n9092), .ZN(n11216) );
  BUF_X1 U7242 ( .A(n9671), .Z(n6685) );
  INV_X1 U7243 ( .A(n9264), .ZN(n9357) );
  NAND2_X1 U7244 ( .A1(n14441), .A2(n9457), .ZN(n11701) );
  INV_X2 U7245 ( .A(n8181), .ZN(n7603) );
  OR3_X1 U7246 ( .A1(n10899), .A2(n15090), .A3(n15168), .ZN(n12933) );
  NAND4_X1 U7247 ( .A1(n9048), .A2(n9047), .A3(n9046), .A4(n9045), .ZN(n13267)
         );
  OR2_X1 U7248 ( .A1(n11106), .A2(n11107), .ZN(n6470) );
  AND2_X1 U7249 ( .A1(n9373), .A2(n9376), .ZN(n6471) );
  INV_X2 U7250 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n14274) );
  INV_X2 U7251 ( .A(n10641), .ZN(n13842) );
  AND4_X4 U7252 ( .A1(n7581), .A2(n7580), .A3(n7579), .A4(n7578), .ZN(n10641)
         );
  OAI21_X2 U7253 ( .B1(n8430), .B2(n8429), .A(n8410), .ZN(n8771) );
  OAI21_X2 U7254 ( .B1(n6691), .B2(n6690), .A(n9704), .ZN(n9712) );
  NAND2_X2 U7255 ( .A1(n9276), .A2(n9275), .ZN(n13575) );
  NOR2_X2 U7256 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8538) );
  OAI22_X2 U7257 ( .A1(n13465), .A2(n9461), .B1(n9431), .B2(n13219), .ZN(
        n13453) );
  NAND2_X2 U7258 ( .A1(n9373), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9372) );
  NAND4_X4 U7259 ( .A1(n7556), .A2(n7485), .A3(n7555), .A4(n7554), .ZN(n7573)
         );
  OAI21_X2 U7260 ( .B1(n11358), .B2(n7076), .A(n7073), .ZN(n11580) );
  NAND2_X2 U7261 ( .A1(n11281), .A2(n9785), .ZN(n11358) );
  XNOR2_X2 U7262 ( .A(n8237), .B(n8236), .ZN(n9665) );
  NAND2_X2 U7263 ( .A1(n8268), .A2(n8272), .ZN(n8237) );
  OR2_X1 U7264 ( .A1(n9018), .A2(n10590), .ZN(n9021) );
  NAND2_X2 U7265 ( .A1(n9017), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n9022) );
  INV_X2 U7266 ( .A(n8978), .ZN(n12008) );
  AND2_X4 U7267 ( .A1(n8482), .A2(n10022), .ZN(n12159) );
  XNOR2_X2 U7268 ( .A(n8295), .B(n13691), .ZN(n14006) );
  OAI21_X2 U7269 ( .B1(n13182), .B2(n7310), .A(n7316), .ZN(n7309) );
  NOR2_X2 U7270 ( .A1(n13184), .A2(n13183), .ZN(n13182) );
  INV_X1 U7271 ( .A(n6471), .ZN(n6472) );
  INV_X1 U7272 ( .A(n6471), .ZN(n6473) );
  INV_X2 U7273 ( .A(n10476), .ZN(n13489) );
  INV_X1 U7274 ( .A(n8482), .ZN(n8632) );
  XNOR2_X2 U7275 ( .A(n8388), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n8665) );
  NAND2_X2 U7276 ( .A1(n8387), .A2(n8386), .ZN(n8388) );
  AOI21_X2 U7277 ( .B1(n11491), .B2(n11489), .A(n11490), .ZN(n13759) );
  NAND2_X2 U7278 ( .A1(n10929), .A2(n10928), .ZN(n11491) );
  BUF_X8 U7279 ( .A(n10922), .Z(n12424) );
  NAND2_X2 U7280 ( .A1(n9658), .A2(n6687), .ZN(n9689) );
  OAI21_X2 U7281 ( .B1(n7684), .B2(n6785), .A(n6787), .ZN(n7718) );
  NAND2_X2 U7282 ( .A1(n7668), .A2(n7667), .ZN(n7684) );
  XNOR2_X2 U7283 ( .A(n6829), .B(n8352), .ZN(n8355) );
  XNOR2_X2 U7284 ( .A(n13082), .B(n13081), .ZN(n12519) );
  NAND2_X2 U7285 ( .A1(n9134), .A2(n9133), .ZN(n11052) );
  AOI21_X2 U7286 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(n14305), .A(n14545), .ZN(
        n14550) );
  NAND2_X1 U7287 ( .A1(n13962), .A2(n13961), .ZN(n13964) );
  CLKBUF_X2 U7288 ( .A(n9721), .Z(n13535) );
  NAND2_X1 U7289 ( .A1(n14161), .A2(n9993), .ZN(n14020) );
  AND2_X1 U7290 ( .A1(n7368), .A2(n13997), .ZN(n7367) );
  NAND2_X1 U7291 ( .A1(n14427), .A2(n11737), .ZN(n12499) );
  NAND2_X1 U7292 ( .A1(n11075), .A2(n11074), .ZN(n11343) );
  NAND2_X1 U7293 ( .A1(n10964), .A2(n12392), .ZN(n12400) );
  NOR2_X1 U7294 ( .A1(n9493), .A2(n7415), .ZN(n7413) );
  INV_X4 U7297 ( .A(n7750), .ZN(n8284) );
  INV_X1 U7298 ( .A(n9687), .ZN(n6476) );
  INV_X4 U7299 ( .A(n6519), .ZN(n12444) );
  CLKBUF_X1 U7300 ( .A(n9187), .Z(n9331) );
  NAND2_X4 U7301 ( .A1(n10453), .A2(n10469), .ZN(n12454) );
  BUF_X2 U7302 ( .A(n8509), .Z(n12145) );
  INV_X2 U7303 ( .A(n8333), .ZN(n7988) );
  NAND2_X4 U7304 ( .A1(n10107), .A2(n13650), .ZN(n10098) );
  INV_X2 U7305 ( .A(n7612), .ZN(n7530) );
  INV_X1 U7306 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7528) );
  AOI211_X1 U7307 ( .C1(n14111), .C2(n14683), .A(n13952), .B(n13951), .ZN(
        n13953) );
  NAND2_X1 U7308 ( .A1(n13947), .A2(n12021), .ZN(n12025) );
  NAND2_X1 U7309 ( .A1(n13700), .A2(n12431), .ZN(n13793) );
  NAND2_X1 U7310 ( .A1(n13982), .A2(n6574), .ZN(n14126) );
  AOI21_X1 U7311 ( .B1(n12015), .B2(n14618), .A(n12014), .ZN(n14110) );
  AOI21_X1 U7312 ( .B1(n7236), .B2(n7237), .A(n7234), .ZN(n7233) );
  AND2_X1 U7313 ( .A1(n6791), .A2(n6790), .ZN(n13405) );
  NAND2_X1 U7314 ( .A1(n8816), .A2(n8815), .ZN(n12949) );
  NAND2_X1 U7315 ( .A1(n8845), .A2(n8844), .ZN(n12137) );
  NAND2_X1 U7316 ( .A1(n6708), .A2(n13433), .ZN(n6791) );
  OR2_X1 U7317 ( .A1(n8842), .A2(n8841), .ZN(n8845) );
  NAND2_X1 U7318 ( .A1(n12827), .A2(n12826), .ZN(n12825) );
  OAI21_X1 U7319 ( .B1(n14021), .B2(n7369), .A(n7367), .ZN(n9927) );
  NAND2_X1 U7320 ( .A1(n7130), .A2(n6549), .ZN(n13424) );
  NAND2_X1 U7321 ( .A1(n8428), .A2(n8427), .ZN(n12578) );
  AOI21_X1 U7322 ( .B1(n8209), .B2(n8208), .A(n8207), .ZN(n8222) );
  NAND2_X1 U7323 ( .A1(n8785), .A2(n8784), .ZN(n12834) );
  NAND2_X1 U7324 ( .A1(n8798), .A2(n8797), .ZN(n8811) );
  OR2_X1 U7325 ( .A1(n14071), .A2(n7338), .ZN(n7339) );
  NAND2_X1 U7326 ( .A1(n9298), .A2(n9297), .ZN(n13401) );
  OAI21_X1 U7327 ( .B1(n11975), .B2(n9986), .A(n9987), .ZN(n14082) );
  NOR2_X1 U7328 ( .A1(n14008), .A2(n14138), .ZN(n13992) );
  AOI21_X1 U7329 ( .B1(n12860), .B2(n12167), .A(n12169), .ZN(n12851) );
  OAI21_X1 U7330 ( .B1(n8783), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n8416), .ZN(
        n8796) );
  NAND2_X1 U7331 ( .A1(n9984), .A2(n9983), .ZN(n11975) );
  NAND2_X1 U7332 ( .A1(n8416), .A2(n8415), .ZN(n8783) );
  NAND2_X1 U7333 ( .A1(n8098), .A2(n8097), .ZN(n14138) );
  NAND2_X1 U7334 ( .A1(n9287), .A2(n9286), .ZN(n13569) );
  NAND2_X1 U7335 ( .A1(n8071), .A2(n10022), .ZN(n8072) );
  NAND2_X1 U7336 ( .A1(n9261), .A2(n9260), .ZN(n13581) );
  OR2_X1 U7337 ( .A1(n11943), .A2(n11948), .ZN(n11945) );
  AND2_X1 U7338 ( .A1(n8138), .A2(n8118), .ZN(n8120) );
  NAND2_X1 U7339 ( .A1(n11365), .A2(n7306), .ZN(n7305) );
  NAND2_X1 U7340 ( .A1(n8028), .A2(n8027), .ZN(n14159) );
  AOI21_X1 U7341 ( .B1(n6713), .B2(n6503), .A(n6712), .ZN(n11707) );
  NAND2_X1 U7342 ( .A1(n8116), .A2(SI_24_), .ZN(n8138) );
  NAND2_X1 U7343 ( .A1(n11343), .A2(n11342), .ZN(n6858) );
  NAND2_X1 U7344 ( .A1(n8038), .A2(n8026), .ZN(n11437) );
  NOR2_X1 U7345 ( .A1(n9534), .A2(n9533), .ZN(n9535) );
  NAND2_X1 U7346 ( .A1(n12400), .A2(n6570), .ZN(n11075) );
  NAND2_X1 U7347 ( .A1(n7958), .A2(n7957), .ZN(n14172) );
  NAND2_X1 U7348 ( .A1(n10710), .A2(n10709), .ZN(n12397) );
  OR2_X2 U7349 ( .A1(n6495), .A2(n14456), .ZN(n14442) );
  NAND2_X1 U7350 ( .A1(n8687), .A2(n8686), .ZN(n12555) );
  NAND2_X1 U7351 ( .A1(n7801), .A2(n7800), .ZN(n14628) );
  OR2_X1 U7352 ( .A1(n7850), .A2(SI_14_), .ZN(n7888) );
  NOR2_X1 U7353 ( .A1(n15401), .A2(n14290), .ZN(n14293) );
  NAND2_X1 U7354 ( .A1(n9119), .A2(n9118), .ZN(n12391) );
  INV_X1 U7355 ( .A(n11512), .ZN(n14732) );
  NAND3_X1 U7356 ( .A1(n6793), .A2(n6792), .A3(n7846), .ZN(n7366) );
  OAI21_X1 U7357 ( .B1(n9865), .B2(P3_U3151), .A(n9864), .ZN(n12629) );
  NOR2_X1 U7358 ( .A1(n14322), .A2(n14286), .ZN(n14288) );
  NOR2_X2 U7359 ( .A1(n11837), .A2(n12925), .ZN(n10675) );
  NOR2_X1 U7360 ( .A1(n8774), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8786) );
  NAND2_X2 U7361 ( .A1(n9423), .A2(n13518), .ZN(n14919) );
  AND2_X1 U7362 ( .A1(n9490), .A2(n9489), .ZN(n7415) );
  XNOR2_X1 U7363 ( .A(n6653), .B(n13268), .ZN(n10363) );
  AND3_X1 U7364 ( .A1(n7647), .A2(n7646), .A3(n7645), .ZN(n14718) );
  NAND2_X1 U7365 ( .A1(n9056), .A2(n9055), .ZN(n10530) );
  CLKBUF_X1 U7366 ( .A(n9758), .Z(n9883) );
  INV_X4 U7367 ( .A(n9705), .ZN(n9686) );
  BUF_X1 U7368 ( .A(n11019), .Z(n6493) );
  BUF_X2 U7370 ( .A(n13098), .Z(n6725) );
  AND2_X1 U7371 ( .A1(n6917), .A2(n6795), .ZN(n6794) );
  INV_X4 U7372 ( .A(n12453), .ZN(n10922) );
  CLKBUF_X1 U7373 ( .A(n9475), .Z(n14950) );
  AOI21_X1 U7374 ( .B1(n6494), .B2(n7792), .A(n6587), .ZN(n6917) );
  CLKBUF_X1 U7375 ( .A(n12148), .Z(n8867) );
  AND2_X1 U7376 ( .A1(n9470), .A2(n9432), .ZN(n10212) );
  NOR2_X1 U7377 ( .A1(n6727), .A2(n11773), .ZN(n9475) );
  NAND2_X2 U7378 ( .A1(n6490), .A2(n10022), .ZN(n7670) );
  NAND2_X4 U7379 ( .A1(n13079), .A2(n7272), .ZN(n8482) );
  INV_X1 U7380 ( .A(n10469), .ZN(n10456) );
  AND2_X1 U7381 ( .A1(n6921), .A2(n6918), .ZN(n6494) );
  NAND2_X2 U7382 ( .A1(n9469), .A2(n6472), .ZN(n9478) );
  NAND2_X1 U7383 ( .A1(n8325), .A2(n14206), .ZN(n10079) );
  NAND3_X1 U7384 ( .A1(n14210), .A2(n9950), .A3(n11987), .ZN(n10469) );
  NAND2_X1 U7385 ( .A1(n8425), .A2(n8426), .ZN(n7272) );
  NAND2_X2 U7386 ( .A1(n12008), .A2(n8979), .ZN(n9671) );
  NAND2_X1 U7387 ( .A1(n8419), .A2(n6830), .ZN(n13079) );
  NAND2_X1 U7388 ( .A1(n9936), .A2(n11421), .ZN(n10453) );
  NAND2_X1 U7389 ( .A1(n6473), .A2(n10216), .ZN(n6727) );
  NAND2_X1 U7390 ( .A1(n14200), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7516) );
  MUX2_X1 U7391 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8418), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n8419) );
  NAND2_X1 U7392 ( .A1(n7517), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7518) );
  NAND2_X1 U7393 ( .A1(n7540), .A2(n7539), .ZN(n11421) );
  XNOR2_X1 U7394 ( .A(n8351), .B(n13065), .ZN(n8353) );
  AND2_X1 U7395 ( .A1(n8332), .A2(n6524), .ZN(n11987) );
  OR2_X1 U7396 ( .A1(n9375), .A2(n6606), .ZN(n9376) );
  AND2_X1 U7397 ( .A1(n9374), .A2(n9238), .ZN(n10216) );
  NAND2_X1 U7398 ( .A1(n13068), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8351) );
  XNOR2_X1 U7399 ( .A(n8327), .B(P1_IR_REG_26__SCAN_IN), .ZN(n14210) );
  NAND2_X1 U7400 ( .A1(n6738), .A2(n6735), .ZN(n13650) );
  NAND2_X1 U7401 ( .A1(n7539), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7537) );
  XNOR2_X1 U7402 ( .A(n7545), .B(n7544), .ZN(n8333) );
  XNOR2_X1 U7403 ( .A(n7217), .B(P1_IR_REG_22__SCAN_IN), .ZN(n10010) );
  NAND2_X1 U7404 ( .A1(n8975), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8977) );
  INV_X2 U7405 ( .A(n13070), .ZN(n13076) );
  NOR2_X1 U7406 ( .A1(n6737), .A2(n6736), .ZN(n6735) );
  AND2_X1 U7407 ( .A1(n8904), .A2(n8854), .ZN(n8940) );
  NAND2_X1 U7408 ( .A1(n8450), .A2(n8449), .ZN(n8666) );
  NAND2_X1 U7409 ( .A1(n6955), .A2(n7299), .ZN(n8422) );
  NAND2_X2 U7410 ( .A1(n10022), .A2(P2_U3088), .ZN(n13652) );
  AND2_X2 U7411 ( .A1(n9371), .A2(n9405), .ZN(n11773) );
  NAND2_X1 U7412 ( .A1(n7791), .A2(SI_10_), .ZN(n7814) );
  NAND2_X1 U7413 ( .A1(n7538), .A2(n7547), .ZN(n7539) );
  NAND2_X1 U7414 ( .A1(n6478), .A2(n6729), .ZN(n6738) );
  AND2_X1 U7415 ( .A1(n7542), .A2(n7544), .ZN(n7538) );
  NAND2_X1 U7416 ( .A1(n8985), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8984) );
  NAND2_X2 U7417 ( .A1(n8119), .A2(P2_U3088), .ZN(n13643) );
  NAND2_X2 U7418 ( .A1(n8119), .A2(P3_U3151), .ZN(n13078) );
  INV_X1 U7419 ( .A(n8859), .ZN(n6955) );
  AND2_X1 U7420 ( .A1(n6477), .A2(n9369), .ZN(n8972) );
  OAI21_X1 U7421 ( .B1(n7612), .B2(n10021), .A(n7560), .ZN(n7561) );
  NOR2_X1 U7422 ( .A1(n7546), .A2(n7551), .ZN(n7218) );
  NOR2_X1 U7423 ( .A1(n9130), .A2(n7318), .ZN(n7317) );
  NOR2_X1 U7424 ( .A1(n7955), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n7542) );
  AND2_X1 U7425 ( .A1(n7299), .A2(n6607), .ZN(n6753) );
  NOR2_X1 U7426 ( .A1(n9104), .A2(n6936), .ZN(n9369) );
  AND2_X1 U7427 ( .A1(n8350), .A2(n7300), .ZN(n7299) );
  NAND2_X1 U7428 ( .A1(n7397), .A2(n7514), .ZN(n7396) );
  CLKBUF_X1 U7429 ( .A(n9013), .Z(n9029) );
  AND4_X1 U7430 ( .A1(n9406), .A2(n9387), .A3(n8969), .A4(n8968), .ZN(n8970)
         );
  AND3_X1 U7431 ( .A1(n8963), .A2(n8964), .A3(n8962), .ZN(n9366) );
  AND4_X1 U7432 ( .A1(n7507), .A2(n7506), .A3(n7505), .A4(n7504), .ZN(n7508)
         );
  AND2_X1 U7433 ( .A1(n14274), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14272) );
  AND3_X1 U7434 ( .A1(n6953), .A2(n6952), .A3(n8684), .ZN(n6954) );
  AND4_X1 U7435 ( .A1(n8348), .A2(n8909), .A3(n8907), .A4(n8854), .ZN(n8420)
         );
  AND2_X1 U7436 ( .A1(n8967), .A2(n8966), .ZN(n9230) );
  NOR2_X1 U7437 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n7401) );
  NOR2_X1 U7438 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n8478) );
  INV_X4 U7439 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  OR2_X1 U7440 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6487) );
  INV_X4 U7441 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7442 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8854) );
  INV_X1 U7443 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7526) );
  INV_X1 U7444 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7527) );
  NOR2_X1 U7445 ( .A1(P3_IR_REG_11__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n8342) );
  NOR2_X1 U7446 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n8343) );
  NOR2_X1 U7447 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_6__SCAN_IN), .ZN(
        n8344) );
  NOR2_X1 U7448 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n6736) );
  INV_X1 U7449 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n7501) );
  INV_X1 U7450 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9406) );
  INV_X1 U7451 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9387) );
  INV_X1 U7452 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10039) );
  INV_X1 U7453 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n7608) );
  INV_X4 U7454 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X2 U7455 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n7403) );
  AND2_X1 U7456 ( .A1(n8974), .A2(n6546), .ZN(n6477) );
  NAND2_X1 U7457 ( .A1(n9369), .A2(n6546), .ZN(n6478) );
  AND3_X2 U7458 ( .A1(n8988), .A2(n9230), .A3(n8970), .ZN(n6546) );
  OR2_X1 U7459 ( .A1(n9195), .A2(n9007), .ZN(n9008) );
  CLKBUF_X1 U7460 ( .A(n9195), .Z(n6709) );
  NOR2_X1 U7461 ( .A1(n11010), .A2(n11153), .ZN(n11005) );
  AOI22_X1 U7462 ( .A1(n9187), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n10289), .B2(
        n9239), .ZN(n6949) );
  INV_X2 U7463 ( .A(n9663), .ZN(n9187) );
  INV_X1 U7464 ( .A(n14020), .ZN(n6479) );
  NAND2_X1 U7465 ( .A1(n9992), .A2(n7363), .ZN(n6480) );
  CLKBUF_X1 U7466 ( .A(n14636), .Z(n6481) );
  AND2_X1 U7467 ( .A1(n9894), .A2(n9895), .ZN(n6482) );
  NAND2_X1 U7468 ( .A1(n9992), .A2(n7363), .ZN(n14161) );
  NAND2_X1 U7469 ( .A1(n9970), .A2(n9969), .ZN(n14636) );
  NAND2_X2 U7470 ( .A1(n8978), .A2(n8979), .ZN(n9018) );
  NAND2_X2 U7471 ( .A1(n7072), .A2(n9832), .ZN(n9836) );
  NOR2_X2 U7472 ( .A1(n10673), .A2(n9769), .ZN(n10671) );
  NOR2_X2 U7473 ( .A1(n10671), .A2(n9771), .ZN(n10781) );
  NAND2_X1 U7474 ( .A1(n12613), .A2(n12614), .ZN(n7070) );
  XNOR2_X2 U7475 ( .A(n12059), .B(n12060), .ZN(n13805) );
  AND3_X2 U7476 ( .A1(n7401), .A2(n7402), .A3(n7400), .ZN(n8988) );
  INV_X8 U7477 ( .A(n7530), .ZN(n8119) );
  NAND2_X1 U7478 ( .A1(n7718), .A2(n7717), .ZN(n7739) );
  OR2_X1 U7479 ( .A1(n10071), .A2(n9664), .ZN(n9093) );
  NOR2_X2 U7480 ( .A1(n9130), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n9231) );
  OR2_X1 U7481 ( .A1(n9548), .A2(n9547), .ZN(n6508) );
  NAND2_X1 U7482 ( .A1(n11807), .A2(n6486), .ZN(n6483) );
  AND2_X1 U7483 ( .A1(n6483), .A2(n6484), .ZN(n7388) );
  OR2_X1 U7484 ( .A1(n6485), .A2(n9980), .ZN(n6484) );
  INV_X1 U7485 ( .A(n7389), .ZN(n6485) );
  AND2_X1 U7486 ( .A1(n11808), .A2(n7389), .ZN(n6486) );
  NOR2_X2 U7487 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n7558) );
  NAND4_X4 U7488 ( .A1(n9020), .A2(n9022), .A3(n9021), .A4(n9023), .ZN(n9477)
         );
  AND2_X2 U7489 ( .A1(n7744), .A2(n7508), .ZN(n6488) );
  INV_X1 U7490 ( .A(n6488), .ZN(n7903) );
  INV_X4 U7491 ( .A(n9687), .ZN(n9705) );
  INV_X1 U7492 ( .A(n9647), .ZN(n9687) );
  NAND2_X2 U7493 ( .A1(n9977), .A2(n9976), .ZN(n11650) );
  NOR2_X4 U7494 ( .A1(n14442), .A2(n14443), .ZN(n11702) );
  XNOR2_X2 U7495 ( .A(n11119), .B(n13842), .ZN(n11111) );
  NAND2_X1 U7496 ( .A1(n8325), .A2(n14206), .ZN(n6489) );
  NAND2_X1 U7497 ( .A1(n8325), .A2(n14206), .ZN(n6490) );
  NOR2_X4 U7498 ( .A1(n8328), .A2(n7394), .ZN(n7532) );
  NAND2_X2 U7499 ( .A1(n7558), .A2(n7502), .ZN(n7588) );
  NAND2_X1 U7500 ( .A1(n12527), .A2(n7522), .ZN(n6491) );
  NAND2_X1 U7501 ( .A1(n6489), .A2(n6720), .ZN(n7644) );
  OAI211_X1 U7502 ( .C1(n10079), .C2(n13847), .A(n7571), .B(n7570), .ZN(n11019) );
  OR2_X1 U7503 ( .A1(n13543), .A2(n13133), .ZN(n9356) );
  XOR2_X1 U7504 ( .A(n13241), .B(n13537), .Z(n9746) );
  NAND2_X1 U7505 ( .A1(n11600), .A2(n11599), .ZN(n7252) );
  OAI21_X1 U7506 ( .B1(n7127), .B2(n7123), .A(n7118), .ZN(n13353) );
  NOR2_X1 U7507 ( .A1(n7123), .A2(n7121), .ZN(n7120) );
  INV_X2 U7508 ( .A(n9664), .ZN(n9679) );
  INV_X2 U7509 ( .A(n7670), .ZN(n8282) );
  NOR2_X1 U7510 ( .A1(n7385), .A2(n7384), .ZN(n7383) );
  INV_X1 U7511 ( .A(n9532), .ZN(n6692) );
  INV_X1 U7512 ( .A(n9642), .ZN(n6700) );
  INV_X1 U7513 ( .A(n9655), .ZN(n6694) );
  NOR2_X1 U7514 ( .A1(n7149), .A2(n7153), .ZN(n7148) );
  INV_X1 U7515 ( .A(n8443), .ZN(n7153) );
  INV_X1 U7516 ( .A(n8458), .ZN(n7149) );
  NAND2_X1 U7517 ( .A1(n6783), .A2(n7901), .ZN(n7947) );
  OR2_X1 U7518 ( .A1(n7900), .A2(n7899), .ZN(n7901) );
  NAND2_X1 U7519 ( .A1(n6989), .A2(n14223), .ZN(n14224) );
  NAND2_X1 U7520 ( .A1(n14268), .A2(n14222), .ZN(n6989) );
  INV_X1 U7521 ( .A(n9760), .ZN(n9761) );
  OR2_X1 U7522 ( .A1(n12966), .A2(n12828), .ZN(n12341) );
  AND2_X1 U7523 ( .A1(n12624), .A2(n9831), .ZN(n12335) );
  INV_X1 U7524 ( .A(n13047), .ZN(n6978) );
  OR2_X1 U7525 ( .A1(n6750), .A2(n6749), .ZN(n6748) );
  INV_X1 U7526 ( .A(n6752), .ZN(n6749) );
  AND2_X1 U7527 ( .A1(n8679), .A2(n6551), .ZN(n6750) );
  AND2_X1 U7528 ( .A1(n8883), .A2(n12274), .ZN(n7284) );
  OR2_X1 U7529 ( .A1(n12673), .A2(n15134), .ZN(n12234) );
  NAND2_X1 U7530 ( .A1(n6804), .A2(n6803), .ZN(n12229) );
  INV_X1 U7531 ( .A(n15091), .ZN(n6804) );
  NAND2_X1 U7532 ( .A1(n9759), .A2(n10676), .ZN(n12217) );
  INV_X1 U7533 ( .A(n7157), .ZN(n7156) );
  OAI21_X1 U7534 ( .B1(n8624), .B2(n7158), .A(n8383), .ZN(n7157) );
  OAI21_X1 U7535 ( .B1(n8366), .B2(n7146), .A(n8527), .ZN(n7140) );
  NAND2_X1 U7536 ( .A1(n10058), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8369) );
  INV_X1 U7537 ( .A(n13175), .ZN(n6865) );
  NAND2_X1 U7538 ( .A1(n12515), .A2(n6854), .ZN(n6853) );
  INV_X1 U7539 ( .A(n12516), .ZN(n6854) );
  NAND2_X1 U7540 ( .A1(n7113), .A2(n6528), .ZN(n7112) );
  OR2_X1 U7541 ( .A1(n9157), .A2(n6553), .ZN(n7113) );
  OR2_X1 U7542 ( .A1(n13331), .A2(n7446), .ZN(n7100) );
  INV_X1 U7543 ( .A(n6936), .ZN(n6934) );
  AND2_X1 U7544 ( .A1(n11860), .A2(n6555), .ZN(n7259) );
  NOR2_X1 U7545 ( .A1(n14051), .A2(n7346), .ZN(n7345) );
  INV_X1 U7546 ( .A(n9921), .ZN(n7346) );
  INV_X1 U7547 ( .A(n11421), .ZN(n9937) );
  NOR2_X1 U7548 ( .A1(n14511), .A2(n6886), .ZN(n6885) );
  INV_X1 U7549 ( .A(n6887), .ZN(n6886) );
  NAND2_X1 U7550 ( .A1(n6932), .A2(n8154), .ZN(n8172) );
  NAND2_X1 U7551 ( .A1(n8139), .A2(n6566), .ZN(n6932) );
  NOR2_X1 U7552 ( .A1(n6526), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n7270) );
  NAND2_X1 U7553 ( .A1(n7615), .A2(n7634), .ZN(n7632) );
  OAI21_X1 U7554 ( .B1(n8119), .B2(n10018), .A(n7584), .ZN(n7631) );
  NAND2_X1 U7555 ( .A1(n8119), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7584) );
  XNOR2_X1 U7556 ( .A(n14228), .B(n15028), .ZN(n14264) );
  NAND2_X1 U7557 ( .A1(n15102), .A2(n12217), .ZN(n9766) );
  NAND2_X1 U7558 ( .A1(n6673), .A2(n6672), .ZN(n11882) );
  INV_X1 U7559 ( .A(n11885), .ZN(n6672) );
  INV_X1 U7560 ( .A(n8867), .ZN(n8789) );
  INV_X1 U7561 ( .A(n8510), .ZN(n8793) );
  BUF_X1 U7562 ( .A(n8778), .Z(n8865) );
  AND2_X1 U7563 ( .A1(n8353), .A2(n8355), .ZN(n8509) );
  OR2_X1 U7564 ( .A1(n11550), .A2(n11551), .ZN(n7008) );
  NOR2_X1 U7565 ( .A1(n12744), .A2(n7041), .ZN(n7039) );
  NOR2_X1 U7566 ( .A1(n14375), .A2(n12731), .ZN(n14391) );
  NAND2_X1 U7567 ( .A1(n6757), .A2(n6761), .ZN(n12896) );
  NAND2_X1 U7568 ( .A1(n12920), .A2(n6764), .ZN(n6757) );
  NAND2_X1 U7569 ( .A1(n8482), .A2(n10022), .ZN(n8760) );
  NAND2_X1 U7570 ( .A1(n6475), .A2(n6976), .ZN(n8485) );
  OR2_X1 U7571 ( .A1(n13017), .A2(n8840), .ZN(n7489) );
  NAND2_X1 U7572 ( .A1(n8902), .A2(n14415), .ZN(n8903) );
  INV_X1 U7573 ( .A(n8529), .ZN(n8814) );
  INV_X1 U7574 ( .A(n7301), .ZN(n7300) );
  AND2_X1 U7575 ( .A1(n8349), .A2(n8420), .ZN(n8350) );
  NAND2_X1 U7576 ( .A1(n10087), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8382) );
  NAND2_X1 U7577 ( .A1(n8559), .A2(n8373), .ZN(n7165) );
  NAND2_X1 U7578 ( .A1(n10056), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8367) );
  NAND2_X1 U7579 ( .A1(n9365), .A2(n9364), .ZN(n13537) );
  AND2_X1 U7580 ( .A1(n9356), .A2(n9354), .ZN(n13332) );
  AND2_X1 U7581 ( .A1(n7128), .A2(n9723), .ZN(n7127) );
  INV_X1 U7582 ( .A(n7469), .ZN(n7468) );
  OAI21_X1 U7583 ( .B1(n7471), .B2(n13391), .A(n7473), .ZN(n7469) );
  NOR2_X1 U7584 ( .A1(n13405), .A2(n9296), .ZN(n13390) );
  NOR2_X1 U7585 ( .A1(n7477), .A2(n7476), .ZN(n7475) );
  INV_X1 U7586 ( .A(n9459), .ZN(n7476) );
  OAI21_X1 U7587 ( .B1(n7088), .B2(n7090), .A(n7086), .ZN(n9142) );
  AOI21_X1 U7588 ( .B1(n7089), .B2(n7092), .A(n7087), .ZN(n7086) );
  AND2_X1 U7589 ( .A1(n9116), .A2(n9115), .ZN(n10991) );
  INV_X2 U7590 ( .A(n10098), .ZN(n9239) );
  AND2_X1 U7591 ( .A1(n9731), .A2(n9442), .ZN(n7465) );
  NAND2_X1 U7592 ( .A1(n9378), .A2(n9377), .ZN(n14886) );
  AND2_X1 U7593 ( .A1(n7450), .A2(n9746), .ZN(n7438) );
  NAND2_X1 U7594 ( .A1(n7444), .A2(n7443), .ZN(n7442) );
  NAND2_X1 U7595 ( .A1(n7448), .A2(n7446), .ZN(n7443) );
  OAI21_X1 U7596 ( .B1(n7450), .B2(n9746), .A(n7447), .ZN(n7444) );
  INV_X1 U7597 ( .A(n13344), .ZN(n13543) );
  NAND2_X1 U7598 ( .A1(n9333), .A2(n9332), .ZN(n13547) );
  AND2_X1 U7599 ( .A1(n8988), .A2(n9230), .ZN(n9370) );
  NAND2_X1 U7600 ( .A1(n11593), .A2(n7252), .ZN(n7249) );
  NAND2_X1 U7601 ( .A1(n6595), .A2(n7252), .ZN(n7248) );
  OR2_X1 U7602 ( .A1(n11505), .A2(n7251), .ZN(n7250) );
  NAND2_X1 U7603 ( .A1(n8239), .A2(n8238), .ZN(n13929) );
  OR2_X1 U7604 ( .A1(n9665), .A2(n7670), .ZN(n8239) );
  NAND2_X1 U7605 ( .A1(n12475), .A2(n8294), .ZN(n12024) );
  NAND2_X1 U7606 ( .A1(n14126), .A2(n12019), .ZN(n13962) );
  AOI21_X1 U7607 ( .B1(n7372), .B2(n13983), .A(n6557), .ZN(n7370) );
  INV_X1 U7608 ( .A(n7372), .ZN(n7371) );
  NAND2_X1 U7609 ( .A1(n7992), .A2(n7991), .ZN(n14062) );
  INV_X1 U7610 ( .A(n14048), .ZN(n14051) );
  OR2_X1 U7611 ( .A1(n14511), .A2(n13807), .ZN(n9915) );
  INV_X1 U7612 ( .A(n6492), .ZN(n7990) );
  INV_X1 U7613 ( .A(n10079), .ZN(n7989) );
  NOR2_X1 U7614 ( .A1(n7218), .A2(n14199), .ZN(n7217) );
  NAND2_X1 U7615 ( .A1(n6897), .A2(n6895), .ZN(n7767) );
  AOI21_X1 U7616 ( .B1(n6898), .B2(n6900), .A(n6896), .ZN(n6895) );
  INV_X1 U7617 ( .A(n7762), .ZN(n6896) );
  NAND2_X1 U7618 ( .A1(n15394), .A2(n14279), .ZN(n14281) );
  OAI21_X1 U7619 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n14244), .A(n14243), .ZN(
        n14258) );
  INV_X1 U7620 ( .A(n12887), .ZN(n12862) );
  AND2_X1 U7621 ( .A1(P3_U3897), .A2(n13079), .ZN(n15078) );
  AOI21_X1 U7622 ( .B1(n13635), .B2(n8282), .A(n8281), .ZN(n14091) );
  INV_X1 U7623 ( .A(n9497), .ZN(n6705) );
  OAI21_X1 U7624 ( .B1(n7650), .B2(n7649), .A(n7648), .ZN(n7680) );
  INV_X1 U7625 ( .A(n7703), .ZN(n7177) );
  OR2_X1 U7626 ( .A1(n7753), .A2(n7207), .ZN(n7206) );
  INV_X1 U7627 ( .A(n7751), .ZN(n7207) );
  NOR2_X1 U7628 ( .A1(n7754), .A2(n7751), .ZN(n7208) );
  INV_X1 U7629 ( .A(n9558), .ZN(n6683) );
  AOI21_X1 U7630 ( .B1(n7202), .B2(n7200), .A(n7199), .ZN(n7198) );
  NAND2_X1 U7631 ( .A1(n7195), .A2(n7844), .ZN(n7193) );
  AND2_X1 U7632 ( .A1(n7984), .A2(n7216), .ZN(n7215) );
  INV_X1 U7633 ( .A(n7943), .ZN(n7216) );
  AND2_X1 U7634 ( .A1(n14048), .A2(n8000), .ZN(n8004) );
  AND2_X1 U7635 ( .A1(n7985), .A2(n7213), .ZN(n7212) );
  NAND2_X1 U7636 ( .A1(n7214), .A2(n7943), .ZN(n7213) );
  AND2_X1 U7637 ( .A1(n14072), .A2(n7982), .ZN(n7985) );
  NAND2_X1 U7638 ( .A1(n6586), .A2(n7412), .ZN(n7408) );
  NAND2_X1 U7639 ( .A1(n8073), .A2(n7181), .ZN(n7178) );
  NAND2_X1 U7640 ( .A1(n7423), .A2(n6561), .ZN(n7422) );
  INV_X1 U7641 ( .A(n9651), .ZN(n7427) );
  INV_X1 U7642 ( .A(n9657), .ZN(n6689) );
  NOR2_X1 U7643 ( .A1(n12160), .A2(n12161), .ZN(n7297) );
  AND2_X1 U7644 ( .A1(n12938), .A2(n12164), .ZN(n12162) );
  INV_X1 U7645 ( .A(n8400), .ZN(n7152) );
  INV_X1 U7646 ( .A(n9200), .ZN(n7105) );
  AND2_X1 U7647 ( .A1(n7491), .A2(n6907), .ZN(n6904) );
  NAND2_X1 U7648 ( .A1(n6908), .A2(n8115), .ZN(n6907) );
  INV_X1 U7649 ( .A(n8093), .ZN(n6908) );
  XNOR2_X1 U7650 ( .A(n12624), .B(n9838), .ZN(n9828) );
  OR2_X1 U7651 ( .A1(n8472), .A2(n10745), .ZN(n8473) );
  OR2_X1 U7652 ( .A1(n8510), .A2(n15113), .ZN(n8474) );
  INV_X1 U7653 ( .A(n10908), .ZN(n7033) );
  NOR2_X1 U7654 ( .A1(n10757), .A2(n10726), .ZN(n7031) );
  NAND2_X1 U7655 ( .A1(n14994), .A2(n6567), .ZN(n10843) );
  NOR2_X1 U7656 ( .A1(n14380), .A2(n8471), .ZN(n7041) );
  NOR2_X1 U7657 ( .A1(n6506), .A2(n6968), .ZN(n6963) );
  OR2_X1 U7658 ( .A1(n12578), .A2(n12829), .ZN(n12349) );
  OR2_X1 U7659 ( .A1(n12834), .A2(n12654), .ZN(n8794) );
  NOR2_X1 U7660 ( .A1(n8788), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8802) );
  INV_X1 U7661 ( .A(n12826), .ZN(n8891) );
  NOR2_X1 U7662 ( .A1(n12207), .A2(n6822), .ZN(n6821) );
  INV_X1 U7663 ( .A(n8888), .ZN(n6822) );
  NAND2_X1 U7664 ( .A1(n6761), .A2(n6759), .ZN(n6758) );
  INV_X1 U7665 ( .A(n6764), .ZN(n6759) );
  NAND2_X1 U7666 ( .A1(n6538), .A2(n6760), .ZN(n6756) );
  INV_X1 U7667 ( .A(n6761), .ZN(n6760) );
  NOR2_X1 U7668 ( .A1(n6763), .A2(n12921), .ZN(n7287) );
  OR2_X1 U7669 ( .A1(n12666), .A2(n11836), .ZN(n12273) );
  XNOR2_X1 U7670 ( .A(n12670), .B(n6766), .ZN(n11409) );
  XNOR2_X1 U7671 ( .A(n9772), .B(n15088), .ZN(n15093) );
  AND2_X1 U7672 ( .A1(n11034), .A2(n11194), .ZN(n6972) );
  OR2_X1 U7673 ( .A1(n8414), .A2(n11912), .ZN(n8416) );
  INV_X1 U7674 ( .A(n8382), .ZN(n7158) );
  NAND2_X1 U7675 ( .A1(n10082), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8380) );
  NAND2_X1 U7676 ( .A1(n10073), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8378) );
  NAND2_X1 U7677 ( .A1(n10068), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8376) );
  INV_X1 U7678 ( .A(n8367), .ZN(n7146) );
  INV_X1 U7679 ( .A(n8369), .ZN(n7142) );
  AND2_X1 U7680 ( .A1(n9120), .A2(n8956), .ZN(n9151) );
  NOR2_X1 U7681 ( .A1(n9319), .A2(n7126), .ZN(n7125) );
  INV_X1 U7682 ( .A(n6521), .ZN(n7126) );
  NAND2_X1 U7683 ( .A1(n9462), .A2(n9463), .ZN(n7464) );
  NAND2_X1 U7684 ( .A1(n13331), .A2(n7102), .ZN(n7101) );
  NOR2_X1 U7685 ( .A1(n9746), .A2(n7103), .ZN(n7102) );
  NOR2_X1 U7686 ( .A1(n6502), .A2(n9386), .ZN(n7097) );
  AND2_X1 U7687 ( .A1(n13537), .A2(n14945), .ZN(n6943) );
  NOR2_X1 U7688 ( .A1(n13332), .A2(n13354), .ZN(n7450) );
  NOR2_X1 U7689 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n8967) );
  INV_X1 U7690 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n7319) );
  AOI21_X1 U7691 ( .B1(n12101), .B2(n12098), .A(n13669), .ZN(n7236) );
  INV_X1 U7692 ( .A(n12101), .ZN(n7237) );
  INV_X1 U7693 ( .A(n7230), .ZN(n7229) );
  NOR2_X1 U7694 ( .A1(n13967), .A2(n6874), .ZN(n6873) );
  INV_X1 U7695 ( .A(n6875), .ZN(n6874) );
  INV_X1 U7696 ( .A(n9997), .ZN(n7355) );
  INV_X1 U7697 ( .A(n14022), .ZN(n9994) );
  NOR2_X1 U7698 ( .A1(n14518), .A2(n11900), .ZN(n6887) );
  NOR2_X1 U7699 ( .A1(n11688), .A2(n11659), .ZN(n7326) );
  INV_X1 U7700 ( .A(n9978), .ZN(n7328) );
  INV_X1 U7701 ( .A(n6523), .ZN(n7379) );
  NOR2_X1 U7702 ( .A1(n9907), .A2(n9971), .ZN(n7334) );
  INV_X1 U7703 ( .A(n9972), .ZN(n7336) );
  NAND2_X1 U7704 ( .A1(n14732), .A2(n11494), .ZN(n6881) );
  NAND2_X1 U7705 ( .A1(n6550), .A2(n9902), .ZN(n7360) );
  NAND2_X1 U7706 ( .A1(n9894), .A2(n9895), .ZN(n6660) );
  AOI21_X1 U7707 ( .B1(n7342), .B2(n7341), .A(n6580), .ZN(n7340) );
  INV_X1 U7708 ( .A(n7345), .ZN(n7341) );
  NAND2_X1 U7709 ( .A1(n8226), .A2(n8225), .ZN(n8234) );
  NAND2_X1 U7710 ( .A1(n8173), .A2(SI_26_), .ZN(n8174) );
  NAND2_X1 U7711 ( .A1(n6929), .A2(n6924), .ZN(n8171) );
  NAND2_X1 U7712 ( .A1(n7513), .A2(n7399), .ZN(n7398) );
  INV_X1 U7713 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n7399) );
  OR2_X1 U7714 ( .A1(n8095), .A2(SI_22_), .ZN(n8070) );
  AND2_X1 U7715 ( .A1(n8025), .A2(n6628), .ZN(n7375) );
  OAI21_X1 U7716 ( .B1(n8023), .B2(n8022), .A(n8021), .ZN(n8024) );
  INV_X1 U7717 ( .A(n6916), .ZN(n6915) );
  OAI21_X1 U7718 ( .B1(n15327), .B2(n7946), .A(n7976), .ZN(n6916) );
  INV_X1 U7719 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n7536) );
  INV_X1 U7720 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n7271) );
  INV_X1 U7721 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n7504) );
  INV_X1 U7722 ( .A(n7790), .ZN(n6920) );
  AOI21_X1 U7723 ( .B1(n7793), .B2(n6923), .A(n6922), .ZN(n6921) );
  INV_X1 U7724 ( .A(n7814), .ZN(n6922) );
  INV_X1 U7725 ( .A(n7789), .ZN(n6923) );
  XNOR2_X1 U7726 ( .A(n7835), .B(SI_11_), .ZN(n7837) );
  INV_X1 U7727 ( .A(n7687), .ZN(n6785) );
  AOI21_X1 U7728 ( .B1(n7687), .B2(n6789), .A(n6788), .ZN(n6787) );
  INV_X1 U7729 ( .A(n7713), .ZN(n6788) );
  INV_X1 U7730 ( .A(n7683), .ZN(n6789) );
  AND2_X2 U7731 ( .A1(n6782), .A2(n6780), .ZN(n7612) );
  INV_X1 U7732 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n6781) );
  XNOR2_X1 U7733 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n14271) );
  NAND2_X1 U7734 ( .A1(n6657), .A2(n6991), .ZN(n14221) );
  NAND2_X1 U7735 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n6992), .ZN(n6991) );
  INV_X1 U7736 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6992) );
  XNOR2_X1 U7737 ( .A(n14224), .B(n15009), .ZN(n14265) );
  OAI21_X1 U7738 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n14238), .A(n14237), .ZN(
        n14262) );
  AOI21_X1 U7739 ( .B1(n7068), .B2(n9850), .A(n6584), .ZN(n7065) );
  OR2_X1 U7740 ( .A1(n12641), .A2(n9850), .ZN(n7066) );
  AOI21_X1 U7741 ( .B1(n7075), .B2(n7074), .A(n6577), .ZN(n7073) );
  INV_X1 U7742 ( .A(n11357), .ZN(n7074) );
  AND2_X1 U7743 ( .A1(n9851), .A2(n7069), .ZN(n7068) );
  OR2_X1 U7744 ( .A1(n12641), .A2(n9850), .ZN(n7069) );
  NAND2_X1 U7745 ( .A1(n9761), .A2(n8498), .ZN(n9763) );
  NOR2_X1 U7746 ( .A1(n11579), .A2(n6507), .ZN(n7053) );
  INV_X1 U7747 ( .A(n12665), .ZN(n12280) );
  NAND2_X1 U7748 ( .A1(n9830), .A2(n9831), .ZN(n7072) );
  NAND2_X1 U7749 ( .A1(n9794), .A2(n7060), .ZN(n7059) );
  NAND2_X1 U7750 ( .A1(n11581), .A2(n9794), .ZN(n7055) );
  XNOR2_X1 U7751 ( .A(n9777), .B(n15088), .ZN(n9773) );
  NAND2_X1 U7752 ( .A1(n12544), .A2(n9807), .ZN(n7048) );
  OR2_X1 U7753 ( .A1(n11926), .A2(n6534), .ZN(n7050) );
  XNOR2_X1 U7754 ( .A(n7295), .B(n8454), .ZN(n12197) );
  INV_X1 U7755 ( .A(n8865), .ZN(n8830) );
  OAI21_X1 U7756 ( .B1(n8510), .B2(P3_REG3_REG_3__SCAN_IN), .A(n8513), .ZN(
        n6806) );
  INV_X1 U7757 ( .A(n12148), .ZN(n6739) );
  XNOR2_X1 U7758 ( .A(n10843), .B(n10824), .ZN(n15016) );
  NAND2_X1 U7759 ( .A1(n15016), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n15015) );
  NAND2_X1 U7760 ( .A1(n7001), .A2(n7000), .ZN(n15072) );
  OR2_X1 U7761 ( .A1(n12678), .A2(n12690), .ZN(n6770) );
  AOI21_X1 U7762 ( .B1(n12736), .B2(n12735), .A(n12734), .ZN(n14353) );
  AND2_X1 U7763 ( .A1(n12726), .A2(n7011), .ZN(n7012) );
  INV_X1 U7764 ( .A(n14359), .ZN(n7011) );
  OR2_X1 U7765 ( .A1(n12706), .A2(n12707), .ZN(n7015) );
  INV_X1 U7766 ( .A(n12726), .ZN(n7014) );
  OR2_X1 U7767 ( .A1(n12706), .A2(n7013), .ZN(n6773) );
  OR2_X1 U7768 ( .A1(n14359), .A2(n12707), .ZN(n7013) );
  XNOR2_X1 U7769 ( .A(n12753), .B(n12755), .ZN(n14367) );
  NAND2_X1 U7770 ( .A1(n14367), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n14366) );
  AND2_X1 U7771 ( .A1(n12349), .A2(n12350), .ZN(n12813) );
  NAND2_X1 U7772 ( .A1(n8892), .A2(n8891), .ZN(n12824) );
  INV_X1 U7773 ( .A(n12822), .ZN(n8892) );
  NOR2_X1 U7774 ( .A1(n12335), .A2(n6819), .ZN(n6818) );
  NAND2_X1 U7775 ( .A1(n6741), .A2(n6554), .ZN(n12841) );
  NAND2_X1 U7776 ( .A1(n12851), .A2(n6742), .ZN(n6741) );
  OR2_X1 U7777 ( .A1(n12624), .A2(n12656), .ZN(n6742) );
  INV_X1 U7778 ( .A(n12336), .ZN(n12840) );
  AND2_X1 U7779 ( .A1(n12170), .A2(n12333), .ZN(n12854) );
  OR2_X1 U7780 ( .A1(n12169), .A2(n12168), .ZN(n12864) );
  AOI21_X1 U7781 ( .B1(n12866), .B2(n8793), .A(n8769), .ZN(n12874) );
  AOI21_X1 U7782 ( .B1(n12900), .B2(n6532), .A(n6825), .ZN(n6824) );
  OR2_X1 U7783 ( .A1(n12635), .A2(n12911), .ZN(n12311) );
  OR2_X1 U7784 ( .A1(n12896), .A2(n12897), .ZN(n6980) );
  NAND2_X1 U7785 ( .A1(n6956), .A2(n6629), .ZN(n12920) );
  NAND2_X1 U7786 ( .A1(n11915), .A2(n6630), .ZN(n6956) );
  NAND2_X1 U7787 ( .A1(n12929), .A2(n6765), .ZN(n12928) );
  OR2_X1 U7788 ( .A1(n6747), .A2(n6533), .ZN(n6746) );
  INV_X1 U7789 ( .A(n6748), .ZN(n6747) );
  NAND2_X1 U7790 ( .A1(n6745), .A2(n6748), .ZN(n11844) );
  NAND2_X1 U7791 ( .A1(n11760), .A2(n6533), .ZN(n6745) );
  NAND2_X1 U7792 ( .A1(n12182), .A2(n7284), .ZN(n6810) );
  NOR2_X1 U7793 ( .A1(n12287), .A2(n6535), .ZN(n7282) );
  INV_X1 U7794 ( .A(n7284), .ZN(n6811) );
  NAND2_X1 U7795 ( .A1(n11763), .A2(n7284), .ZN(n7283) );
  NAND2_X1 U7796 ( .A1(n11765), .A2(n11764), .ZN(n11763) );
  AOI21_X1 U7797 ( .B1(n6572), .B2(n11329), .A(n7279), .ZN(n7278) );
  NOR2_X1 U7798 ( .A1(n8879), .A2(n15161), .ZN(n7279) );
  INV_X1 U7799 ( .A(n8879), .ZN(n7281) );
  NOR2_X1 U7800 ( .A1(n11329), .A2(n11516), .ZN(n7280) );
  INV_X1 U7801 ( .A(n12257), .ZN(n8616) );
  INV_X1 U7802 ( .A(n15103), .ZN(n12927) );
  NAND2_X1 U7803 ( .A1(n8801), .A2(n8800), .ZN(n9848) );
  AND2_X1 U7804 ( .A1(n8863), .A2(n12370), .ZN(n15104) );
  CLKBUF_X1 U7805 ( .A(n8920), .Z(n8914) );
  NAND2_X1 U7806 ( .A1(n7166), .A2(n7167), .ZN(n8842) );
  AOI21_X1 U7807 ( .B1(n7168), .B2(n8810), .A(n6646), .ZN(n7167) );
  NOR2_X1 U7808 ( .A1(n8424), .A2(n8423), .ZN(n8425) );
  NAND2_X1 U7809 ( .A1(n8421), .A2(n6734), .ZN(n8426) );
  NOR2_X1 U7810 ( .A1(P3_IR_REG_27__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n8423) );
  NAND2_X1 U7811 ( .A1(n8759), .A2(n8407), .ZN(n8430) );
  AND2_X1 U7812 ( .A1(n8402), .A2(n8401), .ZN(n8443) );
  NAND2_X1 U7813 ( .A1(n8730), .A2(n8398), .ZN(n8459) );
  NAND2_X1 U7814 ( .A1(n8459), .A2(n8458), .ZN(n8461) );
  NAND2_X1 U7815 ( .A1(n8728), .A2(n8727), .ZN(n8730) );
  INV_X1 U7816 ( .A(n8695), .ZN(n7173) );
  OR2_X1 U7817 ( .A1(n8681), .A2(n8391), .ZN(n7174) );
  AND2_X1 U7818 ( .A1(n8382), .A2(n8381), .ZN(n8624) );
  NAND2_X1 U7819 ( .A1(n8611), .A2(n8380), .ZN(n8625) );
  NAND2_X1 U7820 ( .A1(n8625), .A2(n8624), .ZN(n8627) );
  NOR2_X1 U7821 ( .A1(n8571), .A2(n7164), .ZN(n7163) );
  INV_X1 U7822 ( .A(n8374), .ZN(n7164) );
  NAND2_X1 U7823 ( .A1(n8372), .A2(n8371), .ZN(n8559) );
  AND2_X1 U7824 ( .A1(n8369), .A2(n8368), .ZN(n8527) );
  NAND2_X1 U7825 ( .A1(n8367), .A2(n8365), .ZN(n8514) );
  NAND2_X1 U7826 ( .A1(n8364), .A2(n8363), .ZN(n8515) );
  NAND2_X1 U7827 ( .A1(n6848), .A2(n6847), .ZN(n8480) );
  NAND2_X1 U7828 ( .A1(n7294), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6847) );
  OAI21_X1 U7829 ( .B1(n6849), .B2(n8612), .A(P3_IR_REG_1__SCAN_IN), .ZN(n6848) );
  INV_X1 U7830 ( .A(n13122), .ZN(n7312) );
  OR2_X1 U7831 ( .A1(n12499), .A2(n12500), .ZN(n6867) );
  NOR2_X1 U7832 ( .A1(n9746), .A2(n7332), .ZN(n7331) );
  NAND2_X1 U7833 ( .A1(n9744), .A2(n13354), .ZN(n7332) );
  INV_X1 U7834 ( .A(n9696), .ZN(n9745) );
  AND2_X1 U7835 ( .A1(n9353), .A2(n9352), .ZN(n13133) );
  INV_X1 U7836 ( .A(n9671), .ZN(n9246) );
  OR2_X1 U7837 ( .A1(n9176), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n9201) );
  OR2_X1 U7838 ( .A1(n7129), .A2(n9319), .ZN(n7128) );
  NOR2_X1 U7839 ( .A1(n13380), .A2(n6569), .ZN(n7129) );
  AND2_X1 U7840 ( .A1(n13401), .A2(n13246), .ZN(n9467) );
  NAND2_X1 U7841 ( .A1(n13380), .A2(n7472), .ZN(n7471) );
  INV_X1 U7842 ( .A(n9467), .ZN(n7472) );
  NOR2_X1 U7843 ( .A1(n13395), .A2(n13396), .ZN(n13394) );
  AND2_X1 U7844 ( .A1(n13575), .A2(n13248), .ZN(n9466) );
  NOR2_X1 U7845 ( .A1(n13413), .A2(n13406), .ZN(n6790) );
  OR2_X1 U7846 ( .A1(n9229), .A2(n7133), .ZN(n7131) );
  NAND2_X1 U7847 ( .A1(n7137), .A2(n7138), .ZN(n7133) );
  OR2_X1 U7848 ( .A1(n6560), .A2(n7134), .ZN(n7132) );
  INV_X1 U7849 ( .A(n7138), .ZN(n7134) );
  NAND2_X1 U7850 ( .A1(n7137), .A2(n9250), .ZN(n7136) );
  OR2_X1 U7851 ( .A1(n13600), .A2(n13218), .ZN(n7083) );
  NAND2_X1 U7852 ( .A1(n7479), .A2(n7478), .ZN(n13501) );
  AOI21_X1 U7853 ( .B1(n7480), .B2(n11708), .A(n6548), .ZN(n7478) );
  NAND2_X1 U7854 ( .A1(n13501), .A2(n13500), .ZN(n13499) );
  NOR2_X1 U7855 ( .A1(n13515), .A2(n7481), .ZN(n7480) );
  INV_X1 U7856 ( .A(n9458), .ZN(n7481) );
  OR2_X1 U7857 ( .A1(n11701), .A2(n11708), .ZN(n11699) );
  INV_X1 U7858 ( .A(n7112), .ZN(n7110) );
  AOI21_X1 U7859 ( .B1(n7109), .B2(n7115), .A(n7107), .ZN(n7106) );
  INV_X1 U7860 ( .A(n9725), .ZN(n7107) );
  NAND2_X1 U7861 ( .A1(n11267), .A2(n11270), .ZN(n7117) );
  NAND2_X1 U7862 ( .A1(n9453), .A2(n9452), .ZN(n11316) );
  NAND2_X1 U7863 ( .A1(n7456), .A2(n7455), .ZN(n9453) );
  AND2_X1 U7864 ( .A1(n7457), .A2(n6605), .ZN(n7455) );
  INV_X1 U7865 ( .A(n9734), .ZN(n11270) );
  NAND2_X1 U7866 ( .A1(n10990), .A2(n10991), .ZN(n10989) );
  NAND2_X1 U7867 ( .A1(n11159), .A2(n9440), .ZN(n7466) );
  NAND2_X1 U7868 ( .A1(n9037), .A2(n9036), .ZN(n10507) );
  XNOR2_X1 U7869 ( .A(n14906), .B(n13267), .ZN(n10508) );
  NAND2_X1 U7870 ( .A1(n10264), .A2(n9476), .ZN(n10263) );
  CLKBUF_X1 U7871 ( .A(n10212), .Z(n9471) );
  NAND2_X1 U7872 ( .A1(n13538), .A2(n7096), .ZN(n7095) );
  INV_X1 U7873 ( .A(n7098), .ZN(n7096) );
  INV_X1 U7874 ( .A(n7445), .ZN(n7441) );
  INV_X1 U7875 ( .A(n13542), .ZN(n6718) );
  OR2_X1 U7876 ( .A1(n11547), .A2(n9664), .ZN(n9261) );
  OR2_X1 U7877 ( .A1(n11437), .A2(n9664), .ZN(n9252) );
  OR2_X1 U7878 ( .A1(n10089), .A2(n9664), .ZN(n9134) );
  NAND2_X1 U7879 ( .A1(n10218), .A2(n10217), .ZN(n14945) );
  INV_X1 U7880 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7320) );
  OR2_X1 U7881 ( .A1(n9064), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n9090) );
  OR2_X1 U7882 ( .A1(n9040), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n9051) );
  INV_X1 U7883 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9024) );
  OR2_X1 U7884 ( .A1(n8061), .A2(n12105), .ZN(n8077) );
  OR2_X1 U7885 ( .A1(n7971), .A2(n7960), .ZN(n7994) );
  NAND2_X1 U7886 ( .A1(n7226), .A2(n7229), .ZN(n7223) );
  AND2_X1 U7887 ( .A1(n13784), .A2(n7227), .ZN(n7226) );
  NAND2_X1 U7888 ( .A1(n7230), .A2(n7228), .ZN(n7227) );
  INV_X1 U7889 ( .A(n13736), .ZN(n7228) );
  NAND2_X1 U7890 ( .A1(n13792), .A2(n12440), .ZN(n13658) );
  AOI21_X1 U7891 ( .B1(n7248), .B2(n7249), .A(n7246), .ZN(n7245) );
  INV_X1 U7892 ( .A(n11602), .ZN(n7246) );
  INV_X1 U7893 ( .A(n7259), .ZN(n7258) );
  AOI21_X1 U7894 ( .B1(n7259), .B2(n7257), .A(n6588), .ZN(n7256) );
  INV_X1 U7895 ( .A(n11857), .ZN(n7257) );
  NAND2_X1 U7896 ( .A1(n11858), .A2(n11857), .ZN(n7260) );
  NAND2_X1 U7897 ( .A1(n7260), .A2(n7259), .ZN(n11902) );
  NAND2_X1 U7898 ( .A1(n13723), .A2(n13724), .ZN(n13722) );
  NOR2_X1 U7899 ( .A1(n8232), .A2(n8229), .ZN(n6889) );
  INV_X1 U7900 ( .A(n8229), .ZN(n6888) );
  NAND2_X1 U7901 ( .A1(n7183), .A2(n7182), .ZN(n8230) );
  NAND2_X1 U7902 ( .A1(n13964), .A2(n7376), .ZN(n13947) );
  AND2_X1 U7903 ( .A1(n13940), .A2(n12020), .ZN(n7376) );
  AND2_X1 U7904 ( .A1(n10004), .A2(n9930), .ZN(n7372) );
  NAND2_X1 U7905 ( .A1(n9929), .A2(n9928), .ZN(n13974) );
  INV_X1 U7906 ( .A(n13997), .ZN(n6661) );
  NAND2_X1 U7907 ( .A1(n14021), .A2(n6527), .ZN(n14005) );
  OR2_X1 U7908 ( .A1(n14159), .A2(n14058), .ZN(n14041) );
  NAND2_X1 U7909 ( .A1(n14071), .A2(n7345), .ZN(n7344) );
  OR2_X1 U7910 ( .A1(n11949), .A2(n13719), .ZN(n11976) );
  NAND2_X1 U7911 ( .A1(n11945), .A2(n6564), .ZN(n11971) );
  AND4_X1 U7912 ( .A1(n7913), .A2(n7912), .A3(n7911), .A4(n7910), .ZN(n13714)
         );
  NOR2_X1 U7913 ( .A1(n11870), .A2(n7390), .ZN(n7389) );
  INV_X1 U7914 ( .A(n9982), .ZN(n7390) );
  AND4_X1 U7915 ( .A1(n7867), .A2(n7866), .A3(n7865), .A4(n7864), .ZN(n13807)
         );
  NAND2_X1 U7916 ( .A1(n7347), .A2(n7350), .ZN(n11869) );
  INV_X1 U7917 ( .A(n7351), .ZN(n7350) );
  OAI21_X1 U7918 ( .B1(n14475), .B2(n7352), .A(n11870), .ZN(n7351) );
  AND2_X1 U7919 ( .A1(n9915), .A2(n7914), .ZN(n14475) );
  NAND2_X1 U7920 ( .A1(n11817), .A2(n9914), .ZN(n14476) );
  NAND2_X1 U7921 ( .A1(n14476), .A2(n14475), .ZN(n14474) );
  NAND2_X1 U7922 ( .A1(n6470), .A2(n6523), .ZN(n14617) );
  NAND2_X1 U7923 ( .A1(n7772), .A2(n7771), .ZN(n11674) );
  INV_X1 U7924 ( .A(n7360), .ZN(n7361) );
  INV_X1 U7925 ( .A(n14055), .ZN(n14631) );
  NAND2_X1 U7926 ( .A1(n8043), .A2(n8042), .ZN(n14151) );
  AND2_X1 U7927 ( .A1(n14033), .A2(n9991), .ZN(n7363) );
  NAND2_X1 U7928 ( .A1(n7859), .A2(n7858), .ZN(n14511) );
  NAND2_X1 U7929 ( .A1(n9932), .A2(n9931), .ZN(n14618) );
  AND2_X1 U7930 ( .A1(n14655), .A2(n10459), .ZN(n14755) );
  AND2_X1 U7931 ( .A1(n14730), .A2(n14743), .ZN(n14691) );
  NAND2_X1 U7932 ( .A1(n7395), .A2(n7535), .ZN(n7394) );
  INV_X1 U7933 ( .A(n7396), .ZN(n7395) );
  NAND2_X1 U7934 ( .A1(n8120), .A2(n8121), .ZN(n8139) );
  INV_X1 U7935 ( .A(n8069), .ZN(n6909) );
  NAND2_X1 U7936 ( .A1(n6797), .A2(n8070), .ZN(n9274) );
  AND2_X1 U7937 ( .A1(n8089), .A2(n8085), .ZN(n6797) );
  INV_X1 U7938 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n7544) );
  NAND2_X1 U7939 ( .A1(n7951), .A2(n7950), .ZN(n7987) );
  INV_X1 U7940 ( .A(n7952), .ZN(n7950) );
  AND2_X1 U7941 ( .A1(n6914), .A2(n7946), .ZN(n7978) );
  NAND2_X1 U7942 ( .A1(n7366), .A2(n7849), .ZN(n7871) );
  NAND2_X1 U7943 ( .A1(n7767), .A2(n7766), .ZN(n7790) );
  INV_X1 U7944 ( .A(n6899), .ZN(n6898) );
  NAND2_X1 U7945 ( .A1(n7611), .A2(n7610), .ZN(n7616) );
  XNOR2_X1 U7946 ( .A(n6655), .B(n14272), .ZN(n14275) );
  INV_X1 U7947 ( .A(n14271), .ZN(n6655) );
  XNOR2_X1 U7948 ( .A(n14221), .B(n6990), .ZN(n14268) );
  INV_X1 U7949 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n6990) );
  NAND2_X1 U7950 ( .A1(n15397), .A2(n14282), .ZN(n14283) );
  AOI21_X1 U7951 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n14246), .A(n14245), .ZN(
        n14303) );
  AND2_X1 U7952 ( .A1(n13216), .A2(n12508), .ZN(n7315) );
  NAND2_X1 U7953 ( .A1(n9837), .A2(n12601), .ZN(n7052) );
  NAND2_X1 U7954 ( .A1(n8773), .A2(n8772), .ZN(n12966) );
  NAND2_X1 U7955 ( .A1(n9768), .A2(n9767), .ZN(n9769) );
  NAND2_X1 U7956 ( .A1(n9766), .A2(n9777), .ZN(n9768) );
  NAND2_X1 U7957 ( .A1(n8762), .A2(n8761), .ZN(n12865) );
  OR2_X1 U7958 ( .A1(n11004), .A2(n8760), .ZN(n8762) );
  AOI21_X1 U7959 ( .B1(n7046), .B2(n6534), .A(n7043), .ZN(n7042) );
  NAND2_X1 U7960 ( .A1(n6537), .A2(n7044), .ZN(n7043) );
  NAND2_X1 U7961 ( .A1(n8720), .A2(n8719), .ZN(n12930) );
  OR2_X1 U7962 ( .A1(n10429), .A2(n8760), .ZN(n8720) );
  INV_X1 U7963 ( .A(n12661), .ZN(n12912) );
  NAND2_X1 U7964 ( .A1(n8747), .A2(n8746), .ZN(n12877) );
  OR2_X1 U7965 ( .A1(n10880), .A2(n8760), .ZN(n8747) );
  AND2_X1 U7966 ( .A1(n9856), .A2(n15112), .ZN(n12649) );
  OAI21_X2 U7967 ( .B1(n9854), .B2(n9853), .A(n9852), .ZN(n12642) );
  INV_X1 U7968 ( .A(n12649), .ZN(n12634) );
  INV_X1 U7969 ( .A(n12642), .ZN(n12637) );
  AND3_X1 U7970 ( .A1(n10738), .A2(n12370), .A3(n8482), .ZN(n15103) );
  NAND2_X1 U7971 ( .A1(n8755), .A2(n8754), .ZN(n12887) );
  XNOR2_X1 U7972 ( .A(n8560), .B(P3_IR_REG_6__SCAN_IN), .ZN(n10858) );
  NAND2_X1 U7973 ( .A1(n7008), .A2(n7010), .ZN(n11788) );
  NAND2_X1 U7974 ( .A1(n7008), .A2(n7007), .ZN(n7009) );
  AND2_X1 U7975 ( .A1(n7010), .A2(n12680), .ZN(n7007) );
  NOR2_X1 U7976 ( .A1(n11789), .A2(n8674), .ZN(n12676) );
  NAND2_X1 U7977 ( .A1(n6844), .A2(n15069), .ZN(n6843) );
  XNOR2_X1 U7978 ( .A(n12758), .B(n6845), .ZN(n6844) );
  INV_X1 U7979 ( .A(n12757), .ZN(n6845) );
  INV_X1 U7980 ( .A(n7039), .ZN(n7036) );
  NAND2_X1 U7981 ( .A1(n7038), .A2(n7040), .ZN(n7037) );
  OR2_X1 U7982 ( .A1(n12745), .A2(n14390), .ZN(n7040) );
  INV_X1 U7983 ( .A(n12933), .ZN(n14402) );
  AND2_X1 U7984 ( .A1(n8847), .A2(n8846), .ZN(n9888) );
  OAI21_X1 U7985 ( .B1(n6975), .B2(n6836), .A(n6834), .ZN(n6832) );
  NAND2_X1 U7986 ( .A1(n6835), .A2(n12922), .ZN(n6834) );
  NAND2_X1 U7987 ( .A1(n15183), .A2(n15150), .ZN(n13003) );
  INV_X1 U7988 ( .A(n9848), .ZN(n13022) );
  NAND2_X1 U7989 ( .A1(n8457), .A2(n8456), .ZN(n13047) );
  NAND2_X1 U7990 ( .A1(n8422), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8418) );
  OAI21_X1 U7991 ( .B1(n8811), .B2(n8810), .A(n8812), .ZN(n8826) );
  CLKBUF_X1 U7992 ( .A(n8898), .Z(n8454) );
  NAND2_X1 U7993 ( .A1(n7305), .A2(n6575), .ZN(n14427) );
  INV_X1 U7994 ( .A(n14425), .ZN(n7304) );
  OR2_X1 U7995 ( .A1(n10484), .A2(n10483), .ZN(n10485) );
  OR2_X1 U7996 ( .A1(n10077), .A2(n9664), .ZN(n6868) );
  NAND2_X1 U7997 ( .A1(n6866), .A2(n6867), .ZN(n13174) );
  NAND2_X1 U7998 ( .A1(n6862), .A2(n6861), .ZN(n6866) );
  INV_X1 U7999 ( .A(n12501), .ZN(n6861) );
  INV_X1 U8000 ( .A(n12502), .ZN(n6862) );
  INV_X1 U8001 ( .A(n13401), .ZN(n13563) );
  NAND2_X1 U8002 ( .A1(n9321), .A2(n9320), .ZN(n13553) );
  NAND2_X1 U8003 ( .A1(n9204), .A2(n9203), .ZN(n13611) );
  NAND2_X1 U8004 ( .A1(n7442), .A2(n7433), .ZN(n13540) );
  NAND2_X1 U8005 ( .A1(n7436), .A2(n7434), .ZN(n7433) );
  NAND2_X1 U8006 ( .A1(n7440), .A2(n7445), .ZN(n7436) );
  OAI21_X1 U8007 ( .B1(n13539), .B2(n14903), .A(n9429), .ZN(n9434) );
  NAND2_X1 U8008 ( .A1(n7093), .A2(n7098), .ZN(n13539) );
  AND2_X1 U8009 ( .A1(n9344), .A2(n9343), .ZN(n13344) );
  OAI21_X1 U8010 ( .B1(n13336), .B2(n13337), .A(n13335), .ZN(n13541) );
  OR2_X1 U8011 ( .A1(n10065), .A2(n9664), .ZN(n9080) );
  AND2_X1 U8012 ( .A1(n14919), .A2(n9432), .ZN(n14916) );
  INV_X1 U8013 ( .A(n10216), .ZN(n9432) );
  NOR2_X1 U8014 ( .A1(n7264), .A2(n13817), .ZN(n7262) );
  NOR2_X1 U8015 ( .A1(n7267), .A2(n7265), .ZN(n7264) );
  INV_X1 U8016 ( .A(n7268), .ZN(n7265) );
  NAND2_X1 U8017 ( .A1(n7268), .A2(n7269), .ZN(n7266) );
  NAND2_X1 U8018 ( .A1(n8141), .A2(n8140), .ZN(n14125) );
  NAND2_X1 U8019 ( .A1(n14673), .A2(n10467), .ZN(n13815) );
  OAI21_X1 U8020 ( .B1(n7499), .B2(n11828), .A(n8337), .ZN(n6892) );
  NAND2_X1 U8021 ( .A1(n8205), .A2(n8204), .ZN(n13821) );
  NAND2_X1 U8022 ( .A1(n8187), .A2(n8186), .ZN(n13956) );
  XNOR2_X1 U8023 ( .A(n6871), .B(n14091), .ZN(n14089) );
  NOR2_X1 U8024 ( .A1(n13929), .A2(n14096), .ZN(n6870) );
  AND2_X1 U8025 ( .A1(n12486), .A2(n13935), .ZN(n14100) );
  NAND2_X1 U8026 ( .A1(n8211), .A2(n8210), .ZN(n14104) );
  NAND2_X1 U8027 ( .A1(n12041), .A2(n8282), .ZN(n8211) );
  NAND2_X1 U8028 ( .A1(n7749), .A2(n7748), .ZN(n11589) );
  XNOR2_X1 U8029 ( .A(n14275), .B(n10313), .ZN(n15409) );
  OAI21_X1 U8030 ( .B1(n14550), .B2(n14551), .A(n6996), .ZN(n6995) );
  INV_X1 U8031 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6996) );
  NAND2_X1 U8032 ( .A1(n14343), .A2(n6997), .ZN(n15380) );
  INV_X1 U8033 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n6998) );
  NOR2_X1 U8034 ( .A1(n9506), .A2(n9503), .ZN(n7418) );
  INV_X1 U8035 ( .A(n9503), .ZN(n7417) );
  NAND2_X1 U8036 ( .A1(n9529), .A2(n6511), .ZN(n7425) );
  INV_X1 U8037 ( .A(n7702), .ZN(n7175) );
  NOR2_X1 U8038 ( .A1(n7177), .A2(n7702), .ZN(n7176) );
  NAND2_X1 U8039 ( .A1(n9542), .A2(n6510), .ZN(n7430) );
  NAND2_X1 U8040 ( .A1(n7725), .A2(n7726), .ZN(n7724) );
  AOI21_X1 U8041 ( .B1(n7208), .B2(n7206), .A(n7205), .ZN(n7204) );
  NAND2_X1 U8042 ( .A1(n7802), .A2(n7201), .ZN(n7200) );
  NOR2_X1 U8043 ( .A1(n7201), .A2(n7802), .ZN(n7202) );
  INV_X1 U8044 ( .A(n9559), .ZN(n6675) );
  AND2_X1 U8045 ( .A1(n7196), .A2(n7194), .ZN(n7192) );
  AND2_X1 U8046 ( .A1(n8005), .A2(n7211), .ZN(n7210) );
  NAND2_X1 U8047 ( .A1(n7212), .A2(n7215), .ZN(n7211) );
  INV_X1 U8048 ( .A(n9623), .ZN(n6697) );
  INV_X1 U8049 ( .A(n9639), .ZN(n7423) );
  INV_X1 U8050 ( .A(n9635), .ZN(n6721) );
  INV_X1 U8051 ( .A(n9636), .ZN(n6722) );
  NAND2_X1 U8052 ( .A1(n7180), .A2(n7179), .ZN(n8101) );
  NAND2_X1 U8053 ( .A1(n8074), .A2(n8075), .ZN(n7179) );
  NOR2_X1 U8054 ( .A1(n9644), .A2(n9643), .ZN(n9645) );
  NAND2_X1 U8055 ( .A1(n7186), .A2(n7185), .ZN(n8144) );
  NAND2_X1 U8056 ( .A1(n8126), .A2(n8128), .ZN(n7185) );
  NOR2_X1 U8057 ( .A1(n7893), .A2(n7892), .ZN(n7897) );
  NAND2_X1 U8058 ( .A1(n7189), .A2(n7188), .ZN(n8190) );
  NAND2_X1 U8059 ( .A1(n8167), .A2(n8169), .ZN(n7188) );
  NAND2_X1 U8060 ( .A1(n7366), .A2(n7364), .ZN(n7896) );
  NOR2_X1 U8061 ( .A1(n6558), .A2(n7365), .ZN(n7364) );
  INV_X1 U8062 ( .A(n7849), .ZN(n7365) );
  MUX2_X1 U8063 ( .A(n12204), .B(n12203), .S(n12370), .Z(n12360) );
  NAND2_X1 U8064 ( .A1(n7027), .A2(n10824), .ZN(n7026) );
  INV_X1 U8065 ( .A(n7028), .ZN(n7027) );
  NAND2_X1 U8066 ( .A1(n15023), .A2(n7028), .ZN(n7025) );
  AND2_X1 U8067 ( .A1(n15005), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7028) );
  AND2_X1 U8068 ( .A1(n9848), .A2(n12811), .ZN(n12166) );
  NAND2_X1 U8069 ( .A1(n11762), .A2(n14407), .ZN(n6752) );
  INV_X1 U8070 ( .A(n8521), .ZN(n6971) );
  INV_X1 U8071 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n6953) );
  INV_X1 U8072 ( .A(n9656), .ZN(n6688) );
  INV_X1 U8073 ( .A(n9356), .ZN(n7103) );
  AND2_X1 U8074 ( .A1(n13505), .A2(n6947), .ZN(n6946) );
  AND2_X1 U8075 ( .A1(n9430), .A2(n6948), .ZN(n6947) );
  NAND2_X1 U8076 ( .A1(n6902), .A2(n6901), .ZN(n8214) );
  NAND2_X1 U8077 ( .A1(n13821), .A2(n8212), .ZN(n6901) );
  NAND2_X1 U8078 ( .A1(n14104), .A2(n8256), .ZN(n6902) );
  NAND2_X1 U8079 ( .A1(n8120), .A2(n6930), .ZN(n6929) );
  NOR2_X1 U8080 ( .A1(n6928), .A2(n6931), .ZN(n6930) );
  INV_X1 U8081 ( .A(n6925), .ZN(n6924) );
  OAI21_X1 U8082 ( .B1(n8138), .B2(n6928), .A(n6926), .ZN(n6925) );
  INV_X1 U8083 ( .A(n6927), .ZN(n6926) );
  OAI21_X1 U8084 ( .B1(n6933), .B2(n6928), .A(n15310), .ZN(n6927) );
  INV_X1 U8085 ( .A(n8150), .ZN(n6933) );
  INV_X1 U8086 ( .A(n7837), .ZN(n6918) );
  OAI21_X1 U8087 ( .B1(n7631), .B2(SI_2_), .A(n6726), .ZN(n6852) );
  OAI21_X1 U8088 ( .B1(n7612), .B2(n10039), .A(n6728), .ZN(n7613) );
  NAND2_X1 U8089 ( .A1(n7612), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6728) );
  INV_X1 U8090 ( .A(n11515), .ZN(n7077) );
  NAND2_X1 U8091 ( .A1(n6541), .A2(n7297), .ZN(n7296) );
  NOR2_X1 U8092 ( .A1(n12132), .A2(n12131), .ZN(n7298) );
  NAND2_X1 U8093 ( .A1(n6739), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8490) );
  OR2_X1 U8094 ( .A1(n14972), .A2(n6778), .ZN(n7018) );
  NAND2_X1 U8095 ( .A1(n6779), .A2(n7019), .ZN(n6778) );
  INV_X1 U8096 ( .A(n10821), .ZN(n6779) );
  INV_X1 U8097 ( .A(n7026), .ZN(n7019) );
  OAI21_X1 U8098 ( .B1(n14999), .B2(n7024), .A(n7021), .ZN(n7020) );
  NAND2_X1 U8099 ( .A1(n15023), .A2(n7023), .ZN(n7024) );
  INV_X1 U8100 ( .A(n7022), .ZN(n7021) );
  OAI21_X1 U8101 ( .B1(n7026), .B2(n7023), .A(n7025), .ZN(n7022) );
  AOI21_X1 U8102 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n10866), .A(n10865), .ZN(
        n10868) );
  AND2_X1 U8103 ( .A1(n6771), .A2(n6773), .ZN(n12730) );
  NOR2_X1 U8104 ( .A1(n7012), .A2(n14349), .ZN(n6771) );
  INV_X1 U8105 ( .A(n12350), .ZN(n7291) );
  OR2_X1 U8106 ( .A1(n9848), .A2(n12811), .ZN(n12354) );
  INV_X1 U8107 ( .A(n12652), .ZN(n12811) );
  NOR2_X1 U8108 ( .A1(n12334), .A2(n6814), .ZN(n6813) );
  INV_X1 U8109 ( .A(n6821), .ZN(n6814) );
  NAND2_X1 U8110 ( .A1(n6817), .A2(n12333), .ZN(n6816) );
  INV_X1 U8111 ( .A(n6818), .ZN(n6817) );
  AND2_X1 U8112 ( .A1(n8749), .A2(n8748), .ZN(n8764) );
  INV_X1 U8113 ( .A(n12311), .ZN(n6826) );
  INV_X1 U8114 ( .A(n12320), .ZN(n6825) );
  NOR2_X1 U8115 ( .A1(n12913), .A2(n6765), .ZN(n6764) );
  AOI21_X1 U8116 ( .B1(n6499), .B2(n6763), .A(n6762), .ZN(n6761) );
  NOR2_X1 U8117 ( .A1(n13055), .A2(n12924), .ZN(n6762) );
  AND2_X1 U8118 ( .A1(n8721), .A2(n15330), .ZN(n8735) );
  INV_X1 U8119 ( .A(n6961), .ZN(n6960) );
  NOR2_X1 U8120 ( .A1(n6961), .A2(n8563), .ZN(n6959) );
  OR2_X1 U8121 ( .A1(n12671), .A2(n15144), .ZN(n12244) );
  INV_X1 U8122 ( .A(n12651), .ZN(n8840) );
  NAND2_X1 U8123 ( .A1(n12368), .A2(n12369), .ZN(n12198) );
  NAND2_X1 U8124 ( .A1(n8347), .A2(n7302), .ZN(n7301) );
  INV_X1 U8125 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n7302) );
  INV_X1 U8126 ( .A(n8812), .ZN(n7169) );
  NOR2_X1 U8127 ( .A1(n8349), .A2(n8612), .ZN(n6734) );
  INV_X1 U8128 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8905) );
  NOR2_X1 U8129 ( .A1(P3_IR_REG_23__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), .ZN(
        n7078) );
  AOI21_X1 U8130 ( .B1(n8443), .B2(n7152), .A(n7151), .ZN(n7150) );
  INV_X1 U8131 ( .A(n8402), .ZN(n7151) );
  NAND2_X1 U8132 ( .A1(n8403), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8405) );
  INV_X1 U8133 ( .A(n8373), .ZN(n7161) );
  OR2_X1 U8134 ( .A1(n8592), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8593) );
  NAND2_X1 U8135 ( .A1(n10062), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8371) );
  NAND4_X1 U8136 ( .A1(n8503), .A2(n8517), .A3(n7294), .A4(n7293), .ZN(n8531)
         );
  INV_X1 U8137 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n7293) );
  INV_X1 U8138 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7294) );
  NOR2_X1 U8139 ( .A1(n9122), .A2(n9121), .ZN(n9120) );
  NOR2_X1 U8140 ( .A1(n9223), .A2(n8997), .ZN(n8959) );
  INV_X1 U8141 ( .A(n7125), .ZN(n7121) );
  NAND2_X1 U8142 ( .A1(n7474), .A2(n13196), .ZN(n7473) );
  INV_X1 U8143 ( .A(n7471), .ZN(n7470) );
  NOR2_X1 U8144 ( .A1(n9278), .A2(n9277), .ZN(n9301) );
  INV_X1 U8145 ( .A(n13424), .ZN(n6708) );
  NAND2_X1 U8146 ( .A1(n13586), .A2(n9259), .ZN(n7138) );
  AND2_X1 U8147 ( .A1(n11702), .A2(n6944), .ZN(n13469) );
  AND2_X1 U8148 ( .A1(n6946), .A2(n6945), .ZN(n6944) );
  NAND2_X1 U8149 ( .A1(n9128), .A2(n7085), .ZN(n7091) );
  INV_X1 U8150 ( .A(n9116), .ZN(n7085) );
  OR2_X1 U8151 ( .A1(n9109), .A2(n9108), .ZN(n9122) );
  AND2_X1 U8152 ( .A1(n9469), .A2(n10208), .ZN(n9672) );
  INV_X1 U8153 ( .A(n7453), .ZN(n7449) );
  NOR2_X1 U8154 ( .A1(n13470), .A2(n13586), .ZN(n13458) );
  NAND2_X1 U8155 ( .A1(n11702), .A2(n6946), .ZN(n13507) );
  OAI21_X1 U8156 ( .B1(n7106), .B2(n7105), .A(n6509), .ZN(n6712) );
  INV_X1 U8157 ( .A(n11267), .ZN(n6713) );
  NAND2_X1 U8158 ( .A1(n6941), .A2(n6940), .ZN(n14896) );
  INV_X1 U8159 ( .A(n14895), .ZN(n6941) );
  NAND2_X1 U8160 ( .A1(n11160), .A2(n14930), .ZN(n14895) );
  NOR2_X1 U8161 ( .A1(n7829), .A2(n7828), .ZN(n7861) );
  OR2_X1 U8162 ( .A1(n7184), .A2(n8214), .ZN(n7182) );
  NOR2_X1 U8163 ( .A1(n14133), .A2(n14125), .ZN(n6875) );
  INV_X1 U8164 ( .A(n9925), .ZN(n7369) );
  OR2_X1 U8165 ( .A1(n14503), .A2(n13714), .ZN(n9917) );
  NOR2_X1 U8166 ( .A1(n7908), .A2(n13806), .ZN(n7925) );
  INV_X1 U8167 ( .A(n9915), .ZN(n7352) );
  NOR2_X1 U8168 ( .A1(n7352), .A2(n7349), .ZN(n7348) );
  INV_X1 U8169 ( .A(n9914), .ZN(n7349) );
  NOR2_X1 U8170 ( .A1(n7756), .A2(n10176), .ZN(n7780) );
  INV_X1 U8171 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7705) );
  AND2_X1 U8172 ( .A1(n9963), .A2(n9903), .ZN(n7358) );
  INV_X1 U8173 ( .A(n8299), .ZN(n9893) );
  NOR2_X1 U8174 ( .A1(n6884), .A2(n14503), .ZN(n6883) );
  INV_X1 U8175 ( .A(n6885), .ZN(n6884) );
  NAND2_X1 U8176 ( .A1(n7386), .A2(n8274), .ZN(n7385) );
  INV_X1 U8177 ( .A(n8233), .ZN(n7384) );
  INV_X1 U8178 ( .A(n8278), .ZN(n7382) );
  NAND2_X1 U8179 ( .A1(n6905), .A2(n6632), .ZN(n6903) );
  NAND2_X1 U8180 ( .A1(n6904), .A2(n7375), .ZN(n6719) );
  NAND2_X1 U8181 ( .A1(n7987), .A2(n7986), .ZN(n8023) );
  INV_X1 U8182 ( .A(n7947), .ZN(n7934) );
  INV_X1 U8183 ( .A(n6494), .ZN(n6796) );
  XNOR2_X1 U8184 ( .A(n7848), .B(SI_12_), .ZN(n7846) );
  NAND2_X1 U8185 ( .A1(n7684), .A2(n6787), .ZN(n6786) );
  NAND2_X1 U8186 ( .A1(n6787), .A2(n6785), .ZN(n6784) );
  NAND2_X1 U8187 ( .A1(n6798), .A2(SI_4_), .ZN(n7663) );
  NAND2_X1 U8188 ( .A1(n6652), .A2(n7631), .ZN(n7611) );
  NAND2_X1 U8189 ( .A1(n14226), .A2(n14227), .ZN(n14228) );
  AOI22_X1 U8190 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14233), .B1(n14284), .B2(
        n14232), .ZN(n14234) );
  INV_X1 U8191 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14233) );
  INV_X1 U8192 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n15330) );
  OR2_X1 U8193 ( .A1(n8737), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8468) );
  NOR2_X1 U8194 ( .A1(n8468), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8749) );
  NAND2_X1 U8195 ( .A1(n7070), .A2(n6571), .ZN(n12569) );
  NAND2_X1 U8196 ( .A1(n9807), .A2(n9804), .ZN(n7044) );
  NOR2_X1 U8197 ( .A1(n7490), .A2(n7047), .ZN(n7046) );
  INV_X1 U8198 ( .A(n12112), .ZN(n7047) );
  AND2_X1 U8199 ( .A1(n12580), .A2(n9841), .ZN(n12602) );
  OR2_X1 U8200 ( .A1(n8473), .A2(n8355), .ZN(n8476) );
  NAND2_X1 U8201 ( .A1(n6739), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8477) );
  OR2_X1 U8202 ( .A1(n8688), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8705) );
  NOR2_X1 U8203 ( .A1(n8705), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8721) );
  OAI22_X1 U8204 ( .A1(n8778), .A2(n10765), .B1(n10766), .B2(n12148), .ZN(
        n6802) );
  NAND2_X1 U8205 ( .A1(n8480), .A2(n6529), .ZN(n7032) );
  OAI22_X1 U8206 ( .A1(n7030), .A2(n7029), .B1(n7031), .B2(n10757), .ZN(n10760) );
  INV_X1 U8207 ( .A(n8480), .ZN(n7030) );
  NAND2_X1 U8208 ( .A1(n6529), .A2(n10740), .ZN(n7029) );
  OR2_X1 U8209 ( .A1(n10834), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n6777) );
  NAND2_X1 U8210 ( .A1(n10844), .A2(n15015), .ZN(n10847) );
  NOR2_X1 U8211 ( .A1(n11373), .A2(n6634), .ZN(n11374) );
  OR2_X1 U8212 ( .A1(n15046), .A2(n15047), .ZN(n7002) );
  XNOR2_X1 U8213 ( .A(n11378), .B(n6837), .ZN(n15059) );
  NAND2_X1 U8214 ( .A1(n11377), .A2(n6838), .ZN(n11378) );
  NAND2_X1 U8215 ( .A1(n6839), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n6838) );
  OAI21_X1 U8216 ( .B1(n15075), .B2(n15074), .A(n15073), .ZN(n15077) );
  AND2_X1 U8217 ( .A1(n15072), .A2(n11375), .ZN(n11549) );
  INV_X1 U8218 ( .A(n11556), .ZN(n11565) );
  NAND2_X1 U8219 ( .A1(n11557), .A2(n11558), .ZN(n11561) );
  NAND2_X1 U8220 ( .A1(n11561), .A2(n11560), .ZN(n11790) );
  INV_X1 U8221 ( .A(n7005), .ZN(n7003) );
  AOI21_X1 U8222 ( .B1(n11553), .B2(n6516), .A(n7006), .ZN(n7005) );
  NOR2_X1 U8223 ( .A1(n11787), .A2(n12688), .ZN(n7006) );
  NAND2_X1 U8224 ( .A1(n11790), .A2(n6840), .ZN(n12679) );
  NAND2_X1 U8225 ( .A1(n11793), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n6840) );
  NAND2_X1 U8226 ( .A1(n6770), .A2(n12715), .ZN(n12724) );
  NOR2_X1 U8227 ( .A1(n12739), .A2(n14351), .ZN(n14370) );
  XNOR2_X1 U8228 ( .A(n12730), .B(n14365), .ZN(n14374) );
  NOR2_X1 U8229 ( .A1(n14374), .A2(n8738), .ZN(n14375) );
  NAND2_X1 U8230 ( .A1(n14366), .A2(n12756), .ZN(n14386) );
  INV_X1 U8231 ( .A(n12753), .ZN(n12754) );
  AOI21_X1 U8232 ( .B1(n7039), .B2(n14390), .A(n6645), .ZN(n7038) );
  OAI21_X1 U8233 ( .B1(n12786), .B2(n12785), .A(n12199), .ZN(n12769) );
  OAI21_X1 U8234 ( .B1(n12822), .B2(n6831), .A(n7290), .ZN(n12801) );
  AOI21_X1 U8235 ( .B1(n12813), .B2(n7292), .A(n7291), .ZN(n7290) );
  NAND2_X1 U8236 ( .A1(n12813), .A2(n8891), .ZN(n6831) );
  INV_X1 U8237 ( .A(n12346), .ZN(n7292) );
  AND2_X1 U8238 ( .A1(n12353), .A2(n12354), .ZN(n12800) );
  NAND2_X1 U8239 ( .A1(n12825), .A2(n8794), .ZN(n12812) );
  NOR2_X1 U8240 ( .A1(n12813), .A2(n6967), .ZN(n6966) );
  INV_X1 U8241 ( .A(n8794), .ZN(n6967) );
  AOI21_X1 U8242 ( .B1(n12841), .B2(n12336), .A(n6740), .ZN(n12827) );
  AND2_X1 U8243 ( .A1(n12966), .A2(n12655), .ZN(n6740) );
  AOI21_X1 U8244 ( .B1(n12817), .B2(n8793), .A(n8358), .ZN(n12829) );
  NAND2_X1 U8245 ( .A1(n8764), .A2(n8763), .ZN(n8766) );
  AND2_X1 U8246 ( .A1(n6756), .A2(n6977), .ZN(n6755) );
  AOI21_X1 U8247 ( .B1(n6497), .B2(n12897), .A(n6592), .ZN(n6977) );
  NAND2_X1 U8248 ( .A1(n7286), .A2(n7288), .ZN(n12901) );
  AOI21_X1 U8249 ( .B1(n12913), .B2(n7289), .A(n12315), .ZN(n7288) );
  INV_X1 U8250 ( .A(n12304), .ZN(n7289) );
  AOI21_X1 U8251 ( .B1(n6522), .B2(n6811), .A(n6809), .ZN(n6808) );
  INV_X1 U8252 ( .A(n12296), .ZN(n6809) );
  AND2_X1 U8253 ( .A1(n12291), .A2(n12303), .ZN(n12290) );
  AOI21_X1 U8254 ( .B1(n6496), .B2(n6747), .A(n6635), .ZN(n6744) );
  AND2_X1 U8255 ( .A1(n6751), .A2(n6551), .ZN(n11778) );
  NAND2_X1 U8256 ( .A1(n11760), .A2(n12182), .ZN(n6751) );
  OR2_X1 U8257 ( .A1(n8643), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8659) );
  AOI21_X1 U8258 ( .B1(n7278), .B2(n7280), .A(n7277), .ZN(n7276) );
  AND2_X1 U8259 ( .A1(n12273), .A2(n12265), .ZN(n12272) );
  OR2_X1 U8260 ( .A1(n8618), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8643) );
  NOR2_X1 U8261 ( .A1(n8565), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8582) );
  INV_X1 U8262 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n15301) );
  AND2_X1 U8263 ( .A1(n8582), .A2(n15301), .ZN(n8602) );
  INV_X1 U8264 ( .A(n11409), .ZN(n12246) );
  NAND2_X1 U8265 ( .A1(n11184), .A2(n8563), .ZN(n11410) );
  OR2_X1 U8266 ( .A1(n8552), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8565) );
  NAND2_X1 U8267 ( .A1(n6520), .A2(n11185), .ZN(n11184) );
  INV_X1 U8268 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n15288) );
  NAND2_X1 U8269 ( .A1(n11037), .A2(n12228), .ZN(n11036) );
  INV_X1 U8270 ( .A(n11034), .ZN(n12228) );
  NAND2_X1 U8271 ( .A1(n12234), .A2(n12236), .ZN(n11034) );
  NAND2_X1 U8272 ( .A1(n11193), .A2(n8521), .ZN(n11035) );
  NAND2_X1 U8273 ( .A1(n12226), .A2(n12229), .ZN(n11194) );
  AND2_X1 U8274 ( .A1(n15092), .A2(n8508), .ZN(n11195) );
  NAND2_X1 U8275 ( .A1(n11195), .A2(n11194), .ZN(n11193) );
  NAND2_X1 U8276 ( .A1(n6799), .A2(n8505), .ZN(n15088) );
  NAND2_X1 U8277 ( .A1(n9766), .A2(n8874), .ZN(n15087) );
  INV_X1 U8278 ( .A(n15093), .ZN(n12179) );
  AND2_X1 U8279 ( .A1(n8901), .A2(n10891), .ZN(n15110) );
  NAND2_X1 U8280 ( .A1(n12808), .A2(n12813), .ZN(n12810) );
  NAND2_X1 U8281 ( .A1(n12824), .A2(n12346), .ZN(n12808) );
  OR2_X1 U8282 ( .A1(n12901), .A2(n12900), .ZN(n12991) );
  OR2_X1 U8283 ( .A1(n15111), .A2(n12384), .ZN(n15169) );
  NAND2_X1 U8284 ( .A1(n11030), .A2(n12211), .ZN(n15168) );
  INV_X1 U8285 ( .A(n15169), .ZN(n15164) );
  INV_X1 U8286 ( .A(n8873), .ZN(n10681) );
  NAND2_X1 U8287 ( .A1(n8918), .A2(n8917), .ZN(n10893) );
  AND2_X1 U8288 ( .A1(n7299), .A2(n6828), .ZN(n6827) );
  INV_X1 U8289 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n6828) );
  NAND2_X1 U8290 ( .A1(n8796), .A2(n8795), .ZN(n8798) );
  NAND2_X1 U8291 ( .A1(n8745), .A2(n8405), .ZN(n8757) );
  NAND2_X1 U8292 ( .A1(n8757), .A2(n8756), .ZN(n8759) );
  NAND2_X1 U8293 ( .A1(n8405), .A2(n8404), .ZN(n8743) );
  OR2_X1 U8294 ( .A1(n8403), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8404) );
  NAND2_X1 U8295 ( .A1(n8714), .A2(n8396), .ZN(n8728) );
  AND2_X1 U8296 ( .A1(n8398), .A2(n8397), .ZN(n8727) );
  AOI21_X1 U8297 ( .B1(n6625), .B2(n8391), .A(n7171), .ZN(n7170) );
  INV_X1 U8298 ( .A(n8394), .ZN(n7171) );
  AND2_X1 U8299 ( .A1(n8396), .A2(n8395), .ZN(n8711) );
  NAND2_X1 U8300 ( .A1(n8712), .A2(n8711), .ZN(n8714) );
  INV_X1 U8301 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8700) );
  INV_X1 U8302 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8684) );
  INV_X1 U8303 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8449) );
  INV_X1 U8304 ( .A(n8654), .ZN(n8450) );
  AOI21_X1 U8305 ( .B1(n7156), .B2(n7158), .A(n6637), .ZN(n7154) );
  NOR2_X1 U8306 ( .A1(n8593), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n8629) );
  NAND2_X1 U8307 ( .A1(n8591), .A2(n8378), .ZN(n8609) );
  AND2_X1 U8308 ( .A1(n8380), .A2(n8379), .ZN(n8608) );
  NAND2_X1 U8309 ( .A1(n8609), .A2(n8608), .ZN(n8611) );
  OAI21_X1 U8310 ( .B1(n8559), .B2(n7162), .A(n7159), .ZN(n8589) );
  AOI21_X1 U8311 ( .B1(n7163), .B2(n7161), .A(n7160), .ZN(n7159) );
  INV_X1 U8312 ( .A(n7163), .ZN(n7162) );
  INV_X1 U8313 ( .A(n8376), .ZN(n7160) );
  AND2_X1 U8314 ( .A1(n8378), .A2(n8377), .ZN(n8588) );
  NAND2_X1 U8315 ( .A1(n8589), .A2(n8588), .ZN(n8591) );
  NAND2_X1 U8316 ( .A1(n7143), .A2(n7141), .ZN(n8545) );
  AOI21_X1 U8317 ( .B1(n7145), .B2(n7146), .A(n7142), .ZN(n7141) );
  INV_X1 U8318 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8546) );
  NOR2_X2 U8319 ( .A1(n8531), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n8530) );
  NAND2_X1 U8320 ( .A1(n8361), .A2(n8360), .ZN(n8502) );
  INV_X1 U8321 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8503) );
  AND2_X1 U8322 ( .A1(n10708), .A2(n10615), .ZN(n10620) );
  NOR2_X1 U8323 ( .A1(n11730), .A2(n7307), .ZN(n7306) );
  INV_X1 U8324 ( .A(n11364), .ZN(n7307) );
  OR2_X1 U8325 ( .A1(n11728), .A2(n11727), .ZN(n11729) );
  AND2_X1 U8326 ( .A1(n13107), .A2(n13104), .ZN(n7324) );
  AND2_X1 U8327 ( .A1(n13099), .A2(n13096), .ZN(n13160) );
  NOR2_X1 U8328 ( .A1(n12500), .A2(n12501), .ZN(n6860) );
  CLKBUF_X1 U8329 ( .A(n10601), .Z(n10490) );
  CLKBUF_X1 U8330 ( .A(n10619), .Z(n10700) );
  AND2_X1 U8331 ( .A1(n13228), .A2(n13099), .ZN(n13100) );
  OR2_X1 U8332 ( .A1(n10219), .A2(n10107), .ZN(n14420) );
  CLKBUF_X1 U8333 ( .A(n8996), .Z(n9667) );
  OR2_X1 U8334 ( .A1(n14810), .A2(n14809), .ZN(n14812) );
  OR2_X1 U8335 ( .A1(n10422), .A2(n10421), .ZN(n10797) );
  OR2_X1 U8336 ( .A1(n14829), .A2(n14830), .ZN(n14827) );
  NAND2_X1 U8337 ( .A1(n13635), .A2(n9679), .ZN(n9681) );
  INV_X1 U8338 ( .A(n7438), .ZN(n7435) );
  NAND2_X1 U8339 ( .A1(n7447), .A2(n7446), .ZN(n7445) );
  NAND2_X1 U8340 ( .A1(n7100), .A2(n7094), .ZN(n7093) );
  AND2_X1 U8341 ( .A1(n7101), .A2(n7097), .ZN(n7094) );
  NAND2_X1 U8342 ( .A1(n7104), .A2(n7099), .ZN(n7098) );
  AND2_X1 U8343 ( .A1(n9346), .A2(n9336), .ZN(n13350) );
  NOR2_X1 U8344 ( .A1(n13365), .A2(n13547), .ZN(n13349) );
  NOR2_X1 U8345 ( .A1(n13397), .A2(n13558), .ZN(n13384) );
  NAND2_X1 U8346 ( .A1(n13384), .A2(n13371), .ZN(n13365) );
  NOR2_X1 U8347 ( .A1(n13429), .A2(n13569), .ZN(n13415) );
  AOI21_X1 U8348 ( .B1(n7462), .B2(n7460), .A(n6583), .ZN(n7459) );
  INV_X1 U8349 ( .A(n9463), .ZN(n7460) );
  NOR2_X1 U8350 ( .A1(n13434), .A2(n13433), .ZN(n13436) );
  NAND2_X1 U8351 ( .A1(n6951), .A2(n6950), .ZN(n13429) );
  INV_X1 U8352 ( .A(n6791), .ZN(n13423) );
  NAND2_X1 U8353 ( .A1(n13469), .A2(n9431), .ZN(n13470) );
  AOI22_X1 U8354 ( .A1(n13512), .A2(n9228), .B1(n13607), .B2(n13185), .ZN(
        n13496) );
  NAND2_X1 U8355 ( .A1(n11702), .A2(n9430), .ZN(n13522) );
  NAND2_X1 U8356 ( .A1(n9168), .A2(n8957), .ZN(n9206) );
  NAND2_X1 U8357 ( .A1(n7111), .A2(n7112), .ZN(n11467) );
  NAND2_X1 U8358 ( .A1(n11267), .A2(n7114), .ZN(n7111) );
  OAI21_X1 U8359 ( .B1(n11316), .B2(n9454), .A(n6576), .ZN(n11471) );
  AOI21_X1 U8360 ( .B1(n7087), .B2(n7458), .A(n6565), .ZN(n7457) );
  INV_X1 U8361 ( .A(n9450), .ZN(n7458) );
  NAND2_X1 U8362 ( .A1(n11209), .A2(n6498), .ZN(n11272) );
  NAND2_X1 U8363 ( .A1(n11209), .A2(n11249), .ZN(n11208) );
  AND2_X1 U8364 ( .A1(n11217), .A2(n10999), .ZN(n11209) );
  OR2_X1 U8365 ( .A1(n9096), .A2(n9095), .ZN(n9109) );
  NAND2_X1 U8366 ( .A1(n14894), .A2(n9443), .ZN(n11215) );
  NOR2_X1 U8367 ( .A1(n10529), .A2(n10530), .ZN(n11160) );
  NAND2_X1 U8368 ( .A1(n10980), .A2(n10360), .ZN(n10506) );
  INV_X1 U8369 ( .A(n6653), .ZN(n10980) );
  AND2_X1 U8370 ( .A1(n10944), .A2(n10214), .ZN(n10360) );
  NOR2_X1 U8371 ( .A1(n9469), .A2(n11773), .ZN(n10373) );
  AND2_X1 U8372 ( .A1(n9404), .A2(n9400), .ZN(n14920) );
  INV_X1 U8373 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8983) );
  INV_X1 U8374 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8976) );
  NOR2_X1 U8375 ( .A1(n8974), .A2(n13637), .ZN(n6729) );
  INV_X1 U8376 ( .A(n8985), .ZN(n6737) );
  OR2_X1 U8377 ( .A1(n9396), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n9392) );
  OR2_X1 U8378 ( .A1(n9405), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n9394) );
  INV_X1 U8379 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8962) );
  INV_X1 U8380 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8964) );
  NAND2_X1 U8381 ( .A1(n7320), .A2(n7319), .ZN(n7318) );
  AND2_X1 U8382 ( .A1(n7319), .A2(n8989), .ZN(n8990) );
  AND2_X1 U8383 ( .A1(n9106), .A2(n9130), .ZN(n10415) );
  AND2_X1 U8384 ( .A1(n9065), .A2(n9090), .ZN(n10347) );
  NAND2_X1 U8385 ( .A1(n8076), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8107) );
  INV_X1 U8386 ( .A(n13668), .ZN(n7234) );
  OR2_X1 U8387 ( .A1(n7706), .A2(n7705), .ZN(n7732) );
  INV_X1 U8388 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7731) );
  INV_X1 U8389 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7828) );
  OR2_X1 U8390 ( .A1(n7732), .A2(n7731), .ZN(n7756) );
  NAND2_X1 U8391 ( .A1(n13687), .A2(n12099), .ZN(n12100) );
  NAND2_X1 U8392 ( .A1(n12100), .A2(n12101), .ZN(n13667) );
  INV_X1 U8393 ( .A(n10580), .ZN(n7238) );
  NAND2_X1 U8394 ( .A1(n10639), .A2(n7240), .ZN(n7241) );
  INV_X1 U8395 ( .A(n10642), .ZN(n7240) );
  INV_X2 U8396 ( .A(n12452), .ZN(n12446) );
  INV_X1 U8397 ( .A(n8260), .ZN(n8255) );
  AND4_X1 U8398 ( .A1(n7629), .A2(n7628), .A3(n7627), .A4(n7626), .ZN(n13728)
         );
  INV_X1 U8399 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10176) );
  INV_X1 U8400 ( .A(n14104), .ZN(n12478) );
  AND2_X1 U8401 ( .A1(n13992), .A2(n6599), .ZN(n13944) );
  NAND2_X1 U8402 ( .A1(n13992), .A2(n6873), .ZN(n13965) );
  NAND2_X1 U8403 ( .A1(n13992), .A2(n13981), .ZN(n13976) );
  AOI21_X1 U8404 ( .B1(n9998), .B2(n7355), .A(n6582), .ZN(n7353) );
  NOR2_X1 U8405 ( .A1(n14151), .A2(n14041), .ZN(n14027) );
  NOR2_X1 U8406 ( .A1(n14033), .A2(n7343), .ZN(n7342) );
  INV_X1 U8407 ( .A(n9923), .ZN(n7343) );
  AND2_X1 U8408 ( .A1(n8045), .A2(n8012), .ZN(n14036) );
  NAND2_X1 U8409 ( .A1(n7981), .A2(n7980), .ZN(n13734) );
  OR2_X1 U8410 ( .A1(n11976), .A2(n13734), .ZN(n14070) );
  NAND2_X1 U8411 ( .A1(n11945), .A2(n9918), .ZN(n11969) );
  AOI21_X1 U8412 ( .B1(n7389), .B2(n14475), .A(n6581), .ZN(n7387) );
  OR2_X1 U8413 ( .A1(n7878), .A2(n7862), .ZN(n7908) );
  NAND2_X1 U8414 ( .A1(n11692), .A2(n6887), .ZN(n14481) );
  AOI21_X1 U8415 ( .B1(n9979), .B2(n7328), .A(n6578), .ZN(n7327) );
  NAND2_X1 U8416 ( .A1(n11692), .A2(n14337), .ZN(n11809) );
  AOI21_X1 U8417 ( .B1(n9910), .B2(n7379), .A(n7378), .ZN(n7377) );
  INV_X1 U8418 ( .A(n9910), .ZN(n7380) );
  AND2_X1 U8419 ( .A1(n11652), .A2(n14526), .ZN(n11692) );
  NAND2_X1 U8420 ( .A1(n7780), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7807) );
  NAND2_X1 U8421 ( .A1(n14617), .A2(n9910), .ZN(n14619) );
  NOR2_X1 U8422 ( .A1(n6878), .A2(n6881), .ZN(n6877) );
  NAND2_X1 U8423 ( .A1(n10005), .A2(n6879), .ZN(n6878) );
  AOI21_X1 U8424 ( .B1(n11107), .B2(n7336), .A(n6579), .ZN(n7335) );
  NOR2_X1 U8425 ( .A1(n14660), .A2(n14724), .ZN(n11179) );
  NAND2_X1 U8426 ( .A1(n7362), .A2(n9902), .ZN(n11173) );
  AND2_X1 U8427 ( .A1(n14681), .A2(n14711), .ZN(n14678) );
  NAND2_X1 U8428 ( .A1(n6660), .A2(n6659), .ZN(n6658) );
  INV_X1 U8429 ( .A(n11005), .ZN(n6659) );
  NAND2_X1 U8430 ( .A1(n11010), .A2(n14694), .ZN(n8299) );
  NAND2_X1 U8431 ( .A1(n9992), .A2(n9991), .ZN(n14040) );
  OAI211_X1 U8432 ( .C1(n11987), .C2(n9939), .A(n14210), .B(n9938), .ZN(n10461) );
  AND2_X1 U8433 ( .A1(n10472), .A2(n10469), .ZN(n11232) );
  INV_X1 U8434 ( .A(n7218), .ZN(n8321) );
  INV_X1 U8435 ( .A(n11881), .ZN(n9950) );
  XNOR2_X1 U8436 ( .A(n8234), .B(n8233), .ZN(n12043) );
  XNOR2_X1 U8437 ( .A(n8222), .B(n8221), .ZN(n12041) );
  INV_X1 U8438 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7514) );
  INV_X1 U8439 ( .A(n7398), .ZN(n7397) );
  XNOR2_X1 U8440 ( .A(n8209), .B(n8176), .ZN(n13648) );
  XNOR2_X1 U8441 ( .A(n8172), .B(n8155), .ZN(n13651) );
  NAND2_X1 U8442 ( .A1(n6913), .A2(n6912), .ZN(n7948) );
  AOI22_X1 U8443 ( .A1(n6542), .A2(n6915), .B1(n6500), .B2(n7488), .ZN(n6912)
         );
  INV_X1 U8444 ( .A(n7503), .ZN(n7219) );
  NOR2_X1 U8445 ( .A1(n6526), .A2(n7588), .ZN(n7220) );
  NAND2_X1 U8446 ( .A1(n6919), .A2(n6921), .ZN(n7838) );
  NAND2_X1 U8447 ( .A1(n6920), .A2(n7793), .ZN(n6919) );
  OR2_X1 U8448 ( .A1(n7661), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n7719) );
  AND2_X1 U8449 ( .A1(n7664), .A2(n7638), .ZN(n10019) );
  OAI21_X1 U8450 ( .B1(n7612), .B2(P2_DATAO_REG_0__SCAN_IN), .A(n6723), .ZN(
        n7565) );
  NAND2_X1 U8451 ( .A1(n9024), .A2(n7612), .ZN(n6723) );
  NAND2_X1 U8452 ( .A1(n6983), .A2(n6981), .ZN(n14270) );
  NAND2_X1 U8453 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n6982), .ZN(n6981) );
  INV_X1 U8454 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6982) );
  XNOR2_X1 U8455 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), 
        .ZN(n14269) );
  NAND2_X1 U8456 ( .A1(n14325), .A2(n14295), .ZN(n14297) );
  AOI21_X1 U8457 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n14240), .A(n14239), .ZN(
        n14260) );
  OAI22_X1 U8458 ( .A1(n14303), .A2(n14249), .B1(P1_ADDR_REG_13__SCAN_IN), 
        .B2(n14248), .ZN(n14306) );
  AND2_X1 U8459 ( .A1(n8938), .A2(n8937), .ZN(n8939) );
  AND2_X1 U8460 ( .A1(n7065), .A2(n7063), .ZN(n7062) );
  INV_X1 U8461 ( .A(n7068), .ZN(n7063) );
  NAND2_X1 U8462 ( .A1(n7065), .A2(n7067), .ZN(n7064) );
  OR2_X1 U8463 ( .A1(n9851), .A2(n9850), .ZN(n7067) );
  NAND2_X1 U8464 ( .A1(n8829), .A2(n8828), .ZN(n12538) );
  NAND2_X1 U8465 ( .A1(n11358), .A2(n11357), .ZN(n11356) );
  NAND2_X1 U8466 ( .A1(n6667), .A2(n9764), .ZN(n9765) );
  INV_X1 U8467 ( .A(n9763), .ZN(n6667) );
  NAND2_X1 U8468 ( .A1(n7070), .A2(n9822), .ZN(n12571) );
  AOI21_X1 U8469 ( .B1(n7059), .B2(n12666), .A(n7057), .ZN(n7056) );
  NOR2_X1 U8470 ( .A1(n7060), .A2(n9794), .ZN(n7057) );
  AOI21_X1 U8471 ( .B1(n12833), .B2(n8793), .A(n8792), .ZN(n12842) );
  OR2_X1 U8472 ( .A1(n10518), .A2(n8760), .ZN(n8734) );
  NAND2_X1 U8473 ( .A1(n11356), .A2(n9789), .ZN(n11514) );
  INV_X1 U8474 ( .A(n7072), .ZN(n7071) );
  NAND2_X1 U8475 ( .A1(n9830), .A2(n9832), .ZN(n12620) );
  NAND2_X1 U8476 ( .A1(n8432), .A2(n8431), .ZN(n12624) );
  NAND2_X1 U8477 ( .A1(n7055), .A2(n9795), .ZN(n11833) );
  INV_X1 U8478 ( .A(n7059), .ZN(n7054) );
  INV_X1 U8479 ( .A(n12660), .ZN(n12924) );
  NOR2_X1 U8480 ( .A1(n7487), .A2(n7486), .ZN(n9811) );
  NAND2_X1 U8481 ( .A1(n8466), .A2(n8465), .ZN(n12635) );
  OR2_X1 U8482 ( .A1(n10574), .A2(n8760), .ZN(n8466) );
  XNOR2_X1 U8483 ( .A(n12118), .B(n12528), .ZN(n12112) );
  AND2_X1 U8484 ( .A1(n7050), .A2(n7049), .ZN(n12110) );
  AND2_X1 U8485 ( .A1(n7048), .A2(n6537), .ZN(n12111) );
  AND2_X1 U8486 ( .A1(n9892), .A2(n13063), .ZN(n12380) );
  NAND2_X1 U8487 ( .A1(n12376), .A2(n12381), .ZN(n6664) );
  OR2_X1 U8488 ( .A1(n12376), .A2(n15111), .ZN(n6665) );
  NAND4_X1 U8489 ( .A1(n8824), .A2(n8823), .A3(n8822), .A4(n8821), .ZN(n12773)
         );
  NAND4_X1 U8490 ( .A1(n8526), .A2(n8525), .A3(n8524), .A4(n8523), .ZN(n12673)
         );
  NAND3_X1 U8491 ( .A1(n6805), .A2(n8512), .A3(n8511), .ZN(n15091) );
  NAND2_X1 U8492 ( .A1(n6739), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8512) );
  OR2_X1 U8493 ( .A1(n10732), .A2(n10911), .ZN(n10774) );
  NAND2_X1 U8494 ( .A1(n7032), .A2(n10740), .ZN(n10741) );
  AND2_X1 U8495 ( .A1(n14971), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n14972) );
  AOI21_X1 U8496 ( .B1(n10842), .B2(n10814), .A(n14993), .ZN(n15014) );
  NAND2_X1 U8497 ( .A1(n10860), .A2(n10861), .ZN(n10864) );
  NAND2_X1 U8498 ( .A1(n10864), .A2(n10863), .ZN(n11377) );
  XNOR2_X1 U8499 ( .A(n11374), .B(n6837), .ZN(n15046) );
  INV_X1 U8500 ( .A(n7002), .ZN(n15045) );
  XNOR2_X1 U8501 ( .A(n11549), .B(n11565), .ZN(n11376) );
  NOR2_X1 U8502 ( .A1(n11376), .A2(n11395), .ZN(n11550) );
  XNOR2_X1 U8503 ( .A(n12679), .B(n12688), .ZN(n11792) );
  AND2_X1 U8504 ( .A1(n11788), .A2(n11787), .ZN(n12675) );
  INV_X1 U8505 ( .A(n6770), .ZN(n12705) );
  NAND2_X1 U8506 ( .A1(n6772), .A2(n6773), .ZN(n14360) );
  INV_X1 U8507 ( .A(n7012), .ZN(n6772) );
  NAND2_X1 U8508 ( .A1(n6775), .A2(n15082), .ZN(n6774) );
  XNOR2_X1 U8509 ( .A(n14391), .B(n14390), .ZN(n6775) );
  AND2_X1 U8510 ( .A1(n12466), .A2(n8835), .ZN(n12777) );
  AND2_X1 U8511 ( .A1(n8834), .A2(n8820), .ZN(n12791) );
  AND2_X1 U8512 ( .A1(n12790), .A2(n12789), .ZN(n12951) );
  AOI21_X1 U8513 ( .B1(n12793), .B2(n12815), .A(n12788), .ZN(n12789) );
  OR2_X1 U8514 ( .A1(n12784), .A2(n12922), .ZN(n12790) );
  NAND2_X1 U8515 ( .A1(n6768), .A2(n6767), .ZN(n12957) );
  NAND2_X1 U8516 ( .A1(n6769), .A2(n6964), .ZN(n6768) );
  AOI21_X1 U8517 ( .B1(n12958), .B2(n12815), .A(n12814), .ZN(n6767) );
  AOI21_X1 U8518 ( .B1(n12812), .B2(n12813), .A(n12922), .ZN(n6769) );
  AND2_X1 U8519 ( .A1(n12824), .A2(n12823), .ZN(n12961) );
  INV_X1 U8520 ( .A(n6815), .ZN(n12839) );
  AOI21_X1 U8521 ( .B1(n6820), .B2(n6818), .A(n12334), .ZN(n6815) );
  NAND2_X1 U8522 ( .A1(n6820), .A2(n12206), .ZN(n12855) );
  NAND2_X1 U8523 ( .A1(n8889), .A2(n8888), .ZN(n12863) );
  NAND2_X1 U8524 ( .A1(n6980), .A2(n6497), .ZN(n12884) );
  AOI21_X1 U8525 ( .B1(n12920), .B2(n12921), .A(n6499), .ZN(n12909) );
  NAND2_X1 U8526 ( .A1(n12928), .A2(n12304), .ZN(n12914) );
  OAI21_X1 U8527 ( .B1(n11760), .B2(n6747), .A(n6496), .ZN(n11843) );
  OAI21_X1 U8528 ( .B1(n11765), .B2(n6811), .A(n6522), .ZN(n11847) );
  NAND2_X1 U8529 ( .A1(n11763), .A2(n12274), .ZN(n11782) );
  OAI21_X1 U8530 ( .B1(n8880), .B2(n7280), .A(n7278), .ZN(n11536) );
  NAND2_X1 U8531 ( .A1(n8880), .A2(n8879), .ZN(n11438) );
  INV_X1 U8532 ( .A(n15112), .ZN(n14400) );
  NAND2_X1 U8533 ( .A1(n12144), .A2(n12143), .ZN(n12938) );
  INV_X1 U8534 ( .A(n12938), .ZN(n13010) );
  NAND2_X1 U8535 ( .A1(n6974), .A2(n6973), .ZN(n9887) );
  INV_X1 U8536 ( .A(n12538), .ZN(n13017) );
  INV_X1 U8537 ( .A(n12578), .ZN(n13026) );
  INV_X2 U8538 ( .A(n15173), .ZN(n15175) );
  AND2_X1 U8539 ( .A1(n10723), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13063) );
  INV_X1 U8540 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13065) );
  INV_X1 U8541 ( .A(n9879), .ZN(n10881) );
  NAND2_X1 U8542 ( .A1(n8444), .A2(n8443), .ZN(n8446) );
  NAND2_X1 U8543 ( .A1(n8461), .A2(n8400), .ZN(n8444) );
  INV_X1 U8544 ( .A(SI_16_), .ZN(n15247) );
  INV_X1 U8545 ( .A(SI_15_), .ZN(n15224) );
  NAND2_X1 U8546 ( .A1(n7174), .A2(n6625), .ZN(n8698) );
  NAND2_X1 U8547 ( .A1(n7174), .A2(n8392), .ZN(n8696) );
  INV_X1 U8548 ( .A(SI_14_), .ZN(n15263) );
  INV_X1 U8549 ( .A(SI_11_), .ZN(n15315) );
  NAND2_X1 U8550 ( .A1(n8627), .A2(n8382), .ZN(n8637) );
  NAND2_X1 U8551 ( .A1(n7165), .A2(n7163), .ZN(n8574) );
  NAND2_X1 U8552 ( .A1(n7165), .A2(n8374), .ZN(n8572) );
  NAND2_X1 U8553 ( .A1(n7144), .A2(n8367), .ZN(n8528) );
  NAND2_X1 U8554 ( .A1(n8515), .A2(n8366), .ZN(n7144) );
  INV_X1 U8555 ( .A(SI_1_), .ZN(n7562) );
  CLKBUF_X1 U8556 ( .A(n10710), .Z(n10711) );
  NAND2_X1 U8557 ( .A1(n12400), .A2(n10968), .ZN(n10969) );
  NAND2_X1 U8558 ( .A1(n7303), .A2(n10482), .ZN(n14784) );
  AOI22_X1 U8559 ( .A1(n9187), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n9239), .B2(
        n10333), .ZN(n9042) );
  OAI21_X1 U8560 ( .B1(n13163), .B2(n7323), .A(n7321), .ZN(n13137) );
  AOI21_X1 U8561 ( .B1(n7324), .B2(n7322), .A(n6545), .ZN(n7321) );
  NAND2_X1 U8562 ( .A1(n7324), .A2(n14428), .ZN(n7323) );
  NOR2_X1 U8563 ( .A1(n13100), .A2(n14782), .ZN(n7322) );
  OAI22_X1 U8564 ( .A1(n9664), .A2(n10023), .B1(n10314), .B2(n10098), .ZN(
        n7082) );
  AND2_X1 U8565 ( .A1(n12514), .A2(n12513), .ZN(n6855) );
  NAND2_X1 U8566 ( .A1(n6858), .A2(n11344), .ZN(n11347) );
  INV_X1 U8567 ( .A(n6864), .ZN(n13173) );
  AOI21_X1 U8568 ( .B1(n13123), .B2(n7314), .A(n7312), .ZN(n7311) );
  NAND2_X1 U8569 ( .A1(n7315), .A2(n13123), .ZN(n7313) );
  NAND2_X1 U8570 ( .A1(n9179), .A2(n9178), .ZN(n14456) );
  AND2_X1 U8571 ( .A1(n14428), .A2(n13489), .ZN(n13225) );
  AND2_X1 U8572 ( .A1(n10222), .A2(n10209), .ZN(n14430) );
  NAND2_X1 U8573 ( .A1(n12040), .A2(n10607), .ZN(n10702) );
  NAND2_X1 U8574 ( .A1(n12499), .A2(n12500), .ZN(n6863) );
  INV_X1 U8575 ( .A(n13210), .ZN(n14787) );
  OR2_X1 U8576 ( .A1(n9747), .A2(n9469), .ZN(n9748) );
  XNOR2_X1 U8577 ( .A(n7330), .B(n9432), .ZN(n9747) );
  NAND2_X1 U8578 ( .A1(n9246), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9035) );
  OR2_X1 U8579 ( .A1(n9019), .A2(n10591), .ZN(n9020) );
  AND2_X1 U8580 ( .A1(n14843), .A2(n14842), .ZN(n14845) );
  NAND2_X1 U8581 ( .A1(n13320), .A2(n13523), .ZN(n13532) );
  XNOR2_X1 U8582 ( .A(n13325), .B(n13319), .ZN(n13320) );
  NAND2_X1 U8583 ( .A1(n7122), .A2(n9722), .ZN(n13355) );
  NAND2_X1 U8584 ( .A1(n7124), .A2(n7127), .ZN(n7122) );
  NAND2_X1 U8585 ( .A1(n6710), .A2(n13364), .ZN(n13551) );
  NAND2_X1 U8586 ( .A1(n6711), .A2(n14886), .ZN(n6710) );
  XNOR2_X1 U8587 ( .A(n13362), .B(n13363), .ZN(n6711) );
  NAND2_X1 U8588 ( .A1(n7124), .A2(n7128), .ZN(n13362) );
  NOR2_X1 U8589 ( .A1(n13394), .A2(n9467), .ZN(n13381) );
  OR2_X1 U8590 ( .A1(n13394), .A2(n7471), .ZN(n13379) );
  OAI21_X1 U8591 ( .B1(n13390), .B2(n13391), .A(n6521), .ZN(n13376) );
  OR2_X1 U8592 ( .A1(n11913), .A2(n9664), .ZN(n9298) );
  INV_X1 U8593 ( .A(n13581), .ZN(n13450) );
  NAND2_X1 U8594 ( .A1(n7131), .A2(n7132), .ZN(n13442) );
  NAND2_X1 U8595 ( .A1(n7461), .A2(n9463), .ZN(n13440) );
  NAND2_X1 U8596 ( .A1(n7135), .A2(n7137), .ZN(n13454) );
  NAND2_X1 U8597 ( .A1(n13499), .A2(n9459), .ZN(n13485) );
  OR2_X1 U8598 ( .A1(n10915), .A2(n9664), .ZN(n8995) );
  NAND2_X1 U8599 ( .A1(n9006), .A2(n9005), .ZN(n13600) );
  NAND2_X1 U8600 ( .A1(n11699), .A2(n7480), .ZN(n13516) );
  OAI21_X1 U8601 ( .B1(n11267), .B2(n7108), .A(n7106), .ZN(n14433) );
  AND2_X1 U8602 ( .A1(n7117), .A2(n7116), .ZN(n11312) );
  INV_X1 U8603 ( .A(n9157), .ZN(n7116) );
  INV_X1 U8604 ( .A(n14916), .ZN(n14898) );
  NAND2_X1 U8605 ( .A1(n9451), .A2(n9450), .ZN(n11046) );
  NAND2_X1 U8606 ( .A1(n10989), .A2(n9116), .ZN(n11204) );
  NAND2_X1 U8607 ( .A1(n7466), .A2(n9442), .ZN(n14892) );
  INV_X1 U8608 ( .A(n10267), .ZN(n10944) );
  NAND2_X1 U8609 ( .A1(n14919), .A2(n14907), .ZN(n13472) );
  NAND2_X1 U8610 ( .A1(n7095), .A2(n6942), .ZN(n7451) );
  NOR2_X1 U8611 ( .A1(n13541), .A2(n6716), .ZN(n13544) );
  NAND2_X1 U8612 ( .A1(n6718), .A2(n6717), .ZN(n6716) );
  NAND2_X1 U8613 ( .A1(n13543), .A2(n14945), .ZN(n6717) );
  AND2_X1 U8614 ( .A1(n9273), .A2(n9274), .ZN(n11772) );
  INV_X1 U8615 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10916) );
  INV_X1 U8616 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10631) );
  INV_X1 U8617 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10635) );
  INV_X1 U8618 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10695) );
  INV_X1 U8619 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10430) );
  INV_X1 U8620 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10228) );
  INV_X1 U8621 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10088) );
  INV_X1 U8622 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10084) );
  INV_X1 U8623 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10076) );
  INV_X1 U8624 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10070) );
  INV_X1 U8625 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10064) );
  INV_X1 U8626 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10062) );
  INV_X1 U8627 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10058) );
  INV_X1 U8628 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10060) );
  INV_X1 U8629 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10024) );
  NAND2_X1 U8630 ( .A1(n11594), .A2(n11593), .ZN(n11645) );
  NAND2_X1 U8631 ( .A1(n7224), .A2(n7222), .ZN(n13680) );
  AND2_X1 U8632 ( .A1(n7223), .A2(n12083), .ZN(n7222) );
  NAND2_X1 U8633 ( .A1(n7244), .A2(n7248), .ZN(n11601) );
  OR2_X1 U8634 ( .A1(n13722), .A2(n7249), .ZN(n7244) );
  NAND2_X1 U8635 ( .A1(n7253), .A2(n7256), .ZN(n11958) );
  OR2_X1 U8636 ( .A1(n11858), .A2(n7258), .ZN(n7253) );
  NAND2_X1 U8637 ( .A1(n7942), .A2(n7941), .ZN(n13719) );
  NAND2_X1 U8638 ( .A1(n13680), .A2(n6681), .ZN(n13775) );
  NAND2_X1 U8639 ( .A1(n12079), .A2(n6682), .ZN(n6681) );
  INV_X1 U8640 ( .A(n12084), .ZN(n6682) );
  AOI21_X1 U8641 ( .B1(n7256), .B2(n7258), .A(n6559), .ZN(n7254) );
  NAND2_X1 U8642 ( .A1(n7874), .A2(n7873), .ZN(n14518) );
  INV_X1 U8643 ( .A(n11656), .ZN(n14526) );
  AND2_X1 U8644 ( .A1(n7260), .A2(n6555), .ZN(n11859) );
  OR2_X1 U8645 ( .A1(n10581), .A2(n10580), .ZN(n7243) );
  NAND2_X1 U8646 ( .A1(n7242), .A2(n7241), .ZN(n10919) );
  NAND2_X1 U8647 ( .A1(n7225), .A2(n7230), .ZN(n13783) );
  NAND2_X1 U8648 ( .A1(n13710), .A2(n13736), .ZN(n7225) );
  AND2_X1 U8649 ( .A1(n8288), .A2(n8324), .ZN(n6893) );
  INV_X1 U8650 ( .A(n13728), .ZN(n13840) );
  INV_X1 U8651 ( .A(n11010), .ZN(n13843) );
  INV_X1 U8652 ( .A(n13929), .ZN(n14094) );
  NAND2_X1 U8653 ( .A1(n12013), .A2(n12012), .ZN(n12014) );
  NAND2_X1 U8654 ( .A1(n13964), .A2(n12020), .ZN(n13949) );
  AOI21_X1 U8655 ( .B1(n13943), .B2(n14618), .A(n13942), .ZN(n14114) );
  NAND2_X1 U8656 ( .A1(n13974), .A2(n7372), .ZN(n12011) );
  AND2_X1 U8657 ( .A1(n14000), .A2(n9999), .ZN(n13984) );
  NAND2_X1 U8658 ( .A1(n14005), .A2(n9925), .ZN(n13989) );
  AND2_X1 U8659 ( .A1(n14021), .A2(n9924), .ZN(n14007) );
  NAND2_X1 U8660 ( .A1(n7344), .A2(n9923), .ZN(n14034) );
  NAND2_X1 U8661 ( .A1(n7344), .A2(n7342), .ZN(n14156) );
  OR2_X1 U8662 ( .A1(n11437), .A2(n7670), .ZN(n8028) );
  NAND2_X1 U8663 ( .A1(n14071), .A2(n9921), .ZN(n14049) );
  NAND2_X1 U8664 ( .A1(n7391), .A2(n9982), .ZN(n11868) );
  OR2_X1 U8665 ( .A1(n14473), .A2(n14475), .ZN(n7391) );
  NAND2_X1 U8666 ( .A1(n14474), .A2(n9915), .ZN(n11871) );
  AND2_X1 U8667 ( .A1(n12444), .A2(n10003), .ZN(n14480) );
  NAND2_X1 U8668 ( .A1(n7329), .A2(n9978), .ZN(n11686) );
  NAND2_X1 U8669 ( .A1(n11650), .A2(n11651), .ZN(n7329) );
  AND2_X1 U8670 ( .A1(n6470), .A2(n9908), .ZN(n11424) );
  OR2_X1 U8671 ( .A1(n12490), .A2(n7988), .ZN(n14065) );
  NAND2_X1 U8672 ( .A1(n6481), .A2(n14637), .ZN(n7337) );
  NAND2_X1 U8673 ( .A1(n7362), .A2(n7361), .ZN(n7359) );
  INV_X1 U8674 ( .A(n14677), .ZN(n14488) );
  NAND2_X1 U8675 ( .A1(n14665), .A2(n14480), .ZN(n14083) );
  INV_X1 U8676 ( .A(n14065), .ZN(n14683) );
  AND2_X1 U8677 ( .A1(n14665), .A2(n10465), .ZN(n14677) );
  INV_X1 U8678 ( .A(n14083), .ZN(n14662) );
  AND2_X2 U8679 ( .A1(n11255), .A2(n11254), .ZN(n14776) );
  NAND2_X1 U8680 ( .A1(n14089), .A2(n14679), .ZN(n14090) );
  NOR2_X1 U8681 ( .A1(n14100), .A2(n14099), .ZN(n14101) );
  OR2_X1 U8682 ( .A1(n9950), .A2(n14210), .ZN(n10042) );
  AOI21_X1 U8683 ( .B1(n9274), .B2(n8096), .A(n6530), .ZN(n11827) );
  INV_X1 U8684 ( .A(n10010), .ZN(n14215) );
  OR2_X1 U8685 ( .A1(n8040), .A2(n6910), .ZN(n8041) );
  NAND2_X1 U8686 ( .A1(n7232), .A2(n7231), .ZN(n7540) );
  NAND2_X1 U8687 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n7547), .ZN(n7231) );
  NAND2_X1 U8688 ( .A1(n7543), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7545) );
  INV_X1 U8689 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10637) );
  INV_X1 U8690 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10597) );
  INV_X1 U8691 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10633) );
  INV_X1 U8692 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10685) );
  INV_X1 U8693 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10227) );
  INV_X1 U8694 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10087) );
  NAND2_X1 U8695 ( .A1(n7794), .A2(n7793), .ZN(n7815) );
  INV_X1 U8696 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10082) );
  INV_X1 U8697 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10073) );
  OAI21_X1 U8698 ( .B1(n7718), .B2(n6900), .A(n6898), .ZN(n7763) );
  NAND2_X1 U8699 ( .A1(n7739), .A2(n6869), .ZN(n7743) );
  NOR2_X1 U8700 ( .A1(n7742), .A2(n6900), .ZN(n6869) );
  INV_X1 U8701 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10068) );
  OAI21_X1 U8702 ( .B1(n7717), .B2(n7718), .A(n7739), .ZN(n10071) );
  INV_X1 U8703 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10040) );
  NAND2_X1 U8704 ( .A1(n7688), .A2(n7687), .ZN(n7714) );
  NAND2_X1 U8705 ( .A1(n7684), .A2(n7683), .ZN(n7688) );
  INV_X1 U8706 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10025) );
  INV_X1 U8707 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10020) );
  INV_X1 U8708 ( .A(n14272), .ZN(n14273) );
  NOR2_X1 U8709 ( .A1(n14276), .A2(n15408), .ZN(n14319) );
  OAI21_X1 U8710 ( .B1(n14278), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n15404), .ZN(
        n15395) );
  XNOR2_X1 U8711 ( .A(n6656), .B(n14281), .ZN(n15399) );
  XNOR2_X1 U8712 ( .A(n14283), .B(n13272), .ZN(n14324) );
  NOR2_X1 U8713 ( .A1(n14324), .A2(n14323), .ZN(n14322) );
  XNOR2_X1 U8714 ( .A(n14293), .B(n6999), .ZN(n14327) );
  INV_X1 U8715 ( .A(n14294), .ZN(n6999) );
  NAND2_X1 U8716 ( .A1(n14327), .A2(n14326), .ZN(n14325) );
  NOR2_X1 U8717 ( .A1(n14301), .A2(n14302), .ZN(n14538) );
  OAI21_X1 U8718 ( .B1(n14543), .B2(n14542), .A(n6985), .ZN(n6984) );
  INV_X1 U8719 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6985) );
  NAND2_X1 U8720 ( .A1(n14553), .A2(n6993), .ZN(n14559) );
  INV_X1 U8721 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n6994) );
  INV_X1 U8722 ( .A(n7315), .ZN(n7310) );
  NOR2_X1 U8723 ( .A1(n12604), .A2(n7051), .ZN(n12561) );
  INV_X1 U8724 ( .A(n6669), .ZN(n6668) );
  OAI21_X1 U8725 ( .B1(n13022), .B2(n12649), .A(n12648), .ZN(n6669) );
  AOI21_X1 U8726 ( .B1(n6842), .B2(n6641), .A(n12761), .ZN(n6841) );
  AND2_X1 U8727 ( .A1(n7034), .A2(n6843), .ZN(n6650) );
  AND2_X1 U8728 ( .A1(n6974), .A2(n8871), .ZN(n12474) );
  NAND2_X1 U8729 ( .A1(n6833), .A2(n6644), .ZN(n9889) );
  OAI21_X1 U8730 ( .B1(n11832), .B2(n13076), .A(n7273), .ZN(P3_U3268) );
  NOR2_X1 U8731 ( .A1(n13078), .A2(n15265), .ZN(n7274) );
  NOR2_X1 U8732 ( .A1(n9434), .A2(n9433), .ZN(n9474) );
  AND2_X1 U8733 ( .A1(n13536), .A2(n14916), .ZN(n9433) );
  INV_X1 U8734 ( .A(n6679), .ZN(n6678) );
  OAI21_X1 U8735 ( .B1(n6872), .B2(n13803), .A(n13666), .ZN(n6679) );
  NAND2_X1 U8736 ( .A1(n7266), .A2(n13795), .ZN(n7263) );
  NAND2_X1 U8737 ( .A1(n6589), .A2(n8324), .ZN(n6894) );
  INV_X1 U8738 ( .A(n6988), .ZN(n14330) );
  XNOR2_X1 U8739 ( .A(n15391), .B(n15393), .ZN(n6732) );
  INV_X1 U8740 ( .A(n7309), .ZN(n13202) );
  INV_X1 U8741 ( .A(n14647), .ZN(n6879) );
  CLKBUF_X3 U8742 ( .A(n8119), .Z(n6720) );
  NAND2_X1 U8743 ( .A1(n8889), .A2(n6821), .ZN(n6820) );
  NAND2_X1 U8744 ( .A1(n8353), .A2(n8354), .ZN(n8778) );
  OR2_X1 U8745 ( .A1(n6939), .A2(n11353), .ZN(n6495) );
  INV_X1 U8746 ( .A(n13354), .ZN(n7119) );
  INV_X1 U8747 ( .A(n12897), .ZN(n12900) );
  AND2_X1 U8748 ( .A1(n12311), .A2(n12316), .ZN(n12897) );
  INV_X1 U8749 ( .A(n9746), .ZN(n7446) );
  AND2_X1 U8750 ( .A1(n6746), .A2(n12287), .ZN(n6496) );
  AND2_X1 U8751 ( .A1(n12885), .A2(n6979), .ZN(n6497) );
  AND2_X1 U8752 ( .A1(n6938), .A2(n11249), .ZN(n6498) );
  AND2_X1 U8753 ( .A1(n12930), .A2(n12661), .ZN(n6499) );
  INV_X1 U8754 ( .A(n9628), .ZN(n7412) );
  AND2_X1 U8755 ( .A1(n7946), .A2(n15327), .ZN(n6500) );
  OR2_X1 U8756 ( .A1(n8859), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n6501) );
  INV_X1 U8757 ( .A(n12921), .ZN(n6765) );
  AND2_X1 U8758 ( .A1(n9746), .A2(n7103), .ZN(n6502) );
  AND2_X1 U8759 ( .A1(n7109), .A2(n9200), .ZN(n6503) );
  INV_X2 U8760 ( .A(n9647), .ZN(n9514) );
  NAND2_X1 U8761 ( .A1(n6905), .A2(n6910), .ZN(n7374) );
  NAND2_X1 U8762 ( .A1(n12669), .A2(n9786), .ZN(n6504) );
  AND2_X1 U8763 ( .A1(n7631), .A2(SI_2_), .ZN(n6505) );
  NOR2_X1 U8764 ( .A1(n13022), .A2(n12811), .ZN(n6506) );
  NOR2_X1 U8765 ( .A1(n9795), .A2(n12666), .ZN(n6507) );
  AOI21_X1 U8766 ( .B1(n13466), .B2(n7139), .A(n6594), .ZN(n7137) );
  OR2_X1 U8767 ( .A1(n14443), .A2(n11709), .ZN(n6509) );
  AND2_X1 U8768 ( .A1(n9539), .A2(n9538), .ZN(n6510) );
  AND2_X1 U8769 ( .A1(n9527), .A2(n9526), .ZN(n6511) );
  AND2_X1 U8770 ( .A1(n6498), .A2(n6937), .ZN(n6512) );
  NAND2_X1 U8771 ( .A1(n9310), .A2(n9309), .ZN(n13558) );
  INV_X1 U8772 ( .A(n13575), .ZN(n6950) );
  NAND2_X1 U8773 ( .A1(n11581), .A2(n7054), .ZN(n6513) );
  AND2_X1 U8774 ( .A1(n8596), .A2(n8595), .ZN(n11383) );
  INV_X1 U8775 ( .A(n11383), .ZN(n6839) );
  AND2_X1 U8776 ( .A1(n7283), .A2(n7285), .ZN(n6514) );
  NAND2_X1 U8777 ( .A1(n6640), .A2(n6907), .ZN(n6515) );
  AND2_X1 U8778 ( .A1(n11787), .A2(n12688), .ZN(n6516) );
  AND2_X1 U8779 ( .A1(n10746), .A2(n10739), .ZN(n15082) );
  OR3_X1 U8780 ( .A1(n14660), .A2(n14647), .A3(n6881), .ZN(n6517) );
  INV_X1 U8781 ( .A(n8154), .ZN(n6928) );
  AND2_X1 U8782 ( .A1(n15082), .A2(n7035), .ZN(n6518) );
  INV_X1 U8783 ( .A(n14886), .ZN(n7099) );
  NAND3_X1 U8784 ( .A1(n8507), .A2(n8506), .A3(n6801), .ZN(n9772) );
  NAND2_X2 U8785 ( .A1(n9043), .A2(n9042), .ZN(n14906) );
  AND2_X1 U8786 ( .A1(n11129), .A2(n8551), .ZN(n6520) );
  INV_X1 U8787 ( .A(n9128), .ZN(n7092) );
  OR2_X1 U8788 ( .A1(n13563), .A2(n13246), .ZN(n6521) );
  INV_X1 U8789 ( .A(n9795), .ZN(n7060) );
  NAND2_X1 U8790 ( .A1(n10785), .A2(n8498), .ZN(n8874) );
  AND2_X1 U8791 ( .A1(n7282), .A2(n6810), .ZN(n6522) );
  AND2_X1 U8792 ( .A1(n11423), .A2(n9908), .ZN(n6523) );
  NAND2_X1 U8793 ( .A1(n9241), .A2(n9240), .ZN(n13591) );
  NAND2_X1 U8794 ( .A1(n9681), .A2(n9680), .ZN(n9707) );
  INV_X1 U8795 ( .A(n9018), .ZN(n9264) );
  OR2_X1 U8796 ( .A1(n8328), .A2(n7398), .ZN(n6524) );
  OR2_X1 U8797 ( .A1(n8328), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n6525) );
  NAND2_X1 U8798 ( .A1(n12825), .A2(n6966), .ZN(n6964) );
  OAI211_X1 U8799 ( .C1(n8529), .C2(SI_3_), .A(n8520), .B(n8519), .ZN(n15129)
         );
  NAND2_X1 U8800 ( .A1(n7536), .A2(n7271), .ZN(n6526) );
  INV_X1 U8801 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8963) );
  AND2_X1 U8802 ( .A1(n14006), .A2(n9924), .ZN(n6527) );
  OR2_X1 U8803 ( .A1(n11353), .A2(n11077), .ZN(n6528) );
  AND2_X1 U8804 ( .A1(n8479), .A2(n7033), .ZN(n6529) );
  AND2_X1 U8805 ( .A1(n6906), .A2(n8093), .ZN(n6530) );
  INV_X1 U8806 ( .A(n9767), .ZN(n10674) );
  NAND2_X1 U8807 ( .A1(n8497), .A2(n8873), .ZN(n9767) );
  AND2_X1 U8808 ( .A1(n13992), .A2(n6875), .ZN(n6531) );
  NOR2_X1 U8809 ( .A1(n8886), .A2(n6826), .ZN(n6532) );
  AND2_X1 U8810 ( .A1(n12182), .A2(n6752), .ZN(n6533) );
  OR2_X1 U8811 ( .A1(n9800), .A2(n12926), .ZN(n6534) );
  AND2_X1 U8812 ( .A1(n14407), .A2(n12664), .ZN(n6535) );
  NAND2_X1 U8813 ( .A1(n14018), .A2(n9997), .ZN(n14004) );
  AND2_X1 U8814 ( .A1(n6964), .A2(n6965), .ZN(n6536) );
  OAI211_X1 U8815 ( .C1(n8529), .C2(n7562), .A(n8485), .B(n8484), .ZN(n8498)
         );
  OR2_X1 U8816 ( .A1(n12662), .A2(n9806), .ZN(n6537) );
  INV_X1 U8817 ( .A(n9722), .ZN(n7123) );
  AND2_X1 U8818 ( .A1(n6497), .A2(n6758), .ZN(n6538) );
  NOR2_X1 U8819 ( .A1(n9229), .A2(n7139), .ZN(n6539) );
  AND2_X1 U8820 ( .A1(n13983), .A2(n9999), .ZN(n6540) );
  OR2_X1 U8821 ( .A1(n12938), .A2(n12153), .ZN(n6541) );
  OR2_X1 U8822 ( .A1(n7488), .A2(n15327), .ZN(n6542) );
  NAND2_X1 U8823 ( .A1(n8178), .A2(n8177), .ZN(n14112) );
  INV_X1 U8824 ( .A(n14112), .ZN(n6872) );
  NAND2_X1 U8825 ( .A1(n9219), .A2(n9218), .ZN(n13607) );
  INV_X1 U8826 ( .A(n13607), .ZN(n6948) );
  INV_X1 U8827 ( .A(n14998), .ZN(n7023) );
  NAND2_X1 U8828 ( .A1(n7842), .A2(n7841), .ZN(n11900) );
  OR2_X1 U8829 ( .A1(n13505), .A2(n13253), .ZN(n6543) );
  NAND2_X1 U8830 ( .A1(n8995), .A2(n8994), .ZN(n13595) );
  INV_X1 U8831 ( .A(n13595), .ZN(n6945) );
  XOR2_X1 U8832 ( .A(n13535), .B(n13240), .Z(n6544) );
  AND3_X1 U8833 ( .A1(n13132), .A2(n13225), .A3(n13243), .ZN(n6545) );
  INV_X1 U8834 ( .A(n12206), .ZN(n6819) );
  AND2_X1 U8835 ( .A1(n12312), .A2(n12314), .ZN(n12913) );
  INV_X1 U8836 ( .A(n12913), .ZN(n6763) );
  AND2_X1 U8837 ( .A1(n12500), .A2(n12501), .ZN(n6547) );
  AND2_X1 U8838 ( .A1(n13607), .A2(n13254), .ZN(n6548) );
  OR2_X1 U8839 ( .A1(n13450), .A2(n13249), .ZN(n6549) );
  OR2_X1 U8840 ( .A1(n13839), .A2(n11494), .ZN(n6550) );
  INV_X1 U8841 ( .A(n7804), .ZN(n7201) );
  INV_X1 U8842 ( .A(n8075), .ZN(n7181) );
  NAND2_X1 U8843 ( .A1(n12281), .A2(n12665), .ZN(n6551) );
  OR2_X1 U8844 ( .A1(n11497), .A2(n11512), .ZN(n6552) );
  AND2_X1 U8845 ( .A1(n11353), .A2(n11077), .ZN(n6553) );
  NAND2_X1 U8846 ( .A1(n9166), .A2(n9165), .ZN(n11353) );
  OR2_X1 U8847 ( .A1(n12975), .A2(n9831), .ZN(n6554) );
  NAND2_X1 U8848 ( .A1(n11855), .A2(n11856), .ZN(n6555) );
  AND2_X1 U8849 ( .A1(n12670), .A2(n15149), .ZN(n6556) );
  INV_X1 U8850 ( .A(n13433), .ZN(n13425) );
  XNOR2_X1 U8851 ( .A(n13575), .B(n13248), .ZN(n13433) );
  NAND2_X1 U8852 ( .A1(n8503), .A2(n8478), .ZN(n8516) );
  AND2_X1 U8853 ( .A1(n14125), .A2(n13958), .ZN(n6557) );
  NOR2_X1 U8854 ( .A1(n7868), .A2(SI_13_), .ZN(n6558) );
  INV_X1 U8855 ( .A(n14133), .ZN(n13981) );
  NAND2_X1 U8856 ( .A1(n8125), .A2(n8124), .ZN(n14133) );
  AND2_X1 U8857 ( .A1(n11955), .A2(n11957), .ZN(n6559) );
  AND2_X1 U8858 ( .A1(n13455), .A2(n7136), .ZN(n6560) );
  AND2_X1 U8859 ( .A1(n9638), .A2(n9637), .ZN(n6561) );
  OR2_X1 U8860 ( .A1(n9663), .A2(n10024), .ZN(n6562) );
  INV_X1 U8861 ( .A(n13967), .ZN(n14117) );
  NAND2_X1 U8862 ( .A1(n8157), .A2(n8156), .ZN(n13967) );
  OR2_X1 U8863 ( .A1(n6837), .A2(n11374), .ZN(n6563) );
  INV_X1 U8864 ( .A(n7776), .ZN(n7205) );
  AND2_X1 U8865 ( .A1(n9919), .A2(n9918), .ZN(n6564) );
  AND2_X1 U8866 ( .A1(n11052), .A2(n13260), .ZN(n6565) );
  NAND2_X1 U8867 ( .A1(n7906), .A2(n7905), .ZN(n14503) );
  AND2_X1 U8868 ( .A1(n8138), .A2(n6933), .ZN(n6566) );
  OR2_X1 U8869 ( .A1(n10842), .A2(n10841), .ZN(n6567) );
  AND2_X1 U8870 ( .A1(n11345), .A2(n11344), .ZN(n6568) );
  NAND2_X1 U8871 ( .A1(n7715), .A2(SI_7_), .ZN(n7738) );
  INV_X1 U8872 ( .A(n7738), .ZN(n6900) );
  AND2_X1 U8873 ( .A1(n13391), .A2(n6521), .ZN(n6569) );
  INV_X1 U8874 ( .A(n7984), .ZN(n7214) );
  INV_X1 U8875 ( .A(n7115), .ZN(n7114) );
  NAND2_X1 U8876 ( .A1(n6528), .A2(n11270), .ZN(n7115) );
  AND2_X1 U8877 ( .A1(n10971), .A2(n10968), .ZN(n6570) );
  AND2_X1 U8878 ( .A1(n9824), .A2(n9822), .ZN(n6571) );
  OR2_X1 U8879 ( .A1(n7281), .A2(n11516), .ZN(n6572) );
  AND2_X1 U8880 ( .A1(n7071), .A2(n9832), .ZN(n6573) );
  AND2_X1 U8881 ( .A1(n10001), .A2(n10000), .ZN(n6574) );
  NAND2_X1 U8882 ( .A1(n8228), .A2(n8227), .ZN(n14096) );
  INV_X1 U8883 ( .A(n8563), .ZN(n6962) );
  INV_X1 U8884 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8909) );
  INV_X1 U8885 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n7547) );
  INV_X1 U8886 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7535) );
  INV_X1 U8887 ( .A(n7490), .ZN(n7049) );
  NOR2_X1 U8888 ( .A1(n12926), .A2(n9803), .ZN(n7490) );
  AND2_X1 U8889 ( .A1(n7304), .A2(n11729), .ZN(n6575) );
  OR2_X1 U8890 ( .A1(n14464), .A2(n11077), .ZN(n6576) );
  NOR2_X1 U8891 ( .A1(n9790), .A2(n12668), .ZN(n6577) );
  NOR2_X1 U8892 ( .A1(n11900), .A2(n13833), .ZN(n6578) );
  NOR2_X1 U8893 ( .A1(n11589), .A2(n13836), .ZN(n6579) );
  NOR2_X1 U8894 ( .A1(n14159), .A2(n14056), .ZN(n6580) );
  NOR2_X1 U8895 ( .A1(n14503), .A2(n13831), .ZN(n6581) );
  AND2_X1 U8896 ( .A1(n8295), .A2(n13691), .ZN(n6582) );
  AND2_X1 U8897 ( .A1(n13450), .A2(n9465), .ZN(n6583) );
  AND2_X1 U8898 ( .A1(n12578), .A2(n12653), .ZN(n6968) );
  NOR2_X1 U8899 ( .A1(n9851), .A2(n7066), .ZN(n6584) );
  XNOR2_X1 U8900 ( .A(n13098), .B(n10267), .ZN(n10247) );
  INV_X1 U8901 ( .A(n7448), .ZN(n7447) );
  OAI22_X1 U8902 ( .A1(n13332), .A2(n7449), .B1(n13344), .B2(n13133), .ZN(
        n7448) );
  NAND2_X1 U8903 ( .A1(n13982), .A2(n10000), .ZN(n6585) );
  AND2_X1 U8904 ( .A1(n9627), .A2(n9626), .ZN(n6586) );
  INV_X1 U8905 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8347) );
  INV_X1 U8906 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10018) );
  AND2_X1 U8907 ( .A1(n7836), .A2(n15315), .ZN(n6587) );
  INV_X1 U8908 ( .A(n7090), .ZN(n7089) );
  NAND2_X1 U8909 ( .A1(n7091), .A2(n9129), .ZN(n7090) );
  INV_X1 U8910 ( .A(n7109), .ZN(n7108) );
  NOR2_X1 U8911 ( .A1(n9185), .A2(n7110), .ZN(n7109) );
  NAND2_X1 U8912 ( .A1(n11903), .A2(n11901), .ZN(n6588) );
  INV_X1 U8913 ( .A(n7316), .ZN(n7314) );
  NAND2_X1 U8914 ( .A1(n12511), .A2(n12512), .ZN(n7316) );
  NOR2_X1 U8915 ( .A1(n8319), .A2(n8318), .ZN(n6589) );
  AND4_X1 U8916 ( .A1(n8490), .A2(n8489), .A3(n8488), .A4(n8487), .ZN(n6590)
         );
  INV_X1 U8917 ( .A(n6590), .ZN(n8497) );
  AND2_X1 U8918 ( .A1(n12089), .A2(n12090), .ZN(n6591) );
  INV_X1 U8919 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n6849) );
  AND2_X1 U8920 ( .A1(n6978), .A2(n12659), .ZN(n6592) );
  AND3_X1 U8921 ( .A1(n12531), .A2(n12535), .A3(n12642), .ZN(n6593) );
  NOR2_X1 U8922 ( .A1(n9431), .A2(n13251), .ZN(n6594) );
  NAND2_X1 U8923 ( .A1(n7250), .A2(n11644), .ZN(n6595) );
  OR2_X1 U8924 ( .A1(n14732), .A2(n13838), .ZN(n6596) );
  OR2_X1 U8925 ( .A1(n12624), .A2(n9831), .ZN(n12333) );
  INV_X1 U8926 ( .A(n9731), .ZN(n14891) );
  XNOR2_X1 U8927 ( .A(n14112), .B(n12463), .ZN(n13940) );
  OR2_X1 U8928 ( .A1(n6510), .A2(n9542), .ZN(n6597) );
  OR2_X1 U8929 ( .A1(n9651), .A2(n7428), .ZN(n6598) );
  AND2_X1 U8930 ( .A1(n6873), .A2(n6872), .ZN(n6599) );
  OR2_X1 U8931 ( .A1(n9620), .A2(n6601), .ZN(n6600) );
  AND2_X1 U8932 ( .A1(n9618), .A2(n9617), .ZN(n6601) );
  NOR2_X1 U8933 ( .A1(n12191), .A2(n12162), .ZN(n6602) );
  AND2_X1 U8934 ( .A1(n7078), .A2(n8909), .ZN(n6603) );
  OR2_X1 U8935 ( .A1(n7046), .A2(n9807), .ZN(n6604) );
  NAND2_X1 U8936 ( .A1(n14955), .A2(n13259), .ZN(n6605) );
  AND2_X1 U8937 ( .A1(n7320), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6606) );
  NOR2_X1 U8938 ( .A1(P3_IR_REG_28__SCAN_IN), .A2(P3_IR_REG_29__SCAN_IN), .ZN(
        n6607) );
  AND2_X1 U8939 ( .A1(n13974), .A2(n9930), .ZN(n6608) );
  NAND2_X1 U8940 ( .A1(n12673), .A2(n8537), .ZN(n6609) );
  AND2_X1 U8941 ( .A1(n7374), .A2(n7373), .ZN(n6610) );
  AND2_X1 U8942 ( .A1(n12840), .A2(n6816), .ZN(n6611) );
  OR2_X1 U8943 ( .A1(n7427), .A2(n9652), .ZN(n6612) );
  OR2_X1 U8944 ( .A1(n9555), .A2(n9554), .ZN(n6613) );
  OR2_X1 U8945 ( .A1(n9529), .A2(n6511), .ZN(n6614) );
  NAND2_X1 U8946 ( .A1(n8127), .A2(n7187), .ZN(n6615) );
  NOR2_X1 U8947 ( .A1(n7412), .A2(n6586), .ZN(n6616) );
  AND2_X1 U8948 ( .A1(n7015), .A2(n7014), .ZN(n6617) );
  OR2_X1 U8949 ( .A1(n6915), .A2(n6500), .ZN(n6618) );
  INV_X1 U8950 ( .A(n7076), .ZN(n7075) );
  NAND2_X1 U8951 ( .A1(n7077), .A2(n9789), .ZN(n7076) );
  OR2_X1 U8952 ( .A1(n7423), .A2(n6561), .ZN(n6619) );
  INV_X1 U8953 ( .A(n7463), .ZN(n7462) );
  NAND2_X1 U8954 ( .A1(n10920), .A2(n10921), .ZN(n6620) );
  OR2_X1 U8955 ( .A1(n9553), .A2(n7407), .ZN(n6621) );
  INV_X1 U8956 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8974) );
  NAND2_X1 U8957 ( .A1(n7184), .A2(n8214), .ZN(n6622) );
  NAND2_X1 U8958 ( .A1(n8168), .A2(n7190), .ZN(n6623) );
  INV_X1 U8959 ( .A(n15053), .ZN(n6837) );
  NOR2_X1 U8960 ( .A1(n8602), .A2(n8583), .ZN(n6624) );
  AND2_X1 U8961 ( .A1(n7173), .A2(n8392), .ZN(n6625) );
  INV_X1 U8962 ( .A(n15149), .ZN(n6766) );
  INV_X1 U8963 ( .A(SI_17_), .ZN(n15327) );
  INV_X1 U8964 ( .A(n8039), .ZN(n6910) );
  AND2_X1 U8965 ( .A1(n11702), .A2(n6947), .ZN(n6626) );
  AND4_X1 U8966 ( .A1(n8648), .A2(n8647), .A3(n8646), .A4(n8645), .ZN(n11834)
         );
  INV_X1 U8967 ( .A(n12263), .ZN(n7277) );
  NAND2_X1 U8968 ( .A1(n7388), .A2(n7387), .ZN(n11947) );
  NAND2_X1 U8969 ( .A1(n12991), .A2(n12311), .ZN(n12883) );
  NOR2_X1 U8970 ( .A1(n8094), .A2(n6909), .ZN(n6627) );
  INV_X1 U8971 ( .A(n13445), .ZN(n6951) );
  INV_X1 U8972 ( .A(n7824), .ZN(n7199) );
  NOR2_X1 U8973 ( .A1(n8036), .A2(n8039), .ZN(n6628) );
  NAND2_X1 U8974 ( .A1(n7305), .A2(n11729), .ZN(n14424) );
  NAND2_X1 U8975 ( .A1(n8479), .A2(n8480), .ZN(n10753) );
  INV_X1 U8976 ( .A(n10753), .ZN(n6976) );
  OR2_X1 U8977 ( .A1(n13007), .A2(n12926), .ZN(n6629) );
  OR2_X1 U8978 ( .A1(n12118), .A2(n12662), .ZN(n6630) );
  OR2_X1 U8979 ( .A1(n11926), .A2(n9804), .ZN(n12544) );
  INV_X1 U8980 ( .A(n12655), .ZN(n12828) );
  AND2_X1 U8981 ( .A1(n11699), .A2(n9458), .ZN(n6631) );
  INV_X1 U8982 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n6952) );
  AND2_X1 U8983 ( .A1(n6907), .A2(n6910), .ZN(n6632) );
  AND2_X1 U8984 ( .A1(n7391), .A2(n7389), .ZN(n6633) );
  AND2_X1 U8985 ( .A1(n6839), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n6634) );
  NOR2_X1 U8986 ( .A1(n12555), .A2(n11916), .ZN(n6635) );
  INV_X1 U8987 ( .A(n9386), .ZN(n7104) );
  NAND2_X1 U8988 ( .A1(n9385), .A2(n9384), .ZN(n9386) );
  OR2_X1 U8989 ( .A1(n7903), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n6636) );
  INV_X1 U8990 ( .A(n6836), .ZN(n6835) );
  NAND2_X1 U8991 ( .A1(n8871), .A2(n15183), .ZN(n6836) );
  AND2_X1 U8992 ( .A1(n10227), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n6637) );
  NAND2_X1 U8993 ( .A1(n6867), .A2(n6863), .ZN(n12502) );
  INV_X1 U8994 ( .A(n7843), .ZN(n7195) );
  OR2_X1 U8995 ( .A1(n13352), .A2(n13210), .ZN(n6638) );
  AND2_X1 U8996 ( .A1(n6980), .A2(n6979), .ZN(n6639) );
  NAND2_X1 U8997 ( .A1(n6627), .A2(n8115), .ZN(n6640) );
  INV_X1 U8998 ( .A(n13479), .ZN(n7477) );
  INV_X1 U8999 ( .A(n14428), .ZN(n14782) );
  AND2_X1 U9000 ( .A1(n10222), .A2(n10221), .ZN(n14428) );
  NAND2_X1 U9001 ( .A1(n7359), .A2(n9903), .ZN(n11139) );
  NAND2_X1 U9002 ( .A1(n11365), .A2(n11364), .ZN(n11731) );
  NAND2_X1 U9003 ( .A1(n7337), .A2(n9972), .ZN(n11098) );
  AOI21_X1 U9004 ( .B1(n11195), .B2(n6972), .A(n6970), .ZN(n11128) );
  XNOR2_X1 U9005 ( .A(n8913), .B(P3_IR_REG_26__SCAN_IN), .ZN(n8936) );
  INV_X1 U9006 ( .A(n8936), .ZN(n6671) );
  INV_X1 U9007 ( .A(n8121), .ZN(n6931) );
  INV_X1 U9008 ( .A(n11658), .ZN(n7378) );
  NAND2_X1 U9009 ( .A1(n8940), .A2(n8905), .ZN(n8943) );
  NAND2_X1 U9010 ( .A1(n9792), .A2(n9791), .ZN(n11581) );
  AND2_X1 U9011 ( .A1(n15082), .A2(n7037), .ZN(n6641) );
  INV_X1 U9012 ( .A(SI_20_), .ZN(n15324) );
  AND2_X1 U9013 ( .A1(n11692), .A2(n6885), .ZN(n6642) );
  AND2_X1 U9014 ( .A1(n11356), .A2(n7075), .ZN(n6643) );
  OR2_X1 U9015 ( .A1(n15183), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n6644) );
  INV_X1 U9016 ( .A(n6535), .ZN(n7285) );
  INV_X1 U9017 ( .A(n6880), .ZN(n14646) );
  NOR2_X1 U9018 ( .A1(n14660), .A2(n6881), .ZN(n6880) );
  INV_X1 U9019 ( .A(n11553), .ZN(n7010) );
  NAND2_X1 U9020 ( .A1(n7002), .A2(n6563), .ZN(n7001) );
  INV_X1 U9021 ( .A(n8454), .ZN(n12163) );
  AND3_X1 U9022 ( .A1(n14755), .A2(n10466), .A3(n10464), .ZN(n13795) );
  INV_X1 U9023 ( .A(n11052), .ZN(n6938) );
  NAND3_X1 U9024 ( .A1(n8496), .A2(n8495), .A3(n8494), .ZN(n8873) );
  INV_X1 U9025 ( .A(n14934), .ZN(n6940) );
  NAND2_X1 U9026 ( .A1(n9147), .A2(n9146), .ZN(n14955) );
  INV_X1 U9027 ( .A(n14955), .ZN(n6937) );
  AND2_X1 U9028 ( .A1(n12744), .A2(n7041), .ZN(n6645) );
  INV_X1 U9029 ( .A(n14961), .ZN(n13614) );
  INV_X1 U9030 ( .A(n15071), .ZN(n7000) );
  AND2_X1 U9031 ( .A1(n8862), .A2(n12196), .ZN(n12922) );
  NAND2_X1 U9032 ( .A1(n7038), .A2(n7036), .ZN(n7035) );
  AND2_X1 U9033 ( .A1(n14209), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6646) );
  NOR2_X1 U9034 ( .A1(n8825), .A2(n7169), .ZN(n7168) );
  AND2_X1 U9035 ( .A1(n10576), .A2(n7221), .ZN(n6647) );
  INV_X1 U9036 ( .A(n6727), .ZN(n9472) );
  AND2_X1 U9037 ( .A1(n7243), .A2(n10638), .ZN(n6648) );
  AND2_X1 U9038 ( .A1(n7032), .A2(n7031), .ZN(n6649) );
  NAND2_X1 U9039 ( .A1(n6987), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n6986) );
  OR2_X1 U9040 ( .A1(n10506), .A2(n14906), .ZN(n10529) );
  NOR2_X2 U9041 ( .A1(n14328), .A2(n14298), .ZN(n14331) );
  NAND2_X1 U9042 ( .A1(n13344), .A2(n13349), .ZN(n13340) );
  NAND2_X1 U9043 ( .A1(n13450), .A2(n13458), .ZN(n13445) );
  NAND2_X1 U9044 ( .A1(n14543), .A2(n14542), .ZN(n14541) );
  NAND2_X1 U9045 ( .A1(n14550), .A2(n14551), .ZN(n14549) );
  NAND2_X2 U9046 ( .A1(n6949), .A2(n9031), .ZN(n6653) );
  NAND4_X1 U9047 ( .A1(n13538), .A2(n7100), .A3(n7097), .A4(n7101), .ZN(n6942)
         );
  INV_X1 U9048 ( .A(n12378), .ZN(n6666) );
  NAND2_X1 U9049 ( .A1(n8771), .A2(n8770), .ZN(n8413) );
  NAND2_X1 U9050 ( .A1(n7147), .A2(n7150), .ZN(n8403) );
  NAND2_X1 U9051 ( .A1(n7155), .A2(n7154), .ZN(n8653) );
  NAND2_X1 U9052 ( .A1(n7172), .A2(n7170), .ZN(n8712) );
  NAND2_X1 U9053 ( .A1(n8390), .A2(n8389), .ZN(n8681) );
  NAND2_X1 U9054 ( .A1(n6663), .A2(n12377), .ZN(n12386) );
  AOI21_X1 U9055 ( .B1(n12801), .B2(n12354), .A(n12166), .ZN(n12786) );
  OAI21_X1 U9056 ( .B1(n7298), .B2(n7296), .A(n6602), .ZN(n7295) );
  NAND2_X1 U9057 ( .A1(n13153), .A2(n13152), .ZN(n13151) );
  NOR2_X2 U9058 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n9013) );
  NOR2_X1 U9059 ( .A1(n13204), .A2(n13205), .ZN(n6857) );
  INV_X1 U9060 ( .A(n7008), .ZN(n11554) );
  INV_X1 U9061 ( .A(n14391), .ZN(n6842) );
  INV_X1 U9062 ( .A(n7082), .ZN(n6714) );
  NOR2_X1 U9063 ( .A1(n12676), .A2(n12677), .ZN(n12678) );
  NAND2_X1 U9064 ( .A1(n7009), .A2(n7004), .ZN(n11789) );
  NOR2_X1 U9065 ( .A1(n14997), .A2(n7028), .ZN(n10823) );
  INV_X1 U9066 ( .A(n10970), .ZN(n10971) );
  NAND3_X1 U9067 ( .A1(n6841), .A2(n6650), .A3(n6846), .ZN(P3_U3201) );
  OAI21_X1 U9068 ( .B1(n7717), .B2(n6900), .A(n7742), .ZN(n6899) );
  OAI21_X1 U9069 ( .B1(n12499), .B2(n6547), .A(n6865), .ZN(n6703) );
  NAND2_X1 U9070 ( .A1(n6651), .A2(n7566), .ZN(n7583) );
  INV_X1 U9071 ( .A(n7568), .ZN(n6651) );
  NAND2_X1 U9072 ( .A1(n7564), .A2(n7582), .ZN(n7568) );
  AND2_X1 U9073 ( .A1(n7611), .A2(n7586), .ZN(n10017) );
  INV_X1 U9074 ( .A(n7585), .ZN(n6652) );
  NAND2_X1 U9075 ( .A1(n9231), .A2(n9370), .ZN(n9374) );
  NAND2_X1 U9076 ( .A1(n7583), .A2(n7582), .ZN(n7633) );
  NAND2_X1 U9077 ( .A1(n10621), .A2(n10620), .ZN(n10710) );
  NAND3_X1 U9078 ( .A1(n13113), .A2(n13112), .A3(n6638), .ZN(P2_U3186) );
  NAND2_X1 U9079 ( .A1(n6702), .A2(n6859), .ZN(n6864) );
  NAND2_X1 U9080 ( .A1(n10478), .A2(n10477), .ZN(n7303) );
  OAI21_X1 U9081 ( .B1(n13182), .B2(n7313), .A(n7311), .ZN(n13204) );
  NOR2_X2 U9082 ( .A1(n13212), .A2(n6855), .ZN(n13153) );
  NAND2_X1 U9083 ( .A1(n6654), .A2(n10618), .ZN(n10703) );
  NAND2_X1 U9084 ( .A1(n10617), .A2(n10610), .ZN(n6654) );
  OR2_X1 U9085 ( .A1(n7688), .A2(n7687), .ZN(n7689) );
  NAND2_X1 U9086 ( .A1(n10603), .A2(n12033), .ZN(n12040) );
  NAND2_X1 U9087 ( .A1(n13158), .A2(n13092), .ZN(n13097) );
  INV_X1 U9088 ( .A(n7561), .ZN(n7563) );
  INV_X1 U9089 ( .A(n10703), .ZN(n10611) );
  NAND2_X1 U9090 ( .A1(n7664), .A2(n7663), .ZN(n7668) );
  OAI211_X1 U9091 ( .C1(n13108), .C2(n13107), .A(n13147), .B(n14428), .ZN(
        n13113) );
  NAND2_X1 U9092 ( .A1(n9446), .A2(n9445), .ZN(n10988) );
  OAI21_X1 U9093 ( .B1(n13247), .B2(n13569), .A(n13412), .ZN(n13395) );
  OAI22_X4 U9094 ( .A1(n13361), .A2(n9468), .B1(n13167), .B2(n13371), .ZN(
        n13348) );
  NAND2_X1 U9095 ( .A1(n7454), .A2(n7087), .ZN(n7456) );
  NAND2_X1 U9096 ( .A1(n13483), .A2(n9460), .ZN(n13465) );
  OAI21_X1 U9097 ( .B1(n11471), .B2(n9455), .A(n9456), .ZN(n14439) );
  NAND2_X1 U9098 ( .A1(n14539), .A2(n14537), .ZN(n14543) );
  INV_X1 U9099 ( .A(n14280), .ZN(n6656) );
  OAI21_X1 U9100 ( .B1(n14557), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n14310), .ZN(
        n14345) );
  NAND2_X1 U9101 ( .A1(n14301), .A2(n14302), .ZN(n14540) );
  NAND2_X1 U9102 ( .A1(n6995), .A2(n14549), .ZN(n14555) );
  OAI21_X1 U9103 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(n14277), .A(n14318), .ZN(
        n15406) );
  OAI21_X1 U9104 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n15383), .A(n15382), .ZN(
        n15392) );
  OAI21_X1 U9105 ( .B1(n14555), .B2(n14554), .A(n6994), .ZN(n6993) );
  NAND2_X1 U9106 ( .A1(n6988), .A2(n6986), .ZN(n14301) );
  NAND2_X1 U9107 ( .A1(n6984), .A2(n14541), .ZN(n14547) );
  NAND2_X1 U9108 ( .A1(n14270), .A2(n14269), .ZN(n6657) );
  NAND2_X1 U9109 ( .A1(n14271), .A2(n14272), .ZN(n6983) );
  NAND2_X1 U9110 ( .A1(n15395), .A2(n15396), .ZN(n15394) );
  OAI21_X1 U9111 ( .B1(n14345), .B2(n14344), .A(n6998), .ZN(n6997) );
  XNOR2_X1 U9112 ( .A(n10530), .B(n13098), .ZN(n12032) );
  OR2_X1 U9113 ( .A1(n14331), .A2(n14332), .ZN(n6988) );
  XNOR2_X1 U9114 ( .A(n15392), .B(n6732), .ZN(SUB_1596_U4) );
  NAND2_X1 U9115 ( .A1(n13499), .A2(n7475), .ZN(n13483) );
  INV_X1 U9116 ( .A(n9451), .ZN(n7454) );
  NAND2_X1 U9117 ( .A1(n10504), .A2(n10503), .ZN(n10502) );
  NAND2_X1 U9118 ( .A1(n6658), .A2(n9957), .ZN(n11112) );
  NAND2_X1 U9119 ( .A1(n14106), .A2(n12475), .ZN(n12477) );
  INV_X1 U9120 ( .A(n13998), .ZN(n6662) );
  NAND2_X1 U9121 ( .A1(n6911), .A2(n6915), .ZN(n7393) );
  NAND2_X1 U9122 ( .A1(n12023), .A2(n12022), .ZN(n14106) );
  NAND2_X2 U9123 ( .A1(n14000), .A2(n6540), .ZN(n13982) );
  NAND2_X2 U9124 ( .A1(n6662), .A2(n6661), .ZN(n14000) );
  NAND2_X1 U9125 ( .A1(n8024), .A2(n15324), .ZN(n8025) );
  NAND3_X1 U9126 ( .A1(n6666), .A2(n6665), .A3(n6664), .ZN(n6663) );
  NAND2_X1 U9127 ( .A1(n8665), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8390) );
  NAND2_X1 U9128 ( .A1(n8413), .A2(n8412), .ZN(n8414) );
  NAND2_X1 U9129 ( .A1(n6670), .A2(n6668), .ZN(P3_U3180) );
  NAND2_X1 U9130 ( .A1(n12643), .A2(n12642), .ZN(n6670) );
  AOI21_X2 U9131 ( .B1(n8911), .B2(n8916), .A(n6671), .ZN(n8920) );
  NAND2_X1 U9132 ( .A1(n9827), .A2(n9826), .ZN(n9830) );
  AOI21_X2 U9133 ( .B1(n11023), .B2(n11022), .A(n9779), .ZN(n11060) );
  NOR2_X2 U9134 ( .A1(n10886), .A2(n10887), .ZN(n10885) );
  NAND2_X1 U9135 ( .A1(n11882), .A2(n9797), .ZN(n11923) );
  INV_X1 U9136 ( .A(n11884), .ZN(n6673) );
  NAND3_X1 U9137 ( .A1(n9837), .A2(n12601), .A3(n12828), .ZN(n12556) );
  NAND2_X1 U9138 ( .A1(n8717), .A2(n6952), .ZN(n8462) );
  NAND3_X1 U9139 ( .A1(n9646), .A2(n6696), .A3(n6598), .ZN(n7426) );
  NAND2_X1 U9140 ( .A1(n7419), .A2(n7422), .ZN(n9644) );
  NAND2_X1 U9141 ( .A1(n7429), .A2(n7430), .ZN(n9548) );
  NAND2_X1 U9142 ( .A1(n6676), .A2(n6675), .ZN(n6674) );
  OAI22_X2 U9143 ( .A1(n9504), .A2(n7418), .B1(n7417), .B2(n9505), .ZN(n9512)
         );
  NAND2_X1 U9144 ( .A1(n9712), .A2(n9711), .ZN(n9718) );
  NOR2_X1 U9145 ( .A1(n6686), .A2(n6616), .ZN(n7410) );
  NAND2_X1 U9146 ( .A1(n6677), .A2(n6674), .ZN(n9581) );
  INV_X1 U9147 ( .A(n9560), .ZN(n6676) );
  NAND2_X1 U9148 ( .A1(n6684), .A2(n6683), .ZN(n6677) );
  NAND2_X1 U9149 ( .A1(n6680), .A2(n6678), .ZN(P1_U3214) );
  NAND2_X1 U9150 ( .A1(n13660), .A2(n13795), .ZN(n6680) );
  NAND2_X2 U9151 ( .A1(n6488), .A2(n7494), .ZN(n8328) );
  AOI21_X2 U9152 ( .B1(n13775), .B2(n13774), .A(n6591), .ZN(n13689) );
  NAND2_X1 U9153 ( .A1(n7255), .A2(n7254), .ZN(n11998) );
  NAND2_X1 U9154 ( .A1(n11750), .A2(n11749), .ZN(n11858) );
  NAND2_X1 U9155 ( .A1(n7247), .A2(n7245), .ZN(n11677) );
  NAND2_X1 U9156 ( .A1(n7424), .A2(n7425), .ZN(n9534) );
  NAND2_X1 U9157 ( .A1(n9560), .A2(n9559), .ZN(n6684) );
  INV_X1 U9158 ( .A(n9496), .ZN(n6730) );
  NAND3_X1 U9159 ( .A1(n9536), .A2(n9537), .A3(n6597), .ZN(n7429) );
  NAND2_X1 U9160 ( .A1(n7426), .A2(n6612), .ZN(n9657) );
  NAND2_X1 U9161 ( .A1(n7431), .A2(n7432), .ZN(n9625) );
  OAI22_X1 U9162 ( .A1(n9689), .A2(n9688), .B1(n9693), .B2(n9692), .ZN(n6691)
         );
  NOR2_X1 U9163 ( .A1(n9625), .A2(n9624), .ZN(n6686) );
  NAND2_X1 U9164 ( .A1(n6689), .A2(n6688), .ZN(n6687) );
  NAND2_X1 U9165 ( .A1(n6698), .A2(n6697), .ZN(n7411) );
  NAND3_X1 U9166 ( .A1(n9477), .A2(n9647), .A3(n10214), .ZN(n9480) );
  NAND2_X1 U9167 ( .A1(n6695), .A2(n6694), .ZN(n9658) );
  NAND2_X1 U9168 ( .A1(n6693), .A2(n6692), .ZN(n9537) );
  OR2_X1 U9169 ( .A1(n9512), .A2(n9511), .ZN(n7483) );
  NAND2_X1 U9170 ( .A1(n9685), .A2(n9684), .ZN(n6690) );
  NAND2_X1 U9171 ( .A1(n9534), .A2(n9533), .ZN(n6693) );
  NAND2_X1 U9172 ( .A1(n9657), .A2(n9656), .ZN(n6695) );
  NAND2_X1 U9173 ( .A1(n6701), .A2(n6700), .ZN(n6696) );
  AOI21_X1 U9174 ( .B1(n9548), .B2(n9547), .A(n9545), .ZN(n9546) );
  NAND2_X1 U9175 ( .A1(n9625), .A2(n9624), .ZN(n6698) );
  OAI21_X1 U9176 ( .B1(n9751), .B2(n6699), .A(n9750), .ZN(n9755) );
  AOI21_X1 U9177 ( .B1(n9749), .B2(n9472), .A(n9748), .ZN(n6699) );
  NAND2_X1 U9178 ( .A1(n6722), .A2(n6721), .ZN(n7421) );
  NAND2_X1 U9179 ( .A1(n9644), .A2(n9643), .ZN(n6701) );
  AND2_X2 U9180 ( .A1(n6864), .A2(n12505), .ZN(n13184) );
  INV_X1 U9181 ( .A(n6703), .ZN(n6702) );
  NAND2_X1 U9182 ( .A1(n10619), .A2(n10618), .ZN(n10621) );
  NAND3_X1 U9183 ( .A1(n12040), .A2(n10611), .A3(n10607), .ZN(n10619) );
  NAND2_X1 U9184 ( .A1(n9620), .A2(n6601), .ZN(n7432) );
  NAND3_X1 U9185 ( .A1(n9549), .A2(n6621), .A3(n6508), .ZN(n7406) );
  NAND3_X1 U9186 ( .A1(n7420), .A2(n7421), .A3(n6619), .ZN(n7419) );
  NAND2_X1 U9187 ( .A1(n6707), .A2(n6704), .ZN(n9504) );
  NAND2_X1 U9188 ( .A1(n6706), .A2(n6705), .ZN(n6704) );
  INV_X1 U9189 ( .A(n9498), .ZN(n6706) );
  NAND2_X1 U9190 ( .A1(n6731), .A2(n6730), .ZN(n6707) );
  NAND2_X1 U9191 ( .A1(n9103), .A2(n9726), .ZN(n10990) );
  NAND2_X1 U9192 ( .A1(n9077), .A2(n9076), .ZN(n14884) );
  NAND2_X2 U9193 ( .A1(n6714), .A2(n6562), .ZN(n10267) );
  NOR2_X2 U9194 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n6715) );
  NAND2_X1 U9195 ( .A1(n7084), .A2(n7083), .ZN(n13480) );
  NAND2_X4 U9196 ( .A1(n10098), .A2(n6720), .ZN(n9664) );
  NAND3_X1 U9197 ( .A1(n6935), .A2(n6546), .A3(n6934), .ZN(n8985) );
  NAND2_X1 U9198 ( .A1(n11706), .A2(n9214), .ZN(n13512) );
  NAND2_X1 U9199 ( .A1(n13496), .A2(n6543), .ZN(n7084) );
  NAND2_X1 U9200 ( .A1(n7081), .A2(n9089), .ZN(n11223) );
  NAND2_X1 U9201 ( .A1(n7080), .A2(n9049), .ZN(n10526) );
  NAND2_X1 U9202 ( .A1(n7896), .A2(n7895), .ZN(n6783) );
  NAND3_X1 U9203 ( .A1(n6719), .A2(n6903), .A3(n6515), .ZN(n8116) );
  NAND2_X1 U9204 ( .A1(n6914), .A2(n6500), .ZN(n7392) );
  NAND3_X1 U9205 ( .A1(n7303), .A2(n10486), .A3(n10482), .ZN(n10489) );
  XNOR2_X1 U9206 ( .A(n14906), .B(n13098), .ZN(n10484) );
  XNOR2_X2 U9207 ( .A(n7616), .B(n7632), .ZN(n10038) );
  NAND2_X1 U9208 ( .A1(n13151), .A2(n6853), .ZN(n13082) );
  OR2_X2 U9209 ( .A1(n9488), .A2(n9487), .ZN(n7416) );
  AND2_X2 U9210 ( .A1(n9475), .A2(n9469), .ZN(n9647) );
  OAI211_X1 U9211 ( .C1(n12540), .C2(n12541), .A(n6724), .B(n12539), .ZN(
        P3_U3160) );
  NAND2_X1 U9212 ( .A1(n12540), .A2(n6593), .ZN(n6724) );
  NAND2_X1 U9213 ( .A1(n9792), .A2(n7053), .ZN(n7058) );
  NOR2_X2 U9214 ( .A1(n8859), .A2(n7301), .ZN(n8904) );
  NAND2_X1 U9215 ( .A1(n13239), .A2(n7324), .ZN(n13147) );
  NAND2_X1 U9216 ( .A1(n7309), .A2(n13124), .ZN(n6856) );
  OAI21_X2 U9217 ( .B1(n12640), .B2(n9850), .A(n7068), .ZN(n12540) );
  NAND2_X1 U9218 ( .A1(n7058), .A2(n7056), .ZN(n11884) );
  NOR2_X2 U9219 ( .A1(n8715), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n8717) );
  NAND2_X1 U9220 ( .A1(n8451), .A2(n8700), .ZN(n8715) );
  AND2_X2 U9221 ( .A1(n13239), .A2(n13104), .ZN(n13108) );
  INV_X1 U9222 ( .A(n7632), .ZN(n6726) );
  NAND2_X1 U9223 ( .A1(n7409), .A2(n7408), .ZN(n9636) );
  OAI21_X2 U9224 ( .B1(n7416), .B2(n7413), .A(n7414), .ZN(n9498) );
  NAND2_X2 U9225 ( .A1(n9080), .A2(n9079), .ZN(n14934) );
  NAND2_X1 U9226 ( .A1(n7411), .A2(n7410), .ZN(n7409) );
  OR2_X1 U9227 ( .A1(n9671), .A2(n9016), .ZN(n9023) );
  NOR2_X2 U9228 ( .A1(n9477), .A2(n10214), .ZN(n9476) );
  NAND2_X1 U9229 ( .A1(n9498), .A2(n9497), .ZN(n6731) );
  XNOR2_X1 U9230 ( .A(n14288), .B(n14289), .ZN(n15402) );
  NAND2_X1 U9231 ( .A1(n14555), .A2(n14554), .ZN(n14553) );
  NAND2_X1 U9232 ( .A1(n14345), .A2(n14344), .ZN(n14343) );
  NOR2_X1 U9233 ( .A1(n14547), .A2(n14546), .ZN(n14545) );
  NAND2_X1 U9234 ( .A1(n14331), .A2(n14332), .ZN(n6987) );
  NOR2_X1 U9235 ( .A1(n15381), .A2(n15380), .ZN(n15383) );
  NAND2_X1 U9236 ( .A1(n7235), .A2(n7233), .ZN(n13671) );
  XNOR2_X1 U9237 ( .A(n6733), .B(n12444), .ZN(n10918) );
  OAI22_X1 U9238 ( .A1(n14705), .A2(n12454), .B1(n10641), .B2(n12453), .ZN(
        n6733) );
  NOR2_X1 U9239 ( .A1(n10581), .A2(n10642), .ZN(n7239) );
  NOR2_X1 U9240 ( .A1(n10576), .A2(n7221), .ZN(n10575) );
  NAND2_X1 U9241 ( .A1(n8346), .A2(n8530), .ZN(n8859) );
  NAND2_X1 U9242 ( .A1(n12762), .A2(n15078), .ZN(n6846) );
  NAND4_X2 U9243 ( .A1(n9013), .A2(n7405), .A3(n7404), .A4(n7403), .ZN(n9104)
         );
  NAND2_X1 U9244 ( .A1(n7466), .A2(n7465), .ZN(n14894) );
  OAI21_X1 U9245 ( .B1(n13453), .B2(n7463), .A(n7459), .ZN(n13434) );
  NAND2_X2 U9246 ( .A1(n8472), .A2(n8355), .ZN(n12148) );
  NAND2_X1 U9247 ( .A1(n11760), .A2(n6496), .ZN(n6743) );
  NAND2_X1 U9248 ( .A1(n6743), .A2(n6744), .ZN(n11915) );
  NAND2_X1 U9249 ( .A1(n6955), .A2(n6753), .ZN(n13068) );
  NAND2_X1 U9250 ( .A1(n12920), .A2(n6538), .ZN(n6754) );
  NAND2_X1 U9251 ( .A1(n6754), .A2(n6755), .ZN(n12872) );
  NAND3_X1 U9252 ( .A1(n6520), .A2(n11409), .A3(n6960), .ZN(n6958) );
  NAND4_X1 U9253 ( .A1(n14393), .A2(n14392), .A3(n14394), .A4(n6774), .ZN(
        P3_U3200) );
  NAND2_X1 U9254 ( .A1(n10834), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n6776) );
  XNOR2_X2 U9255 ( .A(n8504), .B(n8503), .ZN(n10834) );
  NAND3_X1 U9256 ( .A1(n6777), .A2(n10758), .A3(n6776), .ZN(n10819) );
  NAND2_X1 U9257 ( .A1(n6777), .A2(n6776), .ZN(n10759) );
  XNOR2_X1 U9258 ( .A(n10820), .B(n10837), .ZN(n14971) );
  NOR2_X1 U9259 ( .A1(n14972), .A2(n10821), .ZN(n14999) );
  NAND4_X1 U9260 ( .A1(n7526), .A2(n6781), .A3(P1_ADDR_REG_19__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n6780) );
  NAND4_X1 U9261 ( .A1(n7529), .A2(n7527), .A3(n7528), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n6782) );
  INV_X2 U9262 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7529) );
  OR2_X2 U9263 ( .A1(n7947), .A2(n7488), .ZN(n6914) );
  NAND3_X1 U9264 ( .A1(n6786), .A2(n6898), .A3(n6784), .ZN(n6897) );
  OR2_X2 U9265 ( .A1(n8024), .A2(n15324), .ZN(n7491) );
  NAND2_X1 U9266 ( .A1(n6494), .A2(n7765), .ZN(n6795) );
  NAND2_X1 U9267 ( .A1(n6794), .A2(n6796), .ZN(n6792) );
  NAND2_X1 U9268 ( .A1(n7767), .A2(n6794), .ZN(n6793) );
  OAI21_X1 U9269 ( .B1(n7767), .B2(n6796), .A(n6794), .ZN(n7847) );
  NAND2_X1 U9270 ( .A1(n8070), .A2(n8089), .ZN(n9272) );
  OAI21_X1 U9271 ( .B1(n6798), .B2(SI_4_), .A(n7663), .ZN(n7635) );
  MUX2_X1 U9272 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n7530), .Z(n6798) );
  INV_X1 U9273 ( .A(n6800), .ZN(n6799) );
  OAI22_X1 U9274 ( .A1(n8760), .A2(n10028), .B1(SI_2_), .B2(n8529), .ZN(n6800)
         );
  NAND2_X2 U9275 ( .A1(n8482), .A2(n6720), .ZN(n8529) );
  INV_X1 U9276 ( .A(n6802), .ZN(n6801) );
  INV_X1 U9277 ( .A(n15129), .ZN(n6803) );
  INV_X1 U9278 ( .A(n6806), .ZN(n6805) );
  NAND2_X1 U9279 ( .A1(n11765), .A2(n6522), .ZN(n6807) );
  NAND2_X1 U9280 ( .A1(n6807), .A2(n6808), .ZN(n11918) );
  NAND2_X1 U9281 ( .A1(n8889), .A2(n6813), .ZN(n6812) );
  NAND2_X1 U9282 ( .A1(n6812), .A2(n6611), .ZN(n8890) );
  NAND2_X1 U9283 ( .A1(n12901), .A2(n6532), .ZN(n6823) );
  NAND2_X1 U9284 ( .A1(n6823), .A2(n6824), .ZN(n12876) );
  NAND2_X1 U9285 ( .A1(n6955), .A2(n6827), .ZN(n6830) );
  NAND2_X1 U9286 ( .A1(n6832), .A2(n8903), .ZN(n6833) );
  AND2_X1 U9287 ( .A1(n8903), .A2(n8871), .ZN(n6973) );
  INV_X1 U9288 ( .A(n7631), .ZN(n7630) );
  NAND2_X1 U9289 ( .A1(n6850), .A2(n7634), .ZN(n7637) );
  OAI21_X1 U9290 ( .B1(n7633), .B2(n6505), .A(n6851), .ZN(n6850) );
  INV_X1 U9291 ( .A(n6852), .ZN(n6851) );
  AND2_X2 U9292 ( .A1(n6857), .A2(n6856), .ZN(n13212) );
  NAND2_X2 U9293 ( .A1(n6858), .A2(n6568), .ZN(n11365) );
  NAND2_X2 U9294 ( .A1(n13163), .A2(n13100), .ZN(n13239) );
  NAND2_X2 U9295 ( .A1(n13097), .A2(n13160), .ZN(n13163) );
  NAND2_X1 U9296 ( .A1(n12499), .A2(n6860), .ZN(n6859) );
  XNOR2_X1 U9297 ( .A(n10961), .B(n10962), .ZN(n10721) );
  XNOR2_X1 U9298 ( .A(n14946), .B(n6725), .ZN(n10961) );
  NAND2_X2 U9299 ( .A1(n6868), .A2(n9107), .ZN(n14946) );
  NAND2_X1 U9300 ( .A1(n12484), .A2(n12485), .ZN(n13935) );
  NAND2_X1 U9301 ( .A1(n12484), .A2(n6870), .ZN(n6871) );
  INV_X1 U9302 ( .A(n14660), .ZN(n6876) );
  NAND2_X1 U9303 ( .A1(n6877), .A2(n6876), .ZN(n11427) );
  XNOR2_X2 U9304 ( .A(n6882), .B(n7535), .ZN(n14206) );
  OAI21_X2 U9305 ( .B1(n8328), .B2(n7396), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6882) );
  NAND2_X1 U9306 ( .A1(n11692), .A2(n6883), .ZN(n11949) );
  OAI22_X1 U9307 ( .A1(n8230), .A2(n6889), .B1(n8231), .B2(n6888), .ZN(n8260)
         );
  OAI211_X1 U9308 ( .C1(n8320), .C2(n6894), .A(n6891), .B(n6890), .ZN(P1_U3242) );
  NAND3_X1 U9309 ( .A1(n8320), .A2(n8291), .A3(n6893), .ZN(n6890) );
  INV_X1 U9310 ( .A(n6892), .ZN(n6891) );
  NAND2_X1 U9311 ( .A1(n7375), .A2(n7491), .ZN(n7373) );
  INV_X1 U9312 ( .A(n7491), .ZN(n6905) );
  NAND3_X1 U9313 ( .A1(n7374), .A2(n7373), .A3(n6627), .ZN(n6906) );
  NAND3_X1 U9314 ( .A1(n7374), .A2(n7373), .A3(n8069), .ZN(n8095) );
  OR2_X1 U9315 ( .A1(n7947), .A2(n6542), .ZN(n6911) );
  NAND2_X1 U9316 ( .A1(n7947), .A2(n6618), .ZN(n6913) );
  NAND2_X1 U9317 ( .A1(n7790), .A2(n7789), .ZN(n7794) );
  NAND2_X1 U9318 ( .A1(n8139), .A2(n8138), .ZN(n8151) );
  NOR2_X1 U9319 ( .A1(n9104), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n6935) );
  NAND2_X1 U9320 ( .A1(n9366), .A2(n8965), .ZN(n6936) );
  NAND2_X1 U9321 ( .A1(n11209), .A2(n6512), .ZN(n6939) );
  INV_X1 U9322 ( .A(n6939), .ZN(n11317) );
  NOR2_X2 U9323 ( .A1(n14896), .A2(n11216), .ZN(n11217) );
  NOR2_X2 U9324 ( .A1(n13536), .A2(n6943), .ZN(n13538) );
  NAND4_X1 U9325 ( .A1(n6954), .A2(n8340), .A3(n8341), .A4(n8339), .ZN(n8345)
         );
  NAND2_X1 U9326 ( .A1(n6958), .A2(n6957), .ZN(n11328) );
  AOI21_X1 U9327 ( .B1(n6959), .B2(n11409), .A(n6556), .ZN(n6957) );
  NOR2_X1 U9328 ( .A1(n11185), .A2(n6962), .ZN(n6961) );
  NAND2_X1 U9329 ( .A1(n6964), .A2(n6963), .ZN(n8809) );
  INV_X1 U9330 ( .A(n6968), .ZN(n6965) );
  NAND2_X1 U9331 ( .A1(n11034), .A2(n6971), .ZN(n6969) );
  NAND2_X1 U9332 ( .A1(n6969), .A2(n6609), .ZN(n6970) );
  INV_X1 U9333 ( .A(n8872), .ZN(n6975) );
  NAND2_X1 U9334 ( .A1(n6975), .A2(n15106), .ZN(n6974) );
  INV_X1 U9335 ( .A(n6980), .ZN(n12895) );
  NAND2_X1 U9336 ( .A1(n13051), .A2(n12911), .ZN(n6979) );
  NAND2_X1 U9337 ( .A1(n8516), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8518) );
  NAND2_X1 U9338 ( .A1(n8531), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8532) );
  NAND2_X1 U9339 ( .A1(n8859), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8860) );
  NAND2_X1 U9340 ( .A1(n6501), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8856) );
  NAND2_X1 U9341 ( .A1(n8857), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8855) );
  NAND2_X1 U9342 ( .A1(n8943), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8906) );
  NAND2_X1 U9343 ( .A1(n7079), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8913) );
  NAND2_X1 U9344 ( .A1(n8912), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8910) );
  NAND2_X1 U9345 ( .A1(n8699), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8701) );
  OAI21_X1 U9346 ( .B1(n8638), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8640) );
  AOI21_X1 U9347 ( .B1(n11554), .B2(n6516), .A(n7003), .ZN(n7004) );
  INV_X1 U9348 ( .A(n7015), .ZN(n12725) );
  NAND2_X1 U9349 ( .A1(n7016), .A2(n7018), .ZN(n15018) );
  INV_X1 U9350 ( .A(n7020), .ZN(n7016) );
  NOR2_X1 U9351 ( .A1(n7020), .A2(n7017), .ZN(n15017) );
  NAND2_X1 U9352 ( .A1(n7018), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7017) );
  NOR2_X1 U9353 ( .A1(n14999), .A2(n14998), .ZN(n14997) );
  NAND2_X1 U9354 ( .A1(n14391), .A2(n6518), .ZN(n7034) );
  NAND2_X1 U9355 ( .A1(n11923), .A2(n6604), .ZN(n7045) );
  AND2_X1 U9356 ( .A1(n7052), .A2(n12655), .ZN(n7051) );
  NAND2_X1 U9357 ( .A1(n12640), .A2(n7062), .ZN(n7061) );
  OAI211_X1 U9358 ( .C1(n12640), .C2(n7064), .A(n12642), .B(n7061), .ZN(n9873)
         );
  NAND2_X1 U9359 ( .A1(n12640), .A2(n12641), .ZN(n12639) );
  NAND2_X1 U9360 ( .A1(n8940), .A2(n7078), .ZN(n8912) );
  NAND2_X1 U9361 ( .A1(n8940), .A2(n6603), .ZN(n7079) );
  XNOR2_X1 U9362 ( .A(n8453), .B(n8452), .ZN(n8898) );
  XNOR2_X1 U9363 ( .A(n8910), .B(n8909), .ZN(n8916) );
  NAND2_X1 U9364 ( .A1(n10526), .A2(n10525), .ZN(n9062) );
  NAND2_X1 U9365 ( .A1(n10507), .A2(n10508), .ZN(n7080) );
  NAND2_X1 U9366 ( .A1(n11223), .A2(n9727), .ZN(n9103) );
  NAND2_X1 U9367 ( .A1(n14884), .A2(n14891), .ZN(n7081) );
  NAND2_X1 U9368 ( .A1(n10098), .A2(n10022), .ZN(n9663) );
  INV_X1 U9369 ( .A(n11047), .ZN(n7087) );
  INV_X1 U9370 ( .A(n10989), .ZN(n7088) );
  OAI21_X1 U9371 ( .B1(n10989), .B2(n7092), .A(n7089), .ZN(n11048) );
  NAND2_X1 U9372 ( .A1(n13390), .A2(n7125), .ZN(n7124) );
  AOI21_X1 U9373 ( .B1(n13390), .B2(n7120), .A(n7119), .ZN(n7118) );
  NAND3_X1 U9374 ( .A1(n7132), .A2(n13441), .A3(n7131), .ZN(n7130) );
  NAND2_X1 U9375 ( .A1(n9229), .A2(n13466), .ZN(n7135) );
  AND2_X1 U9376 ( .A1(n13595), .A2(n13186), .ZN(n7139) );
  INV_X1 U9377 ( .A(n7140), .ZN(n7145) );
  NAND2_X1 U9378 ( .A1(n8515), .A2(n7145), .ZN(n7143) );
  NAND2_X1 U9379 ( .A1(n8459), .A2(n7148), .ZN(n7147) );
  NAND2_X1 U9380 ( .A1(n8625), .A2(n7156), .ZN(n7155) );
  NAND2_X1 U9381 ( .A1(n8811), .A2(n7168), .ZN(n7166) );
  NAND2_X1 U9382 ( .A1(n8681), .A2(n6625), .ZN(n7172) );
  OAI22_X1 U9383 ( .A1(n7704), .A2(n7176), .B1(n7703), .B2(n7175), .ZN(n7725)
         );
  NAND3_X1 U9384 ( .A1(n8060), .A2(n8059), .A3(n7178), .ZN(n7180) );
  NAND3_X1 U9385 ( .A1(n8195), .A2(n8194), .A3(n6622), .ZN(n7183) );
  INV_X1 U9386 ( .A(n8213), .ZN(n7184) );
  NAND3_X1 U9387 ( .A1(n8106), .A2(n8105), .A3(n6615), .ZN(n7186) );
  INV_X1 U9388 ( .A(n8126), .ZN(n7187) );
  NAND3_X1 U9389 ( .A1(n8149), .A2(n8148), .A3(n6623), .ZN(n7189) );
  INV_X1 U9390 ( .A(n8167), .ZN(n7190) );
  NAND2_X1 U9391 ( .A1(n7191), .A2(n7192), .ZN(n7922) );
  NAND3_X1 U9392 ( .A1(n7827), .A2(n7193), .A3(n7826), .ZN(n7191) );
  NAND2_X1 U9393 ( .A1(n7843), .A2(n7845), .ZN(n7194) );
  AND2_X1 U9394 ( .A1(n14475), .A2(n7884), .ZN(n7196) );
  OAI21_X1 U9395 ( .B1(n7803), .B2(n7202), .A(n7200), .ZN(n7823) );
  NAND2_X1 U9396 ( .A1(n7197), .A2(n7198), .ZN(n7822) );
  NAND2_X1 U9397 ( .A1(n7803), .A2(n7200), .ZN(n7197) );
  OAI21_X1 U9398 ( .B1(n7752), .B2(n7208), .A(n7206), .ZN(n7775) );
  NAND2_X1 U9399 ( .A1(n7203), .A2(n7204), .ZN(n7774) );
  NAND2_X1 U9400 ( .A1(n7752), .A2(n7206), .ZN(n7203) );
  NAND2_X1 U9401 ( .A1(n7983), .A2(n7212), .ZN(n7209) );
  NAND2_X1 U9402 ( .A1(n7209), .A2(n7210), .ZN(n8009) );
  NAND3_X1 U9403 ( .A1(n7508), .A2(n7220), .A3(n7219), .ZN(n7546) );
  NOR2_X1 U9404 ( .A1(n10575), .A2(n6647), .ZN(n13857) );
  NAND2_X1 U9405 ( .A1(n10457), .A2(n10458), .ZN(n7221) );
  NAND2_X1 U9406 ( .A1(n13710), .A2(n7226), .ZN(n7224) );
  OAI21_X1 U9407 ( .B1(n13710), .B2(n7229), .A(n7226), .ZN(n13782) );
  OAI21_X1 U9408 ( .B1(n13710), .B2(n13737), .A(n13736), .ZN(n13735) );
  AOI21_X1 U9409 ( .B1(n13737), .B2(n13736), .A(n12075), .ZN(n7230) );
  OAI21_X1 U9410 ( .B1(n7538), .B2(n14199), .A(P1_IR_REG_20__SCAN_IN), .ZN(
        n7232) );
  NAND2_X1 U9411 ( .A1(n13687), .A2(n7236), .ZN(n7235) );
  NAND2_X1 U9412 ( .A1(n7239), .A2(n7238), .ZN(n7242) );
  AND3_X2 U9413 ( .A1(n7241), .A2(n7242), .A3(n6620), .ZN(n10929) );
  INV_X1 U9414 ( .A(n7243), .ZN(n10640) );
  NAND2_X1 U9415 ( .A1(n13722), .A2(n7248), .ZN(n7247) );
  INV_X1 U9416 ( .A(n11593), .ZN(n7251) );
  NAND2_X1 U9417 ( .A1(n13722), .A2(n11505), .ZN(n11594) );
  NAND2_X1 U9418 ( .A1(n11858), .A2(n7256), .ZN(n7255) );
  NAND2_X1 U9419 ( .A1(n13657), .A2(n7262), .ZN(n7261) );
  OAI211_X1 U9420 ( .C1(n13657), .C2(n7263), .A(n7261), .B(n12465), .ZN(
        P1_U3220) );
  NOR2_X1 U9421 ( .A1(n12458), .A2(n12451), .ZN(n7267) );
  NAND2_X1 U9422 ( .A1(n12458), .A2(n12451), .ZN(n7268) );
  INV_X1 U9423 ( .A(n12458), .ZN(n7269) );
  NAND3_X1 U9424 ( .A1(n7744), .A2(n7270), .A3(n7508), .ZN(n7955) );
  INV_X2 U9425 ( .A(n7272), .ZN(n14348) );
  MUX2_X1 U9426 ( .A(n10745), .B(n10726), .S(n14348), .Z(n10727) );
  MUX2_X1 U9427 ( .A(n10730), .B(n10731), .S(n14348), .Z(n10902) );
  MUX2_X1 U9428 ( .A(n10765), .B(n10766), .S(n14348), .Z(n10768) );
  MUX2_X1 U9429 ( .A(n10806), .B(n10807), .S(n14348), .Z(n10808) );
  MUX2_X1 U9430 ( .A(P3_REG1_REG_4__SCAN_IN), .B(P3_REG2_REG_4__SCAN_IN), .S(
        n14348), .Z(n10813) );
  MUX2_X1 U9431 ( .A(n10815), .B(n10816), .S(n14348), .Z(n10817) );
  MUX2_X1 U9432 ( .A(P3_REG1_REG_6__SCAN_IN), .B(P3_REG2_REG_6__SCAN_IN), .S(
        n14348), .Z(n10852) );
  MUX2_X1 U9433 ( .A(P3_REG1_REG_7__SCAN_IN), .B(P3_REG2_REG_7__SCAN_IN), .S(
        n14348), .Z(n10856) );
  MUX2_X1 U9434 ( .A(P3_REG1_REG_8__SCAN_IN), .B(P3_REG2_REG_8__SCAN_IN), .S(
        n14348), .Z(n11381) );
  MUX2_X1 U9435 ( .A(n15185), .B(n15047), .S(n14348), .Z(n11386) );
  MUX2_X1 U9436 ( .A(n11387), .B(n11388), .S(n14348), .Z(n11389) );
  MUX2_X1 U9437 ( .A(n11394), .B(n11395), .S(n14348), .Z(n11566) );
  MUX2_X1 U9438 ( .A(P3_REG1_REG_12__SCAN_IN), .B(P3_REG2_REG_12__SCAN_IN), 
        .S(n14348), .Z(n11794) );
  MUX2_X1 U9439 ( .A(P3_REG1_REG_13__SCAN_IN), .B(P3_REG2_REG_13__SCAN_IN), 
        .S(n14348), .Z(n12687) );
  MUX2_X1 U9440 ( .A(P3_REG1_REG_15__SCAN_IN), .B(P3_REG2_REG_15__SCAN_IN), 
        .S(n14348), .Z(n12718) );
  MUX2_X1 U9441 ( .A(P3_REG1_REG_16__SCAN_IN), .B(P3_REG2_REG_16__SCAN_IN), 
        .S(n14348), .Z(n12737) );
  MUX2_X1 U9442 ( .A(P3_REG1_REG_17__SCAN_IN), .B(P3_REG2_REG_17__SCAN_IN), 
        .S(n14348), .Z(n12740) );
  MUX2_X1 U9443 ( .A(P3_REG1_REG_18__SCAN_IN), .B(P3_REG2_REG_18__SCAN_IN), 
        .S(n14348), .Z(n14383) );
  MUX2_X1 U9444 ( .A(n12714), .B(n12715), .S(n14348), .Z(n12716) );
  NAND2_X1 U9445 ( .A1(n10746), .A2(n7272), .ZN(n15036) );
  AOI21_X1 U9446 ( .B1(n14348), .B2(P3_STATE_REG_SCAN_IN), .A(n7274), .ZN(
        n7273) );
  NAND2_X1 U9447 ( .A1(n7275), .A2(n7276), .ZN(n8881) );
  NAND2_X1 U9448 ( .A1(n8880), .A2(n7278), .ZN(n7275) );
  NAND2_X1 U9449 ( .A1(n12929), .A2(n7287), .ZN(n7286) );
  CLKBUF_X1 U9450 ( .A(n13182), .Z(n7308) );
  NOR2_X1 U9451 ( .A1(n7308), .A2(n12509), .ZN(n13217) );
  NAND2_X1 U9452 ( .A1(n9370), .A2(n7317), .ZN(n9373) );
  AND4_X2 U9453 ( .A1(n7524), .A2(n7523), .A3(n7496), .A4(n7525), .ZN(n11010)
         );
  NAND2_X1 U9454 ( .A1(n7325), .A2(n7327), .ZN(n11807) );
  NAND2_X1 U9455 ( .A1(n11650), .A2(n7326), .ZN(n7325) );
  NAND4_X1 U9456 ( .A1(n9745), .A2(n6544), .A3(n13332), .A4(n7331), .ZN(n7330)
         );
  NAND2_X1 U9457 ( .A1(n14636), .A2(n7334), .ZN(n7333) );
  NAND2_X1 U9458 ( .A1(n7333), .A2(n7335), .ZN(n11422) );
  INV_X1 U9459 ( .A(n7342), .ZN(n7338) );
  NAND2_X1 U9460 ( .A1(n7339), .A2(n7340), .ZN(n14023) );
  NAND2_X1 U9461 ( .A1(n11817), .A2(n7348), .ZN(n7347) );
  NAND2_X1 U9462 ( .A1(n7354), .A2(n7353), .ZN(n13998) );
  NAND3_X1 U9463 ( .A1(n6479), .A2(n9994), .A3(n9998), .ZN(n7354) );
  NAND2_X1 U9464 ( .A1(n9995), .A2(n9994), .ZN(n14018) );
  NAND2_X1 U9465 ( .A1(n14651), .A2(n9963), .ZN(n7362) );
  NAND3_X1 U9466 ( .A1(n7357), .A2(n7356), .A3(n6596), .ZN(n14638) );
  NAND3_X1 U9467 ( .A1(n6552), .A2(n9903), .A3(n7360), .ZN(n7356) );
  NAND3_X1 U9468 ( .A1(n14651), .A2(n7358), .A3(n6552), .ZN(n7357) );
  OR2_X2 U9469 ( .A1(n6527), .A2(n7369), .ZN(n7368) );
  NAND2_X1 U9470 ( .A1(n7491), .A2(n8025), .ZN(n8037) );
  NAND2_X1 U9471 ( .A1(n11971), .A2(n9920), .ZN(n14073) );
  OAI21_X1 U9472 ( .B1(n6470), .B2(n7380), .A(n7377), .ZN(n9911) );
  OAI21_X2 U9473 ( .B1(n14082), .B2(n9990), .A(n9989), .ZN(n14050) );
  NAND2_X1 U9474 ( .A1(n8279), .A2(n7381), .ZN(n13635) );
  AOI21_X1 U9475 ( .B1(n8234), .B2(n7383), .A(n7382), .ZN(n7381) );
  NAND2_X1 U9476 ( .A1(n8234), .A2(n8233), .ZN(n8268) );
  INV_X1 U9477 ( .A(n8273), .ZN(n7386) );
  NAND3_X1 U9478 ( .A1(n7393), .A2(SI_18_), .A3(n7392), .ZN(n7986) );
  NAND2_X1 U9479 ( .A1(n7949), .A2(n7986), .ZN(n7953) );
  NOR2_X2 U9480 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n7400) );
  NOR2_X2 U9481 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n7402) );
  NOR2_X2 U9482 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n7404) );
  NOR2_X2 U9483 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n7405) );
  NAND2_X1 U9484 ( .A1(n7406), .A2(n6613), .ZN(n9560) );
  INV_X1 U9485 ( .A(n9554), .ZN(n7407) );
  NAND2_X1 U9486 ( .A1(n9493), .A2(n7415), .ZN(n7414) );
  AOI21_X1 U9487 ( .B1(n9512), .B2(n9511), .A(n9509), .ZN(n9510) );
  NAND2_X1 U9488 ( .A1(n9634), .A2(n9633), .ZN(n7420) );
  NAND3_X1 U9489 ( .A1(n9525), .A2(n6614), .A3(n9524), .ZN(n7424) );
  INV_X1 U9490 ( .A(n9652), .ZN(n7428) );
  NAND3_X1 U9491 ( .A1(n9616), .A2(n9615), .A3(n6600), .ZN(n7431) );
  AOI21_X1 U9492 ( .B1(n13348), .B2(n7119), .A(n7453), .ZN(n13330) );
  NAND2_X1 U9493 ( .A1(n13348), .A2(n7435), .ZN(n7434) );
  NAND4_X1 U9494 ( .A1(n7442), .A2(n7439), .A3(n14961), .A4(n7437), .ZN(n7452)
         );
  NAND2_X1 U9495 ( .A1(n13348), .A2(n7438), .ZN(n7437) );
  NAND2_X1 U9496 ( .A1(n7441), .A2(n7440), .ZN(n7439) );
  INV_X1 U9497 ( .A(n13348), .ZN(n7440) );
  NAND2_X1 U9498 ( .A1(n7452), .A2(n7451), .ZN(n13620) );
  AND2_X1 U9499 ( .A1(n13547), .A2(n13243), .ZN(n7453) );
  NAND2_X1 U9500 ( .A1(n7456), .A2(n7457), .ZN(n11271) );
  OR2_X1 U9501 ( .A1(n13453), .A2(n9462), .ZN(n7461) );
  NAND2_X1 U9502 ( .A1(n9464), .A2(n7464), .ZN(n7463) );
  NAND2_X1 U9503 ( .A1(n13395), .A2(n7470), .ZN(n7467) );
  NAND2_X1 U9504 ( .A1(n7467), .A2(n7468), .ZN(n13361) );
  INV_X1 U9505 ( .A(n13558), .ZN(n7474) );
  NAND2_X1 U9506 ( .A1(n11701), .A2(n7480), .ZN(n7479) );
  OR2_X1 U9507 ( .A1(n9671), .A2(n10378), .ZN(n9011) );
  NAND2_X1 U9508 ( .A1(n8920), .A2(n8919), .ZN(n8923) );
  AND3_X1 U9509 ( .A1(n9874), .A2(n10893), .A3(n9875), .ZN(n9862) );
  CLKBUF_X1 U9510 ( .A(n11923), .Z(n11926) );
  INV_X1 U9511 ( .A(n12469), .ZN(n8902) );
  CLKBUF_X1 U9512 ( .A(n9761), .Z(n10670) );
  NAND2_X1 U9513 ( .A1(n8898), .A2(n10881), .ZN(n9758) );
  OAI211_X2 U9514 ( .C1(n9874), .C2(n12195), .A(n9758), .B(n9757), .ZN(n9760)
         );
  NAND2_X1 U9515 ( .A1(n8809), .A2(n8808), .ZN(n12783) );
  NAND2_X1 U9516 ( .A1(n9887), .A2(n15175), .ZN(n8955) );
  INV_X1 U9517 ( .A(n8353), .ZN(n8472) );
  NAND4_X2 U9518 ( .A1(n7607), .A2(n7606), .A3(n7605), .A4(n7604), .ZN(n13841)
         );
  OR2_X1 U9519 ( .A1(n7624), .A2(n10135), .ZN(n7606) );
  INV_X1 U9520 ( .A(n11194), .ZN(n12175) );
  INV_X1 U9521 ( .A(n8355), .ZN(n8354) );
  CLKBUF_X1 U9522 ( .A(n10489), .Z(n14780) );
  NAND2_X1 U9523 ( .A1(n7623), .A2(n7622), .ZN(n7650) );
  INV_X1 U9524 ( .A(n8422), .ZN(n8424) );
  CLKBUF_X1 U9525 ( .A(n13192), .Z(n13194) );
  OAI21_X1 U9526 ( .B1(n9130), .B2(n9367), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n9368) );
  NAND2_X1 U9527 ( .A1(n9962), .A2(n9961), .ZN(n14658) );
  NAND2_X2 U9528 ( .A1(n8987), .A2(n8986), .ZN(n9130) );
  NAND2_X1 U9529 ( .A1(n10578), .A2(n10579), .ZN(n10638) );
  NAND2_X1 U9530 ( .A1(n9718), .A2(n9717), .ZN(n9719) );
  INV_X1 U9531 ( .A(n14679), .ZN(n14699) );
  NAND2_X1 U9532 ( .A1(n14679), .A2(n7988), .ZN(n11235) );
  AOI21_X1 U9533 ( .B1(n9374), .B2(P2_IR_REG_31__SCAN_IN), .A(n7320), .ZN(
        n9375) );
  INV_X1 U9534 ( .A(n9520), .ZN(n9523) );
  NAND2_X1 U9535 ( .A1(n9390), .A2(n6478), .ZN(n13654) );
  OR2_X4 U9536 ( .A1(n10453), .A2(n10456), .ZN(n12453) );
  NAND4_X2 U9537 ( .A1(n9035), .A2(n9034), .A3(n9033), .A4(n9032), .ZN(n13268)
         );
  NAND4_X2 U9538 ( .A1(n9011), .A2(n9010), .A3(n9009), .A4(n9008), .ZN(n13270)
         );
  NAND2_X1 U9539 ( .A1(n14095), .A2(n14618), .ZN(n14102) );
  OAI21_X2 U9540 ( .B1(n9608), .B2(n9607), .A(n9606), .ZN(n9614) );
  XNOR2_X1 U9541 ( .A(n12480), .B(n12024), .ZN(n12015) );
  AND3_X2 U9542 ( .A1(n10897), .A2(n9885), .A3(n9884), .ZN(n15183) );
  INV_X1 U9543 ( .A(n15183), .ZN(n9886) );
  OR2_X1 U9544 ( .A1(n9888), .A2(n13003), .ZN(n7482) );
  INV_X1 U9545 ( .A(n14052), .ZN(n14069) );
  NOR2_X1 U9546 ( .A1(n14070), .A2(n14172), .ZN(n14052) );
  INV_X1 U9547 ( .A(n9919), .ZN(n11974) );
  OR2_X1 U9548 ( .A1(n10079), .A2(n13868), .ZN(n7484) );
  NAND2_X1 U9549 ( .A1(n8181), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n7485) );
  INV_X1 U9550 ( .A(n11828), .ZN(n8324) );
  NOR2_X1 U9551 ( .A1(n9810), .A2(n12591), .ZN(n7486) );
  AND2_X1 U9552 ( .A1(n9809), .A2(n12660), .ZN(n7487) );
  NAND2_X1 U9553 ( .A1(n7945), .A2(n7944), .ZN(n7488) );
  OR2_X1 U9554 ( .A1(n9237), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n7492) );
  AND2_X1 U9555 ( .A1(n9702), .A2(n9701), .ZN(n7493) );
  INV_X1 U9556 ( .A(n12287), .ZN(n8884) );
  INV_X1 U9557 ( .A(n12662), .ZN(n12926) );
  AND4_X1 U9558 ( .A1(n7512), .A2(n7511), .A3(n7510), .A4(n7509), .ZN(n7494)
         );
  INV_X1 U9559 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n14199) );
  OR2_X1 U9560 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10906), .ZN(n7495) );
  INV_X1 U9561 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8601) );
  NAND2_X1 U9562 ( .A1(n8240), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7496) );
  INV_X1 U9563 ( .A(P3_U3897), .ZN(n12658) );
  INV_X2 U9564 ( .A(n8240), .ZN(n7624) );
  INV_X1 U9565 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8907) );
  AND2_X1 U9566 ( .A1(n15110), .A2(n15169), .ZN(n12988) );
  INV_X1 U9567 ( .A(n9907), .ZN(n11107) );
  INV_X1 U9568 ( .A(n10403), .ZN(n10476) );
  NAND2_X1 U9569 ( .A1(n7936), .A2(SI_16_), .ZN(n7946) );
  OR4_X1 U9570 ( .A1(n14924), .A2(n14420), .A3(n13650), .A4(n10208), .ZN(n7497) );
  OR2_X1 U9571 ( .A1(n13540), .A2(n13528), .ZN(n7498) );
  XNOR2_X1 U9572 ( .A(n14096), .B(n13820), .ZN(n12481) );
  INV_X1 U9573 ( .A(n12481), .ZN(n12476) );
  NOR2_X1 U9574 ( .A1(n8317), .A2(n8316), .ZN(n7499) );
  NAND2_X2 U9575 ( .A1(n14673), .A2(n12490), .ZN(n14665) );
  INV_X1 U9576 ( .A(n9897), .ZN(n7597) );
  NAND2_X1 U9577 ( .A1(n8284), .A2(n7597), .ZN(n7598) );
  MUX2_X1 U9578 ( .A(n7621), .B(n7620), .S(n14676), .Z(n7622) );
  INV_X1 U9579 ( .A(n9521), .ZN(n9522) );
  AND2_X1 U9580 ( .A1(n8004), .A2(n8003), .ZN(n8005) );
  NOR2_X1 U9581 ( .A1(n9683), .A2(n9696), .ZN(n9697) );
  NOR2_X1 U9582 ( .A1(n7898), .A2(n15263), .ZN(n7892) );
  AND2_X1 U9583 ( .A1(n10820), .A2(n14976), .ZN(n10821) );
  NAND2_X1 U9584 ( .A1(n11836), .A2(n11834), .ZN(n8649) );
  INV_X1 U9585 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n7500) );
  OR2_X1 U9586 ( .A1(n9799), .A2(n12547), .ZN(n9806) );
  INV_X1 U9587 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8349) );
  INV_X1 U9588 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n15282) );
  INV_X1 U9589 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n11927) );
  NAND2_X1 U9590 ( .A1(n8500), .A2(n8499), .ZN(n15094) );
  INV_X1 U9591 ( .A(n14783), .ZN(n10486) );
  AND2_X1 U9592 ( .A1(n13558), .A2(n13196), .ZN(n9319) );
  INV_X1 U9593 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9121) );
  INV_X1 U9594 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9069) );
  INV_X1 U9595 ( .A(n13591), .ZN(n9431) );
  NAND2_X1 U9596 ( .A1(n11591), .A2(n11592), .ZN(n11593) );
  AND2_X1 U9597 ( .A1(n11506), .A2(n11507), .ZN(n11505) );
  INV_X1 U9598 ( .A(n8077), .ZN(n8076) );
  INV_X1 U9599 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7806) );
  NOR2_X1 U9600 ( .A1(n8011), .A2(n8010), .ZN(n8044) );
  AND2_X1 U9601 ( .A1(n7925), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7959) );
  INV_X1 U9602 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7652) );
  INV_X1 U9603 ( .A(n14062), .ZN(n10006) );
  INV_X1 U9604 ( .A(n11589), .ZN(n10005) );
  INV_X1 U9605 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n7513) );
  INV_X1 U9606 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n8385) );
  NOR2_X1 U9607 ( .A1(n14263), .A2(n14262), .ZN(n14239) );
  INV_X1 U9608 ( .A(n11579), .ZN(n9791) );
  INV_X1 U9609 ( .A(n10785), .ZN(n9764) );
  AND2_X1 U9610 ( .A1(n9774), .A2(n15091), .ZN(n9775) );
  INV_X1 U9611 ( .A(n12656), .ZN(n9831) );
  INV_X1 U9612 ( .A(n12211), .ZN(n9756) );
  OR2_X1 U9613 ( .A1(n8766), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8774) );
  NAND2_X1 U9614 ( .A1(n8735), .A2(n15282), .ZN(n8737) );
  NAND2_X2 U9615 ( .A1(n8472), .A2(n8354), .ZN(n8510) );
  OAI21_X1 U9616 ( .B1(n12769), .B2(n8893), .A(n12201), .ZN(n12132) );
  NAND2_X1 U9617 ( .A1(n12772), .A2(n12771), .ZN(n12770) );
  NOR2_X1 U9618 ( .A1(n8659), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8672) );
  INV_X1 U9619 ( .A(n11326), .ZN(n12252) );
  OR2_X1 U9620 ( .A1(n8935), .A2(n8934), .ZN(n9875) );
  NAND2_X1 U9621 ( .A1(n11538), .A2(n12171), .ZN(n11537) );
  INV_X2 U9622 ( .A(n12364), .ZN(n12370) );
  OAI21_X1 U9623 ( .B1(n12137), .B2(n12136), .A(n12135), .ZN(n12155) );
  INV_X1 U9624 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8408) );
  NAND2_X1 U9625 ( .A1(n8653), .A2(n8384), .ZN(n8387) );
  INV_X1 U9626 ( .A(n11348), .ZN(n11345) );
  NAND2_X1 U9627 ( .A1(n13088), .A2(n13087), .ZN(n13089) );
  OR2_X1 U9628 ( .A1(n9311), .A2(n13168), .ZN(n9322) );
  AND2_X1 U9629 ( .A1(n8959), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9242) );
  OR2_X1 U9630 ( .A1(n9221), .A2(n9220), .ZN(n9223) );
  NAND2_X1 U9631 ( .A1(n9242), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9262) );
  INV_X1 U9632 ( .A(n13611), .ZN(n9430) );
  NAND2_X1 U9633 ( .A1(n13242), .A2(n13231), .ZN(n9385) );
  INV_X1 U9634 ( .A(n11702), .ZN(n14444) );
  INV_X1 U9635 ( .A(n11747), .ZN(n11748) );
  OR2_X1 U9636 ( .A1(n8179), .A2(n13663), .ZN(n8198) );
  OR2_X1 U9637 ( .A1(n8107), .A2(n13754), .ZN(n8130) );
  NAND2_X1 U9638 ( .A1(n7959), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n7971) );
  OR2_X1 U9639 ( .A1(n7807), .A2(n7806), .ZN(n7829) );
  OR2_X1 U9640 ( .A1(n8130), .A2(n8129), .ZN(n8160) );
  NAND2_X1 U9641 ( .A1(n8044), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8061) );
  NAND2_X1 U9642 ( .A1(n9967), .A2(n9966), .ZN(n11138) );
  NAND2_X1 U9643 ( .A1(n14052), .A2(n10006), .ZN(n14058) );
  OR2_X1 U9644 ( .A1(n7839), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n7840) );
  INV_X1 U9645 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n7502) );
  OR2_X1 U9646 ( .A1(n14233), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n14232) );
  NOR2_X1 U9647 ( .A1(n14259), .A2(n14258), .ZN(n14245) );
  NAND2_X1 U9648 ( .A1(n8602), .A2(n8601), .ZN(n8618) );
  AND2_X1 U9649 ( .A1(n9847), .A2(n9845), .ZN(n12581) );
  NAND2_X1 U9650 ( .A1(n8786), .A2(n12607), .ZN(n8788) );
  INV_X1 U9651 ( .A(n15102), .ZN(n12212) );
  INV_X1 U9652 ( .A(n12552), .ZN(n12632) );
  OR2_X1 U9653 ( .A1(n9861), .A2(n10722), .ZN(n9854) );
  INV_X1 U9654 ( .A(n12145), .ZN(n8831) );
  INV_X1 U9655 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n14220) );
  AND2_X1 U9656 ( .A1(n10737), .A2(n10735), .ZN(n10746) );
  NAND2_X1 U9657 ( .A1(n11406), .A2(n12246), .ZN(n11405) );
  INV_X1 U9658 ( .A(n15104), .ZN(n12925) );
  INV_X1 U9659 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8352) );
  AND2_X1 U9660 ( .A1(n8400), .A2(n8399), .ZN(n8458) );
  INV_X1 U9661 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8612) );
  AND2_X1 U9662 ( .A1(n8371), .A2(n8370), .ZN(n8544) );
  AND2_X1 U9663 ( .A1(n8363), .A2(n8362), .ZN(n8501) );
  AND2_X1 U9664 ( .A1(n9151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n9168) );
  OR3_X1 U9665 ( .A1(n9262), .A2(n13206), .A3(n13154), .ZN(n9278) );
  NAND2_X1 U9666 ( .A1(n9477), .A2(n10214), .ZN(n10405) );
  NAND2_X1 U9667 ( .A1(n11772), .A2(n9679), .ZN(n9276) );
  OR2_X1 U9668 ( .A1(n14815), .A2(n14814), .ZN(n14817) );
  AND2_X1 U9669 ( .A1(n10108), .A2(n13644), .ZN(n10116) );
  INV_X1 U9670 ( .A(n9707), .ZN(n13319) );
  INV_X1 U9671 ( .A(n13469), .ZN(n13490) );
  AND2_X1 U9672 ( .A1(n10257), .A2(n9421), .ZN(n10206) );
  OR2_X1 U9673 ( .A1(n9379), .A2(n10219), .ZN(n14422) );
  AND2_X1 U9674 ( .A1(n9672), .A2(n11773), .ZN(n10354) );
  INV_X1 U9675 ( .A(n9738), .ZN(n13500) );
  INV_X1 U9676 ( .A(n11353), .ZN(n14464) );
  INV_X1 U9677 ( .A(n13654), .ZN(n9404) );
  INV_X1 U9678 ( .A(n9394), .ZN(n9388) );
  NAND2_X1 U9679 ( .A1(n11999), .A2(n12000), .ZN(n12056) );
  NAND2_X1 U9680 ( .A1(n11746), .A2(n11748), .ZN(n11749) );
  AND2_X1 U9681 ( .A1(n13681), .A2(n13679), .ZN(n12083) );
  XNOR2_X1 U9682 ( .A(n10577), .B(n6519), .ZN(n10579) );
  INV_X1 U9683 ( .A(n13830), .ZN(n13741) );
  AND2_X1 U9684 ( .A1(n11678), .A2(n11675), .ZN(n11676) );
  OR2_X1 U9685 ( .A1(n13778), .A2(n14053), .ZN(n13808) );
  AND2_X1 U9686 ( .A1(n8198), .A2(n8180), .ZN(n13945) );
  OR2_X1 U9687 ( .A1(n7994), .A2(n7993), .ZN(n8011) );
  INV_X1 U9688 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14222) );
  OR2_X1 U9689 ( .A1(n10147), .A2(n10148), .ZN(n10174) );
  INV_X1 U9690 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n13806) );
  NAND2_X1 U9691 ( .A1(n13956), .A2(n14482), .ZN(n12012) );
  INV_X1 U9692 ( .A(n13992), .ZN(n13978) );
  AND2_X1 U9693 ( .A1(n8335), .A2(n13859), .ZN(n14482) );
  INV_X1 U9694 ( .A(n14755), .ZN(n14723) );
  INV_X1 U9695 ( .A(n9971), .ZN(n14637) );
  INV_X1 U9696 ( .A(n9899), .ZN(n14669) );
  OR2_X1 U9697 ( .A1(n10464), .A2(n13859), .ZN(n14055) );
  AOI21_X1 U9698 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(n14242), .A(n14241), .ZN(
        n14300) );
  XOR2_X1 U9699 ( .A(n12659), .B(n9817), .Z(n12563) );
  INV_X1 U9700 ( .A(n11030), .ZN(n12384) );
  OR2_X1 U9701 ( .A1(n8510), .A2(n12791), .ZN(n8822) );
  NAND2_X1 U9702 ( .A1(n8936), .A2(n8939), .ZN(n9892) );
  INV_X1 U9703 ( .A(n15036), .ZN(n15069) );
  INV_X1 U9704 ( .A(n12922), .ZN(n15106) );
  INV_X1 U9705 ( .A(n12902), .ZN(n12935) );
  AND3_X1 U9706 ( .A1(n8581), .A2(n8580), .A3(n8579), .ZN(n15149) );
  OR2_X1 U9707 ( .A1(n9855), .A2(n15111), .ZN(n15112) );
  NOR2_X1 U9708 ( .A1(n9877), .A2(n9876), .ZN(n10897) );
  INV_X1 U9709 ( .A(n12988), .ZN(n14415) );
  OR2_X1 U9710 ( .A1(n9866), .A2(n8948), .ZN(n8949) );
  INV_X1 U9711 ( .A(n15168), .ZN(n15150) );
  INV_X1 U9712 ( .A(n13063), .ZN(n10090) );
  INV_X1 U9713 ( .A(n11824), .ZN(n9750) );
  OR2_X1 U9714 ( .A1(n10109), .A2(n10115), .ZN(n14862) );
  INV_X1 U9715 ( .A(n14862), .ZN(n14878) );
  AND2_X1 U9716 ( .A1(n10116), .A2(n10115), .ZN(n14875) );
  INV_X1 U9717 ( .A(n10403), .ZN(n13523) );
  INV_X1 U9718 ( .A(n9736), .ZN(n11708) );
  INV_X1 U9719 ( .A(n13472), .ZN(n14890) );
  NAND2_X1 U9720 ( .A1(n14927), .A2(n9422), .ZN(n13518) );
  INV_X1 U9721 ( .A(n13528), .ZN(n14900) );
  INV_X1 U9722 ( .A(n14945), .ZN(n14958) );
  AND2_X1 U9723 ( .A1(n10257), .A2(n10256), .ZN(n10356) );
  OR2_X1 U9724 ( .A1(n9471), .A2(n14950), .ZN(n14961) );
  AND2_X1 U9725 ( .A1(n9402), .A2(n9401), .ZN(n10204) );
  NAND2_X1 U9726 ( .A1(n9388), .A2(n9387), .ZN(n9396) );
  AND2_X1 U9727 ( .A1(n9177), .A2(n9201), .ZN(n14866) );
  AND2_X1 U9728 ( .A1(n10466), .A2(n11233), .ZN(n13769) );
  AND2_X1 U9729 ( .A1(n13769), .A2(n14631), .ZN(n13810) );
  AND2_X1 U9730 ( .A1(n8068), .A2(n8067), .ZN(n13691) );
  OR2_X1 U9731 ( .A1(n10388), .A2(n10387), .ZN(n10434) );
  INV_X1 U9732 ( .A(n13920), .ZN(n14606) );
  INV_X1 U9733 ( .A(n9916), .ZN(n11870) );
  OR2_X1 U9734 ( .A1(n11235), .A2(n10463), .ZN(n14673) );
  AND2_X1 U9735 ( .A1(n9951), .A2(n10042), .ZN(n11254) );
  INV_X1 U9736 ( .A(n14618), .ZN(n14690) );
  INV_X1 U9737 ( .A(n14691), .ZN(n14759) );
  INV_X1 U9738 ( .A(n11254), .ZN(n11236) );
  NAND2_X1 U9739 ( .A1(n14231), .A2(n14230), .ZN(n14284) );
  AND2_X1 U9740 ( .A1(n10737), .A2(n10736), .ZN(n15068) );
  INV_X1 U9741 ( .A(n10675), .ZN(n12608) );
  INV_X1 U9742 ( .A(n12629), .ZN(n12645) );
  INV_X1 U9743 ( .A(n11834), .ZN(n12666) );
  INV_X1 U9744 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n15009) );
  INV_X1 U9745 ( .A(n15082), .ZN(n15063) );
  NOR2_X1 U9746 ( .A1(n8951), .A2(n8953), .ZN(n8954) );
  AND2_X1 U9747 ( .A1(n8950), .A2(n8949), .ZN(n15173) );
  NAND2_X1 U9748 ( .A1(n15175), .A2(n15150), .ZN(n13059) );
  NOR2_X1 U9749 ( .A1(n8914), .A2(n10090), .ZN(n10548) );
  INV_X1 U9750 ( .A(SI_18_), .ZN(n15252) );
  INV_X1 U9751 ( .A(SI_12_), .ZN(n15312) );
  NAND2_X1 U9752 ( .A1(n10494), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14789) );
  AND2_X1 U9753 ( .A1(n10207), .A2(n13518), .ZN(n13210) );
  INV_X1 U9754 ( .A(n14873), .ZN(n14822) );
  INV_X1 U9755 ( .A(n14919), .ZN(n13531) );
  NAND2_X1 U9756 ( .A1(n14919), .A2(n9473), .ZN(n13528) );
  NAND2_X1 U9757 ( .A1(n10356), .A2(n10355), .ZN(n14969) );
  NAND2_X1 U9758 ( .A1(n10258), .A2(n10356), .ZN(n14962) );
  OR2_X1 U9759 ( .A1(n14924), .A2(n14920), .ZN(n14921) );
  AND2_X1 U9760 ( .A1(n10200), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14927) );
  INV_X1 U9761 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10688) );
  INV_X1 U9762 ( .A(n14151), .ZN(n14029) );
  INV_X1 U9763 ( .A(n13795), .ZN(n13817) );
  NAND2_X1 U9764 ( .A1(n8166), .A2(n8165), .ZN(n13822) );
  INV_X1 U9765 ( .A(n14591), .ZN(n14611) );
  INV_X1 U9766 ( .A(n14587), .ZN(n14615) );
  INV_X1 U9767 ( .A(n14665), .ZN(n14087) );
  INV_X1 U9768 ( .A(n14776), .ZN(n14773) );
  OR2_X1 U9769 ( .A1(n14181), .A2(n14180), .ZN(n14198) );
  INV_X1 U9770 ( .A(n14761), .ZN(n14760) );
  AND2_X2 U9771 ( .A1(n11255), .A2(n11236), .ZN(n14761) );
  AND2_X1 U9772 ( .A1(n8326), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10472) );
  INV_X1 U9773 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10913) );
  INV_X1 U9774 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10517) );
  AND2_X1 U9775 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10102), .ZN(P2_U3947) );
  NAND2_X1 U9776 ( .A1(n9474), .A2(n7498), .ZN(P2_U3236) );
  NOR2_X1 U9777 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n7507) );
  NOR2_X1 U9778 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n7506) );
  NOR2_X1 U9779 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n7505) );
  NOR3_X1 U9780 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .A3(
        P1_IR_REG_23__SCAN_IN), .ZN(n7512) );
  NOR2_X1 U9781 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n7511) );
  NOR2_X1 U9782 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n7510) );
  NOR2_X1 U9783 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n7509) );
  NOR2_X1 U9784 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n7515) );
  NAND2_X1 U9785 ( .A1(n7532), .A2(n7515), .ZN(n14200) );
  XNOR2_X2 U9786 ( .A(n7516), .B(P1_IR_REG_30__SCAN_IN), .ZN(n7520) );
  INV_X1 U9787 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n7533) );
  NAND2_X1 U9788 ( .A1(n7532), .A2(n7533), .ZN(n7517) );
  XNOR2_X2 U9789 ( .A(n7518), .B(P1_IR_REG_29__SCAN_IN), .ZN(n7519) );
  AND2_X2 U9790 ( .A1(n7520), .A2(n7519), .ZN(n8181) );
  INV_X1 U9791 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11151) );
  OR2_X1 U9792 ( .A1(n7603), .A2(n11151), .ZN(n7525) );
  INV_X2 U9793 ( .A(n7520), .ZN(n12527) );
  AND2_X4 U9794 ( .A1(n7519), .A2(n12527), .ZN(n8240) );
  INV_X2 U9795 ( .A(n7519), .ZN(n7522) );
  NAND2_X4 U9796 ( .A1(n7522), .A2(n7521), .ZN(n8246) );
  INV_X1 U9797 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n11152) );
  OR2_X1 U9798 ( .A1(n8246), .A2(n11152), .ZN(n7524) );
  NAND2_X4 U9799 ( .A1(n12527), .A2(n7522), .ZN(n8248) );
  NAND2_X1 U9800 ( .A1(n7693), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n7523) );
  INV_X1 U9801 ( .A(SI_0_), .ZN(n10034) );
  NOR2_X1 U9802 ( .A1(n6720), .A2(n10034), .ZN(n7531) );
  INV_X1 U9803 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8491) );
  XNOR2_X1 U9804 ( .A(n7531), .B(n8491), .ZN(n14217) );
  OR2_X2 U9805 ( .A1(n7532), .A2(n14199), .ZN(n7534) );
  XNOR2_X2 U9806 ( .A(n7534), .B(n7533), .ZN(n8325) );
  MUX2_X1 U9807 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14217), .S(n10079), .Z(n14694)
         );
  XNOR2_X2 U9808 ( .A(n7537), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9936) );
  NAND2_X1 U9809 ( .A1(n8299), .A2(n10453), .ZN(n7541) );
  INV_X1 U9810 ( .A(n14694), .ZN(n11153) );
  NAND2_X1 U9811 ( .A1(n13843), .A2(n11153), .ZN(n8298) );
  NAND2_X1 U9812 ( .A1(n7541), .A2(n8298), .ZN(n7572) );
  INV_X1 U9813 ( .A(n7542), .ZN(n7543) );
  NOR2_X1 U9814 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n7550) );
  INV_X1 U9815 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n7549) );
  INV_X1 U9816 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n7548) );
  NAND4_X1 U9817 ( .A1(n7550), .A2(n7549), .A3(n7548), .A4(n7547), .ZN(n7551)
         );
  NAND2_X1 U9818 ( .A1(n8333), .A2(n14215), .ZN(n10002) );
  NAND2_X1 U9819 ( .A1(n7988), .A2(n10010), .ZN(n11237) );
  NAND2_X1 U9820 ( .A1(n10002), .A2(n11237), .ZN(n8252) );
  MUX2_X1 U9821 ( .A(n11421), .B(n9936), .S(n8252), .Z(n7552) );
  INV_X1 U9822 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10154) );
  OR2_X1 U9823 ( .A1(n8246), .A2(n10154), .ZN(n7556) );
  INV_X1 U9824 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7553) );
  OR2_X1 U9825 ( .A1(n6491), .A2(n7553), .ZN(n7555) );
  NAND2_X1 U9826 ( .A1(n8240), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7554) );
  INV_X2 U9827 ( .A(n7573), .ZN(n11150) );
  NAND2_X1 U9828 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n7557) );
  MUX2_X1 U9829 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7557), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n7559) );
  NAND2_X1 U9830 ( .A1(n7559), .A2(n6487), .ZN(n13847) );
  INV_X1 U9831 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10021) );
  OR2_X1 U9832 ( .A1(n7644), .A2(n10021), .ZN(n7571) );
  INV_X1 U9833 ( .A(n8119), .ZN(n10022) );
  NAND2_X1 U9834 ( .A1(n7612), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7560) );
  NAND2_X1 U9835 ( .A1(n7561), .A2(SI_1_), .ZN(n7582) );
  NAND2_X1 U9836 ( .A1(n7563), .A2(n7562), .ZN(n7564) );
  NOR2_X1 U9837 ( .A1(n7565), .A2(n10034), .ZN(n7566) );
  INV_X1 U9838 ( .A(n7566), .ZN(n7567) );
  NAND2_X1 U9839 ( .A1(n7568), .A2(n7567), .ZN(n7569) );
  NAND2_X1 U9840 ( .A1(n7583), .A2(n7569), .ZN(n10023) );
  OR2_X1 U9841 ( .A1(n7670), .A2(n10023), .ZN(n7570) );
  NAND2_X1 U9842 ( .A1(n11150), .A2(n6493), .ZN(n9895) );
  NAND3_X1 U9843 ( .A1(n7572), .A2(n8284), .A3(n9895), .ZN(n7596) );
  OAI21_X1 U9844 ( .B1(n7573), .B2(n7552), .A(n6493), .ZN(n7576) );
  NAND2_X1 U9845 ( .A1(n7573), .A2(n7552), .ZN(n7574) );
  INV_X1 U9846 ( .A(n11019), .ZN(n14698) );
  NAND2_X1 U9847 ( .A1(n7574), .A2(n14698), .ZN(n7575) );
  NAND2_X1 U9848 ( .A1(n7576), .A2(n7575), .ZN(n7595) );
  NAND2_X1 U9849 ( .A1(n8240), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7581) );
  INV_X1 U9850 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10645) );
  OR2_X1 U9851 ( .A1(n7603), .A2(n10645), .ZN(n7580) );
  INV_X1 U9852 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7577) );
  OR2_X1 U9853 ( .A1(n8248), .A2(n7577), .ZN(n7579) );
  INV_X1 U9854 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10156) );
  OR2_X1 U9855 ( .A1(n8246), .A2(n10156), .ZN(n7578) );
  NAND2_X1 U9856 ( .A1(n7633), .A2(SI_2_), .ZN(n7610) );
  OAI21_X1 U9857 ( .B1(n7633), .B2(SI_2_), .A(n7610), .ZN(n7585) );
  NAND2_X1 U9858 ( .A1(n7585), .A2(n7630), .ZN(n7586) );
  NAND2_X1 U9859 ( .A1(n8282), .A2(n10017), .ZN(n7592) );
  OR2_X1 U9860 ( .A1(n6492), .A2(n10018), .ZN(n7590) );
  NAND2_X1 U9861 ( .A1(n6487), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7587) );
  MUX2_X1 U9862 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7587), .S(
        P1_IR_REG_2__SCAN_IN), .Z(n7589) );
  NAND2_X1 U9863 ( .A1(n7589), .A2(n7588), .ZN(n13868) );
  AND2_X1 U9864 ( .A1(n7590), .A2(n7484), .ZN(n7591) );
  NAND2_X2 U9865 ( .A1(n7592), .A2(n7591), .ZN(n11119) );
  INV_X2 U9866 ( .A(n11119), .ZN(n14705) );
  NAND2_X1 U9867 ( .A1(n13842), .A2(n14705), .ZN(n7599) );
  NAND2_X1 U9868 ( .A1(n10641), .A2(n11119), .ZN(n9897) );
  AND2_X1 U9869 ( .A1(n7599), .A2(n9897), .ZN(n7594) );
  NAND2_X1 U9870 ( .A1(n7573), .A2(n14698), .ZN(n9894) );
  NAND3_X1 U9871 ( .A1(n9893), .A2(n7750), .A3(n9894), .ZN(n7593) );
  NAND4_X1 U9872 ( .A1(n7596), .A2(n7595), .A3(n7594), .A4(n7593), .ZN(n7602)
         );
  OAI21_X1 U9873 ( .B1(n7599), .B2(n8284), .A(n7598), .ZN(n7600) );
  INV_X1 U9874 ( .A(n7600), .ZN(n7601) );
  NAND2_X1 U9875 ( .A1(n7602), .A2(n7601), .ZN(n7619) );
  NAND2_X1 U9876 ( .A1(n7693), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n7607) );
  INV_X1 U9877 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10135) );
  INV_X1 U9878 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n14674) );
  OR2_X1 U9879 ( .A1(n8246), .A2(n14674), .ZN(n7605) );
  OR2_X1 U9880 ( .A1(n7603), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7604) );
  NAND2_X1 U9881 ( .A1(n7588), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7609) );
  XNOR2_X1 U9882 ( .A(n7609), .B(n7608), .ZN(n13879) );
  NAND2_X1 U9883 ( .A1(n7613), .A2(SI_3_), .ZN(n7634) );
  INV_X1 U9884 ( .A(n7613), .ZN(n7614) );
  INV_X1 U9885 ( .A(SI_3_), .ZN(n10026) );
  NAND2_X1 U9886 ( .A1(n7614), .A2(n10026), .ZN(n7615) );
  NAND2_X1 U9887 ( .A1(n10038), .A2(n8282), .ZN(n7618) );
  OR2_X1 U9888 ( .A1(n6492), .A2(n10039), .ZN(n7617) );
  OAI211_X1 U9889 ( .C1(n10079), .C2(n13879), .A(n7618), .B(n7617), .ZN(n14676) );
  XNOR2_X1 U9890 ( .A(n13841), .B(n14676), .ZN(n9899) );
  NAND2_X1 U9891 ( .A1(n7619), .A2(n9899), .ZN(n7623) );
  NAND2_X1 U9892 ( .A1(n13841), .A2(n7750), .ZN(n7621) );
  INV_X1 U9893 ( .A(n13841), .ZN(n9960) );
  NAND2_X1 U9894 ( .A1(n9960), .A2(n7552), .ZN(n7620) );
  INV_X2 U9895 ( .A(n8246), .ZN(n7651) );
  NAND2_X1 U9896 ( .A1(n7651), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7629) );
  INV_X1 U9897 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10136) );
  OR2_X1 U9898 ( .A1(n7624), .A2(n10136), .ZN(n7628) );
  NAND2_X1 U9899 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n7653) );
  OAI21_X1 U9900 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n7653), .ZN(n14656) );
  OR2_X1 U9901 ( .A1(n7603), .A2(n14656), .ZN(n7627) );
  INV_X1 U9902 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7625) );
  OR2_X1 U9903 ( .A1(n8248), .A2(n7625), .ZN(n7626) );
  INV_X1 U9904 ( .A(SI_2_), .ZN(n10029) );
  INV_X1 U9905 ( .A(n7635), .ZN(n7636) );
  NAND2_X1 U9906 ( .A1(n7637), .A2(n7636), .ZN(n7664) );
  OR2_X1 U9907 ( .A1(n7637), .A2(n7636), .ZN(n7638) );
  NAND2_X1 U9908 ( .A1(n8282), .A2(n10019), .ZN(n7647) );
  OR2_X1 U9909 ( .A1(n7588), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n7640) );
  NAND2_X1 U9910 ( .A1(n7640), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7639) );
  MUX2_X1 U9911 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7639), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n7643) );
  INV_X1 U9912 ( .A(n7640), .ZN(n7642) );
  INV_X1 U9913 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n7641) );
  NAND2_X1 U9914 ( .A1(n7642), .A2(n7641), .ZN(n7661) );
  NAND2_X1 U9915 ( .A1(n7643), .A2(n7661), .ZN(n14575) );
  OR2_X1 U9916 ( .A1(n10079), .A2(n14575), .ZN(n7646) );
  OR2_X1 U9917 ( .A1(n6492), .A2(n10020), .ZN(n7645) );
  MUX2_X1 U9918 ( .A(n13728), .B(n14718), .S(n7750), .Z(n7649) );
  INV_X1 U9919 ( .A(n14718), .ZN(n13765) );
  MUX2_X1 U9920 ( .A(n13840), .B(n13765), .S(n8284), .Z(n7648) );
  NAND2_X1 U9921 ( .A1(n7650), .A2(n7649), .ZN(n7678) );
  NAND2_X1 U9922 ( .A1(n7680), .A2(n7678), .ZN(n7673) );
  NAND2_X1 U9923 ( .A1(n7651), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7659) );
  OR2_X1 U9924 ( .A1(n7624), .A2(n14768), .ZN(n7658) );
  NOR2_X1 U9925 ( .A1(n7653), .A2(n7652), .ZN(n7694) );
  INV_X1 U9926 ( .A(n7694), .ZN(n7696) );
  NAND2_X1 U9927 ( .A1(n7653), .A2(n7652), .ZN(n7654) );
  NAND2_X1 U9928 ( .A1(n7696), .A2(n7654), .ZN(n13726) );
  OR2_X1 U9929 ( .A1(n7603), .A2(n13726), .ZN(n7657) );
  INV_X1 U9930 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7655) );
  OR2_X1 U9931 ( .A1(n8248), .A2(n7655), .ZN(n7656) );
  NAND4_X1 U9932 ( .A1(n7659), .A2(n7658), .A3(n7657), .A4(n7656), .ZN(n13839)
         );
  NAND2_X1 U9933 ( .A1(n7661), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7660) );
  MUX2_X1 U9934 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7660), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n7662) );
  NAND2_X1 U9935 ( .A1(n7662), .A2(n7719), .ZN(n10198) );
  MUX2_X1 U9936 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n8119), .Z(n7665) );
  NAND2_X1 U9937 ( .A1(n7665), .A2(SI_5_), .ZN(n7683) );
  OAI21_X1 U9938 ( .B1(n7665), .B2(SI_5_), .A(n7683), .ZN(n7666) );
  INV_X1 U9939 ( .A(n7666), .ZN(n7667) );
  OR2_X1 U9940 ( .A1(n7668), .A2(n7667), .ZN(n7669) );
  NAND2_X1 U9941 ( .A1(n7684), .A2(n7669), .ZN(n10063) );
  OR2_X1 U9942 ( .A1(n10063), .A2(n7670), .ZN(n7672) );
  OR2_X1 U9943 ( .A1(n6492), .A2(n10025), .ZN(n7671) );
  OAI211_X1 U9944 ( .C1(n10079), .C2(n10198), .A(n7672), .B(n7671), .ZN(n14724) );
  MUX2_X1 U9945 ( .A(n13839), .B(n14724), .S(n8284), .Z(n7676) );
  NAND2_X1 U9946 ( .A1(n7673), .A2(n7676), .ZN(n7675) );
  MUX2_X1 U9947 ( .A(n14724), .B(n13839), .S(n8284), .Z(n7674) );
  NAND2_X1 U9948 ( .A1(n7675), .A2(n7674), .ZN(n7682) );
  INV_X1 U9949 ( .A(n7676), .ZN(n7677) );
  AND2_X1 U9950 ( .A1(n7678), .A2(n7677), .ZN(n7679) );
  NAND2_X1 U9951 ( .A1(n7680), .A2(n7679), .ZN(n7681) );
  NAND2_X1 U9952 ( .A1(n7682), .A2(n7681), .ZN(n7704) );
  MUX2_X1 U9953 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n8119), .Z(n7685) );
  NAND2_X1 U9954 ( .A1(n7685), .A2(SI_6_), .ZN(n7713) );
  OAI21_X1 U9955 ( .B1(SI_6_), .B2(n7685), .A(n7713), .ZN(n7686) );
  INV_X1 U9956 ( .A(n7686), .ZN(n7687) );
  NAND2_X1 U9957 ( .A1(n7714), .A2(n7689), .ZN(n10065) );
  OR2_X1 U9958 ( .A1(n10065), .A2(n7670), .ZN(n7692) );
  NAND2_X1 U9959 ( .A1(n7719), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7690) );
  XNOR2_X1 U9960 ( .A(n7690), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10161) );
  AOI22_X1 U9961 ( .A1(n7990), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n7989), .B2(
        n10161), .ZN(n7691) );
  NAND2_X1 U9962 ( .A1(n7692), .A2(n7691), .ZN(n11512) );
  NAND2_X1 U9963 ( .A1(n7693), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n7701) );
  INV_X1 U9964 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10141) );
  OR2_X1 U9965 ( .A1(n7624), .A2(n10141), .ZN(n7700) );
  INV_X1 U9966 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n11144) );
  OR2_X1 U9967 ( .A1(n8246), .A2(n11144), .ZN(n7699) );
  NAND2_X1 U9968 ( .A1(n7694), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7706) );
  INV_X1 U9969 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7695) );
  NAND2_X1 U9970 ( .A1(n7696), .A2(n7695), .ZN(n7697) );
  NAND2_X1 U9971 ( .A1(n7706), .A2(n7697), .ZN(n11481) );
  OR2_X1 U9972 ( .A1(n7603), .A2(n11481), .ZN(n7698) );
  NAND4_X1 U9973 ( .A1(n7701), .A2(n7700), .A3(n7699), .A4(n7698), .ZN(n13838)
         );
  MUX2_X1 U9974 ( .A(n11512), .B(n13838), .S(n8284), .Z(n7703) );
  MUX2_X1 U9975 ( .A(n13838), .B(n11512), .S(n8284), .Z(n7702) );
  NAND2_X1 U9976 ( .A1(n8240), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7712) );
  INV_X1 U9977 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10162) );
  OR2_X1 U9978 ( .A1(n8246), .A2(n10162), .ZN(n7711) );
  NAND2_X1 U9979 ( .A1(n7706), .A2(n7705), .ZN(n7707) );
  NAND2_X1 U9980 ( .A1(n7732), .A2(n7707), .ZN(n11642) );
  OR2_X1 U9981 ( .A1(n7603), .A2(n11642), .ZN(n7710) );
  INV_X1 U9982 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7708) );
  OR2_X1 U9983 ( .A1(n8248), .A2(n7708), .ZN(n7709) );
  NAND4_X1 U9984 ( .A1(n7712), .A2(n7711), .A3(n7710), .A4(n7709), .ZN(n13837)
         );
  MUX2_X1 U9985 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n8119), .Z(n7715) );
  OAI21_X1 U9986 ( .B1(SI_7_), .B2(n7715), .A(n7738), .ZN(n7716) );
  INV_X1 U9987 ( .A(n7716), .ZN(n7717) );
  OR2_X1 U9988 ( .A1(n10071), .A2(n7670), .ZN(n7722) );
  OAI21_X1 U9989 ( .B1(n7719), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7720) );
  XNOR2_X1 U9990 ( .A(n7720), .B(P1_IR_REG_7__SCAN_IN), .ZN(n13890) );
  AOI22_X1 U9991 ( .A1(n7990), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7989), .B2(
        n13890), .ZN(n7721) );
  NAND2_X1 U9992 ( .A1(n7722), .A2(n7721), .ZN(n14647) );
  MUX2_X1 U9993 ( .A(n13837), .B(n14647), .S(n8284), .Z(n7726) );
  MUX2_X1 U9994 ( .A(n13837), .B(n14647), .S(n8212), .Z(n7723) );
  NAND2_X1 U9995 ( .A1(n7724), .A2(n7723), .ZN(n7730) );
  INV_X1 U9996 ( .A(n7725), .ZN(n7728) );
  INV_X1 U9997 ( .A(n7726), .ZN(n7727) );
  NAND2_X1 U9998 ( .A1(n7728), .A2(n7727), .ZN(n7729) );
  NAND2_X1 U9999 ( .A1(n7730), .A2(n7729), .ZN(n7752) );
  NAND2_X1 U10000 ( .A1(n7693), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n7737) );
  INV_X1 U10001 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10127) );
  OR2_X1 U10002 ( .A1(n7624), .A2(n10127), .ZN(n7736) );
  NAND2_X1 U10003 ( .A1(n7732), .A2(n7731), .ZN(n7733) );
  NAND2_X1 U10004 ( .A1(n7756), .A2(n7733), .ZN(n11604) );
  OR2_X1 U10005 ( .A1(n7603), .A2(n11604), .ZN(n7735) );
  INV_X1 U10006 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n11101) );
  OR2_X1 U10007 ( .A1(n8246), .A2(n11101), .ZN(n7734) );
  NAND4_X1 U10008 ( .A1(n7737), .A2(n7736), .A3(n7735), .A4(n7734), .ZN(n13836) );
  MUX2_X1 U10009 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n8119), .Z(n7740) );
  NAND2_X1 U10010 ( .A1(n7740), .A2(SI_8_), .ZN(n7762) );
  OAI21_X1 U10011 ( .B1(SI_8_), .B2(n7740), .A(n7762), .ZN(n7741) );
  INV_X1 U10012 ( .A(n7741), .ZN(n7742) );
  NAND2_X1 U10013 ( .A1(n7763), .A2(n7743), .ZN(n10077) );
  OR2_X1 U10014 ( .A1(n10077), .A2(n7670), .ZN(n7749) );
  INV_X1 U10015 ( .A(n7744), .ZN(n7746) );
  NAND2_X1 U10016 ( .A1(n7746), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7745) );
  MUX2_X1 U10017 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7745), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n7747) );
  NOR2_X1 U10018 ( .A1(n7746), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n7797) );
  INV_X1 U10019 ( .A(n7797), .ZN(n7769) );
  NAND2_X1 U10020 ( .A1(n7747), .A2(n7769), .ZN(n10178) );
  INV_X1 U10021 ( .A(n10178), .ZN(n10152) );
  AOI22_X1 U10022 ( .A1(n7990), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7989), .B2(
        n10152), .ZN(n7748) );
  MUX2_X1 U10024 ( .A(n13836), .B(n11589), .S(n8212), .Z(n7753) );
  MUX2_X1 U10025 ( .A(n13836), .B(n11589), .S(n8284), .Z(n7751) );
  INV_X1 U10026 ( .A(n7753), .ZN(n7754) );
  NAND2_X1 U10027 ( .A1(n7693), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7761) );
  INV_X1 U10028 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7755) );
  OR2_X1 U10029 ( .A1(n7624), .A2(n7755), .ZN(n7760) );
  INV_X1 U10030 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n11430) );
  OR2_X1 U10031 ( .A1(n8246), .A2(n11430), .ZN(n7759) );
  INV_X1 U10032 ( .A(n7780), .ZN(n7782) );
  NAND2_X1 U10033 ( .A1(n7756), .A2(n10176), .ZN(n7757) );
  NAND2_X1 U10034 ( .A1(n7782), .A2(n7757), .ZN(n11680) );
  OR2_X1 U10035 ( .A1(n7603), .A2(n11680), .ZN(n7758) );
  NAND4_X1 U10036 ( .A1(n7761), .A2(n7760), .A3(n7759), .A4(n7758), .ZN(n13835) );
  MUX2_X1 U10037 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n8119), .Z(n7764) );
  NAND2_X1 U10038 ( .A1(n7764), .A2(SI_9_), .ZN(n7789) );
  OAI21_X1 U10039 ( .B1(SI_9_), .B2(n7764), .A(n7789), .ZN(n7765) );
  INV_X1 U10040 ( .A(n7765), .ZN(n7766) );
  OR2_X1 U10041 ( .A1(n7767), .A2(n7766), .ZN(n7768) );
  NAND2_X1 U10042 ( .A1(n7790), .A2(n7768), .ZN(n10085) );
  OR2_X1 U10043 ( .A1(n10085), .A2(n7670), .ZN(n7772) );
  NAND2_X1 U10044 ( .A1(n7769), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7770) );
  XNOR2_X1 U10045 ( .A(n7770), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10384) );
  AOI22_X1 U10046 ( .A1(n7990), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7989), .B2(
        n10384), .ZN(n7771) );
  MUX2_X1 U10047 ( .A(n13835), .B(n11674), .S(n8284), .Z(n7776) );
  MUX2_X1 U10048 ( .A(n13835), .B(n11674), .S(n8212), .Z(n7773) );
  NAND2_X1 U10049 ( .A1(n7774), .A2(n7773), .ZN(n7779) );
  INV_X1 U10050 ( .A(n7775), .ZN(n7777) );
  NAND2_X1 U10051 ( .A1(n7777), .A2(n7205), .ZN(n7778) );
  NAND2_X1 U10052 ( .A1(n7779), .A2(n7778), .ZN(n7803) );
  NAND2_X1 U10053 ( .A1(n8240), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7788) );
  INV_X1 U10054 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10441) );
  OR2_X1 U10055 ( .A1(n8246), .A2(n10441), .ZN(n7787) );
  INV_X1 U10056 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7781) );
  NAND2_X1 U10057 ( .A1(n7782), .A2(n7781), .ZN(n7783) );
  NAND2_X1 U10058 ( .A1(n7807), .A2(n7783), .ZN(n14624) );
  OR2_X1 U10059 ( .A1(n7603), .A2(n14624), .ZN(n7786) );
  INV_X1 U10060 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7784) );
  OR2_X1 U10061 ( .A1(n8248), .A2(n7784), .ZN(n7785) );
  NAND4_X1 U10062 ( .A1(n7788), .A2(n7787), .A3(n7786), .A4(n7785), .ZN(n13834) );
  MUX2_X1 U10063 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n8119), .Z(n7791) );
  OAI21_X1 U10064 ( .B1(SI_10_), .B2(n7791), .A(n7814), .ZN(n7792) );
  INV_X1 U10065 ( .A(n7792), .ZN(n7793) );
  OR2_X1 U10066 ( .A1(n7794), .A2(n7793), .ZN(n7795) );
  NAND2_X1 U10067 ( .A1(n7815), .A2(n7795), .ZN(n10089) );
  OR2_X1 U10068 ( .A1(n10089), .A2(n7670), .ZN(n7801) );
  INV_X1 U10069 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n7796) );
  AND2_X1 U10070 ( .A1(n7797), .A2(n7796), .ZN(n7817) );
  INV_X1 U10071 ( .A(n7817), .ZN(n7798) );
  NAND2_X1 U10072 ( .A1(n7798), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7799) );
  XNOR2_X1 U10073 ( .A(n7799), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10432) );
  AOI22_X1 U10074 ( .A1(n7990), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7989), 
        .B2(n10432), .ZN(n7800) );
  MUX2_X1 U10075 ( .A(n13834), .B(n14628), .S(n8212), .Z(n7804) );
  MUX2_X1 U10076 ( .A(n13834), .B(n14628), .S(n8284), .Z(n7802) );
  NAND2_X1 U10077 ( .A1(n7651), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7813) );
  INV_X1 U10078 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7805) );
  OR2_X1 U10079 ( .A1(n7624), .A2(n7805), .ZN(n7812) );
  NAND2_X1 U10080 ( .A1(n7807), .A2(n7806), .ZN(n7808) );
  NAND2_X1 U10081 ( .A1(n7829), .A2(n7808), .ZN(n11862) );
  OR2_X1 U10082 ( .A1(n7603), .A2(n11862), .ZN(n7811) );
  INV_X1 U10083 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7809) );
  OR2_X1 U10084 ( .A1(n8248), .A2(n7809), .ZN(n7810) );
  NAND4_X1 U10085 ( .A1(n7813), .A2(n7812), .A3(n7811), .A4(n7810), .ZN(n14630) );
  MUX2_X1 U10086 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n8119), .Z(n7835) );
  XNOR2_X1 U10087 ( .A(n7838), .B(n7837), .ZN(n10226) );
  NAND2_X1 U10088 ( .A1(n10226), .A2(n8282), .ZN(n7820) );
  INV_X1 U10089 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n7816) );
  NAND2_X1 U10090 ( .A1(n7817), .A2(n7816), .ZN(n7839) );
  NAND2_X1 U10091 ( .A1(n7839), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7818) );
  XNOR2_X1 U10092 ( .A(n7818), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10445) );
  AOI22_X1 U10093 ( .A1(n7990), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7989), 
        .B2(n10445), .ZN(n7819) );
  NAND2_X1 U10094 ( .A1(n7820), .A2(n7819), .ZN(n11656) );
  MUX2_X1 U10095 ( .A(n14630), .B(n11656), .S(n8284), .Z(n7824) );
  MUX2_X1 U10096 ( .A(n14630), .B(n11656), .S(n8212), .Z(n7821) );
  NAND2_X1 U10097 ( .A1(n7822), .A2(n7821), .ZN(n7827) );
  INV_X1 U10098 ( .A(n7823), .ZN(n7825) );
  NAND2_X1 U10099 ( .A1(n7825), .A2(n7199), .ZN(n7826) );
  NAND2_X1 U10100 ( .A1(n7693), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7834) );
  INV_X1 U10101 ( .A(n7861), .ZN(n7876) );
  NAND2_X1 U10102 ( .A1(n7829), .A2(n7828), .ZN(n7830) );
  NAND2_X1 U10103 ( .A1(n7876), .A2(n7830), .ZN(n11907) );
  OR2_X1 U10104 ( .A1(n7603), .A2(n11907), .ZN(n7833) );
  INV_X1 U10105 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10540) );
  OR2_X1 U10106 ( .A1(n7624), .A2(n10540), .ZN(n7832) );
  INV_X1 U10107 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11693) );
  OR2_X1 U10108 ( .A1(n8246), .A2(n11693), .ZN(n7831) );
  NAND4_X1 U10109 ( .A1(n7834), .A2(n7833), .A3(n7832), .A4(n7831), .ZN(n13833) );
  INV_X1 U10110 ( .A(n7835), .ZN(n7836) );
  MUX2_X1 U10111 ( .A(n8385), .B(n10430), .S(n6720), .Z(n7848) );
  XNOR2_X1 U10112 ( .A(n7847), .B(n7846), .ZN(n10399) );
  NAND2_X1 U10113 ( .A1(n10399), .A2(n8282), .ZN(n7842) );
  NAND2_X1 U10114 ( .A1(n7840), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7853) );
  XNOR2_X1 U10115 ( .A(n7853), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10650) );
  AOI22_X1 U10116 ( .A1(n7990), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7989), 
        .B2(n10650), .ZN(n7841) );
  MUX2_X1 U10117 ( .A(n13833), .B(n11900), .S(n8212), .Z(n7844) );
  MUX2_X1 U10118 ( .A(n13833), .B(n11900), .S(n8284), .Z(n7843) );
  INV_X1 U10119 ( .A(n7844), .ZN(n7845) );
  NAND2_X1 U10120 ( .A1(n7848), .A2(n15312), .ZN(n7849) );
  MUX2_X1 U10121 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n6720), .Z(n7868) );
  NAND2_X1 U10122 ( .A1(n7868), .A2(SI_13_), .ZN(n7894) );
  NAND2_X1 U10123 ( .A1(n7896), .A2(n7894), .ZN(n7850) );
  NAND2_X1 U10124 ( .A1(n7850), .A2(SI_14_), .ZN(n7851) );
  NAND2_X1 U10125 ( .A1(n7888), .A2(n7851), .ZN(n7891) );
  MUX2_X1 U10126 ( .A(n10685), .B(n10695), .S(n6720), .Z(n7898) );
  INV_X1 U10127 ( .A(n7898), .ZN(n7890) );
  XNOR2_X1 U10128 ( .A(n7891), .B(n7890), .ZN(n10684) );
  NAND2_X1 U10129 ( .A1(n10684), .A2(n8282), .ZN(n7859) );
  INV_X1 U10130 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n7852) );
  NAND2_X1 U10131 ( .A1(n7853), .A2(n7852), .ZN(n7854) );
  NAND2_X1 U10132 ( .A1(n7854), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7872) );
  INV_X1 U10133 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n7855) );
  NAND2_X1 U10134 ( .A1(n7872), .A2(n7855), .ZN(n7856) );
  NAND2_X1 U10135 ( .A1(n7856), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7857) );
  XNOR2_X1 U10136 ( .A(n7857), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10663) );
  AOI22_X1 U10137 ( .A1(n7990), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7989), 
        .B2(n10663), .ZN(n7858) );
  NAND2_X1 U10138 ( .A1(n7693), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7867) );
  INV_X1 U10139 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n14485) );
  OR2_X1 U10140 ( .A1(n8246), .A2(n14485), .ZN(n7866) );
  INV_X1 U10141 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7860) );
  OR2_X1 U10142 ( .A1(n7624), .A2(n7860), .ZN(n7865) );
  NAND2_X1 U10143 ( .A1(n7861), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7878) );
  INV_X1 U10144 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7862) );
  NAND2_X1 U10145 ( .A1(n7878), .A2(n7862), .ZN(n7863) );
  NAND2_X1 U10146 ( .A1(n7908), .A2(n7863), .ZN(n14484) );
  OR2_X1 U10147 ( .A1(n7603), .A2(n14484), .ZN(n7864) );
  NAND2_X1 U10148 ( .A1(n14511), .A2(n13807), .ZN(n7914) );
  INV_X1 U10149 ( .A(n7868), .ZN(n7869) );
  XNOR2_X1 U10150 ( .A(n7869), .B(SI_13_), .ZN(n7870) );
  XNOR2_X1 U10151 ( .A(n7871), .B(n7870), .ZN(n10516) );
  NAND2_X1 U10152 ( .A1(n10516), .A2(n8282), .ZN(n7874) );
  XNOR2_X1 U10153 ( .A(n7872), .B(P1_IR_REG_13__SCAN_IN), .ZN(n14592) );
  AOI22_X1 U10154 ( .A1(n7990), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7989), 
        .B2(n14592), .ZN(n7873) );
  INV_X1 U10155 ( .A(n14518), .ZN(n11959) );
  INV_X1 U10156 ( .A(n8212), .ZN(n8256) );
  NAND2_X1 U10157 ( .A1(n7693), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n7882) );
  INV_X1 U10158 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10652) );
  OR2_X1 U10159 ( .A1(n7624), .A2(n10652), .ZN(n7881) );
  INV_X1 U10160 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7875) );
  NAND2_X1 U10161 ( .A1(n7876), .A2(n7875), .ZN(n7877) );
  NAND2_X1 U10162 ( .A1(n7878), .A2(n7877), .ZN(n11965) );
  OR2_X1 U10163 ( .A1(n7603), .A2(n11965), .ZN(n7880) );
  INV_X1 U10164 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11813) );
  OR2_X1 U10165 ( .A1(n8246), .A2(n11813), .ZN(n7879) );
  NAND4_X1 U10166 ( .A1(n7882), .A2(n7881), .A3(n7880), .A4(n7879), .ZN(n14483) );
  MUX2_X1 U10167 ( .A(n14483), .B(n14518), .S(n8284), .Z(n7919) );
  NAND2_X1 U10168 ( .A1(n14483), .A2(n8256), .ZN(n7883) );
  OAI211_X1 U10169 ( .C1(n11959), .C2(n8256), .A(n7919), .B(n7883), .ZN(n7884)
         );
  MUX2_X1 U10170 ( .A(n10633), .B(n10635), .S(n6720), .Z(n7885) );
  NAND2_X1 U10171 ( .A1(n7885), .A2(n15224), .ZN(n7945) );
  INV_X1 U10172 ( .A(n7885), .ZN(n7886) );
  NAND2_X1 U10173 ( .A1(n7886), .A2(SI_15_), .ZN(n7887) );
  NAND2_X1 U10174 ( .A1(n7945), .A2(n7887), .ZN(n7893) );
  AND2_X1 U10175 ( .A1(n7888), .A2(n7893), .ZN(n7889) );
  OAI21_X1 U10176 ( .B1(n7891), .B2(n7890), .A(n7889), .ZN(n7902) );
  AND2_X1 U10177 ( .A1(n7894), .A2(n7897), .ZN(n7895) );
  INV_X1 U10178 ( .A(n7897), .ZN(n7900) );
  NAND2_X1 U10179 ( .A1(n7898), .A2(n15263), .ZN(n7899) );
  NAND2_X1 U10180 ( .A1(n7902), .A2(n7934), .ZN(n10632) );
  NAND2_X1 U10181 ( .A1(n10632), .A2(n8282), .ZN(n7906) );
  NAND2_X1 U10182 ( .A1(n7903), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7904) );
  XNOR2_X1 U10183 ( .A(n7904), .B(P1_IR_REG_15__SCAN_IN), .ZN(n11300) );
  AOI22_X1 U10184 ( .A1(n7990), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7989), 
        .B2(n11300), .ZN(n7905) );
  NAND2_X1 U10185 ( .A1(n7693), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n7913) );
  INV_X1 U10186 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11875) );
  OR2_X1 U10187 ( .A1(n8246), .A2(n11875), .ZN(n7912) );
  INV_X1 U10188 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7907) );
  OR2_X1 U10189 ( .A1(n7624), .A2(n7907), .ZN(n7911) );
  INV_X1 U10190 ( .A(n7925), .ZN(n7927) );
  NAND2_X1 U10191 ( .A1(n7908), .A2(n13806), .ZN(n7909) );
  NAND2_X1 U10192 ( .A1(n7927), .A2(n7909), .ZN(n13812) );
  OR2_X1 U10193 ( .A1(n7603), .A2(n13812), .ZN(n7910) );
  AOI21_X1 U10194 ( .B1(n9917), .B2(n9915), .A(n7750), .ZN(n7916) );
  NAND2_X1 U10195 ( .A1(n14503), .A2(n13714), .ZN(n8296) );
  AOI21_X1 U10196 ( .B1(n8296), .B2(n7914), .A(n8256), .ZN(n7915) );
  NOR2_X1 U10197 ( .A1(n7916), .A2(n7915), .ZN(n7921) );
  INV_X1 U10198 ( .A(n14475), .ZN(n14472) );
  INV_X1 U10199 ( .A(n14483), .ZN(n12003) );
  NAND2_X1 U10200 ( .A1(n12003), .A2(n8256), .ZN(n7917) );
  OAI21_X1 U10201 ( .B1(n14518), .B2(n8256), .A(n7917), .ZN(n7918) );
  OR3_X1 U10202 ( .A1(n14472), .A2(n7919), .A3(n7918), .ZN(n7920) );
  NAND3_X1 U10203 ( .A1(n7922), .A2(n7921), .A3(n7920), .ZN(n7924) );
  MUX2_X1 U10204 ( .A(n8296), .B(n9917), .S(n8212), .Z(n7923) );
  NAND2_X1 U10205 ( .A1(n7924), .A2(n7923), .ZN(n7983) );
  INV_X1 U10206 ( .A(n7959), .ZN(n7969) );
  INV_X1 U10207 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7926) );
  NAND2_X1 U10208 ( .A1(n7927), .A2(n7926), .ZN(n7928) );
  NAND2_X1 U10209 ( .A1(n7969), .A2(n7928), .ZN(n13717) );
  OR2_X1 U10210 ( .A1(n13717), .A2(n7603), .ZN(n7933) );
  INV_X1 U10211 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11297) );
  OR2_X1 U10212 ( .A1(n8246), .A2(n11297), .ZN(n7932) );
  INV_X1 U10213 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n11291) );
  OR2_X1 U10214 ( .A1(n7624), .A2(n11291), .ZN(n7931) );
  INV_X1 U10215 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n7929) );
  OR2_X1 U10216 ( .A1(n8248), .A2(n7929), .ZN(n7930) );
  NAND4_X1 U10217 ( .A1(n7933), .A2(n7932), .A3(n7931), .A4(n7930), .ZN(n13830) );
  NAND2_X1 U10218 ( .A1(n7934), .A2(n7945), .ZN(n7938) );
  MUX2_X1 U10219 ( .A(n10597), .B(n10631), .S(n6720), .Z(n7935) );
  NAND2_X1 U10220 ( .A1(n7935), .A2(n15247), .ZN(n7944) );
  INV_X1 U10221 ( .A(n7935), .ZN(n7936) );
  AND2_X1 U10222 ( .A1(n7944), .A2(n7946), .ZN(n7937) );
  XNOR2_X1 U10223 ( .A(n7938), .B(n7937), .ZN(n10596) );
  NAND2_X1 U10224 ( .A1(n10596), .A2(n8282), .ZN(n7942) );
  NAND2_X1 U10225 ( .A1(n6636), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7939) );
  MUX2_X1 U10226 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7939), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n7940) );
  NAND2_X1 U10227 ( .A1(n7940), .A2(n7546), .ZN(n11616) );
  INV_X1 U10228 ( .A(n11616), .ZN(n11293) );
  AOI22_X1 U10229 ( .A1(n7990), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7989), 
        .B2(n11293), .ZN(n7941) );
  MUX2_X1 U10230 ( .A(n13830), .B(n13719), .S(n8284), .Z(n7984) );
  MUX2_X1 U10231 ( .A(n13830), .B(n13719), .S(n8212), .Z(n7943) );
  MUX2_X1 U10232 ( .A(n10637), .B(n10688), .S(n6720), .Z(n7976) );
  NAND2_X1 U10233 ( .A1(n7948), .A2(n15252), .ZN(n7949) );
  INV_X1 U10234 ( .A(n7953), .ZN(n7951) );
  MUX2_X1 U10235 ( .A(n10913), .B(n10916), .S(n6720), .Z(n7952) );
  NAND2_X1 U10236 ( .A1(n7953), .A2(n7952), .ZN(n7954) );
  NAND2_X1 U10237 ( .A1(n7987), .A2(n7954), .ZN(n10915) );
  OR2_X1 U10238 ( .A1(n10915), .A2(n7670), .ZN(n7958) );
  NAND2_X1 U10239 ( .A1(n7955), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7956) );
  XNOR2_X1 U10240 ( .A(n7956), .B(P1_IR_REG_18__SCAN_IN), .ZN(n13916) );
  AOI22_X1 U10241 ( .A1(n7990), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n7989), 
        .B2(n13916), .ZN(n7957) );
  INV_X1 U10242 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14080) );
  INV_X1 U10243 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n7960) );
  NAND2_X1 U10244 ( .A1(n7971), .A2(n7960), .ZN(n7961) );
  NAND2_X1 U10245 ( .A1(n7994), .A2(n7961), .ZN(n14079) );
  OR2_X1 U10246 ( .A1(n14079), .A2(n7603), .ZN(n7967) );
  INV_X1 U10247 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n7962) );
  OR2_X1 U10248 ( .A1(n7624), .A2(n7962), .ZN(n7965) );
  INV_X1 U10249 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n7963) );
  OR2_X1 U10250 ( .A1(n8248), .A2(n7963), .ZN(n7964) );
  AND2_X1 U10251 ( .A1(n7965), .A2(n7964), .ZN(n7966) );
  OAI211_X1 U10252 ( .C1(n8246), .C2(n14080), .A(n7967), .B(n7966), .ZN(n13829) );
  OR2_X1 U10253 ( .A1(n14172), .A2(n13829), .ZN(n9989) );
  NAND2_X1 U10254 ( .A1(n14172), .A2(n13829), .ZN(n9988) );
  NAND2_X1 U10255 ( .A1(n9989), .A2(n9988), .ZN(n14072) );
  INV_X1 U10256 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n7968) );
  NAND2_X1 U10257 ( .A1(n7969), .A2(n7968), .ZN(n7970) );
  NAND2_X1 U10258 ( .A1(n7971), .A2(n7970), .ZN(n13742) );
  OR2_X1 U10259 ( .A1(n13742), .A2(n7603), .ZN(n7975) );
  NAND2_X1 U10260 ( .A1(n8240), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7974) );
  NAND2_X1 U10261 ( .A1(n7693), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n7973) );
  INV_X1 U10262 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n11978) );
  OR2_X1 U10263 ( .A1(n8246), .A2(n11978), .ZN(n7972) );
  NAND4_X1 U10264 ( .A1(n7975), .A2(n7974), .A3(n7973), .A4(n7972), .ZN(n14074) );
  XNOR2_X1 U10265 ( .A(n7976), .B(SI_17_), .ZN(n7977) );
  XNOR2_X1 U10266 ( .A(n7978), .B(n7977), .ZN(n10636) );
  NAND2_X1 U10267 ( .A1(n10636), .A2(n8282), .ZN(n7981) );
  NAND2_X1 U10268 ( .A1(n7546), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7979) );
  XNOR2_X1 U10269 ( .A(n7979), .B(P1_IR_REG_17__SCAN_IN), .ZN(n11614) );
  AOI22_X1 U10270 ( .A1(n7990), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7989), 
        .B2(n11614), .ZN(n7980) );
  MUX2_X1 U10271 ( .A(n14074), .B(n13734), .S(n8212), .Z(n8001) );
  NAND2_X1 U10272 ( .A1(n13734), .A2(n14074), .ZN(n9987) );
  NAND2_X1 U10273 ( .A1(n8001), .A2(n9987), .ZN(n7982) );
  MUX2_X1 U10274 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n6720), .Z(n8019) );
  XNOR2_X1 U10275 ( .A(n8019), .B(SI_19_), .ZN(n8022) );
  XNOR2_X1 U10276 ( .A(n8023), .B(n8022), .ZN(n12009) );
  NAND2_X1 U10277 ( .A1(n12009), .A2(n8282), .ZN(n7992) );
  AOI22_X1 U10278 ( .A1(n7990), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n7988), 
        .B2(n7989), .ZN(n7991) );
  INV_X1 U10279 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n7993) );
  NAND2_X1 U10280 ( .A1(n7994), .A2(n7993), .ZN(n7995) );
  NAND2_X1 U10281 ( .A1(n8011), .A2(n7995), .ZN(n14060) );
  AOI22_X1 U10282 ( .A1(n7651), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n8240), .B2(
        P1_REG1_REG_19__SCAN_IN), .ZN(n7997) );
  NAND2_X1 U10283 ( .A1(n7693), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n7996) );
  OAI211_X1 U10284 ( .C1(n14060), .C2(n7603), .A(n7997), .B(n7996), .ZN(n14075) );
  XNOR2_X1 U10285 ( .A(n14062), .B(n14075), .ZN(n14048) );
  NAND2_X1 U10286 ( .A1(n13829), .A2(n7750), .ZN(n7999) );
  INV_X1 U10287 ( .A(n13829), .ZN(n14054) );
  NAND2_X1 U10288 ( .A1(n14054), .A2(n8256), .ZN(n7998) );
  MUX2_X1 U10289 ( .A(n7999), .B(n7998), .S(n14172), .Z(n8000) );
  INV_X1 U10290 ( .A(n8001), .ZN(n8002) );
  OR2_X1 U10291 ( .A1(n13734), .A2(n14074), .ZN(n9985) );
  NAND3_X1 U10292 ( .A1(n14072), .A2(n8002), .A3(n9985), .ZN(n8003) );
  NAND2_X1 U10293 ( .A1(n14062), .A2(n7750), .ZN(n8007) );
  OR2_X1 U10294 ( .A1(n14062), .A2(n8212), .ZN(n8006) );
  MUX2_X1 U10295 ( .A(n8007), .B(n8006), .S(n14075), .Z(n8008) );
  NAND2_X1 U10296 ( .A1(n8009), .A2(n8008), .ZN(n8032) );
  INV_X1 U10297 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8010) );
  INV_X1 U10298 ( .A(n8044), .ZN(n8045) );
  NAND2_X1 U10299 ( .A1(n8011), .A2(n8010), .ZN(n8012) );
  NAND2_X1 U10300 ( .A1(n14036), .A2(n8181), .ZN(n8018) );
  INV_X1 U10301 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n8015) );
  NAND2_X1 U10302 ( .A1(n8240), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n8014) );
  NAND2_X1 U10303 ( .A1(n7651), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8013) );
  OAI211_X1 U10304 ( .C1(n8015), .C2(n8248), .A(n8014), .B(n8013), .ZN(n8016)
         );
  INV_X1 U10305 ( .A(n8016), .ZN(n8017) );
  NAND2_X1 U10306 ( .A1(n8018), .A2(n8017), .ZN(n13828) );
  INV_X1 U10307 ( .A(n8019), .ZN(n8020) );
  INV_X1 U10308 ( .A(SI_19_), .ZN(n10687) );
  NAND2_X1 U10309 ( .A1(n8020), .A2(n10687), .ZN(n8021) );
  INV_X1 U10310 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11420) );
  INV_X1 U10311 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11436) );
  MUX2_X1 U10312 ( .A(n11420), .B(n11436), .S(n8119), .Z(n8036) );
  OR2_X1 U10313 ( .A1(n8037), .A2(n8036), .ZN(n8038) );
  NAND2_X1 U10314 ( .A1(n8037), .A2(n8036), .ZN(n8026) );
  OR2_X1 U10315 ( .A1(n6492), .A2(n11420), .ZN(n8027) );
  MUX2_X1 U10316 ( .A(n13828), .B(n14159), .S(n8284), .Z(n8029) );
  INV_X1 U10317 ( .A(n8029), .ZN(n8031) );
  MUX2_X1 U10318 ( .A(n14159), .B(n13828), .S(n8284), .Z(n8030) );
  OAI21_X1 U10319 ( .B1(n8032), .B2(n8031), .A(n8030), .ZN(n8034) );
  NAND2_X1 U10320 ( .A1(n8032), .A2(n8031), .ZN(n8033) );
  NAND2_X1 U10321 ( .A1(n8034), .A2(n8033), .ZN(n8055) );
  MUX2_X1 U10322 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n8119), .Z(n8035) );
  NAND2_X1 U10323 ( .A1(n8035), .A2(SI_21_), .ZN(n8069) );
  OAI21_X1 U10324 ( .B1(SI_21_), .B2(n8035), .A(n8069), .ZN(n8039) );
  NAND2_X1 U10325 ( .A1(n8038), .A2(n7491), .ZN(n8040) );
  NAND2_X1 U10326 ( .A1(n6610), .A2(n8041), .ZN(n11547) );
  OR2_X1 U10327 ( .A1(n11547), .A2(n7670), .ZN(n8043) );
  INV_X1 U10328 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11544) );
  OR2_X1 U10329 ( .A1(n6492), .A2(n11544), .ZN(n8042) );
  INV_X1 U10330 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n13692) );
  NAND2_X1 U10331 ( .A1(n8045), .A2(n13692), .ZN(n8046) );
  NAND2_X1 U10332 ( .A1(n8061), .A2(n8046), .ZN(n14025) );
  OR2_X1 U10333 ( .A1(n14025), .A2(n7603), .ZN(n8052) );
  INV_X1 U10334 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n8049) );
  NAND2_X1 U10335 ( .A1(n7651), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8048) );
  NAND2_X1 U10336 ( .A1(n8240), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n8047) );
  OAI211_X1 U10337 ( .C1(n8049), .C2(n8248), .A(n8048), .B(n8047), .ZN(n8050)
         );
  INV_X1 U10338 ( .A(n8050), .ZN(n8051) );
  NAND2_X1 U10339 ( .A1(n8052), .A2(n8051), .ZN(n13827) );
  MUX2_X1 U10340 ( .A(n14151), .B(n13827), .S(n8256), .Z(n8056) );
  NAND2_X1 U10341 ( .A1(n8055), .A2(n8056), .ZN(n8054) );
  MUX2_X1 U10342 ( .A(n14151), .B(n13827), .S(n8212), .Z(n8053) );
  NAND2_X1 U10343 ( .A1(n8054), .A2(n8053), .ZN(n8060) );
  INV_X1 U10344 ( .A(n8055), .ZN(n8058) );
  INV_X1 U10345 ( .A(n8056), .ZN(n8057) );
  NAND2_X1 U10346 ( .A1(n8058), .A2(n8057), .ZN(n8059) );
  INV_X1 U10347 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n12105) );
  NAND2_X1 U10348 ( .A1(n8061), .A2(n12105), .ZN(n8062) );
  AND2_X1 U10349 ( .A1(n8077), .A2(n8062), .ZN(n14009) );
  NAND2_X1 U10350 ( .A1(n14009), .A2(n8181), .ZN(n8068) );
  INV_X1 U10351 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n8065) );
  NAND2_X1 U10352 ( .A1(n7651), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8064) );
  NAND2_X1 U10353 ( .A1(n8240), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8063) );
  OAI211_X1 U10354 ( .C1(n8065), .C2(n8248), .A(n8064), .B(n8063), .ZN(n8066)
         );
  INV_X1 U10355 ( .A(n8066), .ZN(n8067) );
  NAND2_X1 U10356 ( .A1(n8095), .A2(SI_22_), .ZN(n8089) );
  INV_X1 U10357 ( .A(n9272), .ZN(n8071) );
  NAND2_X2 U10358 ( .A1(n14216), .A2(n10079), .ZN(n8295) );
  MUX2_X1 U10359 ( .A(n13691), .B(n8295), .S(n8256), .Z(n8075) );
  MUX2_X1 U10360 ( .A(n8295), .B(n13691), .S(n8284), .Z(n8073) );
  INV_X1 U10361 ( .A(n8073), .ZN(n8074) );
  INV_X1 U10362 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n13675) );
  NAND2_X1 U10363 ( .A1(n8077), .A2(n13675), .ZN(n8078) );
  NAND2_X1 U10364 ( .A1(n8107), .A2(n8078), .ZN(n13993) );
  OR2_X1 U10365 ( .A1(n13993), .A2(n7603), .ZN(n8084) );
  INV_X1 U10366 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n8081) );
  NAND2_X1 U10367 ( .A1(n7651), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8080) );
  NAND2_X1 U10368 ( .A1(n8240), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8079) );
  OAI211_X1 U10369 ( .C1(n8081), .C2(n8248), .A(n8080), .B(n8079), .ZN(n8082)
         );
  INV_X1 U10370 ( .A(n8082), .ZN(n8083) );
  NAND2_X1 U10371 ( .A1(n8084), .A2(n8083), .ZN(n13825) );
  INV_X1 U10372 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8409) );
  MUX2_X1 U10373 ( .A(n8408), .B(n8409), .S(n8119), .Z(n9271) );
  INV_X1 U10374 ( .A(n9271), .ZN(n8085) );
  MUX2_X1 U10375 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n6720), .Z(n8086) );
  NAND2_X1 U10376 ( .A1(n8086), .A2(SI_23_), .ZN(n8115) );
  INV_X1 U10377 ( .A(n8086), .ZN(n8087) );
  INV_X1 U10378 ( .A(SI_23_), .ZN(n11311) );
  NAND2_X1 U10379 ( .A1(n8087), .A2(n11311), .ZN(n8088) );
  NAND2_X1 U10380 ( .A1(n8115), .A2(n8088), .ZN(n8092) );
  AND2_X1 U10381 ( .A1(n8089), .A2(n8092), .ZN(n8096) );
  INV_X1 U10382 ( .A(SI_22_), .ZN(n8090) );
  NOR2_X1 U10383 ( .A1(n9271), .A2(n8090), .ZN(n8094) );
  NOR2_X1 U10384 ( .A1(n8085), .A2(SI_22_), .ZN(n8091) );
  NOR2_X1 U10385 ( .A1(n8092), .A2(n8091), .ZN(n8093) );
  NAND2_X1 U10386 ( .A1(n11827), .A2(n8282), .ZN(n8098) );
  INV_X1 U10387 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11830) );
  OR2_X1 U10388 ( .A1(n6492), .A2(n11830), .ZN(n8097) );
  MUX2_X1 U10389 ( .A(n13825), .B(n14138), .S(n8212), .Z(n8102) );
  NAND2_X1 U10390 ( .A1(n8101), .A2(n8102), .ZN(n8100) );
  MUX2_X1 U10391 ( .A(n13825), .B(n14138), .S(n8256), .Z(n8099) );
  NAND2_X1 U10392 ( .A1(n8100), .A2(n8099), .ZN(n8106) );
  INV_X1 U10393 ( .A(n8101), .ZN(n8104) );
  INV_X1 U10394 ( .A(n8102), .ZN(n8103) );
  NAND2_X1 U10395 ( .A1(n8104), .A2(n8103), .ZN(n8105) );
  INV_X1 U10396 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n13754) );
  NAND2_X1 U10397 ( .A1(n8107), .A2(n13754), .ZN(n8108) );
  AND2_X1 U10398 ( .A1(n8130), .A2(n8108), .ZN(n13979) );
  NAND2_X1 U10399 ( .A1(n13979), .A2(n8181), .ZN(n8114) );
  INV_X1 U10400 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n8111) );
  NAND2_X1 U10401 ( .A1(n8240), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8110) );
  NAND2_X1 U10402 ( .A1(n7651), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8109) );
  OAI211_X1 U10403 ( .C1(n8111), .C2(n8248), .A(n8110), .B(n8109), .ZN(n8112)
         );
  INV_X1 U10404 ( .A(n8112), .ZN(n8113) );
  NAND2_X1 U10405 ( .A1(n8114), .A2(n8113), .ZN(n13824) );
  INV_X1 U10406 ( .A(n8116), .ZN(n8117) );
  NAND2_X1 U10407 ( .A1(n8117), .A2(n15287), .ZN(n8118) );
  MUX2_X1 U10408 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n6720), .Z(n8121) );
  INV_X1 U10409 ( .A(n8120), .ZN(n8122) );
  NAND2_X1 U10410 ( .A1(n8122), .A2(n6931), .ZN(n8123) );
  NAND2_X1 U10411 ( .A1(n8139), .A2(n8123), .ZN(n11913) );
  OR2_X1 U10412 ( .A1(n11913), .A2(n7670), .ZN(n8125) );
  INV_X1 U10413 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11880) );
  OR2_X1 U10414 ( .A1(n6492), .A2(n11880), .ZN(n8124) );
  MUX2_X1 U10415 ( .A(n13824), .B(n14133), .S(n8284), .Z(n8127) );
  MUX2_X1 U10416 ( .A(n14133), .B(n13824), .S(n8256), .Z(n8126) );
  INV_X1 U10417 ( .A(n8127), .ZN(n8128) );
  INV_X1 U10418 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8129) );
  NAND2_X1 U10419 ( .A1(n8130), .A2(n8129), .ZN(n8131) );
  AND2_X1 U10420 ( .A1(n8160), .A2(n8131), .ZN(n13703) );
  NAND2_X1 U10421 ( .A1(n13703), .A2(n8181), .ZN(n8137) );
  INV_X1 U10422 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n8134) );
  NAND2_X1 U10423 ( .A1(n8240), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8133) );
  NAND2_X1 U10424 ( .A1(n7651), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8132) );
  OAI211_X1 U10425 ( .C1(n8134), .C2(n8248), .A(n8133), .B(n8132), .ZN(n8135)
         );
  INV_X1 U10426 ( .A(n8135), .ZN(n8136) );
  NAND2_X1 U10427 ( .A1(n8137), .A2(n8136), .ZN(n13823) );
  MUX2_X1 U10428 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n8119), .Z(n8152) );
  XNOR2_X1 U10429 ( .A(n8152), .B(SI_25_), .ZN(n8150) );
  XNOR2_X1 U10430 ( .A(n8151), .B(n8150), .ZN(n11984) );
  NAND2_X1 U10431 ( .A1(n11984), .A2(n8282), .ZN(n8141) );
  INV_X1 U10432 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11990) );
  OR2_X1 U10433 ( .A1(n6492), .A2(n11990), .ZN(n8140) );
  MUX2_X1 U10434 ( .A(n13823), .B(n14125), .S(n8212), .Z(n8145) );
  NAND2_X1 U10435 ( .A1(n8144), .A2(n8145), .ZN(n8143) );
  MUX2_X1 U10436 ( .A(n13823), .B(n14125), .S(n8256), .Z(n8142) );
  NAND2_X1 U10437 ( .A1(n8143), .A2(n8142), .ZN(n8149) );
  INV_X1 U10438 ( .A(n8144), .ZN(n8147) );
  INV_X1 U10439 ( .A(n8145), .ZN(n8146) );
  NAND2_X1 U10440 ( .A1(n8147), .A2(n8146), .ZN(n8148) );
  INV_X1 U10441 ( .A(n8152), .ZN(n8153) );
  INV_X1 U10442 ( .A(SI_25_), .ZN(n15304) );
  NAND2_X1 U10443 ( .A1(n8153), .A2(n15304), .ZN(n8154) );
  MUX2_X1 U10444 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n8119), .Z(n8170) );
  INV_X1 U10445 ( .A(SI_26_), .ZN(n15310) );
  XNOR2_X1 U10446 ( .A(n8170), .B(n15310), .ZN(n8155) );
  NAND2_X1 U10447 ( .A1(n13651), .A2(n8282), .ZN(n8157) );
  INV_X1 U10448 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14211) );
  OR2_X1 U10449 ( .A1(n6492), .A2(n14211), .ZN(n8156) );
  INV_X1 U10450 ( .A(n8160), .ZN(n8158) );
  NAND2_X1 U10451 ( .A1(n8158), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8179) );
  INV_X1 U10452 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8159) );
  NAND2_X1 U10453 ( .A1(n8160), .A2(n8159), .ZN(n8161) );
  NAND2_X1 U10454 ( .A1(n8179), .A2(n8161), .ZN(n13797) );
  OR2_X1 U10455 ( .A1(n13797), .A2(n7603), .ZN(n8166) );
  INV_X1 U10456 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n14188) );
  NAND2_X1 U10457 ( .A1(n8240), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8163) );
  NAND2_X1 U10458 ( .A1(n7651), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8162) );
  OAI211_X1 U10459 ( .C1(n14188), .C2(n8248), .A(n8163), .B(n8162), .ZN(n8164)
         );
  INV_X1 U10460 ( .A(n8164), .ZN(n8165) );
  MUX2_X1 U10461 ( .A(n13967), .B(n13822), .S(n8212), .Z(n8168) );
  MUX2_X1 U10462 ( .A(n13967), .B(n13822), .S(n8256), .Z(n8167) );
  INV_X1 U10463 ( .A(n8168), .ZN(n8169) );
  NAND2_X1 U10464 ( .A1(n8171), .A2(n8170), .ZN(n8175) );
  INV_X1 U10465 ( .A(n8172), .ZN(n8173) );
  NAND2_X1 U10466 ( .A1(n8175), .A2(n8174), .ZN(n8209) );
  INV_X1 U10467 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14209) );
  INV_X1 U10468 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13649) );
  MUX2_X1 U10469 ( .A(n14209), .B(n13649), .S(n8119), .Z(n8206) );
  XNOR2_X1 U10470 ( .A(n8206), .B(SI_27_), .ZN(n8208) );
  INV_X1 U10471 ( .A(n8208), .ZN(n8176) );
  NAND2_X1 U10472 ( .A1(n13648), .A2(n8282), .ZN(n8178) );
  OR2_X1 U10473 ( .A1(n6492), .A2(n14209), .ZN(n8177) );
  INV_X1 U10474 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n13663) );
  NAND2_X1 U10475 ( .A1(n8179), .A2(n13663), .ZN(n8180) );
  NAND2_X1 U10476 ( .A1(n13945), .A2(n8181), .ZN(n8187) );
  INV_X1 U10477 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n8184) );
  NAND2_X1 U10478 ( .A1(n7651), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8183) );
  NAND2_X1 U10479 ( .A1(n8240), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8182) );
  OAI211_X1 U10480 ( .C1(n8184), .C2(n6491), .A(n8183), .B(n8182), .ZN(n8185)
         );
  INV_X1 U10481 ( .A(n8185), .ZN(n8186) );
  MUX2_X1 U10482 ( .A(n14112), .B(n13956), .S(n8256), .Z(n8191) );
  NAND2_X1 U10483 ( .A1(n8190), .A2(n8191), .ZN(n8189) );
  MUX2_X1 U10484 ( .A(n13956), .B(n14112), .S(n8256), .Z(n8188) );
  NAND2_X1 U10485 ( .A1(n8189), .A2(n8188), .ZN(n8195) );
  INV_X1 U10486 ( .A(n8190), .ZN(n8193) );
  INV_X1 U10487 ( .A(n8191), .ZN(n8192) );
  NAND2_X1 U10488 ( .A1(n8193), .A2(n8192), .ZN(n8194) );
  INV_X1 U10489 ( .A(n8198), .ZN(n8196) );
  NAND2_X1 U10490 ( .A1(n8196), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n12487) );
  INV_X1 U10491 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8197) );
  NAND2_X1 U10492 ( .A1(n8198), .A2(n8197), .ZN(n8199) );
  NAND2_X1 U10493 ( .A1(n12487), .A2(n8199), .ZN(n12459) );
  OR2_X1 U10494 ( .A1(n12459), .A2(n7603), .ZN(n8205) );
  INV_X1 U10495 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n8202) );
  NAND2_X1 U10496 ( .A1(n7651), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8201) );
  NAND2_X1 U10497 ( .A1(n8240), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8200) );
  OAI211_X1 U10498 ( .C1(n8202), .C2(n6491), .A(n8201), .B(n8200), .ZN(n8203)
         );
  INV_X1 U10499 ( .A(n8203), .ZN(n8204) );
  INV_X1 U10500 ( .A(SI_27_), .ZN(n15265) );
  NOR2_X1 U10501 ( .A1(n8206), .A2(n15265), .ZN(n8207) );
  MUX2_X1 U10502 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n8119), .Z(n8223) );
  INV_X1 U10503 ( .A(SI_28_), .ZN(n15236) );
  XNOR2_X1 U10504 ( .A(n8223), .B(n15236), .ZN(n8221) );
  INV_X1 U10505 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12042) );
  OR2_X1 U10506 ( .A1(n6492), .A2(n12042), .ZN(n8210) );
  MUX2_X1 U10507 ( .A(n13821), .B(n14104), .S(n8212), .Z(n8213) );
  OR2_X1 U10508 ( .A1(n12487), .A2(n7603), .ZN(n8220) );
  INV_X1 U10509 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n8217) );
  NAND2_X1 U10510 ( .A1(n7651), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8216) );
  NAND2_X1 U10511 ( .A1(n8240), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8215) );
  OAI211_X1 U10512 ( .C1(n8217), .C2(n8248), .A(n8216), .B(n8215), .ZN(n8218)
         );
  INV_X1 U10513 ( .A(n8218), .ZN(n8219) );
  NAND2_X1 U10514 ( .A1(n8220), .A2(n8219), .ZN(n13820) );
  NAND2_X1 U10515 ( .A1(n8222), .A2(n8221), .ZN(n8226) );
  INV_X1 U10516 ( .A(n8223), .ZN(n8224) );
  NAND2_X1 U10517 ( .A1(n8224), .A2(n15236), .ZN(n8225) );
  INV_X1 U10518 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n12134) );
  INV_X1 U10519 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13641) );
  MUX2_X1 U10520 ( .A(n12134), .B(n13641), .S(n8119), .Z(n8235) );
  XNOR2_X1 U10521 ( .A(n8235), .B(SI_29_), .ZN(n8233) );
  NAND2_X1 U10522 ( .A1(n12043), .A2(n8282), .ZN(n8228) );
  OR2_X1 U10523 ( .A1(n6492), .A2(n12134), .ZN(n8227) );
  MUX2_X1 U10524 ( .A(n13820), .B(n14096), .S(n8212), .Z(n8231) );
  MUX2_X1 U10525 ( .A(n13820), .B(n14096), .S(n8256), .Z(n8229) );
  INV_X1 U10526 ( .A(n8231), .ZN(n8232) );
  INV_X1 U10527 ( .A(SI_29_), .ZN(n15285) );
  NAND2_X1 U10528 ( .A1(n8235), .A2(n15285), .ZN(n8272) );
  MUX2_X1 U10529 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n8119), .Z(n8269) );
  XNOR2_X1 U10530 ( .A(n8269), .B(SI_30_), .ZN(n8236) );
  INV_X1 U10531 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12526) );
  OR2_X1 U10532 ( .A1(n6492), .A2(n12526), .ZN(n8238) );
  INV_X1 U10533 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n8243) );
  NAND2_X1 U10534 ( .A1(n7651), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8242) );
  NAND2_X1 U10535 ( .A1(n8240), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8241) );
  OAI211_X1 U10536 ( .C1(n6491), .C2(n8243), .A(n8242), .B(n8241), .ZN(n13819)
         );
  INV_X1 U10537 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n8244) );
  OR2_X1 U10538 ( .A1(n7624), .A2(n8244), .ZN(n8251) );
  INV_X1 U10539 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n8245) );
  OR2_X1 U10540 ( .A1(n8246), .A2(n8245), .ZN(n8250) );
  INV_X1 U10541 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n8247) );
  OR2_X1 U10542 ( .A1(n8248), .A2(n8247), .ZN(n8249) );
  AND3_X1 U10543 ( .A1(n8251), .A2(n8250), .A3(n8249), .ZN(n8283) );
  INV_X1 U10544 ( .A(n8252), .ZN(n8253) );
  OAI22_X1 U10545 ( .A1(n8283), .A2(n8256), .B1(n9936), .B2(n8253), .ZN(n8254)
         );
  AOI22_X1 U10546 ( .A1(n13929), .A2(n8256), .B1(n13819), .B2(n8254), .ZN(
        n8258) );
  NAND2_X1 U10547 ( .A1(n8255), .A2(n8258), .ZN(n8262) );
  INV_X1 U10548 ( .A(n8283), .ZN(n13932) );
  NAND2_X1 U10549 ( .A1(n9936), .A2(n9937), .ZN(n9932) );
  OAI21_X1 U10550 ( .B1(n13932), .B2(n9932), .A(n13819), .ZN(n8257) );
  MUX2_X1 U10551 ( .A(n14094), .B(n8257), .S(n8256), .Z(n8261) );
  INV_X1 U10552 ( .A(n8258), .ZN(n8259) );
  AOI22_X1 U10553 ( .A1(n8262), .A2(n8261), .B1(n8260), .B2(n8259), .ZN(n8320)
         );
  INV_X1 U10554 ( .A(n10453), .ZN(n8263) );
  NAND2_X1 U10555 ( .A1(n8263), .A2(n7988), .ZN(n11006) );
  NAND2_X1 U10556 ( .A1(n9936), .A2(n14215), .ZN(n10464) );
  OAI21_X1 U10557 ( .B1(n14215), .B2(n9937), .A(n10464), .ZN(n8264) );
  NAND2_X1 U10558 ( .A1(n11006), .A2(n8264), .ZN(n8318) );
  INV_X1 U10559 ( .A(n9936), .ZN(n11545) );
  NAND2_X1 U10560 ( .A1(n11545), .A2(n9937), .ZN(n10009) );
  NAND2_X1 U10561 ( .A1(n8318), .A2(n10009), .ZN(n8289) );
  INV_X1 U10562 ( .A(n8289), .ZN(n8288) );
  INV_X1 U10563 ( .A(n8269), .ZN(n8270) );
  INV_X1 U10564 ( .A(SI_30_), .ZN(n15229) );
  NOR2_X1 U10565 ( .A1(n8270), .A2(n15229), .ZN(n8273) );
  MUX2_X1 U10566 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n8119), .Z(n8265) );
  XNOR2_X1 U10567 ( .A(n8265), .B(SI_31_), .ZN(n8271) );
  OAI21_X1 U10568 ( .B1(SI_30_), .B2(n8269), .A(n8272), .ZN(n8266) );
  INV_X1 U10569 ( .A(n8271), .ZN(n8274) );
  NOR2_X1 U10570 ( .A1(n8266), .A2(n8274), .ZN(n8267) );
  NAND2_X1 U10571 ( .A1(n8268), .A2(n8267), .ZN(n8279) );
  OAI21_X1 U10572 ( .B1(n8274), .B2(n15229), .A(n8269), .ZN(n8277) );
  OAI21_X1 U10573 ( .B1(n8271), .B2(SI_30_), .A(n8270), .ZN(n8276) );
  NOR2_X1 U10574 ( .A1(n8273), .A2(n8272), .ZN(n8275) );
  AOI22_X1 U10575 ( .A1(n8277), .A2(n8276), .B1(n8275), .B2(n8274), .ZN(n8278)
         );
  INV_X1 U10576 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n8280) );
  NOR2_X1 U10577 ( .A1(n6492), .A2(n8280), .ZN(n8281) );
  INV_X1 U10578 ( .A(n14091), .ZN(n13930) );
  AND2_X1 U10579 ( .A1(n13930), .A2(n8283), .ZN(n8286) );
  NOR2_X1 U10580 ( .A1(n13930), .A2(n8283), .ZN(n8285) );
  MUX2_X1 U10581 ( .A(n8286), .B(n8285), .S(n8284), .Z(n8287) );
  INV_X1 U10582 ( .A(n8287), .ZN(n8291) );
  INV_X1 U10583 ( .A(n8318), .ZN(n8293) );
  XNOR2_X1 U10584 ( .A(n14091), .B(n13932), .ZN(n8319) );
  INV_X1 U10585 ( .A(n8319), .ZN(n8290) );
  NOR2_X1 U10586 ( .A1(n8290), .A2(n8289), .ZN(n8292) );
  MUX2_X1 U10587 ( .A(n8293), .B(n8292), .S(n8291), .Z(n8317) );
  INV_X1 U10588 ( .A(n13956), .ZN(n12463) );
  NAND2_X1 U10589 ( .A1(n14104), .A2(n13821), .ZN(n12475) );
  OR2_X1 U10590 ( .A1(n14104), .A2(n13821), .ZN(n8294) );
  INV_X1 U10591 ( .A(n13824), .ZN(n13705) );
  XNOR2_X1 U10592 ( .A(n14133), .B(n13705), .ZN(n13983) );
  XNOR2_X1 U10593 ( .A(n14138), .B(n13825), .ZN(n13997) );
  INV_X1 U10594 ( .A(n13828), .ZN(n14056) );
  XNOR2_X1 U10595 ( .A(n14159), .B(n14056), .ZN(n14033) );
  INV_X1 U10596 ( .A(n14072), .ZN(n14081) );
  XNOR2_X1 U10597 ( .A(n13719), .B(n13741), .ZN(n11948) );
  NAND2_X1 U10598 ( .A1(n9985), .A2(n9987), .ZN(n9919) );
  NAND2_X1 U10599 ( .A1(n9917), .A2(n8296), .ZN(n9916) );
  XNOR2_X1 U10600 ( .A(n11900), .B(n13833), .ZN(n11688) );
  INV_X1 U10601 ( .A(n13834), .ZN(n11751) );
  OR2_X1 U10602 ( .A1(n14628), .A2(n11751), .ZN(n11658) );
  NAND2_X1 U10603 ( .A1(n14628), .A2(n11751), .ZN(n8297) );
  NAND2_X1 U10604 ( .A1(n11658), .A2(n8297), .ZN(n14627) );
  XNOR2_X1 U10605 ( .A(n11589), .B(n13836), .ZN(n9907) );
  AND2_X1 U10606 ( .A1(n8299), .A2(n8298), .ZN(n14689) );
  XNOR2_X1 U10607 ( .A(n13840), .B(n13765), .ZN(n9963) );
  NAND4_X1 U10608 ( .A1(n14689), .A2(n6482), .A3(n11111), .A4(n9963), .ZN(
        n8300) );
  XNOR2_X1 U10609 ( .A(n13839), .B(n11494), .ZN(n11172) );
  NOR3_X1 U10610 ( .A1(n8300), .A2(n14669), .A3(n11172), .ZN(n8301) );
  XNOR2_X1 U10611 ( .A(n14647), .B(n13837), .ZN(n9971) );
  XNOR2_X1 U10612 ( .A(n11512), .B(n13838), .ZN(n11140) );
  NAND4_X1 U10613 ( .A1(n9907), .A2(n8301), .A3(n9971), .A4(n11140), .ZN(n8302) );
  NOR2_X1 U10614 ( .A1(n14627), .A2(n8302), .ZN(n8303) );
  XNOR2_X1 U10615 ( .A(n11656), .B(n14630), .ZN(n11659) );
  XNOR2_X1 U10616 ( .A(n11674), .B(n13835), .ZN(n11423) );
  NAND4_X1 U10617 ( .A1(n11688), .A2(n8303), .A3(n11659), .A4(n11423), .ZN(
        n8304) );
  NOR2_X1 U10618 ( .A1(n9916), .A2(n8304), .ZN(n8305) );
  XNOR2_X1 U10619 ( .A(n14518), .B(n14483), .ZN(n11818) );
  NAND4_X1 U10620 ( .A1(n9919), .A2(n14475), .A3(n8305), .A4(n11818), .ZN(
        n8306) );
  OR4_X1 U10621 ( .A1(n14051), .A2(n14081), .A3(n11948), .A4(n8306), .ZN(n8307) );
  NOR2_X1 U10622 ( .A1(n14033), .A2(n8307), .ZN(n8308) );
  XNOR2_X1 U10623 ( .A(n14151), .B(n13827), .ZN(n14022) );
  NAND4_X1 U10624 ( .A1(n13997), .A2(n14006), .A3(n8308), .A4(n14022), .ZN(
        n8309) );
  NOR2_X1 U10625 ( .A1(n13983), .A2(n8309), .ZN(n8310) );
  XNOR2_X1 U10626 ( .A(n13967), .B(n13822), .ZN(n13954) );
  XNOR2_X1 U10627 ( .A(n14125), .B(n13823), .ZN(n10004) );
  NAND4_X1 U10628 ( .A1(n12024), .A2(n8310), .A3(n13954), .A4(n10004), .ZN(
        n8311) );
  NOR3_X1 U10629 ( .A1(n8319), .A2(n13940), .A3(n8311), .ZN(n8313) );
  XNOR2_X1 U10630 ( .A(n13929), .B(n13819), .ZN(n8312) );
  NAND3_X1 U10631 ( .A1(n8313), .A2(n8312), .A3(n12481), .ZN(n8314) );
  XOR2_X1 U10632 ( .A(n7988), .B(n8314), .Z(n8315) );
  NOR2_X1 U10633 ( .A1(n8315), .A2(n10009), .ZN(n8316) );
  OAI21_X1 U10634 ( .B1(n8321), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8323) );
  INV_X1 U10635 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8322) );
  XNOR2_X1 U10636 ( .A(n8323), .B(n8322), .ZN(n8326) );
  INV_X1 U10637 ( .A(n8326), .ZN(n10078) );
  NAND2_X1 U10638 ( .A1(n10078), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11828) );
  INV_X1 U10639 ( .A(n10464), .ZN(n8335) );
  INV_X1 U10640 ( .A(n8325), .ZN(n13859) );
  INV_X1 U10641 ( .A(n14206), .ZN(n14562) );
  NAND2_X1 U10642 ( .A1(n6524), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8327) );
  NAND2_X1 U10643 ( .A1(n8328), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8329) );
  MUX2_X1 U10644 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8329), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n8330) );
  NAND2_X1 U10645 ( .A1(n8330), .A2(n6525), .ZN(n11881) );
  NAND2_X1 U10646 ( .A1(n6525), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8331) );
  MUX2_X1 U10647 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8331), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n8332) );
  NAND2_X1 U10648 ( .A1(n11421), .A2(n8333), .ZN(n8334) );
  NAND2_X1 U10649 ( .A1(n8335), .A2(n8334), .ZN(n11233) );
  NAND4_X1 U10650 ( .A1(n14482), .A2(n14562), .A3(n11232), .A4(n11233), .ZN(
        n8336) );
  OAI211_X1 U10651 ( .C1(n14215), .C2(n11828), .A(n8336), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8337) );
  NAND2_X1 U10652 ( .A1(n8538), .A2(n15288), .ZN(n8552) );
  NAND2_X1 U10653 ( .A1(n8672), .A2(n11927), .ZN(n8688) );
  INV_X1 U10654 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n8748) );
  INV_X1 U10655 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n8763) );
  INV_X1 U10656 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n12607) );
  NAND2_X1 U10657 ( .A1(n8788), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8338) );
  INV_X1 U10658 ( .A(n8802), .ZN(n8803) );
  NAND2_X1 U10659 ( .A1(n8338), .A2(n8803), .ZN(n12817) );
  NOR2_X1 U10660 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_12__SCAN_IN), 
        .ZN(n8341) );
  NOR2_X1 U10661 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), .ZN(
        n8340) );
  NOR2_X1 U10662 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), 
        .ZN(n8339) );
  NAND3_X1 U10663 ( .A1(n8344), .A2(n8343), .A3(n8342), .ZN(n8447) );
  NOR2_X1 U10664 ( .A1(n8345), .A2(n8447), .ZN(n8346) );
  NOR2_X1 U10665 ( .A1(P3_IR_REG_26__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), 
        .ZN(n8348) );
  INV_X1 U10666 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12959) );
  NAND2_X1 U10667 ( .A1(n8789), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8357) );
  NAND2_X1 U10668 ( .A1(n12145), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8356) );
  OAI211_X1 U10669 ( .C1(n8865), .C2(n12959), .A(n8357), .B(n8356), .ZN(n8358)
         );
  INV_X1 U10670 ( .A(n12829), .ZN(n12653) );
  XNOR2_X1 U10671 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8481) );
  NAND2_X1 U10672 ( .A1(n9024), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8493) );
  INV_X1 U10673 ( .A(n8493), .ZN(n8359) );
  NAND2_X1 U10674 ( .A1(n8481), .A2(n8359), .ZN(n8361) );
  NAND2_X1 U10675 ( .A1(n10024), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8360) );
  NAND2_X1 U10676 ( .A1(n10060), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8363) );
  NAND2_X1 U10677 ( .A1(n10018), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8362) );
  NAND2_X1 U10678 ( .A1(n8502), .A2(n8501), .ZN(n8364) );
  INV_X1 U10679 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10056) );
  NAND2_X1 U10680 ( .A1(n10039), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8365) );
  INV_X1 U10681 ( .A(n8514), .ZN(n8366) );
  NAND2_X1 U10682 ( .A1(n10020), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8368) );
  NAND2_X1 U10683 ( .A1(n10025), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8370) );
  NAND2_X1 U10684 ( .A1(n8545), .A2(n8544), .ZN(n8372) );
  NAND2_X1 U10685 ( .A1(n10040), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8373) );
  NAND2_X1 U10686 ( .A1(n10064), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8374) );
  NAND2_X1 U10687 ( .A1(n10070), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8375) );
  NAND2_X1 U10688 ( .A1(n8376), .A2(n8375), .ZN(n8571) );
  NAND2_X1 U10689 ( .A1(n10076), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8377) );
  NAND2_X1 U10690 ( .A1(n10084), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8379) );
  NAND2_X1 U10691 ( .A1(n10088), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8381) );
  NAND2_X1 U10692 ( .A1(n10228), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8383) );
  XNOR2_X1 U10693 ( .A(n10430), .B(P2_DATAO_REG_12__SCAN_IN), .ZN(n8652) );
  INV_X1 U10694 ( .A(n8652), .ZN(n8384) );
  NAND2_X1 U10695 ( .A1(n8385), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8386) );
  NAND2_X1 U10696 ( .A1(n8388), .A2(n10517), .ZN(n8389) );
  AND2_X1 U10697 ( .A1(n10685), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8391) );
  NAND2_X1 U10698 ( .A1(n10695), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8392) );
  NAND2_X1 U10699 ( .A1(n10633), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8394) );
  NAND2_X1 U10700 ( .A1(n10635), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8393) );
  NAND2_X1 U10701 ( .A1(n8394), .A2(n8393), .ZN(n8695) );
  NAND2_X1 U10702 ( .A1(n10597), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8396) );
  NAND2_X1 U10703 ( .A1(n10631), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8395) );
  NAND2_X1 U10704 ( .A1(n10637), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8398) );
  NAND2_X1 U10705 ( .A1(n10688), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8397) );
  NAND2_X1 U10706 ( .A1(n10913), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8400) );
  NAND2_X1 U10707 ( .A1(n10916), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8399) );
  INV_X1 U10708 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n12010) );
  NAND2_X1 U10709 ( .A1(n12010), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8402) );
  INV_X1 U10710 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n12129) );
  NAND2_X1 U10711 ( .A1(n12129), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8401) );
  OR2_X2 U10712 ( .A1(n8743), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8745) );
  NAND2_X1 U10713 ( .A1(n11544), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8407) );
  INV_X1 U10714 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11546) );
  NAND2_X1 U10715 ( .A1(n11546), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8406) );
  AND2_X1 U10716 ( .A1(n8407), .A2(n8406), .ZN(n8756) );
  XNOR2_X1 U10717 ( .A(n8408), .B(P1_DATAO_REG_22__SCAN_IN), .ZN(n8429) );
  NAND2_X1 U10718 ( .A1(n8409), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8410) );
  XNOR2_X1 U10719 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8770) );
  INV_X1 U10720 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8411) );
  NAND2_X1 U10721 ( .A1(n8411), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8412) );
  INV_X1 U10722 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11912) );
  NAND2_X1 U10723 ( .A1(n8414), .A2(n11912), .ZN(n8415) );
  INV_X1 U10724 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11985) );
  XNOR2_X1 U10725 ( .A(n11985), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n8417) );
  XNOR2_X1 U10726 ( .A(n8796), .B(n8417), .ZN(n11725) );
  NAND2_X1 U10727 ( .A1(n8904), .A2(n8420), .ZN(n8421) );
  NAND2_X1 U10728 ( .A1(n11725), .A2(n12159), .ZN(n8428) );
  NAND2_X1 U10729 ( .A1(n8814), .A2(SI_25_), .ZN(n8427) );
  XNOR2_X1 U10730 ( .A(n8430), .B(n8429), .ZN(n11032) );
  NAND2_X1 U10731 ( .A1(n11032), .A2(n12159), .ZN(n8432) );
  NAND2_X1 U10732 ( .A1(n8814), .A2(SI_22_), .ZN(n8431) );
  INV_X1 U10733 ( .A(n12624), .ZN(n12975) );
  NAND2_X1 U10734 ( .A1(n8766), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8433) );
  NAND2_X1 U10735 ( .A1(n8774), .A2(n8433), .ZN(n12856) );
  NAND2_X1 U10736 ( .A1(n12856), .A2(n8793), .ZN(n8439) );
  INV_X1 U10737 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n8436) );
  NAND2_X1 U10738 ( .A1(n8789), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8435) );
  NAND2_X1 U10739 ( .A1(n12145), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8434) );
  OAI211_X1 U10740 ( .C1(n8865), .C2(n8436), .A(n8435), .B(n8434), .ZN(n8437)
         );
  INV_X1 U10741 ( .A(n8437), .ZN(n8438) );
  NAND2_X1 U10742 ( .A1(n8439), .A2(n8438), .ZN(n12656) );
  INV_X1 U10743 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12732) );
  AND2_X1 U10744 ( .A1(n8468), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8440) );
  OR2_X1 U10745 ( .A1(n8440), .A2(n8749), .ZN(n12890) );
  NAND2_X1 U10746 ( .A1(n12890), .A2(n8793), .ZN(n8442) );
  AOI22_X1 U10747 ( .A1(n8830), .A2(P3_REG1_REG_19__SCAN_IN), .B1(n12145), 
        .B2(P3_REG0_REG_19__SCAN_IN), .ZN(n8441) );
  OAI211_X1 U10748 ( .C1(n8867), .C2(n12732), .A(n8442), .B(n8441), .ZN(n12659) );
  INV_X1 U10749 ( .A(n12659), .ZN(n12899) );
  OR2_X1 U10750 ( .A1(n8444), .A2(n8443), .ZN(n8445) );
  NAND2_X1 U10751 ( .A1(n8446), .A2(n8445), .ZN(n10686) );
  NAND2_X1 U10752 ( .A1(n10686), .A2(n12159), .ZN(n8457) );
  AND2_X2 U10753 ( .A1(n8530), .A2(n8546), .ZN(n8576) );
  INV_X1 U10754 ( .A(n8447), .ZN(n8448) );
  NAND2_X1 U10755 ( .A1(n8576), .A2(n8448), .ZN(n8654) );
  NOR2_X2 U10756 ( .A1(n8666), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n8682) );
  NAND2_X1 U10757 ( .A1(n8682), .A2(n8684), .ZN(n8699) );
  INV_X1 U10758 ( .A(n8699), .ZN(n8451) );
  INV_X1 U10759 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8452) );
  NOR2_X1 U10760 ( .A1(n8529), .A2(SI_19_), .ZN(n8455) );
  AOI21_X1 U10761 ( .B1(n8454), .B2(n6475), .A(n8455), .ZN(n8456) );
  OR2_X1 U10762 ( .A1(n8459), .A2(n8458), .ZN(n8460) );
  NAND2_X1 U10763 ( .A1(n8461), .A2(n8460), .ZN(n10574) );
  NAND2_X1 U10764 ( .A1(n8462), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8463) );
  XNOR2_X1 U10765 ( .A(n8463), .B(P3_IR_REG_18__SCAN_IN), .ZN(n14380) );
  NOR2_X1 U10766 ( .A1(n8529), .A2(n15252), .ZN(n8464) );
  AOI21_X1 U10767 ( .B1(n14380), .B2(n6474), .A(n8464), .ZN(n8465) );
  INV_X1 U10768 ( .A(n12635), .ZN(n13051) );
  INV_X1 U10769 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n8471) );
  AOI22_X1 U10770 ( .A1(n8830), .A2(P3_REG1_REG_18__SCAN_IN), .B1(n12145), 
        .B2(P3_REG0_REG_18__SCAN_IN), .ZN(n8470) );
  NAND2_X1 U10771 ( .A1(n8737), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8467) );
  NAND2_X1 U10772 ( .A1(n8468), .A2(n8467), .ZN(n12904) );
  NAND2_X1 U10773 ( .A1(n12904), .A2(n8793), .ZN(n8469) );
  OAI211_X1 U10774 ( .C1(n12148), .C2(n8471), .A(n8470), .B(n8469), .ZN(n12886) );
  INV_X1 U10775 ( .A(n12886), .ZN(n12911) );
  INV_X1 U10776 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10726) );
  INV_X1 U10777 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10745) );
  NAND2_X1 U10778 ( .A1(n8509), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8475) );
  INV_X1 U10779 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n15113) );
  NAND4_X1 U10780 ( .A1(n8477), .A2(n8476), .A3(n8475), .A4(n8474), .ZN(n9759)
         );
  INV_X1 U10781 ( .A(n8478), .ZN(n8479) );
  XNOR2_X1 U10782 ( .A(n8493), .B(n8481), .ZN(n10067) );
  NOR2_X1 U10783 ( .A1(n10067), .A2(n6720), .ZN(n8483) );
  NAND2_X1 U10784 ( .A1(n8483), .A2(n8482), .ZN(n8484) );
  INV_X1 U10785 ( .A(n8498), .ZN(n10676) );
  NAND2_X1 U10786 ( .A1(n12217), .A2(n8874), .ZN(n15105) );
  INV_X1 U10787 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10731) );
  INV_X1 U10788 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n8486) );
  OR2_X1 U10789 ( .A1(n8510), .A2(n8486), .ZN(n8489) );
  NAND2_X1 U10790 ( .A1(n8509), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8488) );
  INV_X1 U10791 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10730) );
  OR2_X1 U10792 ( .A1(n8778), .A2(n10730), .ZN(n8487) );
  NAND2_X1 U10793 ( .A1(n8491), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8492) );
  NAND2_X1 U10794 ( .A1(n8493), .A2(n8492), .ZN(n10033) );
  NAND2_X1 U10795 ( .A1(n12159), .A2(n10033), .ZN(n8496) );
  OR2_X1 U10796 ( .A1(n8529), .A2(n10034), .ZN(n8495) );
  NAND2_X1 U10797 ( .A1(n6474), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n8494) );
  NAND2_X1 U10798 ( .A1(n15105), .A2(n9767), .ZN(n8500) );
  OR2_X1 U10799 ( .A1(n8498), .A2(n9759), .ZN(n8499) );
  XNOR2_X1 U10800 ( .A(n8502), .B(n8501), .ZN(n10028) );
  OR2_X1 U10801 ( .A1(n8478), .A2(n8612), .ZN(n8504) );
  NAND2_X1 U10802 ( .A1(n6475), .A2(n10834), .ZN(n8505) );
  NAND2_X1 U10803 ( .A1(n8509), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8507) );
  INV_X1 U10804 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15226) );
  OR2_X1 U10805 ( .A1(n8510), .A2(n15226), .ZN(n8506) );
  INV_X1 U10806 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10766) );
  INV_X1 U10807 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10765) );
  NAND2_X1 U10808 ( .A1(n15094), .A2(n15093), .ZN(n15092) );
  INV_X1 U10809 ( .A(n15088), .ZN(n10783) );
  OR2_X1 U10810 ( .A1(n9772), .A2(n10783), .ZN(n8508) );
  NAND2_X1 U10811 ( .A1(n8509), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8513) );
  INV_X1 U10812 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10807) );
  INV_X1 U10813 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10806) );
  OR2_X1 U10814 ( .A1(n8778), .A2(n10806), .ZN(n8511) );
  XNOR2_X1 U10815 ( .A(n8515), .B(n8514), .ZN(n10027) );
  NAND2_X1 U10816 ( .A1(n12159), .A2(n10027), .ZN(n8520) );
  INV_X1 U10817 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8517) );
  XNOR2_X1 U10818 ( .A(n8518), .B(n8517), .ZN(n14976) );
  NAND2_X1 U10819 ( .A1(n6474), .A2(n14976), .ZN(n8519) );
  NAND2_X1 U10820 ( .A1(n15091), .A2(n15129), .ZN(n12226) );
  NAND2_X1 U10821 ( .A1(n15091), .A2(n6803), .ZN(n8521) );
  NAND2_X1 U10822 ( .A1(n12145), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8526) );
  INV_X1 U10823 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10822) );
  OR2_X1 U10824 ( .A1(n12148), .A2(n10822), .ZN(n8525) );
  AND2_X1 U10825 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8522) );
  NOR2_X1 U10826 ( .A1(n8538), .A2(n8522), .ZN(n11041) );
  OR2_X1 U10827 ( .A1(n8510), .A2(n11041), .ZN(n8524) );
  INV_X1 U10828 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10841) );
  OR2_X1 U10829 ( .A1(n8778), .A2(n10841), .ZN(n8523) );
  XNOR2_X1 U10830 ( .A(n8528), .B(n8527), .ZN(n10031) );
  OR2_X1 U10831 ( .A1(n8529), .A2(SI_4_), .ZN(n8536) );
  INV_X1 U10832 ( .A(n8530), .ZN(n8534) );
  MUX2_X1 U10833 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8532), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n8533) );
  NAND2_X1 U10834 ( .A1(n8534), .A2(n8533), .ZN(n15005) );
  NAND2_X1 U10835 ( .A1(n6474), .A2(n15005), .ZN(n8535) );
  OAI211_X1 U10836 ( .C1(n8760), .C2(n10031), .A(n8536), .B(n8535), .ZN(n15134) );
  NAND2_X1 U10837 ( .A1(n12673), .A2(n15134), .ZN(n12236) );
  INV_X1 U10838 ( .A(n15134), .ZN(n8537) );
  NAND2_X1 U10839 ( .A1(n12145), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8543) );
  INV_X1 U10840 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n10815) );
  OR2_X1 U10841 ( .A1(n8778), .A2(n10815), .ZN(n8542) );
  OR2_X1 U10842 ( .A1(n15288), .A2(n8538), .ZN(n8539) );
  AND2_X1 U10843 ( .A1(n8552), .A2(n8539), .ZN(n11127) );
  OR2_X1 U10844 ( .A1(n8510), .A2(n11127), .ZN(n8541) );
  INV_X1 U10845 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10816) );
  OR2_X1 U10846 ( .A1(n12148), .A2(n10816), .ZN(n8540) );
  NAND4_X1 U10847 ( .A1(n8543), .A2(n8542), .A3(n8541), .A4(n8540), .ZN(n12672) );
  XNOR2_X1 U10848 ( .A(n8545), .B(n8544), .ZN(n10050) );
  OR2_X1 U10849 ( .A1(n8529), .A2(SI_5_), .ZN(n8549) );
  OR2_X1 U10850 ( .A1(n8530), .A2(n8612), .ZN(n8547) );
  XNOR2_X1 U10851 ( .A(n8547), .B(n8546), .ZN(n15023) );
  NAND2_X1 U10852 ( .A1(n6475), .A2(n15023), .ZN(n8548) );
  OAI211_X1 U10853 ( .C1(n8760), .C2(n10050), .A(n8549), .B(n8548), .ZN(n15139) );
  OR2_X1 U10854 ( .A1(n12672), .A2(n15139), .ZN(n12242) );
  NAND2_X1 U10855 ( .A1(n12672), .A2(n15139), .ZN(n12233) );
  NAND2_X1 U10856 ( .A1(n12242), .A2(n12233), .ZN(n11130) );
  NAND2_X1 U10857 ( .A1(n11128), .A2(n11130), .ZN(n11129) );
  INV_X1 U10858 ( .A(n15139), .ZN(n8550) );
  OR2_X1 U10859 ( .A1(n12672), .A2(n8550), .ZN(n8551) );
  NAND2_X1 U10860 ( .A1(n12145), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8557) );
  INV_X1 U10861 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n10826) );
  OR2_X1 U10862 ( .A1(n12148), .A2(n10826), .ZN(n8556) );
  NAND2_X1 U10863 ( .A1(n8552), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8553) );
  AND2_X1 U10864 ( .A1(n8565), .A2(n8553), .ZN(n11188) );
  OR2_X1 U10865 ( .A1(n8510), .A2(n11188), .ZN(n8555) );
  INV_X1 U10866 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n10845) );
  OR2_X1 U10867 ( .A1(n8865), .A2(n10845), .ZN(n8554) );
  NAND4_X1 U10868 ( .A1(n8557), .A2(n8556), .A3(n8555), .A4(n8554), .ZN(n12671) );
  INV_X1 U10869 ( .A(SI_6_), .ZN(n15331) );
  XNOR2_X1 U10870 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n8558) );
  XNOR2_X1 U10871 ( .A(n8559), .B(n8558), .ZN(n10036) );
  NAND2_X1 U10872 ( .A1(n12159), .A2(n10036), .ZN(n8562) );
  OR2_X1 U10873 ( .A1(n8576), .A2(n8612), .ZN(n8560) );
  NAND2_X1 U10874 ( .A1(n6474), .A2(n10858), .ZN(n8561) );
  OAI211_X1 U10875 ( .C1(n8529), .C2(n15331), .A(n8562), .B(n8561), .ZN(n9780)
         );
  INV_X1 U10876 ( .A(n9780), .ZN(n15144) );
  NAND2_X1 U10877 ( .A1(n12671), .A2(n15144), .ZN(n12243) );
  NAND2_X1 U10878 ( .A1(n12244), .A2(n12243), .ZN(n11185) );
  INV_X1 U10879 ( .A(n11185), .ZN(n12174) );
  NAND2_X1 U10880 ( .A1(n12671), .A2(n9780), .ZN(n8563) );
  NAND2_X1 U10881 ( .A1(n12145), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8570) );
  INV_X1 U10882 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n8564) );
  OR2_X1 U10883 ( .A1(n8778), .A2(n8564), .ZN(n8569) );
  AND2_X1 U10884 ( .A1(n8565), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8566) );
  NOR2_X1 U10885 ( .A1(n8582), .A2(n8566), .ZN(n11415) );
  OR2_X1 U10886 ( .A1(n8510), .A2(n11415), .ZN(n8568) );
  INV_X1 U10887 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11414) );
  OR2_X1 U10888 ( .A1(n8867), .A2(n11414), .ZN(n8567) );
  NAND4_X1 U10889 ( .A1(n8570), .A2(n8569), .A3(n8568), .A4(n8567), .ZN(n12670) );
  NAND2_X1 U10890 ( .A1(n8572), .A2(n8571), .ZN(n8573) );
  NAND2_X1 U10891 ( .A1(n8574), .A2(n8573), .ZN(n10048) );
  NAND2_X1 U10892 ( .A1(n12159), .A2(n10048), .ZN(n8581) );
  OR2_X1 U10893 ( .A1(n8529), .A2(SI_7_), .ZN(n8580) );
  INV_X1 U10894 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8575) );
  NAND2_X1 U10895 ( .A1(n8576), .A2(n8575), .ZN(n8592) );
  NAND2_X1 U10896 ( .A1(n8592), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8578) );
  INV_X1 U10897 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8577) );
  XNOR2_X1 U10898 ( .A(n8578), .B(n8577), .ZN(n15035) );
  NAND2_X1 U10899 ( .A1(n6474), .A2(n15035), .ZN(n8579) );
  INV_X1 U10900 ( .A(n11328), .ZN(n8600) );
  NAND2_X1 U10901 ( .A1(n12145), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8587) );
  NOR2_X1 U10902 ( .A1(n8582), .A2(n15301), .ZN(n8583) );
  OR2_X1 U10903 ( .A1(n8510), .A2(n6624), .ZN(n8586) );
  INV_X1 U10904 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10870) );
  OR2_X1 U10905 ( .A1(n12148), .A2(n10870), .ZN(n8585) );
  INV_X1 U10906 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n10862) );
  OR2_X1 U10907 ( .A1(n8865), .A2(n10862), .ZN(n8584) );
  NAND4_X1 U10908 ( .A1(n8587), .A2(n8586), .A3(n8585), .A4(n8584), .ZN(n12669) );
  INV_X1 U10909 ( .A(SI_8_), .ZN(n15379) );
  OR2_X1 U10910 ( .A1(n8589), .A2(n8588), .ZN(n8590) );
  NAND2_X1 U10911 ( .A1(n8591), .A2(n8590), .ZN(n10053) );
  OR2_X1 U10912 ( .A1(n8760), .A2(n10053), .ZN(n8598) );
  INV_X1 U10913 ( .A(n8629), .ZN(n8596) );
  NAND2_X1 U10914 ( .A1(n8593), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8594) );
  MUX2_X1 U10915 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8594), .S(
        P3_IR_REG_8__SCAN_IN), .Z(n8595) );
  NAND2_X1 U10916 ( .A1(n6475), .A2(n11383), .ZN(n8597) );
  OAI211_X1 U10917 ( .C1(n8529), .C2(n15379), .A(n8598), .B(n8597), .ZN(n9786)
         );
  NOR2_X1 U10918 ( .A1(n12669), .A2(n9786), .ZN(n8599) );
  AOI21_X1 U10919 ( .B1(n8600), .B2(n6504), .A(n8599), .ZN(n11440) );
  NAND2_X1 U10920 ( .A1(n12145), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8607) );
  INV_X1 U10921 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15185) );
  OR2_X1 U10922 ( .A1(n8778), .A2(n15185), .ZN(n8606) );
  OR2_X1 U10923 ( .A1(n8602), .A2(n8601), .ZN(n8603) );
  AND2_X1 U10924 ( .A1(n8618), .A2(n8603), .ZN(n11519) );
  OR2_X1 U10925 ( .A1(n8510), .A2(n11519), .ZN(n8605) );
  INV_X1 U10926 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n15047) );
  OR2_X1 U10927 ( .A1(n8867), .A2(n15047), .ZN(n8604) );
  NAND4_X1 U10928 ( .A1(n8607), .A2(n8606), .A3(n8605), .A4(n8604), .ZN(n12668) );
  OR2_X1 U10929 ( .A1(n8609), .A2(n8608), .ZN(n8610) );
  NAND2_X1 U10930 ( .A1(n8611), .A2(n8610), .ZN(n10049) );
  NAND2_X1 U10931 ( .A1(n12159), .A2(n10049), .ZN(n8615) );
  OR2_X1 U10932 ( .A1(n8629), .A2(n8612), .ZN(n8613) );
  INV_X1 U10933 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8628) );
  XNOR2_X1 U10934 ( .A(n8613), .B(n8628), .ZN(n15053) );
  NAND2_X1 U10935 ( .A1(n6474), .A2(n15053), .ZN(n8614) );
  OAI211_X1 U10936 ( .C1(n8529), .C2(SI_9_), .A(n8615), .B(n8614), .ZN(n15161)
         );
  INV_X1 U10937 ( .A(n15161), .ZN(n11516) );
  XNOR2_X1 U10938 ( .A(n12668), .B(n11516), .ZN(n12257) );
  NAND2_X1 U10939 ( .A1(n11440), .A2(n8616), .ZN(n11439) );
  NAND2_X1 U10940 ( .A1(n12668), .A2(n11516), .ZN(n8617) );
  NAND2_X1 U10941 ( .A1(n11439), .A2(n8617), .ZN(n11538) );
  NAND2_X1 U10942 ( .A1(n12145), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8623) );
  INV_X1 U10943 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11387) );
  OR2_X1 U10944 ( .A1(n8865), .A2(n11387), .ZN(n8622) );
  NAND2_X1 U10945 ( .A1(n8618), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8619) );
  AND2_X1 U10946 ( .A1(n8643), .A2(n8619), .ZN(n11588) );
  OR2_X1 U10947 ( .A1(n8510), .A2(n11588), .ZN(n8621) );
  INV_X1 U10948 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11388) );
  OR2_X1 U10949 ( .A1(n12148), .A2(n11388), .ZN(n8620) );
  NAND4_X1 U10950 ( .A1(n8623), .A2(n8622), .A3(n8621), .A4(n8620), .ZN(n12667) );
  OR2_X1 U10951 ( .A1(n8625), .A2(n8624), .ZN(n8626) );
  NAND2_X1 U10952 ( .A1(n8627), .A2(n8626), .ZN(n10041) );
  NAND2_X1 U10953 ( .A1(n10041), .A2(n12159), .ZN(n8634) );
  INV_X1 U10954 ( .A(SI_10_), .ZN(n15248) );
  NAND2_X1 U10955 ( .A1(n8629), .A2(n8628), .ZN(n8638) );
  NAND2_X1 U10956 ( .A1(n8638), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8631) );
  INV_X1 U10957 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8630) );
  XNOR2_X1 U10958 ( .A(n8631), .B(n8630), .ZN(n11390) );
  AOI22_X1 U10959 ( .A1(n8814), .A2(n15248), .B1(n6474), .B2(n11390), .ZN(
        n8633) );
  NAND2_X1 U10960 ( .A1(n8634), .A2(n8633), .ZN(n15167) );
  OR2_X1 U10961 ( .A1(n12667), .A2(n15167), .ZN(n12270) );
  NAND2_X1 U10962 ( .A1(n12667), .A2(n15167), .ZN(n12263) );
  NAND2_X1 U10963 ( .A1(n12270), .A2(n12263), .ZN(n12171) );
  INV_X1 U10964 ( .A(n15167), .ZN(n11583) );
  NAND2_X1 U10965 ( .A1(n11583), .A2(n12667), .ZN(n8635) );
  NAND2_X1 U10966 ( .A1(n11537), .A2(n8635), .ZN(n11715) );
  XNOR2_X1 U10967 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8636) );
  XNOR2_X1 U10968 ( .A(n8637), .B(n8636), .ZN(n10054) );
  NAND2_X1 U10969 ( .A1(n10054), .A2(n12159), .ZN(n8642) );
  INV_X1 U10970 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8639) );
  XNOR2_X1 U10971 ( .A(n8640), .B(n8639), .ZN(n11556) );
  AOI22_X1 U10972 ( .A1(n8814), .A2(n15315), .B1(n6475), .B2(n11556), .ZN(
        n8641) );
  NAND2_X1 U10973 ( .A1(n8642), .A2(n8641), .ZN(n11836) );
  NAND2_X1 U10974 ( .A1(n12145), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8648) );
  INV_X1 U10975 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n11394) );
  OR2_X1 U10976 ( .A1(n8865), .A2(n11394), .ZN(n8647) );
  NAND2_X1 U10977 ( .A1(n8643), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8644) );
  AND2_X1 U10978 ( .A1(n8659), .A2(n8644), .ZN(n14399) );
  OR2_X1 U10979 ( .A1(n8510), .A2(n14399), .ZN(n8646) );
  INV_X1 U10980 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11395) );
  OR2_X1 U10981 ( .A1(n12148), .A2(n11395), .ZN(n8645) );
  NAND2_X1 U10982 ( .A1(n11715), .A2(n8649), .ZN(n8651) );
  OR2_X1 U10983 ( .A1(n11836), .A2(n11834), .ZN(n8650) );
  NAND2_X1 U10984 ( .A1(n8651), .A2(n8650), .ZN(n11760) );
  XNOR2_X1 U10985 ( .A(n8653), .B(n8652), .ZN(n10074) );
  NAND2_X1 U10986 ( .A1(n10074), .A2(n12159), .ZN(n8658) );
  NAND2_X1 U10987 ( .A1(n8654), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8655) );
  MUX2_X1 U10988 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8655), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n8656) );
  AND2_X1 U10989 ( .A1(n8656), .A2(n8666), .ZN(n11791) );
  AOI22_X1 U10990 ( .A1(n8814), .A2(SI_12_), .B1(n6475), .B2(n11791), .ZN(
        n8657) );
  NAND2_X1 U10991 ( .A1(n8658), .A2(n8657), .ZN(n12281) );
  NAND2_X1 U10992 ( .A1(n12145), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8664) );
  INV_X1 U10993 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11767) );
  OR2_X1 U10994 ( .A1(n8867), .A2(n11767), .ZN(n8663) );
  AND2_X1 U10995 ( .A1(n8659), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8660) );
  NOR2_X1 U10996 ( .A1(n8672), .A2(n8660), .ZN(n11888) );
  OR2_X1 U10997 ( .A1(n8510), .A2(n11888), .ZN(n8662) );
  INV_X1 U10998 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n11559) );
  OR2_X1 U10999 ( .A1(n8778), .A2(n11559), .ZN(n8661) );
  NAND4_X1 U11000 ( .A1(n8664), .A2(n8663), .A3(n8662), .A4(n8661), .ZN(n12665) );
  OR2_X1 U11001 ( .A1(n12281), .A2(n12280), .ZN(n12264) );
  NAND2_X1 U11002 ( .A1(n12281), .A2(n12280), .ZN(n12274) );
  NAND2_X1 U11003 ( .A1(n12264), .A2(n12274), .ZN(n12182) );
  XNOR2_X1 U11004 ( .A(n8665), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n10086) );
  NAND2_X1 U11005 ( .A1(n10086), .A2(n12159), .ZN(n8670) );
  INV_X1 U11006 ( .A(SI_13_), .ZN(n15261) );
  NAND2_X1 U11007 ( .A1(n8666), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8668) );
  INV_X1 U11008 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8667) );
  XNOR2_X1 U11009 ( .A(n8668), .B(n8667), .ZN(n12680) );
  AOI22_X1 U11010 ( .A1(n8814), .A2(n15261), .B1(n6474), .B2(n12680), .ZN(
        n8669) );
  NAND2_X1 U11011 ( .A1(n8670), .A2(n8669), .ZN(n14407) );
  INV_X1 U11012 ( .A(n14407), .ZN(n11932) );
  NAND2_X1 U11013 ( .A1(n12145), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8678) );
  INV_X1 U11014 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n8671) );
  OR2_X1 U11015 ( .A1(n8865), .A2(n8671), .ZN(n8677) );
  OR2_X1 U11016 ( .A1(n8672), .A2(n11927), .ZN(n8673) );
  AND2_X1 U11017 ( .A1(n8673), .A2(n8688), .ZN(n11930) );
  OR2_X1 U11018 ( .A1(n8510), .A2(n11930), .ZN(n8676) );
  INV_X1 U11019 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n8674) );
  OR2_X1 U11020 ( .A1(n12148), .A2(n8674), .ZN(n8675) );
  NAND4_X1 U11021 ( .A1(n8678), .A2(n8677), .A3(n8676), .A4(n8675), .ZN(n12664) );
  NAND2_X1 U11022 ( .A1(n11932), .A2(n12664), .ZN(n8679) );
  INV_X1 U11023 ( .A(n12664), .ZN(n11762) );
  XNOR2_X1 U11024 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n8680) );
  XNOR2_X1 U11025 ( .A(n8681), .B(n8680), .ZN(n10097) );
  NAND2_X1 U11026 ( .A1(n10097), .A2(n12159), .ZN(n8687) );
  INV_X1 U11027 ( .A(n8682), .ZN(n8683) );
  NAND2_X1 U11028 ( .A1(n8683), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8685) );
  XNOR2_X1 U11029 ( .A(n8685), .B(n8684), .ZN(n12700) );
  AOI22_X1 U11030 ( .A1(n8814), .A2(n15263), .B1(n6475), .B2(n12700), .ZN(
        n8686) );
  NAND2_X1 U11031 ( .A1(n8830), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8694) );
  INV_X1 U11032 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n11937) );
  OR2_X1 U11033 ( .A1(n8831), .A2(n11937), .ZN(n8693) );
  NAND2_X1 U11034 ( .A1(n8688), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8689) );
  AND2_X1 U11035 ( .A1(n8705), .A2(n8689), .ZN(n12549) );
  OR2_X1 U11036 ( .A1(n8510), .A2(n12549), .ZN(n8692) );
  INV_X1 U11037 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n8690) );
  OR2_X1 U11038 ( .A1(n12148), .A2(n8690), .ZN(n8691) );
  NAND4_X1 U11039 ( .A1(n8694), .A2(n8693), .A3(n8692), .A4(n8691), .ZN(n12663) );
  XNOR2_X1 U11040 ( .A(n12555), .B(n12663), .ZN(n12287) );
  INV_X1 U11041 ( .A(n12663), .ZN(n11916) );
  NAND2_X1 U11042 ( .A1(n8696), .A2(n8695), .ZN(n8697) );
  NAND2_X1 U11043 ( .A1(n8698), .A2(n8697), .ZN(n10310) );
  OR2_X1 U11044 ( .A1(n10310), .A2(n8760), .ZN(n8703) );
  XNOR2_X1 U11045 ( .A(n8701), .B(n8700), .ZN(n12750) );
  INV_X1 U11046 ( .A(n12750), .ZN(n12735) );
  AOI22_X1 U11047 ( .A1(n8814), .A2(SI_15_), .B1(n6474), .B2(n12735), .ZN(
        n8702) );
  NAND2_X1 U11048 ( .A1(n8703), .A2(n8702), .ZN(n12118) );
  NAND2_X1 U11049 ( .A1(n8830), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8710) );
  INV_X1 U11050 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n8704) );
  OR2_X1 U11051 ( .A1(n8831), .A2(n8704), .ZN(n8709) );
  AND2_X1 U11052 ( .A1(n8705), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8706) );
  NOR2_X1 U11053 ( .A1(n8721), .A2(n8706), .ZN(n12116) );
  OR2_X1 U11054 ( .A1(n8510), .A2(n12116), .ZN(n8708) );
  INV_X1 U11055 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12707) );
  OR2_X1 U11056 ( .A1(n8867), .A2(n12707), .ZN(n8707) );
  NAND4_X1 U11057 ( .A1(n8710), .A2(n8709), .A3(n8708), .A4(n8707), .ZN(n12662) );
  INV_X1 U11058 ( .A(n12118), .ZN(n13007) );
  OR2_X1 U11059 ( .A1(n8712), .A2(n8711), .ZN(n8713) );
  NAND2_X1 U11060 ( .A1(n8714), .A2(n8713), .ZN(n10429) );
  NAND2_X1 U11061 ( .A1(n8715), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8716) );
  MUX2_X1 U11062 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8716), .S(
        P3_IR_REG_16__SCAN_IN), .Z(n8718) );
  INV_X1 U11063 ( .A(n8717), .ZN(n8731) );
  AND2_X1 U11064 ( .A1(n8718), .A2(n8731), .ZN(n14347) );
  AOI22_X1 U11065 ( .A1(n8814), .A2(SI_16_), .B1(n14347), .B2(n6474), .ZN(
        n8719) );
  NOR2_X1 U11066 ( .A1(n8721), .A2(n15330), .ZN(n8722) );
  OR2_X1 U11067 ( .A1(n8735), .A2(n8722), .ZN(n12931) );
  NAND2_X1 U11068 ( .A1(n8793), .A2(n12931), .ZN(n8726) );
  INV_X1 U11069 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13001) );
  OR2_X1 U11070 ( .A1(n8778), .A2(n13001), .ZN(n8725) );
  INV_X1 U11071 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13057) );
  OR2_X1 U11072 ( .A1(n8831), .A2(n13057), .ZN(n8724) );
  INV_X1 U11073 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12727) );
  OR2_X1 U11074 ( .A1(n8867), .A2(n12727), .ZN(n8723) );
  NAND4_X1 U11075 ( .A1(n8726), .A2(n8725), .A3(n8724), .A4(n8723), .ZN(n12661) );
  OR2_X1 U11076 ( .A1(n12930), .A2(n12912), .ZN(n12292) );
  NAND2_X1 U11077 ( .A1(n12930), .A2(n12912), .ZN(n12304) );
  NAND2_X1 U11078 ( .A1(n12292), .A2(n12304), .ZN(n12921) );
  OR2_X1 U11079 ( .A1(n8728), .A2(n8727), .ZN(n8729) );
  NAND2_X1 U11080 ( .A1(n8730), .A2(n8729), .ZN(n10518) );
  NAND2_X1 U11081 ( .A1(n8731), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8732) );
  XNOR2_X1 U11082 ( .A(n8732), .B(P3_IR_REG_17__SCAN_IN), .ZN(n14365) );
  AOI22_X1 U11083 ( .A1(SI_17_), .A2(n8814), .B1(n14365), .B2(n6475), .ZN(
        n8733) );
  NAND2_X1 U11084 ( .A1(n8734), .A2(n8733), .ZN(n12598) );
  OR2_X1 U11085 ( .A1(n8735), .A2(n15282), .ZN(n8736) );
  NAND2_X1 U11086 ( .A1(n8737), .A2(n8736), .ZN(n12915) );
  NAND2_X1 U11087 ( .A1(n12915), .A2(n8793), .ZN(n8742) );
  INV_X1 U11088 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12997) );
  OR2_X1 U11089 ( .A1(n8865), .A2(n12997), .ZN(n8741) );
  NAND2_X1 U11090 ( .A1(n12145), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8740) );
  INV_X1 U11091 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n8738) );
  OR2_X1 U11092 ( .A1(n12148), .A2(n8738), .ZN(n8739) );
  NAND4_X1 U11093 ( .A1(n8742), .A2(n8741), .A3(n8740), .A4(n8739), .ZN(n12660) );
  OR2_X1 U11094 ( .A1(n12598), .A2(n12924), .ZN(n12312) );
  NAND2_X1 U11095 ( .A1(n12598), .A2(n12924), .ZN(n12314) );
  INV_X1 U11096 ( .A(n12598), .ZN(n13055) );
  NAND2_X1 U11097 ( .A1(n12635), .A2(n12911), .ZN(n12316) );
  OR2_X1 U11098 ( .A1(n13047), .A2(n12659), .ZN(n12320) );
  NAND2_X1 U11099 ( .A1(n13047), .A2(n12659), .ZN(n12321) );
  NAND2_X1 U11100 ( .A1(n12320), .A2(n12321), .ZN(n12885) );
  NAND2_X1 U11101 ( .A1(n8743), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8744) );
  NAND2_X1 U11102 ( .A1(n8745), .A2(n8744), .ZN(n10880) );
  NAND2_X1 U11103 ( .A1(n8814), .A2(SI_20_), .ZN(n8746) );
  NOR2_X1 U11104 ( .A1(n8749), .A2(n8748), .ZN(n8750) );
  OR2_X1 U11105 ( .A1(n8764), .A2(n8750), .ZN(n12878) );
  NAND2_X1 U11106 ( .A1(n12878), .A2(n8793), .ZN(n8755) );
  INV_X1 U11107 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12982) );
  NAND2_X1 U11108 ( .A1(n8789), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8752) );
  NAND2_X1 U11109 ( .A1(n12145), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8751) );
  OAI211_X1 U11110 ( .C1(n8865), .C2(n12982), .A(n8752), .B(n8751), .ZN(n8753)
         );
  INV_X1 U11111 ( .A(n8753), .ZN(n8754) );
  XNOR2_X1 U11112 ( .A(n12877), .B(n12862), .ZN(n12871) );
  AOI22_X1 U11113 ( .A1(n12872), .A2(n12871), .B1(n12887), .B2(n12877), .ZN(
        n12860) );
  OR2_X1 U11114 ( .A1(n8757), .A2(n8756), .ZN(n8758) );
  NAND2_X1 U11115 ( .A1(n8759), .A2(n8758), .ZN(n11004) );
  NAND2_X1 U11116 ( .A1(n8814), .A2(SI_21_), .ZN(n8761) );
  OR2_X1 U11117 ( .A1(n8764), .A2(n8763), .ZN(n8765) );
  NAND2_X1 U11118 ( .A1(n8766), .A2(n8765), .ZN(n12866) );
  INV_X1 U11119 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12978) );
  NAND2_X1 U11120 ( .A1(n8789), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8768) );
  NAND2_X1 U11121 ( .A1(n12145), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8767) );
  OAI211_X1 U11122 ( .C1(n8865), .C2(n12978), .A(n8768), .B(n8767), .ZN(n8769)
         );
  INV_X1 U11123 ( .A(n12874), .ZN(n12657) );
  NAND2_X1 U11124 ( .A1(n12865), .A2(n12657), .ZN(n12167) );
  NOR2_X1 U11125 ( .A1(n12865), .A2(n12657), .ZN(n12169) );
  XNOR2_X1 U11126 ( .A(n8771), .B(n8770), .ZN(n11309) );
  NAND2_X1 U11127 ( .A1(n11309), .A2(n12159), .ZN(n8773) );
  NAND2_X1 U11128 ( .A1(n8814), .A2(SI_23_), .ZN(n8772) );
  AND2_X1 U11129 ( .A1(n8774), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8775) );
  OR2_X1 U11130 ( .A1(n8775), .A2(n8786), .ZN(n12846) );
  NAND2_X1 U11131 ( .A1(n12846), .A2(n8793), .ZN(n8781) );
  INV_X1 U11132 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12970) );
  NAND2_X1 U11133 ( .A1(n8789), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8777) );
  NAND2_X1 U11134 ( .A1(n12145), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8776) );
  OAI211_X1 U11135 ( .C1(n8778), .C2(n12970), .A(n8777), .B(n8776), .ZN(n8779)
         );
  INV_X1 U11136 ( .A(n8779), .ZN(n8780) );
  NAND2_X1 U11137 ( .A1(n8781), .A2(n8780), .ZN(n12655) );
  NAND2_X1 U11138 ( .A1(n12966), .A2(n12828), .ZN(n8782) );
  NAND2_X1 U11139 ( .A1(n12341), .A2(n8782), .ZN(n12336) );
  XNOR2_X1 U11140 ( .A(n8783), .B(n11880), .ZN(n11577) );
  NAND2_X1 U11141 ( .A1(n11577), .A2(n12159), .ZN(n8785) );
  NAND2_X1 U11142 ( .A1(n8814), .A2(SI_24_), .ZN(n8784) );
  OR2_X1 U11143 ( .A1(n8786), .A2(n12607), .ZN(n8787) );
  NAND2_X1 U11144 ( .A1(n8788), .A2(n8787), .ZN(n12833) );
  INV_X1 U11145 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12964) );
  NAND2_X1 U11146 ( .A1(n8789), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8791) );
  NAND2_X1 U11147 ( .A1(n12145), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8790) );
  OAI211_X1 U11148 ( .C1(n8865), .C2(n12964), .A(n8791), .B(n8790), .ZN(n8792)
         );
  OR2_X1 U11149 ( .A1(n12834), .A2(n12842), .ZN(n12343) );
  NAND2_X1 U11150 ( .A1(n12834), .A2(n12842), .ZN(n12346) );
  NAND2_X1 U11151 ( .A1(n12343), .A2(n12346), .ZN(n12826) );
  INV_X1 U11152 ( .A(n12842), .ZN(n12654) );
  NAND2_X1 U11153 ( .A1(n12578), .A2(n12829), .ZN(n12350) );
  NAND2_X1 U11154 ( .A1(n11985), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8795) );
  NAND2_X1 U11155 ( .A1(n11990), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8797) );
  INV_X1 U11156 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13653) );
  XNOR2_X1 U11157 ( .A(n13653), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n8799) );
  XNOR2_X1 U11158 ( .A(n8811), .B(n8799), .ZN(n11776) );
  NAND2_X1 U11159 ( .A1(n11776), .A2(n12159), .ZN(n8801) );
  NAND2_X1 U11160 ( .A1(n8814), .A2(SI_26_), .ZN(n8800) );
  NAND2_X1 U11161 ( .A1(n8830), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8807) );
  INV_X1 U11162 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13020) );
  OR2_X1 U11163 ( .A1(n8831), .A2(n13020), .ZN(n8806) );
  INV_X1 U11164 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n15325) );
  NAND2_X1 U11165 ( .A1(n15325), .A2(n8802), .ZN(n8819) );
  INV_X1 U11166 ( .A(n8819), .ZN(n8818) );
  AOI21_X1 U11167 ( .B1(P3_REG3_REG_26__SCAN_IN), .B2(n8803), .A(n8818), .ZN(
        n12802) );
  OR2_X1 U11168 ( .A1(n8510), .A2(n12802), .ZN(n8805) );
  INV_X1 U11169 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n12803) );
  OR2_X1 U11170 ( .A1(n8867), .A2(n12803), .ZN(n8804) );
  NAND4_X1 U11171 ( .A1(n8807), .A2(n8806), .A3(n8805), .A4(n8804), .ZN(n12652) );
  NAND2_X1 U11172 ( .A1(n13022), .A2(n12811), .ZN(n8808) );
  AND2_X1 U11173 ( .A1(n14211), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8810) );
  NAND2_X1 U11174 ( .A1(n13653), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8812) );
  XNOR2_X1 U11175 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n8813) );
  XNOR2_X1 U11176 ( .A(n8826), .B(n8813), .ZN(n11831) );
  NAND2_X1 U11177 ( .A1(n11831), .A2(n12159), .ZN(n8816) );
  NAND2_X1 U11178 ( .A1(n8814), .A2(SI_27_), .ZN(n8815) );
  NAND2_X1 U11179 ( .A1(n8830), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8824) );
  INV_X1 U11180 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n8817) );
  OR2_X1 U11181 ( .A1(n8831), .A2(n8817), .ZN(n8823) );
  INV_X1 U11182 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n15303) );
  NAND2_X1 U11183 ( .A1(n15303), .A2(n8818), .ZN(n8834) );
  NAND2_X1 U11184 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(n8819), .ZN(n8820) );
  INV_X1 U11185 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n12792) );
  OR2_X1 U11186 ( .A1(n12148), .A2(n12792), .ZN(n8821) );
  XNOR2_X2 U11187 ( .A(n12949), .B(n12644), .ZN(n12785) );
  INV_X1 U11188 ( .A(n12949), .ZN(n9870) );
  AOI22_X1 U11189 ( .A1(n12783), .A2(n12785), .B1(n12644), .B2(n9870), .ZN(
        n12772) );
  AND2_X1 U11190 ( .A1(n13649), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8825) );
  INV_X1 U11191 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8843) );
  XNOR2_X1 U11192 ( .A(n8843), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n8827) );
  XNOR2_X1 U11193 ( .A(n8842), .B(n8827), .ZN(n13077) );
  NAND2_X1 U11194 ( .A1(n13077), .A2(n12159), .ZN(n8829) );
  OR2_X1 U11195 ( .A1(n8529), .A2(n15236), .ZN(n8828) );
  NAND2_X1 U11196 ( .A1(n8830), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8839) );
  INV_X1 U11197 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13015) );
  OR2_X1 U11198 ( .A1(n8831), .A2(n13015), .ZN(n8838) );
  INV_X1 U11199 ( .A(n8834), .ZN(n8833) );
  INV_X1 U11200 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n8832) );
  NAND2_X1 U11201 ( .A1(n8833), .A2(n8832), .ZN(n12466) );
  NAND2_X1 U11202 ( .A1(n8834), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8835) );
  OR2_X1 U11203 ( .A1(n8510), .A2(n12777), .ZN(n8837) );
  INV_X1 U11204 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n12778) );
  OR2_X1 U11205 ( .A1(n12148), .A2(n12778), .ZN(n8836) );
  NAND4_X1 U11206 ( .A1(n8839), .A2(n8838), .A3(n8837), .A4(n8836), .ZN(n12651) );
  NAND2_X1 U11207 ( .A1(n12538), .A2(n8840), .ZN(n12200) );
  NAND2_X2 U11208 ( .A1(n12201), .A2(n12200), .ZN(n12771) );
  NAND2_X1 U11209 ( .A1(n12770), .A2(n7489), .ZN(n8853) );
  AND2_X1 U11210 ( .A1(n12042), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8841) );
  NAND2_X1 U11211 ( .A1(n8843), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8844) );
  XNOR2_X1 U11212 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n12133) );
  XNOR2_X1 U11213 ( .A(n12137), .B(n12133), .ZN(n13073) );
  NAND2_X1 U11214 ( .A1(n13073), .A2(n12159), .ZN(n8847) );
  OR2_X1 U11215 ( .A1(n8529), .A2(n15285), .ZN(n8846) );
  OR2_X1 U11216 ( .A1(n8510), .A2(n12466), .ZN(n12152) );
  NAND2_X1 U11217 ( .A1(n12145), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8851) );
  INV_X1 U11218 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n8848) );
  OR2_X1 U11219 ( .A1(n8865), .A2(n8848), .ZN(n8850) );
  INV_X1 U11220 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n12468) );
  OR2_X1 U11221 ( .A1(n12148), .A2(n12468), .ZN(n8849) );
  NAND4_X1 U11222 ( .A1(n12152), .A2(n8851), .A3(n8850), .A4(n8849), .ZN(
        n12774) );
  NAND2_X1 U11223 ( .A1(n9888), .A2(n12774), .ZN(n12368) );
  INV_X1 U11224 ( .A(n9888), .ZN(n12472) );
  INV_X1 U11225 ( .A(n12774), .ZN(n8852) );
  NAND2_X1 U11226 ( .A1(n12472), .A2(n8852), .ZN(n12369) );
  XNOR2_X1 U11227 ( .A(n8853), .B(n12198), .ZN(n8872) );
  INV_X1 U11228 ( .A(n8904), .ZN(n8857) );
  XNOR2_X1 U11229 ( .A(n8855), .B(n8854), .ZN(n11030) );
  OR2_X1 U11230 ( .A1(n8454), .A2(n11030), .ZN(n8862) );
  MUX2_X1 U11231 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8856), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n8858) );
  NAND2_X1 U11232 ( .A1(n8858), .A2(n8857), .ZN(n12211) );
  MUX2_X1 U11233 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8860), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n8861) );
  AND2_X1 U11234 ( .A1(n6501), .A2(n8861), .ZN(n9879) );
  NAND2_X1 U11235 ( .A1(n9756), .A2(n9879), .ZN(n12196) );
  INV_X1 U11236 ( .A(n13079), .ZN(n12379) );
  NAND2_X1 U11237 ( .A1(n12379), .A2(n14348), .ZN(n10738) );
  NAND2_X1 U11238 ( .A1(n10738), .A2(n8482), .ZN(n8863) );
  NAND2_X1 U11239 ( .A1(n12384), .A2(n9756), .ZN(n12364) );
  AOI21_X1 U11240 ( .B1(n12379), .B2(P3_B_REG_SCAN_IN), .A(n12925), .ZN(n12764) );
  NAND2_X1 U11241 ( .A1(n12145), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8870) );
  INV_X1 U11242 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n8864) );
  OR2_X1 U11243 ( .A1(n8865), .A2(n8864), .ZN(n8869) );
  INV_X1 U11244 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n8866) );
  OR2_X1 U11245 ( .A1(n8867), .A2(n8866), .ZN(n8868) );
  NAND4_X1 U11246 ( .A1(n12152), .A2(n8870), .A3(n8869), .A4(n8868), .ZN(
        n12650) );
  AOI22_X1 U11247 ( .A1(n12764), .A2(n12650), .B1(n15103), .B2(n12651), .ZN(
        n8871) );
  AND2_X1 U11248 ( .A1(n8873), .A2(n6590), .ZN(n15102) );
  NAND2_X1 U11249 ( .A1(n15087), .A2(n12179), .ZN(n15086) );
  OR2_X1 U11250 ( .A1(n9772), .A2(n15088), .ZN(n12220) );
  NAND2_X1 U11251 ( .A1(n15086), .A2(n12220), .ZN(n11192) );
  NAND2_X1 U11252 ( .A1(n11192), .A2(n12175), .ZN(n8875) );
  NAND2_X1 U11253 ( .A1(n8875), .A2(n12229), .ZN(n11037) );
  NAND2_X1 U11254 ( .A1(n11036), .A2(n12234), .ZN(n11124) );
  INV_X1 U11255 ( .A(n11130), .ZN(n12230) );
  NAND2_X1 U11256 ( .A1(n11124), .A2(n12230), .ZN(n11126) );
  NAND2_X1 U11257 ( .A1(n11126), .A2(n12242), .ZN(n11183) );
  NAND2_X1 U11258 ( .A1(n11183), .A2(n12174), .ZN(n8876) );
  NAND2_X1 U11259 ( .A1(n8876), .A2(n12244), .ZN(n11406) );
  INV_X1 U11260 ( .A(n12670), .ZN(n11330) );
  NAND2_X1 U11261 ( .A1(n11330), .A2(n15149), .ZN(n8877) );
  NAND2_X1 U11262 ( .A1(n11405), .A2(n8877), .ZN(n11327) );
  INV_X1 U11263 ( .A(n9786), .ZN(n15155) );
  OR2_X1 U11264 ( .A1(n12669), .A2(n15155), .ZN(n8879) );
  NAND2_X1 U11265 ( .A1(n12669), .A2(n15155), .ZN(n8878) );
  NAND2_X1 U11266 ( .A1(n8879), .A2(n8878), .ZN(n11326) );
  NAND2_X1 U11267 ( .A1(n11327), .A2(n12252), .ZN(n8880) );
  INV_X1 U11268 ( .A(n12668), .ZN(n11329) );
  NAND2_X1 U11269 ( .A1(n8881), .A2(n12270), .ZN(n11714) );
  NAND2_X1 U11270 ( .A1(n12666), .A2(n11836), .ZN(n12265) );
  NAND2_X1 U11271 ( .A1(n11714), .A2(n12272), .ZN(n8882) );
  NAND2_X1 U11272 ( .A1(n8882), .A2(n12273), .ZN(n11765) );
  INV_X1 U11273 ( .A(n12182), .ZN(n11764) );
  NOR2_X1 U11274 ( .A1(n14407), .A2(n12664), .ZN(n12285) );
  INV_X1 U11275 ( .A(n12285), .ZN(n8883) );
  OR2_X1 U11276 ( .A1(n12555), .A2(n12663), .ZN(n12296) );
  OR2_X1 U11277 ( .A1(n12118), .A2(n12926), .ZN(n12291) );
  NAND2_X1 U11278 ( .A1(n12118), .A2(n12926), .ZN(n12303) );
  NAND2_X1 U11279 ( .A1(n11918), .A2(n12290), .ZN(n8885) );
  NAND2_X1 U11280 ( .A1(n8885), .A2(n12303), .ZN(n12929) );
  INV_X1 U11281 ( .A(n12321), .ZN(n8886) );
  INV_X1 U11282 ( .A(n12876), .ZN(n8887) );
  NAND2_X1 U11283 ( .A1(n8887), .A2(n12875), .ZN(n8889) );
  OR2_X1 U11284 ( .A1(n12877), .A2(n12862), .ZN(n8888) );
  NOR2_X1 U11285 ( .A1(n12865), .A2(n12874), .ZN(n12207) );
  NAND2_X1 U11286 ( .A1(n12865), .A2(n12874), .ZN(n12206) );
  NAND2_X1 U11287 ( .A1(n8890), .A2(n12341), .ZN(n12822) );
  NAND2_X1 U11288 ( .A1(n12949), .A2(n12644), .ZN(n12199) );
  INV_X1 U11289 ( .A(n12200), .ZN(n8893) );
  XOR2_X1 U11290 ( .A(n12198), .B(n12132), .Z(n12469) );
  NAND2_X1 U11291 ( .A1(n12384), .A2(n10881), .ZN(n8894) );
  AOI21_X1 U11292 ( .B1(n12163), .B2(n8894), .A(n9756), .ZN(n8897) );
  NAND2_X1 U11293 ( .A1(n12211), .A2(n10881), .ZN(n8895) );
  AND2_X1 U11294 ( .A1(n11030), .A2(n8895), .ZN(n8896) );
  OR2_X1 U11295 ( .A1(n8897), .A2(n8896), .ZN(n9860) );
  NOR2_X1 U11296 ( .A1(n9883), .A2(n15150), .ZN(n8899) );
  NAND2_X1 U11297 ( .A1(n9860), .A2(n8899), .ZN(n8901) );
  NOR2_X1 U11298 ( .A1(n11030), .A2(n10881), .ZN(n8900) );
  NAND2_X1 U11299 ( .A1(n8454), .A2(n8900), .ZN(n10891) );
  NAND2_X1 U11300 ( .A1(n12163), .A2(n10881), .ZN(n15111) );
  XNOR2_X1 U11301 ( .A(n8921), .B(P3_B_REG_SCAN_IN), .ZN(n8911) );
  INV_X1 U11302 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n8915) );
  NAND2_X1 U11303 ( .A1(n8914), .A2(n8915), .ZN(n8918) );
  NAND2_X1 U11304 ( .A1(n6671), .A2(n8916), .ZN(n8917) );
  INV_X1 U11305 ( .A(n10893), .ZN(n13062) );
  INV_X1 U11306 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n8919) );
  NAND2_X1 U11307 ( .A1(n6671), .A2(n8921), .ZN(n8922) );
  NAND2_X2 U11308 ( .A1(n8923), .A2(n8922), .ZN(n9874) );
  INV_X1 U11309 ( .A(n9874), .ZN(n13064) );
  INV_X1 U11310 ( .A(n8914), .ZN(n8935) );
  NOR2_X1 U11311 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .ZN(
        n8927) );
  NOR4_X1 U11312 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n8926) );
  NOR4_X1 U11313 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n8925) );
  NOR4_X1 U11314 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n8924) );
  NAND4_X1 U11315 ( .A1(n8927), .A2(n8926), .A3(n8925), .A4(n8924), .ZN(n8933)
         );
  NOR4_X1 U11316 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n8931) );
  NOR4_X1 U11317 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n8930) );
  NOR4_X1 U11318 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8929) );
  NOR4_X1 U11319 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n8928) );
  NAND4_X1 U11320 ( .A1(n8931), .A2(n8930), .A3(n8929), .A4(n8928), .ZN(n8932)
         );
  NOR2_X1 U11321 ( .A1(n8933), .A2(n8932), .ZN(n8934) );
  NAND3_X1 U11322 ( .A1(n13062), .A2(n13064), .A3(n9875), .ZN(n9861) );
  INV_X1 U11323 ( .A(n8916), .ZN(n8938) );
  INV_X1 U11324 ( .A(n8921), .ZN(n8937) );
  INV_X1 U11325 ( .A(n8940), .ZN(n8941) );
  NAND2_X1 U11326 ( .A1(n8941), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8942) );
  MUX2_X1 U11327 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8942), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n8944) );
  NAND2_X1 U11328 ( .A1(n8944), .A2(n8943), .ZN(n10723) );
  INV_X1 U11329 ( .A(n12380), .ZN(n10722) );
  INV_X1 U11330 ( .A(n9854), .ZN(n8947) );
  INV_X1 U11331 ( .A(n9883), .ZN(n12381) );
  AND2_X1 U11332 ( .A1(n12381), .A2(n12370), .ZN(n10691) );
  NAND2_X1 U11333 ( .A1(n12211), .A2(n9879), .ZN(n12195) );
  OR3_X1 U11334 ( .A1(n8454), .A2(n11030), .A3(n12195), .ZN(n9857) );
  INV_X1 U11335 ( .A(n9857), .ZN(n8945) );
  OR2_X1 U11336 ( .A1(n10691), .A2(n8945), .ZN(n8946) );
  NAND2_X1 U11337 ( .A1(n8947), .A2(n8946), .ZN(n8950) );
  NAND2_X1 U11338 ( .A1(n9862), .A2(n12380), .ZN(n9866) );
  INV_X1 U11339 ( .A(n9860), .ZN(n8948) );
  NOR2_X1 U11340 ( .A1(n9888), .A2(n13059), .ZN(n8951) );
  INV_X1 U11341 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8952) );
  NOR2_X1 U11342 ( .A1(n15175), .A2(n8952), .ZN(n8953) );
  NAND2_X1 U11343 ( .A1(n8955), .A2(n8954), .ZN(P3_U3456) );
  NAND2_X1 U11344 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9070) );
  NOR2_X1 U11345 ( .A1(n9070), .A2(n9069), .ZN(n9068) );
  NAND2_X1 U11346 ( .A1(n9068), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9096) );
  INV_X1 U11347 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9095) );
  INV_X1 U11348 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9108) );
  AND2_X1 U11349 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n8956) );
  AND2_X1 U11350 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), 
        .ZN(n8957) );
  INV_X1 U11351 ( .A(n9206), .ZN(n8958) );
  NAND2_X1 U11352 ( .A1(n8958), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9221) );
  INV_X1 U11353 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9220) );
  INV_X1 U11354 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8997) );
  INV_X1 U11355 ( .A(n9242), .ZN(n9244) );
  INV_X1 U11356 ( .A(n8959), .ZN(n8999) );
  INV_X1 U11357 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8960) );
  NAND2_X1 U11358 ( .A1(n8999), .A2(n8960), .ZN(n8961) );
  NAND2_X1 U11359 ( .A1(n9244), .A2(n8961), .ZN(n13486) );
  NOR2_X1 U11360 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n8965) );
  NOR2_X1 U11361 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), 
        .ZN(n8966) );
  INV_X1 U11362 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8969) );
  INV_X1 U11363 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8968) );
  AND2_X1 U11364 ( .A1(n8976), .A2(n8983), .ZN(n8971) );
  NAND2_X1 U11365 ( .A1(n8972), .A2(n8971), .ZN(n13638) );
  XNOR2_X2 U11366 ( .A(n8973), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8978) );
  NAND2_X1 U11367 ( .A1(n8972), .A2(n8983), .ZN(n8975) );
  XNOR2_X2 U11368 ( .A(n8977), .B(n8976), .ZN(n8980) );
  INV_X1 U11369 ( .A(n8980), .ZN(n8979) );
  NAND2_X2 U11370 ( .A1(n8980), .A2(n12008), .ZN(n9195) );
  INV_X2 U11371 ( .A(n6709), .ZN(n9324) );
  AOI22_X1 U11372 ( .A1(n9246), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n9324), .B2(
        P2_REG0_REG_18__SCAN_IN), .ZN(n8982) );
  NAND2_X1 U11373 ( .A1(n8980), .A2(n8978), .ZN(n9019) );
  INV_X1 U11374 ( .A(n9019), .ZN(n8996) );
  NAND2_X1 U11375 ( .A1(n9667), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8981) );
  OAI211_X1 U11376 ( .C1(n13486), .C2(n9357), .A(n8982), .B(n8981), .ZN(n13252) );
  INV_X1 U11377 ( .A(n13252), .ZN(n13186) );
  XNOR2_X2 U11378 ( .A(n8984), .B(n8983), .ZN(n10107) );
  INV_X1 U11379 ( .A(n9104), .ZN(n8987) );
  INV_X1 U11380 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n8986) );
  INV_X1 U11381 ( .A(n9130), .ZN(n8992) );
  INV_X1 U11382 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8989) );
  AND2_X1 U11383 ( .A1(n8988), .A2(n8990), .ZN(n8991) );
  NAND2_X1 U11384 ( .A1(n8992), .A2(n8991), .ZN(n9237) );
  NAND2_X1 U11385 ( .A1(n7492), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8993) );
  XNOR2_X1 U11386 ( .A(n8993), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13305) );
  AOI22_X1 U11387 ( .A1(n9331), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n9239), 
        .B2(n13305), .ZN(n8994) );
  INV_X2 U11388 ( .A(n8996), .ZN(n9249) );
  INV_X1 U11389 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13503) );
  NAND2_X1 U11390 ( .A1(n9223), .A2(n8997), .ZN(n8998) );
  NAND2_X1 U11391 ( .A1(n8999), .A2(n8998), .ZN(n13502) );
  OR2_X1 U11392 ( .A1(n13502), .A2(n9357), .ZN(n9003) );
  NAND2_X1 U11393 ( .A1(n9324), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n9001) );
  NAND2_X1 U11394 ( .A1(n9246), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n9000) );
  AND2_X1 U11395 ( .A1(n9001), .A2(n9000), .ZN(n9002) );
  OAI211_X1 U11396 ( .C1(n9249), .C2(n13503), .A(n9003), .B(n9002), .ZN(n13253) );
  INV_X1 U11397 ( .A(n13253), .ZN(n13218) );
  NAND2_X1 U11398 ( .A1(n10636), .A2(n9679), .ZN(n9006) );
  NAND2_X1 U11399 ( .A1(n9237), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9004) );
  XNOR2_X1 U11400 ( .A(n9004), .B(P2_IR_REG_17__SCAN_IN), .ZN(n11624) );
  AOI22_X1 U11401 ( .A1(n9331), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n9239), 
        .B2(n11624), .ZN(n9005) );
  INV_X1 U11402 ( .A(n13600), .ZN(n13505) );
  INV_X1 U11403 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10943) );
  OR2_X1 U11404 ( .A1(n9018), .A2(n10943), .ZN(n9010) );
  INV_X1 U11405 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10947) );
  OR2_X1 U11406 ( .A1(n9019), .A2(n10947), .ZN(n9009) );
  INV_X1 U11407 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9007) );
  NAND2_X1 U11408 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n9012) );
  MUX2_X1 U11409 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9012), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n9015) );
  INV_X1 U11410 ( .A(n9029), .ZN(n9014) );
  NAND2_X1 U11411 ( .A1(n9015), .A2(n9014), .ZN(n10314) );
  XNOR2_X2 U11412 ( .A(n13270), .B(n10267), .ZN(n10264) );
  INV_X1 U11413 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9016) );
  INV_X1 U11414 ( .A(n9195), .ZN(n9017) );
  INV_X1 U11415 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10590) );
  INV_X1 U11416 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10591) );
  INV_X1 U11417 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10316) );
  NAND2_X1 U11418 ( .A1(n6720), .A2(SI_0_), .ZN(n9025) );
  XNOR2_X1 U11419 ( .A(n9025), .B(n9024), .ZN(n13655) );
  MUX2_X1 U11420 ( .A(n10316), .B(n13655), .S(n10098), .Z(n10214) );
  INV_X1 U11421 ( .A(n13270), .ZN(n10244) );
  NAND2_X1 U11422 ( .A1(n10244), .A2(n10267), .ZN(n9026) );
  NAND2_X1 U11423 ( .A1(n10263), .A2(n9026), .ZN(n10364) );
  NAND2_X1 U11424 ( .A1(n10017), .A2(n9679), .ZN(n9031) );
  INV_X1 U11425 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n13637) );
  NOR2_X1 U11426 ( .A1(n9029), .A2(n13637), .ZN(n9027) );
  MUX2_X1 U11427 ( .A(n13637), .B(n9027), .S(P2_IR_REG_2__SCAN_IN), .Z(n9030)
         );
  INV_X1 U11428 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n9028) );
  AND2_X1 U11429 ( .A1(n9029), .A2(n9028), .ZN(n9038) );
  NOR2_X1 U11430 ( .A1(n9030), .A2(n9038), .ZN(n10289) );
  INV_X1 U11431 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10979) );
  OR2_X1 U11432 ( .A1(n9018), .A2(n10979), .ZN(n9034) );
  INV_X1 U11433 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10117) );
  OR2_X1 U11434 ( .A1(n9019), .A2(n10117), .ZN(n9033) );
  OR2_X1 U11435 ( .A1(n9195), .A2(n10398), .ZN(n9032) );
  NAND2_X1 U11436 ( .A1(n10364), .A2(n10363), .ZN(n9037) );
  INV_X1 U11437 ( .A(n13268), .ZN(n10509) );
  NAND2_X1 U11438 ( .A1(n10509), .A2(n6653), .ZN(n9036) );
  NAND2_X1 U11439 ( .A1(n10038), .A2(n9679), .ZN(n9043) );
  INV_X1 U11440 ( .A(n9038), .ZN(n9040) );
  NAND2_X1 U11441 ( .A1(n9040), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9039) );
  MUX2_X1 U11442 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9039), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n9041) );
  AND2_X1 U11443 ( .A1(n9041), .A2(n9051), .ZN(n10333) );
  NAND2_X1 U11444 ( .A1(n9246), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9048) );
  OR2_X1 U11445 ( .A1(n9018), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n9047) );
  INV_X1 U11446 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10290) );
  OR2_X1 U11447 ( .A1(n9249), .A2(n10290), .ZN(n9046) );
  INV_X1 U11448 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9044) );
  OR2_X1 U11449 ( .A1(n9195), .A2(n9044), .ZN(n9045) );
  INV_X1 U11450 ( .A(n13267), .ZN(n10243) );
  NAND2_X1 U11451 ( .A1(n14906), .A2(n10243), .ZN(n9049) );
  NAND2_X1 U11452 ( .A1(n10019), .A2(n9679), .ZN(n9056) );
  NAND2_X1 U11453 ( .A1(n9051), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9050) );
  MUX2_X1 U11454 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9050), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n9054) );
  INV_X1 U11455 ( .A(n9051), .ZN(n9053) );
  INV_X1 U11456 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n9052) );
  NAND2_X1 U11457 ( .A1(n9053), .A2(n9052), .ZN(n9064) );
  NAND2_X1 U11458 ( .A1(n9054), .A2(n9064), .ZN(n14796) );
  INV_X1 U11459 ( .A(n14796), .ZN(n10294) );
  AOI22_X1 U11460 ( .A1(n9187), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n9239), .B2(
        n10294), .ZN(n9055) );
  NAND2_X1 U11461 ( .A1(n9017), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n9060) );
  INV_X1 U11462 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10273) );
  OR2_X1 U11463 ( .A1(n9671), .A2(n10273), .ZN(n9059) );
  OAI21_X1 U11464 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n9070), .ZN(n10954) );
  OR2_X1 U11465 ( .A1(n9018), .A2(n10954), .ZN(n9058) );
  INV_X1 U11466 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10953) );
  OR2_X1 U11467 ( .A1(n9249), .A2(n10953), .ZN(n9057) );
  NAND4_X1 U11468 ( .A1(n9060), .A2(n9059), .A3(n9058), .A4(n9057), .ZN(n13266) );
  XNOR2_X1 U11469 ( .A(n10530), .B(n13266), .ZN(n10525) );
  INV_X1 U11470 ( .A(n13266), .ZN(n11165) );
  NAND2_X1 U11471 ( .A1(n11165), .A2(n10530), .ZN(n9061) );
  NAND2_X1 U11472 ( .A1(n9062), .A2(n9061), .ZN(n11164) );
  OR2_X1 U11473 ( .A1(n10063), .A2(n9664), .ZN(n9067) );
  NAND2_X1 U11474 ( .A1(n9064), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9063) );
  MUX2_X1 U11475 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9063), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n9065) );
  AOI22_X1 U11476 ( .A1(n9187), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n9239), .B2(
        n10347), .ZN(n9066) );
  NAND2_X1 U11477 ( .A1(n9067), .A2(n9066), .ZN(n10602) );
  NAND2_X1 U11478 ( .A1(n9324), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n9075) );
  INV_X1 U11479 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10274) );
  OR2_X1 U11480 ( .A1(n6685), .A2(n10274), .ZN(n9074) );
  INV_X1 U11481 ( .A(n9068), .ZN(n9083) );
  NAND2_X1 U11482 ( .A1(n9070), .A2(n9069), .ZN(n9071) );
  NAND2_X1 U11483 ( .A1(n9083), .A2(n9071), .ZN(n12028) );
  OR2_X1 U11484 ( .A1(n9357), .A2(n12028), .ZN(n9073) );
  INV_X1 U11485 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11168) );
  OR2_X1 U11486 ( .A1(n9249), .A2(n11168), .ZN(n9072) );
  NAND4_X1 U11487 ( .A1(n9075), .A2(n9074), .A3(n9073), .A4(n9072), .ZN(n13265) );
  XNOR2_X1 U11488 ( .A(n10602), .B(n13265), .ZN(n11163) );
  NAND2_X1 U11489 ( .A1(n11164), .A2(n11163), .ZN(n9077) );
  INV_X1 U11490 ( .A(n13265), .ZN(n9441) );
  NAND2_X1 U11491 ( .A1(n10602), .A2(n9441), .ZN(n9076) );
  NAND2_X1 U11492 ( .A1(n9090), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9078) );
  XNOR2_X1 U11493 ( .A(n9078), .B(P2_IR_REG_6__SCAN_IN), .ZN(n13278) );
  AOI22_X1 U11494 ( .A1(n9187), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n9239), .B2(
        n13278), .ZN(n9079) );
  NAND2_X1 U11495 ( .A1(n9246), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9088) );
  INV_X1 U11496 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9081) );
  OR2_X1 U11497 ( .A1(n6709), .A2(n9081), .ZN(n9087) );
  INV_X1 U11498 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9082) );
  NAND2_X1 U11499 ( .A1(n9083), .A2(n9082), .ZN(n9084) );
  NAND2_X1 U11500 ( .A1(n9096), .A2(n9084), .ZN(n14888) );
  OR2_X1 U11501 ( .A1(n9357), .A2(n14888), .ZN(n9086) );
  INV_X1 U11502 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10297) );
  OR2_X1 U11503 ( .A1(n9249), .A2(n10297), .ZN(n9085) );
  NAND4_X1 U11504 ( .A1(n9088), .A2(n9087), .A3(n9086), .A4(n9085), .ZN(n13264) );
  INV_X1 U11505 ( .A(n13264), .ZN(n11166) );
  XNOR2_X1 U11506 ( .A(n14934), .B(n11166), .ZN(n9731) );
  NAND2_X1 U11507 ( .A1(n14934), .A2(n11166), .ZN(n9089) );
  OAI21_X1 U11508 ( .B1(n9090), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9091) );
  XNOR2_X1 U11509 ( .A(n9091), .B(P2_IR_REG_7__SCAN_IN), .ZN(n13293) );
  AOI22_X1 U11510 ( .A1(n9187), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n9239), .B2(
        n13293), .ZN(n9092) );
  NAND2_X1 U11511 ( .A1(n9246), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9101) );
  INV_X1 U11512 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9094) );
  OR2_X1 U11513 ( .A1(n6709), .A2(n9094), .ZN(n9100) );
  NAND2_X1 U11514 ( .A1(n9096), .A2(n9095), .ZN(n9097) );
  NAND2_X1 U11515 ( .A1(n9109), .A2(n9097), .ZN(n11220) );
  OR2_X1 U11516 ( .A1(n9357), .A2(n11220), .ZN(n9099) );
  INV_X1 U11517 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n11227) );
  OR2_X1 U11518 ( .A1(n9249), .A2(n11227), .ZN(n9098) );
  NAND4_X1 U11519 ( .A1(n9101), .A2(n9100), .A3(n9099), .A4(n9098), .ZN(n13263) );
  INV_X1 U11520 ( .A(n13263), .ZN(n9102) );
  OR2_X1 U11521 ( .A1(n11216), .A2(n9102), .ZN(n9727) );
  NAND2_X1 U11522 ( .A1(n11216), .A2(n9102), .ZN(n9726) );
  NAND2_X1 U11523 ( .A1(n9104), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9105) );
  MUX2_X1 U11524 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9105), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n9106) );
  AOI22_X1 U11525 ( .A1(n9187), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n9239), .B2(
        n10415), .ZN(n9107) );
  NAND2_X1 U11526 ( .A1(n9324), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n9114) );
  INV_X1 U11527 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10284) );
  OR2_X1 U11528 ( .A1(n6685), .A2(n10284), .ZN(n9113) );
  NAND2_X1 U11529 ( .A1(n9109), .A2(n9108), .ZN(n9110) );
  NAND2_X1 U11530 ( .A1(n9122), .A2(n9110), .ZN(n10998) );
  OR2_X1 U11531 ( .A1(n9357), .A2(n10998), .ZN(n9112) );
  INV_X1 U11532 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10996) );
  OR2_X1 U11533 ( .A1(n9249), .A2(n10996), .ZN(n9111) );
  NAND4_X1 U11534 ( .A1(n9114), .A2(n9113), .A3(n9112), .A4(n9111), .ZN(n13262) );
  INV_X1 U11535 ( .A(n13262), .ZN(n12393) );
  NAND2_X1 U11536 ( .A1(n14946), .A2(n12393), .ZN(n9116) );
  OR2_X1 U11537 ( .A1(n14946), .A2(n12393), .ZN(n9115) );
  OR2_X1 U11538 ( .A1(n10085), .A2(n9664), .ZN(n9119) );
  NAND2_X1 U11539 ( .A1(n9130), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9117) );
  XNOR2_X1 U11540 ( .A(n9117), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10418) );
  AOI22_X1 U11541 ( .A1(n9187), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n9239), .B2(
        n10418), .ZN(n9118) );
  NAND2_X1 U11542 ( .A1(n9324), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n9127) );
  INV_X1 U11543 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10412) );
  OR2_X1 U11544 ( .A1(n6685), .A2(n10412), .ZN(n9126) );
  INV_X1 U11545 ( .A(n9120), .ZN(n9150) );
  NAND2_X1 U11546 ( .A1(n9122), .A2(n9121), .ZN(n9123) );
  NAND2_X1 U11547 ( .A1(n9150), .A2(n9123), .ZN(n12387) );
  OR2_X1 U11548 ( .A1(n9357), .A2(n12387), .ZN(n9125) );
  INV_X1 U11549 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11207) );
  OR2_X1 U11550 ( .A1(n9249), .A2(n11207), .ZN(n9124) );
  NAND4_X1 U11551 ( .A1(n9127), .A2(n9126), .A3(n9125), .A4(n9124), .ZN(n13261) );
  INV_X1 U11552 ( .A(n13261), .ZN(n9541) );
  OR2_X1 U11553 ( .A1(n12391), .A2(n9541), .ZN(n9128) );
  NAND2_X1 U11554 ( .A1(n12391), .A2(n9541), .ZN(n9129) );
  INV_X1 U11555 ( .A(n9231), .ZN(n9131) );
  NAND2_X1 U11556 ( .A1(n9131), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9132) );
  XNOR2_X1 U11557 ( .A(n9132), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10795) );
  AOI22_X1 U11558 ( .A1(n9187), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n9239), 
        .B2(n10795), .ZN(n9133) );
  NAND2_X1 U11559 ( .A1(n9246), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9140) );
  INV_X1 U11560 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9135) );
  OR2_X1 U11561 ( .A1(n6709), .A2(n9135), .ZN(n9139) );
  INV_X1 U11562 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10423) );
  XNOR2_X1 U11563 ( .A(n9150), .B(n10423), .ZN(n11258) );
  OR2_X1 U11564 ( .A1(n9357), .A2(n11258), .ZN(n9138) );
  INV_X1 U11565 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n9136) );
  OR2_X1 U11566 ( .A1(n9249), .A2(n9136), .ZN(n9137) );
  NAND4_X1 U11567 ( .A1(n9140), .A2(n9139), .A3(n9138), .A4(n9137), .ZN(n13260) );
  XNOR2_X1 U11568 ( .A(n11052), .B(n13260), .ZN(n11047) );
  INV_X1 U11569 ( .A(n13260), .ZN(n11078) );
  NAND2_X1 U11570 ( .A1(n11052), .A2(n11078), .ZN(n9141) );
  NAND2_X1 U11571 ( .A1(n9142), .A2(n9141), .ZN(n11267) );
  NAND2_X1 U11572 ( .A1(n10226), .A2(n9679), .ZN(n9147) );
  INV_X1 U11573 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n9143) );
  AND2_X1 U11574 ( .A1(n9231), .A2(n9143), .ZN(n9159) );
  INV_X1 U11575 ( .A(n9159), .ZN(n9144) );
  NAND2_X1 U11576 ( .A1(n9144), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9145) );
  XNOR2_X1 U11577 ( .A(n9145), .B(P2_IR_REG_11__SCAN_IN), .ZN(n14834) );
  AOI22_X1 U11578 ( .A1(n9187), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n9239), 
        .B2(n14834), .ZN(n9146) );
  NAND2_X1 U11579 ( .A1(n9324), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n9156) );
  INV_X1 U11580 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n9148) );
  OR2_X1 U11581 ( .A1(n6685), .A2(n9148), .ZN(n9155) );
  INV_X1 U11582 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9149) );
  OAI21_X1 U11583 ( .B1(n9150), .B2(n10423), .A(n9149), .ZN(n9152) );
  INV_X1 U11584 ( .A(n9151), .ZN(n9169) );
  NAND2_X1 U11585 ( .A1(n9152), .A2(n9169), .ZN(n11275) );
  OR2_X1 U11586 ( .A1(n9357), .A2(n11275), .ZN(n9154) );
  INV_X1 U11587 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11276) );
  OR2_X1 U11588 ( .A1(n9249), .A2(n11276), .ZN(n9153) );
  NAND4_X1 U11589 ( .A1(n9156), .A2(n9155), .A3(n9154), .A4(n9153), .ZN(n13259) );
  INV_X1 U11590 ( .A(n13259), .ZN(n11313) );
  XNOR2_X1 U11591 ( .A(n14955), .B(n11313), .ZN(n9734) );
  AND2_X1 U11592 ( .A1(n14955), .A2(n11313), .ZN(n9157) );
  NAND2_X1 U11593 ( .A1(n10399), .A2(n9679), .ZN(n9166) );
  INV_X1 U11594 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n9158) );
  AND2_X1 U11595 ( .A1(n9159), .A2(n9158), .ZN(n9163) );
  INV_X1 U11596 ( .A(n9163), .ZN(n9160) );
  NAND2_X1 U11597 ( .A1(n9160), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9161) );
  MUX2_X1 U11598 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9161), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n9164) );
  INV_X1 U11599 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n9162) );
  NAND2_X1 U11600 ( .A1(n9163), .A2(n9162), .ZN(n9176) );
  NAND2_X1 U11601 ( .A1(n9164), .A2(n9176), .ZN(n10799) );
  INV_X1 U11602 ( .A(n10799), .ZN(n14850) );
  AOI22_X1 U11603 ( .A1(n9187), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n9239), 
        .B2(n14850), .ZN(n9165) );
  NAND2_X1 U11604 ( .A1(n9324), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n9174) );
  INV_X1 U11605 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9167) );
  OR2_X1 U11606 ( .A1(n6685), .A2(n9167), .ZN(n9173) );
  INV_X1 U11607 ( .A(n9168), .ZN(n9191) );
  INV_X1 U11608 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n14846) );
  NAND2_X1 U11609 ( .A1(n9169), .A2(n14846), .ZN(n9170) );
  NAND2_X1 U11610 ( .A1(n9191), .A2(n9170), .ZN(n11351) );
  OR2_X1 U11611 ( .A1(n9357), .A2(n11351), .ZN(n9172) );
  INV_X1 U11612 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11318) );
  OR2_X1 U11613 ( .A1(n9249), .A2(n11318), .ZN(n9171) );
  NAND4_X1 U11614 ( .A1(n9174), .A2(n9173), .A3(n9172), .A4(n9171), .ZN(n13258) );
  INV_X1 U11615 ( .A(n13258), .ZN(n11077) );
  NAND2_X1 U11616 ( .A1(n10516), .A2(n9679), .ZN(n9179) );
  NAND2_X1 U11617 ( .A1(n9176), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9175) );
  MUX2_X1 U11618 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9175), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n9177) );
  AOI22_X1 U11619 ( .A1(n9187), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n14866), 
        .B2(n9239), .ZN(n9178) );
  NAND2_X1 U11620 ( .A1(n9324), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n9184) );
  INV_X1 U11621 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9180) );
  OR2_X1 U11622 ( .A1(n6685), .A2(n9180), .ZN(n9183) );
  INV_X1 U11623 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n11368) );
  XNOR2_X1 U11624 ( .A(n9191), .B(n11368), .ZN(n11474) );
  OR2_X1 U11625 ( .A1(n9357), .A2(n11474), .ZN(n9182) );
  INV_X1 U11626 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11475) );
  OR2_X1 U11627 ( .A1(n9249), .A2(n11475), .ZN(n9181) );
  NAND4_X1 U11628 ( .A1(n9184), .A2(n9183), .A3(n9182), .A4(n9181), .ZN(n13257) );
  INV_X1 U11629 ( .A(n13257), .ZN(n14421) );
  NAND2_X1 U11630 ( .A1(n14456), .A2(n14421), .ZN(n9724) );
  INV_X1 U11631 ( .A(n9724), .ZN(n9185) );
  OR2_X1 U11632 ( .A1(n14456), .A2(n14421), .ZN(n9725) );
  NAND2_X1 U11633 ( .A1(n10684), .A2(n9679), .ZN(n9189) );
  NAND2_X1 U11634 ( .A1(n9201), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9186) );
  XNOR2_X1 U11635 ( .A(n9186), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11446) );
  AOI22_X1 U11636 ( .A1(n9239), .A2(n11446), .B1(n9331), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n9188) );
  NAND2_X2 U11637 ( .A1(n9189), .A2(n9188), .ZN(n14443) );
  NAND2_X1 U11638 ( .A1(n9246), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n9199) );
  INV_X1 U11639 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9190) );
  OAI21_X1 U11640 ( .B1(n9191), .B2(n11368), .A(n9190), .ZN(n9192) );
  NAND2_X1 U11641 ( .A1(n9206), .A2(n9192), .ZN(n14436) );
  OR2_X1 U11642 ( .A1(n9357), .A2(n14436), .ZN(n9198) );
  INV_X1 U11643 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n9193) );
  OR2_X1 U11644 ( .A1(n9249), .A2(n9193), .ZN(n9197) );
  INV_X1 U11645 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9194) );
  OR2_X1 U11646 ( .A1(n6709), .A2(n9194), .ZN(n9196) );
  NAND4_X1 U11647 ( .A1(n9199), .A2(n9198), .A3(n9197), .A4(n9196), .ZN(n13256) );
  INV_X1 U11648 ( .A(n13256), .ZN(n11709) );
  NAND2_X1 U11649 ( .A1(n14443), .A2(n11709), .ZN(n9200) );
  INV_X1 U11650 ( .A(n14443), .ZN(n14450) );
  NAND2_X1 U11651 ( .A1(n10632), .A2(n9679), .ZN(n9204) );
  OAI21_X1 U11652 ( .B1(n9201), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9202) );
  XNOR2_X1 U11653 ( .A(n9202), .B(P2_IR_REG_15__SCAN_IN), .ZN(n14872) );
  AOI22_X1 U11654 ( .A1(n14872), .A2(n9239), .B1(n9331), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n9203) );
  INV_X1 U11655 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9205) );
  NAND2_X1 U11656 ( .A1(n9206), .A2(n9205), .ZN(n9207) );
  NAND2_X1 U11657 ( .A1(n9221), .A2(n9207), .ZN(n11742) );
  OR2_X1 U11658 ( .A1(n11742), .A2(n9357), .ZN(n9212) );
  NAND2_X1 U11659 ( .A1(n9324), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n9211) );
  INV_X1 U11660 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9208) );
  OR2_X1 U11661 ( .A1(n6685), .A2(n9208), .ZN(n9210) );
  INV_X1 U11662 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n11704) );
  OR2_X1 U11663 ( .A1(n9249), .A2(n11704), .ZN(n9209) );
  NAND4_X1 U11664 ( .A1(n9212), .A2(n9211), .A3(n9210), .A4(n9209), .ZN(n13255) );
  INV_X1 U11665 ( .A(n13255), .ZN(n14423) );
  NAND2_X1 U11666 ( .A1(n13611), .A2(n14423), .ZN(n9214) );
  OR2_X1 U11667 ( .A1(n13611), .A2(n14423), .ZN(n9213) );
  NAND2_X1 U11668 ( .A1(n9214), .A2(n9213), .ZN(n9736) );
  NAND2_X1 U11669 ( .A1(n11707), .A2(n11708), .ZN(n11706) );
  NAND2_X1 U11670 ( .A1(n10596), .A2(n9679), .ZN(n9219) );
  NAND2_X1 U11671 ( .A1(n9231), .A2(n8988), .ZN(n9215) );
  NAND2_X1 U11672 ( .A1(n9215), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9216) );
  MUX2_X1 U11673 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9216), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n9217) );
  AND2_X1 U11674 ( .A1(n9217), .A2(n9237), .ZN(n11528) );
  AOI22_X1 U11675 ( .A1(n9331), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n9239), 
        .B2(n11528), .ZN(n9218) );
  NAND2_X1 U11676 ( .A1(n9221), .A2(n9220), .ZN(n9222) );
  AND2_X1 U11677 ( .A1(n9223), .A2(n9222), .ZN(n13176) );
  NAND2_X1 U11678 ( .A1(n13176), .A2(n9264), .ZN(n9227) );
  NAND2_X1 U11679 ( .A1(n9324), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n9226) );
  NAND2_X1 U11680 ( .A1(n9246), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n9225) );
  INV_X1 U11681 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13520) );
  OR2_X1 U11682 ( .A1(n9249), .A2(n13520), .ZN(n9224) );
  NAND4_X1 U11683 ( .A1(n9227), .A2(n9226), .A3(n9225), .A4(n9224), .ZN(n13254) );
  NAND2_X1 U11684 ( .A1(n6948), .A2(n13254), .ZN(n9228) );
  INV_X1 U11685 ( .A(n13254), .ZN(n13185) );
  AOI21_X1 U11686 ( .B1(n6945), .B2(n13252), .A(n13480), .ZN(n9229) );
  NAND2_X1 U11687 ( .A1(n12009), .A2(n9679), .ZN(n9241) );
  AND2_X1 U11688 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), 
        .ZN(n9236) );
  INV_X1 U11689 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n9233) );
  INV_X1 U11690 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n9232) );
  NAND3_X1 U11691 ( .A1(n9233), .A2(n9232), .A3(P2_IR_REG_19__SCAN_IN), .ZN(
        n9235) );
  XNOR2_X1 U11692 ( .A(P2_IR_REG_19__SCAN_IN), .B(P2_IR_REG_31__SCAN_IN), .ZN(
        n9234) );
  AOI22_X1 U11693 ( .A1(n9237), .A2(n9236), .B1(n9235), .B2(n9234), .ZN(n9238)
         );
  AOI22_X1 U11694 ( .A1(n9331), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n10216), 
        .B2(n9239), .ZN(n9240) );
  INV_X1 U11695 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n13474) );
  INV_X1 U11696 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9243) );
  NAND2_X1 U11697 ( .A1(n9244), .A2(n9243), .ZN(n9245) );
  NAND2_X1 U11698 ( .A1(n9262), .A2(n9245), .ZN(n13473) );
  OR2_X1 U11699 ( .A1(n13473), .A2(n9357), .ZN(n9248) );
  AOI22_X1 U11700 ( .A1(n9246), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n9324), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n9247) );
  OAI211_X1 U11701 ( .C1(n9249), .C2(n13474), .A(n9248), .B(n9247), .ZN(n13251) );
  XNOR2_X1 U11702 ( .A(n13591), .B(n13251), .ZN(n13466) );
  INV_X1 U11703 ( .A(n13466), .ZN(n9250) );
  NAND2_X1 U11704 ( .A1(n9331), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9251) );
  NAND2_X2 U11705 ( .A1(n9252), .A2(n9251), .ZN(n13586) );
  XNOR2_X1 U11706 ( .A(n9262), .B(P2_REG3_REG_20__SCAN_IN), .ZN(n13459) );
  NAND2_X1 U11707 ( .A1(n13459), .A2(n9264), .ZN(n9258) );
  INV_X1 U11708 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9255) );
  NAND2_X1 U11709 ( .A1(n9324), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n9254) );
  NAND2_X1 U11710 ( .A1(n9667), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n9253) );
  OAI211_X1 U11711 ( .C1(n6685), .C2(n9255), .A(n9254), .B(n9253), .ZN(n9256)
         );
  INV_X1 U11712 ( .A(n9256), .ZN(n9257) );
  NAND2_X1 U11713 ( .A1(n9258), .A2(n9257), .ZN(n13250) );
  XNOR2_X1 U11714 ( .A(n13586), .B(n13250), .ZN(n13455) );
  INV_X1 U11715 ( .A(n13250), .ZN(n9259) );
  NAND2_X1 U11716 ( .A1(n9331), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9260) );
  INV_X1 U11717 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13206) );
  INV_X1 U11718 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13154) );
  OAI21_X1 U11719 ( .B1(n9262), .B2(n13206), .A(n13154), .ZN(n9263) );
  AND2_X1 U11720 ( .A1(n9263), .A2(n9278), .ZN(n13447) );
  NAND2_X1 U11721 ( .A1(n13447), .A2(n9264), .ZN(n9270) );
  INV_X1 U11722 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9267) );
  NAND2_X1 U11723 ( .A1(n9324), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n9266) );
  NAND2_X1 U11724 ( .A1(n9667), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n9265) );
  OAI211_X1 U11725 ( .C1(n6685), .C2(n9267), .A(n9266), .B(n9265), .ZN(n9268)
         );
  INV_X1 U11726 ( .A(n9268), .ZN(n9269) );
  NAND2_X1 U11727 ( .A1(n9270), .A2(n9269), .ZN(n13249) );
  XNOR2_X1 U11728 ( .A(n13581), .B(n13249), .ZN(n13441) );
  INV_X1 U11729 ( .A(n13441), .ZN(n9464) );
  NAND2_X1 U11730 ( .A1(n9272), .A2(n9271), .ZN(n9273) );
  NAND2_X1 U11731 ( .A1(n9331), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n9275) );
  INV_X1 U11732 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9277) );
  INV_X1 U11733 ( .A(n9301), .ZN(n9299) );
  NAND2_X1 U11734 ( .A1(n9278), .A2(n9277), .ZN(n9279) );
  AND2_X1 U11735 ( .A1(n9299), .A2(n9279), .ZN(n13431) );
  NAND2_X1 U11736 ( .A1(n13431), .A2(n9264), .ZN(n9285) );
  INV_X1 U11737 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9282) );
  NAND2_X1 U11738 ( .A1(n9324), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n9281) );
  NAND2_X1 U11739 ( .A1(n9667), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n9280) );
  OAI211_X1 U11740 ( .C1(n6685), .C2(n9282), .A(n9281), .B(n9280), .ZN(n9283)
         );
  INV_X1 U11741 ( .A(n9283), .ZN(n9284) );
  NAND2_X1 U11742 ( .A1(n9285), .A2(n9284), .ZN(n13248) );
  INV_X1 U11743 ( .A(n13248), .ZN(n12517) );
  NOR2_X1 U11744 ( .A1(n13575), .A2(n12517), .ZN(n13406) );
  NAND2_X1 U11745 ( .A1(n11827), .A2(n9679), .ZN(n9287) );
  NAND2_X1 U11746 ( .A1(n9331), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n9286) );
  XNOR2_X1 U11747 ( .A(n9299), .B(P2_REG3_REG_23__SCAN_IN), .ZN(n13418) );
  NAND2_X1 U11748 ( .A1(n13418), .A2(n9264), .ZN(n9293) );
  INV_X1 U11749 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9290) );
  NAND2_X1 U11750 ( .A1(n9324), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n9289) );
  NAND2_X1 U11751 ( .A1(n9667), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n9288) );
  OAI211_X1 U11752 ( .C1(n6685), .C2(n9290), .A(n9289), .B(n9288), .ZN(n9291)
         );
  INV_X1 U11753 ( .A(n9291), .ZN(n9292) );
  NAND2_X1 U11754 ( .A1(n9293), .A2(n9292), .ZN(n13247) );
  INV_X1 U11755 ( .A(n13247), .ZN(n13195) );
  NAND2_X1 U11756 ( .A1(n13569), .A2(n13195), .ZN(n9295) );
  OR2_X1 U11757 ( .A1(n13569), .A2(n13195), .ZN(n9294) );
  NAND2_X1 U11758 ( .A1(n9295), .A2(n9294), .ZN(n13413) );
  INV_X1 U11759 ( .A(n9295), .ZN(n9296) );
  NAND2_X1 U11760 ( .A1(n9331), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n9297) );
  INV_X1 U11761 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13116) );
  INV_X1 U11762 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13197) );
  OAI21_X1 U11763 ( .B1(n9299), .B2(n13116), .A(n13197), .ZN(n9302) );
  AND2_X1 U11764 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(P2_REG3_REG_23__SCAN_IN), 
        .ZN(n9300) );
  NAND2_X1 U11765 ( .A1(n9301), .A2(n9300), .ZN(n9311) );
  NAND2_X1 U11766 ( .A1(n9302), .A2(n9311), .ZN(n13399) );
  OR2_X1 U11767 ( .A1(n13399), .A2(n9357), .ZN(n9308) );
  INV_X1 U11768 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9305) );
  NAND2_X1 U11769 ( .A1(n9324), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9304) );
  NAND2_X1 U11770 ( .A1(n9667), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n9303) );
  OAI211_X1 U11771 ( .C1(n6685), .C2(n9305), .A(n9304), .B(n9303), .ZN(n9306)
         );
  INV_X1 U11772 ( .A(n9306), .ZN(n9307) );
  NAND2_X1 U11773 ( .A1(n9308), .A2(n9307), .ZN(n13246) );
  XNOR2_X1 U11774 ( .A(n13401), .B(n13246), .ZN(n13396) );
  INV_X1 U11775 ( .A(n13396), .ZN(n13391) );
  NAND2_X1 U11776 ( .A1(n11984), .A2(n9679), .ZN(n9310) );
  NAND2_X1 U11777 ( .A1(n9331), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9309) );
  INV_X1 U11778 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13168) );
  NAND2_X1 U11779 ( .A1(n9311), .A2(n13168), .ZN(n9312) );
  AND2_X1 U11780 ( .A1(n9322), .A2(n9312), .ZN(n13385) );
  NAND2_X1 U11781 ( .A1(n13385), .A2(n9264), .ZN(n9318) );
  INV_X1 U11782 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9315) );
  NAND2_X1 U11783 ( .A1(n9324), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n9314) );
  NAND2_X1 U11784 ( .A1(n9667), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n9313) );
  OAI211_X1 U11785 ( .C1(n6685), .C2(n9315), .A(n9314), .B(n9313), .ZN(n9316)
         );
  INV_X1 U11786 ( .A(n9316), .ZN(n9317) );
  NAND2_X1 U11787 ( .A1(n9318), .A2(n9317), .ZN(n13245) );
  INV_X1 U11788 ( .A(n13245), .ZN(n13196) );
  XNOR2_X1 U11789 ( .A(n13558), .B(n13196), .ZN(n13380) );
  INV_X1 U11790 ( .A(n13380), .ZN(n13375) );
  NAND2_X1 U11791 ( .A1(n13651), .A2(n9679), .ZN(n9321) );
  NAND2_X1 U11792 ( .A1(n9331), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9320) );
  INV_X1 U11793 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n13234) );
  NOR2_X1 U11794 ( .A1(n9322), .A2(n13234), .ZN(n9334) );
  INV_X1 U11795 ( .A(n9334), .ZN(n9335) );
  NAND2_X1 U11796 ( .A1(n9322), .A2(n13234), .ZN(n9323) );
  NAND2_X1 U11797 ( .A1(n9335), .A2(n9323), .ZN(n13368) );
  OR2_X1 U11798 ( .A1(n13368), .A2(n9357), .ZN(n9330) );
  INV_X1 U11799 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9327) );
  NAND2_X1 U11800 ( .A1(n9324), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n9326) );
  NAND2_X1 U11801 ( .A1(n9667), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n9325) );
  OAI211_X1 U11802 ( .C1(n6685), .C2(n9327), .A(n9326), .B(n9325), .ZN(n9328)
         );
  INV_X1 U11803 ( .A(n9328), .ZN(n9329) );
  NAND2_X1 U11804 ( .A1(n9330), .A2(n9329), .ZN(n13244) );
  INV_X1 U11805 ( .A(n13244), .ZN(n13167) );
  OR2_X1 U11806 ( .A1(n13553), .A2(n13167), .ZN(n9723) );
  NAND2_X1 U11807 ( .A1(n13553), .A2(n13167), .ZN(n9722) );
  NAND2_X1 U11808 ( .A1(n13648), .A2(n9679), .ZN(n9333) );
  NAND2_X1 U11809 ( .A1(n9331), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9332) );
  AND2_X1 U11810 ( .A1(n9334), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n9345) );
  INV_X1 U11811 ( .A(n9345), .ZN(n9346) );
  INV_X1 U11812 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13109) );
  NAND2_X1 U11813 ( .A1(n9335), .A2(n13109), .ZN(n9336) );
  NAND2_X1 U11814 ( .A1(n13350), .A2(n9264), .ZN(n9342) );
  INV_X1 U11815 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9339) );
  NAND2_X1 U11816 ( .A1(n9667), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n9338) );
  NAND2_X1 U11817 ( .A1(n9324), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9337) );
  OAI211_X1 U11818 ( .C1(n6685), .C2(n9339), .A(n9338), .B(n9337), .ZN(n9340)
         );
  INV_X1 U11819 ( .A(n9340), .ZN(n9341) );
  NAND2_X1 U11820 ( .A1(n9342), .A2(n9341), .ZN(n13243) );
  XNOR2_X1 U11821 ( .A(n13547), .B(n13243), .ZN(n13354) );
  NAND2_X1 U11822 ( .A1(n12041), .A2(n9679), .ZN(n9344) );
  NAND2_X1 U11823 ( .A1(n9331), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9343) );
  NAND2_X1 U11824 ( .A1(n9345), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n9424) );
  INV_X1 U11825 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n13140) );
  NAND2_X1 U11826 ( .A1(n9346), .A2(n13140), .ZN(n9347) );
  NAND2_X1 U11827 ( .A1(n9424), .A2(n9347), .ZN(n13338) );
  OR2_X1 U11828 ( .A1(n13338), .A2(n9357), .ZN(n9353) );
  INV_X1 U11829 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9350) );
  NAND2_X1 U11830 ( .A1(n9324), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n9349) );
  NAND2_X1 U11831 ( .A1(n9667), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n9348) );
  OAI211_X1 U11832 ( .C1(n6685), .C2(n9350), .A(n9349), .B(n9348), .ZN(n9351)
         );
  INV_X1 U11833 ( .A(n9351), .ZN(n9352) );
  NAND2_X1 U11834 ( .A1(n13543), .A2(n13133), .ZN(n9354) );
  INV_X1 U11835 ( .A(n13243), .ZN(n9355) );
  NAND2_X1 U11836 ( .A1(n13547), .A2(n9355), .ZN(n13333) );
  NAND3_X1 U11837 ( .A1(n13353), .A2(n13332), .A3(n13333), .ZN(n13331) );
  OR2_X1 U11838 ( .A1(n9424), .A2(n9357), .ZN(n9363) );
  INV_X1 U11839 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9360) );
  NAND2_X1 U11840 ( .A1(n9324), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9359) );
  NAND2_X1 U11841 ( .A1(n9667), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9358) );
  OAI211_X1 U11842 ( .C1(n6685), .C2(n9360), .A(n9359), .B(n9358), .ZN(n9361)
         );
  INV_X1 U11843 ( .A(n9361), .ZN(n9362) );
  NAND2_X1 U11844 ( .A1(n9363), .A2(n9362), .ZN(n13241) );
  NAND2_X1 U11845 ( .A1(n12043), .A2(n9679), .ZN(n9365) );
  NAND2_X1 U11846 ( .A1(n9331), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n9364) );
  NAND2_X1 U11847 ( .A1(n9370), .A2(n9366), .ZN(n9367) );
  MUX2_X1 U11848 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9368), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n9371) );
  NAND2_X1 U11849 ( .A1(n9369), .A2(n9370), .ZN(n9405) );
  NAND2_X1 U11850 ( .A1(n10216), .A2(n11773), .ZN(n9378) );
  XNOR2_X2 U11851 ( .A(n9372), .B(P2_IR_REG_21__SCAN_IN), .ZN(n9469) );
  INV_X1 U11852 ( .A(n6473), .ZN(n9728) );
  NAND2_X1 U11853 ( .A1(n9469), .A2(n9728), .ZN(n9377) );
  INV_X1 U11854 ( .A(n13133), .ZN(n13242) );
  NAND2_X1 U11855 ( .A1(n9469), .A2(n11773), .ZN(n10219) );
  INV_X1 U11856 ( .A(n14420), .ZN(n13231) );
  INV_X1 U11857 ( .A(n10107), .ZN(n9379) );
  INV_X1 U11858 ( .A(P2_B_REG_SCAN_IN), .ZN(n9398) );
  NOR2_X1 U11859 ( .A1(n13650), .A2(n9398), .ZN(n9380) );
  NOR2_X1 U11860 ( .A1(n14422), .A2(n9380), .ZN(n13321) );
  INV_X1 U11861 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9383) );
  NAND2_X1 U11862 ( .A1(n9667), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9382) );
  NAND2_X1 U11863 ( .A1(n9324), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9381) );
  OAI211_X1 U11864 ( .C1(n6685), .C2(n9383), .A(n9382), .B(n9381), .ZN(n13240)
         );
  NAND2_X1 U11865 ( .A1(n13321), .A2(n13240), .ZN(n9384) );
  NAND2_X1 U11866 ( .A1(n9392), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9389) );
  MUX2_X1 U11867 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9389), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n9390) );
  NAND2_X1 U11868 ( .A1(n9396), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9391) );
  MUX2_X1 U11869 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9391), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n9393) );
  NAND2_X1 U11870 ( .A1(n9393), .A2(n9392), .ZN(n11986) );
  NAND2_X1 U11871 ( .A1(n9394), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9395) );
  MUX2_X1 U11872 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9395), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n9397) );
  NAND2_X1 U11873 ( .A1(n9397), .A2(n9396), .ZN(n11914) );
  XOR2_X1 U11874 ( .A(n11914), .B(n9398), .Z(n9399) );
  NAND2_X1 U11875 ( .A1(n11986), .A2(n9399), .ZN(n9400) );
  INV_X1 U11876 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14923) );
  NAND2_X1 U11877 ( .A1(n14920), .A2(n14923), .ZN(n9402) );
  NAND2_X1 U11878 ( .A1(n13654), .A2(n11914), .ZN(n9401) );
  NAND2_X1 U11879 ( .A1(n9432), .A2(n6473), .ZN(n10208) );
  NOR2_X1 U11880 ( .A1(n10204), .A2(n10354), .ZN(n9408) );
  NOR2_X1 U11881 ( .A1(n11986), .A2(n11914), .ZN(n9403) );
  NAND2_X1 U11882 ( .A1(n9404), .A2(n9403), .ZN(n9891) );
  NAND2_X1 U11883 ( .A1(n9405), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9407) );
  XNOR2_X1 U11884 ( .A(n9407), .B(n9406), .ZN(n9890) );
  AND2_X1 U11885 ( .A1(n9891), .A2(n9890), .ZN(n10200) );
  AND2_X1 U11886 ( .A1(n9408), .A2(n14927), .ZN(n10258) );
  NOR4_X1 U11887 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n9412) );
  NOR4_X1 U11888 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n9411) );
  NOR4_X1 U11889 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9410) );
  NOR4_X1 U11890 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n9409) );
  NAND4_X1 U11891 ( .A1(n9412), .A2(n9411), .A3(n9410), .A4(n9409), .ZN(n9418)
         );
  NOR2_X1 U11892 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n9416) );
  NOR4_X1 U11893 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n9415) );
  NOR4_X1 U11894 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n9414) );
  NOR4_X1 U11895 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n9413) );
  NAND4_X1 U11896 ( .A1(n9416), .A2(n9415), .A3(n9414), .A4(n9413), .ZN(n9417)
         );
  OAI21_X1 U11897 ( .B1(n9418), .B2(n9417), .A(n14920), .ZN(n10257) );
  INV_X1 U11898 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14925) );
  NAND2_X1 U11899 ( .A1(n14920), .A2(n14925), .ZN(n9420) );
  NAND2_X1 U11900 ( .A1(n13654), .A2(n11986), .ZN(n9419) );
  NAND2_X1 U11901 ( .A1(n9420), .A2(n9419), .ZN(n14926) );
  INV_X1 U11902 ( .A(n14926), .ZN(n9421) );
  NAND2_X1 U11903 ( .A1(n10258), .A2(n10206), .ZN(n9423) );
  INV_X1 U11904 ( .A(n9469), .ZN(n11548) );
  NAND2_X1 U11905 ( .A1(n14950), .A2(n11548), .ZN(n10255) );
  INV_X1 U11906 ( .A(n10255), .ZN(n9422) );
  INV_X1 U11907 ( .A(n13537), .ZN(n9427) );
  NAND2_X1 U11908 ( .A1(n10373), .A2(n9728), .ZN(n10218) );
  INV_X1 U11909 ( .A(n10218), .ZN(n14907) );
  INV_X1 U11910 ( .A(n9424), .ZN(n9425) );
  INV_X1 U11911 ( .A(n13518), .ZN(n14905) );
  AOI22_X1 U11912 ( .A1(n9425), .A2(n14905), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n14903), .ZN(n9426) );
  OAI21_X1 U11913 ( .B1(n9427), .B2(n13472), .A(n9426), .ZN(n9428) );
  INV_X1 U11914 ( .A(n9428), .ZN(n9429) );
  INV_X1 U11915 ( .A(n13553), .ZN(n13371) );
  INV_X1 U11916 ( .A(n10602), .ZN(n14930) );
  INV_X1 U11917 ( .A(n14946), .ZN(n10999) );
  INV_X1 U11918 ( .A(n12391), .ZN(n11249) );
  NAND2_X1 U11919 ( .A1(n13563), .A2(n13415), .ZN(n13397) );
  NAND2_X1 U11920 ( .A1(n10373), .A2(n6473), .ZN(n10403) );
  NOR2_X2 U11921 ( .A1(n13537), .A2(n13340), .ZN(n13326) );
  AOI211_X1 U11922 ( .C1(n13537), .C2(n13340), .A(n13105), .B(n13326), .ZN(
        n13536) );
  INV_X1 U11923 ( .A(n10264), .ZN(n9435) );
  INV_X1 U11924 ( .A(n10214), .ZN(n10408) );
  NAND2_X1 U11925 ( .A1(n9477), .A2(n10408), .ZN(n10259) );
  NAND2_X1 U11926 ( .A1(n9435), .A2(n10259), .ZN(n10260) );
  NAND2_X1 U11927 ( .A1(n10244), .A2(n10944), .ZN(n9436) );
  NAND2_X1 U11928 ( .A1(n10260), .A2(n9436), .ZN(n10359) );
  INV_X1 U11929 ( .A(n10363), .ZN(n10358) );
  NAND2_X1 U11930 ( .A1(n10359), .A2(n10358), .ZN(n10357) );
  NAND2_X1 U11931 ( .A1(n10980), .A2(n10509), .ZN(n9437) );
  NAND2_X1 U11932 ( .A1(n10357), .A2(n9437), .ZN(n10504) );
  INV_X1 U11933 ( .A(n10508), .ZN(n10503) );
  OR2_X1 U11934 ( .A1(n14906), .A2(n13267), .ZN(n9438) );
  NAND2_X1 U11935 ( .A1(n10502), .A2(n9438), .ZN(n10523) );
  INV_X1 U11936 ( .A(n10525), .ZN(n10522) );
  NAND2_X1 U11937 ( .A1(n10523), .A2(n10522), .ZN(n10521) );
  OR2_X1 U11938 ( .A1(n13266), .A2(n10530), .ZN(n9439) );
  NAND2_X1 U11939 ( .A1(n10521), .A2(n9439), .ZN(n11159) );
  NAND2_X1 U11940 ( .A1(n10602), .A2(n13265), .ZN(n9440) );
  NAND2_X1 U11941 ( .A1(n14930), .A2(n9441), .ZN(n9442) );
  NAND2_X1 U11942 ( .A1(n14934), .A2(n13264), .ZN(n9443) );
  OR2_X1 U11943 ( .A1(n11216), .A2(n13263), .ZN(n9444) );
  NAND2_X1 U11944 ( .A1(n11215), .A2(n9444), .ZN(n9446) );
  NAND2_X1 U11945 ( .A1(n11216), .A2(n13263), .ZN(n9445) );
  INV_X1 U11946 ( .A(n10991), .ZN(n9447) );
  NAND2_X1 U11947 ( .A1(n10988), .A2(n9447), .ZN(n9449) );
  NAND2_X1 U11948 ( .A1(n14946), .A2(n13262), .ZN(n9448) );
  NAND2_X1 U11949 ( .A1(n9449), .A2(n9448), .ZN(n11201) );
  XNOR2_X1 U11950 ( .A(n12391), .B(n13261), .ZN(n11202) );
  INV_X1 U11951 ( .A(n11202), .ZN(n11203) );
  NAND2_X1 U11952 ( .A1(n11201), .A2(n11203), .ZN(n9451) );
  NAND2_X1 U11953 ( .A1(n12391), .A2(n13261), .ZN(n9450) );
  OR2_X1 U11954 ( .A1(n14955), .A2(n13259), .ZN(n9452) );
  NOR2_X1 U11955 ( .A1(n11353), .A2(n13258), .ZN(n9454) );
  AND2_X1 U11956 ( .A1(n14456), .A2(n13257), .ZN(n9455) );
  OR2_X1 U11957 ( .A1(n14456), .A2(n13257), .ZN(n9456) );
  XNOR2_X1 U11958 ( .A(n14443), .B(n13256), .ZN(n14438) );
  NAND2_X1 U11959 ( .A1(n14443), .A2(n13256), .ZN(n9457) );
  OR2_X1 U11960 ( .A1(n13611), .A2(n13255), .ZN(n9458) );
  XNOR2_X1 U11961 ( .A(n13607), .B(n13254), .ZN(n13515) );
  XNOR2_X1 U11962 ( .A(n13600), .B(n13253), .ZN(n9738) );
  NAND2_X1 U11963 ( .A1(n13600), .A2(n13253), .ZN(n9459) );
  XNOR2_X1 U11964 ( .A(n13595), .B(n13186), .ZN(n13479) );
  OR2_X1 U11965 ( .A1(n13595), .A2(n13252), .ZN(n9460) );
  NOR2_X1 U11966 ( .A1(n13591), .A2(n13251), .ZN(n9461) );
  INV_X1 U11967 ( .A(n13251), .ZN(n13219) );
  AND2_X1 U11968 ( .A1(n13586), .A2(n13250), .ZN(n9462) );
  OR2_X1 U11969 ( .A1(n13586), .A2(n13250), .ZN(n9463) );
  INV_X1 U11970 ( .A(n13249), .ZN(n9465) );
  NOR2_X1 U11971 ( .A1(n13436), .A2(n9466), .ZN(n13414) );
  NAND2_X1 U11972 ( .A1(n13414), .A2(n13413), .ZN(n13412) );
  NOR2_X1 U11973 ( .A1(n13553), .A2(n13244), .ZN(n9468) );
  XNOR2_X1 U11974 ( .A(n9478), .B(n11773), .ZN(n9470) );
  AND2_X1 U11975 ( .A1(n9472), .A2(n9469), .ZN(n10587) );
  OR2_X1 U11976 ( .A1(n9471), .A2(n10587), .ZN(n9473) );
  NAND2_X1 U11977 ( .A1(n9476), .A2(n9514), .ZN(n9481) );
  INV_X1 U11978 ( .A(n9478), .ZN(n10211) );
  INV_X1 U11979 ( .A(n14950), .ZN(n10374) );
  NAND3_X1 U11980 ( .A1(n10405), .A2(n10211), .A3(n10374), .ZN(n9479) );
  NAND3_X1 U11981 ( .A1(n9481), .A2(n9480), .A3(n9479), .ZN(n9486) );
  NAND2_X1 U11982 ( .A1(n13270), .A2(n9647), .ZN(n9483) );
  NAND2_X1 U11983 ( .A1(n9514), .A2(n10267), .ZN(n9482) );
  NAND2_X1 U11984 ( .A1(n9483), .A2(n9482), .ZN(n9485) );
  AOI22_X1 U11985 ( .A1(n13270), .A2(n9514), .B1(n9647), .B2(n10267), .ZN(
        n9484) );
  AOI21_X1 U11986 ( .B1(n9486), .B2(n9485), .A(n9484), .ZN(n9488) );
  NOR2_X1 U11987 ( .A1(n9486), .A2(n9485), .ZN(n9487) );
  NAND2_X1 U11988 ( .A1(n6653), .A2(n9647), .ZN(n9490) );
  NAND2_X1 U11989 ( .A1(n13268), .A2(n9514), .ZN(n9489) );
  NAND2_X1 U11990 ( .A1(n6653), .A2(n9514), .ZN(n9492) );
  NAND2_X1 U11991 ( .A1(n13268), .A2(n9647), .ZN(n9491) );
  NAND2_X1 U11992 ( .A1(n9492), .A2(n9491), .ZN(n9493) );
  NAND2_X1 U11993 ( .A1(n14906), .A2(n9676), .ZN(n9495) );
  NAND2_X1 U11994 ( .A1(n13267), .A2(n9647), .ZN(n9494) );
  NAND2_X1 U11995 ( .A1(n9495), .A2(n9494), .ZN(n9497) );
  AOI22_X1 U11996 ( .A1(n14906), .A2(n6476), .B1(n9676), .B2(n13267), .ZN(
        n9496) );
  NAND2_X1 U11997 ( .A1(n10530), .A2(n6476), .ZN(n9500) );
  NAND2_X1 U11998 ( .A1(n13266), .A2(n9676), .ZN(n9499) );
  NAND2_X1 U11999 ( .A1(n9500), .A2(n9499), .ZN(n9505) );
  NAND2_X1 U12000 ( .A1(n10530), .A2(n9676), .ZN(n9502) );
  NAND2_X1 U12001 ( .A1(n13266), .A2(n6476), .ZN(n9501) );
  NAND2_X1 U12002 ( .A1(n9502), .A2(n9501), .ZN(n9503) );
  INV_X1 U12003 ( .A(n9505), .ZN(n9506) );
  NAND2_X1 U12004 ( .A1(n10602), .A2(n9676), .ZN(n9508) );
  NAND2_X1 U12005 ( .A1(n13265), .A2(n9705), .ZN(n9507) );
  NAND2_X1 U12006 ( .A1(n9508), .A2(n9507), .ZN(n9511) );
  AOI22_X1 U12007 ( .A1(n10602), .A2(n9705), .B1(n9676), .B2(n13265), .ZN(
        n9509) );
  INV_X1 U12008 ( .A(n9510), .ZN(n9513) );
  NAND2_X1 U12009 ( .A1(n9513), .A2(n7483), .ZN(n9520) );
  NAND2_X1 U12010 ( .A1(n14934), .A2(n9705), .ZN(n9516) );
  NAND2_X1 U12011 ( .A1(n13264), .A2(n9686), .ZN(n9515) );
  NAND2_X1 U12012 ( .A1(n9516), .A2(n9515), .ZN(n9521) );
  NAND2_X1 U12013 ( .A1(n9520), .A2(n9521), .ZN(n9519) );
  NAND2_X1 U12014 ( .A1(n14934), .A2(n9686), .ZN(n9517) );
  OAI21_X1 U12015 ( .B1(n11166), .B2(n9686), .A(n9517), .ZN(n9518) );
  NAND2_X1 U12016 ( .A1(n9519), .A2(n9518), .ZN(n9525) );
  NAND2_X1 U12017 ( .A1(n9523), .A2(n9522), .ZN(n9524) );
  NAND2_X1 U12018 ( .A1(n11216), .A2(n9686), .ZN(n9527) );
  NAND2_X1 U12019 ( .A1(n13263), .A2(n9705), .ZN(n9526) );
  AOI22_X1 U12020 ( .A1(n11216), .A2(n9705), .B1(n9686), .B2(n13263), .ZN(
        n9528) );
  INV_X1 U12021 ( .A(n9528), .ZN(n9529) );
  NAND2_X1 U12022 ( .A1(n14946), .A2(n9705), .ZN(n9531) );
  NAND2_X1 U12023 ( .A1(n13262), .A2(n9686), .ZN(n9530) );
  NAND2_X1 U12024 ( .A1(n9531), .A2(n9530), .ZN(n9533) );
  AOI22_X1 U12025 ( .A1(n14946), .A2(n9686), .B1(n9705), .B2(n13262), .ZN(
        n9532) );
  INV_X1 U12026 ( .A(n9535), .ZN(n9536) );
  NAND2_X1 U12027 ( .A1(n12391), .A2(n9686), .ZN(n9539) );
  NAND2_X1 U12028 ( .A1(n13261), .A2(n9705), .ZN(n9538) );
  NAND2_X1 U12029 ( .A1(n12391), .A2(n9705), .ZN(n9540) );
  OAI21_X1 U12030 ( .B1(n9705), .B2(n9541), .A(n9540), .ZN(n9542) );
  NAND2_X1 U12031 ( .A1(n11052), .A2(n9705), .ZN(n9544) );
  NAND2_X1 U12032 ( .A1(n13260), .A2(n9686), .ZN(n9543) );
  NAND2_X1 U12033 ( .A1(n9544), .A2(n9543), .ZN(n9547) );
  AOI22_X1 U12034 ( .A1(n11052), .A2(n9686), .B1(n9705), .B2(n13260), .ZN(
        n9545) );
  INV_X1 U12035 ( .A(n9546), .ZN(n9549) );
  NAND2_X1 U12036 ( .A1(n14955), .A2(n9686), .ZN(n9551) );
  NAND2_X1 U12037 ( .A1(n13259), .A2(n9705), .ZN(n9550) );
  NAND2_X1 U12038 ( .A1(n9551), .A2(n9550), .ZN(n9554) );
  NAND2_X1 U12039 ( .A1(n14955), .A2(n9705), .ZN(n9552) );
  OAI21_X1 U12040 ( .B1(n9705), .B2(n11313), .A(n9552), .ZN(n9553) );
  INV_X1 U12041 ( .A(n9553), .ZN(n9555) );
  NAND2_X1 U12042 ( .A1(n11353), .A2(n9705), .ZN(n9557) );
  NAND2_X1 U12043 ( .A1(n13258), .A2(n9686), .ZN(n9556) );
  NAND2_X1 U12044 ( .A1(n9557), .A2(n9556), .ZN(n9559) );
  AOI22_X1 U12045 ( .A1(n11353), .A2(n9686), .B1(n9705), .B2(n13258), .ZN(
        n9558) );
  NAND2_X1 U12046 ( .A1(n14456), .A2(n9686), .ZN(n9562) );
  NAND2_X1 U12047 ( .A1(n13257), .A2(n9705), .ZN(n9561) );
  NAND2_X1 U12048 ( .A1(n9562), .A2(n9561), .ZN(n9580) );
  AND2_X1 U12049 ( .A1(n13253), .A2(n9705), .ZN(n9563) );
  AOI21_X1 U12050 ( .B1(n13600), .B2(n9686), .A(n9563), .ZN(n9593) );
  NAND2_X1 U12051 ( .A1(n13600), .A2(n9705), .ZN(n9565) );
  NAND2_X1 U12052 ( .A1(n13253), .A2(n9686), .ZN(n9564) );
  NAND2_X1 U12053 ( .A1(n9565), .A2(n9564), .ZN(n9591) );
  NAND2_X1 U12054 ( .A1(n9593), .A2(n9591), .ZN(n9570) );
  AND2_X1 U12055 ( .A1(n13254), .A2(n9705), .ZN(n9566) );
  AOI21_X1 U12056 ( .B1(n13607), .B2(n9686), .A(n9566), .ZN(n9588) );
  NAND2_X1 U12057 ( .A1(n13607), .A2(n9705), .ZN(n9568) );
  NAND2_X1 U12058 ( .A1(n13254), .A2(n9686), .ZN(n9567) );
  NAND2_X1 U12059 ( .A1(n9568), .A2(n9567), .ZN(n9587) );
  NAND2_X1 U12060 ( .A1(n9588), .A2(n9587), .ZN(n9569) );
  NAND2_X1 U12061 ( .A1(n9570), .A2(n9569), .ZN(n9600) );
  AND2_X1 U12062 ( .A1(n13255), .A2(n9705), .ZN(n9571) );
  AOI21_X1 U12063 ( .B1(n13611), .B2(n9686), .A(n9571), .ZN(n9599) );
  NAND2_X1 U12064 ( .A1(n13611), .A2(n9705), .ZN(n9573) );
  NAND2_X1 U12065 ( .A1(n13255), .A2(n9686), .ZN(n9572) );
  NAND2_X1 U12066 ( .A1(n9573), .A2(n9572), .ZN(n9598) );
  AND2_X1 U12067 ( .A1(n9599), .A2(n9598), .ZN(n9574) );
  NOR2_X1 U12068 ( .A1(n9600), .A2(n9574), .ZN(n9582) );
  AND2_X1 U12069 ( .A1(n13256), .A2(n9705), .ZN(n9575) );
  AOI21_X1 U12070 ( .B1(n14443), .B2(n9686), .A(n9575), .ZN(n9584) );
  NAND2_X1 U12071 ( .A1(n14443), .A2(n9705), .ZN(n9577) );
  NAND2_X1 U12072 ( .A1(n13256), .A2(n9686), .ZN(n9576) );
  NAND2_X1 U12073 ( .A1(n9577), .A2(n9576), .ZN(n9583) );
  NAND2_X1 U12074 ( .A1(n9584), .A2(n9583), .ZN(n9578) );
  OAI211_X1 U12075 ( .C1(n9581), .C2(n9580), .A(n9582), .B(n9578), .ZN(n9608)
         );
  AOI22_X1 U12076 ( .A1(n14456), .A2(n9705), .B1(n9686), .B2(n13257), .ZN(
        n9579) );
  AOI21_X1 U12077 ( .B1(n9581), .B2(n9580), .A(n9579), .ZN(n9607) );
  INV_X1 U12078 ( .A(n9582), .ZN(n9604) );
  INV_X1 U12079 ( .A(n9583), .ZN(n9586) );
  INV_X1 U12080 ( .A(n9584), .ZN(n9585) );
  NAND2_X1 U12081 ( .A1(n9586), .A2(n9585), .ZN(n9603) );
  INV_X1 U12082 ( .A(n9587), .ZN(n9590) );
  INV_X1 U12083 ( .A(n9588), .ZN(n9589) );
  NAND2_X1 U12084 ( .A1(n9590), .A2(n9589), .ZN(n9592) );
  NAND3_X1 U12085 ( .A1(n9592), .A2(n13505), .A3(n13218), .ZN(n9597) );
  INV_X1 U12086 ( .A(n9591), .ZN(n9596) );
  INV_X1 U12087 ( .A(n9592), .ZN(n9595) );
  INV_X1 U12088 ( .A(n9593), .ZN(n9594) );
  AOI22_X1 U12089 ( .A1(n9597), .A2(n9596), .B1(n9595), .B2(n9594), .ZN(n9602)
         );
  OR3_X1 U12090 ( .A1(n9600), .A2(n9599), .A3(n9598), .ZN(n9601) );
  OAI211_X1 U12091 ( .C1(n9604), .C2(n9603), .A(n9602), .B(n9601), .ZN(n9605)
         );
  INV_X1 U12092 ( .A(n9605), .ZN(n9606) );
  AND2_X1 U12093 ( .A1(n13252), .A2(n9686), .ZN(n9609) );
  AOI21_X1 U12094 ( .B1(n13595), .B2(n9705), .A(n9609), .ZN(n9613) );
  NAND2_X1 U12095 ( .A1(n13595), .A2(n9686), .ZN(n9611) );
  NAND2_X1 U12096 ( .A1(n13252), .A2(n9705), .ZN(n9610) );
  NAND2_X1 U12097 ( .A1(n9611), .A2(n9610), .ZN(n9612) );
  OAI21_X1 U12098 ( .B1(n9614), .B2(n9613), .A(n9612), .ZN(n9616) );
  NAND2_X1 U12099 ( .A1(n9614), .A2(n9613), .ZN(n9615) );
  NAND2_X1 U12100 ( .A1(n13591), .A2(n9686), .ZN(n9618) );
  NAND2_X1 U12101 ( .A1(n13251), .A2(n9705), .ZN(n9617) );
  NAND2_X1 U12102 ( .A1(n13591), .A2(n9705), .ZN(n9619) );
  OAI21_X1 U12103 ( .B1(n9705), .B2(n13219), .A(n9619), .ZN(n9620) );
  NAND2_X1 U12104 ( .A1(n13586), .A2(n9705), .ZN(n9622) );
  NAND2_X1 U12105 ( .A1(n13250), .A2(n9686), .ZN(n9621) );
  NAND2_X1 U12106 ( .A1(n9622), .A2(n9621), .ZN(n9624) );
  AOI22_X1 U12107 ( .A1(n13586), .A2(n9686), .B1(n9705), .B2(n13250), .ZN(
        n9623) );
  NAND2_X1 U12108 ( .A1(n13581), .A2(n9686), .ZN(n9627) );
  NAND2_X1 U12109 ( .A1(n13249), .A2(n9705), .ZN(n9626) );
  AOI22_X1 U12110 ( .A1(n13581), .A2(n9705), .B1(n9686), .B2(n13249), .ZN(
        n9628) );
  NAND2_X1 U12111 ( .A1(n13575), .A2(n9705), .ZN(n9630) );
  NAND2_X1 U12112 ( .A1(n13248), .A2(n9686), .ZN(n9629) );
  NAND2_X1 U12113 ( .A1(n9630), .A2(n9629), .ZN(n9635) );
  NAND2_X1 U12114 ( .A1(n9636), .A2(n9635), .ZN(n9634) );
  NAND2_X1 U12115 ( .A1(n13575), .A2(n9686), .ZN(n9632) );
  NAND2_X1 U12116 ( .A1(n13248), .A2(n6476), .ZN(n9631) );
  NAND2_X1 U12117 ( .A1(n9632), .A2(n9631), .ZN(n9633) );
  NAND2_X1 U12118 ( .A1(n13569), .A2(n9686), .ZN(n9638) );
  NAND2_X1 U12119 ( .A1(n13247), .A2(n9705), .ZN(n9637) );
  AOI22_X1 U12120 ( .A1(n13569), .A2(n9705), .B1(n9686), .B2(n13247), .ZN(
        n9639) );
  NAND2_X1 U12121 ( .A1(n13401), .A2(n9705), .ZN(n9641) );
  NAND2_X1 U12122 ( .A1(n13246), .A2(n9514), .ZN(n9640) );
  NAND2_X1 U12123 ( .A1(n9641), .A2(n9640), .ZN(n9643) );
  AOI22_X1 U12124 ( .A1(n13401), .A2(n9686), .B1(n9705), .B2(n13246), .ZN(
        n9642) );
  INV_X1 U12125 ( .A(n9645), .ZN(n9646) );
  NAND2_X1 U12126 ( .A1(n13558), .A2(n9676), .ZN(n9649) );
  NAND2_X1 U12127 ( .A1(n13245), .A2(n9705), .ZN(n9648) );
  NAND2_X1 U12128 ( .A1(n9649), .A2(n9648), .ZN(n9652) );
  NAND2_X1 U12129 ( .A1(n13558), .A2(n9705), .ZN(n9650) );
  OAI21_X1 U12130 ( .B1(n9705), .B2(n13196), .A(n9650), .ZN(n9651) );
  NAND2_X1 U12131 ( .A1(n13553), .A2(n6476), .ZN(n9654) );
  NAND2_X1 U12132 ( .A1(n13244), .A2(n9514), .ZN(n9653) );
  NAND2_X1 U12133 ( .A1(n9654), .A2(n9653), .ZN(n9656) );
  AOI22_X1 U12134 ( .A1(n13553), .A2(n9686), .B1(n9705), .B2(n13244), .ZN(
        n9655) );
  NAND2_X1 U12135 ( .A1(n13547), .A2(n9686), .ZN(n9660) );
  NAND2_X1 U12136 ( .A1(n13243), .A2(n9705), .ZN(n9659) );
  NAND2_X1 U12137 ( .A1(n9660), .A2(n9659), .ZN(n9688) );
  AOI22_X1 U12138 ( .A1(n13547), .A2(n9705), .B1(n9686), .B2(n13243), .ZN(
        n9661) );
  AOI21_X1 U12139 ( .B1(n9689), .B2(n9688), .A(n9661), .ZN(n9662) );
  INV_X1 U12140 ( .A(n9662), .ZN(n9685) );
  INV_X1 U12141 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12138) );
  OAI22_X1 U12142 ( .A1(n9665), .A2(n9664), .B1(n9663), .B2(n12138), .ZN(n9666) );
  AOI22_X1 U12143 ( .A1(n9666), .A2(n9676), .B1(n6476), .B2(n13240), .ZN(n9700) );
  INV_X1 U12144 ( .A(n9666), .ZN(n9721) );
  INV_X1 U12145 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9670) );
  NAND2_X1 U12146 ( .A1(n9667), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9669) );
  NAND2_X1 U12147 ( .A1(n9324), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9668) );
  OAI211_X1 U12148 ( .C1(n6685), .C2(n9670), .A(n9669), .B(n9668), .ZN(n13322)
         );
  AND2_X1 U12149 ( .A1(n13322), .A2(n9686), .ZN(n9706) );
  NAND2_X1 U12150 ( .A1(n9472), .A2(n11773), .ZN(n9716) );
  NAND2_X1 U12151 ( .A1(n9716), .A2(n9672), .ZN(n9673) );
  OAI21_X1 U12152 ( .B1(n9706), .B2(n9673), .A(n13240), .ZN(n9674) );
  OAI21_X1 U12153 ( .B1(n9721), .B2(n9686), .A(n9674), .ZN(n9699) );
  AND2_X1 U12154 ( .A1(n13241), .A2(n9705), .ZN(n9675) );
  AOI21_X1 U12155 ( .B1(n13537), .B2(n9514), .A(n9675), .ZN(n9691) );
  NAND2_X1 U12156 ( .A1(n13537), .A2(n9705), .ZN(n9678) );
  NAND2_X1 U12157 ( .A1(n13241), .A2(n9686), .ZN(n9677) );
  NAND2_X1 U12158 ( .A1(n9678), .A2(n9677), .ZN(n9690) );
  AOI22_X1 U12159 ( .A1(n9700), .A2(n9699), .B1(n9691), .B2(n9690), .ZN(n9683)
         );
  NAND2_X1 U12160 ( .A1(n9331), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n9680) );
  INV_X1 U12161 ( .A(n13322), .ZN(n9682) );
  XNOR2_X1 U12162 ( .A(n9707), .B(n9682), .ZN(n9696) );
  INV_X1 U12163 ( .A(n9697), .ZN(n9684) );
  AOI22_X1 U12164 ( .A1(n13543), .A2(n9705), .B1(n9686), .B2(n13242), .ZN(
        n9693) );
  OAI22_X1 U12165 ( .A1(n13344), .A2(n6476), .B1(n13133), .B2(n9514), .ZN(
        n9692) );
  INV_X1 U12166 ( .A(n9690), .ZN(n9695) );
  INV_X1 U12167 ( .A(n9691), .ZN(n9694) );
  AOI22_X1 U12168 ( .A1(n9695), .A2(n9694), .B1(n9693), .B2(n9692), .ZN(n9698)
         );
  AOI21_X1 U12169 ( .B1(n9698), .B2(n9745), .A(n9697), .ZN(n9703) );
  INV_X1 U12170 ( .A(n9699), .ZN(n9702) );
  INV_X1 U12171 ( .A(n9700), .ZN(n9701) );
  NOR2_X1 U12172 ( .A1(n9703), .A2(n7493), .ZN(n9704) );
  AND2_X1 U12173 ( .A1(n9705), .A2(n13322), .ZN(n9709) );
  NOR2_X1 U12174 ( .A1(n9706), .A2(n6476), .ZN(n9708) );
  MUX2_X1 U12175 ( .A(n9709), .B(n9708), .S(n9707), .Z(n9710) );
  INV_X1 U12176 ( .A(n9710), .ZN(n9711) );
  INV_X1 U12177 ( .A(n9718), .ZN(n9749) );
  OAI21_X1 U12178 ( .B1(n9469), .B2(n6473), .A(n9432), .ZN(n9713) );
  OAI21_X1 U12179 ( .B1(n9478), .B2(n11773), .A(n9713), .ZN(n9714) );
  NAND2_X1 U12180 ( .A1(n9749), .A2(n9714), .ZN(n9720) );
  NAND3_X1 U12181 ( .A1(n10216), .A2(n9469), .A3(n9728), .ZN(n9715) );
  NAND2_X1 U12182 ( .A1(n9716), .A2(n9715), .ZN(n9717) );
  NAND2_X1 U12183 ( .A1(n9720), .A2(n9719), .ZN(n9751) );
  NAND2_X1 U12184 ( .A1(n9723), .A2(n9722), .ZN(n13363) );
  NAND2_X1 U12185 ( .A1(n9725), .A2(n9724), .ZN(n11472) );
  XNOR2_X1 U12186 ( .A(n11353), .B(n11077), .ZN(n11315) );
  NAND2_X1 U12187 ( .A1(n9727), .A2(n9726), .ZN(n11224) );
  OAI21_X1 U12188 ( .B1(n9477), .B2(n10408), .A(n10259), .ZN(n10595) );
  AND4_X1 U12189 ( .A1(n10264), .A2(n9728), .A3(n10363), .A4(n10595), .ZN(
        n9729) );
  NAND4_X1 U12190 ( .A1(n11163), .A2(n9729), .A3(n10508), .A4(n10525), .ZN(
        n9730) );
  NOR3_X1 U12191 ( .A1(n11224), .A2(n9731), .A3(n9730), .ZN(n9732) );
  NAND4_X1 U12192 ( .A1(n11047), .A2(n10991), .A3(n9732), .A4(n11202), .ZN(
        n9733) );
  OR4_X1 U12193 ( .A1(n11472), .A2(n11315), .A3(n9734), .A4(n9733), .ZN(n9735)
         );
  NOR2_X1 U12194 ( .A1(n9736), .A2(n9735), .ZN(n9737) );
  NAND4_X1 U12195 ( .A1(n9738), .A2(n9737), .A3(n13515), .A4(n14438), .ZN(
        n9739) );
  NOR2_X1 U12196 ( .A1(n13479), .A2(n9739), .ZN(n9740) );
  NAND4_X1 U12197 ( .A1(n13441), .A2(n9740), .A3(n13455), .A4(n13466), .ZN(
        n9741) );
  NOR2_X1 U12198 ( .A1(n13413), .A2(n9741), .ZN(n9742) );
  NAND3_X1 U12199 ( .A1(n13396), .A2(n9742), .A3(n13433), .ZN(n9743) );
  NOR3_X1 U12200 ( .A1(n13363), .A2(n13380), .A3(n9743), .ZN(n9744) );
  OR2_X1 U12201 ( .A1(n9890), .A2(P2_U3088), .ZN(n11824) );
  INV_X1 U12202 ( .A(n14927), .ZN(n14924) );
  OAI21_X1 U12203 ( .B1(n11824), .B2(n11773), .A(P2_B_REG_SCAN_IN), .ZN(n9752)
         );
  INV_X1 U12204 ( .A(n9752), .ZN(n9753) );
  NAND2_X1 U12205 ( .A1(n7497), .A2(n9753), .ZN(n9754) );
  NAND2_X1 U12206 ( .A1(n9755), .A2(n9754), .ZN(P2_U3328) );
  NAND2_X1 U12207 ( .A1(n9756), .A2(n10881), .ZN(n9757) );
  XNOR2_X1 U12208 ( .A(n12949), .B(n10670), .ZN(n12534) );
  NOR2_X1 U12209 ( .A1(n12534), .A2(n12773), .ZN(n12530) );
  AOI21_X1 U12210 ( .B1(n12534), .B2(n12773), .A(n12530), .ZN(n9851) );
  INV_X2 U12211 ( .A(n9761), .ZN(n9777) );
  XNOR2_X1 U12212 ( .A(n9838), .B(n15134), .ZN(n9776) );
  INV_X1 U12213 ( .A(n9759), .ZN(n10785) );
  OAI21_X1 U12214 ( .B1(n9760), .B2(n9764), .A(n8874), .ZN(n9762) );
  NAND2_X1 U12215 ( .A1(n9762), .A2(n9763), .ZN(n9770) );
  NAND2_X1 U12216 ( .A1(n9770), .A2(n9765), .ZN(n10673) );
  INV_X1 U12217 ( .A(n9770), .ZN(n9771) );
  INV_X1 U12218 ( .A(n9772), .ZN(n10884) );
  XNOR2_X1 U12219 ( .A(n9773), .B(n9772), .ZN(n10782) );
  OAI22_X1 U12220 ( .A1(n10781), .A2(n10782), .B1(n9773), .B2(n9772), .ZN(
        n10886) );
  XNOR2_X1 U12221 ( .A(n9777), .B(n15129), .ZN(n9774) );
  XNOR2_X1 U12222 ( .A(n9774), .B(n15091), .ZN(n10887) );
  NOR2_X1 U12223 ( .A1(n10885), .A2(n9775), .ZN(n10936) );
  XOR2_X1 U12224 ( .A(n12673), .B(n9776), .Z(n10937) );
  NAND2_X1 U12225 ( .A1(n10936), .A2(n10937), .ZN(n10935) );
  OAI21_X1 U12226 ( .B1(n9776), .B2(n12673), .A(n10935), .ZN(n11023) );
  XNOR2_X1 U12227 ( .A(n12528), .B(n15139), .ZN(n9778) );
  XOR2_X1 U12228 ( .A(n12672), .B(n9778), .Z(n11022) );
  NOR2_X1 U12229 ( .A1(n9778), .A2(n12672), .ZN(n9779) );
  XNOR2_X1 U12230 ( .A(n12528), .B(n9780), .ZN(n9781) );
  XNOR2_X1 U12231 ( .A(n9781), .B(n12671), .ZN(n11059) );
  NAND2_X1 U12232 ( .A1(n11060), .A2(n11059), .ZN(n11058) );
  INV_X1 U12233 ( .A(n9781), .ZN(n9782) );
  NAND2_X1 U12234 ( .A1(n9782), .A2(n12671), .ZN(n9783) );
  NAND2_X1 U12235 ( .A1(n11058), .A2(n9783), .ZN(n11283) );
  XNOR2_X1 U12236 ( .A(n12246), .B(n12528), .ZN(n11282) );
  NAND2_X1 U12237 ( .A1(n11283), .A2(n11282), .ZN(n11281) );
  INV_X1 U12238 ( .A(n11282), .ZN(n9784) );
  NAND2_X1 U12239 ( .A1(n9784), .A2(n12670), .ZN(n9785) );
  XNOR2_X1 U12240 ( .A(n12528), .B(n9786), .ZN(n9787) );
  XNOR2_X1 U12241 ( .A(n9787), .B(n12669), .ZN(n11357) );
  INV_X1 U12242 ( .A(n9787), .ZN(n9788) );
  NAND2_X1 U12243 ( .A1(n9788), .A2(n12669), .ZN(n9789) );
  XNOR2_X1 U12244 ( .A(n12528), .B(n15161), .ZN(n9790) );
  XNOR2_X1 U12245 ( .A(n9790), .B(n12668), .ZN(n11515) );
  INV_X1 U12246 ( .A(n11580), .ZN(n9792) );
  XNOR2_X1 U12247 ( .A(n12528), .B(n15167), .ZN(n9793) );
  XNOR2_X1 U12248 ( .A(n9793), .B(n12667), .ZN(n11579) );
  NAND2_X1 U12249 ( .A1(n9793), .A2(n12667), .ZN(n9794) );
  XNOR2_X1 U12250 ( .A(n12528), .B(n11836), .ZN(n9795) );
  XNOR2_X1 U12251 ( .A(n12281), .B(n9838), .ZN(n9796) );
  XOR2_X1 U12252 ( .A(n12665), .B(n9796), .Z(n11885) );
  NAND2_X1 U12253 ( .A1(n9796), .A2(n12280), .ZN(n9797) );
  XNOR2_X1 U12254 ( .A(n14407), .B(n12528), .ZN(n11924) );
  NOR2_X1 U12255 ( .A1(n11924), .A2(n12664), .ZN(n9804) );
  XNOR2_X1 U12256 ( .A(n12555), .B(n12528), .ZN(n9798) );
  NAND2_X1 U12257 ( .A1(n9798), .A2(n12663), .ZN(n9801) );
  INV_X1 U12258 ( .A(n9801), .ZN(n9799) );
  XOR2_X1 U12259 ( .A(n12663), .B(n9798), .Z(n12547) );
  INV_X1 U12260 ( .A(n9806), .ZN(n9802) );
  OR2_X1 U12261 ( .A1(n9804), .A2(n9802), .ZN(n9800) );
  NAND2_X1 U12262 ( .A1(n11924), .A2(n12664), .ZN(n12545) );
  AND2_X1 U12263 ( .A1(n12545), .A2(n9801), .ZN(n9805) );
  OR2_X1 U12264 ( .A1(n9802), .A2(n9805), .ZN(n9803) );
  AND2_X1 U12265 ( .A1(n9805), .A2(n12926), .ZN(n9807) );
  XNOR2_X1 U12266 ( .A(n12930), .B(n10670), .ZN(n12122) );
  NOR2_X1 U12267 ( .A1(n12122), .A2(n12661), .ZN(n12590) );
  XNOR2_X1 U12268 ( .A(n12598), .B(n9838), .ZN(n9808) );
  XNOR2_X1 U12269 ( .A(n9808), .B(n12660), .ZN(n12593) );
  INV_X1 U12270 ( .A(n12593), .ZN(n9810) );
  OR2_X1 U12271 ( .A1(n12590), .A2(n9810), .ZN(n9812) );
  INV_X1 U12272 ( .A(n9808), .ZN(n9809) );
  NAND2_X1 U12273 ( .A1(n12122), .A2(n12661), .ZN(n12591) );
  OAI21_X1 U12274 ( .B1(n12121), .B2(n9812), .A(n9811), .ZN(n12627) );
  XNOR2_X1 U12275 ( .A(n12635), .B(n9838), .ZN(n9813) );
  XNOR2_X1 U12276 ( .A(n9813), .B(n12886), .ZN(n12628) );
  NAND2_X1 U12277 ( .A1(n12627), .A2(n12628), .ZN(n9816) );
  INV_X1 U12278 ( .A(n9813), .ZN(n9814) );
  NAND2_X1 U12279 ( .A1(n9814), .A2(n12886), .ZN(n9815) );
  NAND2_X1 U12280 ( .A1(n9816), .A2(n9815), .ZN(n12562) );
  XNOR2_X1 U12281 ( .A(n13047), .B(n12528), .ZN(n9817) );
  NAND2_X1 U12282 ( .A1(n12562), .A2(n12563), .ZN(n9819) );
  NAND2_X1 U12283 ( .A1(n9817), .A2(n12659), .ZN(n9818) );
  NAND2_X1 U12284 ( .A1(n9819), .A2(n9818), .ZN(n12613) );
  XNOR2_X1 U12285 ( .A(n12877), .B(n9838), .ZN(n9820) );
  XNOR2_X1 U12286 ( .A(n9820), .B(n12887), .ZN(n12614) );
  INV_X1 U12287 ( .A(n9820), .ZN(n9821) );
  NAND2_X1 U12288 ( .A1(n9821), .A2(n12887), .ZN(n9822) );
  XNOR2_X1 U12289 ( .A(n12865), .B(n9838), .ZN(n9823) );
  NAND2_X1 U12290 ( .A1(n9823), .A2(n12874), .ZN(n9825) );
  OAI21_X1 U12291 ( .B1(n9823), .B2(n12874), .A(n9825), .ZN(n12572) );
  INV_X1 U12292 ( .A(n12572), .ZN(n9824) );
  NAND2_X1 U12293 ( .A1(n12569), .A2(n9825), .ZN(n9829) );
  INV_X1 U12294 ( .A(n9829), .ZN(n9827) );
  INV_X1 U12295 ( .A(n9828), .ZN(n9826) );
  NAND2_X1 U12296 ( .A1(n9829), .A2(n9828), .ZN(n9832) );
  INV_X1 U12297 ( .A(n9836), .ZN(n9834) );
  XNOR2_X1 U12298 ( .A(n12966), .B(n12528), .ZN(n9835) );
  INV_X1 U12299 ( .A(n9835), .ZN(n9833) );
  NAND2_X1 U12300 ( .A1(n9834), .A2(n9833), .ZN(n9837) );
  NAND2_X2 U12301 ( .A1(n9836), .A2(n9835), .ZN(n12601) );
  NAND2_X1 U12302 ( .A1(n12556), .A2(n12601), .ZN(n9842) );
  XNOR2_X1 U12303 ( .A(n12834), .B(n9838), .ZN(n9839) );
  NAND2_X1 U12304 ( .A1(n9839), .A2(n12842), .ZN(n12580) );
  INV_X1 U12305 ( .A(n9839), .ZN(n9840) );
  NAND2_X1 U12306 ( .A1(n9840), .A2(n12654), .ZN(n9841) );
  NAND2_X1 U12307 ( .A1(n9842), .A2(n12602), .ZN(n12579) );
  NAND2_X1 U12308 ( .A1(n12579), .A2(n12580), .ZN(n9846) );
  XNOR2_X1 U12309 ( .A(n12578), .B(n12528), .ZN(n9843) );
  NAND2_X1 U12310 ( .A1(n9843), .A2(n12829), .ZN(n9847) );
  INV_X1 U12311 ( .A(n9843), .ZN(n9844) );
  NAND2_X1 U12312 ( .A1(n9844), .A2(n12653), .ZN(n9845) );
  NAND2_X1 U12313 ( .A1(n9846), .A2(n12581), .ZN(n12583) );
  NAND2_X2 U12314 ( .A1(n12583), .A2(n9847), .ZN(n12640) );
  XNOR2_X1 U12315 ( .A(n9848), .B(n10670), .ZN(n9849) );
  NOR2_X1 U12316 ( .A1(n9849), .A2(n12652), .ZN(n9850) );
  AOI21_X1 U12317 ( .B1(n9849), .B2(n12652), .A(n9850), .ZN(n12641) );
  NAND2_X1 U12318 ( .A1(n9860), .A2(n15168), .ZN(n9853) );
  OR2_X1 U12319 ( .A1(n9866), .A2(n9857), .ZN(n9852) );
  NAND2_X1 U12320 ( .A1(n12380), .A2(n15150), .ZN(n9855) );
  OR2_X1 U12321 ( .A1(n9861), .A2(n9855), .ZN(n9856) );
  OAI211_X1 U12322 ( .C1(n12381), .C2(n12364), .A(n9892), .B(n10723), .ZN(
        n9859) );
  NOR2_X1 U12323 ( .A1(n9862), .A2(n9857), .ZN(n9858) );
  AOI211_X1 U12324 ( .C1(n9861), .C2(n9860), .A(n9859), .B(n9858), .ZN(n9865)
         );
  INV_X1 U12325 ( .A(n9862), .ZN(n9863) );
  NAND3_X1 U12326 ( .A1(n10691), .A2(n12380), .A3(n9863), .ZN(n9864) );
  INV_X1 U12327 ( .A(n12791), .ZN(n9868) );
  OR2_X1 U12328 ( .A1(n9866), .A2(n9883), .ZN(n11837) );
  AOI22_X1 U12329 ( .A1(n15104), .A2(n12651), .B1(n12652), .B2(n15103), .ZN(
        n12787) );
  OAI22_X1 U12330 ( .A1(n11837), .A2(n12787), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15303), .ZN(n9867) );
  AOI21_X1 U12331 ( .B1(n12629), .B2(n9868), .A(n9867), .ZN(n9869) );
  OAI21_X1 U12332 ( .B1(n9870), .B2(n12649), .A(n9869), .ZN(n9871) );
  INV_X1 U12333 ( .A(n9871), .ZN(n9872) );
  NAND2_X1 U12334 ( .A1(n9873), .A2(n9872), .ZN(P3_U3154) );
  XNOR2_X1 U12335 ( .A(n9874), .B(n10893), .ZN(n9877) );
  NAND2_X1 U12336 ( .A1(n9875), .A2(n12380), .ZN(n9876) );
  NAND2_X1 U12337 ( .A1(n8454), .A2(n12384), .ZN(n9878) );
  OAI21_X1 U12338 ( .B1(n9879), .B2(n15168), .A(n9878), .ZN(n9880) );
  NAND2_X1 U12339 ( .A1(n9880), .A2(n9883), .ZN(n9881) );
  NAND2_X1 U12340 ( .A1(n9881), .A2(n12364), .ZN(n9882) );
  NAND2_X1 U12341 ( .A1(n9882), .A2(n10893), .ZN(n9885) );
  MUX2_X1 U12342 ( .A(n10891), .B(n9883), .S(n12370), .Z(n10894) );
  NAND2_X1 U12343 ( .A1(n10894), .A2(n13062), .ZN(n9884) );
  NAND2_X1 U12344 ( .A1(n9889), .A2(n7482), .ZN(P3_U3488) );
  INV_X1 U12345 ( .A(n9890), .ZN(n10099) );
  NOR2_X1 U12346 ( .A1(n9891), .A2(n10099), .ZN(n10102) );
  NOR2_X4 U12347 ( .A1(n9892), .A2(n10090), .ZN(P3_U3897) );
  AND2_X2 U12348 ( .A1(n10472), .A2(n10456), .ZN(P1_U4016) );
  NAND2_X1 U12349 ( .A1(n9894), .A2(n9893), .ZN(n9896) );
  NAND2_X1 U12350 ( .A1(n9896), .A2(n9895), .ZN(n11113) );
  NAND2_X1 U12351 ( .A1(n11113), .A2(n11111), .ZN(n9898) );
  NAND2_X1 U12352 ( .A1(n9898), .A2(n9897), .ZN(n14668) );
  NAND2_X1 U12353 ( .A1(n14668), .A2(n9899), .ZN(n9901) );
  NAND2_X1 U12354 ( .A1(n9960), .A2(n14676), .ZN(n9900) );
  NAND2_X1 U12355 ( .A1(n9901), .A2(n9900), .ZN(n14651) );
  NAND2_X1 U12356 ( .A1(n13728), .A2(n13765), .ZN(n9902) );
  NAND2_X1 U12357 ( .A1(n13839), .A2(n11494), .ZN(n9903) );
  INV_X1 U12358 ( .A(n13838), .ZN(n11497) );
  NAND2_X1 U12359 ( .A1(n14638), .A2(n9971), .ZN(n9906) );
  INV_X1 U12360 ( .A(n13837), .ZN(n9904) );
  NAND2_X1 U12361 ( .A1(n14647), .A2(n9904), .ZN(n9905) );
  NAND2_X1 U12362 ( .A1(n9906), .A2(n9905), .ZN(n11106) );
  INV_X1 U12363 ( .A(n13836), .ZN(n11425) );
  OR2_X1 U12364 ( .A1(n11589), .A2(n11425), .ZN(n9908) );
  INV_X1 U12365 ( .A(n11423), .ZN(n9973) );
  INV_X1 U12366 ( .A(n14627), .ZN(n14621) );
  INV_X1 U12367 ( .A(n13835), .ZN(n9909) );
  NAND2_X1 U12368 ( .A1(n11674), .A2(n9909), .ZN(n14616) );
  AND2_X1 U12369 ( .A1(n14621), .A2(n14616), .ZN(n9910) );
  NAND2_X1 U12370 ( .A1(n9911), .A2(n11659), .ZN(n11664) );
  INV_X1 U12371 ( .A(n14630), .ZN(n11906) );
  OR2_X1 U12372 ( .A1(n11656), .A2(n11906), .ZN(n9912) );
  NAND2_X1 U12373 ( .A1(n11664), .A2(n9912), .ZN(n11689) );
  NAND2_X1 U12374 ( .A1(n11689), .A2(n11688), .ZN(n11687) );
  INV_X1 U12375 ( .A(n13833), .ZN(n11962) );
  OR2_X1 U12376 ( .A1(n11900), .A2(n11962), .ZN(n9913) );
  NAND2_X1 U12377 ( .A1(n11687), .A2(n9913), .ZN(n11819) );
  NAND2_X1 U12378 ( .A1(n11819), .A2(n11818), .ZN(n11817) );
  OR2_X1 U12379 ( .A1(n14518), .A2(n12003), .ZN(n9914) );
  NAND2_X1 U12380 ( .A1(n11869), .A2(n9917), .ZN(n11943) );
  NAND2_X1 U12381 ( .A1(n13719), .A2(n13741), .ZN(n9918) );
  INV_X1 U12382 ( .A(n14074), .ZN(n13786) );
  OR2_X1 U12383 ( .A1(n13734), .A2(n13786), .ZN(n9920) );
  NAND2_X1 U12384 ( .A1(n14073), .A2(n14072), .ZN(n14071) );
  OR2_X1 U12385 ( .A1(n14172), .A2(n14054), .ZN(n9921) );
  INV_X1 U12386 ( .A(n14075), .ZN(n9922) );
  NAND2_X1 U12387 ( .A1(n14062), .A2(n9922), .ZN(n9923) );
  NAND2_X1 U12388 ( .A1(n14023), .A2(n14022), .ZN(n14021) );
  NAND2_X1 U12389 ( .A1(n14029), .A2(n13827), .ZN(n9924) );
  INV_X1 U12390 ( .A(n13691), .ZN(n13826) );
  OR2_X1 U12391 ( .A1(n8295), .A2(n13826), .ZN(n9925) );
  INV_X1 U12392 ( .A(n13825), .ZN(n13753) );
  NAND2_X1 U12393 ( .A1(n14138), .A2(n13753), .ZN(n9926) );
  NAND2_X1 U12394 ( .A1(n9927), .A2(n9926), .ZN(n13972) );
  INV_X1 U12395 ( .A(n13972), .ZN(n9929) );
  INV_X1 U12396 ( .A(n13983), .ZN(n9928) );
  NAND2_X1 U12397 ( .A1(n13981), .A2(n13824), .ZN(n9930) );
  OAI21_X1 U12398 ( .B1(n6608), .B2(n10004), .A(n12011), .ZN(n9933) );
  OR2_X1 U12399 ( .A1(n8333), .A2(n10010), .ZN(n9931) );
  NAND2_X1 U12400 ( .A1(n9933), .A2(n14618), .ZN(n14131) );
  NAND2_X1 U12401 ( .A1(n13822), .A2(n14631), .ZN(n9935) );
  NAND2_X1 U12402 ( .A1(n13824), .A2(n14482), .ZN(n9934) );
  NAND2_X1 U12403 ( .A1(n9935), .A2(n9934), .ZN(n14124) );
  INV_X1 U12404 ( .A(n14124), .ZN(n9956) );
  OR2_X2 U12405 ( .A1(n9936), .A2(n14215), .ZN(n14688) );
  NOR2_X4 U12406 ( .A1(n14688), .A2(n9937), .ZN(n14679) );
  INV_X1 U12407 ( .A(n11232), .ZN(n10463) );
  NAND2_X1 U12408 ( .A1(n11881), .A2(P1_B_REG_SCAN_IN), .ZN(n9939) );
  INV_X1 U12409 ( .A(P1_B_REG_SCAN_IN), .ZN(n12488) );
  NAND2_X1 U12410 ( .A1(n9950), .A2(n12488), .ZN(n9938) );
  NAND2_X2 U12411 ( .A1(n11232), .A2(n10461), .ZN(n14687) );
  NOR4_X1 U12412 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n9948) );
  NOR4_X1 U12413 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n9947) );
  OR4_X1 U12414 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n9945) );
  NOR4_X1 U12415 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n9943) );
  NOR4_X1 U12416 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n9942) );
  NOR4_X1 U12417 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9941) );
  NOR4_X1 U12418 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n9940) );
  NAND4_X1 U12419 ( .A1(n9943), .A2(n9942), .A3(n9941), .A4(n9940), .ZN(n9944)
         );
  NOR4_X1 U12420 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n9945), .A4(n9944), .ZN(n9946) );
  AND3_X1 U12421 ( .A1(n9948), .A2(n9947), .A3(n9946), .ZN(n10460) );
  NAND2_X1 U12422 ( .A1(n11232), .A2(n10460), .ZN(n9949) );
  NAND2_X1 U12423 ( .A1(n14687), .A2(n9949), .ZN(n9954) );
  OR2_X1 U12424 ( .A1(n10461), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9951) );
  OR2_X1 U12425 ( .A1(n10461), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9952) );
  OR2_X1 U12426 ( .A1(n11987), .A2(n14210), .ZN(n10045) );
  NAND2_X1 U12427 ( .A1(n9952), .A2(n10045), .ZN(n11231) );
  NOR2_X1 U12428 ( .A1(n11254), .A2(n11231), .ZN(n9953) );
  AND2_X1 U12429 ( .A1(n9954), .A2(n9953), .ZN(n9955) );
  NAND2_X1 U12430 ( .A1(n9955), .A2(n11233), .ZN(n12490) );
  INV_X1 U12431 ( .A(n14665), .ZN(n14644) );
  AOI21_X1 U12432 ( .B1(n14131), .B2(n9956), .A(n14644), .ZN(n10016) );
  NAND2_X1 U12433 ( .A1(n11150), .A2(n14698), .ZN(n9957) );
  INV_X1 U12434 ( .A(n11111), .ZN(n11114) );
  NAND2_X1 U12435 ( .A1(n11112), .A2(n11114), .ZN(n9959) );
  NAND2_X1 U12436 ( .A1(n10641), .A2(n14705), .ZN(n9958) );
  NAND2_X1 U12437 ( .A1(n9959), .A2(n9958), .ZN(n14667) );
  NAND2_X1 U12438 ( .A1(n14667), .A2(n14669), .ZN(n9962) );
  INV_X1 U12439 ( .A(n14676), .ZN(n14711) );
  NAND2_X1 U12440 ( .A1(n9960), .A2(n14711), .ZN(n9961) );
  INV_X1 U12441 ( .A(n9963), .ZN(n14659) );
  NAND2_X1 U12442 ( .A1(n14658), .A2(n14659), .ZN(n9965) );
  NAND2_X1 U12443 ( .A1(n13728), .A2(n14718), .ZN(n9964) );
  NAND2_X1 U12444 ( .A1(n9965), .A2(n9964), .ZN(n11171) );
  NAND2_X1 U12445 ( .A1(n11171), .A2(n11172), .ZN(n9967) );
  INV_X1 U12446 ( .A(n13839), .ZN(n11495) );
  NAND2_X1 U12447 ( .A1(n11495), .A2(n11494), .ZN(n9966) );
  INV_X1 U12448 ( .A(n11140), .ZN(n9968) );
  NAND2_X1 U12449 ( .A1(n11138), .A2(n9968), .ZN(n9970) );
  NAND2_X1 U12450 ( .A1(n14732), .A2(n11497), .ZN(n9969) );
  OR2_X1 U12451 ( .A1(n14647), .A2(n13837), .ZN(n9972) );
  NAND2_X1 U12452 ( .A1(n11422), .A2(n9973), .ZN(n9975) );
  OR2_X1 U12453 ( .A1(n11674), .A2(n13835), .ZN(n9974) );
  NAND2_X1 U12454 ( .A1(n9975), .A2(n9974), .ZN(n14626) );
  NAND2_X1 U12455 ( .A1(n14626), .A2(n14627), .ZN(n9977) );
  OR2_X1 U12456 ( .A1(n14628), .A2(n13834), .ZN(n9976) );
  INV_X1 U12457 ( .A(n11659), .ZN(n11651) );
  OR2_X1 U12458 ( .A1(n11656), .A2(n14630), .ZN(n9978) );
  INV_X1 U12459 ( .A(n11688), .ZN(n9979) );
  INV_X1 U12460 ( .A(n11818), .ZN(n11808) );
  NAND2_X1 U12461 ( .A1(n11807), .A2(n11808), .ZN(n9981) );
  OR2_X1 U12462 ( .A1(n14518), .A2(n14483), .ZN(n9980) );
  NAND2_X1 U12463 ( .A1(n9981), .A2(n9980), .ZN(n14473) );
  INV_X1 U12464 ( .A(n13807), .ZN(n13832) );
  NAND2_X1 U12465 ( .A1(n14511), .A2(n13832), .ZN(n9982) );
  INV_X1 U12466 ( .A(n13714), .ZN(n13831) );
  NAND2_X1 U12467 ( .A1(n11947), .A2(n11948), .ZN(n9984) );
  OR2_X1 U12468 ( .A1(n13719), .A2(n13830), .ZN(n9983) );
  INV_X1 U12469 ( .A(n9985), .ZN(n9986) );
  INV_X1 U12470 ( .A(n9988), .ZN(n9990) );
  NAND2_X1 U12471 ( .A1(n14050), .A2(n14051), .ZN(n9992) );
  OR2_X1 U12472 ( .A1(n14062), .A2(n14075), .ZN(n9991) );
  INV_X1 U12473 ( .A(n14033), .ZN(n14039) );
  NAND2_X1 U12474 ( .A1(n14159), .A2(n13828), .ZN(n9993) );
  INV_X1 U12475 ( .A(n14020), .ZN(n9995) );
  INV_X1 U12476 ( .A(n13827), .ZN(n9996) );
  NAND2_X1 U12477 ( .A1(n14029), .A2(n9996), .ZN(n9997) );
  INV_X1 U12478 ( .A(n14006), .ZN(n9998) );
  NAND2_X1 U12479 ( .A1(n14138), .A2(n13825), .ZN(n9999) );
  NAND2_X1 U12480 ( .A1(n13981), .A2(n13705), .ZN(n10000) );
  INV_X1 U12481 ( .A(n10004), .ZN(n10001) );
  OR2_X1 U12482 ( .A1(n10453), .A2(n10002), .ZN(n10003) );
  NAND2_X1 U12483 ( .A1(n6585), .A2(n10004), .ZN(n14127) );
  AND3_X1 U12484 ( .A1(n14126), .A2(n14662), .A3(n14127), .ZN(n10015) );
  OR2_X1 U12485 ( .A1(n6493), .A2(n14694), .ZN(n11118) );
  NOR2_X1 U12486 ( .A1(n11118), .A2(n11119), .ZN(n14681) );
  NAND2_X1 U12487 ( .A1(n14678), .A2(n14718), .ZN(n14660) );
  NOR2_X1 U12488 ( .A1(n11427), .A2(n11674), .ZN(n14629) );
  INV_X1 U12489 ( .A(n14628), .ZN(n14756) );
  AND2_X1 U12490 ( .A1(n14629), .A2(n14756), .ZN(n11652) );
  INV_X1 U12491 ( .A(n11900), .ZN(n14337) );
  INV_X1 U12492 ( .A(n14503), .ZN(n12057) );
  NAND2_X1 U12493 ( .A1(n8295), .A2(n14027), .ZN(n14008) );
  NAND2_X1 U12494 ( .A1(n14125), .A2(n13976), .ZN(n10007) );
  NAND2_X1 U12495 ( .A1(n10007), .A2(n14679), .ZN(n10008) );
  OR2_X1 U12496 ( .A1(n6531), .A2(n10008), .ZN(n14128) );
  INV_X1 U12497 ( .A(n14673), .ZN(n14643) );
  AOI22_X1 U12498 ( .A1(n13703), .A2(n14643), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n14087), .ZN(n10013) );
  INV_X1 U12499 ( .A(n10009), .ZN(n10011) );
  NAND2_X1 U12500 ( .A1(n10011), .A2(n10010), .ZN(n14655) );
  INV_X1 U12501 ( .A(n14655), .ZN(n10465) );
  NAND2_X1 U12502 ( .A1(n14125), .A2(n14677), .ZN(n10012) );
  OAI211_X1 U12503 ( .C1(n14128), .C2(n14065), .A(n10013), .B(n10012), .ZN(
        n10014) );
  OR3_X1 U12504 ( .A1(n10016), .A2(n10015), .A3(n10014), .ZN(P1_U3268) );
  NAND2_X1 U12505 ( .A1(n10022), .A2(P1_U3086), .ZN(n14208) );
  INV_X1 U12506 ( .A(n14208), .ZN(n11826) );
  INV_X1 U12507 ( .A(n11826), .ZN(n14214) );
  INV_X1 U12508 ( .A(n10017), .ZN(n10061) );
  AND2_X1 U12509 ( .A1(n8119), .A2(P1_U3086), .ZN(n14202) );
  INV_X2 U12510 ( .A(n14202), .ZN(n12044) );
  OAI222_X1 U12511 ( .A1(n14214), .A2(n10061), .B1(n13868), .B2(P1_U3086), 
        .C1(n10018), .C2(n12044), .ZN(P1_U3353) );
  INV_X1 U12512 ( .A(n10019), .ZN(n10059) );
  OAI222_X1 U12513 ( .A1(n14214), .A2(n10059), .B1(n14575), .B2(P1_U3086), 
        .C1(n10020), .C2(n12044), .ZN(P1_U3351) );
  OAI222_X1 U12514 ( .A1(n12044), .A2(n10021), .B1(n13847), .B2(P1_U3086), 
        .C1(n14214), .C2(n10023), .ZN(P1_U3354) );
  OAI222_X1 U12515 ( .A1(n13652), .A2(n10024), .B1(n13643), .B2(n10023), .C1(
        P2_U3088), .C2(n10314), .ZN(P2_U3326) );
  OAI222_X1 U12516 ( .A1(n14214), .A2(n10063), .B1(n10198), .B2(P1_U3086), 
        .C1(n10025), .C2(n12044), .ZN(P1_U3350) );
  NOR2_X1 U12517 ( .A1(n8119), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13070) );
  OAI222_X1 U12518 ( .A1(n13076), .A2(n10027), .B1(n13078), .B2(n10026), .C1(
        n14976), .C2(P3_U3151), .ZN(P3_U3292) );
  INV_X1 U12519 ( .A(n10028), .ZN(n10030) );
  OAI222_X1 U12520 ( .A1(n13076), .A2(n10030), .B1(n13078), .B2(n10029), .C1(
        n10834), .C2(P3_U3151), .ZN(P3_U3293) );
  INV_X1 U12521 ( .A(n10031), .ZN(n10032) );
  INV_X1 U12522 ( .A(SI_4_), .ZN(n15281) );
  OAI222_X1 U12523 ( .A1(n13076), .A2(n10032), .B1(n13078), .B2(n15281), .C1(
        n15005), .C2(P3_U3151), .ZN(P3_U3291) );
  INV_X1 U12524 ( .A(n10033), .ZN(n10035) );
  OAI222_X1 U12525 ( .A1(n6849), .A2(P3_U3151), .B1(n13076), .B2(n10035), .C1(
        n10034), .C2(n13078), .ZN(P3_U3295) );
  INV_X1 U12526 ( .A(n10858), .ZN(n10866) );
  INV_X1 U12527 ( .A(n10036), .ZN(n10037) );
  OAI222_X1 U12528 ( .A1(n10866), .A2(P3_U3151), .B1(n13076), .B2(n10037), 
        .C1(n15331), .C2(n13078), .ZN(P3_U3289) );
  INV_X1 U12529 ( .A(n10038), .ZN(n10057) );
  OAI222_X1 U12530 ( .A1(n12044), .A2(n10039), .B1(n14214), .B2(n10057), .C1(
        P1_U3086), .C2(n13879), .ZN(P1_U3352) );
  INV_X1 U12531 ( .A(n10161), .ZN(n10242) );
  OAI222_X1 U12532 ( .A1(n14214), .A2(n10065), .B1(n10242), .B2(P1_U3086), 
        .C1(n10040), .C2(n12044), .ZN(P1_U3349) );
  OAI222_X1 U12533 ( .A1(n13076), .A2(n10041), .B1(n13078), .B2(n15248), .C1(
        n11390), .C2(P3_U3151), .ZN(P3_U3285) );
  INV_X1 U12534 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10044) );
  INV_X1 U12535 ( .A(n10042), .ZN(n10043) );
  AOI22_X1 U12536 ( .A1(n14687), .A2(n10044), .B1(n10472), .B2(n10043), .ZN(
        P1_U3445) );
  INV_X1 U12537 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10047) );
  INV_X1 U12538 ( .A(n10045), .ZN(n10046) );
  AOI22_X1 U12539 ( .A1(n14687), .A2(n10047), .B1(n10472), .B2(n10046), .ZN(
        P1_U3446) );
  INV_X1 U12540 ( .A(SI_7_), .ZN(n15250) );
  OAI222_X1 U12541 ( .A1(n13076), .A2(n10048), .B1(n13078), .B2(n15250), .C1(
        n15035), .C2(P3_U3151), .ZN(P3_U3288) );
  INV_X1 U12542 ( .A(SI_9_), .ZN(n15268) );
  OAI222_X1 U12543 ( .A1(n13076), .A2(n10049), .B1(n13078), .B2(n15268), .C1(
        n15053), .C2(P3_U3151), .ZN(P3_U3286) );
  INV_X1 U12544 ( .A(n10050), .ZN(n10052) );
  INV_X1 U12545 ( .A(SI_5_), .ZN(n10051) );
  OAI222_X1 U12546 ( .A1(n13076), .A2(n10052), .B1(n13078), .B2(n10051), .C1(
        n15023), .C2(P3_U3151), .ZN(P3_U3290) );
  OAI222_X1 U12547 ( .A1(n13076), .A2(n10053), .B1(n13078), .B2(n15379), .C1(
        n6839), .C2(P3_U3151), .ZN(P3_U3287) );
  OAI222_X1 U12548 ( .A1(n13076), .A2(n10054), .B1(n11556), .B2(P3_U3151), 
        .C1(n13078), .C2(n15315), .ZN(P3_U3284) );
  NAND2_X1 U12549 ( .A1(n9477), .A2(P2_U3947), .ZN(n10055) );
  OAI21_X1 U12550 ( .B1(n8491), .B2(P2_U3947), .A(n10055), .ZN(P2_U3531) );
  INV_X1 U12551 ( .A(n10333), .ZN(n10341) );
  OAI222_X1 U12552 ( .A1(n10341), .A2(P2_U3088), .B1(n13643), .B2(n10057), 
        .C1(n10056), .C2(n13652), .ZN(P2_U3324) );
  OAI222_X1 U12553 ( .A1(P2_U3088), .A2(n14796), .B1(n13643), .B2(n10059), 
        .C1(n10058), .C2(n13652), .ZN(P2_U3323) );
  INV_X1 U12554 ( .A(n10289), .ZN(n10126) );
  OAI222_X1 U12555 ( .A1(P2_U3088), .A2(n10126), .B1(n13643), .B2(n10061), 
        .C1(n10060), .C2(n13652), .ZN(P2_U3325) );
  INV_X1 U12556 ( .A(n10347), .ZN(n10353) );
  OAI222_X1 U12557 ( .A1(P2_U3088), .A2(n10353), .B1(n13643), .B2(n10063), 
        .C1(n10062), .C2(n13652), .ZN(P2_U3322) );
  INV_X1 U12558 ( .A(n13278), .ZN(n10066) );
  OAI222_X1 U12559 ( .A1(P2_U3088), .A2(n10066), .B1(n13643), .B2(n10065), 
        .C1(n10064), .C2(n13652), .ZN(P2_U3321) );
  OAI222_X1 U12560 ( .A1(P3_U3151), .A2(n10753), .B1(n13078), .B2(n7562), .C1(
        n13076), .C2(n10067), .ZN(P3_U3294) );
  INV_X1 U12561 ( .A(n13890), .ZN(n10069) );
  OAI222_X1 U12562 ( .A1(n14214), .A2(n10071), .B1(n10069), .B2(P1_U3086), 
        .C1(n10068), .C2(n12044), .ZN(P1_U3348) );
  INV_X1 U12563 ( .A(n13293), .ZN(n10072) );
  OAI222_X1 U12564 ( .A1(P2_U3088), .A2(n10072), .B1(n13643), .B2(n10071), 
        .C1(n10070), .C2(n13652), .ZN(P2_U3320) );
  OAI222_X1 U12565 ( .A1(n14214), .A2(n10077), .B1(n10178), .B2(P1_U3086), 
        .C1(n10073), .C2(n12044), .ZN(P1_U3347) );
  INV_X1 U12566 ( .A(n10074), .ZN(n10075) );
  INV_X1 U12567 ( .A(n11791), .ZN(n11793) );
  OAI222_X1 U12568 ( .A1(n13076), .A2(n10075), .B1(n11793), .B2(P3_U3151), 
        .C1(n15312), .C2(n13078), .ZN(P3_U3283) );
  INV_X1 U12569 ( .A(n10415), .ZN(n10309) );
  OAI222_X1 U12570 ( .A1(P2_U3088), .A2(n10309), .B1(n13643), .B2(n10077), 
        .C1(n10076), .C2(n13652), .ZN(P2_U3319) );
  OR2_X1 U12571 ( .A1(n10464), .A2(n10078), .ZN(n10080) );
  NAND2_X1 U12572 ( .A1(n10080), .A2(n10079), .ZN(n10150) );
  NOR2_X1 U12573 ( .A1(n11232), .A2(n8324), .ZN(n10149) );
  INV_X1 U12574 ( .A(n10149), .ZN(n10081) );
  AND2_X1 U12575 ( .A1(n10150), .A2(n10081), .ZN(n14587) );
  NOR2_X1 U12576 ( .A1(n14587), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U12577 ( .A(n10384), .ZN(n10083) );
  OAI222_X1 U12578 ( .A1(n14214), .A2(n10085), .B1(n10083), .B2(P1_U3086), 
        .C1(n10082), .C2(n12044), .ZN(P1_U3346) );
  INV_X1 U12579 ( .A(n10418), .ZN(n14821) );
  OAI222_X1 U12580 ( .A1(P2_U3088), .A2(n14821), .B1(n13643), .B2(n10085), 
        .C1(n10084), .C2(n13652), .ZN(P2_U3318) );
  OAI222_X1 U12581 ( .A1(n13076), .A2(n10086), .B1(n13078), .B2(n15261), .C1(
        n12680), .C2(P3_U3151), .ZN(P3_U3282) );
  INV_X1 U12582 ( .A(n10432), .ZN(n10442) );
  OAI222_X1 U12583 ( .A1(n14208), .A2(n10089), .B1(n10442), .B2(P1_U3086), 
        .C1(n10087), .C2(n12044), .ZN(P1_U3345) );
  INV_X1 U12584 ( .A(n10795), .ZN(n10425) );
  OAI222_X1 U12585 ( .A1(P2_U3088), .A2(n10425), .B1(n13643), .B2(n10089), 
        .C1(n10088), .C2(n13652), .ZN(P2_U3317) );
  INV_X1 U12586 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10091) );
  NOR2_X1 U12587 ( .A1(n10548), .A2(n10091), .ZN(P3_U3251) );
  INV_X1 U12588 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10092) );
  NOR2_X1 U12589 ( .A1(n10548), .A2(n10092), .ZN(P3_U3249) );
  INV_X1 U12590 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10093) );
  NOR2_X1 U12591 ( .A1(n10548), .A2(n10093), .ZN(P3_U3250) );
  INV_X1 U12592 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10094) );
  NOR2_X1 U12593 ( .A1(n10548), .A2(n10094), .ZN(P3_U3247) );
  INV_X1 U12594 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10095) );
  NOR2_X1 U12595 ( .A1(n10548), .A2(n10095), .ZN(P3_U3248) );
  INV_X1 U12596 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10096) );
  NOR2_X1 U12597 ( .A1(n10548), .A2(n10096), .ZN(P3_U3259) );
  OAI222_X1 U12598 ( .A1(n13076), .A2(n10097), .B1(n13078), .B2(n15263), .C1(
        n12700), .C2(P3_U3151), .ZN(P3_U3281) );
  OAI21_X1 U12599 ( .B1(n10219), .B2(n10099), .A(n10098), .ZN(n10100) );
  INV_X1 U12600 ( .A(n10100), .ZN(n10101) );
  OR2_X1 U12601 ( .A1(n10102), .A2(n10101), .ZN(n10108) );
  AND2_X1 U12602 ( .A1(n10107), .A2(n10108), .ZN(n14795) );
  AND2_X1 U12603 ( .A1(n14795), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14873) );
  OR2_X1 U12604 ( .A1(n10108), .A2(P2_U3088), .ZN(n14832) );
  INV_X1 U12605 ( .A(n14832), .ZN(n14871) );
  NOR2_X1 U12606 ( .A1(n10979), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10114) );
  INV_X1 U12607 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10378) );
  MUX2_X1 U12608 ( .A(n10378), .B(P2_REG1_REG_1__SCAN_IN), .S(n10314), .Z(
        n10104) );
  AND2_X1 U12609 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n10103) );
  NAND2_X1 U12610 ( .A1(n10104), .A2(n10103), .ZN(n10318) );
  OAI21_X1 U12611 ( .B1(n10378), .B2(n10314), .A(n10318), .ZN(n10105) );
  INV_X1 U12612 ( .A(n10105), .ZN(n10112) );
  INV_X1 U12613 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10370) );
  MUX2_X1 U12614 ( .A(n10370), .B(P2_REG1_REG_2__SCAN_IN), .S(n10289), .Z(
        n10111) );
  MUX2_X1 U12615 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n10370), .S(n10289), .Z(
        n10106) );
  NAND2_X1 U12616 ( .A1(n10106), .A2(n10105), .ZN(n10328) );
  INV_X1 U12617 ( .A(n10328), .ZN(n10110) );
  NOR2_X1 U12618 ( .A1(n10107), .A2(P2_U3088), .ZN(n13644) );
  INV_X1 U12619 ( .A(n10116), .ZN(n10109) );
  INV_X1 U12620 ( .A(n13650), .ZN(n10115) );
  AOI211_X1 U12621 ( .C1(n10112), .C2(n10111), .A(n10110), .B(n14862), .ZN(
        n10113) );
  AOI211_X1 U12622 ( .C1(n14871), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n10114), .B(
        n10113), .ZN(n10125) );
  MUX2_X1 U12623 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10117), .S(n10289), .Z(
        n10120) );
  MUX2_X1 U12624 ( .A(n10947), .B(P2_REG2_REG_1__SCAN_IN), .S(n10314), .Z(
        n10311) );
  AND2_X1 U12625 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n10118) );
  NAND2_X1 U12626 ( .A1(n10311), .A2(n10118), .ZN(n10312) );
  INV_X1 U12627 ( .A(n10314), .ZN(n10321) );
  NAND2_X1 U12628 ( .A1(n10321), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10121) );
  NAND2_X1 U12629 ( .A1(n10312), .A2(n10121), .ZN(n10119) );
  NAND2_X1 U12630 ( .A1(n10120), .A2(n10119), .ZN(n10336) );
  MUX2_X1 U12631 ( .A(n10117), .B(P2_REG2_REG_2__SCAN_IN), .S(n10289), .Z(
        n10122) );
  NAND3_X1 U12632 ( .A1(n10122), .A2(n10312), .A3(n10121), .ZN(n10123) );
  NAND3_X1 U12633 ( .A1(n14875), .A2(n10336), .A3(n10123), .ZN(n10124) );
  OAI211_X1 U12634 ( .C1(n14822), .C2(n10126), .A(n10125), .B(n10124), .ZN(
        P2_U3216) );
  MUX2_X1 U12635 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10127), .S(n10178), .Z(
        n10148) );
  INV_X1 U12636 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10128) );
  MUX2_X1 U12637 ( .A(n10128), .B(P1_REG1_REG_1__SCAN_IN), .S(n13847), .Z(
        n10130) );
  AND2_X1 U12638 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n10129) );
  NAND2_X1 U12639 ( .A1(n10130), .A2(n10129), .ZN(n13851) );
  INV_X1 U12640 ( .A(n13847), .ZN(n13846) );
  NAND2_X1 U12641 ( .A1(n13846), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10131) );
  NAND2_X1 U12642 ( .A1(n13851), .A2(n10131), .ZN(n13862) );
  INV_X1 U12643 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10132) );
  MUX2_X1 U12644 ( .A(n10132), .B(P1_REG1_REG_2__SCAN_IN), .S(n13868), .Z(
        n13863) );
  NAND2_X1 U12645 ( .A1(n13862), .A2(n13863), .ZN(n13877) );
  INV_X1 U12646 ( .A(n13868), .ZN(n10157) );
  NAND2_X1 U12647 ( .A1(n10157), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n13876) );
  NAND2_X1 U12648 ( .A1(n13877), .A2(n13876), .ZN(n10134) );
  MUX2_X1 U12649 ( .A(n10135), .B(P1_REG1_REG_3__SCAN_IN), .S(n13879), .Z(
        n10133) );
  NAND2_X1 U12650 ( .A1(n10134), .A2(n10133), .ZN(n14577) );
  OR2_X1 U12651 ( .A1(n13879), .A2(n10135), .ZN(n14576) );
  NAND2_X1 U12652 ( .A1(n14577), .A2(n14576), .ZN(n10138) );
  MUX2_X1 U12653 ( .A(n10136), .B(P1_REG1_REG_4__SCAN_IN), .S(n14575), .Z(
        n10137) );
  NAND2_X1 U12654 ( .A1(n10138), .A2(n10137), .ZN(n14580) );
  INV_X1 U12655 ( .A(n14575), .ZN(n14574) );
  NAND2_X1 U12656 ( .A1(n14574), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10139) );
  AND2_X1 U12657 ( .A1(n14580), .A2(n10139), .ZN(n10187) );
  INV_X1 U12658 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n14768) );
  MUX2_X1 U12659 ( .A(n14768), .B(P1_REG1_REG_5__SCAN_IN), .S(n10198), .Z(
        n10188) );
  NAND2_X1 U12660 ( .A1(n10187), .A2(n10188), .ZN(n10186) );
  NAND2_X1 U12661 ( .A1(n10198), .A2(n14768), .ZN(n10140) );
  AND2_X1 U12662 ( .A1(n10186), .A2(n10140), .ZN(n10232) );
  MUX2_X1 U12663 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10141), .S(n10161), .Z(
        n10231) );
  NAND2_X1 U12664 ( .A1(n10232), .A2(n10231), .ZN(n13893) );
  NAND2_X1 U12665 ( .A1(n10161), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n13892) );
  NAND2_X1 U12666 ( .A1(n13893), .A2(n13892), .ZN(n10144) );
  INV_X1 U12667 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10142) );
  MUX2_X1 U12668 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n10142), .S(n13890), .Z(
        n10143) );
  NAND2_X1 U12669 ( .A1(n10144), .A2(n10143), .ZN(n13895) );
  NAND2_X1 U12670 ( .A1(n13890), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10145) );
  NAND2_X1 U12671 ( .A1(n13895), .A2(n10145), .ZN(n10147) );
  INV_X1 U12672 ( .A(n10174), .ZN(n10146) );
  AOI21_X1 U12673 ( .B1(n10148), .B2(n10147), .A(n10146), .ZN(n10169) );
  OR2_X1 U12674 ( .A1(n10150), .A2(n10149), .ZN(n14565) );
  NOR2_X2 U12675 ( .A1(n14565), .A2(n14562), .ZN(n14603) );
  INV_X1 U12676 ( .A(n14603), .ZN(n11090) );
  NOR2_X1 U12677 ( .A1(n14565), .A2(n13859), .ZN(n14591) );
  INV_X1 U12678 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n14238) );
  NAND2_X1 U12679 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n11605) );
  OAI21_X1 U12680 ( .B1(n14615), .B2(n14238), .A(n11605), .ZN(n10151) );
  AOI21_X1 U12681 ( .B1(n10152), .B2(n14591), .A(n10151), .ZN(n10168) );
  OR2_X1 U12682 ( .A1(n8325), .A2(n14206), .ZN(n10153) );
  OR2_X1 U12683 ( .A1(n14565), .A2(n10153), .ZN(n13920) );
  MUX2_X1 U12684 ( .A(n10154), .B(P1_REG2_REG_1__SCAN_IN), .S(n13847), .Z(
        n13845) );
  AND2_X1 U12685 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n13858) );
  NAND2_X1 U12686 ( .A1(n13845), .A2(n13858), .ZN(n13844) );
  NAND2_X1 U12687 ( .A1(n13846), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10155) );
  NAND2_X1 U12688 ( .A1(n13844), .A2(n10155), .ZN(n13864) );
  MUX2_X1 U12689 ( .A(n10156), .B(P1_REG2_REG_2__SCAN_IN), .S(n13868), .Z(
        n13865) );
  NAND2_X1 U12690 ( .A1(n13864), .A2(n13865), .ZN(n13882) );
  NAND2_X1 U12691 ( .A1(n10157), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n13881) );
  NAND2_X1 U12692 ( .A1(n13882), .A2(n13881), .ZN(n10159) );
  MUX2_X1 U12693 ( .A(n14674), .B(P1_REG2_REG_3__SCAN_IN), .S(n13879), .Z(
        n10158) );
  NAND2_X1 U12694 ( .A1(n10159), .A2(n10158), .ZN(n14569) );
  OR2_X1 U12695 ( .A1(n13879), .A2(n14674), .ZN(n14568) );
  INV_X1 U12696 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n14664) );
  MUX2_X1 U12697 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n14664), .S(n14575), .Z(
        n14570) );
  AOI21_X1 U12698 ( .B1(n14569), .B2(n14568), .A(n14570), .ZN(n14567) );
  NOR2_X1 U12699 ( .A1(n14575), .A2(n14664), .ZN(n10190) );
  INV_X1 U12700 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n11178) );
  MUX2_X1 U12701 ( .A(n11178), .B(P1_REG2_REG_5__SCAN_IN), .S(n10198), .Z(
        n10189) );
  OAI21_X1 U12702 ( .B1(n14567), .B2(n10190), .A(n10189), .ZN(n10237) );
  INV_X1 U12703 ( .A(n10198), .ZN(n10160) );
  NAND2_X1 U12704 ( .A1(n10160), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10236) );
  MUX2_X1 U12705 ( .A(n11144), .B(P1_REG2_REG_6__SCAN_IN), .S(n10161), .Z(
        n10235) );
  AOI21_X1 U12706 ( .B1(n10237), .B2(n10236), .A(n10235), .ZN(n13898) );
  NOR2_X1 U12707 ( .A1(n10242), .A2(n11144), .ZN(n13897) );
  MUX2_X1 U12708 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10162), .S(n13890), .Z(
        n13896) );
  OAI21_X1 U12709 ( .B1(n13898), .B2(n13897), .A(n13896), .ZN(n13900) );
  NAND2_X1 U12710 ( .A1(n13890), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10164) );
  MUX2_X1 U12711 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n11101), .S(n10178), .Z(
        n10163) );
  AOI21_X1 U12712 ( .B1(n13900), .B2(n10164), .A(n10163), .ZN(n10181) );
  INV_X1 U12713 ( .A(n10181), .ZN(n10166) );
  NAND3_X1 U12714 ( .A1(n13900), .A2(n10164), .A3(n10163), .ZN(n10165) );
  NAND3_X1 U12715 ( .A1(n14606), .A2(n10166), .A3(n10165), .ZN(n10167) );
  OAI211_X1 U12716 ( .C1(n10169), .C2(n11090), .A(n10168), .B(n10167), .ZN(
        P1_U3251) );
  NAND2_X1 U12717 ( .A1(n10178), .A2(n10127), .ZN(n10172) );
  NAND2_X1 U12718 ( .A1(n10174), .A2(n10172), .ZN(n10170) );
  MUX2_X1 U12719 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n7755), .S(n10384), .Z(
        n10171) );
  NAND2_X1 U12720 ( .A1(n10170), .A2(n10171), .ZN(n10386) );
  INV_X1 U12721 ( .A(n10171), .ZN(n10173) );
  NAND3_X1 U12722 ( .A1(n10174), .A2(n10173), .A3(n10172), .ZN(n10175) );
  AND2_X1 U12723 ( .A1(n10386), .A2(n10175), .ZN(n10185) );
  NOR2_X1 U12724 ( .A1(n10176), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11682) );
  INV_X1 U12725 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14240) );
  NOR2_X1 U12726 ( .A1(n14615), .A2(n14240), .ZN(n10177) );
  AOI211_X1 U12727 ( .C1(n14591), .C2(n10384), .A(n11682), .B(n10177), .ZN(
        n10184) );
  NOR2_X1 U12728 ( .A1(n10178), .A2(n11101), .ZN(n10180) );
  MUX2_X1 U12729 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n11430), .S(n10384), .Z(
        n10179) );
  OAI21_X1 U12730 ( .B1(n10181), .B2(n10180), .A(n10179), .ZN(n10381) );
  OR3_X1 U12731 ( .A1(n10181), .A2(n10180), .A3(n10179), .ZN(n10182) );
  NAND3_X1 U12732 ( .A1(n10381), .A2(n14606), .A3(n10182), .ZN(n10183) );
  OAI211_X1 U12733 ( .C1(n10185), .C2(n11090), .A(n10184), .B(n10183), .ZN(
        P1_U3252) );
  OAI21_X1 U12734 ( .B1(n10188), .B2(n10187), .A(n10186), .ZN(n10194) );
  INV_X1 U12735 ( .A(n10237), .ZN(n10192) );
  NOR3_X1 U12736 ( .A1(n14567), .A2(n10190), .A3(n10189), .ZN(n10191) );
  NOR3_X1 U12737 ( .A1(n13920), .A2(n10192), .A3(n10191), .ZN(n10193) );
  AOI21_X1 U12738 ( .B1(n14603), .B2(n10194), .A(n10193), .ZN(n10197) );
  NAND2_X1 U12739 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n13727) );
  INV_X1 U12740 ( .A(n13727), .ZN(n10195) );
  AOI21_X1 U12741 ( .B1(n14587), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10195), .ZN(
        n10196) );
  OAI211_X1 U12742 ( .C1(n10198), .C2(n14611), .A(n10197), .B(n10196), .ZN(
        P1_U3248) );
  NAND2_X1 U12743 ( .A1(n10206), .A2(n10204), .ZN(n10199) );
  NAND2_X1 U12744 ( .A1(n10199), .A2(n10255), .ZN(n10203) );
  INV_X1 U12745 ( .A(n10354), .ZN(n10201) );
  AND2_X1 U12746 ( .A1(n10201), .A2(n10200), .ZN(n10202) );
  NAND2_X1 U12747 ( .A1(n10203), .A2(n10202), .ZN(n10494) );
  NOR2_X1 U12748 ( .A1(n10494), .A2(P2_U3088), .ZN(n10404) );
  NAND2_X1 U12749 ( .A1(n14927), .A2(n10204), .ZN(n14922) );
  INV_X1 U12750 ( .A(n14922), .ZN(n10205) );
  AND2_X1 U12751 ( .A1(n10206), .A2(n10205), .ZN(n10222) );
  NAND2_X1 U12752 ( .A1(n10222), .A2(n14907), .ZN(n10207) );
  INV_X1 U12753 ( .A(n10208), .ZN(n10209) );
  INV_X1 U12754 ( .A(n9477), .ZN(n10210) );
  OAI22_X1 U12755 ( .A1(n10210), .A2(n14420), .B1(n10509), .B2(n14422), .ZN(
        n10265) );
  AOI22_X1 U12756 ( .A1(n14787), .A2(n10267), .B1(n14430), .B2(n10265), .ZN(
        n10225) );
  OR2_X4 U12757 ( .A1(n10212), .A2(n10211), .ZN(n13098) );
  NAND2_X1 U12758 ( .A1(n13270), .A2(n10403), .ZN(n10248) );
  XNOR2_X1 U12759 ( .A(n10247), .B(n10248), .ZN(n10246) );
  NAND2_X1 U12760 ( .A1(n9477), .A2(n10403), .ZN(n10213) );
  NAND2_X1 U12761 ( .A1(n10213), .A2(n10408), .ZN(n10402) );
  NAND2_X1 U12762 ( .A1(n13098), .A2(n10214), .ZN(n10215) );
  NAND2_X1 U12763 ( .A1(n10402), .A2(n10215), .ZN(n10245) );
  XNOR2_X1 U12764 ( .A(n10246), .B(n10245), .ZN(n10223) );
  NAND2_X1 U12765 ( .A1(n10373), .A2(n10216), .ZN(n10217) );
  INV_X1 U12766 ( .A(n10219), .ZN(n10220) );
  NOR2_X1 U12767 ( .A1(n14945), .A2(n10220), .ZN(n10221) );
  NAND2_X1 U12768 ( .A1(n10223), .A2(n14428), .ZN(n10224) );
  OAI211_X1 U12769 ( .C1(n10404), .C2(n10943), .A(n10225), .B(n10224), .ZN(
        P2_U3194) );
  INV_X1 U12770 ( .A(n10226), .ZN(n10229) );
  INV_X1 U12771 ( .A(n10445), .ZN(n10539) );
  OAI222_X1 U12772 ( .A1(n12044), .A2(n10227), .B1(n14208), .B2(n10229), .C1(
        P1_U3086), .C2(n10539), .ZN(P1_U3344) );
  INV_X1 U12773 ( .A(n14834), .ZN(n10230) );
  OAI222_X1 U12774 ( .A1(n10230), .A2(P2_U3088), .B1(n13643), .B2(n10229), 
        .C1(n10228), .C2(n13652), .ZN(P2_U3316) );
  NAND2_X1 U12775 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n11483) );
  OAI211_X1 U12776 ( .C1(n10232), .C2(n10231), .A(n14603), .B(n13893), .ZN(
        n10233) );
  NAND2_X1 U12777 ( .A1(n11483), .A2(n10233), .ZN(n10234) );
  AOI21_X1 U12778 ( .B1(n14587), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n10234), .ZN(
        n10241) );
  INV_X1 U12779 ( .A(n13898), .ZN(n10239) );
  NAND3_X1 U12780 ( .A1(n10237), .A2(n10236), .A3(n10235), .ZN(n10238) );
  NAND3_X1 U12781 ( .A1(n14606), .A2(n10239), .A3(n10238), .ZN(n10240) );
  OAI211_X1 U12782 ( .C1(n14611), .C2(n10242), .A(n10241), .B(n10240), .ZN(
        P1_U3249) );
  OAI22_X1 U12783 ( .A1(n10244), .A2(n14420), .B1(n10243), .B2(n14422), .ZN(
        n10365) );
  AOI22_X1 U12784 ( .A1(n14787), .A2(n6653), .B1(n14430), .B2(n10365), .ZN(
        n10254) );
  NAND2_X1 U12785 ( .A1(n10246), .A2(n10245), .ZN(n10251) );
  INV_X1 U12786 ( .A(n10247), .ZN(n10249) );
  NAND2_X1 U12787 ( .A1(n10249), .A2(n10248), .ZN(n10250) );
  NAND2_X1 U12788 ( .A1(n10251), .A2(n10250), .ZN(n10478) );
  XNOR2_X1 U12789 ( .A(n6653), .B(n13098), .ZN(n10479) );
  NAND2_X1 U12790 ( .A1(n13268), .A2(n13105), .ZN(n10480) );
  XNOR2_X1 U12791 ( .A(n10479), .B(n10480), .ZN(n10477) );
  XNOR2_X1 U12792 ( .A(n10478), .B(n10477), .ZN(n10252) );
  NAND2_X1 U12793 ( .A1(n10252), .A2(n14428), .ZN(n10253) );
  OAI211_X1 U12794 ( .C1(n10404), .C2(n10979), .A(n10254), .B(n10253), .ZN(
        P2_U3209) );
  AND2_X1 U12795 ( .A1(n14926), .A2(n10255), .ZN(n10256) );
  INV_X1 U12796 ( .A(n10259), .ZN(n10262) );
  INV_X1 U12797 ( .A(n10260), .ZN(n10261) );
  AOI21_X1 U12798 ( .B1(n10262), .B2(n10264), .A(n10261), .ZN(n10951) );
  OAI21_X1 U12799 ( .B1(n9476), .B2(n10264), .A(n10263), .ZN(n10266) );
  AOI21_X1 U12800 ( .B1(n10266), .B2(n14886), .A(n10265), .ZN(n10948) );
  AOI211_X1 U12801 ( .C1(n10408), .C2(n10267), .A(n13105), .B(n10360), .ZN(
        n10946) );
  AOI21_X1 U12802 ( .B1(n10267), .B2(n14945), .A(n10946), .ZN(n10268) );
  OAI211_X1 U12803 ( .C1(n10951), .C2(n13614), .A(n10948), .B(n10268), .ZN(
        n10376) );
  INV_X2 U12804 ( .A(n14962), .ZN(n14964) );
  NAND2_X1 U12805 ( .A1(n10376), .A2(n14964), .ZN(n10269) );
  OAI21_X1 U12806 ( .B1(n14964), .B2(n9007), .A(n10269), .ZN(P2_U3433) );
  NAND2_X1 U12807 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n10715) );
  NAND2_X1 U12808 ( .A1(n10289), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10327) );
  NAND2_X1 U12809 ( .A1(n10328), .A2(n10327), .ZN(n10271) );
  MUX2_X1 U12810 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n10515), .S(n10333), .Z(
        n10270) );
  NAND2_X1 U12811 ( .A1(n10271), .A2(n10270), .ZN(n10330) );
  NAND2_X1 U12812 ( .A1(n10333), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10272) );
  NAND2_X1 U12813 ( .A1(n10330), .A2(n10272), .ZN(n14801) );
  MUX2_X1 U12814 ( .A(n10273), .B(P2_REG1_REG_4__SCAN_IN), .S(n14796), .Z(
        n14800) );
  NAND2_X1 U12815 ( .A1(n14801), .A2(n14800), .ZN(n14799) );
  NAND2_X1 U12816 ( .A1(n10294), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10343) );
  NAND2_X1 U12817 ( .A1(n14799), .A2(n10343), .ZN(n10276) );
  MUX2_X1 U12818 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n10274), .S(n10347), .Z(
        n10275) );
  NAND2_X1 U12819 ( .A1(n10276), .A2(n10275), .ZN(n13281) );
  NAND2_X1 U12820 ( .A1(n10347), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n13280) );
  NAND2_X1 U12821 ( .A1(n13281), .A2(n13280), .ZN(n10279) );
  INV_X1 U12822 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10277) );
  MUX2_X1 U12823 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10277), .S(n13278), .Z(
        n10278) );
  NAND2_X1 U12824 ( .A1(n10279), .A2(n10278), .ZN(n13296) );
  NAND2_X1 U12825 ( .A1(n13278), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n13295) );
  NAND2_X1 U12826 ( .A1(n13296), .A2(n13295), .ZN(n10282) );
  INV_X1 U12827 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10280) );
  MUX2_X1 U12828 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10280), .S(n13293), .Z(
        n10281) );
  NAND2_X1 U12829 ( .A1(n10282), .A2(n10281), .ZN(n13298) );
  NAND2_X1 U12830 ( .A1(n13293), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10283) );
  NAND2_X1 U12831 ( .A1(n13298), .A2(n10283), .ZN(n10286) );
  MUX2_X1 U12832 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n10284), .S(n10415), .Z(
        n10285) );
  NAND2_X1 U12833 ( .A1(n10286), .A2(n10285), .ZN(n10411) );
  OAI211_X1 U12834 ( .C1(n10286), .C2(n10285), .A(n14878), .B(n10411), .ZN(
        n10287) );
  NAND2_X1 U12835 ( .A1(n10715), .A2(n10287), .ZN(n10288) );
  AOI21_X1 U12836 ( .B1(n14871), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n10288), .ZN(
        n10308) );
  NAND2_X1 U12837 ( .A1(n10289), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n10335) );
  NAND2_X1 U12838 ( .A1(n10336), .A2(n10335), .ZN(n10292) );
  MUX2_X1 U12839 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10290), .S(n10333), .Z(
        n10291) );
  NAND2_X1 U12840 ( .A1(n10292), .A2(n10291), .ZN(n10338) );
  NAND2_X1 U12841 ( .A1(n10333), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10293) );
  NAND2_X1 U12842 ( .A1(n10338), .A2(n10293), .ZN(n14804) );
  MUX2_X1 U12843 ( .A(n10953), .B(P2_REG2_REG_4__SCAN_IN), .S(n14796), .Z(
        n14803) );
  NAND2_X1 U12844 ( .A1(n14804), .A2(n14803), .ZN(n14802) );
  NAND2_X1 U12845 ( .A1(n10294), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10349) );
  NAND2_X1 U12846 ( .A1(n14802), .A2(n10349), .ZN(n10296) );
  MUX2_X1 U12847 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11168), .S(n10347), .Z(
        n10295) );
  NAND2_X1 U12848 ( .A1(n10296), .A2(n10295), .ZN(n13276) );
  NAND2_X1 U12849 ( .A1(n10347), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n13275) );
  NAND2_X1 U12850 ( .A1(n13276), .A2(n13275), .ZN(n10299) );
  MUX2_X1 U12851 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10297), .S(n13278), .Z(
        n10298) );
  NAND2_X1 U12852 ( .A1(n10299), .A2(n10298), .ZN(n13290) );
  NAND2_X1 U12853 ( .A1(n13278), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n13289) );
  NAND2_X1 U12854 ( .A1(n13290), .A2(n13289), .ZN(n10301) );
  MUX2_X1 U12855 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n11227), .S(n13293), .Z(
        n10300) );
  NAND2_X1 U12856 ( .A1(n10301), .A2(n10300), .ZN(n13292) );
  NAND2_X1 U12857 ( .A1(n13293), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10305) );
  NAND2_X1 U12858 ( .A1(n13292), .A2(n10305), .ZN(n10303) );
  MUX2_X1 U12859 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10996), .S(n10415), .Z(
        n10302) );
  NAND2_X1 U12860 ( .A1(n10303), .A2(n10302), .ZN(n10417) );
  MUX2_X1 U12861 ( .A(n10996), .B(P2_REG2_REG_8__SCAN_IN), .S(n10415), .Z(
        n10304) );
  NAND3_X1 U12862 ( .A1(n13292), .A2(n10305), .A3(n10304), .ZN(n10306) );
  NAND3_X1 U12863 ( .A1(n14875), .A2(n10417), .A3(n10306), .ZN(n10307) );
  OAI211_X1 U12864 ( .C1(n14822), .C2(n10309), .A(n10308), .B(n10307), .ZN(
        P2_U3222) );
  OAI222_X1 U12865 ( .A1(n13076), .A2(n10310), .B1(n13078), .B2(n15224), .C1(
        n12750), .C2(P3_U3151), .ZN(P3_U3280) );
  INV_X1 U12866 ( .A(n14875), .ZN(n14856) );
  NOR2_X1 U12867 ( .A1(n14856), .A2(n10591), .ZN(n14790) );
  AOI22_X1 U12868 ( .A1(n14790), .A2(P2_IR_REG_0__SCAN_IN), .B1(n14875), .B2(
        n10311), .ZN(n10324) );
  INV_X1 U12869 ( .A(n10312), .ZN(n10323) );
  INV_X1 U12870 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10313) );
  OAI22_X1 U12871 ( .A1(n14832), .A2(n10313), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10943), .ZN(n10320) );
  MUX2_X1 U12872 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n10378), .S(n10314), .Z(
        n10315) );
  OAI21_X1 U12873 ( .B1(n9016), .B2(n10316), .A(n10315), .ZN(n10317) );
  AND3_X1 U12874 ( .A1(n14878), .A2(n10318), .A3(n10317), .ZN(n10319) );
  AOI211_X1 U12875 ( .C1(n14873), .C2(n10321), .A(n10320), .B(n10319), .ZN(
        n10322) );
  OAI21_X1 U12876 ( .B1(n10324), .B2(n10323), .A(n10322), .ZN(P2_U3215) );
  INV_X1 U12877 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10325) );
  NOR2_X1 U12878 ( .A1(n14832), .A2(n10325), .ZN(n10332) );
  INV_X1 U12879 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10515) );
  MUX2_X1 U12880 ( .A(n10515), .B(P2_REG1_REG_3__SCAN_IN), .S(n10333), .Z(
        n10326) );
  NAND3_X1 U12881 ( .A1(n10328), .A2(n10327), .A3(n10326), .ZN(n10329) );
  AND3_X1 U12882 ( .A1(n14878), .A2(n10330), .A3(n10329), .ZN(n10331) );
  AOI211_X1 U12883 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(P2_U3088), .A(n10332), 
        .B(n10331), .ZN(n10340) );
  MUX2_X1 U12884 ( .A(n10290), .B(P2_REG2_REG_3__SCAN_IN), .S(n10333), .Z(
        n10334) );
  NAND3_X1 U12885 ( .A1(n10336), .A2(n10335), .A3(n10334), .ZN(n10337) );
  NAND3_X1 U12886 ( .A1(n14875), .A2(n10338), .A3(n10337), .ZN(n10339) );
  OAI211_X1 U12887 ( .C1(n14822), .C2(n10341), .A(n10340), .B(n10339), .ZN(
        P2_U3217) );
  NAND2_X1 U12888 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n12030) );
  INV_X1 U12889 ( .A(n12030), .ZN(n10346) );
  MUX2_X1 U12890 ( .A(n10274), .B(P2_REG1_REG_5__SCAN_IN), .S(n10347), .Z(
        n10342) );
  NAND3_X1 U12891 ( .A1(n14799), .A2(n10343), .A3(n10342), .ZN(n10344) );
  AND3_X1 U12892 ( .A1(n14878), .A2(n13281), .A3(n10344), .ZN(n10345) );
  AOI211_X1 U12893 ( .C1(n14871), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n10346), .B(
        n10345), .ZN(n10352) );
  MUX2_X1 U12894 ( .A(n11168), .B(P2_REG2_REG_5__SCAN_IN), .S(n10347), .Z(
        n10348) );
  NAND3_X1 U12895 ( .A1(n14802), .A2(n10349), .A3(n10348), .ZN(n10350) );
  NAND3_X1 U12896 ( .A1(n14875), .A2(n13276), .A3(n10350), .ZN(n10351) );
  OAI211_X1 U12897 ( .C1(n14822), .C2(n10353), .A(n10352), .B(n10351), .ZN(
        P2_U3219) );
  NOR2_X1 U12898 ( .A1(n14922), .A2(n10354), .ZN(n10355) );
  INV_X2 U12899 ( .A(n14969), .ZN(n13616) );
  OAI21_X1 U12900 ( .B1(n10359), .B2(n10358), .A(n10357), .ZN(n10984) );
  INV_X1 U12901 ( .A(n10984), .ZN(n10368) );
  INV_X1 U12902 ( .A(n10360), .ZN(n10362) );
  INV_X1 U12903 ( .A(n10506), .ZN(n10361) );
  AOI211_X1 U12904 ( .C1(n6653), .C2(n10362), .A(n13489), .B(n10361), .ZN(
        n10983) );
  AOI21_X1 U12905 ( .B1(n6653), .B2(n14945), .A(n10983), .ZN(n10367) );
  XNOR2_X1 U12906 ( .A(n10364), .B(n10363), .ZN(n10366) );
  AOI21_X1 U12907 ( .B1(n10366), .B2(n14886), .A(n10365), .ZN(n10987) );
  OAI211_X1 U12908 ( .C1(n13614), .C2(n10368), .A(n10367), .B(n10987), .ZN(
        n10396) );
  NAND2_X1 U12909 ( .A1(n10396), .A2(n13616), .ZN(n10369) );
  OAI21_X1 U12910 ( .B1(n13616), .B2(n10370), .A(n10369), .ZN(P2_U3501) );
  NOR2_X1 U12911 ( .A1(n9471), .A2(n14886), .ZN(n10371) );
  OR2_X1 U12912 ( .A1(n10595), .A2(n10371), .ZN(n10372) );
  INV_X1 U12913 ( .A(n14422), .ZN(n13233) );
  NAND2_X1 U12914 ( .A1(n13270), .A2(n13233), .ZN(n10401) );
  AND2_X1 U12915 ( .A1(n10372), .A2(n10401), .ZN(n10588) );
  NAND2_X1 U12916 ( .A1(n10408), .A2(n10373), .ZN(n10589) );
  OAI211_X1 U12917 ( .C1(n10595), .C2(n10374), .A(n10588), .B(n10589), .ZN(
        n10393) );
  NAND2_X1 U12918 ( .A1(n10393), .A2(n13616), .ZN(n10375) );
  OAI21_X1 U12919 ( .B1(n13616), .B2(n9016), .A(n10375), .ZN(P2_U3499) );
  NAND2_X1 U12920 ( .A1(n10376), .A2(n13616), .ZN(n10377) );
  OAI21_X1 U12921 ( .B1(n13616), .B2(n10378), .A(n10377), .ZN(P2_U3500) );
  NAND2_X1 U12922 ( .A1(n10384), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10380) );
  MUX2_X1 U12923 ( .A(n10441), .B(P1_REG2_REG_10__SCAN_IN), .S(n10432), .Z(
        n10379) );
  AOI21_X1 U12924 ( .B1(n10381), .B2(n10380), .A(n10379), .ZN(n10449) );
  NAND3_X1 U12925 ( .A1(n10381), .A2(n10380), .A3(n10379), .ZN(n10382) );
  NAND2_X1 U12926 ( .A1(n10382), .A2(n14606), .ZN(n10392) );
  AND2_X1 U12927 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11755) );
  NOR2_X1 U12928 ( .A1(n14611), .A2(n10442), .ZN(n10383) );
  AOI211_X1 U12929 ( .C1(n14587), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n11755), 
        .B(n10383), .ZN(n10391) );
  OR2_X1 U12930 ( .A1(n10384), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n10385) );
  NAND2_X1 U12931 ( .A1(n10386), .A2(n10385), .ZN(n10388) );
  INV_X1 U12932 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n14774) );
  MUX2_X1 U12933 ( .A(n14774), .B(P1_REG1_REG_10__SCAN_IN), .S(n10432), .Z(
        n10387) );
  AOI21_X1 U12934 ( .B1(n10388), .B2(n10387), .A(n11090), .ZN(n10389) );
  NAND2_X1 U12935 ( .A1(n10389), .A2(n10434), .ZN(n10390) );
  OAI211_X1 U12936 ( .C1(n10449), .C2(n10392), .A(n10391), .B(n10390), .ZN(
        P1_U3253) );
  INV_X1 U12937 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10395) );
  NAND2_X1 U12938 ( .A1(n10393), .A2(n14964), .ZN(n10394) );
  OAI21_X1 U12939 ( .B1(n14964), .B2(n10395), .A(n10394), .ZN(P2_U3430) );
  INV_X1 U12940 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10398) );
  NAND2_X1 U12941 ( .A1(n10396), .A2(n14964), .ZN(n10397) );
  OAI21_X1 U12942 ( .B1(n14964), .B2(n10398), .A(n10397), .ZN(P2_U3436) );
  INV_X1 U12943 ( .A(n10399), .ZN(n10431) );
  AOI22_X1 U12944 ( .A1(n10650), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n14202), .ZN(n10400) );
  OAI21_X1 U12945 ( .B1(n10431), .B2(n14208), .A(n10400), .ZN(P1_U3343) );
  INV_X1 U12946 ( .A(n14430), .ZN(n14779) );
  OAI22_X1 U12947 ( .A1(n14782), .A2(n10402), .B1(n14779), .B2(n10401), .ZN(
        n10407) );
  INV_X1 U12948 ( .A(n13225), .ZN(n13201) );
  OAI22_X1 U12949 ( .A1(n13201), .A2(n10405), .B1(n10404), .B2(n10590), .ZN(
        n10406) );
  AOI211_X1 U12950 ( .C1(n10408), .C2(n14787), .A(n10407), .B(n10406), .ZN(
        n10409) );
  INV_X1 U12951 ( .A(n10409), .ZN(P2_U3204) );
  NAND2_X1 U12952 ( .A1(n10415), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10410) );
  NAND2_X1 U12953 ( .A1(n10411), .A2(n10410), .ZN(n14810) );
  MUX2_X1 U12954 ( .A(n10412), .B(P2_REG1_REG_9__SCAN_IN), .S(n10418), .Z(
        n14809) );
  OAI21_X1 U12955 ( .B1(n10418), .B2(P2_REG1_REG_9__SCAN_IN), .A(n14812), .ZN(
        n10414) );
  INV_X1 U12956 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n11057) );
  MUX2_X1 U12957 ( .A(n11057), .B(P2_REG1_REG_10__SCAN_IN), .S(n10795), .Z(
        n10413) );
  NOR2_X1 U12958 ( .A1(n10414), .A2(n10413), .ZN(n10790) );
  AOI211_X1 U12959 ( .C1(n10414), .C2(n10413), .A(n14862), .B(n10790), .ZN(
        n10428) );
  NAND2_X1 U12960 ( .A1(n10415), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10416) );
  NAND2_X1 U12961 ( .A1(n10417), .A2(n10416), .ZN(n14815) );
  MUX2_X1 U12962 ( .A(n11207), .B(P2_REG2_REG_9__SCAN_IN), .S(n10418), .Z(
        n14814) );
  NAND2_X1 U12963 ( .A1(n14821), .A2(n11207), .ZN(n10419) );
  NAND2_X1 U12964 ( .A1(n14817), .A2(n10419), .ZN(n10422) );
  MUX2_X1 U12965 ( .A(n9136), .B(P2_REG2_REG_10__SCAN_IN), .S(n10795), .Z(
        n10421) );
  INV_X1 U12966 ( .A(n10797), .ZN(n10420) );
  AOI211_X1 U12967 ( .C1(n10422), .C2(n10421), .A(n14856), .B(n10420), .ZN(
        n10427) );
  NOR2_X1 U12968 ( .A1(n10423), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10976) );
  AOI21_X1 U12969 ( .B1(n14871), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n10976), 
        .ZN(n10424) );
  OAI21_X1 U12970 ( .B1(n14822), .B2(n10425), .A(n10424), .ZN(n10426) );
  OR3_X1 U12971 ( .A1(n10428), .A2(n10427), .A3(n10426), .ZN(P2_U3224) );
  INV_X1 U12972 ( .A(n14347), .ZN(n12738) );
  OAI222_X1 U12973 ( .A1(n13076), .A2(n10429), .B1(n13078), .B2(n15247), .C1(
        n12738), .C2(P3_U3151), .ZN(P3_U3279) );
  OAI222_X1 U12974 ( .A1(P2_U3088), .A2(n10799), .B1(n13643), .B2(n10431), 
        .C1(n10430), .C2(n13652), .ZN(P2_U3315) );
  MUX2_X1 U12975 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n7805), .S(n10445), .Z(
        n10435) );
  INV_X1 U12976 ( .A(n10435), .ZN(n10439) );
  NAND2_X1 U12977 ( .A1(n10432), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10433) );
  NAND2_X1 U12978 ( .A1(n10434), .A2(n10433), .ZN(n10438) );
  INV_X1 U12979 ( .A(n10438), .ZN(n10436) );
  NAND2_X1 U12980 ( .A1(n10436), .A2(n10435), .ZN(n10543) );
  INV_X1 U12981 ( .A(n10543), .ZN(n10437) );
  AOI21_X1 U12982 ( .B1(n10439), .B2(n10438), .A(n10437), .ZN(n10452) );
  AND2_X1 U12983 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n11864) );
  NOR2_X1 U12984 ( .A1(n14611), .A2(n10539), .ZN(n10440) );
  AOI211_X1 U12985 ( .C1(n14587), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n11864), 
        .B(n10440), .ZN(n10451) );
  INV_X1 U12986 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11654) );
  MUX2_X1 U12987 ( .A(n11654), .B(P1_REG2_REG_11__SCAN_IN), .S(n10445), .Z(
        n10444) );
  NOR2_X1 U12988 ( .A1(n10442), .A2(n10441), .ZN(n10447) );
  INV_X1 U12989 ( .A(n10447), .ZN(n10443) );
  NAND2_X1 U12990 ( .A1(n10444), .A2(n10443), .ZN(n10448) );
  MUX2_X1 U12991 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n11654), .S(n10445), .Z(
        n10446) );
  OAI21_X1 U12992 ( .B1(n10449), .B2(n10447), .A(n10446), .ZN(n10535) );
  OAI211_X1 U12993 ( .C1(n10449), .C2(n10448), .A(n10535), .B(n14606), .ZN(
        n10450) );
  OAI211_X1 U12994 ( .C1(n10452), .C2(n11090), .A(n10451), .B(n10450), .ZN(
        P1_U3254) );
  OR2_X1 U12995 ( .A1(n11010), .A2(n12453), .ZN(n10455) );
  AOI22_X1 U12996 ( .A1(n14694), .A2(n12441), .B1(n10456), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n10454) );
  AND2_X1 U12997 ( .A1(n10455), .A2(n10454), .ZN(n10576) );
  OR2_X4 U12998 ( .A1(n14679), .A2(n12454), .ZN(n12452) );
  OR2_X1 U12999 ( .A1(n11010), .A2(n12452), .ZN(n10458) );
  AOI22_X1 U13000 ( .A1(n10922), .A2(n14694), .B1(n10456), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n10457) );
  OR2_X1 U13001 ( .A1(n14688), .A2(n8333), .ZN(n10459) );
  INV_X1 U13002 ( .A(n11231), .ZN(n10462) );
  OR2_X1 U13003 ( .A1(n10461), .A2(n10460), .ZN(n11230) );
  NAND3_X1 U13004 ( .A1(n10462), .A2(n11254), .A3(n11230), .ZN(n10468) );
  NOR2_X1 U13005 ( .A1(n10468), .A2(n10463), .ZN(n10466) );
  NAND2_X1 U13006 ( .A1(n10466), .A2(n10465), .ZN(n10467) );
  AOI22_X1 U13007 ( .A1(n13810), .A2(n7573), .B1(n13815), .B2(n14694), .ZN(
        n10475) );
  NAND2_X1 U13008 ( .A1(n11235), .A2(n10468), .ZN(n10471) );
  AND2_X1 U13009 ( .A1(n11233), .A2(n10469), .ZN(n10470) );
  NAND2_X1 U13010 ( .A1(n10471), .A2(n10470), .ZN(n10930) );
  INV_X1 U13011 ( .A(n10472), .ZN(n10473) );
  NOR2_X1 U13012 ( .A1(n10930), .A2(n10473), .ZN(n10646) );
  INV_X1 U13013 ( .A(n10646), .ZN(n10583) );
  NAND2_X1 U13014 ( .A1(n10583), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n10474) );
  OAI211_X1 U13015 ( .C1(n13857), .C2(n13817), .A(n10475), .B(n10474), .ZN(
        P1_U3232) );
  INV_X2 U13016 ( .A(n10476), .ZN(n13105) );
  NAND2_X1 U13017 ( .A1(n13266), .A2(n13105), .ZN(n10598) );
  XNOR2_X1 U13018 ( .A(n12032), .B(n10598), .ZN(n10501) );
  NAND3_X1 U13019 ( .A1(n13225), .A2(n13267), .A3(n10484), .ZN(n10500) );
  INV_X1 U13020 ( .A(n10479), .ZN(n10481) );
  NAND2_X1 U13021 ( .A1(n10481), .A2(n10480), .ZN(n10482) );
  AND2_X1 U13022 ( .A1(n13267), .A2(n13489), .ZN(n10483) );
  NAND2_X1 U13023 ( .A1(n10484), .A2(n10483), .ZN(n10487) );
  NAND2_X1 U13024 ( .A1(n10487), .A2(n10485), .ZN(n14783) );
  AND2_X1 U13025 ( .A1(n10501), .A2(n10487), .ZN(n10488) );
  NAND2_X1 U13026 ( .A1(n10489), .A2(n10488), .ZN(n10601) );
  OAI21_X1 U13027 ( .B1(n10501), .B2(n14780), .A(n10490), .ZN(n10491) );
  NAND2_X1 U13028 ( .A1(n10491), .A2(n14428), .ZN(n10499) );
  INV_X1 U13029 ( .A(n10530), .ZN(n10955) );
  NAND2_X1 U13030 ( .A1(n13267), .A2(n13231), .ZN(n10493) );
  NAND2_X1 U13031 ( .A1(n13265), .A2(n13233), .ZN(n10492) );
  NAND2_X1 U13032 ( .A1(n10493), .A2(n10492), .ZN(n10527) );
  AOI22_X1 U13033 ( .A1(n14430), .A2(n10527), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10496) );
  OR2_X1 U13034 ( .A1(n14789), .A2(n10954), .ZN(n10495) );
  OAI211_X1 U13035 ( .C1(n10955), .C2(n13210), .A(n10496), .B(n10495), .ZN(
        n10497) );
  INV_X1 U13036 ( .A(n10497), .ZN(n10498) );
  OAI211_X1 U13037 ( .C1(n10501), .C2(n10500), .A(n10499), .B(n10498), .ZN(
        P2_U3202) );
  OAI21_X1 U13038 ( .B1(n10504), .B2(n10503), .A(n10502), .ZN(n14914) );
  INV_X1 U13039 ( .A(n14914), .ZN(n14911) );
  INV_X1 U13040 ( .A(n10529), .ZN(n10505) );
  AOI211_X1 U13041 ( .C1(n14906), .C2(n10506), .A(n13105), .B(n10505), .ZN(
        n14915) );
  AOI21_X1 U13042 ( .B1(n14906), .B2(n14945), .A(n14915), .ZN(n10511) );
  XNOR2_X1 U13043 ( .A(n10507), .B(n10508), .ZN(n10510) );
  OAI22_X1 U13044 ( .A1(n11165), .A2(n14422), .B1(n10509), .B2(n14420), .ZN(
        n14777) );
  AOI21_X1 U13045 ( .B1(n10510), .B2(n14886), .A(n14777), .ZN(n14909) );
  OAI211_X1 U13046 ( .C1(n13614), .C2(n14911), .A(n10511), .B(n14909), .ZN(
        n10513) );
  NAND2_X1 U13047 ( .A1(n10513), .A2(n14964), .ZN(n10512) );
  OAI21_X1 U13048 ( .B1(n14964), .B2(n9044), .A(n10512), .ZN(P2_U3439) );
  NAND2_X1 U13049 ( .A1(n10513), .A2(n13616), .ZN(n10514) );
  OAI21_X1 U13050 ( .B1(n13616), .B2(n10515), .A(n10514), .ZN(P2_U3502) );
  INV_X1 U13051 ( .A(n10516), .ZN(n10519) );
  INV_X1 U13052 ( .A(n14592), .ZN(n10653) );
  OAI222_X1 U13053 ( .A1(n14208), .A2(n10519), .B1(n10653), .B2(P1_U3086), 
        .C1(n10517), .C2(n12044), .ZN(P1_U3342) );
  INV_X1 U13054 ( .A(n14365), .ZN(n12755) );
  OAI222_X1 U13055 ( .A1(n13076), .A2(n10518), .B1(n13078), .B2(n15327), .C1(
        n12755), .C2(P3_U3151), .ZN(P3_U3278) );
  INV_X1 U13056 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10520) );
  INV_X1 U13057 ( .A(n14866), .ZN(n10800) );
  OAI222_X1 U13058 ( .A1(n13652), .A2(n10520), .B1(n13643), .B2(n10519), .C1(
        P2_U3088), .C2(n10800), .ZN(P2_U3314) );
  INV_X1 U13059 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10533) );
  OAI21_X1 U13060 ( .B1(n10523), .B2(n10522), .A(n10521), .ZN(n10524) );
  INV_X1 U13061 ( .A(n10524), .ZN(n10960) );
  XNOR2_X1 U13062 ( .A(n10526), .B(n10525), .ZN(n10528) );
  AOI21_X1 U13063 ( .B1(n10528), .B2(n14886), .A(n10527), .ZN(n10952) );
  AOI211_X1 U13064 ( .C1(n10530), .C2(n10529), .A(n13105), .B(n11160), .ZN(
        n10957) );
  AOI21_X1 U13065 ( .B1(n10530), .B2(n14945), .A(n10957), .ZN(n10531) );
  OAI211_X1 U13066 ( .C1(n10960), .C2(n13614), .A(n10952), .B(n10531), .ZN(
        n13617) );
  NAND2_X1 U13067 ( .A1(n13617), .A2(n14964), .ZN(n10532) );
  OAI21_X1 U13068 ( .B1(n14964), .B2(n10533), .A(n10532), .ZN(P2_U3442) );
  MUX2_X1 U13069 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n11693), .S(n10650), .Z(
        n10534) );
  INV_X1 U13070 ( .A(n10534), .ZN(n10537) );
  OAI21_X1 U13071 ( .B1(n11654), .B2(n10539), .A(n10535), .ZN(n10536) );
  NOR2_X1 U13072 ( .A1(n10536), .A2(n10537), .ZN(n10656) );
  AOI21_X1 U13073 ( .B1(n10537), .B2(n10536), .A(n10656), .ZN(n10547) );
  INV_X1 U13074 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n14246) );
  NAND2_X1 U13075 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n11905)
         );
  OAI21_X1 U13076 ( .B1(n14615), .B2(n14246), .A(n11905), .ZN(n10538) );
  AOI21_X1 U13077 ( .B1(n10650), .B2(n14591), .A(n10538), .ZN(n10546) );
  NAND2_X1 U13078 ( .A1(n10539), .A2(n7805), .ZN(n10541) );
  MUX2_X1 U13079 ( .A(n10540), .B(P1_REG1_REG_12__SCAN_IN), .S(n10650), .Z(
        n10542) );
  AOI21_X1 U13080 ( .B1(n10543), .B2(n10541), .A(n10542), .ZN(n10651) );
  AND3_X1 U13081 ( .A1(n10543), .A2(n10542), .A3(n10541), .ZN(n10544) );
  OAI21_X1 U13082 ( .B1(n10651), .B2(n10544), .A(n14603), .ZN(n10545) );
  OAI211_X1 U13083 ( .C1(n10547), .C2(n13920), .A(n10546), .B(n10545), .ZN(
        P1_U3255) );
  CLKBUF_X1 U13084 ( .A(n10548), .Z(n10573) );
  INV_X1 U13085 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10549) );
  NOR2_X1 U13086 ( .A1(n10573), .A2(n10549), .ZN(P3_U3235) );
  INV_X1 U13087 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10550) );
  NOR2_X1 U13088 ( .A1(n10573), .A2(n10550), .ZN(P3_U3252) );
  INV_X1 U13089 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10551) );
  NOR2_X1 U13090 ( .A1(n10573), .A2(n10551), .ZN(P3_U3239) );
  INV_X1 U13091 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10552) );
  NOR2_X1 U13092 ( .A1(n10573), .A2(n10552), .ZN(P3_U3246) );
  INV_X1 U13093 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10553) );
  NOR2_X1 U13094 ( .A1(n10573), .A2(n10553), .ZN(P3_U3245) );
  INV_X1 U13095 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10554) );
  NOR2_X1 U13096 ( .A1(n10573), .A2(n10554), .ZN(P3_U3261) );
  INV_X1 U13097 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10555) );
  NOR2_X1 U13098 ( .A1(n10573), .A2(n10555), .ZN(P3_U3260) );
  INV_X1 U13099 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10556) );
  NOR2_X1 U13100 ( .A1(n10573), .A2(n10556), .ZN(P3_U3238) );
  INV_X1 U13101 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10557) );
  NOR2_X1 U13102 ( .A1(n10573), .A2(n10557), .ZN(P3_U3237) );
  INV_X1 U13103 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10558) );
  NOR2_X1 U13104 ( .A1(n10573), .A2(n10558), .ZN(P3_U3236) );
  INV_X1 U13105 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10559) );
  NOR2_X1 U13106 ( .A1(n10573), .A2(n10559), .ZN(P3_U3258) );
  INV_X1 U13107 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10560) );
  NOR2_X1 U13108 ( .A1(n10573), .A2(n10560), .ZN(P3_U3244) );
  INV_X1 U13109 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10561) );
  NOR2_X1 U13110 ( .A1(n10573), .A2(n10561), .ZN(P3_U3243) );
  INV_X1 U13111 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10562) );
  NOR2_X1 U13112 ( .A1(n10573), .A2(n10562), .ZN(P3_U3242) );
  INV_X1 U13113 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10563) );
  NOR2_X1 U13114 ( .A1(n10573), .A2(n10563), .ZN(P3_U3241) );
  INV_X1 U13115 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10564) );
  NOR2_X1 U13116 ( .A1(n10573), .A2(n10564), .ZN(P3_U3240) );
  INV_X1 U13117 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10565) );
  NOR2_X1 U13118 ( .A1(n10573), .A2(n10565), .ZN(P3_U3255) );
  INV_X1 U13119 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10566) );
  NOR2_X1 U13120 ( .A1(n10573), .A2(n10566), .ZN(P3_U3263) );
  INV_X1 U13121 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10567) );
  NOR2_X1 U13122 ( .A1(n10573), .A2(n10567), .ZN(P3_U3262) );
  INV_X1 U13123 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10568) );
  NOR2_X1 U13124 ( .A1(n10573), .A2(n10568), .ZN(P3_U3254) );
  INV_X1 U13125 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10569) );
  NOR2_X1 U13126 ( .A1(n10573), .A2(n10569), .ZN(P3_U3257) );
  INV_X1 U13127 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n10570) );
  NOR2_X1 U13128 ( .A1(n10573), .A2(n10570), .ZN(P3_U3234) );
  INV_X1 U13129 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10571) );
  NOR2_X1 U13130 ( .A1(n10573), .A2(n10571), .ZN(P3_U3253) );
  INV_X1 U13131 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10572) );
  NOR2_X1 U13132 ( .A1(n10573), .A2(n10572), .ZN(P3_U3256) );
  INV_X1 U13133 ( .A(n14380), .ZN(n12748) );
  OAI222_X1 U13134 ( .A1(n13076), .A2(n10574), .B1(n13078), .B2(n15252), .C1(
        n12748), .C2(P3_U3151), .ZN(P3_U3277) );
  AOI21_X1 U13135 ( .B1(n10576), .B2(n12444), .A(n10575), .ZN(n10581) );
  OAI22_X1 U13136 ( .A1(n11150), .A2(n12453), .B1(n14698), .B2(n12454), .ZN(
        n10577) );
  AOI22_X1 U13137 ( .A1(n7573), .A2(n12446), .B1(n10922), .B2(n6493), .ZN(
        n10578) );
  OAI21_X1 U13138 ( .B1(n10579), .B2(n10578), .A(n10638), .ZN(n10580) );
  AOI21_X1 U13139 ( .B1(n10581), .B2(n10580), .A(n10640), .ZN(n10586) );
  INV_X1 U13140 ( .A(n13769), .ZN(n13778) );
  INV_X1 U13141 ( .A(n14482), .ZN(n14053) );
  INV_X1 U13142 ( .A(n13808), .ZN(n10582) );
  AOI22_X1 U13143 ( .A1(n10582), .A2(n13843), .B1(n13815), .B2(n6493), .ZN(
        n10585) );
  NOR2_X1 U13144 ( .A1(n10641), .A2(n14055), .ZN(n11008) );
  AOI22_X1 U13145 ( .A1(n10583), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n11008), 
        .B2(n13769), .ZN(n10584) );
  OAI211_X1 U13146 ( .C1(n10586), .C2(n13817), .A(n10585), .B(n10584), .ZN(
        P1_U3222) );
  NAND2_X1 U13147 ( .A1(n14919), .A2(n10587), .ZN(n14912) );
  OAI21_X1 U13148 ( .B1(n9472), .B2(n10589), .A(n10588), .ZN(n10593) );
  OAI22_X1 U13149 ( .A1(n14919), .A2(n10591), .B1(n10590), .B2(n13518), .ZN(
        n10592) );
  AOI21_X1 U13150 ( .B1(n14919), .B2(n10593), .A(n10592), .ZN(n10594) );
  OAI21_X1 U13151 ( .B1(n10595), .B2(n14912), .A(n10594), .ZN(P2_U3265) );
  INV_X1 U13152 ( .A(n10596), .ZN(n10630) );
  OAI222_X1 U13153 ( .A1(n14208), .A2(n10630), .B1(n11616), .B2(P1_U3086), 
        .C1(n10597), .C2(n12044), .ZN(P1_U3339) );
  INV_X1 U13154 ( .A(n12032), .ZN(n10599) );
  NAND2_X1 U13155 ( .A1(n10599), .A2(n10598), .ZN(n10600) );
  NAND2_X1 U13156 ( .A1(n10601), .A2(n10600), .ZN(n10603) );
  XNOR2_X1 U13157 ( .A(n10602), .B(n6725), .ZN(n10604) );
  NAND2_X1 U13158 ( .A1(n13265), .A2(n13105), .ZN(n10605) );
  XNOR2_X1 U13159 ( .A(n10604), .B(n10605), .ZN(n12033) );
  INV_X1 U13160 ( .A(n10604), .ZN(n10606) );
  NAND2_X1 U13161 ( .A1(n10606), .A2(n10605), .ZN(n10607) );
  XNOR2_X1 U13162 ( .A(n14934), .B(n13098), .ZN(n10608) );
  AND2_X1 U13163 ( .A1(n13264), .A2(n13489), .ZN(n10609) );
  NAND2_X1 U13164 ( .A1(n10608), .A2(n10609), .ZN(n10618) );
  INV_X1 U13165 ( .A(n10608), .ZN(n10617) );
  INV_X1 U13166 ( .A(n10609), .ZN(n10610) );
  XNOR2_X1 U13167 ( .A(n11216), .B(n6725), .ZN(n10707) );
  AND2_X1 U13168 ( .A1(n13263), .A2(n13489), .ZN(n10612) );
  NAND2_X1 U13169 ( .A1(n10707), .A2(n10612), .ZN(n10708) );
  INV_X1 U13170 ( .A(n10707), .ZN(n10614) );
  INV_X1 U13171 ( .A(n10612), .ZN(n10613) );
  NAND2_X1 U13172 ( .A1(n10614), .A2(n10613), .ZN(n10615) );
  INV_X1 U13173 ( .A(n10620), .ZN(n10616) );
  AOI21_X1 U13174 ( .B1(n10700), .B2(n10616), .A(n14782), .ZN(n10623) );
  NOR3_X1 U13175 ( .A1(n13201), .A2(n10617), .A3(n11166), .ZN(n10622) );
  OAI21_X1 U13176 ( .B1(n10623), .B2(n10622), .A(n10711), .ZN(n10629) );
  NAND2_X1 U13177 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n13286) );
  NAND2_X1 U13178 ( .A1(n13264), .A2(n13231), .ZN(n10625) );
  NAND2_X1 U13179 ( .A1(n13262), .A2(n13233), .ZN(n10624) );
  NAND2_X1 U13180 ( .A1(n10625), .A2(n10624), .ZN(n11225) );
  NAND2_X1 U13181 ( .A1(n14430), .A2(n11225), .ZN(n10626) );
  OAI211_X1 U13182 ( .C1(n14789), .C2(n11220), .A(n13286), .B(n10626), .ZN(
        n10627) );
  AOI21_X1 U13183 ( .B1(n11216), .B2(n14787), .A(n10627), .ZN(n10628) );
  NAND2_X1 U13184 ( .A1(n10629), .A2(n10628), .ZN(P2_U3185) );
  INV_X1 U13185 ( .A(n11528), .ZN(n11525) );
  OAI222_X1 U13186 ( .A1(n13652), .A2(n10631), .B1(n13643), .B2(n10630), .C1(
        P2_U3088), .C2(n11525), .ZN(P2_U3311) );
  INV_X1 U13187 ( .A(n10632), .ZN(n10634) );
  INV_X1 U13188 ( .A(n11300), .ZN(n11092) );
  OAI222_X1 U13189 ( .A1(n12044), .A2(n10633), .B1(n14214), .B2(n10634), .C1(
        P1_U3086), .C2(n11092), .ZN(P1_U3340) );
  INV_X1 U13190 ( .A(n14872), .ZN(n11458) );
  OAI222_X1 U13191 ( .A1(n13652), .A2(n10635), .B1(n13643), .B2(n10634), .C1(
        n11458), .C2(P2_U3088), .ZN(P2_U3312) );
  INV_X1 U13192 ( .A(n10636), .ZN(n10689) );
  INV_X1 U13193 ( .A(n11614), .ZN(n13905) );
  OAI222_X1 U13194 ( .A1(n14208), .A2(n10689), .B1(n13905), .B2(P1_U3086), 
        .C1(n10637), .C2(n12044), .ZN(P1_U3338) );
  INV_X1 U13195 ( .A(n10638), .ZN(n10639) );
  OAI22_X1 U13196 ( .A1(n10641), .A2(n12452), .B1(n14705), .B2(n12453), .ZN(
        n10917) );
  XNOR2_X1 U13197 ( .A(n10918), .B(n10917), .ZN(n10642) );
  AOI21_X1 U13198 ( .B1(n6648), .B2(n10642), .A(n10919), .ZN(n10649) );
  OR2_X1 U13199 ( .A1(n11150), .A2(n14053), .ZN(n10644) );
  NAND2_X1 U13200 ( .A1(n13841), .A2(n14631), .ZN(n10643) );
  NAND2_X1 U13201 ( .A1(n10644), .A2(n10643), .ZN(n11115) );
  INV_X1 U13202 ( .A(n13815), .ZN(n13803) );
  OAI22_X1 U13203 ( .A1(n10646), .A2(n10645), .B1(n13803), .B2(n14705), .ZN(
        n10647) );
  AOI21_X1 U13204 ( .B1(n13769), .B2(n11115), .A(n10647), .ZN(n10648) );
  OAI21_X1 U13205 ( .B1(n10649), .B2(n13817), .A(n10648), .ZN(P1_U3237) );
  INV_X1 U13206 ( .A(n10663), .ZN(n11088) );
  AOI22_X1 U13207 ( .A1(n10663), .A2(n7860), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n11088), .ZN(n10655) );
  INV_X1 U13208 ( .A(n10650), .ZN(n10657) );
  AOI21_X1 U13209 ( .B1(n10540), .B2(n10657), .A(n10651), .ZN(n14598) );
  MUX2_X1 U13210 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10652), .S(n14592), .Z(
        n14597) );
  NAND2_X1 U13211 ( .A1(n14598), .A2(n14597), .ZN(n14596) );
  OAI21_X1 U13212 ( .B1(n10653), .B2(n10652), .A(n14596), .ZN(n10654) );
  NOR2_X1 U13213 ( .A1(n10655), .A2(n10654), .ZN(n11087) );
  AOI21_X1 U13214 ( .B1(n10655), .B2(n10654), .A(n11087), .ZN(n10669) );
  NAND2_X1 U13215 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n14592), .ZN(n10659) );
  AOI21_X1 U13216 ( .B1(n11693), .B2(n10657), .A(n10656), .ZN(n14595) );
  MUX2_X1 U13217 ( .A(n11813), .B(P1_REG2_REG_13__SCAN_IN), .S(n14592), .Z(
        n10658) );
  INV_X1 U13218 ( .A(n10658), .ZN(n14594) );
  NAND2_X1 U13219 ( .A1(n14595), .A2(n14594), .ZN(n14593) );
  NAND2_X1 U13220 ( .A1(n10659), .A2(n14593), .ZN(n10661) );
  MUX2_X1 U13221 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n14485), .S(n10663), .Z(
        n10660) );
  NAND2_X1 U13222 ( .A1(n10660), .A2(n10661), .ZN(n11085) );
  OAI211_X1 U13223 ( .C1(n10661), .C2(n10660), .A(n14606), .B(n11085), .ZN(
        n10662) );
  INV_X1 U13224 ( .A(n10662), .ZN(n10667) );
  INV_X1 U13225 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10665) );
  NAND2_X1 U13226 ( .A1(n14591), .A2(n10663), .ZN(n10664) );
  NAND2_X1 U13227 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n12002)
         );
  OAI211_X1 U13228 ( .C1(n10665), .C2(n14615), .A(n10664), .B(n12002), .ZN(
        n10666) );
  NOR2_X1 U13229 ( .A1(n10667), .A2(n10666), .ZN(n10668) );
  OAI21_X1 U13230 ( .B1(n10669), .B2(n11090), .A(n10668), .ZN(P1_U3257) );
  INV_X1 U13231 ( .A(n15105), .ZN(n12176) );
  NOR3_X1 U13232 ( .A1(n12176), .A2(n10670), .A3(n15102), .ZN(n10672) );
  AOI211_X1 U13233 ( .C1(n10674), .C2(n10673), .A(n10672), .B(n10671), .ZN(
        n10680) );
  NOR2_X2 U13234 ( .A1(n11837), .A2(n12927), .ZN(n12552) );
  OAI22_X1 U13235 ( .A1(n12608), .A2(n10884), .B1(n10676), .B2(n12649), .ZN(
        n10677) );
  AOI21_X1 U13236 ( .B1(n12552), .B2(n8497), .A(n10677), .ZN(n10679) );
  NAND2_X1 U13237 ( .A1(n12645), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10787) );
  NAND2_X1 U13238 ( .A1(n10787), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n10678) );
  OAI211_X1 U13239 ( .C1(n10680), .C2(n12637), .A(n10679), .B(n10678), .ZN(
        P3_U3162) );
  NAND2_X1 U13240 ( .A1(n10787), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10683) );
  NAND2_X1 U13241 ( .A1(n8497), .A2(n10681), .ZN(n12213) );
  NAND2_X1 U13242 ( .A1(n12212), .A2(n12213), .ZN(n10690) );
  AOI22_X1 U13243 ( .A1(n12642), .A2(n10690), .B1(n12634), .B2(n8873), .ZN(
        n10682) );
  OAI211_X1 U13244 ( .C1(n10785), .C2(n12608), .A(n10683), .B(n10682), .ZN(
        P3_U3172) );
  INV_X1 U13245 ( .A(n10684), .ZN(n10696) );
  OAI222_X1 U13246 ( .A1(n14208), .A2(n10696), .B1(n11088), .B2(P1_U3086), 
        .C1(n10685), .C2(n12044), .ZN(P1_U3341) );
  OAI222_X1 U13247 ( .A1(P3_U3151), .A2(n8454), .B1(n13078), .B2(n10687), .C1(
        n13076), .C2(n10686), .ZN(P3_U3276) );
  INV_X1 U13248 ( .A(n11624), .ZN(n11632) );
  OAI222_X1 U13249 ( .A1(P2_U3088), .A2(n11632), .B1(n13643), .B2(n10689), 
        .C1(n10688), .C2(n13652), .ZN(P2_U3310) );
  INV_X1 U13250 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10693) );
  INV_X1 U13251 ( .A(n10690), .ZN(n12173) );
  NOR3_X1 U13252 ( .A1(n12173), .A2(n15150), .A3(n10691), .ZN(n10692) );
  AOI21_X1 U13253 ( .B1(n15104), .B2(n9764), .A(n10692), .ZN(n11083) );
  MUX2_X1 U13254 ( .A(n10693), .B(n11083), .S(n15175), .Z(n10694) );
  OAI21_X1 U13255 ( .B1(n10681), .B2(n13059), .A(n10694), .ZN(P3_U3390) );
  INV_X1 U13256 ( .A(n11446), .ZN(n11457) );
  OAI222_X1 U13257 ( .A1(P2_U3088), .A2(n11457), .B1(n13643), .B2(n10696), 
        .C1(n10695), .C2(n13652), .ZN(P2_U3313) );
  NAND2_X1 U13258 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n13271) );
  NAND2_X1 U13259 ( .A1(n13265), .A2(n13231), .ZN(n10698) );
  NAND2_X1 U13260 ( .A1(n13263), .A2(n13233), .ZN(n10697) );
  NAND2_X1 U13261 ( .A1(n10698), .A2(n10697), .ZN(n14885) );
  NAND2_X1 U13262 ( .A1(n14430), .A2(n14885), .ZN(n10699) );
  OAI211_X1 U13263 ( .C1(n14789), .C2(n14888), .A(n13271), .B(n10699), .ZN(
        n10705) );
  INV_X1 U13264 ( .A(n10700), .ZN(n10701) );
  AOI211_X1 U13265 ( .C1(n10703), .C2(n10702), .A(n14782), .B(n10701), .ZN(
        n10704) );
  AOI211_X1 U13266 ( .C1(n14934), .C2(n14787), .A(n10705), .B(n10704), .ZN(
        n10706) );
  INV_X1 U13267 ( .A(n10706), .ZN(P2_U3211) );
  NAND2_X1 U13268 ( .A1(n13262), .A2(n13105), .ZN(n10962) );
  NAND3_X1 U13269 ( .A1(n10707), .A2(n13225), .A3(n13263), .ZN(n10720) );
  AND2_X1 U13270 ( .A1(n10721), .A2(n10708), .ZN(n10709) );
  OAI21_X1 U13271 ( .B1(n10721), .B2(n10711), .A(n12397), .ZN(n10712) );
  NAND2_X1 U13272 ( .A1(n10712), .A2(n14428), .ZN(n10719) );
  NOR2_X1 U13273 ( .A1(n14789), .A2(n10998), .ZN(n10717) );
  NAND2_X1 U13274 ( .A1(n13263), .A2(n13231), .ZN(n10714) );
  NAND2_X1 U13275 ( .A1(n13261), .A2(n13233), .ZN(n10713) );
  AND2_X1 U13276 ( .A1(n10714), .A2(n10713), .ZN(n10993) );
  OAI21_X1 U13277 ( .B1(n14779), .B2(n10993), .A(n10715), .ZN(n10716) );
  AOI211_X1 U13278 ( .C1(n14946), .C2(n14787), .A(n10717), .B(n10716), .ZN(
        n10718) );
  OAI211_X1 U13279 ( .C1(n10721), .C2(n10720), .A(n10719), .B(n10718), .ZN(
        P2_U3193) );
  NOR2_X1 U13280 ( .A1(n10723), .A2(P3_U3151), .ZN(n12377) );
  INV_X1 U13281 ( .A(n12377), .ZN(n12383) );
  NAND2_X1 U13282 ( .A1(n10722), .A2(n12383), .ZN(n10737) );
  NAND2_X1 U13283 ( .A1(n10723), .A2(n12370), .ZN(n10724) );
  AND2_X1 U13284 ( .A1(n8482), .A2(n10724), .ZN(n10735) );
  INV_X1 U13285 ( .A(n10746), .ZN(n10725) );
  MUX2_X1 U13286 ( .A(n12658), .B(n10725), .S(n13079), .Z(n15052) );
  NAND2_X1 U13287 ( .A1(n10727), .A2(n6976), .ZN(n10773) );
  INV_X1 U13288 ( .A(n10727), .ZN(n10728) );
  NAND2_X1 U13289 ( .A1(n10728), .A2(n10753), .ZN(n10729) );
  NAND2_X1 U13290 ( .A1(n10773), .A2(n10729), .ZN(n10732) );
  INV_X1 U13291 ( .A(n10732), .ZN(n10734) );
  NAND2_X1 U13292 ( .A1(n10902), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10911) );
  INV_X1 U13293 ( .A(n10911), .ZN(n10733) );
  OAI21_X1 U13294 ( .B1(n10734), .B2(n10733), .A(n10774), .ZN(n10751) );
  INV_X1 U13295 ( .A(n10735), .ZN(n10736) );
  INV_X1 U13296 ( .A(n15068), .ZN(n15043) );
  INV_X1 U13297 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n14219) );
  OAI22_X1 U13298 ( .A1(n15043), .A2(n14219), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15113), .ZN(n10750) );
  INV_X1 U13299 ( .A(n10738), .ZN(n10739) );
  NOR2_X1 U13300 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n10731), .ZN(n10908) );
  NAND2_X1 U13301 ( .A1(n8478), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10740) );
  AOI21_X1 U13302 ( .B1(n10726), .B2(n10741), .A(n6649), .ZN(n10748) );
  NAND2_X1 U13303 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n6849), .ZN(n10906) );
  INV_X1 U13304 ( .A(n10906), .ZN(n10742) );
  OAI21_X1 U13305 ( .B1(n10753), .B2(n10742), .A(n7495), .ZN(n10744) );
  OR2_X1 U13306 ( .A1(n10744), .A2(n10745), .ZN(n10754) );
  INV_X1 U13307 ( .A(n10754), .ZN(n10743) );
  AOI21_X1 U13308 ( .B1(n10745), .B2(n10744), .A(n10743), .ZN(n10747) );
  OAI22_X1 U13309 ( .A1(n15063), .A2(n10748), .B1(n10747), .B2(n15036), .ZN(
        n10749) );
  AOI211_X1 U13310 ( .C1(n15078), .C2(n10751), .A(n10750), .B(n10749), .ZN(
        n10752) );
  OAI21_X1 U13311 ( .B1(n10753), .B2(n15052), .A(n10752), .ZN(P3_U3183) );
  MUX2_X1 U13312 ( .A(P3_REG1_REG_2__SCAN_IN), .B(n10765), .S(n10834), .Z(
        n10756) );
  NAND2_X1 U13313 ( .A1(n10754), .A2(n7495), .ZN(n10755) );
  NAND2_X1 U13314 ( .A1(n10756), .A2(n10755), .ZN(n10836) );
  OAI21_X1 U13315 ( .B1(n10756), .B2(n10755), .A(n10836), .ZN(n10764) );
  OAI22_X1 U13316 ( .A1(n15043), .A2(n14220), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15226), .ZN(n10763) );
  AND2_X1 U13317 ( .A1(n8478), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10757) );
  INV_X1 U13318 ( .A(n10760), .ZN(n10758) );
  NAND2_X1 U13319 ( .A1(n10760), .A2(n10759), .ZN(n10761) );
  AOI21_X1 U13320 ( .B1(n10819), .B2(n10761), .A(n15063), .ZN(n10762) );
  AOI211_X1 U13321 ( .C1(n15069), .C2(n10764), .A(n10763), .B(n10762), .ZN(
        n10780) );
  INV_X1 U13322 ( .A(n10774), .ZN(n10772) );
  INV_X1 U13323 ( .A(n10773), .ZN(n10771) );
  INV_X1 U13324 ( .A(n10834), .ZN(n10767) );
  NAND2_X1 U13325 ( .A1(n10768), .A2(n10767), .ZN(n14979) );
  INV_X1 U13326 ( .A(n10768), .ZN(n10769) );
  NAND2_X1 U13327 ( .A1(n10769), .A2(n10834), .ZN(n10770) );
  AND2_X1 U13328 ( .A1(n14979), .A2(n10770), .ZN(n10775) );
  NOR3_X1 U13329 ( .A1(n10772), .A2(n10771), .A3(n10775), .ZN(n10778) );
  NAND2_X1 U13330 ( .A1(n10774), .A2(n10773), .ZN(n10776) );
  NAND2_X1 U13331 ( .A1(n10776), .A2(n10775), .ZN(n14980) );
  INV_X1 U13332 ( .A(n14980), .ZN(n10777) );
  OAI21_X1 U13333 ( .B1(n10778), .B2(n10777), .A(n15078), .ZN(n10779) );
  OAI211_X1 U13334 ( .C1(n15052), .C2(n10834), .A(n10780), .B(n10779), .ZN(
        P3_U3184) );
  XOR2_X1 U13335 ( .A(n10782), .B(n10781), .Z(n10789) );
  AOI22_X1 U13336 ( .A1(n10675), .A2(n15091), .B1(n10783), .B2(n12634), .ZN(
        n10784) );
  OAI21_X1 U13337 ( .B1(n10785), .B2(n12632), .A(n10784), .ZN(n10786) );
  AOI21_X1 U13338 ( .B1(n10787), .B2(P3_REG3_REG_2__SCAN_IN), .A(n10786), .ZN(
        n10788) );
  OAI21_X1 U13339 ( .B1(n10789), .B2(n12637), .A(n10788), .ZN(P3_U3177) );
  AOI21_X1 U13340 ( .B1(n10795), .B2(P2_REG1_REG_10__SCAN_IN), .A(n10790), 
        .ZN(n14837) );
  MUX2_X1 U13341 ( .A(n9148), .B(P2_REG1_REG_11__SCAN_IN), .S(n14834), .Z(
        n14836) );
  NOR2_X1 U13342 ( .A1(n14837), .A2(n14836), .ZN(n14835) );
  AOI21_X1 U13343 ( .B1(n14834), .B2(P2_REG1_REG_11__SCAN_IN), .A(n14835), 
        .ZN(n14849) );
  MUX2_X1 U13344 ( .A(n9167), .B(P2_REG1_REG_12__SCAN_IN), .S(n10799), .Z(
        n14848) );
  NAND2_X1 U13345 ( .A1(n14849), .A2(n14848), .ZN(n14847) );
  OAI21_X1 U13346 ( .B1(n14850), .B2(P2_REG1_REG_12__SCAN_IN), .A(n14847), 
        .ZN(n14863) );
  MUX2_X1 U13347 ( .A(n9180), .B(P2_REG1_REG_13__SCAN_IN), .S(n14866), .Z(
        n14864) );
  NOR2_X1 U13348 ( .A1(n14863), .A2(n14864), .ZN(n14861) );
  INV_X1 U13349 ( .A(n14861), .ZN(n10791) );
  NAND2_X1 U13350 ( .A1(n14866), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n10792) );
  INV_X1 U13351 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n14455) );
  MUX2_X1 U13352 ( .A(n14455), .B(P2_REG1_REG_14__SCAN_IN), .S(n11446), .Z(
        n10793) );
  AOI21_X1 U13353 ( .B1(n10791), .B2(n10792), .A(n10793), .ZN(n11455) );
  NAND2_X1 U13354 ( .A1(n10793), .A2(n10792), .ZN(n10794) );
  OAI21_X1 U13355 ( .B1(n14861), .B2(n10794), .A(n14878), .ZN(n10805) );
  NAND2_X1 U13356 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14431)
         );
  NAND2_X1 U13357 ( .A1(n10795), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10796) );
  NAND2_X1 U13358 ( .A1(n10797), .A2(n10796), .ZN(n14829) );
  MUX2_X1 U13359 ( .A(n11276), .B(P2_REG2_REG_11__SCAN_IN), .S(n14834), .Z(
        n14830) );
  OR2_X1 U13360 ( .A1(n14834), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n10798) );
  NAND2_X1 U13361 ( .A1(n14827), .A2(n10798), .ZN(n14843) );
  MUX2_X1 U13362 ( .A(n11318), .B(P2_REG2_REG_12__SCAN_IN), .S(n10799), .Z(
        n14842) );
  AOI21_X1 U13363 ( .B1(n11318), .B2(n10799), .A(n14845), .ZN(n14860) );
  MUX2_X1 U13364 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n11475), .S(n14866), .Z(
        n14859) );
  NAND2_X1 U13365 ( .A1(n14860), .A2(n14859), .ZN(n14858) );
  OAI21_X1 U13366 ( .B1(n11475), .B2(n10800), .A(n14858), .ZN(n11447) );
  XNOR2_X1 U13367 ( .A(n11447), .B(n11457), .ZN(n10801) );
  NAND2_X1 U13368 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n10801), .ZN(n11448) );
  OAI211_X1 U13369 ( .C1(P2_REG2_REG_14__SCAN_IN), .C2(n10801), .A(n14875), 
        .B(n11448), .ZN(n10802) );
  AND2_X1 U13370 ( .A1(n14431), .A2(n10802), .ZN(n10804) );
  AOI22_X1 U13371 ( .A1(n14873), .A2(n11446), .B1(n14871), .B2(
        P2_ADDR_REG_14__SCAN_IN), .ZN(n10803) );
  OAI211_X1 U13372 ( .C1(n11455), .C2(n10805), .A(n10804), .B(n10803), .ZN(
        P2_U3228) );
  XNOR2_X1 U13373 ( .A(n10852), .B(n10858), .ZN(n10854) );
  INV_X1 U13374 ( .A(n15005), .ZN(n10842) );
  INV_X1 U13375 ( .A(n10813), .ZN(n10814) );
  NAND2_X1 U13376 ( .A1(n14980), .A2(n14979), .ZN(n10811) );
  INV_X1 U13377 ( .A(n14976), .ZN(n10837) );
  NAND2_X1 U13378 ( .A1(n10808), .A2(n10837), .ZN(n10812) );
  INV_X1 U13379 ( .A(n10808), .ZN(n10809) );
  NAND2_X1 U13380 ( .A1(n10809), .A2(n14976), .ZN(n10810) );
  AND2_X1 U13381 ( .A1(n10812), .A2(n10810), .ZN(n14977) );
  NAND2_X1 U13382 ( .A1(n10811), .A2(n14977), .ZN(n14982) );
  NAND2_X1 U13383 ( .A1(n14982), .A2(n10812), .ZN(n14991) );
  XNOR2_X1 U13384 ( .A(n10813), .B(n10842), .ZN(n14990) );
  AND2_X1 U13385 ( .A1(n14991), .A2(n14990), .ZN(n14993) );
  INV_X1 U13386 ( .A(n15023), .ZN(n10824) );
  NOR2_X1 U13387 ( .A1(n10817), .A2(n10824), .ZN(n15010) );
  NAND2_X1 U13388 ( .A1(n10817), .A2(n10824), .ZN(n15011) );
  OAI21_X1 U13389 ( .B1(n15014), .B2(n15010), .A(n15011), .ZN(n10855) );
  XOR2_X1 U13390 ( .A(n10854), .B(n10855), .Z(n10851) );
  INV_X1 U13391 ( .A(n15078), .ZN(n15054) );
  INV_X1 U13392 ( .A(n15052), .ZN(n15080) );
  INV_X1 U13393 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n10832) );
  NAND2_X1 U13394 ( .A1(n10834), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10818) );
  NAND2_X1 U13395 ( .A1(n10819), .A2(n10818), .ZN(n10820) );
  MUX2_X1 U13396 ( .A(n10822), .B(P3_REG2_REG_4__SCAN_IN), .S(n15005), .Z(
        n14998) );
  NOR2_X1 U13397 ( .A1(n10824), .A2(n10823), .ZN(n10825) );
  NOR2_X1 U13398 ( .A1(n10825), .A2(n15017), .ZN(n10828) );
  MUX2_X1 U13399 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n10826), .S(n10858), .Z(
        n10827) );
  NOR2_X1 U13400 ( .A1(n10828), .A2(n10827), .ZN(n10865) );
  AOI21_X1 U13401 ( .B1(n10828), .B2(n10827), .A(n10865), .ZN(n10829) );
  INV_X1 U13402 ( .A(n10829), .ZN(n10830) );
  NAND2_X1 U13403 ( .A1(n15082), .A2(n10830), .ZN(n10831) );
  NAND2_X1 U13404 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n11061) );
  OAI211_X1 U13405 ( .C1(n15043), .C2(n10832), .A(n10831), .B(n11061), .ZN(
        n10833) );
  AOI21_X1 U13406 ( .B1(n15080), .B2(n10858), .A(n10833), .ZN(n10850) );
  NAND2_X1 U13407 ( .A1(n10834), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10835) );
  NAND2_X1 U13408 ( .A1(n10836), .A2(n10835), .ZN(n10838) );
  XNOR2_X1 U13409 ( .A(n10838), .B(n10837), .ZN(n14985) );
  NAND2_X1 U13410 ( .A1(n14985), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n10840) );
  NAND2_X1 U13411 ( .A1(n10838), .A2(n14976), .ZN(n10839) );
  NAND2_X1 U13412 ( .A1(n10840), .A2(n10839), .ZN(n14995) );
  MUX2_X1 U13413 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n10841), .S(n15005), .Z(
        n14996) );
  NAND2_X1 U13414 ( .A1(n14995), .A2(n14996), .ZN(n14994) );
  NAND2_X1 U13415 ( .A1(n15023), .A2(n10843), .ZN(n10844) );
  MUX2_X1 U13416 ( .A(n10845), .B(P3_REG1_REG_6__SCAN_IN), .S(n10858), .Z(
        n10846) );
  NAND2_X1 U13417 ( .A1(n10847), .A2(n10846), .ZN(n10857) );
  OAI21_X1 U13418 ( .B1(n10847), .B2(n10846), .A(n10857), .ZN(n10848) );
  NAND2_X1 U13419 ( .A1(n10848), .A2(n15069), .ZN(n10849) );
  OAI211_X1 U13420 ( .C1(n10851), .C2(n15054), .A(n10850), .B(n10849), .ZN(
        P3_U3188) );
  XNOR2_X1 U13421 ( .A(n11381), .B(n11383), .ZN(n11384) );
  INV_X1 U13422 ( .A(n10852), .ZN(n10853) );
  AOI22_X1 U13423 ( .A1(n10855), .A2(n10854), .B1(n10858), .B2(n10853), .ZN(
        n15030) );
  XNOR2_X1 U13424 ( .A(n10856), .B(n15035), .ZN(n15029) );
  OAI22_X1 U13425 ( .A1(n15030), .A2(n15029), .B1(n10856), .B2(n15035), .ZN(
        n11385) );
  XOR2_X1 U13426 ( .A(n11384), .B(n11385), .Z(n10879) );
  OAI21_X1 U13427 ( .B1(n10858), .B2(n10845), .A(n10857), .ZN(n10859) );
  NAND2_X1 U13428 ( .A1(n15035), .A2(n10859), .ZN(n10861) );
  INV_X1 U13429 ( .A(n15035), .ZN(n10867) );
  XNOR2_X1 U13430 ( .A(n10859), .B(n10867), .ZN(n15034) );
  NAND2_X1 U13431 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n15034), .ZN(n10860) );
  MUX2_X1 U13432 ( .A(n10862), .B(P3_REG1_REG_8__SCAN_IN), .S(n11383), .Z(
        n10863) );
  OAI21_X1 U13433 ( .B1(n10864), .B2(n10863), .A(n11377), .ZN(n10877) );
  NOR2_X1 U13434 ( .A1(n15052), .A2(n6839), .ZN(n10876) );
  NOR2_X1 U13435 ( .A1(n10867), .A2(n10868), .ZN(n10869) );
  XOR2_X1 U13436 ( .A(n10868), .B(n15035), .Z(n15032) );
  NOR2_X1 U13437 ( .A1(n11414), .A2(n15032), .ZN(n15031) );
  NOR2_X1 U13438 ( .A1(n10869), .A2(n15031), .ZN(n10872) );
  MUX2_X1 U13439 ( .A(P3_REG2_REG_8__SCAN_IN), .B(n10870), .S(n11383), .Z(
        n10871) );
  NOR2_X1 U13440 ( .A1(n10872), .A2(n10871), .ZN(n11373) );
  AOI21_X1 U13441 ( .B1(n10872), .B2(n10871), .A(n11373), .ZN(n10874) );
  NAND2_X1 U13442 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n11359) );
  NAND2_X1 U13443 ( .A1(n15068), .A2(P3_ADDR_REG_8__SCAN_IN), .ZN(n10873) );
  OAI211_X1 U13444 ( .C1(n15063), .C2(n10874), .A(n11359), .B(n10873), .ZN(
        n10875) );
  AOI211_X1 U13445 ( .C1(n10877), .C2(n15069), .A(n10876), .B(n10875), .ZN(
        n10878) );
  OAI21_X1 U13446 ( .B1(n10879), .B2(n15054), .A(n10878), .ZN(P3_U3190) );
  OAI222_X1 U13447 ( .A1(P3_U3151), .A2(n10881), .B1(n13078), .B2(n15324), 
        .C1(n13076), .C2(n10880), .ZN(P3_U3275) );
  INV_X1 U13448 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n15284) );
  OAI22_X1 U13449 ( .A1(n12649), .A2(n15129), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15284), .ZN(n10882) );
  AOI21_X1 U13450 ( .B1(n10675), .B2(n12673), .A(n10882), .ZN(n10883) );
  OAI21_X1 U13451 ( .B1(n10884), .B2(n12632), .A(n10883), .ZN(n10889) );
  AOI211_X1 U13452 ( .C1(n10887), .C2(n10886), .A(n12637), .B(n10885), .ZN(
        n10888) );
  AOI211_X1 U13453 ( .C1(n15284), .C2(n12629), .A(n10889), .B(n10888), .ZN(
        n10890) );
  INV_X1 U13454 ( .A(n10890), .ZN(P3_U3158) );
  NAND2_X1 U13455 ( .A1(n10891), .A2(n12364), .ZN(n10892) );
  NAND2_X1 U13456 ( .A1(n10892), .A2(n13062), .ZN(n10896) );
  NAND2_X1 U13457 ( .A1(n10894), .A2(n10893), .ZN(n10895) );
  NAND3_X1 U13458 ( .A1(n10897), .A2(n10896), .A3(n10895), .ZN(n10899) );
  NAND2_X2 U13459 ( .A1(n10899), .A2(n15112), .ZN(n15117) );
  INV_X1 U13460 ( .A(n11083), .ZN(n10898) );
  NAND2_X1 U13461 ( .A1(n10898), .A2(n15117), .ZN(n10901) );
  INV_X1 U13462 ( .A(n15111), .ZN(n15090) );
  AOI22_X1 U13463 ( .A1(n14402), .A2(n8873), .B1(n14400), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n10900) );
  OAI211_X1 U13464 ( .C1(n10731), .C2(n15117), .A(n10901), .B(n10900), .ZN(
        P3_U3233) );
  NOR3_X1 U13465 ( .A1(n15069), .A2(n15082), .A3(n15078), .ZN(n10912) );
  INV_X1 U13466 ( .A(n10902), .ZN(n10903) );
  NAND2_X1 U13467 ( .A1(n15078), .A2(n10903), .ZN(n10904) );
  MUX2_X1 U13468 ( .A(n10904), .B(n15052), .S(P3_IR_REG_0__SCAN_IN), .Z(n10910) );
  AOI22_X1 U13469 ( .A1(n15068), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n10905) );
  OAI21_X1 U13470 ( .B1(n10906), .B2(n15036), .A(n10905), .ZN(n10907) );
  AOI21_X1 U13471 ( .B1(n15082), .B2(n10908), .A(n10907), .ZN(n10909) );
  OAI211_X1 U13472 ( .C1(n10912), .C2(n10911), .A(n10910), .B(n10909), .ZN(
        P3_U3182) );
  INV_X1 U13473 ( .A(n13916), .ZN(n14610) );
  OAI222_X1 U13474 ( .A1(n14208), .A2(n10915), .B1(n14610), .B2(P1_U3086), 
        .C1(n10913), .C2(n12044), .ZN(P1_U3337) );
  INV_X1 U13475 ( .A(n13305), .ZN(n10914) );
  OAI222_X1 U13476 ( .A1(n13652), .A2(n10916), .B1(n13643), .B2(n10915), .C1(
        P2_U3088), .C2(n10914), .ZN(P2_U3309) );
  INV_X1 U13477 ( .A(n10917), .ZN(n10921) );
  INV_X1 U13478 ( .A(n10918), .ZN(n10920) );
  NAND2_X1 U13479 ( .A1(n12446), .A2(n13841), .ZN(n10924) );
  NAND2_X1 U13480 ( .A1(n14676), .A2(n12424), .ZN(n10923) );
  NAND2_X1 U13481 ( .A1(n10924), .A2(n10923), .ZN(n11486) );
  NAND2_X1 U13482 ( .A1(n13841), .A2(n12424), .ZN(n10926) );
  NAND2_X1 U13483 ( .A1(n14676), .A2(n12441), .ZN(n10925) );
  NAND2_X1 U13484 ( .A1(n10926), .A2(n10925), .ZN(n10927) );
  XNOR2_X1 U13485 ( .A(n10927), .B(n12444), .ZN(n11487) );
  XOR2_X1 U13486 ( .A(n11486), .B(n11487), .Z(n10928) );
  OAI211_X1 U13487 ( .C1(n10929), .C2(n10928), .A(n11491), .B(n13795), .ZN(
        n10934) );
  INV_X1 U13488 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n13872) );
  NAND2_X1 U13489 ( .A1(n10930), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10931) );
  NAND2_X1 U13490 ( .A1(n10931), .A2(n11828), .ZN(n13798) );
  AOI22_X1 U13491 ( .A1(n14482), .A2(n13842), .B1(n13840), .B2(n14631), .ZN(
        n14670) );
  OAI22_X1 U13492 ( .A1(n14670), .A2(n13778), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13872), .ZN(n10932) );
  AOI21_X1 U13493 ( .B1(n13872), .B2(n13798), .A(n10932), .ZN(n10933) );
  OAI211_X1 U13494 ( .C1(n14711), .C2(n13803), .A(n10934), .B(n10933), .ZN(
        P1_U3218) );
  OAI21_X1 U13495 ( .B1(n10937), .B2(n10936), .A(n10935), .ZN(n10938) );
  NAND2_X1 U13496 ( .A1(n10938), .A2(n12642), .ZN(n10942) );
  NAND2_X1 U13497 ( .A1(n10675), .A2(n12672), .ZN(n10939) );
  NAND2_X1 U13498 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_U3151), .ZN(n15007) );
  OAI211_X1 U13499 ( .C1(n12649), .C2(n15134), .A(n10939), .B(n15007), .ZN(
        n10940) );
  AOI21_X1 U13500 ( .B1(n12552), .B2(n15091), .A(n10940), .ZN(n10941) );
  OAI211_X1 U13501 ( .C1(n11041), .C2(n12645), .A(n10942), .B(n10941), .ZN(
        P3_U3170) );
  OAI22_X1 U13502 ( .A1(n13472), .A2(n10944), .B1(n13518), .B2(n10943), .ZN(
        n10945) );
  AOI21_X1 U13503 ( .B1(n14916), .B2(n10946), .A(n10945), .ZN(n10950) );
  INV_X1 U13504 ( .A(n14919), .ZN(n14903) );
  MUX2_X1 U13505 ( .A(n10948), .B(n10947), .S(n14903), .Z(n10949) );
  OAI211_X1 U13506 ( .C1(n13528), .C2(n10951), .A(n10950), .B(n10949), .ZN(
        P2_U3264) );
  MUX2_X1 U13507 ( .A(n10953), .B(n10952), .S(n14919), .Z(n10959) );
  OAI22_X1 U13508 ( .A1(n13472), .A2(n10955), .B1(n10954), .B2(n13518), .ZN(
        n10956) );
  AOI21_X1 U13509 ( .B1(n10957), .B2(n14916), .A(n10956), .ZN(n10958) );
  OAI211_X1 U13510 ( .C1(n10960), .C2(n13528), .A(n10959), .B(n10958), .ZN(
        P2_U3261) );
  INV_X1 U13511 ( .A(n10961), .ZN(n12394) );
  NAND2_X1 U13512 ( .A1(n12394), .A2(n10962), .ZN(n10963) );
  NAND2_X1 U13513 ( .A1(n12397), .A2(n10963), .ZN(n10964) );
  XNOR2_X1 U13514 ( .A(n12391), .B(n6725), .ZN(n10965) );
  NAND2_X1 U13515 ( .A1(n13261), .A2(n13105), .ZN(n10966) );
  XNOR2_X1 U13516 ( .A(n10965), .B(n10966), .ZN(n12392) );
  INV_X1 U13517 ( .A(n10965), .ZN(n10967) );
  NAND2_X1 U13518 ( .A1(n10967), .A2(n10966), .ZN(n10968) );
  XNOR2_X1 U13519 ( .A(n11052), .B(n13134), .ZN(n11070) );
  NAND2_X1 U13520 ( .A1(n13260), .A2(n13105), .ZN(n11071) );
  XNOR2_X1 U13521 ( .A(n11070), .B(n11071), .ZN(n10970) );
  AOI21_X1 U13522 ( .B1(n10969), .B2(n10970), .A(n14782), .ZN(n10972) );
  NAND2_X1 U13523 ( .A1(n10972), .A2(n11075), .ZN(n10978) );
  NAND2_X1 U13524 ( .A1(n13261), .A2(n13231), .ZN(n10974) );
  NAND2_X1 U13525 ( .A1(n13259), .A2(n13233), .ZN(n10973) );
  NAND2_X1 U13526 ( .A1(n10974), .A2(n10973), .ZN(n11049) );
  NOR2_X1 U13527 ( .A1(n14789), .A2(n11258), .ZN(n10975) );
  AOI211_X1 U13528 ( .C1(n14430), .C2(n11049), .A(n10976), .B(n10975), .ZN(
        n10977) );
  OAI211_X1 U13529 ( .C1(n6938), .C2(n13210), .A(n10978), .B(n10977), .ZN(
        P2_U3189) );
  OAI22_X1 U13530 ( .A1(n14919), .A2(n10117), .B1(n10979), .B2(n13518), .ZN(
        n10982) );
  NOR2_X1 U13531 ( .A1(n13472), .A2(n10980), .ZN(n10981) );
  AOI211_X1 U13532 ( .C1(n10983), .C2(n14916), .A(n10982), .B(n10981), .ZN(
        n10986) );
  NAND2_X1 U13533 ( .A1(n10984), .A2(n14900), .ZN(n10985) );
  OAI211_X1 U13534 ( .C1(n14903), .C2(n10987), .A(n10986), .B(n10985), .ZN(
        P2_U3263) );
  XNOR2_X1 U13535 ( .A(n10988), .B(n10991), .ZN(n14951) );
  INV_X1 U13536 ( .A(n14951), .ZN(n11003) );
  OAI21_X1 U13537 ( .B1(n10991), .B2(n10990), .A(n10989), .ZN(n10992) );
  NAND2_X1 U13538 ( .A1(n10992), .A2(n14886), .ZN(n10994) );
  NAND2_X1 U13539 ( .A1(n10994), .A2(n10993), .ZN(n10995) );
  AOI21_X1 U13540 ( .B1(n14951), .B2(n9471), .A(n10995), .ZN(n14953) );
  MUX2_X1 U13541 ( .A(n10996), .B(n14953), .S(n14919), .Z(n11002) );
  OAI21_X1 U13542 ( .B1(n11217), .B2(n10999), .A(n13523), .ZN(n10997) );
  NOR2_X1 U13543 ( .A1(n10997), .A2(n11209), .ZN(n14948) );
  OAI22_X1 U13544 ( .A1(n10999), .A2(n13472), .B1(n10998), .B2(n13518), .ZN(
        n11000) );
  AOI21_X1 U13545 ( .B1(n14948), .B2(n14916), .A(n11000), .ZN(n11001) );
  OAI211_X1 U13546 ( .C1(n11003), .C2(n14912), .A(n11002), .B(n11001), .ZN(
        P2_U3257) );
  INV_X1 U13547 ( .A(SI_21_), .ZN(n15260) );
  OAI222_X1 U13548 ( .A1(P3_U3151), .A2(n12211), .B1(n13078), .B2(n15260), 
        .C1(n13076), .C2(n11004), .ZN(P3_U3274) );
  XOR2_X1 U13549 ( .A(n11005), .B(n6482), .Z(n14697) );
  INV_X1 U13550 ( .A(n11006), .ZN(n11007) );
  NAND2_X1 U13551 ( .A1(n14665), .A2(n11007), .ZN(n14645) );
  NAND2_X1 U13552 ( .A1(n14480), .A2(n8333), .ZN(n14730) );
  INV_X1 U13553 ( .A(n11008), .ZN(n11015) );
  AOI21_X1 U13554 ( .B1(n6482), .B2(n13843), .A(n14690), .ZN(n11013) );
  NAND2_X1 U13555 ( .A1(n6493), .A2(n14694), .ZN(n11009) );
  NAND2_X1 U13556 ( .A1(n11118), .A2(n11009), .ZN(n14700) );
  XNOR2_X1 U13557 ( .A(n11150), .B(n14700), .ZN(n11011) );
  OAI21_X1 U13558 ( .B1(n11011), .B2(n14690), .A(n11010), .ZN(n11012) );
  OAI21_X1 U13559 ( .B1(n11013), .B2(n14482), .A(n11012), .ZN(n11014) );
  OAI211_X1 U13560 ( .C1(n14697), .C2(n14730), .A(n11015), .B(n11014), .ZN(
        n14701) );
  NAND2_X1 U13561 ( .A1(n14701), .A2(n14665), .ZN(n11021) );
  INV_X1 U13562 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n11016) );
  OAI22_X1 U13563 ( .A1(n14665), .A2(n10154), .B1(n11016), .B2(n14673), .ZN(
        n11018) );
  NOR2_X1 U13564 ( .A1(n14065), .A2(n14699), .ZN(n14491) );
  INV_X1 U13565 ( .A(n14491), .ZN(n11154) );
  NOR2_X1 U13566 ( .A1(n11154), .A2(n14700), .ZN(n11017) );
  AOI211_X1 U13567 ( .C1(n14677), .C2(n6493), .A(n11018), .B(n11017), .ZN(
        n11020) );
  OAI211_X1 U13568 ( .C1(n14697), .C2(n14645), .A(n11021), .B(n11020), .ZN(
        P1_U3292) );
  XOR2_X1 U13569 ( .A(n11023), .B(n11022), .Z(n11028) );
  NAND2_X1 U13570 ( .A1(n10675), .A2(n12671), .ZN(n11024) );
  NAND2_X1 U13571 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(P3_U3151), .ZN(n15026) );
  OAI211_X1 U13572 ( .C1(n12649), .C2(n15139), .A(n11024), .B(n15026), .ZN(
        n11026) );
  NOR2_X1 U13573 ( .A1(n12645), .A2(n11127), .ZN(n11025) );
  AOI211_X1 U13574 ( .C1(n12552), .C2(n12673), .A(n11026), .B(n11025), .ZN(
        n11027) );
  OAI21_X1 U13575 ( .B1(n11028), .B2(n12637), .A(n11027), .ZN(P3_U3167) );
  NOR2_X1 U13576 ( .A1(n13078), .A2(SI_22_), .ZN(n11029) );
  AOI21_X1 U13577 ( .B1(n11030), .B2(P3_STATE_REG_SCAN_IN), .A(n11029), .ZN(
        n11031) );
  OAI21_X1 U13578 ( .B1(n11032), .B2(n13076), .A(n11031), .ZN(n11033) );
  INV_X1 U13579 ( .A(n11033), .ZN(P3_U3273) );
  XNOR2_X1 U13580 ( .A(n11035), .B(n11034), .ZN(n11040) );
  AOI22_X1 U13581 ( .A1(n15104), .A2(n12672), .B1(n15091), .B2(n15103), .ZN(
        n11039) );
  OAI21_X1 U13582 ( .B1(n11037), .B2(n12228), .A(n11036), .ZN(n15137) );
  INV_X1 U13583 ( .A(n15110), .ZN(n12815) );
  NAND2_X1 U13584 ( .A1(n15137), .A2(n12815), .ZN(n11038) );
  OAI211_X1 U13585 ( .C1(n11040), .C2(n12922), .A(n11039), .B(n11038), .ZN(
        n15135) );
  INV_X1 U13586 ( .A(n15135), .ZN(n11045) );
  INV_X2 U13587 ( .A(n15117), .ZN(n15119) );
  OR2_X1 U13588 ( .A1(n15111), .A2(n12211), .ZN(n11766) );
  INV_X1 U13589 ( .A(n11766), .ZN(n15100) );
  NAND2_X1 U13590 ( .A1(n15117), .A2(n15100), .ZN(n15114) );
  INV_X1 U13591 ( .A(n15114), .ZN(n12816) );
  NOR2_X1 U13592 ( .A1(n15117), .A2(n10822), .ZN(n11043) );
  OAI22_X1 U13593 ( .A1(n12933), .A2(n15134), .B1(n11041), .B2(n15112), .ZN(
        n11042) );
  AOI211_X1 U13594 ( .C1(n15137), .C2(n12816), .A(n11043), .B(n11042), .ZN(
        n11044) );
  OAI21_X1 U13595 ( .B1(n11045), .B2(n15119), .A(n11044), .ZN(P3_U3229) );
  XNOR2_X1 U13596 ( .A(n11046), .B(n7087), .ZN(n11261) );
  XNOR2_X1 U13597 ( .A(n11048), .B(n11047), .ZN(n11050) );
  AOI21_X1 U13598 ( .B1(n11050), .B2(n14886), .A(n11049), .ZN(n11266) );
  AOI21_X1 U13599 ( .B1(n11208), .B2(n11052), .A(n13489), .ZN(n11051) );
  AND2_X1 U13600 ( .A1(n11051), .A2(n11272), .ZN(n11264) );
  AOI21_X1 U13601 ( .B1(n11052), .B2(n14945), .A(n11264), .ZN(n11053) );
  OAI211_X1 U13602 ( .C1(n11261), .C2(n13614), .A(n11266), .B(n11053), .ZN(
        n11055) );
  NAND2_X1 U13603 ( .A1(n11055), .A2(n14964), .ZN(n11054) );
  OAI21_X1 U13604 ( .B1(n14964), .B2(n9135), .A(n11054), .ZN(P2_U3460) );
  NAND2_X1 U13605 ( .A1(n11055), .A2(n13616), .ZN(n11056) );
  OAI21_X1 U13606 ( .B1(n13616), .B2(n11057), .A(n11056), .ZN(P2_U3509) );
  OAI211_X1 U13607 ( .C1(n11060), .C2(n11059), .A(n11058), .B(n12642), .ZN(
        n11065) );
  NAND2_X1 U13608 ( .A1(n10675), .A2(n12670), .ZN(n11062) );
  OAI211_X1 U13609 ( .C1(n15144), .C2(n12649), .A(n11062), .B(n11061), .ZN(
        n11063) );
  AOI21_X1 U13610 ( .B1(n12552), .B2(n12672), .A(n11063), .ZN(n11064) );
  OAI211_X1 U13611 ( .C1(n11188), .C2(n12645), .A(n11065), .B(n11064), .ZN(
        P3_U3179) );
  XNOR2_X1 U13612 ( .A(n14955), .B(n13134), .ZN(n11066) );
  NAND2_X1 U13613 ( .A1(n13259), .A2(n13105), .ZN(n11067) );
  NAND2_X1 U13614 ( .A1(n11066), .A2(n11067), .ZN(n11342) );
  INV_X1 U13615 ( .A(n11066), .ZN(n11069) );
  INV_X1 U13616 ( .A(n11067), .ZN(n11068) );
  NAND2_X1 U13617 ( .A1(n11069), .A2(n11068), .ZN(n11344) );
  NAND2_X1 U13618 ( .A1(n11342), .A2(n11344), .ZN(n11076) );
  INV_X1 U13619 ( .A(n11070), .ZN(n11073) );
  INV_X1 U13620 ( .A(n11071), .ZN(n11072) );
  NAND2_X1 U13621 ( .A1(n11073), .A2(n11072), .ZN(n11074) );
  XOR2_X1 U13622 ( .A(n11076), .B(n11343), .Z(n11082) );
  OAI22_X1 U13623 ( .A1(n11078), .A2(n14420), .B1(n11077), .B2(n14422), .ZN(
        n11268) );
  AOI22_X1 U13624 ( .A1(n14430), .A2(n11268), .B1(P2_REG3_REG_11__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11079) );
  OAI21_X1 U13625 ( .B1(n11275), .B2(n14789), .A(n11079), .ZN(n11080) );
  AOI21_X1 U13626 ( .B1(n14955), .B2(n14787), .A(n11080), .ZN(n11081) );
  OAI21_X1 U13627 ( .B1(n11082), .B2(n14782), .A(n11081), .ZN(P2_U3208) );
  MUX2_X1 U13628 ( .A(n10730), .B(n11083), .S(n15183), .Z(n11084) );
  OAI21_X1 U13629 ( .B1(n10681), .B2(n13003), .A(n11084), .ZN(P3_U3459) );
  OAI21_X1 U13630 ( .B1(n14485), .B2(n11088), .A(n11085), .ZN(n11299) );
  XNOR2_X1 U13631 ( .A(n11299), .B(n11300), .ZN(n11086) );
  NOR2_X1 U13632 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n11086), .ZN(n11301) );
  AOI21_X1 U13633 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n11086), .A(n11301), 
        .ZN(n11097) );
  AOI21_X1 U13634 ( .B1(n11088), .B2(n7860), .A(n11087), .ZN(n11288) );
  XOR2_X1 U13635 ( .A(n11288), .B(n11092), .Z(n11089) );
  NOR2_X1 U13636 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n11089), .ZN(n11289) );
  AOI21_X1 U13637 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n11089), .A(n11289), 
        .ZN(n11091) );
  OR2_X1 U13638 ( .A1(n11091), .A2(n11090), .ZN(n11096) );
  NOR2_X1 U13639 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n13806), .ZN(n11094) );
  NOR2_X1 U13640 ( .A1(n14611), .A2(n11092), .ZN(n11093) );
  AOI211_X1 U13641 ( .C1(n14587), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n11094), 
        .B(n11093), .ZN(n11095) );
  OAI211_X1 U13642 ( .C1(n11097), .C2(n13920), .A(n11096), .B(n11095), .ZN(
        P1_U3258) );
  XNOR2_X1 U13643 ( .A(n11098), .B(n11107), .ZN(n11239) );
  INV_X1 U13644 ( .A(n11239), .ZN(n11110) );
  NAND2_X1 U13645 ( .A1(n13835), .A2(n14631), .ZN(n11100) );
  NAND2_X1 U13646 ( .A1(n13837), .A2(n14482), .ZN(n11099) );
  AND2_X1 U13647 ( .A1(n11100), .A2(n11099), .ZN(n11606) );
  MUX2_X1 U13648 ( .A(n11101), .B(n11606), .S(n14665), .Z(n11102) );
  OAI21_X1 U13649 ( .B1(n14673), .B2(n11604), .A(n11102), .ZN(n11105) );
  AOI21_X1 U13650 ( .B1(n6517), .B2(n11589), .A(n14699), .ZN(n11103) );
  NAND2_X1 U13651 ( .A1(n11103), .A2(n11427), .ZN(n11242) );
  NOR2_X1 U13652 ( .A1(n11242), .A2(n14065), .ZN(n11104) );
  AOI211_X1 U13653 ( .C1(n14677), .C2(n11589), .A(n11105), .B(n11104), .ZN(
        n11109) );
  NAND2_X1 U13654 ( .A1(n11106), .A2(n11107), .ZN(n11241) );
  NOR2_X1 U13655 ( .A1(n14087), .A2(n14690), .ZN(n14035) );
  NAND3_X1 U13656 ( .A1(n6470), .A2(n11241), .A3(n14035), .ZN(n11108) );
  OAI211_X1 U13657 ( .C1(n11110), .C2(n14083), .A(n11109), .B(n11108), .ZN(
        P1_U3285) );
  XNOR2_X1 U13658 ( .A(n11112), .B(n11111), .ZN(n14704) );
  XNOR2_X1 U13659 ( .A(n11113), .B(n11114), .ZN(n11117) );
  INV_X1 U13660 ( .A(n11115), .ZN(n11116) );
  OAI21_X1 U13661 ( .B1(n11117), .B2(n14690), .A(n11116), .ZN(n14707) );
  NAND2_X1 U13662 ( .A1(n14707), .A2(n14665), .ZN(n11123) );
  AOI211_X1 U13663 ( .C1(n11119), .C2(n11118), .A(n14699), .B(n14681), .ZN(
        n14706) );
  AOI22_X1 U13664 ( .A1(n14644), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n14643), .ZN(n11120) );
  OAI21_X1 U13665 ( .B1(n14488), .B2(n14705), .A(n11120), .ZN(n11121) );
  AOI21_X1 U13666 ( .B1(n14706), .B2(n14683), .A(n11121), .ZN(n11122) );
  OAI211_X1 U13667 ( .C1(n14704), .C2(n14083), .A(n11123), .B(n11122), .ZN(
        P1_U3291) );
  OR2_X1 U13668 ( .A1(n11124), .A2(n12230), .ZN(n11125) );
  AND2_X1 U13669 ( .A1(n11126), .A2(n11125), .ZN(n15140) );
  INV_X1 U13670 ( .A(n15140), .ZN(n11136) );
  OAI22_X1 U13671 ( .A1(n12933), .A2(n15139), .B1(n11127), .B2(n15112), .ZN(
        n11135) );
  AOI22_X1 U13672 ( .A1(n15103), .A2(n12673), .B1(n12671), .B2(n15104), .ZN(
        n11133) );
  OAI21_X1 U13673 ( .B1(n11128), .B2(n11130), .A(n11129), .ZN(n11131) );
  NAND2_X1 U13674 ( .A1(n11131), .A2(n15106), .ZN(n11132) );
  OAI211_X1 U13675 ( .C1(n15140), .C2(n15110), .A(n11133), .B(n11132), .ZN(
        n15142) );
  MUX2_X1 U13676 ( .A(P3_REG2_REG_5__SCAN_IN), .B(n15142), .S(n15117), .Z(
        n11134) );
  AOI211_X1 U13677 ( .C1(n12816), .C2(n11136), .A(n11135), .B(n11134), .ZN(
        n11137) );
  INV_X1 U13678 ( .A(n11137), .ZN(P3_U3228) );
  XNOR2_X1 U13679 ( .A(n11138), .B(n11140), .ZN(n14729) );
  XNOR2_X1 U13680 ( .A(n11139), .B(n11140), .ZN(n11143) );
  NAND2_X1 U13681 ( .A1(n13837), .A2(n14631), .ZN(n11142) );
  NAND2_X1 U13682 ( .A1(n13839), .A2(n14482), .ZN(n11141) );
  AND2_X1 U13683 ( .A1(n11142), .A2(n11141), .ZN(n11485) );
  OAI21_X1 U13684 ( .B1(n11143), .B2(n14690), .A(n11485), .ZN(n14734) );
  INV_X1 U13685 ( .A(n14734), .ZN(n11145) );
  MUX2_X1 U13686 ( .A(n11145), .B(n11144), .S(n14644), .Z(n11149) );
  OAI211_X1 U13687 ( .C1(n11179), .C2(n14732), .A(n14646), .B(n14679), .ZN(
        n14731) );
  INV_X1 U13688 ( .A(n14731), .ZN(n11147) );
  OAI22_X1 U13689 ( .A1(n14488), .A2(n14732), .B1(n11481), .B2(n14673), .ZN(
        n11146) );
  AOI21_X1 U13690 ( .B1(n11147), .B2(n14683), .A(n11146), .ZN(n11148) );
  OAI211_X1 U13691 ( .C1(n14083), .C2(n14729), .A(n11149), .B(n11148), .ZN(
        P1_U3287) );
  NOR2_X1 U13692 ( .A1(n14035), .A2(n14662), .ZN(n11158) );
  NOR2_X1 U13693 ( .A1(n11150), .A2(n14055), .ZN(n14693) );
  OAI22_X1 U13694 ( .A1(n14665), .A2(n11152), .B1(n11151), .B2(n14673), .ZN(
        n11156) );
  AOI21_X1 U13695 ( .B1(n14488), .B2(n11154), .A(n11153), .ZN(n11155) );
  AOI211_X1 U13696 ( .C1(n14693), .C2(n14665), .A(n11156), .B(n11155), .ZN(
        n11157) );
  OAI21_X1 U13697 ( .B1(n14689), .B2(n11158), .A(n11157), .ZN(P1_U3293) );
  XOR2_X1 U13698 ( .A(n11159), .B(n11163), .Z(n14932) );
  OAI211_X1 U13699 ( .C1(n11160), .C2(n14930), .A(n14895), .B(n13523), .ZN(
        n14928) );
  NOR2_X1 U13700 ( .A1(n14928), .A2(n14898), .ZN(n11162) );
  OAI22_X1 U13701 ( .A1(n13472), .A2(n14930), .B1(n13518), .B2(n12028), .ZN(
        n11161) );
  AOI211_X1 U13702 ( .C1(n14932), .C2(n14900), .A(n11162), .B(n11161), .ZN(
        n11170) );
  XNOR2_X1 U13703 ( .A(n11164), .B(n11163), .ZN(n11167) );
  OAI22_X1 U13704 ( .A1(n11166), .A2(n14422), .B1(n11165), .B2(n14420), .ZN(
        n12029) );
  AOI21_X1 U13705 ( .B1(n11167), .B2(n14886), .A(n12029), .ZN(n14929) );
  MUX2_X1 U13706 ( .A(n11168), .B(n14929), .S(n14919), .Z(n11169) );
  NAND2_X1 U13707 ( .A1(n11170), .A2(n11169), .ZN(P2_U3260) );
  XNOR2_X1 U13708 ( .A(n11171), .B(n11172), .ZN(n11177) );
  INV_X1 U13709 ( .A(n11177), .ZN(n14727) );
  INV_X1 U13710 ( .A(n14730), .ZN(n14750) );
  XNOR2_X1 U13711 ( .A(n11173), .B(n11172), .ZN(n11175) );
  AOI22_X1 U13712 ( .A1(n13840), .A2(n14482), .B1(n14631), .B2(n13838), .ZN(
        n11174) );
  OAI21_X1 U13713 ( .B1(n11175), .B2(n14690), .A(n11174), .ZN(n11176) );
  AOI21_X1 U13714 ( .B1(n11177), .B2(n14750), .A(n11176), .ZN(n14726) );
  MUX2_X1 U13715 ( .A(n11178), .B(n14726), .S(n14665), .Z(n11182) );
  AOI211_X1 U13716 ( .C1(n14724), .C2(n14660), .A(n14699), .B(n11179), .ZN(
        n14722) );
  OAI22_X1 U13717 ( .A1(n14488), .A2(n11494), .B1(n14673), .B2(n13726), .ZN(
        n11180) );
  AOI21_X1 U13718 ( .B1(n14722), .B2(n14683), .A(n11180), .ZN(n11181) );
  OAI211_X1 U13719 ( .C1(n14727), .C2(n14645), .A(n11182), .B(n11181), .ZN(
        P1_U3288) );
  XNOR2_X1 U13720 ( .A(n11183), .B(n11185), .ZN(n15145) );
  OAI211_X1 U13721 ( .C1(n6520), .C2(n11185), .A(n15106), .B(n11184), .ZN(
        n11187) );
  AOI22_X1 U13722 ( .A1(n15104), .A2(n12670), .B1(n12672), .B2(n15103), .ZN(
        n11186) );
  OAI211_X1 U13723 ( .C1(n15145), .C2(n15110), .A(n11187), .B(n11186), .ZN(
        n15147) );
  NAND2_X1 U13724 ( .A1(n15147), .A2(n15117), .ZN(n11191) );
  OAI22_X1 U13725 ( .A1(n12933), .A2(n15144), .B1(n11188), .B2(n15112), .ZN(
        n11189) );
  AOI21_X1 U13726 ( .B1(n15119), .B2(P3_REG2_REG_6__SCAN_IN), .A(n11189), .ZN(
        n11190) );
  OAI211_X1 U13727 ( .C1(n15145), .C2(n15114), .A(n11191), .B(n11190), .ZN(
        P3_U3227) );
  XNOR2_X1 U13728 ( .A(n11194), .B(n11192), .ZN(n15130) );
  AOI22_X1 U13729 ( .A1(n15103), .A2(n9772), .B1(n12673), .B2(n15104), .ZN(
        n11197) );
  OAI211_X1 U13730 ( .C1(n11195), .C2(n11194), .A(n15106), .B(n11193), .ZN(
        n11196) );
  OAI211_X1 U13731 ( .C1(n15130), .C2(n15110), .A(n11197), .B(n11196), .ZN(
        n15132) );
  NAND2_X1 U13732 ( .A1(n15132), .A2(n15117), .ZN(n11200) );
  OAI22_X1 U13733 ( .A1(n12933), .A2(n15129), .B1(n15112), .B2(
        P3_REG3_REG_3__SCAN_IN), .ZN(n11198) );
  AOI21_X1 U13734 ( .B1(n15119), .B2(P3_REG2_REG_3__SCAN_IN), .A(n11198), .ZN(
        n11199) );
  OAI211_X1 U13735 ( .C1(n15130), .C2(n15114), .A(n11200), .B(n11199), .ZN(
        P3_U3230) );
  XNOR2_X1 U13736 ( .A(n11201), .B(n11202), .ZN(n11252) );
  INV_X1 U13737 ( .A(n11252), .ZN(n11214) );
  XNOR2_X1 U13738 ( .A(n11204), .B(n11203), .ZN(n11206) );
  NAND2_X1 U13739 ( .A1(n11252), .A2(n9471), .ZN(n11205) );
  AOI22_X1 U13740 ( .A1(n13231), .A2(n13262), .B1(n13260), .B2(n13233), .ZN(
        n12388) );
  OAI211_X1 U13741 ( .C1(n7099), .C2(n11206), .A(n11205), .B(n12388), .ZN(
        n11250) );
  NAND2_X1 U13742 ( .A1(n11250), .A2(n14919), .ZN(n11213) );
  OAI22_X1 U13743 ( .A1(n14919), .A2(n11207), .B1(n12387), .B2(n13518), .ZN(
        n11211) );
  OAI211_X1 U13744 ( .C1(n11209), .C2(n11249), .A(n13523), .B(n11208), .ZN(
        n11248) );
  NOR2_X1 U13745 ( .A1(n11248), .A2(n14898), .ZN(n11210) );
  AOI211_X1 U13746 ( .C1(n14890), .C2(n12391), .A(n11211), .B(n11210), .ZN(
        n11212) );
  OAI211_X1 U13747 ( .C1(n11214), .C2(n14912), .A(n11213), .B(n11212), .ZN(
        P2_U3256) );
  XOR2_X1 U13748 ( .A(n11224), .B(n11215), .Z(n14944) );
  INV_X1 U13749 ( .A(n11216), .ZN(n14942) );
  INV_X1 U13750 ( .A(n14896), .ZN(n11219) );
  INV_X1 U13751 ( .A(n11217), .ZN(n11218) );
  OAI211_X1 U13752 ( .C1(n14942), .C2(n11219), .A(n11218), .B(n13523), .ZN(
        n14940) );
  NOR2_X1 U13753 ( .A1(n14940), .A2(n14898), .ZN(n11222) );
  OAI22_X1 U13754 ( .A1(n14942), .A2(n13472), .B1(n13518), .B2(n11220), .ZN(
        n11221) );
  AOI211_X1 U13755 ( .C1(n14944), .C2(n14900), .A(n11222), .B(n11221), .ZN(
        n11229) );
  XOR2_X1 U13756 ( .A(n11224), .B(n11223), .Z(n11226) );
  AOI21_X1 U13757 ( .B1(n11226), .B2(n14886), .A(n11225), .ZN(n14941) );
  MUX2_X1 U13758 ( .A(n11227), .B(n14941), .S(n14919), .Z(n11228) );
  NAND2_X1 U13759 ( .A1(n11229), .A2(n11228), .ZN(P2_U3258) );
  AND4_X1 U13760 ( .A1(n11233), .A2(n11232), .A3(n11231), .A4(n11230), .ZN(
        n11234) );
  AND2_X1 U13761 ( .A1(n11235), .A2(n11234), .ZN(n11255) );
  INV_X1 U13762 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n11247) );
  INV_X1 U13763 ( .A(n11237), .ZN(n11238) );
  NAND2_X1 U13764 ( .A1(n11238), .A2(n11421), .ZN(n14743) );
  NAND2_X1 U13765 ( .A1(n11239), .A2(n14759), .ZN(n11245) );
  INV_X1 U13766 ( .A(n11606), .ZN(n11240) );
  AOI21_X1 U13767 ( .B1(n11589), .B2(n14723), .A(n11240), .ZN(n11244) );
  NAND3_X1 U13768 ( .A1(n6470), .A2(n11241), .A3(n14618), .ZN(n11243) );
  NAND4_X1 U13769 ( .A1(n11245), .A2(n11244), .A3(n11243), .A4(n11242), .ZN(
        n11256) );
  NAND2_X1 U13770 ( .A1(n11256), .A2(n14761), .ZN(n11246) );
  OAI21_X1 U13771 ( .B1(n14761), .B2(n11247), .A(n11246), .ZN(P1_U3483) );
  OAI21_X1 U13772 ( .B1(n11249), .B2(n14958), .A(n11248), .ZN(n11251) );
  AOI211_X1 U13773 ( .C1(n14950), .C2(n11252), .A(n11251), .B(n11250), .ZN(
        n11323) );
  NAND2_X1 U13774 ( .A1(n14969), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n11253) );
  OAI21_X1 U13775 ( .B1(n11323), .B2(n14969), .A(n11253), .ZN(P2_U3508) );
  NAND2_X1 U13776 ( .A1(n11256), .A2(n14776), .ZN(n11257) );
  OAI21_X1 U13777 ( .B1(n14776), .B2(n10127), .A(n11257), .ZN(P1_U3536) );
  INV_X1 U13778 ( .A(n11258), .ZN(n11259) );
  AOI22_X1 U13779 ( .A1(n13531), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n11259), 
        .B2(n14905), .ZN(n11260) );
  OAI21_X1 U13780 ( .B1(n6938), .B2(n13472), .A(n11260), .ZN(n11263) );
  NOR2_X1 U13781 ( .A1(n11261), .A2(n13528), .ZN(n11262) );
  AOI211_X1 U13782 ( .C1(n11264), .C2(n14916), .A(n11263), .B(n11262), .ZN(
        n11265) );
  OAI21_X1 U13783 ( .B1(n14903), .B2(n11266), .A(n11265), .ZN(P2_U3255) );
  XNOR2_X1 U13784 ( .A(n11267), .B(n11270), .ZN(n11269) );
  AOI21_X1 U13785 ( .B1(n11269), .B2(n14886), .A(n11268), .ZN(n14957) );
  XNOR2_X1 U13786 ( .A(n11271), .B(n11270), .ZN(n14960) );
  NAND2_X1 U13787 ( .A1(n14955), .A2(n11272), .ZN(n11273) );
  NAND2_X1 U13788 ( .A1(n11273), .A2(n13523), .ZN(n11274) );
  OR2_X1 U13789 ( .A1(n11317), .A2(n11274), .ZN(n14956) );
  OAI22_X1 U13790 ( .A1(n14919), .A2(n11276), .B1(n11275), .B2(n13518), .ZN(
        n11277) );
  AOI21_X1 U13791 ( .B1(n14955), .B2(n14890), .A(n11277), .ZN(n11278) );
  OAI21_X1 U13792 ( .B1(n14956), .B2(n14898), .A(n11278), .ZN(n11279) );
  AOI21_X1 U13793 ( .B1(n14960), .B2(n14900), .A(n11279), .ZN(n11280) );
  OAI21_X1 U13794 ( .B1(n14903), .B2(n14957), .A(n11280), .ZN(P2_U3254) );
  OAI211_X1 U13795 ( .C1(n11283), .C2(n11282), .A(n11281), .B(n12642), .ZN(
        n11287) );
  NAND2_X1 U13796 ( .A1(n10675), .A2(n12669), .ZN(n11284) );
  NAND2_X1 U13797 ( .A1(P3_REG3_REG_7__SCAN_IN), .A2(P3_U3151), .ZN(n15041) );
  OAI211_X1 U13798 ( .C1(n12649), .C2(n6766), .A(n11284), .B(n15041), .ZN(
        n11285) );
  AOI21_X1 U13799 ( .B1(n12552), .B2(n12671), .A(n11285), .ZN(n11286) );
  OAI211_X1 U13800 ( .C1(n11415), .C2(n12645), .A(n11287), .B(n11286), .ZN(
        P3_U3153) );
  NOR2_X1 U13801 ( .A1(n11300), .A2(n11288), .ZN(n11290) );
  NOR2_X1 U13802 ( .A1(n11290), .A2(n11289), .ZN(n11295) );
  MUX2_X1 U13803 ( .A(n11291), .B(P1_REG1_REG_16__SCAN_IN), .S(n11616), .Z(
        n11294) );
  NAND2_X1 U13804 ( .A1(n11293), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n11292) );
  OAI211_X1 U13805 ( .C1(n11293), .C2(P1_REG1_REG_16__SCAN_IN), .A(n11295), 
        .B(n11292), .ZN(n11615) );
  OAI211_X1 U13806 ( .C1(n11295), .C2(n11294), .A(n11615), .B(n14603), .ZN(
        n11308) );
  NAND2_X1 U13807 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n13713)
         );
  NAND2_X1 U13808 ( .A1(n11616), .A2(n11297), .ZN(n11296) );
  OAI21_X1 U13809 ( .B1(n11616), .B2(n11297), .A(n11296), .ZN(n11298) );
  INV_X1 U13810 ( .A(n11298), .ZN(n11304) );
  NOR2_X1 U13811 ( .A1(n11300), .A2(n11299), .ZN(n11302) );
  NOR2_X1 U13812 ( .A1(n11302), .A2(n11301), .ZN(n11303) );
  NAND2_X1 U13813 ( .A1(n11303), .A2(n11304), .ZN(n11612) );
  OAI211_X1 U13814 ( .C1(n11304), .C2(n11303), .A(n14606), .B(n11612), .ZN(
        n11305) );
  NAND2_X1 U13815 ( .A1(n13713), .A2(n11305), .ZN(n11306) );
  AOI21_X1 U13816 ( .B1(n14587), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n11306), 
        .ZN(n11307) );
  OAI211_X1 U13817 ( .C1(n14611), .C2(n11616), .A(n11308), .B(n11307), .ZN(
        P1_U3259) );
  NAND2_X1 U13818 ( .A1(n11309), .A2(n13070), .ZN(n11310) );
  OAI211_X1 U13819 ( .C1(n11311), .C2(n13078), .A(n11310), .B(n12383), .ZN(
        P3_U3272) );
  XNOR2_X1 U13820 ( .A(n11312), .B(n11315), .ZN(n11314) );
  OAI22_X1 U13821 ( .A1(n11313), .A2(n14420), .B1(n14421), .B2(n14422), .ZN(
        n11349) );
  AOI21_X1 U13822 ( .B1(n11314), .B2(n14886), .A(n11349), .ZN(n14463) );
  XNOR2_X1 U13823 ( .A(n11316), .B(n11315), .ZN(n14466) );
  OAI211_X1 U13824 ( .C1(n14464), .C2(n11317), .A(n13523), .B(n6495), .ZN(
        n14462) );
  OAI22_X1 U13825 ( .A1(n14919), .A2(n11318), .B1(n11351), .B2(n13518), .ZN(
        n11319) );
  AOI21_X1 U13826 ( .B1(n11353), .B2(n14890), .A(n11319), .ZN(n11320) );
  OAI21_X1 U13827 ( .B1(n14462), .B2(n14898), .A(n11320), .ZN(n11321) );
  AOI21_X1 U13828 ( .B1(n14466), .B2(n14900), .A(n11321), .ZN(n11322) );
  OAI21_X1 U13829 ( .B1(n13531), .B2(n14463), .A(n11322), .ZN(P2_U3253) );
  INV_X1 U13830 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11325) );
  OR2_X1 U13831 ( .A1(n11323), .A2(n14962), .ZN(n11324) );
  OAI21_X1 U13832 ( .B1(n14964), .B2(n11325), .A(n11324), .ZN(P2_U3457) );
  XNOR2_X1 U13833 ( .A(n11327), .B(n11326), .ZN(n15156) );
  XNOR2_X1 U13834 ( .A(n11328), .B(n12252), .ZN(n11332) );
  OAI22_X1 U13835 ( .A1(n11330), .A2(n12927), .B1(n11329), .B2(n12925), .ZN(
        n11331) );
  AOI21_X1 U13836 ( .B1(n11332), .B2(n15106), .A(n11331), .ZN(n11333) );
  OAI21_X1 U13837 ( .B1(n15110), .B2(n15156), .A(n11333), .ZN(n15158) );
  NAND2_X1 U13838 ( .A1(n15158), .A2(n15117), .ZN(n11336) );
  OAI22_X1 U13839 ( .A1(n12933), .A2(n15155), .B1(n6624), .B2(n15112), .ZN(
        n11334) );
  AOI21_X1 U13840 ( .B1(n15119), .B2(P3_REG2_REG_8__SCAN_IN), .A(n11334), .ZN(
        n11335) );
  OAI211_X1 U13841 ( .C1(n15156), .C2(n15114), .A(n11336), .B(n11335), .ZN(
        P3_U3225) );
  XNOR2_X1 U13842 ( .A(n11353), .B(n13134), .ZN(n11337) );
  NAND2_X1 U13843 ( .A1(n13258), .A2(n13105), .ZN(n11338) );
  NAND2_X1 U13844 ( .A1(n11337), .A2(n11338), .ZN(n11364) );
  INV_X1 U13845 ( .A(n11337), .ZN(n11340) );
  INV_X1 U13846 ( .A(n11338), .ZN(n11339) );
  NAND2_X1 U13847 ( .A1(n11340), .A2(n11339), .ZN(n11341) );
  NAND2_X1 U13848 ( .A1(n11364), .A2(n11341), .ZN(n11348) );
  INV_X1 U13849 ( .A(n11365), .ZN(n11346) );
  AOI21_X1 U13850 ( .B1(n11348), .B2(n11347), .A(n11346), .ZN(n11355) );
  AOI22_X1 U13851 ( .A1(n14430), .A2(n11349), .B1(P2_REG3_REG_12__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11350) );
  OAI21_X1 U13852 ( .B1(n11351), .B2(n14789), .A(n11350), .ZN(n11352) );
  AOI21_X1 U13853 ( .B1(n11353), .B2(n14787), .A(n11352), .ZN(n11354) );
  OAI21_X1 U13854 ( .B1(n11355), .B2(n14782), .A(n11354), .ZN(P2_U3196) );
  OAI211_X1 U13855 ( .C1(n11358), .C2(n11357), .A(n11356), .B(n12642), .ZN(
        n11363) );
  NAND2_X1 U13856 ( .A1(n10675), .A2(n12668), .ZN(n11360) );
  OAI211_X1 U13857 ( .C1(n15155), .C2(n12649), .A(n11360), .B(n11359), .ZN(
        n11361) );
  AOI21_X1 U13858 ( .B1(n12552), .B2(n12670), .A(n11361), .ZN(n11362) );
  OAI211_X1 U13859 ( .C1(n6624), .C2(n12645), .A(n11363), .B(n11362), .ZN(
        P3_U3161) );
  XNOR2_X1 U13860 ( .A(n14456), .B(n13134), .ZN(n11728) );
  NAND2_X1 U13861 ( .A1(n13257), .A2(n13105), .ZN(n11727) );
  XNOR2_X1 U13862 ( .A(n11728), .B(n11727), .ZN(n11730) );
  XNOR2_X1 U13863 ( .A(n11731), .B(n11730), .ZN(n11372) );
  NOR2_X1 U13864 ( .A1(n14789), .A2(n11474), .ZN(n11370) );
  NAND2_X1 U13865 ( .A1(n13256), .A2(n13233), .ZN(n11367) );
  NAND2_X1 U13866 ( .A1(n13258), .A2(n13231), .ZN(n11366) );
  AND2_X1 U13867 ( .A1(n11367), .A2(n11366), .ZN(n11469) );
  OAI22_X1 U13868 ( .A1(n14779), .A2(n11469), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11368), .ZN(n11369) );
  AOI211_X1 U13869 ( .C1(n14456), .C2(n14787), .A(n11370), .B(n11369), .ZN(
        n11371) );
  OAI21_X1 U13870 ( .B1(n11372), .B2(n14782), .A(n11371), .ZN(P2_U3206) );
  MUX2_X1 U13871 ( .A(n11388), .B(P3_REG2_REG_10__SCAN_IN), .S(n11390), .Z(
        n15071) );
  NAND2_X1 U13872 ( .A1(n11390), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n11375) );
  AOI21_X1 U13873 ( .B1(n11395), .B2(n11376), .A(n11550), .ZN(n11404) );
  INV_X1 U13874 ( .A(n11390), .ZN(n15081) );
  NAND2_X1 U13875 ( .A1(n15053), .A2(n11378), .ZN(n11379) );
  NAND2_X1 U13876 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n15059), .ZN(n15058) );
  NAND2_X1 U13877 ( .A1(n11379), .A2(n15058), .ZN(n15067) );
  MUX2_X1 U13878 ( .A(P3_REG1_REG_10__SCAN_IN), .B(n11387), .S(n11390), .Z(
        n15066) );
  NAND2_X1 U13879 ( .A1(n15067), .A2(n15066), .ZN(n15065) );
  OAI21_X1 U13880 ( .B1(n15081), .B2(n11387), .A(n15065), .ZN(n11555) );
  XNOR2_X1 U13881 ( .A(n11555), .B(n11565), .ZN(n11380) );
  NAND2_X1 U13882 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n11380), .ZN(n11557) );
  OAI21_X1 U13883 ( .B1(n11380), .B2(P3_REG1_REG_11__SCAN_IN), .A(n11557), 
        .ZN(n11402) );
  INV_X1 U13884 ( .A(n11381), .ZN(n11382) );
  AOI22_X1 U13885 ( .A1(n11385), .A2(n11384), .B1(n11383), .B2(n11382), .ZN(
        n15050) );
  NOR2_X1 U13886 ( .A1(n11386), .A2(n6837), .ZN(n15048) );
  NOR2_X1 U13887 ( .A1(n15050), .A2(n15048), .ZN(n15075) );
  AND2_X1 U13888 ( .A1(n11386), .A2(n6837), .ZN(n15074) );
  NAND2_X1 U13889 ( .A1(n11389), .A2(n15081), .ZN(n11393) );
  INV_X1 U13890 ( .A(n11389), .ZN(n11391) );
  NAND2_X1 U13891 ( .A1(n11391), .A2(n11390), .ZN(n11392) );
  AND2_X1 U13892 ( .A1(n11393), .A2(n11392), .ZN(n15073) );
  NAND2_X1 U13893 ( .A1(n15077), .A2(n11393), .ZN(n11397) );
  XNOR2_X1 U13894 ( .A(n11566), .B(n11556), .ZN(n11396) );
  NAND2_X1 U13895 ( .A1(n11397), .A2(n11396), .ZN(n11569) );
  OAI21_X1 U13896 ( .B1(n11397), .B2(n11396), .A(n11569), .ZN(n11398) );
  NAND2_X1 U13897 ( .A1(n11398), .A2(n15078), .ZN(n11400) );
  AOI22_X1 U13898 ( .A1(n15068), .A2(P3_ADDR_REG_11__SCAN_IN), .B1(P3_U3151), 
        .B2(P3_REG3_REG_11__SCAN_IN), .ZN(n11399) );
  OAI211_X1 U13899 ( .C1(n15052), .C2(n11556), .A(n11400), .B(n11399), .ZN(
        n11401) );
  AOI21_X1 U13900 ( .B1(n15069), .B2(n11402), .A(n11401), .ZN(n11403) );
  OAI21_X1 U13901 ( .B1(n11404), .B2(n15063), .A(n11403), .ZN(P3_U3193) );
  OAI21_X1 U13902 ( .B1(n11406), .B2(n12246), .A(n11405), .ZN(n15151) );
  INV_X1 U13903 ( .A(n15151), .ZN(n11419) );
  INV_X1 U13904 ( .A(n12671), .ZN(n11408) );
  INV_X1 U13905 ( .A(n12669), .ZN(n11407) );
  OAI22_X1 U13906 ( .A1(n11408), .A2(n12927), .B1(n11407), .B2(n12925), .ZN(
        n11413) );
  XNOR2_X1 U13907 ( .A(n11410), .B(n11409), .ZN(n11411) );
  NOR2_X1 U13908 ( .A1(n11411), .A2(n12922), .ZN(n11412) );
  AOI211_X1 U13909 ( .C1(n12815), .C2(n15151), .A(n11413), .B(n11412), .ZN(
        n15153) );
  MUX2_X1 U13910 ( .A(n11414), .B(n15153), .S(n15117), .Z(n11418) );
  INV_X1 U13911 ( .A(n11415), .ZN(n11416) );
  AOI22_X1 U13912 ( .A1(n14402), .A2(n15149), .B1(n14400), .B2(n11416), .ZN(
        n11417) );
  OAI211_X1 U13913 ( .C1(n11419), .C2(n15114), .A(n11418), .B(n11417), .ZN(
        P3_U3226) );
  OAI222_X1 U13914 ( .A1(n14214), .A2(n11437), .B1(P1_U3086), .B2(n11421), 
        .C1(n11420), .C2(n12044), .ZN(P1_U3335) );
  XNOR2_X1 U13915 ( .A(n11422), .B(n11423), .ZN(n14744) );
  OAI21_X1 U13916 ( .B1(n11424), .B2(n11423), .A(n14617), .ZN(n11426) );
  OAI22_X1 U13917 ( .A1(n11425), .A2(n14053), .B1(n11751), .B2(n14055), .ZN(
        n11683) );
  AOI21_X1 U13918 ( .B1(n11426), .B2(n14618), .A(n11683), .ZN(n14746) );
  INV_X1 U13919 ( .A(n14746), .ZN(n11434) );
  NAND2_X1 U13920 ( .A1(n11427), .A2(n11674), .ZN(n11428) );
  NAND2_X1 U13921 ( .A1(n11428), .A2(n14679), .ZN(n11429) );
  OR2_X1 U13922 ( .A1(n11429), .A2(n14629), .ZN(n14745) );
  OAI22_X1 U13923 ( .A1(n14665), .A2(n11430), .B1(n11680), .B2(n14673), .ZN(
        n11431) );
  AOI21_X1 U13924 ( .B1(n11674), .B2(n14677), .A(n11431), .ZN(n11432) );
  OAI21_X1 U13925 ( .B1(n14745), .B2(n14065), .A(n11432), .ZN(n11433) );
  AOI21_X1 U13926 ( .B1(n11434), .B2(n14665), .A(n11433), .ZN(n11435) );
  OAI21_X1 U13927 ( .B1(n14083), .B2(n14744), .A(n11435), .ZN(P1_U3284) );
  OAI222_X1 U13928 ( .A1(P2_U3088), .A2(n6473), .B1(n13643), .B2(n11437), .C1(
        n11436), .C2(n13652), .ZN(P2_U3307) );
  XNOR2_X1 U13929 ( .A(n11438), .B(n8616), .ZN(n15160) );
  OAI211_X1 U13930 ( .C1(n11440), .C2(n8616), .A(n15106), .B(n11439), .ZN(
        n11442) );
  AOI22_X1 U13931 ( .A1(n15103), .A2(n12669), .B1(n12667), .B2(n15104), .ZN(
        n11441) );
  OAI211_X1 U13932 ( .C1(n15110), .C2(n15160), .A(n11442), .B(n11441), .ZN(
        n15162) );
  NAND2_X1 U13933 ( .A1(n15162), .A2(n15117), .ZN(n11445) );
  OAI22_X1 U13934 ( .A1(n12933), .A2(n15161), .B1(n11519), .B2(n15112), .ZN(
        n11443) );
  AOI21_X1 U13935 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n15119), .A(n11443), .ZN(
        n11444) );
  OAI211_X1 U13936 ( .C1(n15160), .C2(n15114), .A(n11445), .B(n11444), .ZN(
        P3_U3224) );
  NAND2_X1 U13937 ( .A1(n11447), .A2(n11446), .ZN(n11449) );
  NAND2_X1 U13938 ( .A1(n11449), .A2(n11448), .ZN(n11450) );
  NAND2_X1 U13939 ( .A1(n14872), .A2(n11450), .ZN(n11451) );
  XOR2_X1 U13940 ( .A(n14872), .B(n11450), .Z(n14876) );
  NAND2_X1 U13941 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n14876), .ZN(n14874) );
  NAND2_X1 U13942 ( .A1(n11451), .A2(n14874), .ZN(n11453) );
  MUX2_X1 U13943 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n13520), .S(n11528), .Z(
        n11452) );
  NAND2_X1 U13944 ( .A1(n11453), .A2(n11452), .ZN(n11524) );
  OAI211_X1 U13945 ( .C1(n11453), .C2(n11452), .A(n11524), .B(n14875), .ZN(
        n11465) );
  NAND2_X1 U13946 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n13178)
         );
  INV_X1 U13947 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n11454) );
  XNOR2_X1 U13948 ( .A(n11528), .B(n11454), .ZN(n11529) );
  INV_X1 U13949 ( .A(n11455), .ZN(n11456) );
  OAI21_X1 U13950 ( .B1(n14455), .B2(n11457), .A(n11456), .ZN(n11459) );
  NAND2_X1 U13951 ( .A1(n14872), .A2(n11459), .ZN(n11460) );
  XNOR2_X1 U13952 ( .A(n11459), .B(n11458), .ZN(n14879) );
  NAND2_X1 U13953 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n14879), .ZN(n14877) );
  NAND2_X1 U13954 ( .A1(n11460), .A2(n14877), .ZN(n11530) );
  XOR2_X1 U13955 ( .A(n11529), .B(n11530), .Z(n11461) );
  NAND2_X1 U13956 ( .A1(n14878), .A2(n11461), .ZN(n11462) );
  NAND2_X1 U13957 ( .A1(n13178), .A2(n11462), .ZN(n11463) );
  AOI21_X1 U13958 ( .B1(n14871), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n11463), 
        .ZN(n11464) );
  OAI211_X1 U13959 ( .C1(n14822), .C2(n11525), .A(n11465), .B(n11464), .ZN(
        P2_U3230) );
  INV_X1 U13960 ( .A(n11472), .ZN(n11466) );
  XNOR2_X1 U13961 ( .A(n11467), .B(n11466), .ZN(n11468) );
  NAND2_X1 U13962 ( .A1(n11468), .A2(n14886), .ZN(n11470) );
  NAND2_X1 U13963 ( .A1(n11470), .A2(n11469), .ZN(n14460) );
  INV_X1 U13964 ( .A(n14460), .ZN(n11480) );
  XOR2_X1 U13965 ( .A(n11472), .B(n11471), .Z(n14461) );
  AOI21_X1 U13966 ( .B1(n6495), .B2(n14456), .A(n13489), .ZN(n11473) );
  NAND2_X1 U13967 ( .A1(n11473), .A2(n14442), .ZN(n14457) );
  OAI22_X1 U13968 ( .A1(n14919), .A2(n11475), .B1(n11474), .B2(n13518), .ZN(
        n11476) );
  AOI21_X1 U13969 ( .B1(n14456), .B2(n14890), .A(n11476), .ZN(n11477) );
  OAI21_X1 U13970 ( .B1(n14457), .B2(n14898), .A(n11477), .ZN(n11478) );
  AOI21_X1 U13971 ( .B1(n14461), .B2(n14900), .A(n11478), .ZN(n11479) );
  OAI21_X1 U13972 ( .B1(n13531), .B2(n11480), .A(n11479), .ZN(P2_U3252) );
  INV_X1 U13973 ( .A(n11481), .ZN(n11482) );
  NAND2_X1 U13974 ( .A1(n13798), .A2(n11482), .ZN(n11484) );
  OAI211_X1 U13975 ( .C1(n11485), .C2(n13778), .A(n11484), .B(n11483), .ZN(
        n11511) );
  NAND2_X1 U13976 ( .A1(n11487), .A2(n11486), .ZN(n11489) );
  AOI22_X1 U13977 ( .A1(n13840), .A2(n12446), .B1(n12424), .B2(n13765), .ZN(
        n11490) );
  OAI22_X1 U13978 ( .A1(n13728), .A2(n12453), .B1(n14718), .B2(n12454), .ZN(
        n11488) );
  XNOR2_X1 U13979 ( .A(n11488), .B(n12444), .ZN(n13762) );
  NAND3_X1 U13980 ( .A1(n11491), .A2(n11490), .A3(n11489), .ZN(n13760) );
  OAI21_X1 U13981 ( .B1(n13759), .B2(n13762), .A(n13760), .ZN(n13723) );
  NAND2_X1 U13982 ( .A1(n12446), .A2(n13839), .ZN(n11493) );
  NAND2_X1 U13983 ( .A1(n14724), .A2(n12424), .ZN(n11492) );
  NAND2_X1 U13984 ( .A1(n11493), .A2(n11492), .ZN(n11502) );
  OAI22_X1 U13985 ( .A1(n11495), .A2(n12453), .B1(n11494), .B2(n12454), .ZN(
        n11496) );
  XNOR2_X1 U13986 ( .A(n11496), .B(n12444), .ZN(n11501) );
  XOR2_X1 U13987 ( .A(n11502), .B(n11501), .Z(n13724) );
  OAI22_X1 U13988 ( .A1(n14732), .A2(n12453), .B1(n11497), .B2(n12452), .ZN(
        n11592) );
  NAND2_X1 U13989 ( .A1(n11512), .A2(n12441), .ZN(n11499) );
  NAND2_X1 U13990 ( .A1(n13838), .A2(n12424), .ZN(n11498) );
  NAND2_X1 U13991 ( .A1(n11499), .A2(n11498), .ZN(n11500) );
  XNOR2_X1 U13992 ( .A(n11500), .B(n12444), .ZN(n11591) );
  XOR2_X1 U13993 ( .A(n11591), .B(n11592), .Z(n11506) );
  INV_X1 U13994 ( .A(n11501), .ZN(n11504) );
  INV_X1 U13995 ( .A(n11502), .ZN(n11503) );
  NAND2_X1 U13996 ( .A1(n11504), .A2(n11503), .ZN(n11507) );
  INV_X1 U13997 ( .A(n11594), .ZN(n11509) );
  AOI21_X1 U13998 ( .B1(n13722), .B2(n11507), .A(n11506), .ZN(n11508) );
  NOR3_X1 U13999 ( .A1(n11509), .A2(n11508), .A3(n13817), .ZN(n11510) );
  AOI211_X1 U14000 ( .C1(n11512), .C2(n13815), .A(n11511), .B(n11510), .ZN(
        n11513) );
  INV_X1 U14001 ( .A(n11513), .ZN(P1_U3239) );
  AOI21_X1 U14002 ( .B1(n11515), .B2(n11514), .A(n6643), .ZN(n11523) );
  INV_X1 U14003 ( .A(n12667), .ZN(n11518) );
  AOI22_X1 U14004 ( .A1(n12634), .A2(n11516), .B1(P3_REG3_REG_9__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11517) );
  OAI21_X1 U14005 ( .B1(n12608), .B2(n11518), .A(n11517), .ZN(n11521) );
  NOR2_X1 U14006 ( .A1(n12645), .A2(n11519), .ZN(n11520) );
  AOI211_X1 U14007 ( .C1(n12552), .C2(n12669), .A(n11521), .B(n11520), .ZN(
        n11522) );
  OAI21_X1 U14008 ( .B1(n11523), .B2(n12637), .A(n11522), .ZN(P3_U3171) );
  OAI21_X1 U14009 ( .B1(n13520), .B2(n11525), .A(n11524), .ZN(n11527) );
  AOI22_X1 U14010 ( .A1(n11624), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13503), 
        .B2(n11632), .ZN(n11526) );
  NAND2_X1 U14011 ( .A1(n11526), .A2(n11527), .ZN(n11625) );
  OAI211_X1 U14012 ( .C1(n11527), .C2(n11526), .A(n14875), .B(n11625), .ZN(
        n11535) );
  NAND2_X1 U14013 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n13187)
         );
  AOI22_X1 U14014 ( .A1(n11530), .A2(n11529), .B1(P2_REG1_REG_16__SCAN_IN), 
        .B2(n11528), .ZN(n11635) );
  XNOR2_X1 U14015 ( .A(n11624), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n11634) );
  XOR2_X1 U14016 ( .A(n11635), .B(n11634), .Z(n11531) );
  NAND2_X1 U14017 ( .A1(n14878), .A2(n11531), .ZN(n11532) );
  NAND2_X1 U14018 ( .A1(n13187), .A2(n11532), .ZN(n11533) );
  AOI21_X1 U14019 ( .B1(n14871), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n11533), 
        .ZN(n11534) );
  OAI211_X1 U14020 ( .C1(n14822), .C2(n11632), .A(n11535), .B(n11534), .ZN(
        P2_U3231) );
  XNOR2_X1 U14021 ( .A(n11536), .B(n12171), .ZN(n15170) );
  AOI22_X1 U14022 ( .A1(n12666), .A2(n15104), .B1(n15103), .B2(n12668), .ZN(
        n11540) );
  OAI211_X1 U14023 ( .C1(n11538), .C2(n12171), .A(n11537), .B(n15106), .ZN(
        n11539) );
  OAI211_X1 U14024 ( .C1(n15170), .C2(n15110), .A(n11540), .B(n11539), .ZN(
        n15172) );
  NAND2_X1 U14025 ( .A1(n15172), .A2(n15117), .ZN(n11543) );
  OAI22_X1 U14026 ( .A1(n12933), .A2(n15167), .B1(n11588), .B2(n15112), .ZN(
        n11541) );
  AOI21_X1 U14027 ( .B1(n15119), .B2(P3_REG2_REG_10__SCAN_IN), .A(n11541), 
        .ZN(n11542) );
  OAI211_X1 U14028 ( .C1(n15170), .C2(n15114), .A(n11543), .B(n11542), .ZN(
        P3_U3223) );
  OAI222_X1 U14029 ( .A1(n14208), .A2(n11547), .B1(P1_U3086), .B2(n11545), 
        .C1(n11544), .C2(n12044), .ZN(P1_U3334) );
  OAI222_X1 U14030 ( .A1(P2_U3088), .A2(n11548), .B1(n13643), .B2(n11547), 
        .C1(n11546), .C2(n13652), .ZN(P2_U3306) );
  NOR2_X1 U14031 ( .A1(n11565), .A2(n11549), .ZN(n11551) );
  MUX2_X1 U14032 ( .A(P3_REG2_REG_12__SCAN_IN), .B(n11767), .S(n11791), .Z(
        n11553) );
  INV_X1 U14033 ( .A(n11788), .ZN(n11552) );
  AOI21_X1 U14034 ( .B1(n11554), .B2(n11553), .A(n11552), .ZN(n11576) );
  NAND2_X1 U14035 ( .A1(n11556), .A2(n11555), .ZN(n11558) );
  MUX2_X1 U14036 ( .A(n11559), .B(P3_REG1_REG_12__SCAN_IN), .S(n11791), .Z(
        n11560) );
  OAI21_X1 U14037 ( .B1(n11561), .B2(n11560), .A(n11790), .ZN(n11574) );
  INV_X1 U14038 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11562) );
  NOR2_X1 U14039 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11562), .ZN(n11563) );
  AOI21_X1 U14040 ( .B1(n15068), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n11563), 
        .ZN(n11564) );
  OAI21_X1 U14041 ( .B1(n15052), .B2(n11793), .A(n11564), .ZN(n11573) );
  NAND2_X1 U14042 ( .A1(n11566), .A2(n11565), .ZN(n11568) );
  XNOR2_X1 U14043 ( .A(n11794), .B(n11791), .ZN(n11567) );
  NAND3_X1 U14044 ( .A1(n11569), .A2(n11568), .A3(n11567), .ZN(n11797) );
  INV_X1 U14045 ( .A(n11797), .ZN(n11571) );
  AOI21_X1 U14046 ( .B1(n11569), .B2(n11568), .A(n11567), .ZN(n11570) );
  NOR3_X1 U14047 ( .A1(n11571), .A2(n11570), .A3(n15054), .ZN(n11572) );
  AOI211_X1 U14048 ( .C1(n15069), .C2(n11574), .A(n11573), .B(n11572), .ZN(
        n11575) );
  OAI21_X1 U14049 ( .B1(n11576), .B2(n15063), .A(n11575), .ZN(P3_U3194) );
  INV_X1 U14050 ( .A(n11577), .ZN(n11578) );
  INV_X1 U14051 ( .A(SI_24_), .ZN(n15287) );
  OAI222_X1 U14052 ( .A1(P3_U3151), .A2(n8921), .B1(n13076), .B2(n11578), .C1(
        n15287), .C2(n13078), .ZN(P3_U3271) );
  AOI21_X1 U14053 ( .B1(n11580), .B2(n11579), .A(n12637), .ZN(n11582) );
  NAND2_X1 U14054 ( .A1(n11582), .A2(n11581), .ZN(n11587) );
  AOI22_X1 U14055 ( .A1(n12634), .A2(n11583), .B1(P3_REG3_REG_10__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11584) );
  OAI21_X1 U14056 ( .B1(n12608), .B2(n11834), .A(n11584), .ZN(n11585) );
  AOI21_X1 U14057 ( .B1(n12552), .B2(n12668), .A(n11585), .ZN(n11586) );
  OAI211_X1 U14058 ( .C1(n11588), .C2(n12645), .A(n11587), .B(n11586), .ZN(
        P3_U3157) );
  AOI22_X1 U14059 ( .A1(n11589), .A2(n12424), .B1(n12446), .B2(n13836), .ZN(
        n11668) );
  AOI22_X1 U14060 ( .A1(n11589), .A2(n12441), .B1(n12424), .B2(n13836), .ZN(
        n11590) );
  XNOR2_X1 U14061 ( .A(n11590), .B(n12444), .ZN(n11669) );
  XOR2_X1 U14062 ( .A(n11668), .B(n11669), .Z(n11602) );
  AND2_X1 U14063 ( .A1(n12446), .A2(n13837), .ZN(n11595) );
  AOI21_X1 U14064 ( .B1(n14647), .B2(n12424), .A(n11595), .ZN(n11597) );
  AOI22_X1 U14065 ( .A1(n14647), .A2(n12441), .B1(n12424), .B2(n13837), .ZN(
        n11596) );
  XNOR2_X1 U14066 ( .A(n11596), .B(n12444), .ZN(n11598) );
  XOR2_X1 U14067 ( .A(n11597), .B(n11598), .Z(n11644) );
  INV_X1 U14068 ( .A(n11597), .ZN(n11600) );
  INV_X1 U14069 ( .A(n11598), .ZN(n11599) );
  OAI21_X1 U14070 ( .B1(n11602), .B2(n11601), .A(n11677), .ZN(n11603) );
  NAND2_X1 U14071 ( .A1(n11603), .A2(n13795), .ZN(n11610) );
  INV_X1 U14072 ( .A(n11604), .ZN(n11608) );
  OAI21_X1 U14073 ( .B1(n11606), .B2(n13778), .A(n11605), .ZN(n11607) );
  AOI21_X1 U14074 ( .B1(n11608), .B2(n13798), .A(n11607), .ZN(n11609) );
  OAI211_X1 U14075 ( .C1(n10005), .C2(n13803), .A(n11610), .B(n11609), .ZN(
        P1_U3221) );
  OR2_X1 U14076 ( .A1(n11614), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n11611) );
  NAND2_X1 U14077 ( .A1(n11614), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n13915) );
  NAND2_X1 U14078 ( .A1(n11611), .A2(n13915), .ZN(n13911) );
  OAI21_X1 U14079 ( .B1(n11297), .B2(n11616), .A(n11612), .ZN(n13913) );
  XOR2_X1 U14080 ( .A(n13911), .B(n13913), .Z(n11623) );
  NAND2_X1 U14081 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13740)
         );
  NOR2_X1 U14082 ( .A1(n11614), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n11613) );
  AOI21_X1 U14083 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n11614), .A(n11613), 
        .ZN(n11618) );
  OAI21_X1 U14084 ( .B1(n11291), .B2(n11616), .A(n11615), .ZN(n11617) );
  NAND2_X1 U14085 ( .A1(n11617), .A2(n11618), .ZN(n13904) );
  OAI211_X1 U14086 ( .C1(n11618), .C2(n11617), .A(n14603), .B(n13904), .ZN(
        n11619) );
  NAND2_X1 U14087 ( .A1(n13740), .A2(n11619), .ZN(n11621) );
  NOR2_X1 U14088 ( .A1(n14611), .A2(n13905), .ZN(n11620) );
  AOI211_X1 U14089 ( .C1(n14587), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n11621), 
        .B(n11620), .ZN(n11622) );
  OAI21_X1 U14090 ( .B1(n11623), .B2(n13920), .A(n11622), .ZN(P1_U3260) );
  NAND2_X1 U14091 ( .A1(n11624), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n11626) );
  NAND2_X1 U14092 ( .A1(n11626), .A2(n11625), .ZN(n11627) );
  NOR2_X1 U14093 ( .A1(n11627), .A2(n13305), .ZN(n13302) );
  AOI21_X1 U14094 ( .B1(n11627), .B2(n13305), .A(n13302), .ZN(n11628) );
  INV_X1 U14095 ( .A(n11628), .ZN(n11629) );
  NOR2_X1 U14096 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n11629), .ZN(n13303) );
  AOI21_X1 U14097 ( .B1(n11629), .B2(P2_REG2_REG_18__SCAN_IN), .A(n13303), 
        .ZN(n11639) );
  INV_X1 U14098 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n11630) );
  NAND2_X1 U14099 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13220)
         );
  OAI21_X1 U14100 ( .B1(n14832), .B2(n11630), .A(n13220), .ZN(n11631) );
  AOI21_X1 U14101 ( .B1(n13305), .B2(n14873), .A(n11631), .ZN(n11638) );
  INV_X1 U14102 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n11633) );
  OAI22_X1 U14103 ( .A1(n11635), .A2(n11634), .B1(n11633), .B2(n11632), .ZN(
        n13306) );
  XOR2_X1 U14104 ( .A(n13305), .B(n13306), .Z(n11636) );
  NAND2_X1 U14105 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n11636), .ZN(n13308) );
  OAI211_X1 U14106 ( .C1(n11636), .C2(P2_REG1_REG_18__SCAN_IN), .A(n14878), 
        .B(n13308), .ZN(n11637) );
  OAI211_X1 U14107 ( .C1(n11639), .C2(n14856), .A(n11638), .B(n11637), .ZN(
        P2_U3232) );
  NAND2_X1 U14108 ( .A1(n13836), .A2(n14631), .ZN(n11641) );
  NAND2_X1 U14109 ( .A1(n13838), .A2(n14482), .ZN(n11640) );
  AND2_X1 U14110 ( .A1(n11641), .A2(n11640), .ZN(n14639) );
  INV_X1 U14111 ( .A(n11642), .ZN(n14642) );
  NAND2_X1 U14112 ( .A1(n13798), .A2(n14642), .ZN(n11643) );
  NAND2_X1 U14113 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n13887) );
  OAI211_X1 U14114 ( .C1(n14639), .C2(n13778), .A(n11643), .B(n13887), .ZN(
        n11648) );
  XNOR2_X1 U14115 ( .A(n11645), .B(n11644), .ZN(n11646) );
  NOR2_X1 U14116 ( .A1(n11646), .A2(n13817), .ZN(n11647) );
  AOI211_X1 U14117 ( .C1(n14647), .C2(n13815), .A(n11648), .B(n11647), .ZN(
        n11649) );
  INV_X1 U14118 ( .A(n11649), .ZN(P1_U3213) );
  XNOR2_X1 U14119 ( .A(n11650), .B(n11651), .ZN(n14528) );
  OAI21_X1 U14120 ( .B1(n11652), .B2(n14526), .A(n14679), .ZN(n11653) );
  OR2_X1 U14121 ( .A1(n11692), .A2(n11653), .ZN(n14524) );
  OAI22_X1 U14122 ( .A1(n14665), .A2(n11654), .B1(n11862), .B2(n14673), .ZN(
        n11655) );
  AOI21_X1 U14123 ( .B1(n11656), .B2(n14677), .A(n11655), .ZN(n11657) );
  OAI21_X1 U14124 ( .B1(n14524), .B2(n14065), .A(n11657), .ZN(n11666) );
  NOR2_X1 U14125 ( .A1(n11659), .A2(n7378), .ZN(n11660) );
  AOI21_X1 U14126 ( .B1(n14619), .B2(n11660), .A(n14690), .ZN(n11663) );
  NAND2_X1 U14127 ( .A1(n13834), .A2(n14482), .ZN(n11662) );
  NAND2_X1 U14128 ( .A1(n13833), .A2(n14631), .ZN(n11661) );
  NAND2_X1 U14129 ( .A1(n11662), .A2(n11661), .ZN(n11865) );
  AOI21_X1 U14130 ( .B1(n11664), .B2(n11663), .A(n11865), .ZN(n14525) );
  NOR2_X1 U14131 ( .A1(n14525), .A2(n14644), .ZN(n11665) );
  AOI211_X1 U14132 ( .C1(n14528), .C2(n14662), .A(n11666), .B(n11665), .ZN(
        n11667) );
  INV_X1 U14133 ( .A(n11667), .ZN(P1_U3282) );
  INV_X1 U14134 ( .A(n11674), .ZN(n14747) );
  NAND2_X1 U14135 ( .A1(n11669), .A2(n11668), .ZN(n11675) );
  AND2_X1 U14136 ( .A1(n11677), .A2(n11675), .ZN(n11679) );
  NAND2_X1 U14137 ( .A1(n11674), .A2(n12441), .ZN(n11671) );
  NAND2_X1 U14138 ( .A1(n13835), .A2(n12424), .ZN(n11670) );
  NAND2_X1 U14139 ( .A1(n11671), .A2(n11670), .ZN(n11672) );
  XNOR2_X1 U14140 ( .A(n11672), .B(n12444), .ZN(n11746) );
  AND2_X1 U14141 ( .A1(n12446), .A2(n13835), .ZN(n11673) );
  AOI21_X1 U14142 ( .B1(n11674), .B2(n12424), .A(n11673), .ZN(n11747) );
  XNOR2_X1 U14143 ( .A(n11746), .B(n11747), .ZN(n11678) );
  NAND2_X1 U14144 ( .A1(n11677), .A2(n11676), .ZN(n11750) );
  OAI211_X1 U14145 ( .C1(n11679), .C2(n11678), .A(n13795), .B(n11750), .ZN(
        n11685) );
  INV_X1 U14146 ( .A(n13798), .ZN(n13813) );
  NOR2_X1 U14147 ( .A1(n13813), .A2(n11680), .ZN(n11681) );
  AOI211_X1 U14148 ( .C1(n13769), .C2(n11683), .A(n11682), .B(n11681), .ZN(
        n11684) );
  OAI211_X1 U14149 ( .C1(n14747), .C2(n13803), .A(n11685), .B(n11684), .ZN(
        P1_U3231) );
  XNOR2_X1 U14150 ( .A(n11686), .B(n11688), .ZN(n14334) );
  OAI211_X1 U14151 ( .C1(n11689), .C2(n11688), .A(n11687), .B(n14618), .ZN(
        n11691) );
  AOI22_X1 U14152 ( .A1(n14482), .A2(n14630), .B1(n14483), .B2(n14631), .ZN(
        n11690) );
  AND2_X1 U14153 ( .A1(n11691), .A2(n11690), .ZN(n14336) );
  INV_X1 U14154 ( .A(n14336), .ZN(n11697) );
  OAI211_X1 U14155 ( .C1(n11692), .C2(n14337), .A(n14679), .B(n11809), .ZN(
        n14335) );
  OAI22_X1 U14156 ( .A1(n14665), .A2(n11693), .B1(n11907), .B2(n14673), .ZN(
        n11694) );
  AOI21_X1 U14157 ( .B1(n11900), .B2(n14677), .A(n11694), .ZN(n11695) );
  OAI21_X1 U14158 ( .B1(n14335), .B2(n14065), .A(n11695), .ZN(n11696) );
  AOI21_X1 U14159 ( .B1(n11697), .B2(n14665), .A(n11696), .ZN(n11698) );
  OAI21_X1 U14160 ( .B1(n14083), .B2(n14334), .A(n11698), .ZN(P1_U3281) );
  INV_X1 U14161 ( .A(n11699), .ZN(n11700) );
  AOI21_X1 U14162 ( .B1(n11708), .B2(n11701), .A(n11700), .ZN(n13615) );
  AOI21_X1 U14163 ( .B1(n14444), .B2(n13611), .A(n13489), .ZN(n11703) );
  AND2_X1 U14164 ( .A1(n11703), .A2(n13522), .ZN(n13610) );
  OAI22_X1 U14165 ( .A1(n9430), .A2(n13472), .B1(n11704), .B2(n14919), .ZN(
        n11705) );
  AOI21_X1 U14166 ( .B1(n13610), .B2(n14916), .A(n11705), .ZN(n11713) );
  OAI21_X1 U14167 ( .B1(n11708), .B2(n11707), .A(n11706), .ZN(n11710) );
  OAI22_X1 U14168 ( .A1(n13185), .A2(n14422), .B1(n11709), .B2(n14420), .ZN(
        n11740) );
  AOI21_X1 U14169 ( .B1(n11710), .B2(n14886), .A(n11740), .ZN(n13613) );
  OAI21_X1 U14170 ( .B1(n11742), .B2(n13518), .A(n13613), .ZN(n11711) );
  NAND2_X1 U14171 ( .A1(n11711), .A2(n14919), .ZN(n11712) );
  OAI211_X1 U14172 ( .C1(n13615), .C2(n13528), .A(n11713), .B(n11712), .ZN(
        P2_U3250) );
  XOR2_X1 U14173 ( .A(n11714), .B(n12272), .Z(n14397) );
  XNOR2_X1 U14174 ( .A(n11715), .B(n12272), .ZN(n11718) );
  NAND2_X1 U14175 ( .A1(n12665), .A2(n15104), .ZN(n11717) );
  NAND2_X1 U14176 ( .A1(n12667), .A2(n15103), .ZN(n11716) );
  NAND2_X1 U14177 ( .A1(n11717), .A2(n11716), .ZN(n11838) );
  AOI21_X1 U14178 ( .B1(n11718), .B2(n15106), .A(n11838), .ZN(n14396) );
  OAI21_X1 U14179 ( .B1(n14397), .B2(n12988), .A(n14396), .ZN(n11723) );
  INV_X1 U14180 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n11719) );
  OAI22_X1 U14181 ( .A1(n13059), .A2(n11836), .B1(n11719), .B2(n15175), .ZN(
        n11720) );
  AOI21_X1 U14182 ( .B1(n11723), .B2(n15175), .A(n11720), .ZN(n11721) );
  INV_X1 U14183 ( .A(n11721), .ZN(P3_U3423) );
  OAI22_X1 U14184 ( .A1(n13003), .A2(n11836), .B1(n15183), .B2(n11394), .ZN(
        n11722) );
  AOI21_X1 U14185 ( .B1(n11723), .B2(n15183), .A(n11722), .ZN(n11724) );
  INV_X1 U14186 ( .A(n11724), .ZN(P3_U3470) );
  INV_X1 U14187 ( .A(n11725), .ZN(n11726) );
  OAI222_X1 U14188 ( .A1(n13076), .A2(n11726), .B1(P3_U3151), .B2(n8916), .C1(
        n15304), .C2(n13078), .ZN(P3_U3270) );
  NAND2_X1 U14189 ( .A1(n13255), .A2(n13105), .ZN(n12501) );
  NAND2_X1 U14190 ( .A1(n14428), .A2(n12501), .ZN(n11739) );
  NAND2_X1 U14191 ( .A1(n13225), .A2(n13255), .ZN(n11738) );
  XNOR2_X1 U14192 ( .A(n14443), .B(n13134), .ZN(n11732) );
  NAND2_X1 U14193 ( .A1(n13256), .A2(n13105), .ZN(n11733) );
  NAND2_X1 U14194 ( .A1(n11732), .A2(n11733), .ZN(n11737) );
  INV_X1 U14195 ( .A(n11732), .ZN(n11735) );
  INV_X1 U14196 ( .A(n11733), .ZN(n11734) );
  NAND2_X1 U14197 ( .A1(n11735), .A2(n11734), .ZN(n11736) );
  NAND2_X1 U14198 ( .A1(n11737), .A2(n11736), .ZN(n14425) );
  XOR2_X1 U14199 ( .A(n6725), .B(n13611), .Z(n12500) );
  MUX2_X1 U14200 ( .A(n11739), .B(n11738), .S(n12502), .Z(n11745) );
  AOI22_X1 U14201 ( .A1(n14430), .A2(n11740), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11741) );
  OAI21_X1 U14202 ( .B1(n11742), .B2(n14789), .A(n11741), .ZN(n11743) );
  AOI21_X1 U14203 ( .B1(n13611), .B2(n14787), .A(n11743), .ZN(n11744) );
  NAND2_X1 U14204 ( .A1(n11745), .A2(n11744), .ZN(P2_U3213) );
  OAI22_X1 U14205 ( .A1(n14756), .A2(n12454), .B1(n11751), .B2(n12453), .ZN(
        n11752) );
  XNOR2_X1 U14206 ( .A(n11752), .B(n12444), .ZN(n11855) );
  AND2_X1 U14207 ( .A1(n12446), .A2(n13834), .ZN(n11753) );
  AOI21_X1 U14208 ( .B1(n14628), .B2(n12424), .A(n11753), .ZN(n11854) );
  XNOR2_X1 U14209 ( .A(n11855), .B(n11854), .ZN(n11857) );
  XNOR2_X1 U14210 ( .A(n11858), .B(n11857), .ZN(n11759) );
  NAND2_X1 U14211 ( .A1(n13835), .A2(n14482), .ZN(n14622) );
  NOR2_X1 U14212 ( .A1(n13778), .A2(n14622), .ZN(n11754) );
  AOI211_X1 U14213 ( .C1(n13810), .C2(n14630), .A(n11755), .B(n11754), .ZN(
        n11756) );
  OAI21_X1 U14214 ( .B1(n13813), .B2(n14624), .A(n11756), .ZN(n11757) );
  AOI21_X1 U14215 ( .B1(n14628), .B2(n13815), .A(n11757), .ZN(n11758) );
  OAI21_X1 U14216 ( .B1(n11759), .B2(n13817), .A(n11758), .ZN(P1_U3217) );
  XNOR2_X1 U14217 ( .A(n11760), .B(n12182), .ZN(n11761) );
  OAI222_X1 U14218 ( .A1(n12925), .A2(n11762), .B1(n12927), .B2(n11834), .C1(
        n11761), .C2(n12922), .ZN(n14412) );
  INV_X1 U14219 ( .A(n14412), .ZN(n11771) );
  OAI21_X1 U14220 ( .B1(n11765), .B2(n11764), .A(n11763), .ZN(n14414) );
  NAND2_X1 U14221 ( .A1(n15110), .A2(n11766), .ZN(n14395) );
  NAND2_X1 U14222 ( .A1(n15117), .A2(n14395), .ZN(n12902) );
  INV_X1 U14223 ( .A(n12281), .ZN(n14411) );
  NOR2_X1 U14224 ( .A1(n12933), .A2(n14411), .ZN(n11769) );
  OAI22_X1 U14225 ( .A1(n15117), .A2(n11767), .B1(n11888), .B2(n15112), .ZN(
        n11768) );
  AOI211_X1 U14226 ( .C1(n14414), .C2(n12935), .A(n11769), .B(n11768), .ZN(
        n11770) );
  OAI21_X1 U14227 ( .B1(n11771), .B2(n15119), .A(n11770), .ZN(P3_U3221) );
  INV_X1 U14228 ( .A(n11772), .ZN(n11775) );
  INV_X1 U14229 ( .A(n13652), .ZN(n13645) );
  AOI22_X1 U14230 ( .A1(n11773), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n13645), .ZN(n11774) );
  OAI21_X1 U14231 ( .B1(n11775), .B2(n13643), .A(n11774), .ZN(P2_U3305) );
  INV_X1 U14232 ( .A(n11776), .ZN(n11777) );
  OAI222_X1 U14233 ( .A1(n6671), .A2(P3_U3151), .B1(n13078), .B2(n15310), .C1(
        n13076), .C2(n11777), .ZN(P3_U3269) );
  OR2_X1 U14234 ( .A1(n12285), .A2(n6535), .ZN(n12183) );
  XNOR2_X1 U14235 ( .A(n11778), .B(n12183), .ZN(n11779) );
  NAND2_X1 U14236 ( .A1(n11779), .A2(n15106), .ZN(n11781) );
  AOI22_X1 U14237 ( .A1(n15104), .A2(n12663), .B1(n12665), .B2(n15103), .ZN(
        n11780) );
  NAND2_X1 U14238 ( .A1(n11781), .A2(n11780), .ZN(n14410) );
  INV_X1 U14239 ( .A(n14410), .ZN(n11786) );
  INV_X1 U14240 ( .A(n12183), .ZN(n12283) );
  XNOR2_X1 U14241 ( .A(n11782), .B(n12283), .ZN(n14406) );
  NOR2_X1 U14242 ( .A1(n14407), .A2(n12933), .ZN(n11784) );
  OAI22_X1 U14243 ( .A1(n15117), .A2(n8674), .B1(n11930), .B2(n15112), .ZN(
        n11783) );
  AOI211_X1 U14244 ( .C1(n14406), .C2(n12935), .A(n11784), .B(n11783), .ZN(
        n11785) );
  OAI21_X1 U14245 ( .B1(n11786), .B2(n15119), .A(n11785), .ZN(P3_U3220) );
  INV_X1 U14246 ( .A(n12680), .ZN(n12688) );
  NAND2_X1 U14247 ( .A1(n11793), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n11787) );
  AOI21_X1 U14248 ( .B1(n8674), .B2(n11789), .A(n12676), .ZN(n11806) );
  NAND2_X1 U14249 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n11792), .ZN(n12681) );
  OAI21_X1 U14250 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n11792), .A(n12681), 
        .ZN(n11804) );
  NAND2_X1 U14251 ( .A1(n11794), .A2(n11793), .ZN(n11796) );
  XNOR2_X1 U14252 ( .A(n12687), .B(n12688), .ZN(n11795) );
  NAND3_X1 U14253 ( .A1(n11797), .A2(n11796), .A3(n11795), .ZN(n12694) );
  INV_X1 U14254 ( .A(n12694), .ZN(n11799) );
  AOI21_X1 U14255 ( .B1(n11797), .B2(n11796), .A(n11795), .ZN(n11798) );
  OAI21_X1 U14256 ( .B1(n11799), .B2(n11798), .A(n15078), .ZN(n11802) );
  NOR2_X1 U14257 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11927), .ZN(n11800) );
  AOI21_X1 U14258 ( .B1(n15068), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n11800), 
        .ZN(n11801) );
  OAI211_X1 U14259 ( .C1(n15052), .C2(n12680), .A(n11802), .B(n11801), .ZN(
        n11803) );
  AOI21_X1 U14260 ( .B1(n15069), .B2(n11804), .A(n11803), .ZN(n11805) );
  OAI21_X1 U14261 ( .B1(n11806), .B2(n15063), .A(n11805), .ZN(P3_U3195) );
  XNOR2_X1 U14262 ( .A(n11807), .B(n11808), .ZN(n14523) );
  AOI21_X1 U14263 ( .B1(n11809), .B2(n14518), .A(n14699), .ZN(n11810) );
  NAND2_X1 U14264 ( .A1(n11810), .A2(n14481), .ZN(n14519) );
  OR2_X1 U14265 ( .A1(n13807), .A2(n14055), .ZN(n11812) );
  NAND2_X1 U14266 ( .A1(n13833), .A2(n14482), .ZN(n11811) );
  NAND2_X1 U14267 ( .A1(n11812), .A2(n11811), .ZN(n14517) );
  OAI22_X1 U14268 ( .A1(n14665), .A2(n11813), .B1(n11965), .B2(n14673), .ZN(
        n11814) );
  AOI21_X1 U14269 ( .B1(n14665), .B2(n14517), .A(n11814), .ZN(n11816) );
  NAND2_X1 U14270 ( .A1(n14518), .A2(n14677), .ZN(n11815) );
  OAI211_X1 U14271 ( .C1(n14519), .C2(n14065), .A(n11816), .B(n11815), .ZN(
        n11821) );
  OAI21_X1 U14272 ( .B1(n11819), .B2(n11818), .A(n11817), .ZN(n14521) );
  INV_X1 U14273 ( .A(n14035), .ZN(n14068) );
  NOR2_X1 U14274 ( .A1(n14521), .A2(n14068), .ZN(n11820) );
  AOI211_X1 U14275 ( .C1(n14523), .C2(n14662), .A(n11821), .B(n11820), .ZN(
        n11822) );
  INV_X1 U14276 ( .A(n11822), .ZN(P1_U3280) );
  INV_X1 U14277 ( .A(n11827), .ZN(n11825) );
  NAND2_X1 U14278 ( .A1(n13645), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n11823) );
  OAI211_X1 U14279 ( .C1(n11825), .C2(n13643), .A(n11824), .B(n11823), .ZN(
        P2_U3304) );
  NAND2_X1 U14280 ( .A1(n11827), .A2(n11826), .ZN(n11829) );
  OAI211_X1 U14281 ( .C1(n11830), .C2(n12044), .A(n11829), .B(n11828), .ZN(
        P1_U3332) );
  INV_X1 U14282 ( .A(n11831), .ZN(n11832) );
  NAND2_X1 U14283 ( .A1(n6513), .A2(n11833), .ZN(n11835) );
  XNOR2_X1 U14284 ( .A(n11835), .B(n11834), .ZN(n11842) );
  INV_X1 U14285 ( .A(n11836), .ZN(n14403) );
  INV_X1 U14286 ( .A(n11837), .ZN(n12647) );
  AOI22_X1 U14287 ( .A1(n12647), .A2(n11838), .B1(P3_REG3_REG_11__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11839) );
  OAI21_X1 U14288 ( .B1(n12645), .B2(n14399), .A(n11839), .ZN(n11840) );
  AOI21_X1 U14289 ( .B1(n14403), .B2(n12634), .A(n11840), .ZN(n11841) );
  OAI21_X1 U14290 ( .B1(n11842), .B2(n12637), .A(n11841), .ZN(P3_U3176) );
  OAI211_X1 U14291 ( .C1(n11844), .C2(n12287), .A(n11843), .B(n15106), .ZN(
        n11846) );
  AOI22_X1 U14292 ( .A1(n15103), .A2(n12664), .B1(n12662), .B2(n15104), .ZN(
        n11845) );
  NAND2_X1 U14293 ( .A1(n11846), .A2(n11845), .ZN(n11935) );
  INV_X1 U14294 ( .A(n11935), .ZN(n11852) );
  OAI21_X1 U14295 ( .B1(n6514), .B2(n8884), .A(n11847), .ZN(n11936) );
  INV_X1 U14296 ( .A(n12549), .ZN(n11848) );
  AOI22_X1 U14297 ( .A1(n15119), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n14400), 
        .B2(n11848), .ZN(n11849) );
  OAI21_X1 U14298 ( .B1(n12555), .B2(n12933), .A(n11849), .ZN(n11850) );
  AOI21_X1 U14299 ( .B1(n11936), .B2(n12935), .A(n11850), .ZN(n11851) );
  OAI21_X1 U14300 ( .B1(n11852), .B2(n15119), .A(n11851), .ZN(P3_U3219) );
  OAI22_X1 U14301 ( .A1(n14526), .A2(n12453), .B1(n11906), .B2(n12452), .ZN(
        n11893) );
  OAI22_X1 U14302 ( .A1(n14526), .A2(n12454), .B1(n11906), .B2(n12453), .ZN(
        n11853) );
  XNOR2_X1 U14303 ( .A(n11853), .B(n12444), .ZN(n11892) );
  XOR2_X1 U14304 ( .A(n11893), .B(n11892), .Z(n11860) );
  INV_X1 U14305 ( .A(n11854), .ZN(n11856) );
  OAI21_X1 U14306 ( .B1(n11860), .B2(n11859), .A(n11902), .ZN(n11861) );
  NAND2_X1 U14307 ( .A1(n11861), .A2(n13795), .ZN(n11867) );
  NOR2_X1 U14308 ( .A1(n13813), .A2(n11862), .ZN(n11863) );
  AOI211_X1 U14309 ( .C1(n13769), .C2(n11865), .A(n11864), .B(n11863), .ZN(
        n11866) );
  OAI211_X1 U14310 ( .C1(n14526), .C2(n13803), .A(n11867), .B(n11866), .ZN(
        P1_U3236) );
  AOI21_X1 U14311 ( .B1(n11870), .B2(n11868), .A(n6633), .ZN(n14506) );
  OAI211_X1 U14312 ( .C1(n11871), .C2(n11870), .A(n14618), .B(n11869), .ZN(
        n11872) );
  INV_X1 U14313 ( .A(n11872), .ZN(n14507) );
  OR2_X1 U14314 ( .A1(n13807), .A2(n14053), .ZN(n11874) );
  NAND2_X1 U14315 ( .A1(n13830), .A2(n14631), .ZN(n11873) );
  NAND2_X1 U14316 ( .A1(n11874), .A2(n11873), .ZN(n14502) );
  OAI21_X1 U14317 ( .B1(n14507), .B2(n14502), .A(n14665), .ZN(n11879) );
  OAI22_X1 U14318 ( .A1(n14665), .A2(n11875), .B1(n13812), .B2(n14673), .ZN(
        n11877) );
  OAI211_X1 U14319 ( .C1(n6642), .C2(n12057), .A(n11949), .B(n14679), .ZN(
        n14504) );
  NOR2_X1 U14320 ( .A1(n14504), .A2(n14065), .ZN(n11876) );
  AOI211_X1 U14321 ( .C1(n14677), .C2(n14503), .A(n11877), .B(n11876), .ZN(
        n11878) );
  OAI211_X1 U14322 ( .C1(n14506), .C2(n14083), .A(n11879), .B(n11878), .ZN(
        P1_U3278) );
  OAI222_X1 U14323 ( .A1(n14208), .A2(n11913), .B1(P1_U3086), .B2(n11881), 
        .C1(n11880), .C2(n12044), .ZN(P1_U3331) );
  INV_X1 U14324 ( .A(n11882), .ZN(n11883) );
  AOI21_X1 U14325 ( .B1(n11885), .B2(n11884), .A(n11883), .ZN(n11891) );
  AOI22_X1 U14326 ( .A1(n10675), .A2(n12664), .B1(P3_REG3_REG_12__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11887) );
  NAND2_X1 U14327 ( .A1(n12552), .A2(n12666), .ZN(n11886) );
  OAI211_X1 U14328 ( .C1(n12645), .C2(n11888), .A(n11887), .B(n11886), .ZN(
        n11889) );
  AOI21_X1 U14329 ( .B1(n12281), .B2(n12634), .A(n11889), .ZN(n11890) );
  OAI21_X1 U14330 ( .B1(n11891), .B2(n12637), .A(n11890), .ZN(P3_U3164) );
  INV_X1 U14331 ( .A(n11892), .ZN(n11895) );
  INV_X1 U14332 ( .A(n11893), .ZN(n11894) );
  NAND2_X1 U14333 ( .A1(n11895), .A2(n11894), .ZN(n11901) );
  AND2_X1 U14334 ( .A1(n11902), .A2(n11901), .ZN(n11904) );
  NAND2_X1 U14335 ( .A1(n11900), .A2(n12441), .ZN(n11897) );
  NAND2_X1 U14336 ( .A1(n13833), .A2(n12424), .ZN(n11896) );
  NAND2_X1 U14337 ( .A1(n11897), .A2(n11896), .ZN(n11898) );
  XNOR2_X1 U14338 ( .A(n11898), .B(n12444), .ZN(n11955) );
  AND2_X1 U14339 ( .A1(n12446), .A2(n13833), .ZN(n11899) );
  AOI21_X1 U14340 ( .B1(n11900), .B2(n12424), .A(n11899), .ZN(n11956) );
  XNOR2_X1 U14341 ( .A(n11955), .B(n11956), .ZN(n11903) );
  OAI211_X1 U14342 ( .C1(n11904), .C2(n11903), .A(n13795), .B(n11958), .ZN(
        n11911) );
  OAI21_X1 U14343 ( .B1(n13808), .B2(n11906), .A(n11905), .ZN(n11909) );
  NOR2_X1 U14344 ( .A1(n13813), .A2(n11907), .ZN(n11908) );
  AOI211_X1 U14345 ( .C1(n13810), .C2(n14483), .A(n11909), .B(n11908), .ZN(
        n11910) );
  OAI211_X1 U14346 ( .C1(n14337), .C2(n13803), .A(n11911), .B(n11910), .ZN(
        P1_U3224) );
  OAI222_X1 U14347 ( .A1(P2_U3088), .A2(n11914), .B1(n13643), .B2(n11913), 
        .C1(n11912), .C2(n13652), .ZN(P2_U3303) );
  XNOR2_X1 U14348 ( .A(n11915), .B(n12290), .ZN(n11917) );
  OAI22_X1 U14349 ( .A1(n11916), .A2(n12927), .B1(n12912), .B2(n12925), .ZN(
        n12114) );
  AOI21_X1 U14350 ( .B1(n11917), .B2(n15106), .A(n12114), .ZN(n13006) );
  XNOR2_X1 U14351 ( .A(n11918), .B(n12290), .ZN(n13004) );
  INV_X1 U14352 ( .A(n12116), .ZN(n11919) );
  AOI22_X1 U14353 ( .A1(n15119), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n14400), 
        .B2(n11919), .ZN(n11920) );
  OAI21_X1 U14354 ( .B1(n13007), .B2(n12933), .A(n11920), .ZN(n11921) );
  AOI21_X1 U14355 ( .B1(n13004), .B2(n12935), .A(n11921), .ZN(n11922) );
  OAI21_X1 U14356 ( .B1(n13006), .B2(n15119), .A(n11922), .ZN(P3_U3218) );
  XNOR2_X1 U14357 ( .A(n11924), .B(n12664), .ZN(n11925) );
  XNOR2_X1 U14358 ( .A(n11926), .B(n11925), .ZN(n11934) );
  OAI22_X1 U14359 ( .A1(n12632), .A2(n12280), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11927), .ZN(n11928) );
  AOI21_X1 U14360 ( .B1(n10675), .B2(n12663), .A(n11928), .ZN(n11929) );
  OAI21_X1 U14361 ( .B1(n12645), .B2(n11930), .A(n11929), .ZN(n11931) );
  AOI21_X1 U14362 ( .B1(n11932), .B2(n12634), .A(n11931), .ZN(n11933) );
  OAI21_X1 U14363 ( .B1(n11934), .B2(n12637), .A(n11933), .ZN(P3_U3174) );
  AOI21_X1 U14364 ( .B1(n14415), .B2(n11936), .A(n11935), .ZN(n11939) );
  MUX2_X1 U14365 ( .A(n11937), .B(n11939), .S(n15175), .Z(n11938) );
  OAI21_X1 U14366 ( .B1(n13059), .B2(n12555), .A(n11938), .ZN(P3_U3432) );
  INV_X1 U14367 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12683) );
  MUX2_X1 U14368 ( .A(n12683), .B(n11939), .S(n15183), .Z(n11940) );
  OAI21_X1 U14369 ( .B1(n13003), .B2(n12555), .A(n11940), .ZN(P3_U3473) );
  INV_X1 U14370 ( .A(n13717), .ZN(n11946) );
  OR2_X1 U14371 ( .A1(n13714), .A2(n14053), .ZN(n11942) );
  NAND2_X1 U14372 ( .A1(n14074), .A2(n14631), .ZN(n11941) );
  NAND2_X1 U14373 ( .A1(n11942), .A2(n11941), .ZN(n14495) );
  NAND2_X1 U14374 ( .A1(n11943), .A2(n11948), .ZN(n11944) );
  AOI21_X1 U14375 ( .B1(n11945), .B2(n11944), .A(n14690), .ZN(n14499) );
  AOI211_X1 U14376 ( .C1(n14643), .C2(n11946), .A(n14495), .B(n14499), .ZN(
        n11954) );
  XNOR2_X1 U14377 ( .A(n11947), .B(n11948), .ZN(n14501) );
  INV_X1 U14378 ( .A(n11949), .ZN(n11950) );
  INV_X1 U14379 ( .A(n13719), .ZN(n14498) );
  OAI211_X1 U14380 ( .C1(n11950), .C2(n14498), .A(n14679), .B(n11976), .ZN(
        n14497) );
  AOI22_X1 U14381 ( .A1(n13719), .A2(n14677), .B1(n14644), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n11951) );
  OAI21_X1 U14382 ( .B1(n14497), .B2(n14065), .A(n11951), .ZN(n11952) );
  AOI21_X1 U14383 ( .B1(n14501), .B2(n14662), .A(n11952), .ZN(n11953) );
  OAI21_X1 U14384 ( .B1(n11954), .B2(n14087), .A(n11953), .ZN(P1_U3277) );
  INV_X1 U14385 ( .A(n11956), .ZN(n11957) );
  OAI22_X1 U14386 ( .A1(n11959), .A2(n12454), .B1(n12003), .B2(n12453), .ZN(
        n11960) );
  XNOR2_X1 U14387 ( .A(n11960), .B(n12444), .ZN(n11995) );
  AND2_X1 U14388 ( .A1(n12446), .A2(n14483), .ZN(n11961) );
  AOI21_X1 U14389 ( .B1(n14518), .B2(n12424), .A(n11961), .ZN(n11994) );
  XNOR2_X1 U14390 ( .A(n11995), .B(n11994), .ZN(n11997) );
  XNOR2_X1 U14391 ( .A(n11998), .B(n11997), .ZN(n11968) );
  NAND2_X1 U14392 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n14588)
         );
  OAI21_X1 U14393 ( .B1(n13808), .B2(n11962), .A(n14588), .ZN(n11963) );
  AOI21_X1 U14394 ( .B1(n13810), .B2(n13832), .A(n11963), .ZN(n11964) );
  OAI21_X1 U14395 ( .B1(n13813), .B2(n11965), .A(n11964), .ZN(n11966) );
  AOI21_X1 U14396 ( .B1(n14518), .B2(n13815), .A(n11966), .ZN(n11967) );
  OAI21_X1 U14397 ( .B1(n11968), .B2(n13817), .A(n11967), .ZN(P1_U3234) );
  NAND2_X1 U14398 ( .A1(n11969), .A2(n11974), .ZN(n11970) );
  NAND3_X1 U14399 ( .A1(n11971), .A2(n14618), .A3(n11970), .ZN(n11973) );
  AOI22_X1 U14400 ( .A1(n13829), .A2(n14631), .B1(n14482), .B2(n13830), .ZN(
        n11972) );
  NAND2_X1 U14401 ( .A1(n11973), .A2(n11972), .ZN(n14181) );
  INV_X1 U14402 ( .A(n14181), .ZN(n11983) );
  XNOR2_X1 U14403 ( .A(n11975), .B(n11974), .ZN(n14176) );
  AOI21_X1 U14404 ( .B1(n11976), .B2(n13734), .A(n14699), .ZN(n11977) );
  NAND2_X1 U14405 ( .A1(n11977), .A2(n14070), .ZN(n14177) );
  OAI22_X1 U14406 ( .A1(n14665), .A2(n11978), .B1(n13742), .B2(n14673), .ZN(
        n11979) );
  AOI21_X1 U14407 ( .B1(n13734), .B2(n14677), .A(n11979), .ZN(n11980) );
  OAI21_X1 U14408 ( .B1(n14177), .B2(n14065), .A(n11980), .ZN(n11981) );
  AOI21_X1 U14409 ( .B1(n14176), .B2(n14662), .A(n11981), .ZN(n11982) );
  OAI21_X1 U14410 ( .B1(n11983), .B2(n14087), .A(n11982), .ZN(P1_U3276) );
  INV_X1 U14411 ( .A(n11984), .ZN(n11989) );
  OAI222_X1 U14412 ( .A1(n11986), .A2(P2_U3088), .B1(n13643), .B2(n11989), 
        .C1(n11985), .C2(n13652), .ZN(P2_U3302) );
  INV_X1 U14413 ( .A(n11987), .ZN(n11988) );
  OAI222_X1 U14414 ( .A1(n12044), .A2(n11990), .B1(n14214), .B2(n11989), .C1(
        n11988), .C2(P1_U3086), .ZN(P1_U3330) );
  INV_X1 U14415 ( .A(n14511), .ZN(n14489) );
  AOI22_X1 U14416 ( .A1(n14511), .A2(n12441), .B1(n12424), .B2(n13832), .ZN(
        n11991) );
  XOR2_X1 U14417 ( .A(n12444), .B(n11991), .Z(n11993) );
  OAI22_X1 U14418 ( .A1(n14489), .A2(n12453), .B1(n13807), .B2(n12452), .ZN(
        n11992) );
  NOR2_X1 U14419 ( .A1(n11993), .A2(n11992), .ZN(n12054) );
  AOI21_X1 U14420 ( .B1(n11993), .B2(n11992), .A(n12054), .ZN(n12000) );
  INV_X1 U14421 ( .A(n11994), .ZN(n11996) );
  AOI22_X2 U14422 ( .A1(n11998), .A2(n11997), .B1(n11996), .B2(n11995), .ZN(
        n11999) );
  OAI21_X1 U14423 ( .B1(n12000), .B2(n11999), .A(n12056), .ZN(n12001) );
  NAND2_X1 U14424 ( .A1(n12001), .A2(n13795), .ZN(n12007) );
  NOR2_X1 U14425 ( .A1(n13714), .A2(n14055), .ZN(n14477) );
  OAI21_X1 U14426 ( .B1(n13808), .B2(n12003), .A(n12002), .ZN(n12005) );
  NOR2_X1 U14427 ( .A1(n13813), .A2(n14484), .ZN(n12004) );
  AOI211_X1 U14428 ( .C1(n13769), .C2(n14477), .A(n12005), .B(n12004), .ZN(
        n12006) );
  OAI211_X1 U14429 ( .C1(n14489), .C2(n13803), .A(n12007), .B(n12006), .ZN(
        P1_U3215) );
  OAI222_X1 U14430 ( .A1(P2_U3088), .A2(n12008), .B1(n13643), .B2(n9665), .C1(
        n12138), .C2(n13652), .ZN(P2_U3297) );
  INV_X1 U14431 ( .A(n12009), .ZN(n12130) );
  OAI222_X1 U14432 ( .A1(n12044), .A2(n12010), .B1(n14208), .B2(n12130), .C1(
        n8333), .C2(P1_U3086), .ZN(P1_U3336) );
  INV_X1 U14433 ( .A(n13823), .ZN(n13958) );
  INV_X1 U14434 ( .A(n13822), .ZN(n13661) );
  AOI22_X1 U14435 ( .A1(n13955), .A2(n13954), .B1(n13661), .B2(n13967), .ZN(
        n13941) );
  OAI22_X2 U14436 ( .A1(n13941), .A2(n13940), .B1(n6872), .B2(n13956), .ZN(
        n12480) );
  NAND2_X1 U14437 ( .A1(n13820), .A2(n14631), .ZN(n12013) );
  INV_X1 U14438 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n12016) );
  OAI22_X1 U14439 ( .A1(n12459), .A2(n14673), .B1(n12016), .B2(n14665), .ZN(
        n12018) );
  NAND2_X1 U14440 ( .A1(n12478), .A2(n13944), .ZN(n12483) );
  OAI211_X1 U14441 ( .C1(n12478), .C2(n13944), .A(n14679), .B(n12483), .ZN(
        n14107) );
  NOR2_X1 U14442 ( .A1(n14107), .A2(n14065), .ZN(n12017) );
  AOI211_X1 U14443 ( .C1(n14677), .C2(n14104), .A(n12018), .B(n12017), .ZN(
        n12027) );
  NAND2_X1 U14444 ( .A1(n14125), .A2(n13823), .ZN(n12019) );
  INV_X1 U14445 ( .A(n13954), .ZN(n13961) );
  NAND2_X1 U14446 ( .A1(n13967), .A2(n13822), .ZN(n12020) );
  INV_X1 U14447 ( .A(n13940), .ZN(n13950) );
  OR2_X1 U14448 ( .A1(n14112), .A2(n13956), .ZN(n12021) );
  INV_X1 U14449 ( .A(n12025), .ZN(n12023) );
  INV_X1 U14450 ( .A(n12024), .ZN(n12022) );
  NAND2_X1 U14451 ( .A1(n12025), .A2(n12024), .ZN(n14105) );
  NAND3_X1 U14452 ( .A1(n14106), .A2(n14662), .A3(n14105), .ZN(n12026) );
  OAI211_X1 U14453 ( .C1(n14110), .C2(n14644), .A(n12027), .B(n12026), .ZN(
        P1_U3265) );
  INV_X1 U14454 ( .A(n14789), .ZN(n13208) );
  INV_X1 U14455 ( .A(n12028), .ZN(n12038) );
  NAND2_X1 U14456 ( .A1(n14430), .A2(n12029), .ZN(n12031) );
  OAI211_X1 U14457 ( .C1(n13210), .C2(n14930), .A(n12031), .B(n12030), .ZN(
        n12037) );
  INV_X1 U14458 ( .A(n10490), .ZN(n12035) );
  AOI22_X1 U14459 ( .A1(n13225), .A2(n13266), .B1(n14428), .B2(n12032), .ZN(
        n12034) );
  NOR3_X1 U14460 ( .A1(n12035), .A2(n12034), .A3(n12033), .ZN(n12036) );
  AOI211_X1 U14461 ( .C1(n13208), .C2(n12038), .A(n12037), .B(n12036), .ZN(
        n12039) );
  OAI21_X1 U14462 ( .B1(n14782), .B2(n12040), .A(n12039), .ZN(P2_U3199) );
  INV_X1 U14463 ( .A(n12041), .ZN(n13647) );
  OAI222_X1 U14464 ( .A1(n12044), .A2(n12042), .B1(n14208), .B2(n13647), .C1(
        n8325), .C2(P1_U3086), .ZN(P1_U3327) );
  INV_X1 U14465 ( .A(n12043), .ZN(n13642) );
  OAI222_X1 U14466 ( .A1(n14214), .A2(n13642), .B1(n7522), .B2(P1_U3086), .C1(
        n12134), .C2(n12044), .ZN(P1_U3326) );
  OAI22_X1 U14467 ( .A1(n8295), .A2(n12454), .B1(n13691), .B2(n12453), .ZN(
        n12045) );
  XNOR2_X1 U14468 ( .A(n12045), .B(n12444), .ZN(n12049) );
  OR2_X1 U14469 ( .A1(n8295), .A2(n12453), .ZN(n12047) );
  NAND2_X1 U14470 ( .A1(n13826), .A2(n12446), .ZN(n12046) );
  NAND2_X1 U14471 ( .A1(n12047), .A2(n12046), .ZN(n12048) );
  NOR2_X1 U14472 ( .A1(n12049), .A2(n12048), .ZN(n13669) );
  AOI21_X1 U14473 ( .B1(n12049), .B2(n12048), .A(n13669), .ZN(n12101) );
  AND2_X1 U14474 ( .A1(n14075), .A2(n12446), .ZN(n12050) );
  AOI21_X1 U14475 ( .B1(n14062), .B2(n12424), .A(n12050), .ZN(n12084) );
  NAND2_X1 U14476 ( .A1(n14062), .A2(n12441), .ZN(n12052) );
  NAND2_X1 U14477 ( .A1(n14075), .A2(n12424), .ZN(n12051) );
  NAND2_X1 U14478 ( .A1(n12052), .A2(n12051), .ZN(n12053) );
  XNOR2_X1 U14479 ( .A(n12053), .B(n12444), .ZN(n12079) );
  INV_X1 U14480 ( .A(n12054), .ZN(n12055) );
  NAND2_X1 U14481 ( .A1(n12056), .A2(n12055), .ZN(n12059) );
  OAI22_X1 U14482 ( .A1(n12057), .A2(n12454), .B1(n13714), .B2(n12453), .ZN(
        n12058) );
  XOR2_X1 U14483 ( .A(n12444), .B(n12058), .Z(n12060) );
  AOI22_X1 U14484 ( .A1(n14503), .A2(n12424), .B1(n12446), .B2(n13831), .ZN(
        n13804) );
  OAI22_X1 U14485 ( .A1(n13805), .A2(n13804), .B1(n12060), .B2(n12059), .ZN(
        n13711) );
  NAND2_X1 U14486 ( .A1(n13719), .A2(n12441), .ZN(n12062) );
  NAND2_X1 U14487 ( .A1(n13830), .A2(n12424), .ZN(n12061) );
  NAND2_X1 U14488 ( .A1(n12062), .A2(n12061), .ZN(n12063) );
  XNOR2_X1 U14489 ( .A(n12063), .B(n6519), .ZN(n12066) );
  AND2_X1 U14490 ( .A1(n12446), .A2(n13830), .ZN(n12064) );
  AOI21_X1 U14491 ( .B1(n13719), .B2(n12424), .A(n12064), .ZN(n12065) );
  NAND2_X1 U14492 ( .A1(n12066), .A2(n12065), .ZN(n12067) );
  OAI21_X1 U14493 ( .B1(n12066), .B2(n12065), .A(n12067), .ZN(n13712) );
  NOR2_X2 U14494 ( .A1(n13711), .A2(n13712), .ZN(n13710) );
  INV_X1 U14495 ( .A(n12067), .ZN(n13737) );
  NAND2_X1 U14496 ( .A1(n13734), .A2(n12441), .ZN(n12069) );
  NAND2_X1 U14497 ( .A1(n14074), .A2(n12424), .ZN(n12068) );
  NAND2_X1 U14498 ( .A1(n12069), .A2(n12068), .ZN(n12070) );
  XNOR2_X1 U14499 ( .A(n12070), .B(n12444), .ZN(n12074) );
  NAND2_X1 U14500 ( .A1(n13734), .A2(n12424), .ZN(n12072) );
  NAND2_X1 U14501 ( .A1(n14074), .A2(n12446), .ZN(n12071) );
  NAND2_X1 U14502 ( .A1(n12072), .A2(n12071), .ZN(n12073) );
  NOR2_X1 U14503 ( .A1(n12074), .A2(n12073), .ZN(n12075) );
  AOI21_X1 U14504 ( .B1(n12074), .B2(n12073), .A(n12075), .ZN(n13736) );
  NAND2_X1 U14505 ( .A1(n14172), .A2(n12441), .ZN(n12077) );
  NAND2_X1 U14506 ( .A1(n13829), .A2(n12424), .ZN(n12076) );
  NAND2_X1 U14507 ( .A1(n12077), .A2(n12076), .ZN(n12078) );
  XNOR2_X1 U14508 ( .A(n12078), .B(n12444), .ZN(n12080) );
  AOI22_X1 U14509 ( .A1(n14172), .A2(n12424), .B1(n12446), .B2(n13829), .ZN(
        n12081) );
  XNOR2_X1 U14510 ( .A(n12080), .B(n12081), .ZN(n13784) );
  XNOR2_X1 U14511 ( .A(n12079), .B(n12084), .ZN(n13681) );
  INV_X1 U14512 ( .A(n12080), .ZN(n12082) );
  NAND2_X1 U14513 ( .A1(n12082), .A2(n12081), .ZN(n13679) );
  AND2_X1 U14514 ( .A1(n13828), .A2(n12446), .ZN(n12085) );
  AOI21_X1 U14515 ( .B1(n14159), .B2(n12424), .A(n12085), .ZN(n12087) );
  AOI22_X1 U14516 ( .A1(n14159), .A2(n12441), .B1(n12424), .B2(n13828), .ZN(
        n12086) );
  XNOR2_X1 U14517 ( .A(n12086), .B(n12444), .ZN(n12088) );
  XOR2_X1 U14518 ( .A(n12087), .B(n12088), .Z(n13774) );
  INV_X1 U14519 ( .A(n12087), .ZN(n12090) );
  INV_X1 U14520 ( .A(n12088), .ZN(n12089) );
  NAND2_X1 U14521 ( .A1(n14151), .A2(n12441), .ZN(n12092) );
  NAND2_X1 U14522 ( .A1(n13827), .A2(n12424), .ZN(n12091) );
  NAND2_X1 U14523 ( .A1(n12092), .A2(n12091), .ZN(n12093) );
  XNOR2_X1 U14524 ( .A(n12093), .B(n12444), .ZN(n12097) );
  NAND2_X1 U14525 ( .A1(n14151), .A2(n12424), .ZN(n12095) );
  NAND2_X1 U14526 ( .A1(n13827), .A2(n12446), .ZN(n12094) );
  NAND2_X1 U14527 ( .A1(n12095), .A2(n12094), .ZN(n12096) );
  NOR2_X1 U14528 ( .A1(n12097), .A2(n12096), .ZN(n12098) );
  AOI21_X1 U14529 ( .B1(n12097), .B2(n12096), .A(n12098), .ZN(n13688) );
  NAND2_X1 U14530 ( .A1(n13689), .A2(n13688), .ZN(n13687) );
  INV_X1 U14531 ( .A(n12098), .ZN(n12099) );
  OAI21_X1 U14532 ( .B1(n12101), .B2(n12100), .A(n13667), .ZN(n12102) );
  NAND2_X1 U14533 ( .A1(n12102), .A2(n13795), .ZN(n12109) );
  NAND2_X1 U14534 ( .A1(n13825), .A2(n14631), .ZN(n12104) );
  NAND2_X1 U14535 ( .A1(n13827), .A2(n14482), .ZN(n12103) );
  NAND2_X1 U14536 ( .A1(n12104), .A2(n12103), .ZN(n14142) );
  INV_X1 U14537 ( .A(n14009), .ZN(n12106) );
  OAI22_X1 U14538 ( .A1(n12106), .A2(n13813), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12105), .ZN(n12107) );
  AOI21_X1 U14539 ( .B1(n14142), .B2(n13769), .A(n12107), .ZN(n12108) );
  OAI211_X1 U14540 ( .C1(n13803), .C2(n8295), .A(n12109), .B(n12108), .ZN(
        P1_U3235) );
  NAND2_X1 U14541 ( .A1(n12111), .A2(n12110), .ZN(n12113) );
  XNOR2_X1 U14542 ( .A(n12113), .B(n12112), .ZN(n12120) );
  AOI22_X1 U14543 ( .A1(n12647), .A2(n12114), .B1(P3_REG3_REG_15__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12115) );
  OAI21_X1 U14544 ( .B1(n12645), .B2(n12116), .A(n12115), .ZN(n12117) );
  AOI21_X1 U14545 ( .B1(n12118), .B2(n12634), .A(n12117), .ZN(n12119) );
  OAI21_X1 U14546 ( .B1(n12120), .B2(n12637), .A(n12119), .ZN(P3_U3181) );
  XNOR2_X1 U14547 ( .A(n12122), .B(n12661), .ZN(n12123) );
  XNOR2_X1 U14548 ( .A(n12121), .B(n12123), .ZN(n12128) );
  NAND2_X1 U14549 ( .A1(n12629), .A2(n12931), .ZN(n12125) );
  AOI22_X1 U14550 ( .A1(n12552), .A2(n12662), .B1(P3_REG3_REG_16__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12124) );
  OAI211_X1 U14551 ( .C1(n12924), .C2(n12608), .A(n12125), .B(n12124), .ZN(
        n12126) );
  AOI21_X1 U14552 ( .B1(n12930), .B2(n12634), .A(n12126), .ZN(n12127) );
  OAI21_X1 U14553 ( .B1(n12128), .B2(n12637), .A(n12127), .ZN(P3_U3166) );
  OAI222_X1 U14554 ( .A1(n9432), .A2(P2_U3088), .B1(n13643), .B2(n12130), .C1(
        n12129), .C2(n13652), .ZN(P2_U3308) );
  INV_X1 U14555 ( .A(n12368), .ZN(n12131) );
  INV_X1 U14556 ( .A(n12133), .ZN(n12136) );
  NAND2_X1 U14557 ( .A1(n12134), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12135) );
  NAND2_X1 U14558 ( .A1(n12138), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12140) );
  NAND2_X1 U14559 ( .A1(n12526), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12139) );
  NAND2_X1 U14560 ( .A1(n12140), .A2(n12139), .ZN(n12154) );
  OR2_X2 U14561 ( .A1(n12155), .A2(n12154), .ZN(n12157) );
  NAND2_X1 U14562 ( .A1(n12157), .A2(n12140), .ZN(n12142) );
  XNOR2_X1 U14563 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n12141) );
  XNOR2_X1 U14564 ( .A(n12142), .B(n12141), .ZN(n13071) );
  NAND2_X1 U14565 ( .A1(n13071), .A2(n12159), .ZN(n12144) );
  INV_X1 U14566 ( .A(SI_31_), .ZN(n13066) );
  OR2_X1 U14567 ( .A1(n8529), .A2(n13066), .ZN(n12143) );
  NAND2_X1 U14568 ( .A1(n12145), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12151) );
  INV_X1 U14569 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n12146) );
  OR2_X1 U14570 ( .A1(n8865), .A2(n12146), .ZN(n12150) );
  INV_X1 U14571 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n12147) );
  OR2_X1 U14572 ( .A1(n12148), .A2(n12147), .ZN(n12149) );
  NAND4_X1 U14573 ( .A1(n12152), .A2(n12151), .A3(n12150), .A4(n12149), .ZN(
        n12763) );
  INV_X1 U14574 ( .A(n12763), .ZN(n12153) );
  INV_X1 U14575 ( .A(n12369), .ZN(n12161) );
  NAND2_X1 U14576 ( .A1(n12155), .A2(n12154), .ZN(n12156) );
  NAND2_X1 U14577 ( .A1(n12157), .A2(n12156), .ZN(n12542) );
  NOR2_X1 U14578 ( .A1(n8529), .A2(n15229), .ZN(n12158) );
  AOI21_X2 U14579 ( .B1(n12542), .B2(n12159), .A(n12158), .ZN(n13013) );
  AOI21_X1 U14580 ( .B1(n12763), .B2(n12650), .A(n13013), .ZN(n12160) );
  NOR2_X1 U14581 ( .A1(n13010), .A2(n12763), .ZN(n12191) );
  AND2_X1 U14582 ( .A1(n13013), .A2(n12650), .ZN(n12164) );
  INV_X1 U14583 ( .A(n12164), .ZN(n12367) );
  INV_X1 U14584 ( .A(n13013), .ZN(n12942) );
  INV_X1 U14585 ( .A(n12650), .ZN(n12165) );
  NAND2_X1 U14586 ( .A1(n12942), .A2(n12165), .ZN(n12365) );
  NAND2_X1 U14587 ( .A1(n12367), .A2(n12365), .ZN(n12361) );
  INV_X1 U14588 ( .A(n12771), .ZN(n12189) );
  INV_X1 U14589 ( .A(n12166), .ZN(n12353) );
  INV_X1 U14590 ( .A(n12167), .ZN(n12168) );
  INV_X1 U14591 ( .A(n12335), .ZN(n12170) );
  INV_X1 U14592 ( .A(n12171), .ZN(n12172) );
  NAND2_X1 U14593 ( .A1(n12272), .A2(n12172), .ZN(n12262) );
  NAND4_X1 U14594 ( .A1(n12176), .A2(n12175), .A3(n12174), .A4(n12173), .ZN(
        n12178) );
  NAND3_X1 U14595 ( .A1(n12230), .A2(n12228), .A3(n12252), .ZN(n12177) );
  NOR2_X1 U14596 ( .A1(n12178), .A2(n12177), .ZN(n12180) );
  NAND4_X1 U14597 ( .A1(n12180), .A2(n12246), .A3(n12179), .A4(n12257), .ZN(
        n12181) );
  NOR4_X1 U14598 ( .A1(n12183), .A2(n12262), .A3(n12182), .A4(n12181), .ZN(
        n12184) );
  NAND4_X1 U14599 ( .A1(n6765), .A2(n12290), .A3(n8884), .A4(n12184), .ZN(
        n12185) );
  NOR4_X1 U14600 ( .A1(n12885), .A2(n12900), .A3(n6763), .A4(n12185), .ZN(
        n12186) );
  INV_X1 U14601 ( .A(n12871), .ZN(n12875) );
  NAND4_X1 U14602 ( .A1(n12864), .A2(n12854), .A3(n12186), .A4(n12875), .ZN(
        n12187) );
  NOR3_X1 U14603 ( .A1(n12826), .A2(n12336), .A3(n12187), .ZN(n12188) );
  NAND4_X1 U14604 ( .A1(n12189), .A2(n12813), .A3(n12800), .A4(n12188), .ZN(
        n12190) );
  NOR4_X1 U14605 ( .A1(n12361), .A2(n12198), .A3(n12190), .A4(n12785), .ZN(
        n12192) );
  INV_X1 U14606 ( .A(n12191), .ZN(n12372) );
  NAND3_X1 U14607 ( .A1(n12192), .A2(n6541), .A3(n12372), .ZN(n12193) );
  XNOR2_X1 U14608 ( .A(n12193), .B(n8454), .ZN(n12194) );
  OAI22_X1 U14609 ( .A1(n12197), .A2(n12196), .B1(n12195), .B2(n12194), .ZN(
        n12378) );
  INV_X1 U14610 ( .A(n12198), .ZN(n12363) );
  OR2_X1 U14611 ( .A1(n12771), .A2(n12785), .ZN(n12205) );
  NAND2_X1 U14612 ( .A1(n12200), .A2(n12199), .ZN(n12202) );
  NAND2_X1 U14613 ( .A1(n12202), .A2(n12201), .ZN(n12203) );
  NAND2_X1 U14614 ( .A1(n12205), .A2(n12203), .ZN(n12204) );
  INV_X1 U14615 ( .A(n12205), .ZN(n12358) );
  INV_X1 U14616 ( .A(n12854), .ZN(n12332) );
  MUX2_X1 U14617 ( .A(n12207), .B(n6819), .S(n12370), .Z(n12208) );
  INV_X1 U14618 ( .A(n12208), .ZN(n12330) );
  INV_X1 U14619 ( .A(n12213), .ZN(n12210) );
  NAND2_X1 U14620 ( .A1(n8874), .A2(n12364), .ZN(n12209) );
  OAI21_X1 U14621 ( .B1(n15105), .B2(n12210), .A(n12209), .ZN(n12216) );
  NAND2_X1 U14622 ( .A1(n12212), .A2(n12211), .ZN(n12214) );
  NAND3_X1 U14623 ( .A1(n12214), .A2(n12364), .A3(n12213), .ZN(n12215) );
  AOI21_X1 U14624 ( .B1(n12216), .B2(n12215), .A(n15093), .ZN(n12219) );
  MUX2_X1 U14625 ( .A(n12217), .B(n8874), .S(n12370), .Z(n12218) );
  NAND2_X1 U14626 ( .A1(n12219), .A2(n12218), .ZN(n12223) );
  NAND2_X1 U14627 ( .A1(n12229), .A2(n12220), .ZN(n12221) );
  NAND2_X1 U14628 ( .A1(n12221), .A2(n12364), .ZN(n12222) );
  NAND2_X1 U14629 ( .A1(n12223), .A2(n12222), .ZN(n12227) );
  NAND2_X1 U14630 ( .A1(n9772), .A2(n15088), .ZN(n12224) );
  AOI21_X1 U14631 ( .B1(n12226), .B2(n12224), .A(n12364), .ZN(n12225) );
  AOI21_X1 U14632 ( .B1(n12227), .B2(n12226), .A(n12225), .ZN(n12232) );
  OAI21_X1 U14633 ( .B1(n12364), .B2(n12229), .A(n12228), .ZN(n12231) );
  OAI21_X1 U14634 ( .B1(n12232), .B2(n12231), .A(n12230), .ZN(n12241) );
  NAND2_X1 U14635 ( .A1(n12243), .A2(n12233), .ZN(n12235) );
  NAND2_X1 U14636 ( .A1(n12235), .A2(n12364), .ZN(n12240) );
  NOR2_X1 U14637 ( .A1(n12235), .A2(n12234), .ZN(n12238) );
  INV_X1 U14638 ( .A(n12236), .ZN(n12237) );
  MUX2_X1 U14639 ( .A(n12238), .B(n12237), .S(n12370), .Z(n12239) );
  AOI21_X1 U14640 ( .B1(n12241), .B2(n12240), .A(n12239), .ZN(n12248) );
  AOI21_X1 U14641 ( .B1(n12244), .B2(n12242), .A(n12364), .ZN(n12247) );
  MUX2_X1 U14642 ( .A(n12244), .B(n12243), .S(n12370), .Z(n12245) );
  OAI211_X1 U14643 ( .C1(n12248), .C2(n12247), .A(n12246), .B(n12245), .ZN(
        n12253) );
  NAND2_X1 U14644 ( .A1(n15149), .A2(n12370), .ZN(n12250) );
  NAND2_X1 U14645 ( .A1(n6766), .A2(n12364), .ZN(n12249) );
  MUX2_X1 U14646 ( .A(n12250), .B(n12249), .S(n12670), .Z(n12251) );
  NAND3_X1 U14647 ( .A1(n12253), .A2(n12252), .A3(n12251), .ZN(n12258) );
  MUX2_X1 U14648 ( .A(n12669), .B(n12364), .S(n15155), .Z(n12254) );
  INV_X1 U14649 ( .A(n12254), .ZN(n12255) );
  OAI21_X1 U14650 ( .B1(n12364), .B2(n12669), .A(n12255), .ZN(n12256) );
  NAND3_X1 U14651 ( .A1(n12258), .A2(n12257), .A3(n12256), .ZN(n12269) );
  AND2_X1 U14652 ( .A1(n12668), .A2(n15161), .ZN(n12260) );
  NOR2_X1 U14653 ( .A1(n12668), .A2(n15161), .ZN(n12259) );
  MUX2_X1 U14654 ( .A(n12260), .B(n12259), .S(n12370), .Z(n12261) );
  NOR2_X1 U14655 ( .A1(n12262), .A2(n12261), .ZN(n12268) );
  NAND2_X1 U14656 ( .A1(n12272), .A2(n7277), .ZN(n12266) );
  NAND3_X1 U14657 ( .A1(n12266), .A2(n12265), .A3(n12264), .ZN(n12267) );
  AOI22_X1 U14658 ( .A1(n12269), .A2(n12268), .B1(n12370), .B2(n12267), .ZN(
        n12279) );
  INV_X1 U14659 ( .A(n12274), .ZN(n12278) );
  INV_X1 U14660 ( .A(n12270), .ZN(n12271) );
  NAND2_X1 U14661 ( .A1(n12272), .A2(n12271), .ZN(n12275) );
  NAND3_X1 U14662 ( .A1(n12275), .A2(n12274), .A3(n12273), .ZN(n12276) );
  NAND2_X1 U14663 ( .A1(n12276), .A2(n12364), .ZN(n12277) );
  OAI21_X1 U14664 ( .B1(n12279), .B2(n12278), .A(n12277), .ZN(n12284) );
  OR3_X1 U14665 ( .A1(n12281), .A2(n12280), .A3(n12370), .ZN(n12282) );
  NAND3_X1 U14666 ( .A1(n12284), .A2(n12283), .A3(n12282), .ZN(n12289) );
  MUX2_X1 U14667 ( .A(n12285), .B(n6535), .S(n12370), .Z(n12286) );
  INV_X1 U14668 ( .A(n12286), .ZN(n12288) );
  AOI21_X1 U14669 ( .B1(n12289), .B2(n12288), .A(n12287), .ZN(n12294) );
  INV_X1 U14670 ( .A(n12290), .ZN(n12293) );
  AND2_X1 U14671 ( .A1(n12292), .A2(n12291), .ZN(n12295) );
  OAI22_X1 U14672 ( .A1(n12294), .A2(n12293), .B1(n12370), .B2(n12295), .ZN(
        n12302) );
  AND2_X1 U14673 ( .A1(n12555), .A2(n12663), .ZN(n12299) );
  INV_X1 U14674 ( .A(n12295), .ZN(n12297) );
  NOR2_X1 U14675 ( .A1(n12297), .A2(n12296), .ZN(n12298) );
  MUX2_X1 U14676 ( .A(n12299), .B(n12298), .S(n12364), .Z(n12300) );
  INV_X1 U14677 ( .A(n12300), .ZN(n12301) );
  NAND3_X1 U14678 ( .A1(n12302), .A2(n12301), .A3(n12304), .ZN(n12307) );
  NAND2_X1 U14679 ( .A1(n12304), .A2(n12303), .ZN(n12305) );
  NAND2_X1 U14680 ( .A1(n12305), .A2(n12370), .ZN(n12306) );
  NAND2_X1 U14681 ( .A1(n12307), .A2(n12306), .ZN(n12310) );
  OR3_X1 U14682 ( .A1(n12930), .A2(n12912), .A3(n12364), .ZN(n12309) );
  NAND2_X1 U14683 ( .A1(n12897), .A2(n12913), .ZN(n12308) );
  AOI21_X1 U14684 ( .B1(n12310), .B2(n12309), .A(n12308), .ZN(n12324) );
  INV_X1 U14685 ( .A(n12316), .ZN(n12313) );
  OAI211_X1 U14686 ( .C1(n12313), .C2(n12312), .A(n12321), .B(n12311), .ZN(
        n12319) );
  INV_X1 U14687 ( .A(n12314), .ZN(n12315) );
  NAND2_X1 U14688 ( .A1(n12897), .A2(n12315), .ZN(n12317) );
  NAND3_X1 U14689 ( .A1(n12317), .A2(n12320), .A3(n12316), .ZN(n12318) );
  MUX2_X1 U14690 ( .A(n12319), .B(n12318), .S(n12364), .Z(n12323) );
  MUX2_X1 U14691 ( .A(n12321), .B(n12320), .S(n12370), .Z(n12322) );
  OAI211_X1 U14692 ( .C1(n12324), .C2(n12323), .A(n12875), .B(n12322), .ZN(
        n12328) );
  NAND2_X1 U14693 ( .A1(n12887), .A2(n12370), .ZN(n12326) );
  OR2_X1 U14694 ( .A1(n12887), .A2(n12370), .ZN(n12325) );
  MUX2_X1 U14695 ( .A(n12326), .B(n12325), .S(n12877), .Z(n12327) );
  NAND3_X1 U14696 ( .A1(n12864), .A2(n12328), .A3(n12327), .ZN(n12329) );
  NAND2_X1 U14697 ( .A1(n12330), .A2(n12329), .ZN(n12331) );
  NOR2_X1 U14698 ( .A1(n12332), .A2(n12331), .ZN(n12338) );
  INV_X1 U14699 ( .A(n12333), .ZN(n12334) );
  MUX2_X1 U14700 ( .A(n12335), .B(n12334), .S(n12370), .Z(n12337) );
  OR3_X1 U14701 ( .A1(n12338), .A2(n12337), .A3(n12336), .ZN(n12340) );
  NAND3_X1 U14702 ( .A1(n12966), .A2(n12828), .A3(n12370), .ZN(n12339) );
  AND2_X1 U14703 ( .A1(n12340), .A2(n12339), .ZN(n12348) );
  INV_X1 U14704 ( .A(n12341), .ZN(n12342) );
  NAND2_X1 U14705 ( .A1(n12346), .A2(n12342), .ZN(n12344) );
  AND2_X1 U14706 ( .A1(n12344), .A2(n12343), .ZN(n12345) );
  MUX2_X1 U14707 ( .A(n12346), .B(n12345), .S(n12364), .Z(n12347) );
  OAI211_X1 U14708 ( .C1(n12348), .C2(n12826), .A(n12347), .B(n12813), .ZN(
        n12352) );
  MUX2_X1 U14709 ( .A(n12350), .B(n12349), .S(n12370), .Z(n12351) );
  NAND3_X1 U14710 ( .A1(n12800), .A2(n12352), .A3(n12351), .ZN(n12356) );
  MUX2_X1 U14711 ( .A(n12354), .B(n12353), .S(n12370), .Z(n12355) );
  NAND2_X1 U14712 ( .A1(n12356), .A2(n12355), .ZN(n12357) );
  NAND2_X1 U14713 ( .A1(n12358), .A2(n12357), .ZN(n12359) );
  NAND2_X1 U14714 ( .A1(n12360), .A2(n12359), .ZN(n12362) );
  AOI21_X1 U14715 ( .B1(n12363), .B2(n12362), .A(n12361), .ZN(n12371) );
  NAND2_X1 U14716 ( .A1(n12365), .A2(n12364), .ZN(n12366) );
  AOI22_X1 U14717 ( .A1(n12371), .A2(n12368), .B1(n12367), .B2(n12366), .ZN(
        n12375) );
  NAND3_X1 U14718 ( .A1(n12371), .A2(n12370), .A3(n12369), .ZN(n12373) );
  NAND2_X1 U14719 ( .A1(n12373), .A2(n12372), .ZN(n12374) );
  OAI21_X1 U14720 ( .B1(n12375), .B2(n12374), .A(n6541), .ZN(n12376) );
  NAND4_X1 U14721 ( .A1(n12381), .A2(n12380), .A3(n12379), .A4(n15103), .ZN(
        n12382) );
  OAI211_X1 U14722 ( .C1(n12384), .C2(n12383), .A(n12382), .B(P3_B_REG_SCAN_IN), .ZN(n12385) );
  NAND2_X1 U14723 ( .A1(n12386), .A2(n12385), .ZN(P3_U3296) );
  NOR2_X1 U14724 ( .A1(n14789), .A2(n12387), .ZN(n12390) );
  NAND2_X1 U14725 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n14824) );
  OAI21_X1 U14726 ( .B1(n14779), .B2(n12388), .A(n14824), .ZN(n12389) );
  AOI211_X1 U14727 ( .C1(n12391), .C2(n14787), .A(n12390), .B(n12389), .ZN(
        n12399) );
  INV_X1 U14728 ( .A(n12392), .ZN(n12396) );
  OAI22_X1 U14729 ( .A1(n12394), .A2(n14782), .B1(n12393), .B2(n13201), .ZN(
        n12395) );
  NAND3_X1 U14730 ( .A1(n12397), .A2(n12396), .A3(n12395), .ZN(n12398) );
  OAI211_X1 U14731 ( .C1(n12400), .C2(n14782), .A(n12399), .B(n12398), .ZN(
        P2_U3203) );
  NAND2_X1 U14732 ( .A1(n14138), .A2(n12441), .ZN(n12402) );
  NAND2_X1 U14733 ( .A1(n13825), .A2(n12424), .ZN(n12401) );
  NAND2_X1 U14734 ( .A1(n12402), .A2(n12401), .ZN(n12403) );
  XNOR2_X1 U14735 ( .A(n12403), .B(n6519), .ZN(n12405) );
  AND2_X1 U14736 ( .A1(n13825), .A2(n12446), .ZN(n12404) );
  AOI21_X1 U14737 ( .B1(n14138), .B2(n12424), .A(n12404), .ZN(n12406) );
  NAND2_X1 U14738 ( .A1(n12405), .A2(n12406), .ZN(n13747) );
  INV_X1 U14739 ( .A(n12405), .ZN(n12408) );
  INV_X1 U14740 ( .A(n12406), .ZN(n12407) );
  NAND2_X1 U14741 ( .A1(n12408), .A2(n12407), .ZN(n12409) );
  AND2_X1 U14742 ( .A1(n13747), .A2(n12409), .ZN(n13668) );
  NAND2_X1 U14743 ( .A1(n13671), .A2(n13747), .ZN(n12419) );
  NAND2_X1 U14744 ( .A1(n14133), .A2(n12441), .ZN(n12411) );
  NAND2_X1 U14745 ( .A1(n13824), .A2(n12424), .ZN(n12410) );
  NAND2_X1 U14746 ( .A1(n12411), .A2(n12410), .ZN(n12412) );
  XNOR2_X1 U14747 ( .A(n12412), .B(n6519), .ZN(n12414) );
  AND2_X1 U14748 ( .A1(n13824), .A2(n12446), .ZN(n12413) );
  AOI21_X1 U14749 ( .B1(n14133), .B2(n10922), .A(n12413), .ZN(n12415) );
  NAND2_X1 U14750 ( .A1(n12414), .A2(n12415), .ZN(n13697) );
  INV_X1 U14751 ( .A(n12414), .ZN(n12417) );
  INV_X1 U14752 ( .A(n12415), .ZN(n12416) );
  NAND2_X1 U14753 ( .A1(n12417), .A2(n12416), .ZN(n12418) );
  AND2_X1 U14754 ( .A1(n13697), .A2(n12418), .ZN(n13748) );
  NAND2_X1 U14755 ( .A1(n12419), .A2(n13748), .ZN(n13696) );
  NAND2_X1 U14756 ( .A1(n13696), .A2(n13697), .ZN(n12430) );
  NAND2_X1 U14757 ( .A1(n14125), .A2(n12441), .ZN(n12421) );
  NAND2_X1 U14758 ( .A1(n13823), .A2(n10922), .ZN(n12420) );
  NAND2_X1 U14759 ( .A1(n12421), .A2(n12420), .ZN(n12422) );
  XNOR2_X1 U14760 ( .A(n12422), .B(n6519), .ZN(n12425) );
  AND2_X1 U14761 ( .A1(n13823), .A2(n12446), .ZN(n12423) );
  AOI21_X1 U14762 ( .B1(n14125), .B2(n12424), .A(n12423), .ZN(n12426) );
  NAND2_X1 U14763 ( .A1(n12425), .A2(n12426), .ZN(n12431) );
  INV_X1 U14764 ( .A(n12425), .ZN(n12428) );
  INV_X1 U14765 ( .A(n12426), .ZN(n12427) );
  NAND2_X1 U14766 ( .A1(n12428), .A2(n12427), .ZN(n12429) );
  AND2_X1 U14767 ( .A1(n12431), .A2(n12429), .ZN(n13698) );
  NAND2_X1 U14768 ( .A1(n12430), .A2(n13698), .ZN(n13700) );
  NAND2_X1 U14769 ( .A1(n13967), .A2(n12441), .ZN(n12433) );
  NAND2_X1 U14770 ( .A1(n13822), .A2(n10922), .ZN(n12432) );
  NAND2_X1 U14771 ( .A1(n12433), .A2(n12432), .ZN(n12434) );
  XNOR2_X1 U14772 ( .A(n12434), .B(n12444), .ZN(n12438) );
  NAND2_X1 U14773 ( .A1(n13967), .A2(n12424), .ZN(n12436) );
  NAND2_X1 U14774 ( .A1(n13822), .A2(n12446), .ZN(n12435) );
  NAND2_X1 U14775 ( .A1(n12436), .A2(n12435), .ZN(n12437) );
  NOR2_X1 U14776 ( .A1(n12438), .A2(n12437), .ZN(n12439) );
  AOI21_X1 U14777 ( .B1(n12438), .B2(n12437), .A(n12439), .ZN(n13794) );
  NAND2_X1 U14778 ( .A1(n13793), .A2(n13794), .ZN(n13792) );
  INV_X1 U14779 ( .A(n12439), .ZN(n12440) );
  NAND2_X1 U14780 ( .A1(n14112), .A2(n12441), .ZN(n12443) );
  NAND2_X1 U14781 ( .A1(n13956), .A2(n10922), .ZN(n12442) );
  NAND2_X1 U14782 ( .A1(n12443), .A2(n12442), .ZN(n12445) );
  XNOR2_X1 U14783 ( .A(n12445), .B(n12444), .ZN(n12450) );
  NAND2_X1 U14784 ( .A1(n14112), .A2(n10922), .ZN(n12448) );
  NAND2_X1 U14785 ( .A1(n13956), .A2(n12446), .ZN(n12447) );
  NAND2_X1 U14786 ( .A1(n12448), .A2(n12447), .ZN(n12449) );
  NOR2_X1 U14787 ( .A1(n12450), .A2(n12449), .ZN(n12451) );
  AOI21_X1 U14788 ( .B1(n12450), .B2(n12449), .A(n12451), .ZN(n13659) );
  NAND2_X1 U14789 ( .A1(n13658), .A2(n13659), .ZN(n13657) );
  INV_X1 U14790 ( .A(n13821), .ZN(n13662) );
  OAI22_X1 U14791 ( .A1(n12478), .A2(n12453), .B1(n13662), .B2(n12452), .ZN(
        n12457) );
  OAI22_X1 U14792 ( .A1(n12478), .A2(n12454), .B1(n13662), .B2(n12453), .ZN(
        n12455) );
  XNOR2_X1 U14793 ( .A(n12455), .B(n12444), .ZN(n12456) );
  XOR2_X1 U14794 ( .A(n12457), .B(n12456), .Z(n12458) );
  INV_X1 U14795 ( .A(n12459), .ZN(n12460) );
  AOI22_X1 U14796 ( .A1(n12460), .A2(n13798), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12462) );
  NAND2_X1 U14797 ( .A1(n13820), .A2(n13810), .ZN(n12461) );
  OAI211_X1 U14798 ( .C1(n12463), .C2(n13808), .A(n12462), .B(n12461), .ZN(
        n12464) );
  AOI21_X1 U14799 ( .B1(n14104), .B2(n13815), .A(n12464), .ZN(n12465) );
  INV_X1 U14800 ( .A(n12466), .ZN(n12467) );
  NAND2_X1 U14801 ( .A1(n14400), .A2(n12467), .ZN(n12765) );
  OAI21_X1 U14802 ( .B1(n15117), .B2(n12468), .A(n12765), .ZN(n12471) );
  NOR2_X1 U14803 ( .A1(n12469), .A2(n12902), .ZN(n12470) );
  AOI211_X1 U14804 ( .C1(n14402), .C2(n12472), .A(n12471), .B(n12470), .ZN(
        n12473) );
  OAI21_X1 U14805 ( .B1(n12474), .B2(n15119), .A(n12473), .ZN(P3_U3204) );
  XNOR2_X2 U14806 ( .A(n12477), .B(n12476), .ZN(n14103) );
  NOR2_X1 U14807 ( .A1(n12478), .A2(n13821), .ZN(n12479) );
  OAI22_X1 U14808 ( .A1(n12480), .A2(n12479), .B1(n13662), .B2(n14104), .ZN(
        n12482) );
  XNOR2_X1 U14809 ( .A(n12482), .B(n12476), .ZN(n14095) );
  NAND2_X1 U14810 ( .A1(n14095), .A2(n14035), .ZN(n12498) );
  AOI21_X1 U14811 ( .B1(n14096), .B2(n12483), .A(n14699), .ZN(n12486) );
  INV_X1 U14812 ( .A(n14096), .ZN(n12485) );
  INV_X1 U14813 ( .A(n12483), .ZN(n12484) );
  NAND2_X1 U14814 ( .A1(n13821), .A2(n14482), .ZN(n14097) );
  NAND2_X1 U14815 ( .A1(n14096), .A2(n14677), .ZN(n12495) );
  INV_X1 U14816 ( .A(n12487), .ZN(n12493) );
  INV_X1 U14817 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n12491) );
  NOR2_X1 U14818 ( .A1(n14206), .A2(n12488), .ZN(n12489) );
  NOR2_X1 U14819 ( .A1(n14055), .A2(n12489), .ZN(n13931) );
  NAND2_X1 U14820 ( .A1(n13819), .A2(n13931), .ZN(n14098) );
  OAI22_X1 U14821 ( .A1(n14665), .A2(n12491), .B1(n14098), .B2(n12490), .ZN(
        n12492) );
  AOI21_X1 U14822 ( .B1(n12493), .B2(n14643), .A(n12492), .ZN(n12494) );
  OAI211_X1 U14823 ( .C1(n14644), .C2(n14097), .A(n12495), .B(n12494), .ZN(
        n12496) );
  AOI21_X1 U14824 ( .B1(n14100), .B2(n14683), .A(n12496), .ZN(n12497) );
  OAI211_X1 U14825 ( .C1(n14103), .C2(n14083), .A(n12498), .B(n12497), .ZN(
        P1_U3356) );
  XNOR2_X1 U14826 ( .A(n13581), .B(n6725), .ZN(n12515) );
  NAND2_X1 U14827 ( .A1(n13249), .A2(n13105), .ZN(n12516) );
  XNOR2_X1 U14828 ( .A(n13586), .B(n13134), .ZN(n12514) );
  NAND2_X1 U14829 ( .A1(n13250), .A2(n13105), .ZN(n12513) );
  NOR2_X1 U14830 ( .A1(n13219), .A2(n13523), .ZN(n13124) );
  XNOR2_X1 U14831 ( .A(n13607), .B(n13134), .ZN(n12504) );
  NAND2_X1 U14832 ( .A1(n13254), .A2(n13105), .ZN(n12503) );
  NAND2_X1 U14833 ( .A1(n12504), .A2(n12503), .ZN(n12505) );
  OAI21_X1 U14834 ( .B1(n12504), .B2(n12503), .A(n12505), .ZN(n13175) );
  XNOR2_X1 U14835 ( .A(n13600), .B(n13134), .ZN(n12507) );
  NAND2_X1 U14836 ( .A1(n13253), .A2(n13105), .ZN(n12506) );
  NAND2_X1 U14837 ( .A1(n12507), .A2(n12506), .ZN(n12508) );
  OAI21_X1 U14838 ( .B1(n12507), .B2(n12506), .A(n12508), .ZN(n13183) );
  INV_X1 U14839 ( .A(n12508), .ZN(n12509) );
  XNOR2_X1 U14840 ( .A(n13595), .B(n6725), .ZN(n12511) );
  NAND2_X1 U14841 ( .A1(n13252), .A2(n13105), .ZN(n12510) );
  XNOR2_X1 U14842 ( .A(n12511), .B(n12510), .ZN(n13216) );
  INV_X1 U14843 ( .A(n12510), .ZN(n12512) );
  XNOR2_X1 U14844 ( .A(n12514), .B(n12513), .ZN(n13205) );
  XNOR2_X1 U14845 ( .A(n13591), .B(n6725), .ZN(n13123) );
  NAND2_X1 U14846 ( .A1(n13123), .A2(n13124), .ZN(n13122) );
  XNOR2_X1 U14847 ( .A(n12515), .B(n12516), .ZN(n13152) );
  XNOR2_X1 U14848 ( .A(n13575), .B(n6725), .ZN(n13081) );
  NAND2_X1 U14849 ( .A1(n13248), .A2(n13489), .ZN(n12518) );
  NOR2_X2 U14850 ( .A1(n12519), .A2(n12518), .ZN(n13084) );
  INV_X1 U14851 ( .A(n12519), .ZN(n12520) );
  AOI22_X1 U14852 ( .A1(n12520), .A2(n14428), .B1(n13225), .B2(n13248), .ZN(
        n12525) );
  AND2_X1 U14853 ( .A1(n13249), .A2(n13231), .ZN(n12521) );
  AOI21_X1 U14854 ( .B1(n13247), .B2(n13233), .A(n12521), .ZN(n13426) );
  AOI22_X1 U14855 ( .A1(n13208), .A2(n13431), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12522) );
  OAI21_X1 U14856 ( .B1(n13426), .B2(n14779), .A(n12522), .ZN(n12523) );
  AOI21_X1 U14857 ( .B1(n13575), .B2(n14787), .A(n12523), .ZN(n12524) );
  OAI21_X1 U14858 ( .B1(n13084), .B2(n12525), .A(n12524), .ZN(P2_U3207) );
  OAI222_X1 U14859 ( .A1(n14214), .A2(n9665), .B1(n12527), .B2(P1_U3086), .C1(
        n12526), .C2(n12044), .ZN(P1_U3325) );
  XNOR2_X1 U14860 ( .A(n12771), .B(n12528), .ZN(n12535) );
  INV_X1 U14861 ( .A(n12535), .ZN(n12529) );
  NAND2_X1 U14862 ( .A1(n12529), .A2(n12642), .ZN(n12541) );
  INV_X1 U14863 ( .A(n12530), .ZN(n12531) );
  AOI22_X1 U14864 ( .A1(n10675), .A2(n12774), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12533) );
  NAND2_X1 U14865 ( .A1(n12552), .A2(n12773), .ZN(n12532) );
  OAI211_X1 U14866 ( .C1(n12645), .C2(n12777), .A(n12533), .B(n12532), .ZN(
        n12537) );
  NOR4_X1 U14867 ( .A1(n12535), .A2(n12637), .A3(n12534), .A4(n12773), .ZN(
        n12536) );
  AOI211_X1 U14868 ( .C1(n12634), .C2(n12538), .A(n12537), .B(n12536), .ZN(
        n12539) );
  INV_X1 U14869 ( .A(n12542), .ZN(n12543) );
  OAI222_X1 U14870 ( .A1(n8353), .A2(P3_U3151), .B1(n13076), .B2(n12543), .C1(
        n15229), .C2(n13078), .ZN(P3_U3265) );
  NAND2_X1 U14871 ( .A1(n12544), .A2(n12545), .ZN(n12546) );
  XOR2_X1 U14872 ( .A(n12547), .B(n12546), .Z(n12548) );
  NAND2_X1 U14873 ( .A1(n12548), .A2(n12642), .ZN(n12554) );
  INV_X1 U14874 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n15238) );
  OAI22_X1 U14875 ( .A1(n12608), .A2(n12926), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15238), .ZN(n12551) );
  NOR2_X1 U14876 ( .A1(n12645), .A2(n12549), .ZN(n12550) );
  AOI211_X1 U14877 ( .C1(n12552), .C2(n12664), .A(n12551), .B(n12550), .ZN(
        n12553) );
  OAI211_X1 U14878 ( .C1(n12649), .C2(n12555), .A(n12554), .B(n12553), .ZN(
        P3_U3155) );
  INV_X1 U14879 ( .A(n12556), .ZN(n12604) );
  AOI22_X1 U14880 ( .A1(n12654), .A2(n10675), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12558) );
  NAND2_X1 U14881 ( .A1(n12629), .A2(n12846), .ZN(n12557) );
  OAI211_X1 U14882 ( .C1(n9831), .C2(n12632), .A(n12558), .B(n12557), .ZN(
        n12559) );
  AOI21_X1 U14883 ( .B1(n12966), .B2(n12634), .A(n12559), .ZN(n12560) );
  OAI21_X1 U14884 ( .B1(n12561), .B2(n12637), .A(n12560), .ZN(P3_U3156) );
  XNOR2_X1 U14885 ( .A(n12562), .B(n12563), .ZN(n12568) );
  NAND2_X1 U14886 ( .A1(n10675), .A2(n12887), .ZN(n12564) );
  NAND2_X1 U14887 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12760)
         );
  OAI211_X1 U14888 ( .C1(n12632), .C2(n12911), .A(n12564), .B(n12760), .ZN(
        n12566) );
  NOR2_X1 U14889 ( .A1(n13047), .A2(n12649), .ZN(n12565) );
  AOI211_X1 U14890 ( .C1(n12890), .C2(n12629), .A(n12566), .B(n12565), .ZN(
        n12567) );
  OAI21_X1 U14891 ( .B1(n12568), .B2(n12637), .A(n12567), .ZN(P3_U3159) );
  INV_X1 U14892 ( .A(n12569), .ZN(n12570) );
  AOI21_X1 U14893 ( .B1(n12572), .B2(n12571), .A(n12570), .ZN(n12577) );
  NAND2_X1 U14894 ( .A1(n12629), .A2(n12866), .ZN(n12574) );
  AOI22_X1 U14895 ( .A1(n12656), .A2(n10675), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12573) );
  OAI211_X1 U14896 ( .C1(n12862), .C2(n12632), .A(n12574), .B(n12573), .ZN(
        n12575) );
  AOI21_X1 U14897 ( .B1(n12865), .B2(n12634), .A(n12575), .ZN(n12576) );
  OAI21_X1 U14898 ( .B1(n12577), .B2(n12637), .A(n12576), .ZN(P3_U3163) );
  INV_X1 U14899 ( .A(n12579), .ZN(n12605) );
  INV_X1 U14900 ( .A(n12580), .ZN(n12582) );
  NOR3_X1 U14901 ( .A1(n12605), .A2(n12582), .A3(n12581), .ZN(n12585) );
  INV_X1 U14902 ( .A(n12583), .ZN(n12584) );
  OAI21_X1 U14903 ( .B1(n12585), .B2(n12584), .A(n12642), .ZN(n12589) );
  AOI22_X1 U14904 ( .A1(n10675), .A2(n12652), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12586) );
  OAI21_X1 U14905 ( .B1(n12842), .B2(n12632), .A(n12586), .ZN(n12587) );
  AOI21_X1 U14906 ( .B1(n12817), .B2(n12629), .A(n12587), .ZN(n12588) );
  OAI211_X1 U14907 ( .C1(n13026), .C2(n12649), .A(n12589), .B(n12588), .ZN(
        P3_U3165) );
  OR2_X1 U14908 ( .A1(n12121), .A2(n12590), .ZN(n12592) );
  NAND2_X1 U14909 ( .A1(n12592), .A2(n12591), .ZN(n12594) );
  XNOR2_X1 U14910 ( .A(n12594), .B(n12593), .ZN(n12600) );
  NAND2_X1 U14911 ( .A1(n12629), .A2(n12915), .ZN(n12596) );
  AOI22_X1 U14912 ( .A1(n10675), .A2(n12886), .B1(P3_REG3_REG_17__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12595) );
  OAI211_X1 U14913 ( .C1(n12912), .C2(n12632), .A(n12596), .B(n12595), .ZN(
        n12597) );
  AOI21_X1 U14914 ( .B1(n12598), .B2(n12634), .A(n12597), .ZN(n12599) );
  OAI21_X1 U14915 ( .B1(n12600), .B2(n12637), .A(n12599), .ZN(P3_U3168) );
  INV_X1 U14916 ( .A(n12834), .ZN(n13030) );
  INV_X1 U14917 ( .A(n12601), .ZN(n12603) );
  NOR3_X1 U14918 ( .A1(n12604), .A2(n12603), .A3(n12602), .ZN(n12606) );
  OAI21_X1 U14919 ( .B1(n12606), .B2(n12605), .A(n12642), .ZN(n12612) );
  NOR2_X1 U14920 ( .A1(n12828), .A2(n12632), .ZN(n12610) );
  OAI22_X1 U14921 ( .A1(n12829), .A2(n12608), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12607), .ZN(n12609) );
  AOI211_X1 U14922 ( .C1(n12833), .C2(n12629), .A(n12610), .B(n12609), .ZN(
        n12611) );
  OAI211_X1 U14923 ( .C1(n13030), .C2(n12649), .A(n12612), .B(n12611), .ZN(
        P3_U3169) );
  XNOR2_X1 U14924 ( .A(n12613), .B(n12614), .ZN(n12619) );
  NAND2_X1 U14925 ( .A1(n12629), .A2(n12878), .ZN(n12616) );
  AOI22_X1 U14926 ( .A1(n12657), .A2(n10675), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12615) );
  OAI211_X1 U14927 ( .C1(n12899), .C2(n12632), .A(n12616), .B(n12615), .ZN(
        n12617) );
  AOI21_X1 U14928 ( .B1(n12877), .B2(n12634), .A(n12617), .ZN(n12618) );
  OAI21_X1 U14929 ( .B1(n12619), .B2(n12637), .A(n12618), .ZN(P3_U3173) );
  AOI21_X1 U14930 ( .B1(n12656), .B2(n12620), .A(n6573), .ZN(n12626) );
  INV_X1 U14931 ( .A(n12856), .ZN(n12622) );
  OAI22_X1 U14932 ( .A1(n12828), .A2(n12925), .B1(n12874), .B2(n12927), .ZN(
        n12852) );
  AOI22_X1 U14933 ( .A1(n12852), .A2(n12647), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12621) );
  OAI21_X1 U14934 ( .B1(n12622), .B2(n12645), .A(n12621), .ZN(n12623) );
  AOI21_X1 U14935 ( .B1(n12624), .B2(n12634), .A(n12623), .ZN(n12625) );
  OAI21_X1 U14936 ( .B1(n12626), .B2(n12637), .A(n12625), .ZN(P3_U3175) );
  XNOR2_X1 U14937 ( .A(n12627), .B(n12628), .ZN(n12638) );
  NAND2_X1 U14938 ( .A1(n12629), .A2(n12904), .ZN(n12631) );
  AOI22_X1 U14939 ( .A1(n10675), .A2(n12659), .B1(P3_REG3_REG_18__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12630) );
  OAI211_X1 U14940 ( .C1(n12924), .C2(n12632), .A(n12631), .B(n12630), .ZN(
        n12633) );
  AOI21_X1 U14941 ( .B1(n12635), .B2(n12634), .A(n12633), .ZN(n12636) );
  OAI21_X1 U14942 ( .B1(n12638), .B2(n12637), .A(n12636), .ZN(P3_U3178) );
  OAI21_X1 U14943 ( .B1(n12641), .B2(n12640), .A(n12639), .ZN(n12643) );
  OAI22_X1 U14944 ( .A1(n12829), .A2(n12927), .B1(n12644), .B2(n12925), .ZN(
        n12797) );
  OAI22_X1 U14945 ( .A1(n12645), .A2(n12802), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15325), .ZN(n12646) );
  AOI21_X1 U14946 ( .B1(n12797), .B2(n12647), .A(n12646), .ZN(n12648) );
  MUX2_X1 U14947 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12763), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14948 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(n12650), .S(P3_U3897), .Z(
        P3_U3521) );
  MUX2_X1 U14949 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n12774), .S(P3_U3897), .Z(
        P3_U3520) );
  MUX2_X1 U14950 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12651), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14951 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12773), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14952 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12652), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14953 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12653), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14954 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12654), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14955 ( .A(n12655), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12658), .Z(
        P3_U3514) );
  MUX2_X1 U14956 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12656), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14957 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12657), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14958 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12887), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14959 ( .A(n12659), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12658), .Z(
        P3_U3510) );
  MUX2_X1 U14960 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12886), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14961 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12660), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14962 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12661), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14963 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12662), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14964 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12663), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14965 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12664), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14966 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12665), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14967 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12666), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14968 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12667), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14969 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n12668), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U14970 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12669), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14971 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12670), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14972 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12671), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14973 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12672), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14974 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12673), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14975 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n15091), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14976 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n9772), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14977 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n9764), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U14978 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n8497), .S(P3_U3897), .Z(
        P3_U3491) );
  NOR2_X1 U14979 ( .A1(n12688), .A2(n12675), .ZN(n12677) );
  NAND2_X1 U14980 ( .A1(n12700), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12715) );
  OAI21_X1 U14981 ( .B1(n12700), .B2(P3_REG2_REG_14__SCAN_IN), .A(n12715), 
        .ZN(n12690) );
  AOI21_X1 U14982 ( .B1(n12678), .B2(n12690), .A(n12705), .ZN(n12704) );
  NAND2_X1 U14983 ( .A1(n12680), .A2(n12679), .ZN(n12682) );
  NAND2_X1 U14984 ( .A1(n12682), .A2(n12681), .ZN(n12686) );
  INV_X1 U14985 ( .A(n12700), .ZN(n12684) );
  NAND2_X1 U14986 ( .A1(n12684), .A2(n12683), .ZN(n12685) );
  NAND2_X1 U14987 ( .A1(n12700), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12714) );
  AND2_X1 U14988 ( .A1(n12685), .A2(n12714), .ZN(n12692) );
  NAND2_X1 U14989 ( .A1(n12692), .A2(n12686), .ZN(n12708) );
  OAI21_X1 U14990 ( .B1(n12686), .B2(n12692), .A(n12708), .ZN(n12702) );
  INV_X1 U14991 ( .A(n12687), .ZN(n12689) );
  NAND2_X1 U14992 ( .A1(n12689), .A2(n12688), .ZN(n12693) );
  AND2_X1 U14993 ( .A1(n12694), .A2(n12693), .ZN(n12696) );
  INV_X1 U14994 ( .A(n12690), .ZN(n12691) );
  MUX2_X1 U14995 ( .A(n12692), .B(n12691), .S(n14348), .Z(n12695) );
  NAND3_X1 U14996 ( .A1(n12694), .A2(n12693), .A3(n12695), .ZN(n12717) );
  OAI211_X1 U14997 ( .C1(n12696), .C2(n12695), .A(n15078), .B(n12717), .ZN(
        n12699) );
  NOR2_X1 U14998 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15238), .ZN(n12697) );
  AOI21_X1 U14999 ( .B1(n15068), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12697), 
        .ZN(n12698) );
  OAI211_X1 U15000 ( .C1(n15052), .C2(n12700), .A(n12699), .B(n12698), .ZN(
        n12701) );
  AOI21_X1 U15001 ( .B1(n15069), .B2(n12702), .A(n12701), .ZN(n12703) );
  OAI21_X1 U15002 ( .B1(n12704), .B2(n15063), .A(n12703), .ZN(P3_U3196) );
  XNOR2_X1 U15003 ( .A(n12750), .B(n12724), .ZN(n12706) );
  AOI21_X1 U15004 ( .B1(n12707), .B2(n12706), .A(n12725), .ZN(n12723) );
  NAND2_X1 U15005 ( .A1(n12714), .A2(n12708), .ZN(n12749) );
  XNOR2_X1 U15006 ( .A(n12735), .B(n12749), .ZN(n12709) );
  NAND2_X1 U15007 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n12709), .ZN(n12751) );
  OAI21_X1 U15008 ( .B1(n12709), .B2(P3_REG1_REG_15__SCAN_IN), .A(n12751), 
        .ZN(n12713) );
  INV_X1 U15009 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n12710) );
  INV_X1 U15010 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n15227) );
  OAI22_X1 U15011 ( .A1(n15043), .A2(n12710), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15227), .ZN(n12712) );
  NOR2_X1 U15012 ( .A1(n15052), .A2(n12750), .ZN(n12711) );
  AOI211_X1 U15013 ( .C1(n15069), .C2(n12713), .A(n12712), .B(n12711), .ZN(
        n12722) );
  NAND2_X1 U15014 ( .A1(n12717), .A2(n12716), .ZN(n12733) );
  XNOR2_X1 U15015 ( .A(n12733), .B(n12750), .ZN(n12719) );
  NOR2_X1 U15016 ( .A1(n12719), .A2(n12718), .ZN(n12734) );
  AND2_X1 U15017 ( .A1(n12719), .A2(n12718), .ZN(n12720) );
  OAI21_X1 U15018 ( .B1(n12734), .B2(n12720), .A(n15078), .ZN(n12721) );
  OAI211_X1 U15019 ( .C1(n12723), .C2(n15063), .A(n12722), .B(n12721), .ZN(
        P3_U3197) );
  AND2_X1 U15020 ( .A1(n12750), .A2(n12724), .ZN(n12726) );
  NAND2_X1 U15021 ( .A1(n12738), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n12729) );
  NAND2_X1 U15022 ( .A1(n14347), .A2(n12727), .ZN(n12728) );
  NAND2_X1 U15023 ( .A1(n12729), .A2(n12728), .ZN(n14359) );
  INV_X1 U15024 ( .A(n12729), .ZN(n14349) );
  NOR2_X1 U15025 ( .A1(n14365), .A2(n12730), .ZN(n12731) );
  AOI22_X1 U15026 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n14380), .B1(n12748), 
        .B2(n8471), .ZN(n14390) );
  XNOR2_X1 U15027 ( .A(n8454), .B(n12732), .ZN(n12744) );
  INV_X1 U15028 ( .A(n12740), .ZN(n12741) );
  INV_X1 U15029 ( .A(n12733), .ZN(n12736) );
  AOI21_X1 U15030 ( .B1(n12738), .B2(n12737), .A(n14353), .ZN(n12739) );
  NOR2_X1 U15031 ( .A1(n12738), .A2(n12737), .ZN(n14351) );
  XNOR2_X1 U15032 ( .A(n14365), .B(n12740), .ZN(n14369) );
  NAND2_X1 U15033 ( .A1(n14370), .A2(n14369), .ZN(n14368) );
  OAI21_X1 U15034 ( .B1(n14365), .B2(n12741), .A(n14368), .ZN(n12742) );
  INV_X1 U15035 ( .A(n12742), .ZN(n12743) );
  XNOR2_X1 U15036 ( .A(n12742), .B(n12748), .ZN(n14382) );
  NOR2_X1 U15037 ( .A1(n14382), .A2(n14383), .ZN(n14381) );
  AOI21_X1 U15038 ( .B1(n12743), .B2(n14380), .A(n14381), .ZN(n12747) );
  XNOR2_X1 U15039 ( .A(n8454), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12757) );
  INV_X1 U15040 ( .A(n12744), .ZN(n12745) );
  MUX2_X1 U15041 ( .A(n12757), .B(n12745), .S(n14348), .Z(n12746) );
  XNOR2_X1 U15042 ( .A(n12747), .B(n12746), .ZN(n12762) );
  INV_X1 U15043 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12993) );
  AOI22_X1 U15044 ( .A1(P3_REG1_REG_18__SCAN_IN), .A2(n12748), .B1(n14380), 
        .B2(n12993), .ZN(n14387) );
  NAND2_X1 U15045 ( .A1(n12750), .A2(n12749), .ZN(n12752) );
  NAND2_X1 U15046 ( .A1(n12752), .A2(n12751), .ZN(n14356) );
  XNOR2_X1 U15047 ( .A(n14347), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n14355) );
  NOR2_X1 U15048 ( .A1(n14347), .A2(n13001), .ZN(n14350) );
  AOI21_X1 U15049 ( .B1(n14356), .B2(n14355), .A(n14350), .ZN(n12753) );
  NAND2_X1 U15050 ( .A1(n12755), .A2(n12754), .ZN(n12756) );
  NAND2_X1 U15051 ( .A1(n14387), .A2(n14386), .ZN(n14385) );
  OAI21_X1 U15052 ( .B1(n14380), .B2(n12993), .A(n14385), .ZN(n12758) );
  NAND2_X1 U15053 ( .A1(n15068), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12759) );
  OAI211_X1 U15054 ( .C1(n15052), .C2(n8454), .A(n12760), .B(n12759), .ZN(
        n12761) );
  NAND2_X1 U15055 ( .A1(n12764), .A2(n12763), .ZN(n13008) );
  OAI21_X1 U15056 ( .B1(n15119), .B2(n13008), .A(n12765), .ZN(n12767) );
  AOI21_X1 U15057 ( .B1(P3_REG2_REG_31__SCAN_IN), .B2(n15119), .A(n12767), 
        .ZN(n12766) );
  OAI21_X1 U15058 ( .B1(n13010), .B2(n12933), .A(n12766), .ZN(P3_U3202) );
  AOI21_X1 U15059 ( .B1(P3_REG2_REG_30__SCAN_IN), .B2(n15119), .A(n12767), 
        .ZN(n12768) );
  OAI21_X1 U15060 ( .B1(n13013), .B2(n12933), .A(n12768), .ZN(P3_U3203) );
  XOR2_X1 U15061 ( .A(n12771), .B(n12769), .Z(n12946) );
  INV_X1 U15062 ( .A(n12946), .ZN(n12782) );
  OAI211_X1 U15063 ( .C1(n12772), .C2(n12771), .A(n12770), .B(n15106), .ZN(
        n12776) );
  AOI22_X1 U15064 ( .A1(n15104), .A2(n12774), .B1(n12773), .B2(n15103), .ZN(
        n12775) );
  NAND2_X1 U15065 ( .A1(n12776), .A2(n12775), .ZN(n12945) );
  NOR2_X1 U15066 ( .A1(n13017), .A2(n12933), .ZN(n12780) );
  OAI22_X1 U15067 ( .A1(n15117), .A2(n12778), .B1(n12777), .B2(n15112), .ZN(
        n12779) );
  AOI211_X1 U15068 ( .C1(n12945), .C2(n15117), .A(n12780), .B(n12779), .ZN(
        n12781) );
  OAI21_X1 U15069 ( .B1(n12782), .B2(n12902), .A(n12781), .ZN(P3_U3205) );
  XOR2_X1 U15070 ( .A(n12785), .B(n12783), .Z(n12784) );
  XNOR2_X1 U15071 ( .A(n12786), .B(n12785), .ZN(n12793) );
  INV_X1 U15072 ( .A(n12787), .ZN(n12788) );
  OAI22_X1 U15073 ( .A1(n15117), .A2(n12792), .B1(n12791), .B2(n15112), .ZN(
        n12795) );
  INV_X1 U15074 ( .A(n12793), .ZN(n12952) );
  NOR2_X1 U15075 ( .A1(n12952), .A2(n15114), .ZN(n12794) );
  AOI211_X1 U15076 ( .C1(n14402), .C2(n12949), .A(n12795), .B(n12794), .ZN(
        n12796) );
  OAI21_X1 U15077 ( .B1(n12951), .B2(n15119), .A(n12796), .ZN(P3_U3206) );
  XNOR2_X1 U15078 ( .A(n6536), .B(n12800), .ZN(n12799) );
  INV_X1 U15079 ( .A(n12797), .ZN(n12798) );
  OAI21_X1 U15080 ( .B1(n12799), .B2(n12922), .A(n12798), .ZN(n12953) );
  INV_X1 U15081 ( .A(n12953), .ZN(n12807) );
  XNOR2_X1 U15082 ( .A(n12801), .B(n12800), .ZN(n12954) );
  NOR2_X1 U15083 ( .A1(n13022), .A2(n12933), .ZN(n12805) );
  OAI22_X1 U15084 ( .A1(n15117), .A2(n12803), .B1(n12802), .B2(n15112), .ZN(
        n12804) );
  AOI211_X1 U15085 ( .C1(n12954), .C2(n12935), .A(n12805), .B(n12804), .ZN(
        n12806) );
  OAI21_X1 U15086 ( .B1(n12807), .B2(n15119), .A(n12806), .ZN(P3_U3207) );
  OR2_X1 U15087 ( .A1(n12808), .A2(n12813), .ZN(n12809) );
  NAND2_X1 U15088 ( .A1(n12810), .A2(n12809), .ZN(n12958) );
  OAI22_X1 U15089 ( .A1(n12842), .A2(n12927), .B1(n12811), .B2(n12925), .ZN(
        n12814) );
  NAND2_X1 U15090 ( .A1(n12958), .A2(n12816), .ZN(n12819) );
  AOI22_X1 U15091 ( .A1(n12817), .A2(n14400), .B1(n15119), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12818) );
  OAI211_X1 U15092 ( .C1(n13026), .C2(n12933), .A(n12819), .B(n12818), .ZN(
        n12820) );
  AOI21_X1 U15093 ( .B1(n12957), .B2(n15117), .A(n12820), .ZN(n12821) );
  INV_X1 U15094 ( .A(n12821), .ZN(P3_U3208) );
  NAND2_X1 U15095 ( .A1(n12822), .A2(n12826), .ZN(n12823) );
  OAI21_X1 U15096 ( .B1(n12827), .B2(n12826), .A(n12825), .ZN(n12831) );
  OAI22_X1 U15097 ( .A1(n12829), .A2(n12925), .B1(n12828), .B2(n12927), .ZN(
        n12830) );
  AOI21_X1 U15098 ( .B1(n12831), .B2(n15106), .A(n12830), .ZN(n12832) );
  OAI21_X1 U15099 ( .B1(n15110), .B2(n12961), .A(n12832), .ZN(n12962) );
  AOI22_X1 U15100 ( .A1(n12833), .A2(n14400), .B1(n15119), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n12836) );
  NAND2_X1 U15101 ( .A1(n12834), .A2(n14402), .ZN(n12835) );
  OAI211_X1 U15102 ( .C1(n12961), .C2(n15114), .A(n12836), .B(n12835), .ZN(
        n12837) );
  AOI21_X1 U15103 ( .B1(n12962), .B2(n15117), .A(n12837), .ZN(n12838) );
  INV_X1 U15104 ( .A(n12838), .ZN(P3_U3209) );
  XNOR2_X1 U15105 ( .A(n12839), .B(n12840), .ZN(n12967) );
  XNOR2_X1 U15106 ( .A(n12841), .B(n12840), .ZN(n12844) );
  OAI22_X1 U15107 ( .A1(n12842), .A2(n12925), .B1(n9831), .B2(n12927), .ZN(
        n12843) );
  AOI21_X1 U15108 ( .B1(n12844), .B2(n15106), .A(n12843), .ZN(n12845) );
  OAI21_X1 U15109 ( .B1(n15110), .B2(n12967), .A(n12845), .ZN(n12968) );
  AOI22_X1 U15110 ( .A1(n12846), .A2(n14400), .B1(n15119), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n12848) );
  NAND2_X1 U15111 ( .A1(n12966), .A2(n14402), .ZN(n12847) );
  OAI211_X1 U15112 ( .C1(n12967), .C2(n15114), .A(n12848), .B(n12847), .ZN(
        n12849) );
  AOI21_X1 U15113 ( .B1(n12968), .B2(n15117), .A(n12849), .ZN(n12850) );
  INV_X1 U15114 ( .A(n12850), .ZN(P3_U3210) );
  XNOR2_X1 U15115 ( .A(n12851), .B(n12854), .ZN(n12853) );
  AOI21_X1 U15116 ( .B1(n12853), .B2(n15106), .A(n12852), .ZN(n12974) );
  XNOR2_X1 U15117 ( .A(n12855), .B(n12854), .ZN(n12972) );
  AOI22_X1 U15118 ( .A1(n15119), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n14400), 
        .B2(n12856), .ZN(n12857) );
  OAI21_X1 U15119 ( .B1(n12975), .B2(n12933), .A(n12857), .ZN(n12858) );
  AOI21_X1 U15120 ( .B1(n12972), .B2(n12935), .A(n12858), .ZN(n12859) );
  OAI21_X1 U15121 ( .B1(n12974), .B2(n15119), .A(n12859), .ZN(P3_U3211) );
  XNOR2_X1 U15122 ( .A(n12860), .B(n12864), .ZN(n12861) );
  OAI222_X1 U15123 ( .A1(n12927), .A2(n12862), .B1(n12925), .B2(n9831), .C1(
        n12922), .C2(n12861), .ZN(n12976) );
  INV_X1 U15124 ( .A(n12976), .ZN(n12870) );
  XOR2_X1 U15125 ( .A(n12864), .B(n12863), .Z(n12977) );
  INV_X1 U15126 ( .A(n12865), .ZN(n13039) );
  AOI22_X1 U15127 ( .A1(n15119), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n14400), 
        .B2(n12866), .ZN(n12867) );
  OAI21_X1 U15128 ( .B1(n13039), .B2(n12933), .A(n12867), .ZN(n12868) );
  AOI21_X1 U15129 ( .B1(n12977), .B2(n12935), .A(n12868), .ZN(n12869) );
  OAI21_X1 U15130 ( .B1(n12870), .B2(n15119), .A(n12869), .ZN(P3_U3212) );
  XNOR2_X1 U15131 ( .A(n12872), .B(n12871), .ZN(n12873) );
  OAI222_X1 U15132 ( .A1(n12925), .A2(n12874), .B1(n12927), .B2(n12899), .C1(
        n12922), .C2(n12873), .ZN(n12980) );
  INV_X1 U15133 ( .A(n12980), .ZN(n12882) );
  XNOR2_X1 U15134 ( .A(n12876), .B(n12875), .ZN(n12981) );
  INV_X1 U15135 ( .A(n12877), .ZN(n13043) );
  AOI22_X1 U15136 ( .A1(n15119), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n14400), 
        .B2(n12878), .ZN(n12879) );
  OAI21_X1 U15137 ( .B1(n13043), .B2(n12933), .A(n12879), .ZN(n12880) );
  AOI21_X1 U15138 ( .B1(n12981), .B2(n12935), .A(n12880), .ZN(n12881) );
  OAI21_X1 U15139 ( .B1(n12882), .B2(n15119), .A(n12881), .ZN(P3_U3213) );
  XNOR2_X1 U15140 ( .A(n12883), .B(n12885), .ZN(n12985) );
  INV_X1 U15141 ( .A(n12985), .ZN(n12894) );
  OAI211_X1 U15142 ( .C1(n6639), .C2(n12885), .A(n12884), .B(n15106), .ZN(
        n12889) );
  AOI22_X1 U15143 ( .A1(n12887), .A2(n15104), .B1(n15103), .B2(n12886), .ZN(
        n12888) );
  NAND2_X1 U15144 ( .A1(n12889), .A2(n12888), .ZN(n12984) );
  AOI22_X1 U15145 ( .A1(n15119), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n14400), 
        .B2(n12890), .ZN(n12891) );
  OAI21_X1 U15146 ( .B1(n13047), .B2(n12933), .A(n12891), .ZN(n12892) );
  AOI21_X1 U15147 ( .B1(n12984), .B2(n15117), .A(n12892), .ZN(n12893) );
  OAI21_X1 U15148 ( .B1(n12894), .B2(n12902), .A(n12893), .ZN(P3_U3214) );
  AOI21_X1 U15149 ( .B1(n12897), .B2(n12896), .A(n12895), .ZN(n12898) );
  OAI222_X1 U15150 ( .A1(n12927), .A2(n12924), .B1(n12925), .B2(n12899), .C1(
        n12922), .C2(n12898), .ZN(n12990) );
  INV_X1 U15151 ( .A(n12991), .ZN(n12903) );
  AND2_X1 U15152 ( .A1(n12901), .A2(n12900), .ZN(n12989) );
  NOR3_X1 U15153 ( .A1(n12903), .A2(n12989), .A3(n12902), .ZN(n12907) );
  AOI22_X1 U15154 ( .A1(n15119), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n14400), 
        .B2(n12904), .ZN(n12905) );
  OAI21_X1 U15155 ( .B1(n13051), .B2(n12933), .A(n12905), .ZN(n12906) );
  AOI211_X1 U15156 ( .C1(n12990), .C2(n15117), .A(n12907), .B(n12906), .ZN(
        n12908) );
  INV_X1 U15157 ( .A(n12908), .ZN(P3_U3215) );
  XNOR2_X1 U15158 ( .A(n12909), .B(n12913), .ZN(n12910) );
  OAI222_X1 U15159 ( .A1(n12927), .A2(n12912), .B1(n12925), .B2(n12911), .C1(
        n12910), .C2(n12922), .ZN(n12995) );
  INV_X1 U15160 ( .A(n12995), .ZN(n12919) );
  XNOR2_X1 U15161 ( .A(n12914), .B(n12913), .ZN(n12996) );
  AOI22_X1 U15162 ( .A1(n15119), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n14400), 
        .B2(n12915), .ZN(n12916) );
  OAI21_X1 U15163 ( .B1(n13055), .B2(n12933), .A(n12916), .ZN(n12917) );
  AOI21_X1 U15164 ( .B1(n12996), .B2(n12935), .A(n12917), .ZN(n12918) );
  OAI21_X1 U15165 ( .B1(n12919), .B2(n15119), .A(n12918), .ZN(P3_U3216) );
  XNOR2_X1 U15166 ( .A(n12920), .B(n12921), .ZN(n12923) );
  OAI222_X1 U15167 ( .A1(n12927), .A2(n12926), .B1(n12925), .B2(n12924), .C1(
        n12923), .C2(n12922), .ZN(n12999) );
  INV_X1 U15168 ( .A(n12999), .ZN(n12937) );
  OAI21_X1 U15169 ( .B1(n12929), .B2(n6765), .A(n12928), .ZN(n13000) );
  INV_X1 U15170 ( .A(n12930), .ZN(n13060) );
  AOI22_X1 U15171 ( .A1(n15119), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n14400), 
        .B2(n12931), .ZN(n12932) );
  OAI21_X1 U15172 ( .B1(n13060), .B2(n12933), .A(n12932), .ZN(n12934) );
  AOI21_X1 U15173 ( .B1(n13000), .B2(n12935), .A(n12934), .ZN(n12936) );
  OAI21_X1 U15174 ( .B1(n12937), .B2(n15119), .A(n12936), .ZN(P3_U3217) );
  INV_X1 U15175 ( .A(n13003), .ZN(n12941) );
  NAND2_X1 U15176 ( .A1(n12938), .A2(n12941), .ZN(n12940) );
  INV_X1 U15177 ( .A(n13008), .ZN(n12939) );
  NAND2_X1 U15178 ( .A1(n15183), .A2(n12939), .ZN(n12943) );
  OAI211_X1 U15179 ( .C1(n15183), .C2(n12146), .A(n12940), .B(n12943), .ZN(
        P3_U3490) );
  NAND2_X1 U15180 ( .A1(n12942), .A2(n12941), .ZN(n12944) );
  OAI211_X1 U15181 ( .C1(n15183), .C2(n8864), .A(n12944), .B(n12943), .ZN(
        P3_U3489) );
  INV_X1 U15182 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n12947) );
  AOI21_X1 U15183 ( .B1(n12946), .B2(n14415), .A(n12945), .ZN(n13014) );
  MUX2_X1 U15184 ( .A(n12947), .B(n13014), .S(n15183), .Z(n12948) );
  OAI21_X1 U15185 ( .B1(n13017), .B2(n13003), .A(n12948), .ZN(P3_U3487) );
  NAND2_X1 U15186 ( .A1(n12949), .A2(n15150), .ZN(n12950) );
  OAI211_X1 U15187 ( .C1(n12952), .C2(n15169), .A(n12951), .B(n12950), .ZN(
        n13018) );
  MUX2_X1 U15188 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n13018), .S(n15183), .Z(
        P3_U3486) );
  INV_X1 U15189 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12955) );
  AOI21_X1 U15190 ( .B1(n12954), .B2(n14415), .A(n12953), .ZN(n13019) );
  MUX2_X1 U15191 ( .A(n12955), .B(n13019), .S(n15183), .Z(n12956) );
  OAI21_X1 U15192 ( .B1(n13022), .B2(n13003), .A(n12956), .ZN(P3_U3485) );
  AOI21_X1 U15193 ( .B1(n15164), .B2(n12958), .A(n12957), .ZN(n13023) );
  MUX2_X1 U15194 ( .A(n12959), .B(n13023), .S(n15183), .Z(n12960) );
  OAI21_X1 U15195 ( .B1(n13026), .B2(n13003), .A(n12960), .ZN(P3_U3484) );
  INV_X1 U15196 ( .A(n12961), .ZN(n12963) );
  AOI21_X1 U15197 ( .B1(n15164), .B2(n12963), .A(n12962), .ZN(n13027) );
  MUX2_X1 U15198 ( .A(n12964), .B(n13027), .S(n15183), .Z(n12965) );
  OAI21_X1 U15199 ( .B1(n13030), .B2(n13003), .A(n12965), .ZN(P3_U3483) );
  INV_X1 U15200 ( .A(n12966), .ZN(n13034) );
  INV_X1 U15201 ( .A(n12967), .ZN(n12969) );
  AOI21_X1 U15202 ( .B1(n15164), .B2(n12969), .A(n12968), .ZN(n13031) );
  MUX2_X1 U15203 ( .A(n12970), .B(n13031), .S(n15183), .Z(n12971) );
  OAI21_X1 U15204 ( .B1(n13034), .B2(n13003), .A(n12971), .ZN(P3_U3482) );
  NAND2_X1 U15205 ( .A1(n12972), .A2(n14415), .ZN(n12973) );
  OAI211_X1 U15206 ( .C1(n12975), .C2(n15168), .A(n12974), .B(n12973), .ZN(
        n13035) );
  MUX2_X1 U15207 ( .A(P3_REG1_REG_22__SCAN_IN), .B(n13035), .S(n15183), .Z(
        P3_U3481) );
  AOI21_X1 U15208 ( .B1(n12977), .B2(n14415), .A(n12976), .ZN(n13036) );
  MUX2_X1 U15209 ( .A(n12978), .B(n13036), .S(n15183), .Z(n12979) );
  OAI21_X1 U15210 ( .B1(n13039), .B2(n13003), .A(n12979), .ZN(P3_U3480) );
  AOI21_X1 U15211 ( .B1(n14415), .B2(n12981), .A(n12980), .ZN(n13040) );
  MUX2_X1 U15212 ( .A(n12982), .B(n13040), .S(n15183), .Z(n12983) );
  OAI21_X1 U15213 ( .B1(n13043), .B2(n13003), .A(n12983), .ZN(P3_U3479) );
  INV_X1 U15214 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12986) );
  AOI21_X1 U15215 ( .B1(n14415), .B2(n12985), .A(n12984), .ZN(n13044) );
  MUX2_X1 U15216 ( .A(n12986), .B(n13044), .S(n15183), .Z(n12987) );
  OAI21_X1 U15217 ( .B1(n13003), .B2(n13047), .A(n12987), .ZN(P3_U3478) );
  NOR2_X1 U15218 ( .A1(n12989), .A2(n12988), .ZN(n12992) );
  AOI21_X1 U15219 ( .B1(n12992), .B2(n12991), .A(n12990), .ZN(n13048) );
  MUX2_X1 U15220 ( .A(n12993), .B(n13048), .S(n15183), .Z(n12994) );
  OAI21_X1 U15221 ( .B1(n13051), .B2(n13003), .A(n12994), .ZN(P3_U3477) );
  AOI21_X1 U15222 ( .B1(n12996), .B2(n14415), .A(n12995), .ZN(n13052) );
  MUX2_X1 U15223 ( .A(n12997), .B(n13052), .S(n15183), .Z(n12998) );
  OAI21_X1 U15224 ( .B1(n13055), .B2(n13003), .A(n12998), .ZN(P3_U3476) );
  AOI21_X1 U15225 ( .B1(n14415), .B2(n13000), .A(n12999), .ZN(n13056) );
  MUX2_X1 U15226 ( .A(n13001), .B(n13056), .S(n15183), .Z(n13002) );
  OAI21_X1 U15227 ( .B1(n13060), .B2(n13003), .A(n13002), .ZN(P3_U3475) );
  NAND2_X1 U15228 ( .A1(n13004), .A2(n14415), .ZN(n13005) );
  OAI211_X1 U15229 ( .C1(n13007), .C2(n15168), .A(n13006), .B(n13005), .ZN(
        n13061) );
  MUX2_X1 U15230 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n13061), .S(n15183), .Z(
        P3_U3474) );
  NOR2_X1 U15231 ( .A1(n15173), .A2(n13008), .ZN(n13011) );
  AOI21_X1 U15232 ( .B1(n15173), .B2(P3_REG0_REG_31__SCAN_IN), .A(n13011), 
        .ZN(n13009) );
  OAI21_X1 U15233 ( .B1(n13010), .B2(n13059), .A(n13009), .ZN(P3_U3458) );
  AOI21_X1 U15234 ( .B1(n15173), .B2(P3_REG0_REG_30__SCAN_IN), .A(n13011), 
        .ZN(n13012) );
  OAI21_X1 U15235 ( .B1(n13013), .B2(n13059), .A(n13012), .ZN(P3_U3457) );
  MUX2_X1 U15236 ( .A(n13015), .B(n13014), .S(n15175), .Z(n13016) );
  OAI21_X1 U15237 ( .B1(n13017), .B2(n13059), .A(n13016), .ZN(P3_U3455) );
  MUX2_X1 U15238 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n13018), .S(n15175), .Z(
        P3_U3454) );
  MUX2_X1 U15239 ( .A(n13020), .B(n13019), .S(n15175), .Z(n13021) );
  OAI21_X1 U15240 ( .B1(n13022), .B2(n13059), .A(n13021), .ZN(P3_U3453) );
  INV_X1 U15241 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13024) );
  MUX2_X1 U15242 ( .A(n13024), .B(n13023), .S(n15175), .Z(n13025) );
  OAI21_X1 U15243 ( .B1(n13026), .B2(n13059), .A(n13025), .ZN(P3_U3452) );
  INV_X1 U15244 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13028) );
  MUX2_X1 U15245 ( .A(n13028), .B(n13027), .S(n15175), .Z(n13029) );
  OAI21_X1 U15246 ( .B1(n13030), .B2(n13059), .A(n13029), .ZN(P3_U3451) );
  INV_X1 U15247 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13032) );
  MUX2_X1 U15248 ( .A(n13032), .B(n13031), .S(n15175), .Z(n13033) );
  OAI21_X1 U15249 ( .B1(n13034), .B2(n13059), .A(n13033), .ZN(P3_U3450) );
  MUX2_X1 U15250 ( .A(P3_REG0_REG_22__SCAN_IN), .B(n13035), .S(n15175), .Z(
        P3_U3449) );
  INV_X1 U15251 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13037) );
  MUX2_X1 U15252 ( .A(n13037), .B(n13036), .S(n15175), .Z(n13038) );
  OAI21_X1 U15253 ( .B1(n13039), .B2(n13059), .A(n13038), .ZN(P3_U3448) );
  INV_X1 U15254 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13041) );
  MUX2_X1 U15255 ( .A(n13041), .B(n13040), .S(n15175), .Z(n13042) );
  OAI21_X1 U15256 ( .B1(n13043), .B2(n13059), .A(n13042), .ZN(P3_U3447) );
  INV_X1 U15257 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13045) );
  MUX2_X1 U15258 ( .A(n13045), .B(n13044), .S(n15175), .Z(n13046) );
  OAI21_X1 U15259 ( .B1(n13059), .B2(n13047), .A(n13046), .ZN(P3_U3446) );
  INV_X1 U15260 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13049) );
  MUX2_X1 U15261 ( .A(n13049), .B(n13048), .S(n15175), .Z(n13050) );
  OAI21_X1 U15262 ( .B1(n13051), .B2(n13059), .A(n13050), .ZN(P3_U3444) );
  INV_X1 U15263 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13053) );
  MUX2_X1 U15264 ( .A(n13053), .B(n13052), .S(n15175), .Z(n13054) );
  OAI21_X1 U15265 ( .B1(n13055), .B2(n13059), .A(n13054), .ZN(P3_U3441) );
  MUX2_X1 U15266 ( .A(n13057), .B(n13056), .S(n15175), .Z(n13058) );
  OAI21_X1 U15267 ( .B1(n13060), .B2(n13059), .A(n13058), .ZN(P3_U3438) );
  MUX2_X1 U15268 ( .A(P3_REG0_REG_15__SCAN_IN), .B(n13061), .S(n15175), .Z(
        P3_U3435) );
  MUX2_X1 U15269 ( .A(P3_D_REG_1__SCAN_IN), .B(n13062), .S(n13063), .Z(
        P3_U3377) );
  MUX2_X1 U15270 ( .A(P3_D_REG_0__SCAN_IN), .B(n13064), .S(n13063), .Z(
        P3_U3376) );
  NAND3_X1 U15271 ( .A1(n13065), .A2(P3_STATE_REG_SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .ZN(n13067) );
  OAI22_X1 U15272 ( .A1(n13068), .A2(n13067), .B1(n13066), .B2(n13078), .ZN(
        n13069) );
  AOI21_X1 U15273 ( .B1(n13071), .B2(n13070), .A(n13069), .ZN(n13072) );
  INV_X1 U15274 ( .A(n13072), .ZN(P3_U3264) );
  INV_X1 U15275 ( .A(n13073), .ZN(n13075) );
  OAI222_X1 U15276 ( .A1(n13078), .A2(n15285), .B1(n13076), .B2(n13075), .C1(
        P3_U3151), .C2(n8355), .ZN(P3_U3266) );
  INV_X1 U15277 ( .A(n13077), .ZN(n13080) );
  OAI222_X1 U15278 ( .A1(n13076), .A2(n13080), .B1(n13079), .B2(P3_U3151), 
        .C1(n15236), .C2(n13078), .ZN(P3_U3267) );
  INV_X1 U15279 ( .A(n13547), .ZN(n13352) );
  AND2_X1 U15280 ( .A1(n13082), .A2(n13081), .ZN(n13083) );
  NOR2_X2 U15281 ( .A1(n13084), .A2(n13083), .ZN(n13086) );
  XNOR2_X1 U15282 ( .A(n13569), .B(n6725), .ZN(n13087) );
  XNOR2_X1 U15283 ( .A(n13086), .B(n13087), .ZN(n13115) );
  AND2_X1 U15284 ( .A1(n13247), .A2(n13489), .ZN(n13085) );
  NAND2_X1 U15285 ( .A1(n13115), .A2(n13085), .ZN(n13114) );
  INV_X1 U15286 ( .A(n13086), .ZN(n13088) );
  NAND2_X1 U15287 ( .A1(n13114), .A2(n13089), .ZN(n13192) );
  XNOR2_X1 U15288 ( .A(n13401), .B(n13134), .ZN(n13162) );
  NAND2_X1 U15289 ( .A1(n13246), .A2(n13105), .ZN(n13090) );
  NOR2_X1 U15290 ( .A1(n13162), .A2(n13090), .ZN(n13091) );
  AOI21_X1 U15291 ( .B1(n13162), .B2(n13090), .A(n13091), .ZN(n13193) );
  NAND2_X1 U15292 ( .A1(n13192), .A2(n13193), .ZN(n13158) );
  INV_X1 U15293 ( .A(n13091), .ZN(n13092) );
  XNOR2_X1 U15294 ( .A(n13558), .B(n6725), .ZN(n13226) );
  AND2_X1 U15295 ( .A1(n13245), .A2(n13489), .ZN(n13093) );
  NAND2_X1 U15296 ( .A1(n13226), .A2(n13093), .ZN(n13099) );
  INV_X1 U15297 ( .A(n13226), .ZN(n13095) );
  INV_X1 U15298 ( .A(n13093), .ZN(n13094) );
  NAND2_X1 U15299 ( .A1(n13095), .A2(n13094), .ZN(n13096) );
  XNOR2_X1 U15300 ( .A(n13553), .B(n6725), .ZN(n13101) );
  NAND2_X1 U15301 ( .A1(n13244), .A2(n13105), .ZN(n13102) );
  XNOR2_X1 U15302 ( .A(n13101), .B(n13102), .ZN(n13228) );
  INV_X1 U15303 ( .A(n13101), .ZN(n13103) );
  NAND2_X1 U15304 ( .A1(n13103), .A2(n13102), .ZN(n13104) );
  XNOR2_X1 U15305 ( .A(n13547), .B(n13134), .ZN(n13131) );
  NAND2_X1 U15306 ( .A1(n13243), .A2(n13105), .ZN(n13106) );
  NOR2_X1 U15307 ( .A1(n13131), .A2(n13106), .ZN(n13143) );
  AOI21_X1 U15308 ( .B1(n13131), .B2(n13106), .A(n13143), .ZN(n13107) );
  OAI22_X1 U15309 ( .A1(n13133), .A2(n14422), .B1(n13167), .B2(n14420), .ZN(
        n13356) );
  INV_X1 U15310 ( .A(n13350), .ZN(n13110) );
  OAI22_X1 U15311 ( .A1(n13110), .A2(n14789), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13109), .ZN(n13111) );
  AOI21_X1 U15312 ( .B1(n13356), .B2(n14430), .A(n13111), .ZN(n13112) );
  INV_X1 U15313 ( .A(n13114), .ZN(n13121) );
  AOI22_X1 U15314 ( .A1(n13115), .A2(n14428), .B1(n13225), .B2(n13247), .ZN(
        n13120) );
  AOI22_X1 U15315 ( .A1(n13246), .A2(n13233), .B1(n13231), .B2(n13248), .ZN(
        n13409) );
  OAI22_X1 U15316 ( .A1(n13409), .A2(n14779), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13116), .ZN(n13117) );
  AOI21_X1 U15317 ( .B1(n13418), .B2(n13208), .A(n13117), .ZN(n13119) );
  NAND2_X1 U15318 ( .A1(n13569), .A2(n14787), .ZN(n13118) );
  OAI211_X1 U15319 ( .C1(n13121), .C2(n13120), .A(n13119), .B(n13118), .ZN(
        P2_U3188) );
  OAI21_X1 U15320 ( .B1(n13124), .B2(n13123), .A(n13122), .ZN(n13125) );
  XNOR2_X1 U15321 ( .A(n13202), .B(n13125), .ZN(n13130) );
  NOR2_X1 U15322 ( .A1(n14789), .A2(n13473), .ZN(n13128) );
  AND2_X1 U15323 ( .A1(n13252), .A2(n13231), .ZN(n13126) );
  AOI21_X1 U15324 ( .B1(n13250), .B2(n13233), .A(n13126), .ZN(n13467) );
  NAND2_X1 U15325 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13317)
         );
  OAI21_X1 U15326 ( .B1(n13467), .B2(n14779), .A(n13317), .ZN(n13127) );
  AOI211_X1 U15327 ( .C1(n13591), .C2(n14787), .A(n13128), .B(n13127), .ZN(
        n13129) );
  OAI21_X1 U15328 ( .B1(n13130), .B2(n14782), .A(n13129), .ZN(P2_U3191) );
  INV_X1 U15329 ( .A(n13131), .ZN(n13132) );
  NOR2_X1 U15330 ( .A1(n13133), .A2(n13523), .ZN(n13135) );
  XNOR2_X1 U15331 ( .A(n13135), .B(n13134), .ZN(n13136) );
  XNOR2_X1 U15332 ( .A(n13344), .B(n13136), .ZN(n13144) );
  NAND2_X1 U15333 ( .A1(n13137), .A2(n13144), .ZN(n13150) );
  NAND2_X1 U15334 ( .A1(n13241), .A2(n13233), .ZN(n13139) );
  NAND2_X1 U15335 ( .A1(n13243), .A2(n13231), .ZN(n13138) );
  NAND2_X1 U15336 ( .A1(n13139), .A2(n13138), .ZN(n13334) );
  OAI22_X1 U15337 ( .A1(n13338), .A2(n14789), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13140), .ZN(n13142) );
  NOR2_X1 U15338 ( .A1(n13344), .A2(n13210), .ZN(n13141) );
  AOI211_X1 U15339 ( .C1(n14430), .C2(n13334), .A(n13142), .B(n13141), .ZN(
        n13149) );
  INV_X1 U15340 ( .A(n13143), .ZN(n13146) );
  INV_X1 U15341 ( .A(n13144), .ZN(n13145) );
  NAND4_X1 U15342 ( .A1(n13147), .A2(n14428), .A3(n13146), .A4(n13145), .ZN(
        n13148) );
  NAND3_X1 U15343 ( .A1(n13150), .A2(n13149), .A3(n13148), .ZN(P2_U3192) );
  OAI211_X1 U15344 ( .C1(n13153), .C2(n13152), .A(n13151), .B(n14428), .ZN(
        n13157) );
  AOI22_X1 U15345 ( .A1(n13248), .A2(n13233), .B1(n13231), .B2(n13250), .ZN(
        n13443) );
  OAI22_X1 U15346 ( .A1(n13443), .A2(n14779), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13154), .ZN(n13155) );
  AOI21_X1 U15347 ( .B1(n13447), .B2(n13208), .A(n13155), .ZN(n13156) );
  OAI211_X1 U15348 ( .C1(n13450), .C2(n13210), .A(n13157), .B(n13156), .ZN(
        P2_U3195) );
  BUF_X1 U15349 ( .A(n13158), .Z(n13159) );
  INV_X1 U15350 ( .A(n13160), .ZN(n13161) );
  AOI21_X1 U15351 ( .B1(n13159), .B2(n13161), .A(n14782), .ZN(n13165) );
  INV_X1 U15352 ( .A(n13246), .ZN(n13166) );
  NOR3_X1 U15353 ( .A1(n13162), .A2(n13166), .A3(n13201), .ZN(n13164) );
  OAI21_X1 U15354 ( .B1(n13165), .B2(n13164), .A(n13163), .ZN(n13172) );
  OAI22_X1 U15355 ( .A1(n13167), .A2(n14422), .B1(n13166), .B2(n14420), .ZN(
        n13377) );
  INV_X1 U15356 ( .A(n13385), .ZN(n13169) );
  OAI22_X1 U15357 ( .A1(n13169), .A2(n14789), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13168), .ZN(n13170) );
  AOI21_X1 U15358 ( .B1(n13377), .B2(n14430), .A(n13170), .ZN(n13171) );
  OAI211_X1 U15359 ( .C1(n7474), .C2(n13210), .A(n13172), .B(n13171), .ZN(
        P2_U3197) );
  AOI21_X1 U15360 ( .B1(n13175), .B2(n13174), .A(n13173), .ZN(n13181) );
  INV_X1 U15361 ( .A(n13176), .ZN(n13519) );
  OAI22_X1 U15362 ( .A1(n13218), .A2(n14422), .B1(n14423), .B2(n14420), .ZN(
        n13513) );
  NAND2_X1 U15363 ( .A1(n14430), .A2(n13513), .ZN(n13177) );
  OAI211_X1 U15364 ( .C1(n14789), .C2(n13519), .A(n13178), .B(n13177), .ZN(
        n13179) );
  AOI21_X1 U15365 ( .B1(n13607), .B2(n14787), .A(n13179), .ZN(n13180) );
  OAI21_X1 U15366 ( .B1(n13181), .B2(n14782), .A(n13180), .ZN(P2_U3198) );
  AOI21_X1 U15367 ( .B1(n13184), .B2(n13183), .A(n7308), .ZN(n13191) );
  OAI22_X1 U15368 ( .A1(n13186), .A2(n14422), .B1(n13185), .B2(n14420), .ZN(
        n13497) );
  NAND2_X1 U15369 ( .A1(n13497), .A2(n14430), .ZN(n13188) );
  OAI211_X1 U15370 ( .C1(n14789), .C2(n13502), .A(n13188), .B(n13187), .ZN(
        n13189) );
  AOI21_X1 U15371 ( .B1(n13600), .B2(n14787), .A(n13189), .ZN(n13190) );
  OAI21_X1 U15372 ( .B1(n13191), .B2(n14782), .A(n13190), .ZN(P2_U3200) );
  OAI211_X1 U15373 ( .C1(n13194), .C2(n13193), .A(n13159), .B(n14428), .ZN(
        n13200) );
  OAI22_X1 U15374 ( .A1(n13196), .A2(n14422), .B1(n13195), .B2(n14420), .ZN(
        n13392) );
  OAI22_X1 U15375 ( .A1(n13399), .A2(n14789), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13197), .ZN(n13198) );
  AOI21_X1 U15376 ( .B1(n13392), .B2(n14430), .A(n13198), .ZN(n13199) );
  OAI211_X1 U15377 ( .C1(n13563), .C2(n13210), .A(n13200), .B(n13199), .ZN(
        P2_U3201) );
  NOR3_X1 U15378 ( .A1(n13202), .A2(n13219), .A3(n13201), .ZN(n13203) );
  AOI21_X1 U15379 ( .B1(n14428), .B2(n13204), .A(n13203), .ZN(n13215) );
  INV_X1 U15380 ( .A(n13205), .ZN(n13214) );
  INV_X1 U15381 ( .A(n13586), .ZN(n13462) );
  AOI22_X1 U15382 ( .A1(n13249), .A2(n13233), .B1(n13231), .B2(n13251), .ZN(
        n13456) );
  OAI22_X1 U15383 ( .A1(n13456), .A2(n14779), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13206), .ZN(n13207) );
  AOI21_X1 U15384 ( .B1(n13459), .B2(n13208), .A(n13207), .ZN(n13209) );
  OAI21_X1 U15385 ( .B1(n13462), .B2(n13210), .A(n13209), .ZN(n13211) );
  AOI21_X1 U15386 ( .B1(n13212), .B2(n14428), .A(n13211), .ZN(n13213) );
  OAI21_X1 U15387 ( .B1(n13215), .B2(n13214), .A(n13213), .ZN(P2_U3205) );
  XNOR2_X1 U15388 ( .A(n13217), .B(n13216), .ZN(n13224) );
  OAI22_X1 U15389 ( .A1(n13219), .A2(n14422), .B1(n13218), .B2(n14420), .ZN(
        n13481) );
  NAND2_X1 U15390 ( .A1(n13481), .A2(n14430), .ZN(n13221) );
  OAI211_X1 U15391 ( .C1(n14789), .C2(n13486), .A(n13221), .B(n13220), .ZN(
        n13222) );
  AOI21_X1 U15392 ( .B1(n13595), .B2(n14787), .A(n13222), .ZN(n13223) );
  OAI21_X1 U15393 ( .B1(n13224), .B2(n14782), .A(n13223), .ZN(P2_U3210) );
  NAND3_X1 U15394 ( .A1(n13226), .A2(n13225), .A3(n13245), .ZN(n13227) );
  OAI21_X1 U15395 ( .B1(n13163), .B2(n14782), .A(n13227), .ZN(n13230) );
  INV_X1 U15396 ( .A(n13228), .ZN(n13229) );
  NAND2_X1 U15397 ( .A1(n13230), .A2(n13229), .ZN(n13238) );
  AND2_X1 U15398 ( .A1(n13245), .A2(n13231), .ZN(n13232) );
  AOI21_X1 U15399 ( .B1(n13243), .B2(n13233), .A(n13232), .ZN(n13364) );
  NOR2_X1 U15400 ( .A1(n13364), .A2(n14779), .ZN(n13236) );
  OAI22_X1 U15401 ( .A1(n13368), .A2(n14789), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13234), .ZN(n13235) );
  AOI211_X1 U15402 ( .C1(n13553), .C2(n14787), .A(n13236), .B(n13235), .ZN(
        n13237) );
  OAI211_X1 U15403 ( .C1(n13239), .C2(n14782), .A(n13238), .B(n13237), .ZN(
        P2_U3212) );
  INV_X2 U15404 ( .A(P2_U3947), .ZN(n13269) );
  MUX2_X1 U15405 ( .A(n13322), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13269), .Z(
        P2_U3562) );
  MUX2_X1 U15406 ( .A(n13240), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13269), .Z(
        P2_U3561) );
  MUX2_X1 U15407 ( .A(n13241), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13269), .Z(
        P2_U3560) );
  MUX2_X1 U15408 ( .A(n13242), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13269), .Z(
        P2_U3559) );
  MUX2_X1 U15409 ( .A(n13243), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13269), .Z(
        P2_U3558) );
  MUX2_X1 U15410 ( .A(n13244), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13269), .Z(
        P2_U3557) );
  MUX2_X1 U15411 ( .A(n13245), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13269), .Z(
        P2_U3556) );
  MUX2_X1 U15412 ( .A(n13246), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13269), .Z(
        P2_U3555) );
  MUX2_X1 U15413 ( .A(n13247), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13269), .Z(
        P2_U3554) );
  MUX2_X1 U15414 ( .A(n13248), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13269), .Z(
        P2_U3553) );
  MUX2_X1 U15415 ( .A(n13249), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13269), .Z(
        P2_U3552) );
  MUX2_X1 U15416 ( .A(n13250), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13269), .Z(
        P2_U3551) );
  MUX2_X1 U15417 ( .A(n13251), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13269), .Z(
        P2_U3550) );
  MUX2_X1 U15418 ( .A(n13252), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13269), .Z(
        P2_U3549) );
  MUX2_X1 U15419 ( .A(n13253), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13269), .Z(
        P2_U3548) );
  MUX2_X1 U15420 ( .A(n13254), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13269), .Z(
        P2_U3547) );
  MUX2_X1 U15421 ( .A(n13255), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13269), .Z(
        P2_U3546) );
  MUX2_X1 U15422 ( .A(n13256), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13269), .Z(
        P2_U3545) );
  MUX2_X1 U15423 ( .A(n13257), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13269), .Z(
        P2_U3544) );
  MUX2_X1 U15424 ( .A(n13258), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13269), .Z(
        P2_U3543) );
  MUX2_X1 U15425 ( .A(n13259), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13269), .Z(
        P2_U3542) );
  MUX2_X1 U15426 ( .A(n13260), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13269), .Z(
        P2_U3541) );
  MUX2_X1 U15427 ( .A(n13261), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13269), .Z(
        P2_U3540) );
  MUX2_X1 U15428 ( .A(n13262), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13269), .Z(
        P2_U3539) );
  MUX2_X1 U15429 ( .A(n13263), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13269), .Z(
        P2_U3538) );
  MUX2_X1 U15430 ( .A(n13264), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13269), .Z(
        P2_U3537) );
  MUX2_X1 U15431 ( .A(n13265), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13269), .Z(
        P2_U3536) );
  MUX2_X1 U15432 ( .A(n13266), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13269), .Z(
        P2_U3535) );
  MUX2_X1 U15433 ( .A(n13267), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13269), .Z(
        P2_U3534) );
  MUX2_X1 U15434 ( .A(n13268), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13269), .Z(
        P2_U3533) );
  MUX2_X1 U15435 ( .A(n13270), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13269), .Z(
        P2_U3532) );
  INV_X1 U15436 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n13272) );
  OAI21_X1 U15437 ( .B1(n14832), .B2(n13272), .A(n13271), .ZN(n13273) );
  AOI21_X1 U15438 ( .B1(n13278), .B2(n14873), .A(n13273), .ZN(n13285) );
  MUX2_X1 U15439 ( .A(n10297), .B(P2_REG2_REG_6__SCAN_IN), .S(n13278), .Z(
        n13274) );
  NAND3_X1 U15440 ( .A1(n13276), .A2(n13275), .A3(n13274), .ZN(n13277) );
  NAND3_X1 U15441 ( .A1(n14875), .A2(n13290), .A3(n13277), .ZN(n13284) );
  MUX2_X1 U15442 ( .A(n10277), .B(P2_REG1_REG_6__SCAN_IN), .S(n13278), .Z(
        n13279) );
  NAND3_X1 U15443 ( .A1(n13281), .A2(n13280), .A3(n13279), .ZN(n13282) );
  NAND3_X1 U15444 ( .A1(n14878), .A2(n13296), .A3(n13282), .ZN(n13283) );
  NAND3_X1 U15445 ( .A1(n13285), .A2(n13284), .A3(n13283), .ZN(P2_U3220) );
  INV_X1 U15446 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n14289) );
  OAI21_X1 U15447 ( .B1(n14832), .B2(n14289), .A(n13286), .ZN(n13287) );
  AOI21_X1 U15448 ( .B1(n13293), .B2(n14873), .A(n13287), .ZN(n13301) );
  MUX2_X1 U15449 ( .A(n11227), .B(P2_REG2_REG_7__SCAN_IN), .S(n13293), .Z(
        n13288) );
  NAND3_X1 U15450 ( .A1(n13290), .A2(n13289), .A3(n13288), .ZN(n13291) );
  NAND3_X1 U15451 ( .A1(n14875), .A2(n13292), .A3(n13291), .ZN(n13300) );
  MUX2_X1 U15452 ( .A(n10280), .B(P2_REG1_REG_7__SCAN_IN), .S(n13293), .Z(
        n13294) );
  NAND3_X1 U15453 ( .A1(n13296), .A2(n13295), .A3(n13294), .ZN(n13297) );
  NAND3_X1 U15454 ( .A1(n14878), .A2(n13298), .A3(n13297), .ZN(n13299) );
  NAND3_X1 U15455 ( .A1(n13301), .A2(n13300), .A3(n13299), .ZN(P2_U3221) );
  NOR2_X1 U15456 ( .A1(n13303), .A2(n13302), .ZN(n13304) );
  XOR2_X1 U15457 ( .A(n13304), .B(P2_REG2_REG_19__SCAN_IN), .Z(n13314) );
  INV_X1 U15458 ( .A(n13314), .ZN(n13312) );
  NAND2_X1 U15459 ( .A1(n13306), .A2(n13305), .ZN(n13307) );
  NAND2_X1 U15460 ( .A1(n13308), .A2(n13307), .ZN(n13310) );
  INV_X1 U15461 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13309) );
  XNOR2_X1 U15462 ( .A(n13310), .B(n13309), .ZN(n13313) );
  NOR2_X1 U15463 ( .A1(n13313), .A2(n14862), .ZN(n13311) );
  AOI211_X1 U15464 ( .C1(n13312), .C2(n14875), .A(n14873), .B(n13311), .ZN(
        n13316) );
  AOI22_X1 U15465 ( .A1(n13314), .A2(n14875), .B1(n14878), .B2(n13313), .ZN(
        n13315) );
  MUX2_X1 U15466 ( .A(n13316), .B(n13315), .S(n9432), .Z(n13318) );
  OAI211_X1 U15467 ( .C1(n7528), .C2(n14832), .A(n13318), .B(n13317), .ZN(
        P2_U3233) );
  NAND2_X1 U15468 ( .A1(n13535), .A2(n13326), .ZN(n13325) );
  NAND2_X1 U15469 ( .A1(n13322), .A2(n13321), .ZN(n13533) );
  NOR2_X1 U15470 ( .A1(n13531), .A2(n13533), .ZN(n13328) );
  NOR2_X1 U15471 ( .A1(n13319), .A2(n13472), .ZN(n13323) );
  AOI211_X1 U15472 ( .C1(n13531), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13328), 
        .B(n13323), .ZN(n13324) );
  OAI21_X1 U15473 ( .B1(n13532), .B2(n14898), .A(n13324), .ZN(P2_U3234) );
  OAI211_X1 U15474 ( .C1(n13535), .C2(n13326), .A(n13523), .B(n13325), .ZN(
        n13534) );
  NOR2_X1 U15475 ( .A1(n13535), .A2(n13472), .ZN(n13327) );
  AOI211_X1 U15476 ( .C1(n13531), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13328), 
        .B(n13327), .ZN(n13329) );
  OAI21_X1 U15477 ( .B1(n14898), .B2(n13534), .A(n13329), .ZN(P2_U3235) );
  XNOR2_X1 U15478 ( .A(n13330), .B(n13332), .ZN(n13545) );
  NAND2_X1 U15479 ( .A1(n13331), .A2(n14886), .ZN(n13337) );
  AOI21_X1 U15480 ( .B1(n13353), .B2(n13333), .A(n13332), .ZN(n13336) );
  INV_X1 U15481 ( .A(n13334), .ZN(n13335) );
  NOR2_X1 U15482 ( .A1(n13338), .A2(n13518), .ZN(n13339) );
  OAI21_X1 U15483 ( .B1(n13541), .B2(n13339), .A(n14919), .ZN(n13347) );
  INV_X1 U15484 ( .A(n13349), .ZN(n13342) );
  INV_X1 U15485 ( .A(n13340), .ZN(n13341) );
  AOI211_X1 U15486 ( .C1(n13543), .C2(n13342), .A(n13489), .B(n13341), .ZN(
        n13542) );
  INV_X1 U15487 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13343) );
  OAI22_X1 U15488 ( .A1(n13344), .A2(n13472), .B1(n13343), .B2(n14919), .ZN(
        n13345) );
  AOI21_X1 U15489 ( .B1(n13542), .B2(n14916), .A(n13345), .ZN(n13346) );
  OAI211_X1 U15490 ( .C1(n13528), .C2(n13545), .A(n13347), .B(n13346), .ZN(
        P2_U3237) );
  XNOR2_X1 U15491 ( .A(n13348), .B(n7119), .ZN(n13550) );
  AOI211_X1 U15492 ( .C1(n13547), .C2(n13365), .A(n13105), .B(n13349), .ZN(
        n13546) );
  AOI22_X1 U15493 ( .A1(n13350), .A2(n14905), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n14903), .ZN(n13351) );
  OAI21_X1 U15494 ( .B1(n13352), .B2(n13472), .A(n13351), .ZN(n13359) );
  OAI21_X1 U15495 ( .B1(n13355), .B2(n13354), .A(n13353), .ZN(n13357) );
  AOI21_X1 U15496 ( .B1(n13357), .B2(n14886), .A(n13356), .ZN(n13549) );
  NOR2_X1 U15497 ( .A1(n13549), .A2(n14903), .ZN(n13358) );
  AOI211_X1 U15498 ( .C1(n13546), .C2(n14916), .A(n13359), .B(n13358), .ZN(
        n13360) );
  OAI21_X1 U15499 ( .B1(n13550), .B2(n13528), .A(n13360), .ZN(P2_U3238) );
  XOR2_X1 U15500 ( .A(n13363), .B(n13361), .Z(n13555) );
  NAND2_X1 U15501 ( .A1(n13551), .A2(n14919), .ZN(n13374) );
  INV_X1 U15502 ( .A(n13384), .ZN(n13367) );
  INV_X1 U15503 ( .A(n13365), .ZN(n13366) );
  AOI211_X1 U15504 ( .C1(n13553), .C2(n13367), .A(n13489), .B(n13366), .ZN(
        n13552) );
  INV_X1 U15505 ( .A(n13368), .ZN(n13369) );
  AOI22_X1 U15506 ( .A1(n13369), .A2(n14905), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n14903), .ZN(n13370) );
  OAI21_X1 U15507 ( .B1(n13371), .B2(n13472), .A(n13370), .ZN(n13372) );
  AOI21_X1 U15508 ( .B1(n13552), .B2(n14916), .A(n13372), .ZN(n13373) );
  OAI211_X1 U15509 ( .C1(n13555), .C2(n13528), .A(n13374), .B(n13373), .ZN(
        P2_U3239) );
  XNOR2_X1 U15510 ( .A(n13376), .B(n13375), .ZN(n13378) );
  AOI21_X1 U15511 ( .B1(n13378), .B2(n14886), .A(n13377), .ZN(n13560) );
  OAI21_X1 U15512 ( .B1(n13381), .B2(n13380), .A(n13379), .ZN(n13556) );
  NAND2_X1 U15513 ( .A1(n13558), .A2(n13397), .ZN(n13382) );
  NAND2_X1 U15514 ( .A1(n13382), .A2(n13523), .ZN(n13383) );
  NOR2_X1 U15515 ( .A1(n13384), .A2(n13383), .ZN(n13557) );
  NAND2_X1 U15516 ( .A1(n13557), .A2(n14916), .ZN(n13387) );
  AOI22_X1 U15517 ( .A1(n13385), .A2(n14905), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n14903), .ZN(n13386) );
  OAI211_X1 U15518 ( .C1(n7474), .C2(n13472), .A(n13387), .B(n13386), .ZN(
        n13388) );
  AOI21_X1 U15519 ( .B1(n13556), .B2(n14900), .A(n13388), .ZN(n13389) );
  OAI21_X1 U15520 ( .B1(n13560), .B2(n14903), .A(n13389), .ZN(P2_U3240) );
  XNOR2_X1 U15521 ( .A(n13390), .B(n13391), .ZN(n13393) );
  AOI21_X1 U15522 ( .B1(n13393), .B2(n14886), .A(n13392), .ZN(n13567) );
  AOI21_X1 U15523 ( .B1(n13396), .B2(n13395), .A(n13394), .ZN(n13565) );
  OAI211_X1 U15524 ( .C1(n13563), .C2(n13415), .A(n13523), .B(n13397), .ZN(
        n13562) );
  INV_X1 U15525 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13398) );
  OAI22_X1 U15526 ( .A1(n13399), .A2(n13518), .B1(n13398), .B2(n14919), .ZN(
        n13400) );
  AOI21_X1 U15527 ( .B1(n13401), .B2(n14890), .A(n13400), .ZN(n13402) );
  OAI21_X1 U15528 ( .B1(n13562), .B2(n14898), .A(n13402), .ZN(n13403) );
  AOI21_X1 U15529 ( .B1(n13565), .B2(n14900), .A(n13403), .ZN(n13404) );
  OAI21_X1 U15530 ( .B1(n13567), .B2(n14903), .A(n13404), .ZN(P2_U3241) );
  INV_X1 U15531 ( .A(n13405), .ZN(n13408) );
  OAI21_X1 U15532 ( .B1(n13423), .B2(n13406), .A(n13413), .ZN(n13407) );
  AOI21_X1 U15533 ( .B1(n13408), .B2(n13407), .A(n7099), .ZN(n13411) );
  INV_X1 U15534 ( .A(n13409), .ZN(n13410) );
  NOR2_X1 U15535 ( .A1(n13411), .A2(n13410), .ZN(n13573) );
  OAI21_X1 U15536 ( .B1(n13414), .B2(n13413), .A(n13412), .ZN(n13568) );
  INV_X1 U15537 ( .A(n13415), .ZN(n13417) );
  AOI21_X1 U15538 ( .B1(n13429), .B2(n13569), .A(n13489), .ZN(n13416) );
  NAND2_X1 U15539 ( .A1(n13417), .A2(n13416), .ZN(n13572) );
  AOI22_X1 U15540 ( .A1(n13418), .A2(n14905), .B1(n13531), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n13420) );
  NAND2_X1 U15541 ( .A1(n13569), .A2(n14890), .ZN(n13419) );
  OAI211_X1 U15542 ( .C1(n13572), .C2(n14898), .A(n13420), .B(n13419), .ZN(
        n13421) );
  AOI21_X1 U15543 ( .B1(n13568), .B2(n14900), .A(n13421), .ZN(n13422) );
  OAI21_X1 U15544 ( .B1(n13573), .B2(n14903), .A(n13422), .ZN(P2_U3242) );
  AOI211_X1 U15545 ( .C1(n13425), .C2(n13424), .A(n7099), .B(n13423), .ZN(
        n13428) );
  INV_X1 U15546 ( .A(n13426), .ZN(n13427) );
  NOR2_X1 U15547 ( .A1(n13428), .A2(n13427), .ZN(n13577) );
  INV_X1 U15548 ( .A(n13429), .ZN(n13430) );
  AOI211_X1 U15549 ( .C1(n13575), .C2(n13445), .A(n13489), .B(n13430), .ZN(
        n13574) );
  AOI22_X1 U15550 ( .A1(n13531), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n13431), 
        .B2(n14905), .ZN(n13432) );
  OAI21_X1 U15551 ( .B1(n6950), .B2(n13472), .A(n13432), .ZN(n13438) );
  AND2_X1 U15552 ( .A1(n13434), .A2(n13433), .ZN(n13435) );
  OR2_X1 U15553 ( .A1(n13436), .A2(n13435), .ZN(n13578) );
  NOR2_X1 U15554 ( .A1(n13578), .A2(n13528), .ZN(n13437) );
  AOI211_X1 U15555 ( .C1(n13574), .C2(n14916), .A(n13438), .B(n13437), .ZN(
        n13439) );
  OAI21_X1 U15556 ( .B1(n13577), .B2(n14903), .A(n13439), .ZN(P2_U3243) );
  XNOR2_X1 U15557 ( .A(n13440), .B(n13441), .ZN(n13583) );
  XNOR2_X1 U15558 ( .A(n13442), .B(n13441), .ZN(n13444) );
  OAI21_X1 U15559 ( .B1(n13444), .B2(n7099), .A(n13443), .ZN(n13579) );
  INV_X1 U15560 ( .A(n13458), .ZN(n13446) );
  AOI211_X1 U15561 ( .C1(n13581), .C2(n13446), .A(n13105), .B(n6951), .ZN(
        n13580) );
  NAND2_X1 U15562 ( .A1(n13580), .A2(n14916), .ZN(n13449) );
  AOI22_X1 U15563 ( .A1(n13531), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n13447), 
        .B2(n14905), .ZN(n13448) );
  OAI211_X1 U15564 ( .C1(n13450), .C2(n13472), .A(n13449), .B(n13448), .ZN(
        n13451) );
  AOI21_X1 U15565 ( .B1(n13579), .B2(n14919), .A(n13451), .ZN(n13452) );
  OAI21_X1 U15566 ( .B1(n13528), .B2(n13583), .A(n13452), .ZN(P2_U3244) );
  XOR2_X1 U15567 ( .A(n13455), .B(n13453), .Z(n13588) );
  XOR2_X1 U15568 ( .A(n13455), .B(n13454), .Z(n13457) );
  OAI21_X1 U15569 ( .B1(n13457), .B2(n7099), .A(n13456), .ZN(n13584) );
  AOI211_X1 U15570 ( .C1(n13586), .C2(n13470), .A(n13489), .B(n13458), .ZN(
        n13585) );
  NAND2_X1 U15571 ( .A1(n13585), .A2(n14916), .ZN(n13461) );
  AOI22_X1 U15572 ( .A1(n13531), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13459), 
        .B2(n14905), .ZN(n13460) );
  OAI211_X1 U15573 ( .C1(n13462), .C2(n13472), .A(n13461), .B(n13460), .ZN(
        n13463) );
  AOI21_X1 U15574 ( .B1(n13584), .B2(n14919), .A(n13463), .ZN(n13464) );
  OAI21_X1 U15575 ( .B1(n13588), .B2(n13528), .A(n13464), .ZN(P2_U3245) );
  XNOR2_X1 U15576 ( .A(n13465), .B(n13466), .ZN(n13593) );
  XNOR2_X1 U15577 ( .A(n6539), .B(n13466), .ZN(n13468) );
  OAI21_X1 U15578 ( .B1(n13468), .B2(n7099), .A(n13467), .ZN(n13589) );
  NAND2_X1 U15579 ( .A1(n13589), .A2(n14919), .ZN(n13478) );
  INV_X1 U15580 ( .A(n13470), .ZN(n13471) );
  AOI211_X1 U15581 ( .C1(n13591), .C2(n13490), .A(n13105), .B(n13471), .ZN(
        n13590) );
  NOR2_X1 U15582 ( .A1(n9431), .A2(n13472), .ZN(n13476) );
  OAI22_X1 U15583 ( .A1(n14919), .A2(n13474), .B1(n13473), .B2(n13518), .ZN(
        n13475) );
  AOI211_X1 U15584 ( .C1(n13590), .C2(n14916), .A(n13476), .B(n13475), .ZN(
        n13477) );
  OAI211_X1 U15585 ( .C1(n13528), .C2(n13593), .A(n13478), .B(n13477), .ZN(
        P2_U3246) );
  XNOR2_X1 U15586 ( .A(n13480), .B(n13479), .ZN(n13482) );
  AOI21_X1 U15587 ( .B1(n13482), .B2(n14886), .A(n13481), .ZN(n13597) );
  INV_X1 U15588 ( .A(n13483), .ZN(n13484) );
  AOI21_X1 U15589 ( .B1(n7477), .B2(n13485), .A(n13484), .ZN(n13598) );
  INV_X1 U15590 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n13487) );
  OAI22_X1 U15591 ( .A1(n14919), .A2(n13487), .B1(n13486), .B2(n13518), .ZN(
        n13488) );
  AOI21_X1 U15592 ( .B1(n13595), .B2(n14890), .A(n13488), .ZN(n13493) );
  AOI21_X1 U15593 ( .B1(n13595), .B2(n13507), .A(n13489), .ZN(n13491) );
  AND2_X1 U15594 ( .A1(n13491), .A2(n13490), .ZN(n13594) );
  NAND2_X1 U15595 ( .A1(n13594), .A2(n14916), .ZN(n13492) );
  OAI211_X1 U15596 ( .C1(n13598), .C2(n13528), .A(n13493), .B(n13492), .ZN(
        n13494) );
  INV_X1 U15597 ( .A(n13494), .ZN(n13495) );
  OAI21_X1 U15598 ( .B1(n13531), .B2(n13597), .A(n13495), .ZN(P2_U3247) );
  XNOR2_X1 U15599 ( .A(n13496), .B(n13500), .ZN(n13498) );
  AOI21_X1 U15600 ( .B1(n13498), .B2(n14886), .A(n13497), .ZN(n13602) );
  OAI21_X1 U15601 ( .B1(n13501), .B2(n13500), .A(n13499), .ZN(n13603) );
  OAI22_X1 U15602 ( .A1(n14919), .A2(n13503), .B1(n13502), .B2(n13518), .ZN(
        n13504) );
  AOI21_X1 U15603 ( .B1(n13600), .B2(n14890), .A(n13504), .ZN(n13509) );
  OR2_X1 U15604 ( .A1(n6626), .A2(n13505), .ZN(n13506) );
  AND3_X1 U15605 ( .A1(n13507), .A2(n13523), .A3(n13506), .ZN(n13599) );
  NAND2_X1 U15606 ( .A1(n13599), .A2(n14916), .ZN(n13508) );
  OAI211_X1 U15607 ( .C1(n13603), .C2(n13528), .A(n13509), .B(n13508), .ZN(
        n13510) );
  INV_X1 U15608 ( .A(n13510), .ZN(n13511) );
  OAI21_X1 U15609 ( .B1(n13531), .B2(n13602), .A(n13511), .ZN(P2_U3248) );
  XNOR2_X1 U15610 ( .A(n13512), .B(n13515), .ZN(n13514) );
  AOI21_X1 U15611 ( .B1(n13514), .B2(n14886), .A(n13513), .ZN(n13608) );
  INV_X1 U15612 ( .A(n13515), .ZN(n13517) );
  OAI21_X1 U15613 ( .B1(n6631), .B2(n13517), .A(n13516), .ZN(n13604) );
  OAI22_X1 U15614 ( .A1(n14919), .A2(n13520), .B1(n13519), .B2(n13518), .ZN(
        n13521) );
  AOI21_X1 U15615 ( .B1(n13607), .B2(n14890), .A(n13521), .ZN(n13527) );
  NAND2_X1 U15616 ( .A1(n13522), .A2(n13607), .ZN(n13524) );
  NAND2_X1 U15617 ( .A1(n13524), .A2(n13523), .ZN(n13525) );
  NOR2_X1 U15618 ( .A1(n6626), .A2(n13525), .ZN(n13606) );
  NAND2_X1 U15619 ( .A1(n13606), .A2(n14916), .ZN(n13526) );
  OAI211_X1 U15620 ( .C1(n13604), .C2(n13528), .A(n13527), .B(n13526), .ZN(
        n13529) );
  INV_X1 U15621 ( .A(n13529), .ZN(n13530) );
  OAI21_X1 U15622 ( .B1(n13531), .B2(n13608), .A(n13530), .ZN(P2_U3249) );
  OAI211_X1 U15623 ( .C1(n13319), .C2(n14958), .A(n13532), .B(n13533), .ZN(
        n13618) );
  MUX2_X1 U15624 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13618), .S(n13616), .Z(
        P2_U3530) );
  OAI211_X1 U15625 ( .C1(n13535), .C2(n14958), .A(n13534), .B(n13533), .ZN(
        n13619) );
  MUX2_X1 U15626 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13619), .S(n13616), .Z(
        P2_U3529) );
  MUX2_X1 U15627 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13620), .S(n13616), .Z(
        P2_U3528) );
  OAI21_X1 U15628 ( .B1(n13614), .B2(n13545), .A(n13544), .ZN(n13621) );
  MUX2_X1 U15629 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13621), .S(n13616), .Z(
        P2_U3527) );
  AOI21_X1 U15630 ( .B1(n13547), .B2(n14945), .A(n13546), .ZN(n13548) );
  OAI211_X1 U15631 ( .C1(n13614), .C2(n13550), .A(n13549), .B(n13548), .ZN(
        n13622) );
  MUX2_X1 U15632 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13622), .S(n13616), .Z(
        P2_U3526) );
  AOI211_X1 U15633 ( .C1(n13553), .C2(n14945), .A(n13552), .B(n13551), .ZN(
        n13554) );
  OAI21_X1 U15634 ( .B1(n13614), .B2(n13555), .A(n13554), .ZN(n13623) );
  MUX2_X1 U15635 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13623), .S(n13616), .Z(
        P2_U3525) );
  INV_X1 U15636 ( .A(n13556), .ZN(n13561) );
  AOI21_X1 U15637 ( .B1(n13558), .B2(n14945), .A(n13557), .ZN(n13559) );
  OAI211_X1 U15638 ( .C1(n13614), .C2(n13561), .A(n13560), .B(n13559), .ZN(
        n13624) );
  MUX2_X1 U15639 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13624), .S(n13616), .Z(
        P2_U3524) );
  OAI21_X1 U15640 ( .B1(n13563), .B2(n14958), .A(n13562), .ZN(n13564) );
  AOI21_X1 U15641 ( .B1(n13565), .B2(n14961), .A(n13564), .ZN(n13566) );
  NAND2_X1 U15642 ( .A1(n13567), .A2(n13566), .ZN(n13625) );
  MUX2_X1 U15643 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13625), .S(n13616), .Z(
        P2_U3523) );
  NAND2_X1 U15644 ( .A1(n13568), .A2(n14961), .ZN(n13571) );
  NAND2_X1 U15645 ( .A1(n13569), .A2(n14945), .ZN(n13570) );
  NAND4_X1 U15646 ( .A1(n13573), .A2(n13572), .A3(n13571), .A4(n13570), .ZN(
        n13626) );
  MUX2_X1 U15647 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13626), .S(n13616), .Z(
        P2_U3522) );
  AOI21_X1 U15648 ( .B1(n13575), .B2(n14945), .A(n13574), .ZN(n13576) );
  OAI211_X1 U15649 ( .C1(n13614), .C2(n13578), .A(n13577), .B(n13576), .ZN(
        n13627) );
  MUX2_X1 U15650 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13627), .S(n13616), .Z(
        P2_U3521) );
  AOI211_X1 U15651 ( .C1(n13581), .C2(n14945), .A(n13580), .B(n13579), .ZN(
        n13582) );
  OAI21_X1 U15652 ( .B1(n13614), .B2(n13583), .A(n13582), .ZN(n13628) );
  MUX2_X1 U15653 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13628), .S(n13616), .Z(
        P2_U3520) );
  AOI211_X1 U15654 ( .C1(n13586), .C2(n14945), .A(n13585), .B(n13584), .ZN(
        n13587) );
  OAI21_X1 U15655 ( .B1(n13614), .B2(n13588), .A(n13587), .ZN(n13629) );
  MUX2_X1 U15656 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13629), .S(n13616), .Z(
        P2_U3519) );
  AOI211_X1 U15657 ( .C1(n13591), .C2(n14945), .A(n13590), .B(n13589), .ZN(
        n13592) );
  OAI21_X1 U15658 ( .B1(n13614), .B2(n13593), .A(n13592), .ZN(n13630) );
  MUX2_X1 U15659 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13630), .S(n13616), .Z(
        P2_U3518) );
  AOI21_X1 U15660 ( .B1(n13595), .B2(n14945), .A(n13594), .ZN(n13596) );
  OAI211_X1 U15661 ( .C1(n13598), .C2(n13614), .A(n13597), .B(n13596), .ZN(
        n13631) );
  MUX2_X1 U15662 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13631), .S(n13616), .Z(
        P2_U3517) );
  AOI21_X1 U15663 ( .B1(n13600), .B2(n14945), .A(n13599), .ZN(n13601) );
  OAI211_X1 U15664 ( .C1(n13603), .C2(n13614), .A(n13602), .B(n13601), .ZN(
        n13632) );
  MUX2_X1 U15665 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13632), .S(n13616), .Z(
        P2_U3516) );
  NOR2_X1 U15666 ( .A1(n13604), .A2(n13614), .ZN(n13605) );
  AOI211_X1 U15667 ( .C1(n13607), .C2(n14945), .A(n13606), .B(n13605), .ZN(
        n13609) );
  NAND2_X1 U15668 ( .A1(n13609), .A2(n13608), .ZN(n13633) );
  MUX2_X1 U15669 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13633), .S(n13616), .Z(
        P2_U3515) );
  AOI21_X1 U15670 ( .B1(n13611), .B2(n14945), .A(n13610), .ZN(n13612) );
  OAI211_X1 U15671 ( .C1(n13615), .C2(n13614), .A(n13613), .B(n13612), .ZN(
        n13634) );
  MUX2_X1 U15672 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13634), .S(n13616), .Z(
        P2_U3514) );
  MUX2_X1 U15673 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n13617), .S(n13616), .Z(
        P2_U3503) );
  MUX2_X1 U15674 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13618), .S(n14964), .Z(
        P2_U3498) );
  MUX2_X1 U15675 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13619), .S(n14964), .Z(
        P2_U3497) );
  MUX2_X1 U15676 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13620), .S(n14964), .Z(
        P2_U3496) );
  MUX2_X1 U15677 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13621), .S(n14964), .Z(
        P2_U3495) );
  MUX2_X1 U15678 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13622), .S(n14964), .Z(
        P2_U3494) );
  MUX2_X1 U15679 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13623), .S(n14964), .Z(
        P2_U3493) );
  MUX2_X1 U15680 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13624), .S(n14964), .Z(
        P2_U3492) );
  MUX2_X1 U15681 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13625), .S(n14964), .Z(
        P2_U3491) );
  MUX2_X1 U15682 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13626), .S(n14964), .Z(
        P2_U3490) );
  MUX2_X1 U15683 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13627), .S(n14964), .Z(
        P2_U3489) );
  MUX2_X1 U15684 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13628), .S(n14964), .Z(
        P2_U3488) );
  MUX2_X1 U15685 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13629), .S(n14964), .Z(
        P2_U3487) );
  MUX2_X1 U15686 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13630), .S(n14964), .Z(
        P2_U3486) );
  MUX2_X1 U15687 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13631), .S(n14964), .Z(
        P2_U3484) );
  MUX2_X1 U15688 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13632), .S(n14964), .Z(
        P2_U3481) );
  MUX2_X1 U15689 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13633), .S(n14964), .Z(
        P2_U3478) );
  MUX2_X1 U15690 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13634), .S(n14964), .Z(
        P2_U3475) );
  INV_X1 U15691 ( .A(n13635), .ZN(n14204) );
  NOR4_X1 U15692 ( .A1(n13638), .A2(P2_IR_REG_30__SCAN_IN), .A3(n13637), .A4(
        P2_U3088), .ZN(n13639) );
  AOI21_X1 U15693 ( .B1(n13645), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n13639), 
        .ZN(n13640) );
  OAI21_X1 U15694 ( .B1(n14204), .B2(n13643), .A(n13640), .ZN(P2_U3296) );
  OAI222_X1 U15695 ( .A1(P2_U3088), .A2(n8980), .B1(n13643), .B2(n13642), .C1(
        n13641), .C2(n13652), .ZN(P2_U3298) );
  AOI21_X1 U15696 ( .B1(n13645), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13644), 
        .ZN(n13646) );
  OAI21_X1 U15697 ( .B1(n13647), .B2(n13643), .A(n13646), .ZN(P2_U3299) );
  INV_X1 U15698 ( .A(n13648), .ZN(n14207) );
  OAI222_X1 U15699 ( .A1(n13650), .A2(P2_U3088), .B1(n13643), .B2(n14207), 
        .C1(n13649), .C2(n13652), .ZN(P2_U3300) );
  INV_X1 U15700 ( .A(n13651), .ZN(n14213) );
  OAI222_X1 U15701 ( .A1(P2_U3088), .A2(n13654), .B1(n13643), .B2(n14213), 
        .C1(n13653), .C2(n13652), .ZN(P2_U3301) );
  INV_X1 U15702 ( .A(n13655), .ZN(n13656) );
  MUX2_X1 U15703 ( .A(n13656), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  OAI21_X1 U15704 ( .B1(n13659), .B2(n13658), .A(n13657), .ZN(n13660) );
  OAI22_X1 U15705 ( .A1(n13662), .A2(n14055), .B1(n13661), .B2(n14053), .ZN(
        n13942) );
  INV_X1 U15706 ( .A(n13945), .ZN(n13664) );
  OAI22_X1 U15707 ( .A1(n13664), .A2(n13813), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13663), .ZN(n13665) );
  AOI21_X1 U15708 ( .B1(n13942), .B2(n13769), .A(n13665), .ZN(n13666) );
  INV_X1 U15709 ( .A(n14138), .ZN(n13996) );
  INV_X1 U15710 ( .A(n13667), .ZN(n13670) );
  NOR3_X1 U15711 ( .A1(n13670), .A2(n13669), .A3(n13668), .ZN(n13672) );
  INV_X1 U15712 ( .A(n13671), .ZN(n13750) );
  OAI21_X1 U15713 ( .B1(n13672), .B2(n13750), .A(n13795), .ZN(n13678) );
  NAND2_X1 U15714 ( .A1(n13824), .A2(n14631), .ZN(n13674) );
  NAND2_X1 U15715 ( .A1(n13826), .A2(n14482), .ZN(n13673) );
  NAND2_X1 U15716 ( .A1(n13674), .A2(n13673), .ZN(n13990) );
  OAI22_X1 U15717 ( .A1(n13993), .A2(n13813), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13675), .ZN(n13676) );
  AOI21_X1 U15718 ( .B1(n13990), .B2(n13769), .A(n13676), .ZN(n13677) );
  OAI211_X1 U15719 ( .C1(n13996), .C2(n13803), .A(n13678), .B(n13677), .ZN(
        P1_U3216) );
  AND2_X1 U15720 ( .A1(n13782), .A2(n13679), .ZN(n13682) );
  OAI211_X1 U15721 ( .C1(n13682), .C2(n13681), .A(n13795), .B(n13680), .ZN(
        n13686) );
  NAND2_X1 U15722 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13927)
         );
  OAI21_X1 U15723 ( .B1(n14054), .B2(n13808), .A(n13927), .ZN(n13684) );
  NOR2_X1 U15724 ( .A1(n13813), .A2(n14060), .ZN(n13683) );
  AOI211_X1 U15725 ( .C1(n13810), .C2(n13828), .A(n13684), .B(n13683), .ZN(
        n13685) );
  OAI211_X1 U15726 ( .C1(n10006), .C2(n13803), .A(n13686), .B(n13685), .ZN(
        P1_U3219) );
  OAI21_X1 U15727 ( .B1(n13689), .B2(n13688), .A(n13687), .ZN(n13690) );
  NAND2_X1 U15728 ( .A1(n13690), .A2(n13795), .ZN(n13695) );
  OAI22_X1 U15729 ( .A1(n13691), .A2(n14055), .B1(n14056), .B2(n14053), .ZN(
        n14150) );
  OAI22_X1 U15730 ( .A1(n13813), .A2(n14025), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13692), .ZN(n13693) );
  AOI21_X1 U15731 ( .B1(n14150), .B2(n13769), .A(n13693), .ZN(n13694) );
  OAI211_X1 U15732 ( .C1(n14029), .C2(n13803), .A(n13695), .B(n13694), .ZN(
        P1_U3223) );
  INV_X1 U15733 ( .A(n14125), .ZN(n13709) );
  INV_X1 U15734 ( .A(n13696), .ZN(n13751) );
  INV_X1 U15735 ( .A(n13697), .ZN(n13699) );
  NOR3_X1 U15736 ( .A1(n13751), .A2(n13699), .A3(n13698), .ZN(n13702) );
  INV_X1 U15737 ( .A(n13700), .ZN(n13701) );
  OAI21_X1 U15738 ( .B1(n13702), .B2(n13701), .A(n13795), .ZN(n13708) );
  AOI22_X1 U15739 ( .A1(n13703), .A2(n13798), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13704) );
  OAI21_X1 U15740 ( .B1(n13705), .B2(n13808), .A(n13704), .ZN(n13706) );
  AOI21_X1 U15741 ( .B1(n13810), .B2(n13822), .A(n13706), .ZN(n13707) );
  OAI211_X1 U15742 ( .C1(n13709), .C2(n13803), .A(n13708), .B(n13707), .ZN(
        P1_U3225) );
  AOI21_X1 U15743 ( .B1(n13712), .B2(n13711), .A(n13710), .ZN(n13721) );
  OAI21_X1 U15744 ( .B1(n13808), .B2(n13714), .A(n13713), .ZN(n13715) );
  AOI21_X1 U15745 ( .B1(n13810), .B2(n14074), .A(n13715), .ZN(n13716) );
  OAI21_X1 U15746 ( .B1(n13813), .B2(n13717), .A(n13716), .ZN(n13718) );
  AOI21_X1 U15747 ( .B1(n13719), .B2(n13815), .A(n13718), .ZN(n13720) );
  OAI21_X1 U15748 ( .B1(n13721), .B2(n13817), .A(n13720), .ZN(P1_U3226) );
  OAI21_X1 U15749 ( .B1(n13724), .B2(n13723), .A(n13722), .ZN(n13725) );
  NAND2_X1 U15750 ( .A1(n13725), .A2(n13795), .ZN(n13733) );
  AOI22_X1 U15751 ( .A1(n13810), .A2(n13838), .B1(n13815), .B2(n14724), .ZN(
        n13732) );
  INV_X1 U15752 ( .A(n13726), .ZN(n13730) );
  OAI21_X1 U15753 ( .B1(n13808), .B2(n13728), .A(n13727), .ZN(n13729) );
  AOI21_X1 U15754 ( .B1(n13730), .B2(n13798), .A(n13729), .ZN(n13731) );
  NAND3_X1 U15755 ( .A1(n13733), .A2(n13732), .A3(n13731), .ZN(P1_U3227) );
  INV_X1 U15756 ( .A(n13734), .ZN(n14179) );
  INV_X1 U15757 ( .A(n13735), .ZN(n13739) );
  NOR3_X1 U15758 ( .A1(n13710), .A2(n13737), .A3(n13736), .ZN(n13738) );
  OAI21_X1 U15759 ( .B1(n13739), .B2(n13738), .A(n13795), .ZN(n13746) );
  OAI21_X1 U15760 ( .B1(n13808), .B2(n13741), .A(n13740), .ZN(n13744) );
  NOR2_X1 U15761 ( .A1(n13813), .A2(n13742), .ZN(n13743) );
  AOI211_X1 U15762 ( .C1(n13810), .C2(n13829), .A(n13744), .B(n13743), .ZN(
        n13745) );
  OAI211_X1 U15763 ( .C1(n14179), .C2(n13803), .A(n13746), .B(n13745), .ZN(
        P1_U3228) );
  INV_X1 U15764 ( .A(n13747), .ZN(n13749) );
  NOR3_X1 U15765 ( .A1(n13750), .A2(n13749), .A3(n13748), .ZN(n13752) );
  OAI21_X1 U15766 ( .B1(n13752), .B2(n13751), .A(n13795), .ZN(n13758) );
  OAI22_X1 U15767 ( .A1(n13958), .A2(n14055), .B1(n13753), .B2(n14053), .ZN(
        n13973) );
  INV_X1 U15768 ( .A(n13979), .ZN(n13755) );
  OAI22_X1 U15769 ( .A1(n13755), .A2(n13813), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13754), .ZN(n13756) );
  AOI21_X1 U15770 ( .B1(n13973), .B2(n13769), .A(n13756), .ZN(n13757) );
  OAI211_X1 U15771 ( .C1(n13981), .C2(n13803), .A(n13758), .B(n13757), .ZN(
        P1_U3229) );
  INV_X1 U15772 ( .A(n13759), .ZN(n13761) );
  NAND2_X1 U15773 ( .A1(n13761), .A2(n13760), .ZN(n13763) );
  XNOR2_X1 U15774 ( .A(n13763), .B(n13762), .ZN(n13764) );
  NAND2_X1 U15775 ( .A1(n13764), .A2(n13795), .ZN(n13773) );
  AOI22_X1 U15776 ( .A1(n13815), .A2(n13765), .B1(P1_REG3_REG_4__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13772) );
  INV_X1 U15777 ( .A(n14656), .ZN(n13766) );
  NAND2_X1 U15778 ( .A1(n13798), .A2(n13766), .ZN(n13771) );
  NAND2_X1 U15779 ( .A1(n13839), .A2(n14631), .ZN(n13768) );
  NAND2_X1 U15780 ( .A1(n13841), .A2(n14482), .ZN(n13767) );
  NAND2_X1 U15781 ( .A1(n13768), .A2(n13767), .ZN(n14652) );
  NAND2_X1 U15782 ( .A1(n14652), .A2(n13769), .ZN(n13770) );
  NAND4_X1 U15783 ( .A1(n13773), .A2(n13772), .A3(n13771), .A4(n13770), .ZN(
        P1_U3230) );
  XNOR2_X1 U15784 ( .A(n13775), .B(n13774), .ZN(n13781) );
  AND2_X1 U15785 ( .A1(n14075), .A2(n14482), .ZN(n13776) );
  AOI21_X1 U15786 ( .B1(n13827), .B2(n14631), .A(n13776), .ZN(n14157) );
  AOI22_X1 U15787 ( .A1(n13798), .A2(n14036), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13777) );
  OAI21_X1 U15788 ( .B1(n14157), .B2(n13778), .A(n13777), .ZN(n13779) );
  AOI21_X1 U15789 ( .B1(n14159), .B2(n13815), .A(n13779), .ZN(n13780) );
  OAI21_X1 U15790 ( .B1(n13781), .B2(n13817), .A(n13780), .ZN(P1_U3233) );
  INV_X1 U15791 ( .A(n14172), .ZN(n13791) );
  OAI21_X1 U15792 ( .B1(n13784), .B2(n13783), .A(n13782), .ZN(n13785) );
  NAND2_X1 U15793 ( .A1(n13785), .A2(n13795), .ZN(n13790) );
  NAND2_X1 U15794 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14613)
         );
  OAI21_X1 U15795 ( .B1(n13786), .B2(n13808), .A(n14613), .ZN(n13788) );
  NOR2_X1 U15796 ( .A1(n13813), .A2(n14079), .ZN(n13787) );
  AOI211_X1 U15797 ( .C1(n13810), .C2(n14075), .A(n13788), .B(n13787), .ZN(
        n13789) );
  OAI211_X1 U15798 ( .C1(n13791), .C2(n13803), .A(n13790), .B(n13789), .ZN(
        P1_U3238) );
  OAI21_X1 U15799 ( .B1(n13794), .B2(n13793), .A(n13792), .ZN(n13796) );
  NAND2_X1 U15800 ( .A1(n13796), .A2(n13795), .ZN(n13802) );
  INV_X1 U15801 ( .A(n13797), .ZN(n13966) );
  AOI22_X1 U15802 ( .A1(n13966), .A2(n13798), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13799) );
  OAI21_X1 U15803 ( .B1(n13958), .B2(n13808), .A(n13799), .ZN(n13800) );
  AOI21_X1 U15804 ( .B1(n13810), .B2(n13956), .A(n13800), .ZN(n13801) );
  OAI211_X1 U15805 ( .C1(n14117), .C2(n13803), .A(n13802), .B(n13801), .ZN(
        P1_U3240) );
  XNOR2_X1 U15806 ( .A(n13805), .B(n13804), .ZN(n13818) );
  OAI22_X1 U15807 ( .A1(n13808), .A2(n13807), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13806), .ZN(n13809) );
  AOI21_X1 U15808 ( .B1(n13810), .B2(n13830), .A(n13809), .ZN(n13811) );
  OAI21_X1 U15809 ( .B1(n13813), .B2(n13812), .A(n13811), .ZN(n13814) );
  AOI21_X1 U15810 ( .B1(n14503), .B2(n13815), .A(n13814), .ZN(n13816) );
  OAI21_X1 U15811 ( .B1(n13818), .B2(n13817), .A(n13816), .ZN(P1_U3241) );
  MUX2_X1 U15812 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n13932), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U15813 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13819), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U15814 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13820), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15815 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n13821), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15816 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13956), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15817 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n13822), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15818 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n13823), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15819 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n13824), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15820 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n13825), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U15821 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n13826), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U15822 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n13827), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U15823 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13828), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15824 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14075), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15825 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n13829), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U15826 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14074), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U15827 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n13830), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U15828 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13831), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15829 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13832), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15830 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14483), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U15831 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13833), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U15832 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14630), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U15833 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13834), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U15834 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13835), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U15835 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13836), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U15836 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13837), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U15837 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13838), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U15838 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13839), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U15839 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13840), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U15840 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13841), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U15841 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n13842), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U15842 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n7573), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U15843 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n13843), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI211_X1 U15844 ( .C1(n13858), .C2(n13845), .A(n14606), .B(n13844), .ZN(
        n13855) );
  AOI22_X1 U15845 ( .A1(n14587), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n13854) );
  NAND2_X1 U15846 ( .A1(n14591), .A2(n13846), .ZN(n13853) );
  INV_X1 U15847 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n14762) );
  INV_X1 U15848 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n13849) );
  MUX2_X1 U15849 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10128), .S(n13847), .Z(
        n13848) );
  OAI21_X1 U15850 ( .B1(n14762), .B2(n13849), .A(n13848), .ZN(n13850) );
  NAND3_X1 U15851 ( .A1(n14603), .A2(n13851), .A3(n13850), .ZN(n13852) );
  NAND4_X1 U15852 ( .A1(n13855), .A2(n13854), .A3(n13853), .A4(n13852), .ZN(
        P1_U3244) );
  NOR2_X1 U15853 ( .A1(n14206), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n13856) );
  NOR2_X1 U15854 ( .A1(n13856), .A2(n8325), .ZN(n14561) );
  MUX2_X1 U15855 ( .A(n13858), .B(n13857), .S(n14206), .Z(n13860) );
  NAND2_X1 U15856 ( .A1(n13860), .A2(n13859), .ZN(n13861) );
  OAI211_X1 U15857 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n14561), .A(n13861), .B(
        P1_U4016), .ZN(n14585) );
  AOI22_X1 U15858 ( .A1(n14587), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n13871) );
  OAI211_X1 U15859 ( .C1(n13863), .C2(n13862), .A(n14603), .B(n13877), .ZN(
        n13867) );
  OAI211_X1 U15860 ( .C1(n13865), .C2(n13864), .A(n14606), .B(n13882), .ZN(
        n13866) );
  OAI211_X1 U15861 ( .C1(n14611), .C2(n13868), .A(n13867), .B(n13866), .ZN(
        n13869) );
  INV_X1 U15862 ( .A(n13869), .ZN(n13870) );
  NAND3_X1 U15863 ( .A1(n14585), .A2(n13871), .A3(n13870), .ZN(P1_U3245) );
  INV_X1 U15864 ( .A(n13879), .ZN(n13874) );
  OAI22_X1 U15865 ( .A1(n14615), .A2(n14222), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13872), .ZN(n13873) );
  AOI21_X1 U15866 ( .B1(n13874), .B2(n14591), .A(n13873), .ZN(n13886) );
  MUX2_X1 U15867 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10135), .S(n13879), .Z(
        n13875) );
  NAND3_X1 U15868 ( .A1(n13877), .A2(n13876), .A3(n13875), .ZN(n13878) );
  NAND3_X1 U15869 ( .A1(n14603), .A2(n14577), .A3(n13878), .ZN(n13885) );
  MUX2_X1 U15870 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n14674), .S(n13879), .Z(
        n13880) );
  NAND3_X1 U15871 ( .A1(n13882), .A2(n13881), .A3(n13880), .ZN(n13883) );
  NAND3_X1 U15872 ( .A1(n14606), .A2(n14569), .A3(n13883), .ZN(n13884) );
  NAND3_X1 U15873 ( .A1(n13886), .A2(n13885), .A3(n13884), .ZN(P1_U3246) );
  INV_X1 U15874 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n13888) );
  OAI21_X1 U15875 ( .B1(n14615), .B2(n13888), .A(n13887), .ZN(n13889) );
  AOI21_X1 U15876 ( .B1(n13890), .B2(n14591), .A(n13889), .ZN(n13903) );
  MUX2_X1 U15877 ( .A(n10142), .B(P1_REG1_REG_7__SCAN_IN), .S(n13890), .Z(
        n13891) );
  NAND3_X1 U15878 ( .A1(n13893), .A2(n13892), .A3(n13891), .ZN(n13894) );
  NAND3_X1 U15879 ( .A1(n14603), .A2(n13895), .A3(n13894), .ZN(n13902) );
  OR3_X1 U15880 ( .A1(n13898), .A2(n13897), .A3(n13896), .ZN(n13899) );
  NAND3_X1 U15881 ( .A1(n14606), .A2(n13900), .A3(n13899), .ZN(n13901) );
  NAND3_X1 U15882 ( .A1(n13903), .A2(n13902), .A3(n13901), .ZN(P1_U3250) );
  INV_X1 U15883 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n13906) );
  OAI21_X1 U15884 ( .B1(n13906), .B2(n13905), .A(n13904), .ZN(n13907) );
  XOR2_X1 U15885 ( .A(n13916), .B(n13907), .Z(n14604) );
  NAND2_X1 U15886 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n14604), .ZN(n14602) );
  NAND2_X1 U15887 ( .A1(n13907), .A2(n13916), .ZN(n13908) );
  NAND2_X1 U15888 ( .A1(n14602), .A2(n13908), .ZN(n13910) );
  INV_X1 U15889 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n13909) );
  XNOR2_X1 U15890 ( .A(n13910), .B(n13909), .ZN(n13924) );
  INV_X1 U15891 ( .A(n13924), .ZN(n13922) );
  INV_X1 U15892 ( .A(n13911), .ZN(n13912) );
  NAND2_X1 U15893 ( .A1(n13913), .A2(n13912), .ZN(n13914) );
  NAND2_X1 U15894 ( .A1(n13915), .A2(n13914), .ZN(n13917) );
  XOR2_X1 U15895 ( .A(n13916), .B(n13917), .Z(n14607) );
  NAND2_X1 U15896 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n14607), .ZN(n14605) );
  NAND2_X1 U15897 ( .A1(n13917), .A2(n13916), .ZN(n13918) );
  NAND2_X1 U15898 ( .A1(n14605), .A2(n13918), .ZN(n13919) );
  XOR2_X1 U15899 ( .A(n13919), .B(P1_REG2_REG_19__SCAN_IN), .Z(n13923) );
  NOR2_X1 U15900 ( .A1(n13923), .A2(n13920), .ZN(n13921) );
  AOI211_X1 U15901 ( .C1(n13922), .C2(n14603), .A(n14591), .B(n13921), .ZN(
        n13926) );
  AOI22_X1 U15902 ( .A1(n13924), .A2(n14603), .B1(n14606), .B2(n13923), .ZN(
        n13925) );
  MUX2_X1 U15903 ( .A(n13926), .B(n13925), .S(n8333), .Z(n13928) );
  OAI211_X1 U15904 ( .C1(n7529), .C2(n14615), .A(n13928), .B(n13927), .ZN(
        P1_U3262) );
  NAND2_X1 U15905 ( .A1(n14089), .A2(n14491), .ZN(n13934) );
  NAND2_X1 U15906 ( .A1(n13932), .A2(n13931), .ZN(n14092) );
  NOR2_X1 U15907 ( .A1(n14644), .A2(n14092), .ZN(n13938) );
  AOI21_X1 U15908 ( .B1(n14087), .B2(P1_REG2_REG_31__SCAN_IN), .A(n13938), 
        .ZN(n13933) );
  OAI211_X1 U15909 ( .C1(n14091), .C2(n14488), .A(n13934), .B(n13933), .ZN(
        P1_U3263) );
  XNOR2_X1 U15910 ( .A(n14094), .B(n13935), .ZN(n13936) );
  NAND2_X1 U15911 ( .A1(n13936), .A2(n14679), .ZN(n14093) );
  NOR2_X1 U15912 ( .A1(n14094), .A2(n14488), .ZN(n13937) );
  AOI211_X1 U15913 ( .C1(n14087), .C2(P1_REG2_REG_30__SCAN_IN), .A(n13938), 
        .B(n13937), .ZN(n13939) );
  OAI21_X1 U15914 ( .B1(n14065), .B2(n14093), .A(n13939), .ZN(P1_U3264) );
  XNOR2_X1 U15915 ( .A(n13941), .B(n13940), .ZN(n13943) );
  AOI211_X1 U15916 ( .C1(n14112), .C2(n13965), .A(n14699), .B(n13944), .ZN(
        n14111) );
  AOI22_X1 U15917 ( .A1(n13945), .A2(n14643), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n14087), .ZN(n13946) );
  OAI21_X1 U15918 ( .B1(n6872), .B2(n14488), .A(n13946), .ZN(n13952) );
  INV_X1 U15919 ( .A(n13947), .ZN(n13948) );
  AOI21_X1 U15920 ( .B1(n13950), .B2(n13949), .A(n13948), .ZN(n14115) );
  NOR2_X1 U15921 ( .A1(n14115), .A2(n14083), .ZN(n13951) );
  OAI21_X1 U15922 ( .B1(n14644), .B2(n14114), .A(n13953), .ZN(P1_U3266) );
  XNOR2_X1 U15923 ( .A(n13955), .B(n13954), .ZN(n13960) );
  NAND2_X1 U15924 ( .A1(n13956), .A2(n14631), .ZN(n13957) );
  OAI21_X1 U15925 ( .B1(n13958), .B2(n14053), .A(n13957), .ZN(n13959) );
  AOI21_X1 U15926 ( .B1(n13960), .B2(n14618), .A(n13959), .ZN(n14121) );
  OR2_X1 U15927 ( .A1(n13962), .A2(n13961), .ZN(n13963) );
  AND2_X1 U15928 ( .A1(n13964), .A2(n13963), .ZN(n14119) );
  OAI211_X1 U15929 ( .C1(n14117), .C2(n6531), .A(n14679), .B(n13965), .ZN(
        n14116) );
  AOI22_X1 U15930 ( .A1(n13966), .A2(n14643), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n14087), .ZN(n13969) );
  NAND2_X1 U15931 ( .A1(n13967), .A2(n14677), .ZN(n13968) );
  OAI211_X1 U15932 ( .C1(n14116), .C2(n14065), .A(n13969), .B(n13968), .ZN(
        n13970) );
  AOI21_X1 U15933 ( .B1(n14119), .B2(n14662), .A(n13970), .ZN(n13971) );
  OAI21_X1 U15934 ( .B1(n14121), .B2(n14644), .A(n13971), .ZN(P1_U3267) );
  AOI21_X1 U15935 ( .B1(n13972), .B2(n13983), .A(n14690), .ZN(n13975) );
  AOI21_X1 U15936 ( .B1(n13975), .B2(n13974), .A(n13973), .ZN(n14135) );
  INV_X1 U15937 ( .A(n13976), .ZN(n13977) );
  AOI211_X1 U15938 ( .C1(n14133), .C2(n13978), .A(n14699), .B(n13977), .ZN(
        n14132) );
  AOI22_X1 U15939 ( .A1(n13979), .A2(n14643), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n14087), .ZN(n13980) );
  OAI21_X1 U15940 ( .B1(n13981), .B2(n14488), .A(n13980), .ZN(n13987) );
  OAI21_X1 U15941 ( .B1(n13984), .B2(n13983), .A(n13982), .ZN(n13985) );
  INV_X1 U15942 ( .A(n13985), .ZN(n14136) );
  NOR2_X1 U15943 ( .A1(n14136), .A2(n14083), .ZN(n13986) );
  AOI211_X1 U15944 ( .C1(n14132), .C2(n14683), .A(n13987), .B(n13986), .ZN(
        n13988) );
  OAI21_X1 U15945 ( .B1(n14087), .B2(n14135), .A(n13988), .ZN(P1_U3269) );
  XNOR2_X1 U15946 ( .A(n13989), .B(n13997), .ZN(n13991) );
  AOI21_X1 U15947 ( .B1(n13991), .B2(n14618), .A(n13990), .ZN(n14140) );
  AOI211_X1 U15948 ( .C1(n14138), .C2(n14008), .A(n14699), .B(n13992), .ZN(
        n14137) );
  INV_X1 U15949 ( .A(n13993), .ZN(n13994) );
  AOI22_X1 U15950 ( .A1(n13994), .A2(n14643), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n14087), .ZN(n13995) );
  OAI21_X1 U15951 ( .B1(n13996), .B2(n14488), .A(n13995), .ZN(n14002) );
  NAND2_X1 U15952 ( .A1(n13998), .A2(n13997), .ZN(n13999) );
  NAND2_X1 U15953 ( .A1(n14000), .A2(n13999), .ZN(n14141) );
  NOR2_X1 U15954 ( .A1(n14141), .A2(n14083), .ZN(n14001) );
  AOI211_X1 U15955 ( .C1(n14137), .C2(n14683), .A(n14002), .B(n14001), .ZN(
        n14003) );
  OAI21_X1 U15956 ( .B1(n14140), .B2(n14644), .A(n14003), .ZN(P1_U3270) );
  XNOR2_X1 U15957 ( .A(n14004), .B(n14006), .ZN(n14148) );
  OAI21_X1 U15958 ( .B1(n14007), .B2(n14006), .A(n14005), .ZN(n14146) );
  OAI211_X1 U15959 ( .C1(n8295), .C2(n14027), .A(n14679), .B(n14008), .ZN(
        n14144) );
  INV_X1 U15960 ( .A(n8295), .ZN(n14014) );
  INV_X1 U15961 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n14012) );
  AND2_X1 U15962 ( .A1(n14009), .A2(n14643), .ZN(n14010) );
  OAI21_X1 U15963 ( .B1(n14142), .B2(n14010), .A(n14665), .ZN(n14011) );
  OAI21_X1 U15964 ( .B1(n14665), .B2(n14012), .A(n14011), .ZN(n14013) );
  AOI21_X1 U15965 ( .B1(n14014), .B2(n14677), .A(n14013), .ZN(n14015) );
  OAI21_X1 U15966 ( .B1(n14144), .B2(n14065), .A(n14015), .ZN(n14016) );
  AOI21_X1 U15967 ( .B1(n14146), .B2(n14035), .A(n14016), .ZN(n14017) );
  OAI21_X1 U15968 ( .B1(n14148), .B2(n14083), .A(n14017), .ZN(P1_U3271) );
  INV_X1 U15969 ( .A(n14018), .ZN(n14019) );
  AOI21_X1 U15970 ( .B1(n14022), .B2(n14020), .A(n14019), .ZN(n14154) );
  OAI211_X1 U15971 ( .C1(n14023), .C2(n14022), .A(n14021), .B(n14618), .ZN(
        n14152) );
  INV_X1 U15972 ( .A(n14150), .ZN(n14024) );
  OAI211_X1 U15973 ( .C1(n14673), .C2(n14025), .A(n14152), .B(n14024), .ZN(
        n14026) );
  NAND2_X1 U15974 ( .A1(n14026), .A2(n14665), .ZN(n14032) );
  AOI211_X1 U15975 ( .C1(n14151), .C2(n14041), .A(n14699), .B(n14027), .ZN(
        n14149) );
  INV_X1 U15976 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n14028) );
  OAI22_X1 U15977 ( .A1(n14029), .A2(n14488), .B1(n14028), .B2(n14665), .ZN(
        n14030) );
  AOI21_X1 U15978 ( .B1(n14149), .B2(n14683), .A(n14030), .ZN(n14031) );
  OAI211_X1 U15979 ( .C1(n14154), .C2(n14083), .A(n14032), .B(n14031), .ZN(
        P1_U3272) );
  NAND2_X1 U15980 ( .A1(n14034), .A2(n14033), .ZN(n14155) );
  NAND3_X1 U15981 ( .A1(n14156), .A2(n14155), .A3(n14035), .ZN(n14047) );
  AOI22_X1 U15982 ( .A1(P1_REG2_REG_20__SCAN_IN), .A2(n14644), .B1(n14036), 
        .B2(n14643), .ZN(n14037) );
  OAI21_X1 U15983 ( .B1(n14157), .B2(n14087), .A(n14037), .ZN(n14038) );
  AOI21_X1 U15984 ( .B1(n14159), .B2(n14677), .A(n14038), .ZN(n14046) );
  NAND2_X1 U15985 ( .A1(n14040), .A2(n14039), .ZN(n14160) );
  NAND3_X1 U15986 ( .A1(n6480), .A2(n14160), .A3(n14662), .ZN(n14045) );
  AOI21_X1 U15987 ( .B1(n14159), .B2(n14058), .A(n14699), .ZN(n14042) );
  NAND2_X1 U15988 ( .A1(n14042), .A2(n14041), .ZN(n14162) );
  INV_X1 U15989 ( .A(n14162), .ZN(n14043) );
  NAND2_X1 U15990 ( .A1(n14043), .A2(n14683), .ZN(n14044) );
  NAND4_X1 U15991 ( .A1(n14047), .A2(n14046), .A3(n14045), .A4(n14044), .ZN(
        P1_U3273) );
  XNOR2_X1 U15992 ( .A(n14049), .B(n14048), .ZN(n14170) );
  XNOR2_X1 U15993 ( .A(n14050), .B(n14051), .ZN(n14168) );
  AOI21_X1 U15994 ( .B1(n14062), .B2(n14069), .A(n14699), .ZN(n14059) );
  OAI22_X1 U15995 ( .A1(n14056), .A2(n14055), .B1(n14054), .B2(n14053), .ZN(
        n14057) );
  AOI21_X1 U15996 ( .B1(n14059), .B2(n14058), .A(n14057), .ZN(n14166) );
  INV_X1 U15997 ( .A(n14060), .ZN(n14061) );
  AOI22_X1 U15998 ( .A1(n14644), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14061), 
        .B2(n14643), .ZN(n14064) );
  NAND2_X1 U15999 ( .A1(n14062), .A2(n14677), .ZN(n14063) );
  OAI211_X1 U16000 ( .C1(n14166), .C2(n14065), .A(n14064), .B(n14063), .ZN(
        n14066) );
  AOI21_X1 U16001 ( .B1(n14168), .B2(n14662), .A(n14066), .ZN(n14067) );
  OAI21_X1 U16002 ( .B1(n14170), .B2(n14068), .A(n14067), .ZN(P1_U3274) );
  AOI211_X1 U16003 ( .C1(n14172), .C2(n14070), .A(n14699), .B(n14052), .ZN(
        n14171) );
  OAI211_X1 U16004 ( .C1(n14073), .C2(n14072), .A(n14071), .B(n14618), .ZN(
        n14077) );
  AOI22_X1 U16005 ( .A1(n14075), .A2(n14631), .B1(n14482), .B2(n14074), .ZN(
        n14076) );
  AND2_X1 U16006 ( .A1(n14077), .A2(n14076), .ZN(n14174) );
  INV_X1 U16007 ( .A(n14174), .ZN(n14078) );
  AOI21_X1 U16008 ( .B1(n14171), .B2(n8333), .A(n14078), .ZN(n14088) );
  OAI22_X1 U16009 ( .A1(n14665), .A2(n14080), .B1(n14079), .B2(n14673), .ZN(
        n14085) );
  XNOR2_X1 U16010 ( .A(n14082), .B(n14081), .ZN(n14175) );
  NOR2_X1 U16011 ( .A1(n14175), .A2(n14083), .ZN(n14084) );
  AOI211_X1 U16012 ( .C1(n14677), .C2(n14172), .A(n14085), .B(n14084), .ZN(
        n14086) );
  OAI21_X1 U16013 ( .B1(n14088), .B2(n14087), .A(n14086), .ZN(P1_U3275) );
  OAI211_X1 U16014 ( .C1(n14091), .C2(n14755), .A(n14090), .B(n14092), .ZN(
        n14182) );
  MUX2_X1 U16015 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14182), .S(n14776), .Z(
        P1_U3559) );
  OAI211_X1 U16016 ( .C1(n14094), .C2(n14755), .A(n14093), .B(n14092), .ZN(
        n14183) );
  MUX2_X1 U16017 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14183), .S(n14776), .Z(
        P1_U3558) );
  OAI211_X1 U16018 ( .C1(n12485), .C2(n14755), .A(n14098), .B(n14097), .ZN(
        n14099) );
  OAI211_X1 U16019 ( .C1(n14103), .C2(n14691), .A(n14102), .B(n14101), .ZN(
        n14184) );
  MUX2_X1 U16020 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14184), .S(n14776), .Z(
        P1_U3557) );
  NAND2_X1 U16021 ( .A1(n14104), .A2(n14723), .ZN(n14109) );
  NAND3_X1 U16022 ( .A1(n14106), .A2(n14759), .A3(n14105), .ZN(n14108) );
  NAND4_X1 U16023 ( .A1(n14110), .A2(n14109), .A3(n14108), .A4(n14107), .ZN(
        n14185) );
  MUX2_X1 U16024 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14185), .S(n14776), .Z(
        P1_U3556) );
  AOI21_X1 U16025 ( .B1(n14112), .B2(n14723), .A(n14111), .ZN(n14113) );
  OAI211_X1 U16026 ( .C1(n14691), .C2(n14115), .A(n14114), .B(n14113), .ZN(
        n14186) );
  MUX2_X1 U16027 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14186), .S(n14776), .Z(
        P1_U3555) );
  INV_X1 U16028 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n14122) );
  OAI21_X1 U16029 ( .B1(n14117), .B2(n14755), .A(n14116), .ZN(n14118) );
  AOI21_X1 U16030 ( .B1(n14119), .B2(n14759), .A(n14118), .ZN(n14120) );
  AND2_X1 U16031 ( .A1(n14121), .A2(n14120), .ZN(n14187) );
  MUX2_X1 U16032 ( .A(n14122), .B(n14187), .S(n14776), .Z(n14123) );
  INV_X1 U16033 ( .A(n14123), .ZN(P1_U3554) );
  AOI21_X1 U16034 ( .B1(n14125), .B2(n14723), .A(n14124), .ZN(n14130) );
  NAND3_X1 U16035 ( .A1(n14127), .A2(n14126), .A3(n14759), .ZN(n14129) );
  NAND4_X1 U16036 ( .A1(n14131), .A2(n14130), .A3(n14129), .A4(n14128), .ZN(
        n14190) );
  MUX2_X1 U16037 ( .A(n14190), .B(P1_REG1_REG_25__SCAN_IN), .S(n14773), .Z(
        P1_U3553) );
  AOI21_X1 U16038 ( .B1(n14133), .B2(n14723), .A(n14132), .ZN(n14134) );
  OAI211_X1 U16039 ( .C1(n14691), .C2(n14136), .A(n14135), .B(n14134), .ZN(
        n14191) );
  MUX2_X1 U16040 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14191), .S(n14776), .Z(
        P1_U3552) );
  AOI21_X1 U16041 ( .B1(n14138), .B2(n14723), .A(n14137), .ZN(n14139) );
  OAI211_X1 U16042 ( .C1(n14691), .C2(n14141), .A(n14140), .B(n14139), .ZN(
        n14192) );
  MUX2_X1 U16043 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14192), .S(n14776), .Z(
        P1_U3551) );
  INV_X1 U16044 ( .A(n14142), .ZN(n14143) );
  OAI211_X1 U16045 ( .C1(n14755), .C2(n8295), .A(n14144), .B(n14143), .ZN(
        n14145) );
  AOI21_X1 U16046 ( .B1(n14146), .B2(n14618), .A(n14145), .ZN(n14147) );
  OAI21_X1 U16047 ( .B1(n14691), .B2(n14148), .A(n14147), .ZN(n14193) );
  MUX2_X1 U16048 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14193), .S(n14776), .Z(
        P1_U3550) );
  AOI211_X1 U16049 ( .C1(n14151), .C2(n14723), .A(n14150), .B(n14149), .ZN(
        n14153) );
  OAI211_X1 U16050 ( .C1(n14154), .C2(n14691), .A(n14153), .B(n14152), .ZN(
        n14194) );
  MUX2_X1 U16051 ( .A(n14194), .B(P1_REG1_REG_21__SCAN_IN), .S(n14773), .Z(
        P1_U3549) );
  NAND3_X1 U16052 ( .A1(n14156), .A2(n14618), .A3(n14155), .ZN(n14165) );
  INV_X1 U16053 ( .A(n14157), .ZN(n14158) );
  AOI21_X1 U16054 ( .B1(n14159), .B2(n14723), .A(n14158), .ZN(n14164) );
  NAND3_X1 U16055 ( .A1(n6480), .A2(n14160), .A3(n14759), .ZN(n14163) );
  NAND4_X1 U16056 ( .A1(n14165), .A2(n14164), .A3(n14163), .A4(n14162), .ZN(
        n14195) );
  MUX2_X1 U16057 ( .A(n14195), .B(P1_REG1_REG_20__SCAN_IN), .S(n14773), .Z(
        P1_U3548) );
  OAI21_X1 U16058 ( .B1(n10006), .B2(n14755), .A(n14166), .ZN(n14167) );
  AOI21_X1 U16059 ( .B1(n14168), .B2(n14759), .A(n14167), .ZN(n14169) );
  OAI21_X1 U16060 ( .B1(n14170), .B2(n14690), .A(n14169), .ZN(n14196) );
  MUX2_X1 U16061 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14196), .S(n14776), .Z(
        P1_U3547) );
  AOI21_X1 U16062 ( .B1(n14172), .B2(n14723), .A(n14171), .ZN(n14173) );
  OAI211_X1 U16063 ( .C1(n14691), .C2(n14175), .A(n14174), .B(n14173), .ZN(
        n14197) );
  MUX2_X1 U16064 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14197), .S(n14776), .Z(
        P1_U3546) );
  NAND2_X1 U16065 ( .A1(n14176), .A2(n14759), .ZN(n14178) );
  OAI211_X1 U16066 ( .C1(n14179), .C2(n14755), .A(n14178), .B(n14177), .ZN(
        n14180) );
  MUX2_X1 U16067 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14198), .S(n14776), .Z(
        P1_U3545) );
  MUX2_X1 U16068 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14182), .S(n14761), .Z(
        P1_U3527) );
  MUX2_X1 U16069 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14183), .S(n14761), .Z(
        P1_U3526) );
  MUX2_X1 U16070 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14184), .S(n14761), .Z(
        P1_U3525) );
  MUX2_X1 U16071 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14185), .S(n14761), .Z(
        P1_U3524) );
  MUX2_X1 U16072 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14186), .S(n14761), .Z(
        P1_U3523) );
  MUX2_X1 U16073 ( .A(n14188), .B(n14187), .S(n14761), .Z(n14189) );
  INV_X1 U16074 ( .A(n14189), .ZN(P1_U3522) );
  MUX2_X1 U16075 ( .A(n14190), .B(P1_REG0_REG_25__SCAN_IN), .S(n14760), .Z(
        P1_U3521) );
  MUX2_X1 U16076 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14191), .S(n14761), .Z(
        P1_U3520) );
  MUX2_X1 U16077 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14192), .S(n14761), .Z(
        P1_U3519) );
  MUX2_X1 U16078 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14193), .S(n14761), .Z(
        P1_U3518) );
  MUX2_X1 U16079 ( .A(n14194), .B(P1_REG0_REG_21__SCAN_IN), .S(n14760), .Z(
        P1_U3517) );
  MUX2_X1 U16080 ( .A(n14195), .B(P1_REG0_REG_20__SCAN_IN), .S(n14760), .Z(
        P1_U3516) );
  MUX2_X1 U16081 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14196), .S(n14761), .Z(
        P1_U3515) );
  MUX2_X1 U16082 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14197), .S(n14761), .Z(
        P1_U3513) );
  MUX2_X1 U16083 ( .A(n14198), .B(P1_REG0_REG_17__SCAN_IN), .S(n14760), .Z(
        P1_U3510) );
  NOR4_X1 U16084 ( .A1(n14200), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), 
        .A4(n14199), .ZN(n14201) );
  AOI21_X1 U16085 ( .B1(n14202), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14201), 
        .ZN(n14203) );
  OAI21_X1 U16086 ( .B1(n14204), .B2(n14208), .A(n14203), .ZN(P1_U3324) );
  OAI222_X1 U16087 ( .A1(n12044), .A2(n14209), .B1(n14208), .B2(n14207), .C1(
        n14206), .C2(P1_U3086), .ZN(P1_U3328) );
  INV_X1 U16088 ( .A(n14210), .ZN(n14212) );
  OAI222_X1 U16089 ( .A1(n14214), .A2(n14213), .B1(P1_U3086), .B2(n14212), 
        .C1(n14211), .C2(n12044), .ZN(P1_U3329) );
  MUX2_X1 U16090 ( .A(n14216), .B(n14215), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  MUX2_X1 U16091 ( .A(n14217), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16092 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n14255) );
  XNOR2_X1 U16093 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n14309) );
  INV_X1 U16094 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14253) );
  INV_X1 U16095 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14251) );
  XOR2_X1 U16096 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .Z(n14307) );
  INV_X1 U16097 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14218) );
  XOR2_X1 U16098 ( .A(n14246), .B(n14218), .Z(n14259) );
  INV_X1 U16099 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14244) );
  XNOR2_X1 U16100 ( .A(n14240), .B(P3_ADDR_REG_9__SCAN_IN), .ZN(n14263) );
  XNOR2_X1 U16101 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n14291) );
  NAND2_X1 U16102 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n14221), .ZN(n14223) );
  NAND2_X1 U16103 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n14224), .ZN(n14227) );
  INV_X1 U16104 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n14225) );
  NAND2_X1 U16105 ( .A1(n14265), .A2(n14225), .ZN(n14226) );
  NAND2_X1 U16106 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n14228), .ZN(n14231) );
  INV_X1 U16107 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n15028) );
  INV_X1 U16108 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14229) );
  NAND2_X1 U16109 ( .A1(n14264), .A2(n14229), .ZN(n14230) );
  INV_X1 U16110 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n15044) );
  NAND2_X1 U16111 ( .A1(n14234), .A2(n15044), .ZN(n14236) );
  XNOR2_X1 U16112 ( .A(n14234), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n14287) );
  NAND2_X1 U16113 ( .A1(n14287), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n14235) );
  NAND2_X1 U16114 ( .A1(n14236), .A2(n14235), .ZN(n14292) );
  NAND2_X1 U16115 ( .A1(n14291), .A2(n14292), .ZN(n14237) );
  NAND2_X1 U16116 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n14260), .ZN(n14242) );
  NOR2_X1 U16117 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n14260), .ZN(n14241) );
  XNOR2_X1 U16118 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n14299) );
  NAND2_X1 U16119 ( .A1(n14300), .A2(n14299), .ZN(n14243) );
  INV_X1 U16120 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n14247) );
  NOR2_X1 U16121 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n14247), .ZN(n14249) );
  INV_X1 U16122 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14248) );
  NOR2_X1 U16123 ( .A1(n14307), .A2(n14306), .ZN(n14250) );
  AOI21_X1 U16124 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n14251), .A(n14250), 
        .ZN(n14257) );
  OR2_X1 U16125 ( .A1(n14253), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n14252) );
  AOI22_X1 U16126 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14253), .B1(n14257), 
        .B2(n14252), .ZN(n14308) );
  NAND2_X1 U16127 ( .A1(n14309), .A2(n14308), .ZN(n14254) );
  OAI21_X1 U16128 ( .B1(P3_ADDR_REG_16__SCAN_IN), .B2(n14255), .A(n14254), 
        .ZN(n14311) );
  XNOR2_X1 U16129 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14311), .ZN(n14312) );
  XNOR2_X1 U16130 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14312), .ZN(n14344) );
  XOR2_X1 U16131 ( .A(P3_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .Z(n14256) );
  XNOR2_X1 U16132 ( .A(n14257), .B(n14256), .ZN(n14554) );
  XOR2_X1 U16133 ( .A(n14259), .B(n14258), .Z(n14542) );
  XNOR2_X1 U16134 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(n14260), .ZN(n14261) );
  XNOR2_X1 U16135 ( .A(n14261), .B(P3_ADDR_REG_10__SCAN_IN), .ZN(n14332) );
  XOR2_X1 U16136 ( .A(n14263), .B(n14262), .Z(n14296) );
  XNOR2_X1 U16137 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n14264), .ZN(n14280) );
  XNOR2_X1 U16138 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n14265), .ZN(n14267) );
  INV_X1 U16139 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n14266) );
  NAND2_X1 U16140 ( .A1(n14267), .A2(n14266), .ZN(n14279) );
  XNOR2_X1 U16141 ( .A(P2_ADDR_REG_4__SCAN_IN), .B(n14267), .ZN(n15396) );
  XNOR2_X1 U16142 ( .A(n14268), .B(P1_ADDR_REG_3__SCAN_IN), .ZN(n15405) );
  XOR2_X1 U16143 ( .A(n14270), .B(n14269), .Z(n14320) );
  NOR2_X1 U16144 ( .A1(n14275), .A2(n10313), .ZN(n14276) );
  OAI21_X1 U16145 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n14274), .A(n14273), .ZN(
        n15400) );
  NAND2_X1 U16146 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15400), .ZN(n15410) );
  NOR2_X1 U16147 ( .A1(n15410), .A2(n15409), .ZN(n15408) );
  NOR2_X1 U16148 ( .A1(n14320), .A2(n14319), .ZN(n14277) );
  NAND2_X1 U16149 ( .A1(n14320), .A2(n14319), .ZN(n14318) );
  NOR2_X1 U16150 ( .A1(n15405), .A2(n15406), .ZN(n14278) );
  NAND2_X1 U16151 ( .A1(n15405), .A2(n15406), .ZN(n15404) );
  NAND2_X1 U16152 ( .A1(n14280), .A2(n14281), .ZN(n14282) );
  INV_X1 U16153 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15398) );
  NAND2_X1 U16154 ( .A1(n15399), .A2(n15398), .ZN(n15397) );
  NOR2_X1 U16155 ( .A1(n14283), .A2(n13272), .ZN(n14286) );
  XNOR2_X1 U16156 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n14285) );
  XOR2_X1 U16157 ( .A(n14285), .B(n14284), .Z(n14323) );
  NOR2_X1 U16158 ( .A1(n14288), .A2(n14289), .ZN(n14290) );
  XNOR2_X1 U16159 ( .A(n14287), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n15403) );
  NOR2_X1 U16160 ( .A1(n15403), .A2(n15402), .ZN(n15401) );
  XNOR2_X1 U16161 ( .A(n14292), .B(n14291), .ZN(n14294) );
  NAND2_X1 U16162 ( .A1(n14293), .A2(n14294), .ZN(n14295) );
  INV_X1 U16163 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14326) );
  NOR2_X1 U16164 ( .A1(n14296), .A2(n14297), .ZN(n14298) );
  XNOR2_X1 U16165 ( .A(n14297), .B(n14296), .ZN(n14329) );
  INV_X1 U16166 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14826) );
  NOR2_X1 U16167 ( .A1(n14329), .A2(n14826), .ZN(n14328) );
  XOR2_X1 U16168 ( .A(n14300), .B(n14299), .Z(n14302) );
  INV_X1 U16169 ( .A(n14538), .ZN(n14539) );
  INV_X1 U16170 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14831) );
  NAND2_X1 U16171 ( .A1(n14831), .A2(n14540), .ZN(n14537) );
  XNOR2_X1 U16172 ( .A(P1_ADDR_REG_13__SCAN_IN), .B(P3_ADDR_REG_13__SCAN_IN), 
        .ZN(n14304) );
  XNOR2_X1 U16173 ( .A(n14304), .B(n14303), .ZN(n14546) );
  NAND2_X1 U16174 ( .A1(n14547), .A2(n14546), .ZN(n14305) );
  XNOR2_X1 U16175 ( .A(n14307), .B(n14306), .ZN(n14551) );
  XNOR2_X1 U16176 ( .A(n14309), .B(n14308), .ZN(n14558) );
  NOR2_X1 U16177 ( .A1(n14559), .A2(n14558), .ZN(n14557) );
  NAND2_X1 U16178 ( .A1(n14559), .A2(n14558), .ZN(n14310) );
  NOR2_X1 U16179 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14311), .ZN(n14315) );
  INV_X1 U16180 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14313) );
  NOR2_X1 U16181 ( .A1(n14313), .A2(n14312), .ZN(n14314) );
  NOR2_X1 U16182 ( .A1(n14315), .A2(n14314), .ZN(n15385) );
  INV_X1 U16183 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n15387) );
  XNOR2_X1 U16184 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(n15387), .ZN(n15384) );
  XOR2_X1 U16185 ( .A(n15385), .B(n15384), .Z(n15381) );
  NAND2_X1 U16186 ( .A1(n15381), .A2(n15380), .ZN(n15382) );
  OAI21_X1 U16187 ( .B1(n15380), .B2(n15381), .A(n15382), .ZN(n14316) );
  XNOR2_X1 U16188 ( .A(n14316), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16189 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14317) );
  OAI21_X1 U16190 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14317), 
        .ZN(U28) );
  INV_X1 U16191 ( .A(P3_RD_REG_SCAN_IN), .ZN(n15296) );
  OAI221_X1 U16192 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(n7526), .C2(n7527), .A(n15296), .ZN(U29) );
  OAI21_X1 U16193 ( .B1(n14320), .B2(n14319), .A(n14318), .ZN(n14321) );
  XNOR2_X1 U16194 ( .A(n14321), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  AOI21_X1 U16195 ( .B1(n14324), .B2(n14323), .A(n14322), .ZN(SUB_1596_U57) );
  OAI21_X1 U16196 ( .B1(n14327), .B2(n14326), .A(n14325), .ZN(SUB_1596_U55) );
  AOI21_X1 U16197 ( .B1(n14329), .B2(n14826), .A(n14328), .ZN(SUB_1596_U54) );
  AOI21_X1 U16198 ( .B1(n14332), .B2(n14331), .A(n14330), .ZN(n14333) );
  XOR2_X1 U16199 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n14333), .Z(SUB_1596_U70)
         );
  INV_X1 U16200 ( .A(n14334), .ZN(n14340) );
  NOR2_X1 U16201 ( .A1(n14334), .A2(n14743), .ZN(n14339) );
  OAI211_X1 U16202 ( .C1(n14337), .C2(n14755), .A(n14336), .B(n14335), .ZN(
        n14338) );
  AOI211_X1 U16203 ( .C1(n14340), .C2(n14750), .A(n14339), .B(n14338), .ZN(
        n14342) );
  INV_X1 U16204 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14341) );
  AOI22_X1 U16205 ( .A1(n14761), .A2(n14342), .B1(n14341), .B2(n14760), .ZN(
        P1_U3495) );
  AOI22_X1 U16206 ( .A1(n14776), .A2(n14342), .B1(n10540), .B2(n14773), .ZN(
        P1_U3540) );
  OAI21_X1 U16207 ( .B1(n14345), .B2(n14344), .A(n14343), .ZN(n14346) );
  XNOR2_X1 U16208 ( .A(n14346), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(SUB_1596_U63)
         );
  AOI22_X1 U16209 ( .A1(n15080), .A2(n14347), .B1(n15068), .B2(
        P3_ADDR_REG_16__SCAN_IN), .ZN(n14364) );
  MUX2_X1 U16210 ( .A(n14350), .B(n14349), .S(n14348), .Z(n14352) );
  NOR2_X1 U16211 ( .A1(n14352), .A2(n14351), .ZN(n14354) );
  XOR2_X1 U16212 ( .A(n14354), .B(n14353), .Z(n14358) );
  XNOR2_X1 U16213 ( .A(n14356), .B(n14355), .ZN(n14357) );
  AOI22_X1 U16214 ( .A1(n14358), .A2(n15078), .B1(n15069), .B2(n14357), .ZN(
        n14363) );
  NAND2_X1 U16215 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(P3_U3151), .ZN(n14362)
         );
  OAI221_X1 U16216 ( .B1(n14360), .B2(n6617), .C1(n14360), .C2(n14359), .A(
        n15082), .ZN(n14361) );
  NAND4_X1 U16217 ( .A1(n14364), .A2(n14363), .A3(n14362), .A4(n14361), .ZN(
        P3_U3198) );
  AOI22_X1 U16218 ( .A1(n15080), .A2(n14365), .B1(n15068), .B2(
        P3_ADDR_REG_17__SCAN_IN), .ZN(n14379) );
  OAI21_X1 U16219 ( .B1(P3_REG1_REG_17__SCAN_IN), .B2(n14367), .A(n14366), 
        .ZN(n14373) );
  OAI211_X1 U16220 ( .C1(n14370), .C2(n14369), .A(n14368), .B(n15078), .ZN(
        n14371) );
  INV_X1 U16221 ( .A(n14371), .ZN(n14372) );
  AOI21_X1 U16222 ( .B1(n15069), .B2(n14373), .A(n14372), .ZN(n14378) );
  NAND2_X1 U16223 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(P3_U3151), .ZN(n14377)
         );
  OAI221_X1 U16224 ( .B1(n14375), .B2(n8738), .C1(n14375), .C2(n14374), .A(
        n15082), .ZN(n14376) );
  NAND4_X1 U16225 ( .A1(n14379), .A2(n14378), .A3(n14377), .A4(n14376), .ZN(
        P3_U3199) );
  AOI22_X1 U16226 ( .A1(n15080), .A2(n14380), .B1(n15068), .B2(
        P3_ADDR_REG_18__SCAN_IN), .ZN(n14394) );
  AOI21_X1 U16227 ( .B1(n14383), .B2(n14382), .A(n14381), .ZN(n14384) );
  INV_X1 U16228 ( .A(n14384), .ZN(n14389) );
  OAI21_X1 U16229 ( .B1(n14387), .B2(n14386), .A(n14385), .ZN(n14388) );
  AOI22_X1 U16230 ( .A1(n14389), .A2(n15078), .B1(n15069), .B2(n14388), .ZN(
        n14393) );
  NAND2_X1 U16231 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(P3_U3151), .ZN(n14392)
         );
  INV_X1 U16232 ( .A(n14395), .ZN(n14398) );
  OAI21_X1 U16233 ( .B1(n14398), .B2(n14397), .A(n14396), .ZN(n14404) );
  INV_X1 U16234 ( .A(n14399), .ZN(n14401) );
  AOI222_X1 U16235 ( .A1(n14404), .A2(n15117), .B1(n14403), .B2(n14402), .C1(
        n14401), .C2(n14400), .ZN(n14405) );
  OAI21_X1 U16236 ( .B1(n15117), .B2(n11395), .A(n14405), .ZN(P3_U3222) );
  AND2_X1 U16237 ( .A1(n14406), .A2(n14415), .ZN(n14409) );
  NOR2_X1 U16238 ( .A1(n14407), .A2(n15168), .ZN(n14408) );
  NOR3_X1 U16239 ( .A1(n14410), .A2(n14409), .A3(n14408), .ZN(n14417) );
  AOI22_X1 U16240 ( .A1(n15183), .A2(n14417), .B1(n8671), .B2(n9886), .ZN(
        P3_U3472) );
  NOR2_X1 U16241 ( .A1(n14411), .A2(n15168), .ZN(n14413) );
  AOI211_X1 U16242 ( .C1(n14415), .C2(n14414), .A(n14413), .B(n14412), .ZN(
        n14419) );
  AOI22_X1 U16243 ( .A1(n15183), .A2(n14419), .B1(n11559), .B2(n9886), .ZN(
        P3_U3471) );
  INV_X1 U16244 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14416) );
  AOI22_X1 U16245 ( .A1(n15175), .A2(n14417), .B1(n14416), .B2(n15173), .ZN(
        P3_U3429) );
  INV_X1 U16246 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14418) );
  AOI22_X1 U16247 ( .A1(n15175), .A2(n14419), .B1(n14418), .B2(n15173), .ZN(
        P3_U3426) );
  OAI22_X1 U16248 ( .A1(n14423), .A2(n14422), .B1(n14421), .B2(n14420), .ZN(
        n14434) );
  NAND2_X1 U16249 ( .A1(n14424), .A2(n14425), .ZN(n14426) );
  NAND2_X1 U16250 ( .A1(n14427), .A2(n14426), .ZN(n14429) );
  AOI222_X1 U16251 ( .A1(n14787), .A2(n14443), .B1(n14434), .B2(n14430), .C1(
        n14429), .C2(n14428), .ZN(n14432) );
  OAI211_X1 U16252 ( .C1(n14789), .C2(n14436), .A(n14432), .B(n14431), .ZN(
        P2_U3187) );
  XOR2_X1 U16253 ( .A(n14438), .B(n14433), .Z(n14435) );
  AOI21_X1 U16254 ( .B1(n14435), .B2(n14886), .A(n14434), .ZN(n14451) );
  INV_X1 U16255 ( .A(n14436), .ZN(n14437) );
  AOI222_X1 U16256 ( .A1(n14443), .A2(n14890), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(n14903), .C1(n14437), .C2(n14905), .ZN(n14448) );
  NAND2_X1 U16257 ( .A1(n14439), .A2(n14438), .ZN(n14440) );
  AND2_X1 U16258 ( .A1(n14441), .A2(n14440), .ZN(n14454) );
  AOI21_X1 U16259 ( .B1(n14443), .B2(n14442), .A(n13489), .ZN(n14445) );
  NAND2_X1 U16260 ( .A1(n14445), .A2(n14444), .ZN(n14449) );
  NOR2_X1 U16261 ( .A1(n14449), .A2(n14898), .ZN(n14446) );
  AOI21_X1 U16262 ( .B1(n14454), .B2(n14900), .A(n14446), .ZN(n14447) );
  OAI211_X1 U16263 ( .C1(n14903), .C2(n14451), .A(n14448), .B(n14447), .ZN(
        P2_U3251) );
  OAI21_X1 U16264 ( .B1(n14450), .B2(n14958), .A(n14449), .ZN(n14453) );
  INV_X1 U16265 ( .A(n14451), .ZN(n14452) );
  AOI211_X1 U16266 ( .C1(n14454), .C2(n14961), .A(n14453), .B(n14452), .ZN(
        n14467) );
  AOI22_X1 U16267 ( .A1(n13616), .A2(n14467), .B1(n14455), .B2(n14969), .ZN(
        P2_U3513) );
  INV_X1 U16268 ( .A(n14456), .ZN(n14458) );
  OAI21_X1 U16269 ( .B1(n14458), .B2(n14958), .A(n14457), .ZN(n14459) );
  AOI211_X1 U16270 ( .C1(n14461), .C2(n14961), .A(n14460), .B(n14459), .ZN(
        n14469) );
  AOI22_X1 U16271 ( .A1(n13616), .A2(n14469), .B1(n9180), .B2(n14969), .ZN(
        P2_U3512) );
  OAI211_X1 U16272 ( .C1(n14464), .C2(n14958), .A(n14463), .B(n14462), .ZN(
        n14465) );
  AOI21_X1 U16273 ( .B1(n14466), .B2(n14961), .A(n14465), .ZN(n14471) );
  AOI22_X1 U16274 ( .A1(n13616), .A2(n14471), .B1(n9167), .B2(n14969), .ZN(
        P2_U3511) );
  AOI22_X1 U16275 ( .A1(n14964), .A2(n14467), .B1(n9194), .B2(n14962), .ZN(
        P2_U3472) );
  INV_X1 U16276 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n14468) );
  AOI22_X1 U16277 ( .A1(n14964), .A2(n14469), .B1(n14468), .B2(n14962), .ZN(
        P2_U3469) );
  INV_X1 U16278 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14470) );
  AOI22_X1 U16279 ( .A1(n14964), .A2(n14471), .B1(n14470), .B2(n14962), .ZN(
        P2_U3466) );
  XNOR2_X1 U16280 ( .A(n14473), .B(n14472), .ZN(n14509) );
  OAI211_X1 U16281 ( .C1(n14476), .C2(n14475), .A(n14474), .B(n14618), .ZN(
        n14479) );
  INV_X1 U16282 ( .A(n14477), .ZN(n14478) );
  NAND2_X1 U16283 ( .A1(n14479), .A2(n14478), .ZN(n14516) );
  AOI21_X1 U16284 ( .B1(n14480), .B2(n14509), .A(n14516), .ZN(n14494) );
  XNOR2_X1 U16285 ( .A(n14511), .B(n14481), .ZN(n14513) );
  INV_X1 U16286 ( .A(n14513), .ZN(n14492) );
  AND2_X1 U16287 ( .A1(n14483), .A2(n14482), .ZN(n14510) );
  OAI22_X1 U16288 ( .A1(n14665), .A2(n14485), .B1(n14484), .B2(n14673), .ZN(
        n14486) );
  AOI21_X1 U16289 ( .B1(n14510), .B2(n14665), .A(n14486), .ZN(n14487) );
  OAI21_X1 U16290 ( .B1(n14489), .B2(n14488), .A(n14487), .ZN(n14490) );
  AOI21_X1 U16291 ( .B1(n14492), .B2(n14491), .A(n14490), .ZN(n14493) );
  OAI21_X1 U16292 ( .B1(n14644), .B2(n14494), .A(n14493), .ZN(P1_U3279) );
  INV_X1 U16293 ( .A(n14495), .ZN(n14496) );
  OAI211_X1 U16294 ( .C1(n14498), .C2(n14755), .A(n14497), .B(n14496), .ZN(
        n14500) );
  AOI211_X1 U16295 ( .C1(n14501), .C2(n14759), .A(n14500), .B(n14499), .ZN(
        n14529) );
  AOI22_X1 U16296 ( .A1(n14776), .A2(n14529), .B1(n11291), .B2(n14773), .ZN(
        P1_U3544) );
  AOI21_X1 U16297 ( .B1(n14503), .B2(n14723), .A(n14502), .ZN(n14505) );
  OAI211_X1 U16298 ( .C1(n14506), .C2(n14691), .A(n14505), .B(n14504), .ZN(
        n14508) );
  NOR2_X1 U16299 ( .A1(n14508), .A2(n14507), .ZN(n14531) );
  AOI22_X1 U16300 ( .A1(n14776), .A2(n14531), .B1(n7907), .B2(n14773), .ZN(
        P1_U3543) );
  AND2_X1 U16301 ( .A1(n14509), .A2(n14759), .ZN(n14515) );
  AOI21_X1 U16302 ( .B1(n14511), .B2(n14723), .A(n14510), .ZN(n14512) );
  OAI21_X1 U16303 ( .B1(n14513), .B2(n14699), .A(n14512), .ZN(n14514) );
  NOR3_X1 U16304 ( .A1(n14516), .A2(n14515), .A3(n14514), .ZN(n14533) );
  AOI22_X1 U16305 ( .A1(n14776), .A2(n14533), .B1(n7860), .B2(n14773), .ZN(
        P1_U3542) );
  AOI21_X1 U16306 ( .B1(n14518), .B2(n14723), .A(n14517), .ZN(n14520) );
  OAI211_X1 U16307 ( .C1(n14521), .C2(n14690), .A(n14520), .B(n14519), .ZN(
        n14522) );
  AOI21_X1 U16308 ( .B1(n14523), .B2(n14759), .A(n14522), .ZN(n14535) );
  AOI22_X1 U16309 ( .A1(n14776), .A2(n14535), .B1(n10652), .B2(n14773), .ZN(
        P1_U3541) );
  OAI211_X1 U16310 ( .C1(n14526), .C2(n14755), .A(n14525), .B(n14524), .ZN(
        n14527) );
  AOI21_X1 U16311 ( .B1(n14528), .B2(n14759), .A(n14527), .ZN(n14536) );
  AOI22_X1 U16312 ( .A1(n14776), .A2(n14536), .B1(n7805), .B2(n14773), .ZN(
        P1_U3539) );
  AOI22_X1 U16313 ( .A1(n14761), .A2(n14529), .B1(n7929), .B2(n14760), .ZN(
        P1_U3507) );
  INV_X1 U16314 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n14530) );
  AOI22_X1 U16315 ( .A1(n14761), .A2(n14531), .B1(n14530), .B2(n14760), .ZN(
        P1_U3504) );
  INV_X1 U16316 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14532) );
  AOI22_X1 U16317 ( .A1(n14761), .A2(n14533), .B1(n14532), .B2(n14760), .ZN(
        P1_U3501) );
  INV_X1 U16318 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14534) );
  AOI22_X1 U16319 ( .A1(n14761), .A2(n14535), .B1(n14534), .B2(n14760), .ZN(
        P1_U3498) );
  AOI22_X1 U16320 ( .A1(n14761), .A2(n14536), .B1(n7809), .B2(n14760), .ZN(
        P1_U3492) );
  OAI222_X1 U16321 ( .A1(n14831), .A2(n14540), .B1(n14831), .B2(n14539), .C1(
        n14538), .C2(n14537), .ZN(SUB_1596_U69) );
  OAI21_X1 U16322 ( .B1(n14543), .B2(n14542), .A(n14541), .ZN(n14544) );
  XNOR2_X1 U16323 ( .A(n14544), .B(P2_ADDR_REG_12__SCAN_IN), .ZN(SUB_1596_U68)
         );
  AOI21_X1 U16324 ( .B1(n14547), .B2(n14546), .A(n14545), .ZN(n14548) );
  XOR2_X1 U16325 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n14548), .Z(SUB_1596_U67)
         );
  OAI21_X1 U16326 ( .B1(n14551), .B2(n14550), .A(n14549), .ZN(n14552) );
  XNOR2_X1 U16327 ( .A(n14552), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  OAI21_X1 U16328 ( .B1(n14555), .B2(n14554), .A(n14553), .ZN(n14556) );
  XNOR2_X1 U16329 ( .A(n14556), .B(P2_ADDR_REG_15__SCAN_IN), .ZN(SUB_1596_U65)
         );
  AOI21_X1 U16330 ( .B1(n14559), .B2(n14558), .A(n14557), .ZN(n14560) );
  XOR2_X1 U16331 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n14560), .Z(SUB_1596_U64)
         );
  OAI21_X1 U16332 ( .B1(n14562), .B2(P1_REG1_REG_0__SCAN_IN), .A(n14561), .ZN(
        n14563) );
  XOR2_X1 U16333 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14563), .Z(n14566) );
  AOI22_X1 U16334 ( .A1(n14587), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14564) );
  OAI21_X1 U16335 ( .B1(n14566), .B2(n14565), .A(n14564), .ZN(P1_U3243) );
  INV_X1 U16336 ( .A(n14567), .ZN(n14572) );
  NAND3_X1 U16337 ( .A1(n14570), .A2(n14569), .A3(n14568), .ZN(n14571) );
  NAND3_X1 U16338 ( .A1(n14606), .A2(n14572), .A3(n14571), .ZN(n14584) );
  AND2_X1 U16339 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n14573) );
  AOI21_X1 U16340 ( .B1(n14587), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n14573), .ZN(
        n14583) );
  NAND2_X1 U16341 ( .A1(n14591), .A2(n14574), .ZN(n14582) );
  MUX2_X1 U16342 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10136), .S(n14575), .Z(
        n14578) );
  NAND3_X1 U16343 ( .A1(n14578), .A2(n14577), .A3(n14576), .ZN(n14579) );
  NAND3_X1 U16344 ( .A1(n14603), .A2(n14580), .A3(n14579), .ZN(n14581) );
  AND4_X1 U16345 ( .A1(n14584), .A2(n14583), .A3(n14582), .A4(n14581), .ZN(
        n14586) );
  NAND2_X1 U16346 ( .A1(n14586), .A2(n14585), .ZN(P1_U3247) );
  NAND2_X1 U16347 ( .A1(n14587), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n14589) );
  NAND2_X1 U16348 ( .A1(n14589), .A2(n14588), .ZN(n14590) );
  AOI21_X1 U16349 ( .B1(n14592), .B2(n14591), .A(n14590), .ZN(n14601) );
  OAI211_X1 U16350 ( .C1(n14595), .C2(n14594), .A(n14593), .B(n14606), .ZN(
        n14600) );
  OAI211_X1 U16351 ( .C1(n14598), .C2(n14597), .A(n14596), .B(n14603), .ZN(
        n14599) );
  NAND3_X1 U16352 ( .A1(n14601), .A2(n14600), .A3(n14599), .ZN(P1_U3256) );
  OAI211_X1 U16353 ( .C1(n14604), .C2(P1_REG1_REG_18__SCAN_IN), .A(n14603), 
        .B(n14602), .ZN(n14609) );
  OAI211_X1 U16354 ( .C1(n14607), .C2(P1_REG2_REG_18__SCAN_IN), .A(n14606), 
        .B(n14605), .ZN(n14608) );
  OAI211_X1 U16355 ( .C1(n14611), .C2(n14610), .A(n14609), .B(n14608), .ZN(
        n14612) );
  INV_X1 U16356 ( .A(n14612), .ZN(n14614) );
  OAI211_X1 U16357 ( .C1(n15387), .C2(n14615), .A(n14614), .B(n14613), .ZN(
        P1_U3261) );
  AND2_X1 U16358 ( .A1(n14617), .A2(n14616), .ZN(n14620) );
  OAI211_X1 U16359 ( .C1(n14621), .C2(n14620), .A(n14619), .B(n14618), .ZN(
        n14623) );
  AND2_X1 U16360 ( .A1(n14623), .A2(n14622), .ZN(n14754) );
  INV_X1 U16361 ( .A(n14624), .ZN(n14625) );
  AOI222_X1 U16362 ( .A1(n14628), .A2(n14677), .B1(n14625), .B2(n14643), .C1(
        P1_REG2_REG_10__SCAN_IN), .C2(n14644), .ZN(n14635) );
  XNOR2_X1 U16363 ( .A(n14626), .B(n14627), .ZN(n14758) );
  XNOR2_X1 U16364 ( .A(n14629), .B(n14628), .ZN(n14632) );
  AOI22_X1 U16365 ( .A1(n14632), .A2(n14679), .B1(n14631), .B2(n14630), .ZN(
        n14753) );
  INV_X1 U16366 ( .A(n14753), .ZN(n14633) );
  AOI22_X1 U16367 ( .A1(n14758), .A2(n14662), .B1(n14683), .B2(n14633), .ZN(
        n14634) );
  OAI211_X1 U16368 ( .C1(n14644), .C2(n14754), .A(n14635), .B(n14634), .ZN(
        P1_U3283) );
  XNOR2_X1 U16369 ( .A(n6481), .B(n14637), .ZN(n14741) );
  XNOR2_X1 U16370 ( .A(n14638), .B(n14637), .ZN(n14640) );
  OAI21_X1 U16371 ( .B1(n14640), .B2(n14690), .A(n14639), .ZN(n14641) );
  AOI21_X1 U16372 ( .B1(n14750), .B2(n14741), .A(n14641), .ZN(n14738) );
  AOI222_X1 U16373 ( .A1(n14647), .A2(n14677), .B1(P1_REG2_REG_7__SCAN_IN), 
        .B2(n14644), .C1(n14643), .C2(n14642), .ZN(n14650) );
  INV_X1 U16374 ( .A(n14645), .ZN(n14684) );
  OAI211_X1 U16375 ( .C1(n6880), .C2(n6879), .A(n14679), .B(n6517), .ZN(n14737) );
  INV_X1 U16376 ( .A(n14737), .ZN(n14648) );
  AOI22_X1 U16377 ( .A1(n14741), .A2(n14684), .B1(n14683), .B2(n14648), .ZN(
        n14649) );
  OAI211_X1 U16378 ( .C1(n14644), .C2(n14738), .A(n14650), .B(n14649), .ZN(
        P1_U3286) );
  XNOR2_X1 U16379 ( .A(n14651), .B(n14659), .ZN(n14654) );
  INV_X1 U16380 ( .A(n14652), .ZN(n14653) );
  OAI21_X1 U16381 ( .B1(n14654), .B2(n14690), .A(n14653), .ZN(n14719) );
  OAI22_X1 U16382 ( .A1(n14673), .A2(n14656), .B1(n14718), .B2(n14655), .ZN(
        n14657) );
  NOR2_X1 U16383 ( .A1(n14719), .A2(n14657), .ZN(n14666) );
  XNOR2_X1 U16384 ( .A(n14658), .B(n14659), .ZN(n14721) );
  OAI211_X1 U16385 ( .C1(n14678), .C2(n14718), .A(n14679), .B(n14660), .ZN(
        n14717) );
  INV_X1 U16386 ( .A(n14717), .ZN(n14661) );
  AOI22_X1 U16387 ( .A1(n14721), .A2(n14662), .B1(n14683), .B2(n14661), .ZN(
        n14663) );
  OAI221_X1 U16388 ( .B1(n14644), .B2(n14666), .C1(n14665), .C2(n14664), .A(
        n14663), .ZN(P1_U3289) );
  XNOR2_X1 U16389 ( .A(n14667), .B(n14669), .ZN(n14715) );
  XNOR2_X1 U16390 ( .A(n14668), .B(n14669), .ZN(n14671) );
  OAI21_X1 U16391 ( .B1(n14671), .B2(n14690), .A(n14670), .ZN(n14672) );
  AOI21_X1 U16392 ( .B1(n14715), .B2(n14750), .A(n14672), .ZN(n14712) );
  OAI22_X1 U16393 ( .A1(n14665), .A2(n14674), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14673), .ZN(n14675) );
  AOI21_X1 U16394 ( .B1(n14677), .B2(n14676), .A(n14675), .ZN(n14686) );
  INV_X1 U16395 ( .A(n14678), .ZN(n14680) );
  OAI211_X1 U16396 ( .C1(n14711), .C2(n14681), .A(n14680), .B(n14679), .ZN(
        n14710) );
  INV_X1 U16397 ( .A(n14710), .ZN(n14682) );
  AOI22_X1 U16398 ( .A1(n14715), .A2(n14684), .B1(n14683), .B2(n14682), .ZN(
        n14685) );
  OAI211_X1 U16399 ( .C1(n14644), .C2(n14712), .A(n14686), .B(n14685), .ZN(
        P1_U3290) );
  AND2_X1 U16400 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14687), .ZN(P1_U3294) );
  AND2_X1 U16401 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14687), .ZN(P1_U3295) );
  AND2_X1 U16402 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14687), .ZN(P1_U3296) );
  AND2_X1 U16403 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14687), .ZN(P1_U3297) );
  AND2_X1 U16404 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14687), .ZN(P1_U3298) );
  AND2_X1 U16405 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14687), .ZN(P1_U3299) );
  AND2_X1 U16406 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14687), .ZN(P1_U3300) );
  AND2_X1 U16407 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14687), .ZN(P1_U3301) );
  AND2_X1 U16408 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14687), .ZN(P1_U3302) );
  AND2_X1 U16409 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14687), .ZN(P1_U3303) );
  AND2_X1 U16410 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14687), .ZN(P1_U3304) );
  AND2_X1 U16411 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14687), .ZN(P1_U3305) );
  AND2_X1 U16412 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14687), .ZN(P1_U3306) );
  AND2_X1 U16413 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14687), .ZN(P1_U3307) );
  AND2_X1 U16414 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14687), .ZN(P1_U3308) );
  AND2_X1 U16415 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14687), .ZN(P1_U3309) );
  AND2_X1 U16416 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14687), .ZN(P1_U3310) );
  AND2_X1 U16417 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14687), .ZN(P1_U3311) );
  AND2_X1 U16418 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14687), .ZN(P1_U3312) );
  AND2_X1 U16419 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14687), .ZN(P1_U3313) );
  AND2_X1 U16420 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14687), .ZN(P1_U3314) );
  AND2_X1 U16421 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14687), .ZN(P1_U3315) );
  AND2_X1 U16422 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14687), .ZN(P1_U3316) );
  AND2_X1 U16423 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14687), .ZN(P1_U3317) );
  AND2_X1 U16424 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14687), .ZN(P1_U3318) );
  AND2_X1 U16425 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14687), .ZN(P1_U3319) );
  AND2_X1 U16426 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14687), .ZN(P1_U3320) );
  AND2_X1 U16427 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14687), .ZN(P1_U3321) );
  AND2_X1 U16428 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14687), .ZN(P1_U3322) );
  AND2_X1 U16429 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14687), .ZN(P1_U3323) );
  INV_X1 U16430 ( .A(n14688), .ZN(n14695) );
  AOI21_X1 U16431 ( .B1(n14691), .B2(n14690), .A(n14689), .ZN(n14692) );
  AOI211_X1 U16432 ( .C1(n14695), .C2(n14694), .A(n14693), .B(n14692), .ZN(
        n14763) );
  INV_X1 U16433 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n14696) );
  AOI22_X1 U16434 ( .A1(n14761), .A2(n14763), .B1(n14696), .B2(n14760), .ZN(
        P1_U3459) );
  INV_X1 U16435 ( .A(n14743), .ZN(n14742) );
  INV_X1 U16436 ( .A(n14697), .ZN(n14703) );
  OAI22_X1 U16437 ( .A1(n14700), .A2(n14699), .B1(n14755), .B2(n14698), .ZN(
        n14702) );
  AOI211_X1 U16438 ( .C1(n14742), .C2(n14703), .A(n14702), .B(n14701), .ZN(
        n14764) );
  AOI22_X1 U16439 ( .A1(n14761), .A2(n14764), .B1(n7553), .B2(n14760), .ZN(
        P1_U3462) );
  AOI21_X1 U16440 ( .B1(n14730), .B2(n14743), .A(n14704), .ZN(n14709) );
  NOR2_X1 U16441 ( .A1(n14755), .A2(n14705), .ZN(n14708) );
  NOR4_X1 U16442 ( .A1(n14709), .A2(n14708), .A3(n14707), .A4(n14706), .ZN(
        n14765) );
  AOI22_X1 U16443 ( .A1(n14761), .A2(n14765), .B1(n7577), .B2(n14760), .ZN(
        P1_U3465) );
  OAI21_X1 U16444 ( .B1(n14711), .B2(n14755), .A(n14710), .ZN(n14714) );
  INV_X1 U16445 ( .A(n14712), .ZN(n14713) );
  AOI211_X1 U16446 ( .C1(n14742), .C2(n14715), .A(n14714), .B(n14713), .ZN(
        n14766) );
  INV_X1 U16447 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n14716) );
  AOI22_X1 U16448 ( .A1(n14761), .A2(n14766), .B1(n14716), .B2(n14760), .ZN(
        P1_U3468) );
  OAI21_X1 U16449 ( .B1(n14718), .B2(n14755), .A(n14717), .ZN(n14720) );
  AOI211_X1 U16450 ( .C1(n14721), .C2(n14759), .A(n14720), .B(n14719), .ZN(
        n14767) );
  AOI22_X1 U16451 ( .A1(n14761), .A2(n14767), .B1(n7625), .B2(n14760), .ZN(
        P1_U3471) );
  AOI21_X1 U16452 ( .B1(n14724), .B2(n14723), .A(n14722), .ZN(n14725) );
  OAI211_X1 U16453 ( .C1(n14743), .C2(n14727), .A(n14726), .B(n14725), .ZN(
        n14728) );
  INV_X1 U16454 ( .A(n14728), .ZN(n14769) );
  AOI22_X1 U16455 ( .A1(n14761), .A2(n14769), .B1(n7655), .B2(n14760), .ZN(
        P1_U3474) );
  AOI21_X1 U16456 ( .B1(n14730), .B2(n14743), .A(n14729), .ZN(n14735) );
  OAI21_X1 U16457 ( .B1(n14732), .B2(n14755), .A(n14731), .ZN(n14733) );
  NOR3_X1 U16458 ( .A1(n14735), .A2(n14734), .A3(n14733), .ZN(n14770) );
  INV_X1 U16459 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14736) );
  AOI22_X1 U16460 ( .A1(n14761), .A2(n14770), .B1(n14736), .B2(n14760), .ZN(
        P1_U3477) );
  OAI21_X1 U16461 ( .B1(n6879), .B2(n14755), .A(n14737), .ZN(n14740) );
  INV_X1 U16462 ( .A(n14738), .ZN(n14739) );
  AOI211_X1 U16463 ( .C1(n14742), .C2(n14741), .A(n14740), .B(n14739), .ZN(
        n14771) );
  AOI22_X1 U16464 ( .A1(n14761), .A2(n14771), .B1(n7708), .B2(n14760), .ZN(
        P1_U3480) );
  INV_X1 U16465 ( .A(n14744), .ZN(n14751) );
  NOR2_X1 U16466 ( .A1(n14744), .A2(n14743), .ZN(n14749) );
  OAI211_X1 U16467 ( .C1(n14747), .C2(n14755), .A(n14746), .B(n14745), .ZN(
        n14748) );
  AOI211_X1 U16468 ( .C1(n14751), .C2(n14750), .A(n14749), .B(n14748), .ZN(
        n14772) );
  INV_X1 U16469 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14752) );
  AOI22_X1 U16470 ( .A1(n14761), .A2(n14772), .B1(n14752), .B2(n14760), .ZN(
        P1_U3486) );
  OAI211_X1 U16471 ( .C1(n14756), .C2(n14755), .A(n14754), .B(n14753), .ZN(
        n14757) );
  AOI21_X1 U16472 ( .B1(n14759), .B2(n14758), .A(n14757), .ZN(n14775) );
  AOI22_X1 U16473 ( .A1(n14761), .A2(n14775), .B1(n7784), .B2(n14760), .ZN(
        P1_U3489) );
  AOI22_X1 U16474 ( .A1(n14776), .A2(n14763), .B1(n14762), .B2(n14773), .ZN(
        P1_U3528) );
  AOI22_X1 U16475 ( .A1(n14776), .A2(n14764), .B1(n10128), .B2(n14773), .ZN(
        P1_U3529) );
  AOI22_X1 U16476 ( .A1(n14776), .A2(n14765), .B1(n10132), .B2(n14773), .ZN(
        P1_U3530) );
  AOI22_X1 U16477 ( .A1(n14776), .A2(n14766), .B1(n10135), .B2(n14773), .ZN(
        P1_U3531) );
  AOI22_X1 U16478 ( .A1(n14776), .A2(n14767), .B1(n10136), .B2(n14773), .ZN(
        P1_U3532) );
  AOI22_X1 U16479 ( .A1(n14776), .A2(n14769), .B1(n14768), .B2(n14773), .ZN(
        P1_U3533) );
  AOI22_X1 U16480 ( .A1(n14776), .A2(n14770), .B1(n10141), .B2(n14773), .ZN(
        P1_U3534) );
  AOI22_X1 U16481 ( .A1(n14776), .A2(n14771), .B1(n10142), .B2(n14773), .ZN(
        P1_U3535) );
  AOI22_X1 U16482 ( .A1(n14776), .A2(n14772), .B1(n7755), .B2(n14773), .ZN(
        P1_U3537) );
  AOI22_X1 U16483 ( .A1(n14776), .A2(n14775), .B1(n14774), .B2(n14773), .ZN(
        P1_U3538) );
  NOR2_X1 U16484 ( .A1(n14871), .A2(P2_U3947), .ZN(P2_U3087) );
  INV_X1 U16485 ( .A(n14777), .ZN(n14778) );
  INV_X1 U16486 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n14904) );
  OAI22_X1 U16487 ( .A1(n14779), .A2(n14778), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14904), .ZN(n14786) );
  INV_X1 U16488 ( .A(n14780), .ZN(n14781) );
  AOI211_X1 U16489 ( .C1(n14784), .C2(n14783), .A(n14782), .B(n14781), .ZN(
        n14785) );
  AOI211_X1 U16490 ( .C1(n14906), .C2(n14787), .A(n14786), .B(n14785), .ZN(
        n14788) );
  OAI21_X1 U16491 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n14789), .A(n14788), .ZN(
        P2_U3190) );
  AOI21_X1 U16492 ( .B1(n14878), .B2(P2_REG1_REG_0__SCAN_IN), .A(n14790), .ZN(
        n14794) );
  AOI22_X1 U16493 ( .A1(n14871), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n14793) );
  OAI22_X1 U16494 ( .A1(n14856), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n14862), .ZN(n14791) );
  OAI21_X1 U16495 ( .B1(n14873), .B2(n14791), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n14792) );
  OAI211_X1 U16496 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n14794), .A(n14793), .B(
        n14792), .ZN(P2_U3214) );
  INV_X1 U16497 ( .A(n14795), .ZN(n14797) );
  OAI21_X1 U16498 ( .B1(n14797), .B2(n14796), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n14798) );
  OAI21_X1 U16499 ( .B1(P2_STATE_REG_SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n14798), .ZN(n14808) );
  OAI211_X1 U16500 ( .C1(n14801), .C2(n14800), .A(n14878), .B(n14799), .ZN(
        n14807) );
  OAI211_X1 U16501 ( .C1(n14804), .C2(n14803), .A(n14875), .B(n14802), .ZN(
        n14806) );
  NAND2_X1 U16502 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14871), .ZN(n14805) );
  NAND4_X1 U16503 ( .A1(n14808), .A2(n14807), .A3(n14806), .A4(n14805), .ZN(
        P2_U3218) );
  NAND2_X1 U16504 ( .A1(n14810), .A2(n14809), .ZN(n14811) );
  NAND2_X1 U16505 ( .A1(n14812), .A2(n14811), .ZN(n14813) );
  NAND2_X1 U16506 ( .A1(n14813), .A2(n14878), .ZN(n14820) );
  NAND2_X1 U16507 ( .A1(n14815), .A2(n14814), .ZN(n14816) );
  NAND2_X1 U16508 ( .A1(n14817), .A2(n14816), .ZN(n14818) );
  NAND2_X1 U16509 ( .A1(n14818), .A2(n14875), .ZN(n14819) );
  OAI211_X1 U16510 ( .C1(n14822), .C2(n14821), .A(n14820), .B(n14819), .ZN(
        n14823) );
  INV_X1 U16511 ( .A(n14823), .ZN(n14825) );
  OAI211_X1 U16512 ( .C1(n14826), .C2(n14832), .A(n14825), .B(n14824), .ZN(
        P2_U3223) );
  INV_X1 U16513 ( .A(n14827), .ZN(n14828) );
  AOI21_X1 U16514 ( .B1(n14830), .B2(n14829), .A(n14828), .ZN(n14841) );
  OAI22_X1 U16515 ( .A1(n14832), .A2(n14831), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9149), .ZN(n14833) );
  AOI21_X1 U16516 ( .B1(n14834), .B2(n14873), .A(n14833), .ZN(n14840) );
  AOI211_X1 U16517 ( .C1(n14837), .C2(n14836), .A(n14862), .B(n14835), .ZN(
        n14838) );
  INV_X1 U16518 ( .A(n14838), .ZN(n14839) );
  OAI211_X1 U16519 ( .C1(n14841), .C2(n14856), .A(n14840), .B(n14839), .ZN(
        P2_U3225) );
  NOR2_X1 U16520 ( .A1(n14843), .A2(n14842), .ZN(n14844) );
  NOR2_X1 U16521 ( .A1(n14845), .A2(n14844), .ZN(n14857) );
  NOR2_X1 U16522 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14846), .ZN(n14854) );
  OAI21_X1 U16523 ( .B1(n14849), .B2(n14848), .A(n14847), .ZN(n14851) );
  AOI22_X1 U16524 ( .A1(n14851), .A2(n14878), .B1(n14850), .B2(n14873), .ZN(
        n14852) );
  INV_X1 U16525 ( .A(n14852), .ZN(n14853) );
  AOI211_X1 U16526 ( .C1(P2_ADDR_REG_12__SCAN_IN), .C2(n14871), .A(n14854), 
        .B(n14853), .ZN(n14855) );
  OAI21_X1 U16527 ( .B1(n14857), .B2(n14856), .A(n14855), .ZN(P2_U3226) );
  AOI22_X1 U16528 ( .A1(n14871), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3088), .ZN(n14870) );
  OAI211_X1 U16529 ( .C1(n14860), .C2(n14859), .A(n14858), .B(n14875), .ZN(
        n14869) );
  AOI211_X1 U16530 ( .C1(n14864), .C2(n14863), .A(n14862), .B(n14861), .ZN(
        n14865) );
  INV_X1 U16531 ( .A(n14865), .ZN(n14868) );
  NAND2_X1 U16532 ( .A1(n14866), .A2(n14873), .ZN(n14867) );
  NAND4_X1 U16533 ( .A1(n14870), .A2(n14869), .A3(n14868), .A4(n14867), .ZN(
        P2_U3227) );
  AOI22_X1 U16534 ( .A1(n14871), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n14883) );
  NAND2_X1 U16535 ( .A1(n14873), .A2(n14872), .ZN(n14882) );
  OAI211_X1 U16536 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n14876), .A(n14875), 
        .B(n14874), .ZN(n14881) );
  OAI211_X1 U16537 ( .C1(n14879), .C2(P2_REG1_REG_15__SCAN_IN), .A(n14878), 
        .B(n14877), .ZN(n14880) );
  NAND4_X1 U16538 ( .A1(n14883), .A2(n14882), .A3(n14881), .A4(n14880), .ZN(
        P2_U3229) );
  XNOR2_X1 U16539 ( .A(n14884), .B(n14891), .ZN(n14887) );
  AOI21_X1 U16540 ( .B1(n14887), .B2(n14886), .A(n14885), .ZN(n14936) );
  INV_X1 U16541 ( .A(n14888), .ZN(n14889) );
  AOI222_X1 U16542 ( .A1(n14934), .A2(n14890), .B1(P2_REG2_REG_6__SCAN_IN), 
        .B2(n14903), .C1(n14889), .C2(n14905), .ZN(n14902) );
  NAND2_X1 U16543 ( .A1(n14892), .A2(n14891), .ZN(n14893) );
  AND2_X1 U16544 ( .A1(n14894), .A2(n14893), .ZN(n14939) );
  AOI21_X1 U16545 ( .B1(n14895), .B2(n14934), .A(n13489), .ZN(n14897) );
  NAND2_X1 U16546 ( .A1(n14897), .A2(n14896), .ZN(n14935) );
  NOR2_X1 U16547 ( .A1(n14935), .A2(n14898), .ZN(n14899) );
  AOI21_X1 U16548 ( .B1(n14939), .B2(n14900), .A(n14899), .ZN(n14901) );
  OAI211_X1 U16549 ( .C1(n14903), .C2(n14936), .A(n14902), .B(n14901), .ZN(
        P2_U3259) );
  INV_X1 U16550 ( .A(n9471), .ZN(n14910) );
  AOI22_X1 U16551 ( .A1(n14907), .A2(n14906), .B1(n14905), .B2(n14904), .ZN(
        n14908) );
  OAI211_X1 U16552 ( .C1(n14911), .C2(n14910), .A(n14909), .B(n14908), .ZN(
        n14917) );
  INV_X1 U16553 ( .A(n14912), .ZN(n14913) );
  AOI222_X1 U16554 ( .A1(n14917), .A2(n14919), .B1(n14916), .B2(n14915), .C1(
        n14914), .C2(n14913), .ZN(n14918) );
  OAI21_X1 U16555 ( .B1(n14919), .B2(n10290), .A(n14918), .ZN(P2_U3262) );
  AND2_X1 U16556 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14921), .ZN(P2_U3266) );
  AND2_X1 U16557 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14921), .ZN(P2_U3267) );
  AND2_X1 U16558 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14921), .ZN(P2_U3268) );
  AND2_X1 U16559 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14921), .ZN(P2_U3269) );
  AND2_X1 U16560 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14921), .ZN(P2_U3270) );
  AND2_X1 U16561 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14921), .ZN(P2_U3271) );
  AND2_X1 U16562 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14921), .ZN(P2_U3272) );
  AND2_X1 U16563 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14921), .ZN(P2_U3273) );
  AND2_X1 U16564 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14921), .ZN(P2_U3274) );
  AND2_X1 U16565 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14921), .ZN(P2_U3275) );
  AND2_X1 U16566 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14921), .ZN(P2_U3276) );
  AND2_X1 U16567 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14921), .ZN(P2_U3277) );
  AND2_X1 U16568 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14921), .ZN(P2_U3278) );
  AND2_X1 U16569 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14921), .ZN(P2_U3279) );
  AND2_X1 U16570 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14921), .ZN(P2_U3280) );
  AND2_X1 U16571 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14921), .ZN(P2_U3281) );
  AND2_X1 U16572 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14921), .ZN(P2_U3282) );
  AND2_X1 U16573 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14921), .ZN(P2_U3283) );
  AND2_X1 U16574 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14921), .ZN(P2_U3284) );
  AND2_X1 U16575 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14921), .ZN(P2_U3285) );
  AND2_X1 U16576 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14921), .ZN(P2_U3286) );
  AND2_X1 U16577 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14921), .ZN(P2_U3287) );
  AND2_X1 U16578 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14921), .ZN(P2_U3288) );
  AND2_X1 U16579 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14921), .ZN(P2_U3289) );
  AND2_X1 U16580 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14921), .ZN(P2_U3290) );
  AND2_X1 U16581 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14921), .ZN(P2_U3291) );
  AND2_X1 U16582 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14921), .ZN(P2_U3292) );
  AND2_X1 U16583 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14921), .ZN(P2_U3293) );
  AND2_X1 U16584 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14921), .ZN(P2_U3294) );
  AND2_X1 U16585 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14921), .ZN(P2_U3295) );
  OAI21_X1 U16586 ( .B1(n14927), .B2(n14923), .A(n14922), .ZN(P2_U3416) );
  AOI22_X1 U16587 ( .A1(n14927), .A2(n14926), .B1(n14925), .B2(n14924), .ZN(
        P2_U3417) );
  OAI211_X1 U16588 ( .C1(n14930), .C2(n14958), .A(n14929), .B(n14928), .ZN(
        n14931) );
  AOI21_X1 U16589 ( .B1(n14932), .B2(n14961), .A(n14931), .ZN(n14965) );
  INV_X1 U16590 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n14933) );
  AOI22_X1 U16591 ( .A1(n14964), .A2(n14965), .B1(n14933), .B2(n14962), .ZN(
        P2_U3445) );
  OAI21_X1 U16592 ( .B1(n6940), .B2(n14958), .A(n14935), .ZN(n14938) );
  INV_X1 U16593 ( .A(n14936), .ZN(n14937) );
  AOI211_X1 U16594 ( .C1(n14939), .C2(n14961), .A(n14938), .B(n14937), .ZN(
        n14966) );
  AOI22_X1 U16595 ( .A1(n14964), .A2(n14966), .B1(n9081), .B2(n14962), .ZN(
        P2_U3448) );
  OAI211_X1 U16596 ( .C1(n14942), .C2(n14958), .A(n14941), .B(n14940), .ZN(
        n14943) );
  AOI21_X1 U16597 ( .B1(n14944), .B2(n14961), .A(n14943), .ZN(n14967) );
  AOI22_X1 U16598 ( .A1(n14964), .A2(n14967), .B1(n9094), .B2(n14962), .ZN(
        P2_U3451) );
  AND2_X1 U16599 ( .A1(n14946), .A2(n14945), .ZN(n14947) );
  OR2_X1 U16600 ( .A1(n14948), .A2(n14947), .ZN(n14949) );
  AOI21_X1 U16601 ( .B1(n14951), .B2(n14950), .A(n14949), .ZN(n14952) );
  AND2_X1 U16602 ( .A1(n14953), .A2(n14952), .ZN(n14968) );
  INV_X1 U16603 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n14954) );
  AOI22_X1 U16604 ( .A1(n14964), .A2(n14968), .B1(n14954), .B2(n14962), .ZN(
        P2_U3454) );
  OAI211_X1 U16605 ( .C1(n6937), .C2(n14958), .A(n14957), .B(n14956), .ZN(
        n14959) );
  AOI21_X1 U16606 ( .B1(n14961), .B2(n14960), .A(n14959), .ZN(n14970) );
  INV_X1 U16607 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n14963) );
  AOI22_X1 U16608 ( .A1(n14964), .A2(n14970), .B1(n14963), .B2(n14962), .ZN(
        P2_U3463) );
  AOI22_X1 U16609 ( .A1(n13616), .A2(n14965), .B1(n10274), .B2(n14969), .ZN(
        P2_U3504) );
  AOI22_X1 U16610 ( .A1(n13616), .A2(n14966), .B1(n10277), .B2(n14969), .ZN(
        P2_U3505) );
  AOI22_X1 U16611 ( .A1(n13616), .A2(n14967), .B1(n10280), .B2(n14969), .ZN(
        P2_U3506) );
  AOI22_X1 U16612 ( .A1(n13616), .A2(n14968), .B1(n10284), .B2(n14969), .ZN(
        P2_U3507) );
  AOI22_X1 U16613 ( .A1(n13616), .A2(n14970), .B1(n9148), .B2(n14969), .ZN(
        P2_U3510) );
  NOR2_X1 U16614 ( .A1(P3_U3897), .A2(n15068), .ZN(P3_U3150) );
  NOR2_X1 U16615 ( .A1(n14971), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n14973) );
  NOR2_X1 U16616 ( .A1(n14973), .A2(n14972), .ZN(n14989) );
  NOR2_X1 U16617 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15284), .ZN(n14974) );
  AOI21_X1 U16618 ( .B1(n15068), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n14974), .ZN(
        n14975) );
  OAI21_X1 U16619 ( .B1(n15052), .B2(n14976), .A(n14975), .ZN(n14984) );
  INV_X1 U16620 ( .A(n14977), .ZN(n14978) );
  NAND3_X1 U16621 ( .A1(n14980), .A2(n14979), .A3(n14978), .ZN(n14981) );
  AOI21_X1 U16622 ( .B1(n14982), .B2(n14981), .A(n15054), .ZN(n14983) );
  NOR2_X1 U16623 ( .A1(n14984), .A2(n14983), .ZN(n14988) );
  XNOR2_X1 U16624 ( .A(n14985), .B(P3_REG1_REG_3__SCAN_IN), .ZN(n14986) );
  NAND2_X1 U16625 ( .A1(n15069), .A2(n14986), .ZN(n14987) );
  OAI211_X1 U16626 ( .C1(n14989), .C2(n15063), .A(n14988), .B(n14987), .ZN(
        P3_U3185) );
  NOR2_X1 U16627 ( .A1(n14991), .A2(n14990), .ZN(n14992) );
  OAI21_X1 U16628 ( .B1(n14993), .B2(n14992), .A(n15078), .ZN(n15004) );
  OAI21_X1 U16629 ( .B1(n14996), .B2(n14995), .A(n14994), .ZN(n15002) );
  AOI21_X1 U16630 ( .B1(n14999), .B2(n14998), .A(n14997), .ZN(n15000) );
  INV_X1 U16631 ( .A(n15000), .ZN(n15001) );
  AOI22_X1 U16632 ( .A1(n15069), .A2(n15002), .B1(n15082), .B2(n15001), .ZN(
        n15003) );
  OAI211_X1 U16633 ( .C1(n15052), .C2(n15005), .A(n15004), .B(n15003), .ZN(
        n15006) );
  INV_X1 U16634 ( .A(n15006), .ZN(n15008) );
  OAI211_X1 U16635 ( .C1(n15009), .C2(n15043), .A(n15008), .B(n15007), .ZN(
        P3_U3186) );
  INV_X1 U16636 ( .A(n15010), .ZN(n15012) );
  NAND2_X1 U16637 ( .A1(n15012), .A2(n15011), .ZN(n15013) );
  XNOR2_X1 U16638 ( .A(n15014), .B(n15013), .ZN(n15025) );
  OAI21_X1 U16639 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n15016), .A(n15015), .ZN(
        n15021) );
  AOI21_X1 U16640 ( .B1(n15018), .B2(n10816), .A(n15017), .ZN(n15019) );
  NOR2_X1 U16641 ( .A1(n15063), .A2(n15019), .ZN(n15020) );
  AOI21_X1 U16642 ( .B1(n15069), .B2(n15021), .A(n15020), .ZN(n15022) );
  OAI21_X1 U16643 ( .B1(n15023), .B2(n15052), .A(n15022), .ZN(n15024) );
  AOI21_X1 U16644 ( .B1(n15025), .B2(n15078), .A(n15024), .ZN(n15027) );
  OAI211_X1 U16645 ( .C1(n15028), .C2(n15043), .A(n15027), .B(n15026), .ZN(
        P3_U3187) );
  XNOR2_X1 U16646 ( .A(n15030), .B(n15029), .ZN(n15040) );
  AOI21_X1 U16647 ( .B1(n11414), .B2(n15032), .A(n15031), .ZN(n15033) );
  NOR2_X1 U16648 ( .A1(n15033), .A2(n15063), .ZN(n15039) );
  XNOR2_X1 U16649 ( .A(n15034), .B(n8564), .ZN(n15037) );
  OAI22_X1 U16650 ( .A1(n15037), .A2(n15036), .B1(n15035), .B2(n15052), .ZN(
        n15038) );
  AOI211_X1 U16651 ( .C1(n15040), .C2(n15078), .A(n15039), .B(n15038), .ZN(
        n15042) );
  OAI211_X1 U16652 ( .C1(n15044), .C2(n15043), .A(n15042), .B(n15041), .ZN(
        P3_U3189) );
  AOI21_X1 U16653 ( .B1(n15047), .B2(n15046), .A(n15045), .ZN(n15064) );
  NOR2_X1 U16654 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8601), .ZN(n15057) );
  INV_X1 U16655 ( .A(n15074), .ZN(n15051) );
  OR2_X1 U16656 ( .A1(n15048), .A2(n15074), .ZN(n15049) );
  AOI22_X1 U16657 ( .A1(n15075), .A2(n15051), .B1(n15050), .B2(n15049), .ZN(
        n15055) );
  OAI22_X1 U16658 ( .A1(n15055), .A2(n15054), .B1(n15053), .B2(n15052), .ZN(
        n15056) );
  AOI211_X1 U16659 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n15068), .A(n15057), .B(
        n15056), .ZN(n15062) );
  OAI21_X1 U16660 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n15059), .A(n15058), .ZN(
        n15060) );
  NAND2_X1 U16661 ( .A1(n15060), .A2(n15069), .ZN(n15061) );
  OAI211_X1 U16662 ( .C1(n15064), .C2(n15063), .A(n15062), .B(n15061), .ZN(
        P3_U3191) );
  INV_X1 U16663 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n15267) );
  OAI21_X1 U16664 ( .B1(n15067), .B2(n15066), .A(n15065), .ZN(n15070) );
  AOI22_X1 U16665 ( .A1(n15070), .A2(n15069), .B1(n15068), .B2(
        P3_ADDR_REG_10__SCAN_IN), .ZN(n15085) );
  OAI21_X1 U16666 ( .B1(n7001), .B2(n7000), .A(n15072), .ZN(n15083) );
  OR3_X1 U16667 ( .A1(n15075), .A2(n15074), .A3(n15073), .ZN(n15076) );
  NAND2_X1 U16668 ( .A1(n15077), .A2(n15076), .ZN(n15079) );
  AOI222_X1 U16669 ( .A1(n15083), .A2(n15082), .B1(n15081), .B2(n15080), .C1(
        n15079), .C2(n15078), .ZN(n15084) );
  OAI211_X1 U16670 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n15267), .A(n15085), .B(
        n15084), .ZN(P3_U3192) );
  OAI21_X1 U16671 ( .B1(n15087), .B2(n12179), .A(n15086), .ZN(n15127) );
  NOR2_X1 U16672 ( .A1(n15088), .A2(n15168), .ZN(n15126) );
  INV_X1 U16673 ( .A(n15126), .ZN(n15089) );
  OAI22_X1 U16674 ( .A1(n15090), .A2(n15089), .B1(n15112), .B2(n15226), .ZN(
        n15099) );
  INV_X1 U16675 ( .A(n15127), .ZN(n15098) );
  AOI22_X1 U16676 ( .A1(n15103), .A2(n9764), .B1(n15091), .B2(n15104), .ZN(
        n15097) );
  OAI21_X1 U16677 ( .B1(n15094), .B2(n15093), .A(n15092), .ZN(n15095) );
  NAND2_X1 U16678 ( .A1(n15095), .A2(n15106), .ZN(n15096) );
  OAI211_X1 U16679 ( .C1(n15098), .C2(n15110), .A(n15097), .B(n15096), .ZN(
        n15125) );
  AOI211_X1 U16680 ( .C1(n15100), .C2(n15127), .A(n15099), .B(n15125), .ZN(
        n15101) );
  AOI22_X1 U16681 ( .A1(n15119), .A2(n10766), .B1(n15101), .B2(n15117), .ZN(
        P3_U3231) );
  AND2_X1 U16682 ( .A1(n8498), .A2(n15150), .ZN(n15122) );
  XNOR2_X1 U16683 ( .A(n15105), .B(n15102), .ZN(n15120) );
  AOI22_X1 U16684 ( .A1(n15104), .A2(n9772), .B1(n8497), .B2(n15103), .ZN(
        n15109) );
  XNOR2_X1 U16685 ( .A(n15105), .B(n9767), .ZN(n15107) );
  NAND2_X1 U16686 ( .A1(n15107), .A2(n15106), .ZN(n15108) );
  OAI211_X1 U16687 ( .C1(n15120), .C2(n15110), .A(n15109), .B(n15108), .ZN(
        n15121) );
  AOI21_X1 U16688 ( .B1(n15122), .B2(n15111), .A(n15121), .ZN(n15118) );
  OAI22_X1 U16689 ( .A1(n15114), .A2(n15120), .B1(n15113), .B2(n15112), .ZN(
        n15115) );
  INV_X1 U16690 ( .A(n15115), .ZN(n15116) );
  OAI221_X1 U16691 ( .B1(n15119), .B2(n15118), .C1(n15117), .C2(n10726), .A(
        n15116), .ZN(P3_U3232) );
  INV_X1 U16692 ( .A(n15120), .ZN(n15123) );
  AOI211_X1 U16693 ( .C1(n15164), .C2(n15123), .A(n15122), .B(n15121), .ZN(
        n15176) );
  INV_X1 U16694 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15124) );
  AOI22_X1 U16695 ( .A1(n15175), .A2(n15176), .B1(n15124), .B2(n15173), .ZN(
        P3_U3393) );
  AOI211_X1 U16696 ( .C1(n15164), .C2(n15127), .A(n15126), .B(n15125), .ZN(
        n15177) );
  INV_X1 U16697 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15128) );
  AOI22_X1 U16698 ( .A1(n15175), .A2(n15177), .B1(n15128), .B2(n15173), .ZN(
        P3_U3396) );
  OAI22_X1 U16699 ( .A1(n15130), .A2(n15169), .B1(n15168), .B2(n15129), .ZN(
        n15131) );
  NOR2_X1 U16700 ( .A1(n15132), .A2(n15131), .ZN(n15178) );
  INV_X1 U16701 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15133) );
  AOI22_X1 U16702 ( .A1(n15175), .A2(n15178), .B1(n15133), .B2(n15173), .ZN(
        P3_U3399) );
  NOR2_X1 U16703 ( .A1(n15134), .A2(n15168), .ZN(n15136) );
  AOI211_X1 U16704 ( .C1(n15164), .C2(n15137), .A(n15136), .B(n15135), .ZN(
        n15179) );
  INV_X1 U16705 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15138) );
  AOI22_X1 U16706 ( .A1(n15175), .A2(n15179), .B1(n15138), .B2(n15173), .ZN(
        P3_U3402) );
  OAI22_X1 U16707 ( .A1(n15140), .A2(n15169), .B1(n15168), .B2(n15139), .ZN(
        n15141) );
  NOR2_X1 U16708 ( .A1(n15142), .A2(n15141), .ZN(n15180) );
  INV_X1 U16709 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15143) );
  AOI22_X1 U16710 ( .A1(n15175), .A2(n15180), .B1(n15143), .B2(n15173), .ZN(
        P3_U3405) );
  OAI22_X1 U16711 ( .A1(n15145), .A2(n15169), .B1(n15144), .B2(n15168), .ZN(
        n15146) );
  NOR2_X1 U16712 ( .A1(n15147), .A2(n15146), .ZN(n15181) );
  INV_X1 U16713 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15148) );
  AOI22_X1 U16714 ( .A1(n15175), .A2(n15181), .B1(n15148), .B2(n15173), .ZN(
        P3_U3408) );
  AOI22_X1 U16715 ( .A1(n15151), .A2(n15164), .B1(n15150), .B2(n15149), .ZN(
        n15152) );
  AND2_X1 U16716 ( .A1(n15153), .A2(n15152), .ZN(n15182) );
  INV_X1 U16717 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15154) );
  AOI22_X1 U16718 ( .A1(n15175), .A2(n15182), .B1(n15154), .B2(n15173), .ZN(
        P3_U3411) );
  OAI22_X1 U16719 ( .A1(n15156), .A2(n15169), .B1(n15155), .B2(n15168), .ZN(
        n15157) );
  NOR2_X1 U16720 ( .A1(n15158), .A2(n15157), .ZN(n15184) );
  INV_X1 U16721 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15159) );
  AOI22_X1 U16722 ( .A1(n15175), .A2(n15184), .B1(n15159), .B2(n15173), .ZN(
        P3_U3414) );
  INV_X1 U16723 ( .A(n15160), .ZN(n15165) );
  NOR2_X1 U16724 ( .A1(n15161), .A2(n15168), .ZN(n15163) );
  AOI211_X1 U16725 ( .C1(n15165), .C2(n15164), .A(n15163), .B(n15162), .ZN(
        n15186) );
  INV_X1 U16726 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15166) );
  AOI22_X1 U16727 ( .A1(n15175), .A2(n15186), .B1(n15166), .B2(n15173), .ZN(
        P3_U3417) );
  OAI22_X1 U16728 ( .A1(n15170), .A2(n15169), .B1(n15168), .B2(n15167), .ZN(
        n15171) );
  NOR2_X1 U16729 ( .A1(n15172), .A2(n15171), .ZN(n15187) );
  INV_X1 U16730 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15174) );
  AOI22_X1 U16731 ( .A1(n15175), .A2(n15187), .B1(n15174), .B2(n15173), .ZN(
        P3_U3420) );
  AOI22_X1 U16732 ( .A1(n15183), .A2(n15176), .B1(n10745), .B2(n9886), .ZN(
        P3_U3460) );
  AOI22_X1 U16733 ( .A1(n15183), .A2(n15177), .B1(n10765), .B2(n9886), .ZN(
        P3_U3461) );
  AOI22_X1 U16734 ( .A1(n15183), .A2(n15178), .B1(n10806), .B2(n9886), .ZN(
        P3_U3462) );
  AOI22_X1 U16735 ( .A1(n15183), .A2(n15179), .B1(n10841), .B2(n9886), .ZN(
        P3_U3463) );
  AOI22_X1 U16736 ( .A1(n15183), .A2(n15180), .B1(n10815), .B2(n9886), .ZN(
        P3_U3464) );
  AOI22_X1 U16737 ( .A1(n15183), .A2(n15181), .B1(n10845), .B2(n9886), .ZN(
        P3_U3465) );
  AOI22_X1 U16738 ( .A1(n15183), .A2(n15182), .B1(n8564), .B2(n9886), .ZN(
        P3_U3466) );
  AOI22_X1 U16739 ( .A1(n15183), .A2(n15184), .B1(n10862), .B2(n9886), .ZN(
        P3_U3467) );
  AOI22_X1 U16740 ( .A1(n15183), .A2(n15186), .B1(n15185), .B2(n9886), .ZN(
        P3_U3468) );
  AOI22_X1 U16741 ( .A1(n15183), .A2(n15187), .B1(n11387), .B2(n9886), .ZN(
        P3_U3469) );
  AOI22_X1 U16742 ( .A1(SI_23_), .A2(keyinput_f9), .B1(SI_25_), .B2(
        keyinput_f7), .ZN(n15188) );
  OAI221_X1 U16743 ( .B1(SI_23_), .B2(keyinput_f9), .C1(SI_25_), .C2(
        keyinput_f7), .A(n15188), .ZN(n15195) );
  AOI22_X1 U16744 ( .A1(SI_24_), .A2(keyinput_f8), .B1(P3_REG3_REG_23__SCAN_IN), .B2(keyinput_f38), .ZN(n15189) );
  OAI221_X1 U16745 ( .B1(SI_24_), .B2(keyinput_f8), .C1(
        P3_REG3_REG_23__SCAN_IN), .C2(keyinput_f38), .A(n15189), .ZN(n15194)
         );
  AOI22_X1 U16746 ( .A1(keyinput_f0), .A2(P3_WR_REG_SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(keyinput_f44), .ZN(n15190) );
  OAI221_X1 U16747 ( .B1(keyinput_f0), .B2(P3_WR_REG_SCAN_IN), .C1(
        P3_REG3_REG_1__SCAN_IN), .C2(keyinput_f44), .A(n15190), .ZN(n15193) );
  AOI22_X1 U16748 ( .A1(SI_20_), .A2(keyinput_f12), .B1(
        P3_REG3_REG_19__SCAN_IN), .B2(keyinput_f41), .ZN(n15191) );
  OAI221_X1 U16749 ( .B1(SI_20_), .B2(keyinput_f12), .C1(
        P3_REG3_REG_19__SCAN_IN), .C2(keyinput_f41), .A(n15191), .ZN(n15192)
         );
  NOR4_X1 U16750 ( .A1(n15195), .A2(n15194), .A3(n15193), .A4(n15192), .ZN(
        n15222) );
  XNOR2_X1 U16751 ( .A(P3_REG3_REG_0__SCAN_IN), .B(keyinput_f54), .ZN(n15202)
         );
  AOI22_X1 U16752 ( .A1(P3_STATE_REG_SCAN_IN), .A2(keyinput_f34), .B1(n15331), 
        .B2(keyinput_f26), .ZN(n15196) );
  OAI221_X1 U16753 ( .B1(P3_STATE_REG_SCAN_IN), .B2(keyinput_f34), .C1(n15331), 
        .C2(keyinput_f26), .A(n15196), .ZN(n15201) );
  AOI22_X1 U16754 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(keyinput_f52), .B1(
        P3_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .ZN(n15197) );
  OAI221_X1 U16755 ( .B1(P3_REG3_REG_4__SCAN_IN), .B2(keyinput_f52), .C1(
        P3_REG3_REG_26__SCAN_IN), .C2(keyinput_f62), .A(n15197), .ZN(n15200)
         );
  AOI22_X1 U16756 ( .A1(P3_REG3_REG_11__SCAN_IN), .A2(keyinput_f58), .B1(
        P3_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .ZN(n15198) );
  OAI221_X1 U16757 ( .B1(P3_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .C1(
        P3_REG3_REG_28__SCAN_IN), .C2(keyinput_f42), .A(n15198), .ZN(n15199)
         );
  NOR4_X1 U16758 ( .A1(n15202), .A2(n15201), .A3(n15200), .A4(n15199), .ZN(
        n15221) );
  AOI22_X1 U16759 ( .A1(SI_19_), .A2(keyinput_f13), .B1(
        P3_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .ZN(n15203) );
  OAI221_X1 U16760 ( .B1(SI_19_), .B2(keyinput_f13), .C1(
        P3_REG3_REG_18__SCAN_IN), .C2(keyinput_f60), .A(n15203), .ZN(n15210)
         );
  AOI22_X1 U16761 ( .A1(SI_11_), .A2(keyinput_f21), .B1(P3_REG3_REG_6__SCAN_IN), .B2(keyinput_f61), .ZN(n15204) );
  OAI221_X1 U16762 ( .B1(SI_11_), .B2(keyinput_f21), .C1(
        P3_REG3_REG_6__SCAN_IN), .C2(keyinput_f61), .A(n15204), .ZN(n15209) );
  AOI22_X1 U16763 ( .A1(SI_5_), .A2(keyinput_f27), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(keyinput_f40), .ZN(n15205) );
  OAI221_X1 U16764 ( .B1(SI_5_), .B2(keyinput_f27), .C1(P3_REG3_REG_3__SCAN_IN), .C2(keyinput_f40), .A(n15205), .ZN(n15208) );
  AOI22_X1 U16765 ( .A1(P3_REG3_REG_22__SCAN_IN), .A2(keyinput_f57), .B1(
        P3_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .ZN(n15206) );
  OAI221_X1 U16766 ( .B1(P3_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .C1(
        P3_REG3_REG_24__SCAN_IN), .C2(keyinput_f51), .A(n15206), .ZN(n15207)
         );
  NOR4_X1 U16767 ( .A1(n15210), .A2(n15209), .A3(n15208), .A4(n15207), .ZN(
        n15220) );
  AOI22_X1 U16768 ( .A1(SI_22_), .A2(keyinput_f10), .B1(
        P3_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .ZN(n15211) );
  OAI221_X1 U16769 ( .B1(SI_22_), .B2(keyinput_f10), .C1(
        P3_REG3_REG_27__SCAN_IN), .C2(keyinput_f36), .A(n15211), .ZN(n15218)
         );
  AOI22_X1 U16770 ( .A1(SI_3_), .A2(keyinput_f29), .B1(SI_4_), .B2(
        keyinput_f28), .ZN(n15212) );
  OAI221_X1 U16771 ( .B1(SI_3_), .B2(keyinput_f29), .C1(SI_4_), .C2(
        keyinput_f28), .A(n15212), .ZN(n15217) );
  AOI22_X1 U16772 ( .A1(SI_2_), .A2(keyinput_f30), .B1(P3_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .ZN(n15213) );
  OAI221_X1 U16773 ( .B1(SI_2_), .B2(keyinput_f30), .C1(
        P3_REG3_REG_12__SCAN_IN), .C2(keyinput_f46), .A(n15213), .ZN(n15216)
         );
  AOI22_X1 U16774 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(keyinput_f53), .B1(
        P3_REG3_REG_17__SCAN_IN), .B2(keyinput_f50), .ZN(n15214) );
  OAI221_X1 U16775 ( .B1(P3_REG3_REG_9__SCAN_IN), .B2(keyinput_f53), .C1(
        P3_REG3_REG_17__SCAN_IN), .C2(keyinput_f50), .A(n15214), .ZN(n15215)
         );
  NOR4_X1 U16776 ( .A1(n15218), .A2(n15217), .A3(n15216), .A4(n15215), .ZN(
        n15219) );
  NAND4_X1 U16777 ( .A1(n15222), .A2(n15221), .A3(n15220), .A4(n15219), .ZN(
        n15278) );
  INV_X1 U16778 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n15313) );
  AOI22_X1 U16779 ( .A1(n15313), .A2(keyinput_f35), .B1(keyinput_f17), .B2(
        n15224), .ZN(n15223) );
  OAI221_X1 U16780 ( .B1(n15313), .B2(keyinput_f35), .C1(n15224), .C2(
        keyinput_f17), .A(n15223), .ZN(n15234) );
  AOI22_X1 U16781 ( .A1(n15227), .A2(keyinput_f63), .B1(keyinput_f59), .B2(
        n15226), .ZN(n15225) );
  OAI221_X1 U16782 ( .B1(n15227), .B2(keyinput_f63), .C1(n15226), .C2(
        keyinput_f59), .A(n15225), .ZN(n15233) );
  AOI22_X1 U16783 ( .A1(n13066), .A2(keyinput_f1), .B1(keyinput_f2), .B2(
        n15229), .ZN(n15228) );
  OAI221_X1 U16784 ( .B1(n13066), .B2(keyinput_f1), .C1(n15229), .C2(
        keyinput_f2), .A(n15228), .ZN(n15232) );
  AOI22_X1 U16785 ( .A1(n15330), .A2(keyinput_f48), .B1(keyinput_f49), .B2(
        n15288), .ZN(n15230) );
  OAI221_X1 U16786 ( .B1(n15330), .B2(keyinput_f48), .C1(n15288), .C2(
        keyinput_f49), .A(n15230), .ZN(n15231) );
  NOR4_X1 U16787 ( .A1(n15234), .A2(n15233), .A3(n15232), .A4(n15231), .ZN(
        n15276) );
  AOI22_X1 U16788 ( .A1(n15312), .A2(keyinput_f20), .B1(n15236), .B2(
        keyinput_f4), .ZN(n15235) );
  OAI221_X1 U16789 ( .B1(n15312), .B2(keyinput_f20), .C1(n15236), .C2(
        keyinput_f4), .A(n15235), .ZN(n15245) );
  AOI22_X1 U16790 ( .A1(n7562), .A2(keyinput_f31), .B1(n15238), .B2(
        keyinput_f37), .ZN(n15237) );
  OAI221_X1 U16791 ( .B1(n7562), .B2(keyinput_f31), .C1(n15238), .C2(
        keyinput_f37), .A(n15237), .ZN(n15244) );
  AOI22_X1 U16792 ( .A1(SI_26_), .A2(keyinput_f6), .B1(n15301), .B2(
        keyinput_f43), .ZN(n15239) );
  OAI221_X1 U16793 ( .B1(SI_26_), .B2(keyinput_f6), .C1(n15301), .C2(
        keyinput_f43), .A(n15239), .ZN(n15243) );
  XNOR2_X1 U16794 ( .A(P3_REG3_REG_20__SCAN_IN), .B(keyinput_f55), .ZN(n15241)
         );
  XNOR2_X1 U16795 ( .A(SI_0_), .B(keyinput_f32), .ZN(n15240) );
  NAND2_X1 U16796 ( .A1(n15241), .A2(n15240), .ZN(n15242) );
  NOR4_X1 U16797 ( .A1(n15245), .A2(n15244), .A3(n15243), .A4(n15242), .ZN(
        n15275) );
  AOI22_X1 U16798 ( .A1(n15248), .A2(keyinput_f22), .B1(n15247), .B2(
        keyinput_f16), .ZN(n15246) );
  OAI221_X1 U16799 ( .B1(n15248), .B2(keyinput_f22), .C1(n15247), .C2(
        keyinput_f16), .A(n15246), .ZN(n15258) );
  AOI22_X1 U16800 ( .A1(n15250), .A2(keyinput_f25), .B1(n11927), .B2(
        keyinput_f56), .ZN(n15249) );
  OAI221_X1 U16801 ( .B1(n15250), .B2(keyinput_f25), .C1(n11927), .C2(
        keyinput_f56), .A(n15249), .ZN(n15257) );
  INV_X1 U16802 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n15253) );
  AOI22_X1 U16803 ( .A1(n15253), .A2(keyinput_f47), .B1(keyinput_f14), .B2(
        n15252), .ZN(n15251) );
  OAI221_X1 U16804 ( .B1(n15253), .B2(keyinput_f47), .C1(n15252), .C2(
        keyinput_f14), .A(n15251), .ZN(n15256) );
  AOI22_X1 U16805 ( .A1(n8763), .A2(keyinput_f45), .B1(keyinput_f33), .B2(
        n15296), .ZN(n15254) );
  OAI221_X1 U16806 ( .B1(n8763), .B2(keyinput_f45), .C1(n15296), .C2(
        keyinput_f33), .A(n15254), .ZN(n15255) );
  NOR4_X1 U16807 ( .A1(n15258), .A2(n15257), .A3(n15256), .A4(n15255), .ZN(
        n15274) );
  AOI22_X1 U16808 ( .A1(n15261), .A2(keyinput_f19), .B1(n15260), .B2(
        keyinput_f11), .ZN(n15259) );
  OAI221_X1 U16809 ( .B1(n15261), .B2(keyinput_f19), .C1(n15260), .C2(
        keyinput_f11), .A(n15259), .ZN(n15272) );
  AOI22_X1 U16810 ( .A1(n15263), .A2(keyinput_f18), .B1(keyinput_f3), .B2(
        n15285), .ZN(n15262) );
  OAI221_X1 U16811 ( .B1(n15263), .B2(keyinput_f18), .C1(n15285), .C2(
        keyinput_f3), .A(n15262), .ZN(n15271) );
  AOI22_X1 U16812 ( .A1(n15327), .A2(keyinput_f15), .B1(n15265), .B2(
        keyinput_f5), .ZN(n15264) );
  OAI221_X1 U16813 ( .B1(n15327), .B2(keyinput_f15), .C1(n15265), .C2(
        keyinput_f5), .A(n15264), .ZN(n15270) );
  AOI22_X1 U16814 ( .A1(n15268), .A2(keyinput_f23), .B1(n15267), .B2(
        keyinput_f39), .ZN(n15266) );
  OAI221_X1 U16815 ( .B1(n15268), .B2(keyinput_f23), .C1(n15267), .C2(
        keyinput_f39), .A(n15266), .ZN(n15269) );
  NOR4_X1 U16816 ( .A1(n15272), .A2(n15271), .A3(n15270), .A4(n15269), .ZN(
        n15273) );
  NAND4_X1 U16817 ( .A1(n15276), .A2(n15275), .A3(n15274), .A4(n15273), .ZN(
        n15277) );
  OAI22_X1 U16818 ( .A1(n15278), .A2(n15277), .B1(keyinput_f24), .B2(SI_8_), 
        .ZN(n15279) );
  AOI21_X1 U16819 ( .B1(keyinput_f24), .B2(SI_8_), .A(n15279), .ZN(n15378) );
  AOI22_X1 U16820 ( .A1(n15282), .A2(keyinput_g50), .B1(keyinput_g28), .B2(
        n15281), .ZN(n15280) );
  OAI221_X1 U16821 ( .B1(n15282), .B2(keyinput_g50), .C1(n15281), .C2(
        keyinput_g28), .A(n15280), .ZN(n15294) );
  AOI22_X1 U16822 ( .A1(n15285), .A2(keyinput_g3), .B1(n15284), .B2(
        keyinput_g40), .ZN(n15283) );
  OAI221_X1 U16823 ( .B1(n15285), .B2(keyinput_g3), .C1(n15284), .C2(
        keyinput_g40), .A(n15283), .ZN(n15293) );
  AOI22_X1 U16824 ( .A1(n15288), .A2(keyinput_g49), .B1(keyinput_g8), .B2(
        n15287), .ZN(n15286) );
  OAI221_X1 U16825 ( .B1(n15288), .B2(keyinput_g49), .C1(n15287), .C2(
        keyinput_g8), .A(n15286), .ZN(n15292) );
  INV_X1 U16826 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n15290) );
  AOI22_X1 U16827 ( .A1(P3_U3151), .A2(keyinput_g34), .B1(keyinput_g52), .B2(
        n15290), .ZN(n15289) );
  OAI221_X1 U16828 ( .B1(P3_U3151), .B2(keyinput_g34), .C1(n15290), .C2(
        keyinput_g52), .A(n15289), .ZN(n15291) );
  NOR4_X1 U16829 ( .A1(n15294), .A2(n15293), .A3(n15292), .A4(n15291), .ZN(
        n15339) );
  INV_X1 U16830 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n15297) );
  AOI22_X1 U16831 ( .A1(n15297), .A2(keyinput_g38), .B1(keyinput_g33), .B2(
        n15296), .ZN(n15295) );
  OAI221_X1 U16832 ( .B1(n15297), .B2(keyinput_g38), .C1(n15296), .C2(
        keyinput_g33), .A(n15295), .ZN(n15308) );
  AOI22_X1 U16833 ( .A1(P3_REG3_REG_0__SCAN_IN), .A2(keyinput_g54), .B1(
        P3_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .ZN(n15298) );
  OAI221_X1 U16834 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .C1(
        P3_REG3_REG_14__SCAN_IN), .C2(keyinput_g37), .A(n15298), .ZN(n15307)
         );
  INV_X1 U16835 ( .A(P3_WR_REG_SCAN_IN), .ZN(n15300) );
  AOI22_X1 U16836 ( .A1(n15301), .A2(keyinput_g43), .B1(keyinput_g0), .B2(
        n15300), .ZN(n15299) );
  OAI221_X1 U16837 ( .B1(n15301), .B2(keyinput_g43), .C1(n15300), .C2(
        keyinput_g0), .A(n15299), .ZN(n15306) );
  AOI22_X1 U16838 ( .A1(n15304), .A2(keyinput_g7), .B1(n15303), .B2(
        keyinput_g36), .ZN(n15302) );
  OAI221_X1 U16839 ( .B1(n15304), .B2(keyinput_g7), .C1(n15303), .C2(
        keyinput_g36), .A(n15302), .ZN(n15305) );
  NOR4_X1 U16840 ( .A1(n15308), .A2(n15307), .A3(n15306), .A4(n15305), .ZN(
        n15338) );
  AOI22_X1 U16841 ( .A1(n15310), .A2(keyinput_g6), .B1(n8763), .B2(
        keyinput_g45), .ZN(n15309) );
  OAI221_X1 U16842 ( .B1(n15310), .B2(keyinput_g6), .C1(n8763), .C2(
        keyinput_g45), .A(n15309), .ZN(n15322) );
  AOI22_X1 U16843 ( .A1(n15313), .A2(keyinput_g35), .B1(keyinput_g20), .B2(
        n15312), .ZN(n15311) );
  OAI221_X1 U16844 ( .B1(n15313), .B2(keyinput_g35), .C1(n15312), .C2(
        keyinput_g20), .A(n15311), .ZN(n15321) );
  INV_X1 U16845 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n15316) );
  AOI22_X1 U16846 ( .A1(n15316), .A2(keyinput_g58), .B1(keyinput_g21), .B2(
        n15315), .ZN(n15314) );
  OAI221_X1 U16847 ( .B1(n15316), .B2(keyinput_g58), .C1(n15315), .C2(
        keyinput_g21), .A(n15314), .ZN(n15320) );
  XNOR2_X1 U16848 ( .A(SI_2_), .B(keyinput_g30), .ZN(n15318) );
  XNOR2_X1 U16849 ( .A(SI_14_), .B(keyinput_g18), .ZN(n15317) );
  NAND2_X1 U16850 ( .A1(n15318), .A2(n15317), .ZN(n15319) );
  NOR4_X1 U16851 ( .A1(n15322), .A2(n15321), .A3(n15320), .A4(n15319), .ZN(
        n15337) );
  AOI22_X1 U16852 ( .A1(n15325), .A2(keyinput_g62), .B1(keyinput_g12), .B2(
        n15324), .ZN(n15323) );
  OAI221_X1 U16853 ( .B1(n15325), .B2(keyinput_g62), .C1(n15324), .C2(
        keyinput_g12), .A(n15323), .ZN(n15335) );
  AOI22_X1 U16854 ( .A1(n15327), .A2(keyinput_g15), .B1(n8601), .B2(
        keyinput_g53), .ZN(n15326) );
  OAI221_X1 U16855 ( .B1(n15327), .B2(keyinput_g15), .C1(n8601), .C2(
        keyinput_g53), .A(n15326), .ZN(n15334) );
  AOI22_X1 U16856 ( .A1(n8832), .A2(keyinput_g42), .B1(keyinput_g31), .B2(
        n7562), .ZN(n15328) );
  OAI221_X1 U16857 ( .B1(n8832), .B2(keyinput_g42), .C1(n7562), .C2(
        keyinput_g31), .A(n15328), .ZN(n15333) );
  AOI22_X1 U16858 ( .A1(n15331), .A2(keyinput_g26), .B1(n15330), .B2(
        keyinput_g48), .ZN(n15329) );
  OAI221_X1 U16859 ( .B1(n15331), .B2(keyinput_g26), .C1(n15330), .C2(
        keyinput_g48), .A(n15329), .ZN(n15332) );
  NOR4_X1 U16860 ( .A1(n15335), .A2(n15334), .A3(n15333), .A4(n15332), .ZN(
        n15336) );
  NAND4_X1 U16861 ( .A1(n15339), .A2(n15338), .A3(n15337), .A4(n15336), .ZN(
        n15376) );
  AOI22_X1 U16862 ( .A1(SI_18_), .A2(keyinput_g14), .B1(
        P3_REG3_REG_24__SCAN_IN), .B2(keyinput_g51), .ZN(n15340) );
  OAI221_X1 U16863 ( .B1(SI_18_), .B2(keyinput_g14), .C1(
        P3_REG3_REG_24__SCAN_IN), .C2(keyinput_g51), .A(n15340), .ZN(n15347)
         );
  AOI22_X1 U16864 ( .A1(SI_23_), .A2(keyinput_g9), .B1(P3_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .ZN(n15341) );
  OAI221_X1 U16865 ( .B1(SI_23_), .B2(keyinput_g9), .C1(
        P3_REG3_REG_19__SCAN_IN), .C2(keyinput_g41), .A(n15341), .ZN(n15346)
         );
  AOI22_X1 U16866 ( .A1(SI_0_), .A2(keyinput_g32), .B1(SI_19_), .B2(
        keyinput_g13), .ZN(n15342) );
  OAI221_X1 U16867 ( .B1(SI_0_), .B2(keyinput_g32), .C1(SI_19_), .C2(
        keyinput_g13), .A(n15342), .ZN(n15345) );
  AOI22_X1 U16868 ( .A1(SI_27_), .A2(keyinput_g5), .B1(SI_28_), .B2(
        keyinput_g4), .ZN(n15343) );
  OAI221_X1 U16869 ( .B1(SI_27_), .B2(keyinput_g5), .C1(SI_28_), .C2(
        keyinput_g4), .A(n15343), .ZN(n15344) );
  NOR4_X1 U16870 ( .A1(n15347), .A2(n15346), .A3(n15345), .A4(n15344), .ZN(
        n15374) );
  XOR2_X1 U16871 ( .A(SI_30_), .B(keyinput_g2), .Z(n15354) );
  AOI22_X1 U16872 ( .A1(P3_REG3_REG_13__SCAN_IN), .A2(keyinput_g56), .B1(
        P3_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .ZN(n15348) );
  OAI221_X1 U16873 ( .B1(P3_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .C1(
        P3_REG3_REG_18__SCAN_IN), .C2(keyinput_g60), .A(n15348), .ZN(n15353)
         );
  AOI22_X1 U16874 ( .A1(P3_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(SI_13_), .B2(keyinput_g19), .ZN(n15349) );
  OAI221_X1 U16875 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(
        SI_13_), .C2(keyinput_g19), .A(n15349), .ZN(n15352) );
  AOI22_X1 U16876 ( .A1(P3_REG3_REG_1__SCAN_IN), .A2(keyinput_g44), .B1(
        P3_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .ZN(n15350) );
  OAI221_X1 U16877 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(keyinput_g44), .C1(
        P3_REG3_REG_22__SCAN_IN), .C2(keyinput_g57), .A(n15350), .ZN(n15351)
         );
  NOR4_X1 U16878 ( .A1(n15354), .A2(n15353), .A3(n15352), .A4(n15351), .ZN(
        n15373) );
  AOI22_X1 U16879 ( .A1(SI_5_), .A2(keyinput_g27), .B1(P3_REG3_REG_6__SCAN_IN), 
        .B2(keyinput_g61), .ZN(n15355) );
  OAI221_X1 U16880 ( .B1(SI_5_), .B2(keyinput_g27), .C1(P3_REG3_REG_6__SCAN_IN), .C2(keyinput_g61), .A(n15355), .ZN(n15362) );
  AOI22_X1 U16881 ( .A1(SI_16_), .A2(keyinput_g16), .B1(
        P3_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .ZN(n15356) );
  OAI221_X1 U16882 ( .B1(SI_16_), .B2(keyinput_g16), .C1(
        P3_REG3_REG_15__SCAN_IN), .C2(keyinput_g63), .A(n15356), .ZN(n15361)
         );
  AOI22_X1 U16883 ( .A1(SI_10_), .A2(keyinput_g22), .B1(
        P3_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .ZN(n15357) );
  OAI221_X1 U16884 ( .B1(SI_10_), .B2(keyinput_g22), .C1(
        P3_REG3_REG_12__SCAN_IN), .C2(keyinput_g46), .A(n15357), .ZN(n15360)
         );
  AOI22_X1 U16885 ( .A1(SI_7_), .A2(keyinput_g25), .B1(P3_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .ZN(n15358) );
  OAI221_X1 U16886 ( .B1(SI_7_), .B2(keyinput_g25), .C1(
        P3_REG3_REG_20__SCAN_IN), .C2(keyinput_g55), .A(n15358), .ZN(n15359)
         );
  NOR4_X1 U16887 ( .A1(n15362), .A2(n15361), .A3(n15360), .A4(n15359), .ZN(
        n15372) );
  AOI22_X1 U16888 ( .A1(SI_15_), .A2(keyinput_g17), .B1(SI_9_), .B2(
        keyinput_g23), .ZN(n15363) );
  OAI221_X1 U16889 ( .B1(SI_15_), .B2(keyinput_g17), .C1(SI_9_), .C2(
        keyinput_g23), .A(n15363), .ZN(n15370) );
  AOI22_X1 U16890 ( .A1(SI_22_), .A2(keyinput_g10), .B1(
        P3_REG3_REG_25__SCAN_IN), .B2(keyinput_g47), .ZN(n15364) );
  OAI221_X1 U16891 ( .B1(SI_22_), .B2(keyinput_g10), .C1(
        P3_REG3_REG_25__SCAN_IN), .C2(keyinput_g47), .A(n15364), .ZN(n15369)
         );
  AOI22_X1 U16892 ( .A1(SI_3_), .A2(keyinput_g29), .B1(SI_21_), .B2(
        keyinput_g11), .ZN(n15365) );
  OAI221_X1 U16893 ( .B1(SI_3_), .B2(keyinput_g29), .C1(SI_21_), .C2(
        keyinput_g11), .A(n15365), .ZN(n15368) );
  AOI22_X1 U16894 ( .A1(SI_31_), .A2(keyinput_g1), .B1(P3_REG3_REG_10__SCAN_IN), .B2(keyinput_g39), .ZN(n15366) );
  OAI221_X1 U16895 ( .B1(SI_31_), .B2(keyinput_g1), .C1(
        P3_REG3_REG_10__SCAN_IN), .C2(keyinput_g39), .A(n15366), .ZN(n15367)
         );
  NOR4_X1 U16896 ( .A1(n15370), .A2(n15369), .A3(n15368), .A4(n15367), .ZN(
        n15371) );
  NAND4_X1 U16897 ( .A1(n15374), .A2(n15373), .A3(n15372), .A4(n15371), .ZN(
        n15375) );
  OAI22_X1 U16898 ( .A1(keyinput_g24), .A2(n15379), .B1(n15376), .B2(n15375), 
        .ZN(n15377) );
  AOI211_X1 U16899 ( .C1(keyinput_g24), .C2(n15379), .A(n15378), .B(n15377), 
        .ZN(n15393) );
  NOR2_X1 U16900 ( .A1(n15385), .A2(n15384), .ZN(n15386) );
  AOI21_X1 U16901 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n15387), .A(n15386), 
        .ZN(n15390) );
  XNOR2_X1 U16902 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n15388) );
  XNOR2_X1 U16903 ( .A(n15388), .B(n7529), .ZN(n15389) );
  XNOR2_X1 U16904 ( .A(n15390), .B(n15389), .ZN(n15391) );
  OAI21_X1 U16905 ( .B1(n15396), .B2(n15395), .A(n15394), .ZN(SUB_1596_U59) );
  OAI21_X1 U16906 ( .B1(n15399), .B2(n15398), .A(n15397), .ZN(SUB_1596_U58) );
  XOR2_X1 U16907 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15400), .Z(SUB_1596_U53) );
  AOI21_X1 U16908 ( .B1(n15403), .B2(n15402), .A(n15401), .ZN(SUB_1596_U56) );
  OAI21_X1 U16909 ( .B1(n15406), .B2(n15405), .A(n15404), .ZN(n15407) );
  XNOR2_X1 U16910 ( .A(n15407), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  AOI21_X1 U16911 ( .B1(n15410), .B2(n15409), .A(n15408), .ZN(SUB_1596_U5) );
  CLKBUF_X1 U7236 ( .A(n9514), .Z(n9676) );
  CLKBUF_X2 U7295 ( .A(n9777), .Z(n9838) );
  CLKBUF_X1 U7296 ( .A(n7750), .Z(n8212) );
  CLKBUF_X2 U7369 ( .A(n9777), .Z(n12528) );
  CLKBUF_X1 U10023 ( .A(n7520), .Z(n7521) );
endmodule

