

module b14_C_SARLock_k_128_10 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4857, n4858, n4859, n4860, n4861, n4862;

  INV_X1 U2393 ( .A(n3887), .ZN(n2763) );
  INV_X1 U2394 ( .A(n3571), .ZN(n3578) );
  NAND2_X1 U2395 ( .A1(n3042), .A2(n3811), .ZN(n3097) );
  INV_X1 U2396 ( .A(IR_REG_4__SCAN_IN), .ZN(n2374) );
  OAI21_X1 U2397 ( .B1(n3692), .B2(n3462), .A(n3441), .ZN(n4026) );
  CLKBUF_X3 U2398 ( .A(n2572), .Z(n3576) );
  NOR4_X2 U2399 ( .A1(n3766), .A2(n4083), .A3(n3765), .A4(n3764), .ZN(n3785)
         );
  AOI21_X2 U2400 ( .B1(n3097), .B2(n3096), .A(n3818), .ZN(n3245) );
  INV_X4 U2401 ( .A(n2609), .ZN(n3725) );
  NAND2_X1 U2402 ( .A1(n3469), .A2(n3832), .ZN(n4183) );
  NAND2_X1 U2403 ( .A1(n3503), .A2(n3502), .ZN(n3511) );
  AND3_X1 U2404 ( .A1(n2982), .A2(n2246), .A3(n2984), .ZN(n2245) );
  AOI21_X1 U2405 ( .B1(n2916), .B2(n2915), .A(n3804), .ZN(n2932) );
  AND2_X1 U2406 ( .A1(n2842), .A2(n2600), .ZN(n2605) );
  NAND2_X1 U2407 ( .A1(n3230), .A2(n3229), .ZN(n3231) );
  AND2_X2 U2408 ( .A1(n2537), .A2(n2740), .ZN(n3571) );
  AND2_X2 U2409 ( .A1(n2742), .A2(n3859), .ZN(n4510) );
  NAND4_X1 U2410 ( .A1(n2661), .A2(n2660), .A3(n2659), .A4(n2658), .ZN(n3885)
         );
  NAND3_X1 U2411 ( .A1(n2337), .A2(n2583), .A3(n2582), .ZN(n3887) );
  BUF_X2 U2412 ( .A(n2543), .Z(n3445) );
  NAND2_X1 U2413 ( .A1(n2603), .A2(n2602), .ZN(n2757) );
  XNOR2_X1 U2414 ( .A(n2387), .B(IR_REG_30__SCAN_IN), .ZN(n2291) );
  INV_X1 U2419 ( .A(n2363), .ZN(n2326) );
  AND2_X1 U2420 ( .A1(n3638), .A2(n2274), .ZN(n2273) );
  NAND2_X1 U2421 ( .A1(n2276), .A2(n3510), .ZN(n2274) );
  INV_X1 U2422 ( .A(IR_REG_26__SCAN_IN), .ZN(n2414) );
  OAI21_X1 U2423 ( .B1(n2686), .B2(n2253), .A(n2250), .ZN(n2981) );
  NOR2_X1 U2424 ( .A1(n2269), .A2(n3516), .ZN(n2268) );
  INV_X1 U2425 ( .A(n2271), .ZN(n2269) );
  NAND2_X1 U2426 ( .A1(n2517), .A2(n3859), .ZN(n2740) );
  NOR2_X1 U2427 ( .A1(IR_REG_15__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2341)
         );
  NOR2_X1 U2428 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2353)
         );
  NOR2_X1 U2429 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2352)
         );
  NOR2_X1 U2430 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2351)
         );
  NAND2_X1 U2431 ( .A1(n2786), .A2(REG3_REG_7__SCAN_IN), .ZN(n2903) );
  INV_X1 U2433 ( .A(n2159), .ZN(n2609) );
  NAND2_X1 U2434 ( .A1(n2466), .A2(n2465), .ZN(n2468) );
  NAND2_X1 U2435 ( .A1(n2511), .A2(n2475), .ZN(n2699) );
  XNOR2_X1 U2436 ( .A(n3924), .B(n2215), .ZN(n4427) );
  INV_X1 U2437 ( .A(n4472), .ZN(n2215) );
  XNOR2_X1 U2438 ( .A(n2207), .B(n4472), .ZN(n4425) );
  AOI21_X1 U2439 ( .B1(n2151), .B2(n2301), .A(n2294), .ZN(n2293) );
  INV_X1 U2440 ( .A(n3747), .ZN(n2294) );
  INV_X1 U2441 ( .A(n4162), .ZN(n2297) );
  XNOR2_X1 U2442 ( .A(n2468), .B(n4360), .ZN(n4358) );
  NOR2_X1 U2443 ( .A1(n4442), .A2(n4443), .ZN(n4441) );
  INV_X1 U2444 ( .A(n3202), .ZN(n2314) );
  INV_X1 U2445 ( .A(n4331), .ZN(n2263) );
  INV_X1 U2446 ( .A(n3657), .ZN(n2288) );
  AOI21_X1 U2447 ( .B1(n2286), .B2(n2171), .A(n3626), .ZN(n2285) );
  INV_X1 U2448 ( .A(n2291), .ZN(n2290) );
  NAND2_X1 U2449 ( .A1(n2187), .A2(n2186), .ZN(n2328) );
  INV_X1 U2450 ( .A(IR_REG_5__SCAN_IN), .ZN(n2187) );
  INV_X1 U2451 ( .A(IR_REG_6__SCAN_IN), .ZN(n2186) );
  NOR2_X1 U2452 ( .A1(n4379), .A2(n2178), .ZN(n3190) );
  INV_X1 U2453 ( .A(n2303), .ZN(n2302) );
  OR2_X1 U2454 ( .A1(n2564), .A2(n2559), .ZN(n2630) );
  INV_X1 U2455 ( .A(IR_REG_28__SCAN_IN), .ZN(n2417) );
  AND2_X1 U2456 ( .A1(n2152), .A2(n2333), .ZN(n2332) );
  NOR2_X1 U2457 ( .A1(n2163), .A2(IR_REG_25__SCAN_IN), .ZN(n2333) );
  NOR2_X1 U2458 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2344)
         );
  INV_X1 U2459 ( .A(IR_REG_11__SCAN_IN), .ZN(n4737) );
  INV_X1 U2460 ( .A(n3689), .ZN(n2280) );
  NAND2_X1 U2461 ( .A1(n3669), .A2(n3672), .ZN(n3619) );
  OR2_X1 U2462 ( .A1(n2981), .A2(n2980), .ZN(n2982) );
  NOR2_X1 U2463 ( .A1(n3609), .A2(n2265), .ZN(n2264) );
  AOI21_X1 U2464 ( .B1(n2268), .B2(n2272), .A(n2176), .ZN(n2267) );
  NAND2_X1 U2465 ( .A1(n2251), .A2(n2772), .ZN(n2255) );
  AOI21_X1 U2466 ( .B1(n2285), .B2(n2287), .A(n2282), .ZN(n2281) );
  INV_X1 U2467 ( .A(n3627), .ZN(n2282) );
  INV_X1 U2468 ( .A(n2285), .ZN(n2283) );
  INV_X1 U2469 ( .A(n3531), .ZN(n3566) );
  CLKBUF_X1 U2470 ( .A(n2542), .Z(n3729) );
  INV_X1 U2471 ( .A(n3412), .ZN(n3462) );
  OR2_X1 U2472 ( .A1(n4369), .A2(n2707), .ZN(n2708) );
  XNOR2_X1 U2473 ( .A(n3175), .B(n2209), .ZN(n2702) );
  OAI21_X1 U2474 ( .B1(n2948), .B2(n4476), .A(n4374), .ZN(n3175) );
  NAND2_X1 U2475 ( .A1(n2702), .A2(REG2_REG_10__SCAN_IN), .ZN(n3176) );
  OR2_X1 U2476 ( .A1(n3195), .A2(n3194), .ZN(n3919) );
  NAND2_X1 U2477 ( .A1(n4426), .A2(n3925), .ZN(n3926) );
  NAND2_X1 U2478 ( .A1(n2206), .A2(n4472), .ZN(n3937) );
  INV_X1 U2479 ( .A(n2207), .ZN(n2206) );
  NOR2_X1 U2480 ( .A1(n3452), .A2(n2307), .ZN(n2306) );
  INV_X1 U2481 ( .A(n3442), .ZN(n2307) );
  AND2_X1 U2482 ( .A1(n3443), .A2(REG3_REG_27__SCAN_IN), .ZN(n3454) );
  AND2_X1 U2483 ( .A1(n3436), .A2(n3428), .ZN(n4033) );
  AOI22_X1 U2484 ( .A1(n4038), .A2(n3426), .B1(n3603), .B2(n3551), .ZN(n4021)
         );
  NAND2_X1 U2485 ( .A1(n3393), .A2(REG3_REG_20__SCAN_IN), .ZN(n3398) );
  INV_X1 U2486 ( .A(n2299), .ZN(n2298) );
  OAI21_X1 U2487 ( .B1(n3750), .B2(n2300), .A(n3748), .ZN(n2299) );
  OR2_X1 U2488 ( .A1(n4168), .A2(n2302), .ZN(n2300) );
  NAND2_X1 U2489 ( .A1(n2304), .A2(n4164), .ZN(n2303) );
  AOI21_X1 U2490 ( .B1(n4182), .B2(n3386), .A(n3385), .ZN(n4162) );
  OAI21_X1 U2491 ( .B1(n3508), .B2(n3641), .A(n3380), .ZN(n4182) );
  OR2_X1 U2492 ( .A1(n3316), .A2(n2325), .ZN(n2324) );
  NOR2_X1 U2493 ( .A1(n3875), .A2(n3256), .ZN(n2325) );
  NOR2_X1 U2494 ( .A1(n3235), .A2(n3779), .ZN(n3316) );
  NAND2_X1 U2495 ( .A1(n2315), .A2(n3103), .ZN(n3147) );
  NAND2_X1 U2496 ( .A1(n2862), .A2(n2319), .ZN(n2318) );
  NOR2_X1 U2497 ( .A1(n2927), .A2(n2320), .ZN(n2319) );
  AND2_X1 U2498 ( .A1(n2893), .A2(n2892), .ZN(n2951) );
  INV_X1 U2499 ( .A(n3886), .ZN(n2804) );
  INV_X1 U2500 ( .A(n2841), .ZN(n2188) );
  AND2_X1 U2501 ( .A1(n2536), .A2(n2519), .ZN(n2742) );
  NAND2_X1 U2502 ( .A1(n2518), .A2(n4468), .ZN(n2734) );
  AND2_X1 U2503 ( .A1(n3974), .A2(n3973), .ZN(n4212) );
  NAND2_X1 U2504 ( .A1(n3219), .A2(n4487), .ZN(n4508) );
  INV_X1 U2505 ( .A(n2404), .ZN(n2560) );
  AND2_X1 U2506 ( .A1(n2152), .A2(n2331), .ZN(n2330) );
  INV_X1 U2507 ( .A(IR_REG_25__SCAN_IN), .ZN(n2331) );
  NOR2_X1 U2508 ( .A1(n2397), .A2(IR_REG_21__SCAN_IN), .ZN(n2411) );
  XNOR2_X1 U2509 ( .A(n2383), .B(n2382), .ZN(n3859) );
  NAND2_X1 U2510 ( .A1(n2381), .A2(IR_REG_31__SCAN_IN), .ZN(n2383) );
  OR2_X1 U2511 ( .A1(n3318), .A2(IR_REG_14__SCAN_IN), .ZN(n3319) );
  NAND2_X1 U2512 ( .A1(n3679), .A2(n3547), .ZN(n3600) );
  AND2_X1 U2513 ( .A1(n3601), .A2(n3599), .ZN(n3547) );
  INV_X1 U2514 ( .A(n4335), .ZN(n3704) );
  NAND2_X1 U2515 ( .A1(n2219), .A2(n2216), .ZN(n2496) );
  NAND2_X1 U2516 ( .A1(n4359), .A2(REG1_REG_4__SCAN_IN), .ZN(n2220) );
  OAI21_X1 U2517 ( .B1(n4358), .B2(n2203), .A(n2200), .ZN(n2501) );
  AOI21_X1 U2518 ( .B1(n2469), .B2(n2202), .A(n2201), .ZN(n2200) );
  INV_X1 U2519 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2202) );
  OAI21_X1 U2520 ( .B1(n2479), .B2(n2198), .A(n2195), .ZN(n2511) );
  XNOR2_X1 U2521 ( .A(n2699), .B(n2895), .ZN(n2476) );
  NAND2_X1 U2522 ( .A1(n2476), .A2(REG2_REG_8__SCAN_IN), .ZN(n2700) );
  NAND2_X1 U2523 ( .A1(n4375), .A2(n4376), .ZN(n4374) );
  OR2_X1 U2524 ( .A1(n4356), .A2(n4314), .ZN(n4449) );
  AOI21_X1 U2525 ( .B1(n4435), .B2(n4434), .A(n4433), .ZN(n4440) );
  XNOR2_X1 U2526 ( .A(n2205), .B(n2180), .ZN(n2204) );
  OR2_X1 U2527 ( .A1(n4441), .A2(n2181), .ZN(n2205) );
  INV_X1 U2528 ( .A(n4398), .ZN(n4445) );
  NAND2_X1 U2529 ( .A1(n4435), .A2(n2156), .ZN(n2228) );
  NOR2_X1 U2530 ( .A1(n4212), .A2(n2185), .ZN(n4224) );
  NOR2_X1 U2531 ( .A1(n3974), .A2(n3973), .ZN(n2185) );
  NAND2_X1 U2532 ( .A1(n2308), .A2(n3453), .ZN(n3965) );
  NAND2_X1 U2533 ( .A1(n2312), .A2(n2311), .ZN(n2308) );
  NOR2_X1 U2534 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2340)
         );
  NOR2_X1 U2535 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2339)
         );
  NOR2_X1 U2536 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2350)
         );
  AOI21_X1 U2537 ( .B1(n3566), .B2(n3887), .A(n2649), .ZN(n2650) );
  AND2_X1 U2538 ( .A1(n3756), .A2(n4022), .ZN(n3846) );
  OR2_X1 U2539 ( .A1(n3890), .A2(n4527), .ZN(n2431) );
  NAND2_X1 U2540 ( .A1(n3905), .A2(n2463), .ZN(n2464) );
  INV_X1 U2541 ( .A(IR_REG_13__SCAN_IN), .ZN(n4738) );
  NOR2_X1 U2542 ( .A1(n4411), .A2(n3923), .ZN(n3924) );
  OR2_X1 U2543 ( .A1(n4416), .A2(n2208), .ZN(n2207) );
  AND2_X1 U2544 ( .A1(n3936), .A2(REG2_REG_15__SCAN_IN), .ZN(n2208) );
  AND2_X1 U2545 ( .A1(n3753), .A2(n4005), .ZN(n3853) );
  NOR2_X1 U2546 ( .A1(n3410), .A2(n4835), .ZN(n3419) );
  NOR2_X1 U2547 ( .A1(n4183), .A2(n3835), .ZN(n4059) );
  OAI21_X1 U2548 ( .B1(n3146), .B2(n2314), .A(n2175), .ZN(n2313) );
  OR2_X1 U2549 ( .A1(n3885), .A2(n2823), .ZN(n3798) );
  NAND2_X1 U2550 ( .A1(n2763), .A2(n2604), .ZN(n3792) );
  INV_X1 U2551 ( .A(IR_REG_18__SCAN_IN), .ZN(n2343) );
  NOR2_X1 U2552 ( .A1(n3381), .A2(IR_REG_17__SCAN_IN), .ZN(n3370) );
  INV_X1 U2553 ( .A(n2354), .ZN(n3381) );
  OAI21_X1 U2554 ( .B1(n3296), .B2(n3295), .A(n3294), .ZN(n3498) );
  INV_X1 U2555 ( .A(n2761), .ZN(n2803) );
  XNOR2_X1 U2556 ( .A(n2548), .B(n3571), .ZN(n2642) );
  INV_X1 U2557 ( .A(n3553), .ZN(n2289) );
  AOI21_X1 U2558 ( .B1(n2273), .B2(n2155), .A(n2174), .ZN(n2271) );
  INV_X1 U2559 ( .A(n3510), .ZN(n2275) );
  INV_X1 U2560 ( .A(n2273), .ZN(n2272) );
  OR2_X1 U2561 ( .A1(n3531), .A2(n2525), .ZN(n2531) );
  AOI22_X1 U2562 ( .A1(n2529), .A2(IR_REG_0__SCAN_IN), .B1(n3561), .B2(n2188), 
        .ZN(n2530) );
  AOI21_X1 U2563 ( .B1(n2261), .B2(n2260), .A(n2259), .ZN(n2258) );
  INV_X1 U2564 ( .A(n3671), .ZN(n2259) );
  INV_X1 U2565 ( .A(n2264), .ZN(n2260) );
  NAND2_X1 U2566 ( .A1(n3087), .A2(REG3_REG_12__SCAN_IN), .ZN(n3129) );
  NAND2_X1 U2567 ( .A1(n2415), .A2(n2153), .ZN(n2192) );
  NAND2_X1 U2568 ( .A1(n2640), .A2(n2641), .ZN(n2242) );
  OR2_X1 U2569 ( .A1(n2650), .A2(n2651), .ZN(n2241) );
  NAND2_X1 U2570 ( .A1(n3511), .A2(n3510), .ZN(n3700) );
  AOI22_X1 U2571 ( .A1(n3901), .A2(n3900), .B1(n4324), .B2(REG1_REG_2__SCAN_IN), .ZN(n2433) );
  XNOR2_X1 U2572 ( .A(n2464), .B(n2493), .ZN(n2488) );
  NOR2_X1 U2573 ( .A1(n2497), .A2(n2222), .ZN(n2221) );
  NAND2_X1 U2574 ( .A1(n2218), .A2(n2217), .ZN(n2216) );
  INV_X1 U2575 ( .A(n2497), .ZN(n2217) );
  INV_X1 U2576 ( .A(n2224), .ZN(n2218) );
  INV_X1 U2577 ( .A(n2503), .ZN(n2201) );
  NAND2_X1 U2578 ( .A1(n2501), .A2(n2470), .ZN(n2471) );
  NOR2_X1 U2579 ( .A1(n2363), .A2(n2328), .ZN(n2439) );
  INV_X1 U2580 ( .A(IR_REG_7__SCAN_IN), .ZN(n2441) );
  NAND2_X1 U2581 ( .A1(n2227), .A2(REG1_REG_8__SCAN_IN), .ZN(n2226) );
  OR2_X1 U2582 ( .A1(n3186), .A2(n3187), .ZN(n2213) );
  XNOR2_X1 U2583 ( .A(n3190), .B(n4474), .ZN(n4390) );
  NOR2_X1 U2584 ( .A1(n4390), .A2(n4633), .ZN(n4389) );
  NOR2_X1 U2585 ( .A1(n3168), .A2(n3167), .ZN(n3171) );
  INV_X1 U2586 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3184) );
  NAND2_X1 U2587 ( .A1(n3919), .A2(n2238), .ZN(n2240) );
  NOR2_X1 U2588 ( .A1(n2239), .A2(n4406), .ZN(n2238) );
  INV_X1 U2589 ( .A(n3918), .ZN(n2239) );
  AND2_X1 U2590 ( .A1(n3920), .A2(n4406), .ZN(n3921) );
  NOR2_X1 U2591 ( .A1(n3933), .A2(n3934), .ZN(n3935) );
  NOR2_X1 U2592 ( .A1(n4401), .A2(n3921), .ZN(n4413) );
  NOR2_X1 U2593 ( .A1(n4413), .A2(n4412), .ZN(n4411) );
  NAND2_X1 U2594 ( .A1(n4427), .A2(n4774), .ZN(n4426) );
  INV_X1 U2595 ( .A(n2310), .ZN(n2309) );
  OAI21_X1 U2596 ( .B1(n3452), .B2(n2311), .A(n3964), .ZN(n2310) );
  AND2_X1 U2597 ( .A1(n3451), .A2(n2172), .ZN(n2311) );
  NAND2_X1 U2598 ( .A1(n4013), .A2(n3450), .ZN(n3451) );
  AND2_X1 U2599 ( .A1(n4109), .A2(n4127), .ZN(n4090) );
  NOR2_X1 U2600 ( .A1(n3373), .A2(n4333), .ZN(n3387) );
  OR3_X1 U2601 ( .A1(n3355), .A2(n3354), .A3(n3353), .ZN(n3373) );
  AND2_X1 U2602 ( .A1(n3343), .A2(n3707), .ZN(n3344) );
  NAND2_X1 U2603 ( .A1(n3874), .A2(n3335), .ZN(n2323) );
  AND2_X1 U2604 ( .A1(n3640), .A2(n3707), .ZN(n3336) );
  NAND2_X1 U2605 ( .A1(n3247), .A2(REG3_REG_15__SCAN_IN), .ZN(n3355) );
  INV_X1 U2606 ( .A(n3246), .ZN(n3779) );
  AND2_X1 U2607 ( .A1(n3241), .A2(n3238), .ZN(n3778) );
  OR2_X1 U2608 ( .A1(n3041), .A2(n3815), .ZN(n3042) );
  OR2_X1 U2609 ( .A1(n2903), .A2(n2902), .ZN(n2937) );
  AND2_X1 U2610 ( .A1(n2679), .A2(n2678), .ZN(n2867) );
  NOR2_X1 U2611 ( .A1(n2720), .A2(n2719), .ZN(n2786) );
  NAND2_X1 U2612 ( .A1(n2676), .A2(REG3_REG_5__SCAN_IN), .ZN(n2720) );
  INV_X1 U2613 ( .A(n2857), .ZN(n2860) );
  AND2_X1 U2614 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2676) );
  INV_X1 U2615 ( .A(n4188), .ZN(n4172) );
  NAND2_X1 U2616 ( .A1(n3792), .A2(n3795), .ZN(n2615) );
  AND2_X1 U2617 ( .A1(n2621), .A2(n4314), .ZN(n4188) );
  OR2_X1 U2618 ( .A1(n4314), .A2(n2614), .ZN(n4185) );
  AND2_X1 U2619 ( .A1(n2598), .A2(n2188), .ZN(n2843) );
  AND2_X1 U2620 ( .A1(n2619), .A2(n3863), .ZN(n4190) );
  INV_X1 U2621 ( .A(n4185), .ZN(n4169) );
  AND2_X1 U2622 ( .A1(n2630), .A2(n2627), .ZN(n2737) );
  INV_X1 U2623 ( .A(n4217), .ZN(n4207) );
  AND2_X1 U2624 ( .A1(n2742), .A2(n2618), .ZN(n4217) );
  NAND2_X1 U2625 ( .A1(n4030), .A2(n4015), .ZN(n4014) );
  NOR2_X1 U2626 ( .A1(n4072), .A2(n4050), .ZN(n4049) );
  INV_X1 U2627 ( .A(n3551), .ZN(n4050) );
  INV_X1 U2628 ( .A(n3200), .ZN(n3201) );
  AND2_X1 U2629 ( .A1(n3111), .A2(n3145), .ZN(n3139) );
  OR2_X1 U2630 ( .A1(n2966), .A2(n3047), .ZN(n3062) );
  INV_X1 U2632 ( .A(n3098), .ZN(n3099) );
  NAND2_X1 U2634 ( .A1(n2964), .A2(n2963), .ZN(n2966) );
  NAND2_X1 U2635 ( .A1(n2189), .A2(n2863), .ZN(n2921) );
  AND2_X1 U2636 ( .A1(n2744), .A2(n2536), .ZN(n4521) );
  INV_X1 U2637 ( .A(n2636), .ZN(n2738) );
  AND3_X1 U2638 ( .A1(n2632), .A2(n2631), .A3(n2630), .ZN(n2637) );
  INV_X1 U2639 ( .A(n4521), .ZN(n4487) );
  OAI21_X1 U2640 ( .B1(n2392), .B2(n2336), .A(n2391), .ZN(n2420) );
  AND2_X1 U2641 ( .A1(n2389), .A2(IR_REG_29__SCAN_IN), .ZN(n2392) );
  AND2_X1 U2642 ( .A1(n2332), .A2(n2417), .ZN(n2329) );
  XNOR2_X1 U2643 ( .A(n2362), .B(n2346), .ZN(n2671) );
  NAND2_X1 U2644 ( .A1(n2397), .A2(IR_REG_31__SCAN_IN), .ZN(n2399) );
  AND2_X1 U2645 ( .A1(n3070), .A2(n3127), .ZN(n3188) );
  INV_X1 U2646 ( .A(IR_REG_3__SCAN_IN), .ZN(n2372) );
  CLKBUF_X1 U2647 ( .A(n2370), .Z(n2371) );
  XNOR2_X1 U2648 ( .A(n2428), .B(n2427), .ZN(n3902) );
  NOR2_X1 U2649 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2426)
         );
  XNOR2_X1 U2650 ( .A(n2214), .B(IR_REG_1__SCAN_IN), .ZN(n3890) );
  AND2_X1 U2651 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2214)
         );
  AOI21_X1 U2652 ( .B1(n2154), .B2(n2281), .A(n2173), .ZN(n2279) );
  INV_X1 U2653 ( .A(n4066), .ZN(n4073) );
  NAND2_X1 U2654 ( .A1(n2975), .A2(n2977), .ZN(n2246) );
  AND2_X1 U2655 ( .A1(n3468), .A2(n3467), .ZN(n3737) );
  AND2_X1 U2656 ( .A1(n3953), .A2(n3455), .ZN(n3980) );
  AND3_X1 U2657 ( .A1(n3397), .A2(n3396), .A3(n3395), .ZN(n4139) );
  INV_X1 U2658 ( .A(n2284), .ZN(n3630) );
  OAI21_X1 U2659 ( .B1(n3600), .B2(n2171), .A(n2286), .ZN(n2284) );
  NAND2_X1 U2660 ( .A1(n2716), .A2(n2715), .ZN(n2773) );
  NAND2_X1 U2661 ( .A1(n2270), .A2(n2271), .ZN(n3650) );
  OR2_X1 U2662 ( .A1(n3511), .A2(n2272), .ZN(n2270) );
  AOI21_X1 U2663 ( .B1(n3600), .B2(n3554), .A(n3553), .ZN(n3656) );
  NAND2_X1 U2664 ( .A1(n2686), .A2(n2668), .ZN(n2716) );
  INV_X1 U2665 ( .A(n3047), .ZN(n3055) );
  NAND2_X1 U2666 ( .A1(n2248), .A2(n2975), .ZN(n2249) );
  OR2_X1 U2667 ( .A1(n2976), .A2(n2977), .ZN(n2248) );
  NAND2_X1 U2668 ( .A1(n2653), .A2(IR_REG_0__SCAN_IN), .ZN(n2528) );
  NAND2_X1 U2669 ( .A1(n2257), .A2(n2261), .ZN(n3670) );
  NAND2_X1 U2670 ( .A1(n2150), .A2(n2264), .ZN(n2257) );
  NAND2_X1 U2671 ( .A1(n2241), .A2(n2652), .ZN(n2751) );
  INV_X1 U2672 ( .A(n3683), .ZN(n4327) );
  OR2_X1 U2673 ( .A1(n2585), .A2(n2579), .ZN(n4335) );
  INV_X1 U2674 ( .A(n3712), .ZN(n4337) );
  OAI21_X1 U2675 ( .B1(n2686), .B2(n2256), .A(n2254), .ZN(n2887) );
  INV_X1 U2676 ( .A(n2255), .ZN(n2254) );
  OAI21_X1 U2677 ( .B1(n3600), .B2(n2283), .A(n2281), .ZN(n3691) );
  INV_X1 U2678 ( .A(n4342), .ZN(n3710) );
  NAND2_X1 U2679 ( .A1(n3433), .A2(n3432), .ZN(n4045) );
  NAND2_X1 U2680 ( .A1(n3425), .A2(n3424), .ZN(n4068) );
  INV_X1 U2681 ( .A(n4085), .ZN(n4044) );
  INV_X1 U2682 ( .A(n4139), .ZN(n4100) );
  INV_X1 U2683 ( .A(n4173), .ZN(n4326) );
  INV_X1 U2684 ( .A(n2951), .ZN(n3881) );
  NAND4_X1 U2685 ( .A1(n2791), .A2(n2790), .A3(n2789), .A4(n2788), .ZN(n3882)
         );
  INV_X1 U2686 ( .A(n2867), .ZN(n3884) );
  OR2_X1 U2687 ( .A1(n2609), .A2(n2768), .ZN(n2610) );
  CLKBUF_X1 U2688 ( .A(n2597), .Z(n3888) );
  INV_X1 U2689 ( .A(n4323), .ZN(n2493) );
  NAND2_X1 U2690 ( .A1(n4358), .A2(REG2_REG_4__SCAN_IN), .ZN(n2199) );
  XNOR2_X1 U2691 ( .A(n2471), .B(n2482), .ZN(n2479) );
  NAND2_X1 U2692 ( .A1(n2700), .A2(n2701), .ZN(n4375) );
  AND2_X1 U2693 ( .A1(n2225), .A2(n2226), .ZN(n4371) );
  NOR2_X1 U2694 ( .A1(n2709), .A2(n3124), .ZN(n3186) );
  NAND2_X1 U2695 ( .A1(n3176), .A2(n3177), .ZN(n4385) );
  NAND2_X1 U2696 ( .A1(n4385), .A2(n4386), .ZN(n4384) );
  AND2_X1 U2697 ( .A1(n2213), .A2(n2212), .ZN(n4379) );
  INV_X1 U2698 ( .A(n4380), .ZN(n2212) );
  INV_X1 U2699 ( .A(n2213), .ZN(n4381) );
  NOR2_X1 U2700 ( .A1(n3921), .A2(n2237), .ZN(n4401) );
  NAND2_X1 U2701 ( .A1(n2240), .A2(REG1_REG_14__SCAN_IN), .ZN(n2237) );
  NAND2_X1 U2702 ( .A1(n2236), .A2(n2240), .ZN(n4403) );
  INV_X1 U2703 ( .A(n3921), .ZN(n2236) );
  NOR2_X1 U2704 ( .A1(n4400), .A2(n4641), .ZN(n4399) );
  NAND2_X1 U2705 ( .A1(n2211), .A2(n2210), .ZN(n4400) );
  NAND2_X1 U2706 ( .A1(n3933), .A2(n3934), .ZN(n2210) );
  INV_X1 U2707 ( .A(n3935), .ZN(n2211) );
  AOI22_X1 U2708 ( .A1(n2232), .A2(n4434), .B1(n3945), .B2(n2179), .ZN(n2231)
         );
  OR2_X1 U2709 ( .A1(n4434), .A2(n2235), .ZN(n2234) );
  INV_X1 U2710 ( .A(n3945), .ZN(n2235) );
  OR2_X1 U2711 ( .A1(n3454), .A2(n3444), .ZN(n3999) );
  XOR2_X1 U2712 ( .A(n4007), .B(n4004), .Z(n4230) );
  NAND2_X1 U2713 ( .A1(n4090), .A2(n4091), .ZN(n4243) );
  NAND2_X1 U2714 ( .A1(n2295), .A2(n2298), .ZN(n4116) );
  NAND2_X1 U2715 ( .A1(n2297), .A2(n2296), .ZN(n2295) );
  NAND2_X1 U2716 ( .A1(n4161), .A2(n2303), .ZN(n4137) );
  INV_X1 U2717 ( .A(n2324), .ZN(n3334) );
  NAND2_X1 U2718 ( .A1(n3147), .A2(n3146), .ZN(n3203) );
  NOR2_X1 U2719 ( .A1(n2321), .A2(n2317), .ZN(n2316) );
  INV_X1 U2720 ( .A(n2322), .ZN(n2317) );
  AND2_X1 U2721 ( .A1(n4350), .A2(n3950), .ZN(n4179) );
  NAND2_X1 U2722 ( .A1(n2318), .A2(n2322), .ZN(n2929) );
  AND2_X1 U2723 ( .A1(n4350), .A2(n2818), .ZN(n4107) );
  AND2_X1 U2724 ( .A1(n4179), .A2(n4510), .ZN(n4461) );
  AND2_X1 U2725 ( .A1(n4350), .A2(n2741), .ZN(n4459) );
  INV_X1 U2726 ( .A(n4461), .ZN(n4195) );
  OR2_X1 U2727 ( .A1(n2734), .A2(n2628), .ZN(n4197) );
  NAND2_X1 U2728 ( .A1(n2188), .A2(n2742), .ZN(n4478) );
  INV_X1 U2729 ( .A(n4197), .ZN(n4457) );
  AND2_X2 U2730 ( .A1(n2637), .A2(n2636), .ZN(n4537) );
  INV_X1 U2731 ( .A(n4537), .ZN(n4534) );
  AND2_X1 U2732 ( .A1(n4214), .A2(n4213), .ZN(n4348) );
  NAND2_X1 U2733 ( .A1(n2184), .A2(n2183), .ZN(n4280) );
  NAND2_X1 U2734 ( .A1(n4224), .A2(n4510), .ZN(n2184) );
  NOR2_X1 U2735 ( .A1(n4223), .A2(n2165), .ZN(n2183) );
  AND2_X2 U2736 ( .A1(n2637), .A2(n2738), .ZN(n4524) );
  NAND2_X1 U2737 ( .A1(n2564), .A2(n2575), .ZN(n4467) );
  NAND2_X1 U2738 ( .A1(n2391), .A2(IR_REG_31__SCAN_IN), .ZN(n2387) );
  XNOR2_X1 U2739 ( .A(n2355), .B(IR_REG_26__SCAN_IN), .ZN(n2404) );
  NAND2_X1 U2740 ( .A1(n2348), .A2(IR_REG_31__SCAN_IN), .ZN(n2349) );
  INV_X1 U2741 ( .A(n2536), .ZN(n4315) );
  INV_X1 U2742 ( .A(n2519), .ZN(n2517) );
  XNOR2_X1 U2743 ( .A(n2535), .B(IR_REG_19__SCAN_IN), .ZN(n4316) );
  XNOR2_X1 U2744 ( .A(n3341), .B(n3340), .ZN(n4472) );
  INV_X1 U2745 ( .A(n3188), .ZN(n4475) );
  NAND2_X1 U2746 ( .A1(n2199), .A2(n2469), .ZN(n2502) );
  AOI21_X1 U2747 ( .B1(n2161), .B2(n4440), .A(n4439), .ZN(n4447) );
  AOI21_X1 U2748 ( .B1(n2204), .B2(n4445), .A(n3951), .ZN(n3952) );
  NAND2_X1 U2749 ( .A1(n2234), .A2(n2231), .ZN(n2230) );
  MUX2_X1 U2750 ( .A(n3484), .B(n3489), .S(n4537), .Z(n3488) );
  MUX2_X1 U2751 ( .A(n4804), .B(n3489), .S(n4524), .Z(n3491) );
  INV_X2 U2752 ( .A(n2572), .ZN(n3561) );
  AND2_X1 U2753 ( .A1(n2266), .A2(n2267), .ZN(n2150) );
  AND2_X1 U2754 ( .A1(n2298), .A2(n2177), .ZN(n2151) );
  OAI21_X1 U2755 ( .B1(n3999), .B2(n3462), .A(n3449), .ZN(n3873) );
  AND4_X1 U2756 ( .A1(n2353), .A2(n2352), .A3(n2351), .A4(n2350), .ZN(n2152)
         );
  AND2_X1 U2757 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2153)
         );
  NOR2_X2 U2758 ( .A1(n2157), .A2(n3966), .ZN(n3974) );
  AND2_X1 U2759 ( .A1(n2283), .A2(n2280), .ZN(n2154) );
  INV_X1 U2760 ( .A(n4150), .ZN(n2304) );
  AND2_X1 U2761 ( .A1(n2275), .A2(n3701), .ZN(n2155) );
  NAND2_X1 U2762 ( .A1(n2242), .A2(n2645), .ZN(n2748) );
  AND2_X1 U2763 ( .A1(n2231), .A2(n2233), .ZN(n2156) );
  OR2_X1 U2764 ( .A1(n4014), .A2(n3996), .ZN(n2157) );
  AND2_X1 U2765 ( .A1(n3797), .A2(n3794), .ZN(n2158) );
  INV_X1 U2766 ( .A(IR_REG_31__SCAN_IN), .ZN(n3170) );
  XNOR2_X1 U2767 ( .A(n2399), .B(n2398), .ZN(n2519) );
  INV_X1 U2768 ( .A(IR_REG_0__SCAN_IN), .ZN(n4547) );
  AOI22_X1 U2769 ( .A1(n4021), .A2(n3435), .B1(n2190), .B2(n4045), .ZN(n4004)
         );
  AND2_X1 U2770 ( .A1(n2291), .A2(n2420), .ZN(n2159) );
  AND2_X1 U2771 ( .A1(n3554), .A2(n3553), .ZN(n2160) );
  OR2_X1 U2772 ( .A1(n4435), .A2(n4434), .ZN(n2161) );
  OR2_X1 U2773 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2162) );
  OR2_X1 U2774 ( .A1(IR_REG_26__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2163)
         );
  INV_X1 U2775 ( .A(n3452), .ZN(n3453) );
  NOR2_X1 U2776 ( .A1(n2363), .A2(IR_REG_5__SCAN_IN), .ZN(n2365) );
  INV_X1 U2777 ( .A(n2420), .ZN(n2520) );
  NAND4_X1 U2778 ( .A1(n2547), .A2(n2546), .A3(n2545), .A4(n2544), .ZN(n2597)
         );
  INV_X1 U2779 ( .A(n2287), .ZN(n2286) );
  OAI22_X1 U2780 ( .A1(n2160), .A2(n2288), .B1(n3553), .B2(n3554), .ZN(n2287)
         );
  AND2_X1 U2781 ( .A1(n3103), .A2(n3202), .ZN(n2164) );
  AND2_X1 U2782 ( .A1(n4222), .A2(n4508), .ZN(n2165) );
  AND2_X1 U2783 ( .A1(n3600), .A2(n2160), .ZN(n2166) );
  INV_X1 U2784 ( .A(n2301), .ZN(n2296) );
  OR2_X1 U2785 ( .A1(n3750), .A2(n2302), .ZN(n2301) );
  AND4_X1 U2786 ( .A1(n2342), .A2(n2341), .A3(n2340), .A4(n2339), .ZN(n2167)
         );
  NAND2_X1 U2787 ( .A1(n2401), .A2(n2360), .ZN(n2518) );
  AND2_X1 U2788 ( .A1(n2281), .A2(n2280), .ZN(n2168) );
  INV_X1 U2789 ( .A(n2262), .ZN(n2261) );
  OAI22_X1 U2790 ( .A1(n3609), .A2(n2263), .B1(n3528), .B2(n3529), .ZN(n2262)
         );
  NAND2_X1 U2791 ( .A1(n3880), .A2(n3047), .ZN(n2169) );
  INV_X1 U2792 ( .A(n2715), .ZN(n2256) );
  OR2_X1 U2793 ( .A1(n2717), .A2(n4606), .ZN(n2170) );
  NAND2_X1 U2794 ( .A1(n2290), .A2(n2520), .ZN(n2542) );
  XNOR2_X1 U2795 ( .A(n2349), .B(IR_REG_24__SCAN_IN), .ZN(n2401) );
  CLKBUF_X3 U2796 ( .A(n2607), .Z(n3412) );
  NOR2_X1 U2797 ( .A1(n3657), .A2(n2289), .ZN(n2171) );
  NAND2_X1 U2798 ( .A1(n2326), .A2(n2327), .ZN(n2696) );
  AOI21_X1 U2799 ( .B1(n2150), .B2(n4330), .A(n4331), .ZN(n3608) );
  OR2_X1 U2800 ( .A1(n4026), .A2(n4010), .ZN(n2172) );
  INV_X1 U2801 ( .A(n3701), .ZN(n2276) );
  NAND2_X1 U2802 ( .A1(n4162), .A2(n4168), .ZN(n4161) );
  AND2_X1 U2803 ( .A1(n3568), .A2(n3567), .ZN(n2173) );
  INV_X1 U2804 ( .A(n4322), .ZN(n2482) );
  INV_X1 U2805 ( .A(n4164), .ZN(n4328) );
  NOR2_X1 U2806 ( .A1(n3513), .A2(n3512), .ZN(n2174) );
  NAND2_X1 U2807 ( .A1(n3215), .A2(n3201), .ZN(n2175) );
  INV_X1 U2808 ( .A(n2277), .ZN(n3699) );
  OR2_X1 U2809 ( .A1(n3511), .A2(n3510), .ZN(n2277) );
  INV_X1 U2810 ( .A(n3970), .ZN(n3971) );
  AND2_X1 U2811 ( .A1(n3518), .A2(n3517), .ZN(n2176) );
  NAND2_X1 U2812 ( .A1(n4100), .A2(n4122), .ZN(n2177) );
  INV_X1 U2814 ( .A(n3773), .ZN(n2321) );
  XNOR2_X1 U2815 ( .A(n2413), .B(n2412), .ZN(n2536) );
  INV_X1 U2816 ( .A(n4330), .ZN(n2265) );
  NAND2_X1 U2817 ( .A1(n2249), .A2(n2982), .ZN(n2983) );
  INV_X1 U2818 ( .A(n2193), .ZN(n3257) );
  NOR2_X1 U2819 ( .A1(n3221), .A2(n3243), .ZN(n2193) );
  AND2_X1 U2820 ( .A1(n3188), .A2(REG1_REG_11__SCAN_IN), .ZN(n2178) );
  INV_X1 U2821 ( .A(n4032), .ZN(n2190) );
  AND2_X1 U2822 ( .A1(n4469), .A2(REG1_REG_18__SCAN_IN), .ZN(n2179) );
  OR2_X1 U2823 ( .A1(n4356), .A2(n4353), .ZN(n4433) );
  OR2_X1 U2824 ( .A1(n2836), .A2(n2860), .ZN(n2871) );
  INV_X1 U2825 ( .A(n2871), .ZN(n2189) );
  INV_X1 U2826 ( .A(n2233), .ZN(n2232) );
  OR2_X1 U2827 ( .A1(n3945), .A2(n2179), .ZN(n2233) );
  INV_X1 U2828 ( .A(n4319), .ZN(n2209) );
  INV_X1 U2829 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2222) );
  INV_X1 U2830 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2197) );
  XOR2_X1 U2831 ( .A(n3950), .B(REG2_REG_19__SCAN_IN), .Z(n2180) );
  AND2_X1 U2832 ( .A1(n4469), .A2(REG2_REG_18__SCAN_IN), .ZN(n2181) );
  AND2_X1 U2833 ( .A1(n2220), .A2(n2224), .ZN(n2182) );
  NAND2_X1 U2835 ( .A1(n2415), .A2(IR_REG_31__SCAN_IN), .ZN(n2449) );
  NAND2_X1 U2837 ( .A1(n2416), .A2(n2192), .ZN(n2191) );
  NOR2_X1 U2838 ( .A1(n4153), .A2(n4152), .ZN(n4154) );
  AND3_X2 U2841 ( .A1(n2326), .A2(n2167), .A3(n2327), .ZN(n2354) );
  NAND2_X1 U2842 ( .A1(n3344), .A2(n3641), .ZN(n3486) );
  NAND2_X1 U2843 ( .A1(n2194), .A2(n2472), .ZN(n2512) );
  NAND2_X1 U2844 ( .A1(n2479), .A2(REG2_REG_6__SCAN_IN), .ZN(n2194) );
  AOI21_X1 U2845 ( .B1(n2472), .B2(n2197), .A(n2196), .ZN(n2195) );
  INV_X1 U2846 ( .A(n2474), .ZN(n2196) );
  INV_X1 U2847 ( .A(n2472), .ZN(n2198) );
  INV_X1 U2848 ( .A(n2469), .ZN(n2203) );
  OAI22_X1 U2849 ( .A1(n3932), .A2(n3931), .B1(n4318), .B2(
        REG2_REG_13__SCAN_IN), .ZN(n3933) );
  NAND2_X1 U2850 ( .A1(n3178), .A2(n4384), .ZN(n3179) );
  NAND2_X1 U2851 ( .A1(n4425), .A2(n3348), .ZN(n4424) );
  NAND2_X1 U2856 ( .A1(n4359), .A2(n2221), .ZN(n2219) );
  XNOR2_X1 U2857 ( .A(n2223), .B(n4322), .ZN(n2480) );
  NAND3_X1 U2858 ( .A1(n2216), .A2(n2170), .A3(n2219), .ZN(n2223) );
  INV_X1 U2859 ( .A(n2223), .ZN(n2437) );
  NAND2_X1 U2860 ( .A1(n2435), .A2(n2467), .ZN(n2224) );
  INV_X1 U2861 ( .A(n2706), .ZN(n2225) );
  NOR2_X1 U2862 ( .A1(n2706), .A2(n2226), .ZN(n2705) );
  NAND2_X1 U2863 ( .A1(n2225), .A2(n2227), .ZN(n2450) );
  NAND2_X1 U2864 ( .A1(n2446), .A2(n2895), .ZN(n2227) );
  OAI211_X1 U2865 ( .C1(n4435), .C2(n2230), .A(n4429), .B(n2228), .ZN(n2229)
         );
  NAND2_X1 U2866 ( .A1(n3952), .A2(n2229), .ZN(U3259) );
  NAND2_X1 U2867 ( .A1(n3919), .A2(n3918), .ZN(n3920) );
  NAND4_X1 U2868 ( .A1(n2242), .A2(n2645), .A3(n2652), .A4(n2241), .ZN(n2749)
         );
  OAI22_X1 U2869 ( .A1(n2572), .A2(n2596), .B1(n2846), .B2(n3577), .ZN(n2548)
         );
  NAND2_X4 U2870 ( .A1(n2518), .A2(n2740), .ZN(n3577) );
  NAND2_X2 U2871 ( .A1(n2518), .A2(n2526), .ZN(n2572) );
  INV_X1 U2872 ( .A(IR_REG_0__SCAN_IN), .ZN(n2244) );
  INV_X1 U2873 ( .A(IR_REG_1__SCAN_IN), .ZN(n2243) );
  NAND3_X1 U2874 ( .A1(n2427), .A2(n2244), .A3(n2243), .ZN(n2370) );
  INV_X2 U2875 ( .A(IR_REG_2__SCAN_IN), .ZN(n2427) );
  NAND2_X1 U2876 ( .A1(n2247), .A2(n2245), .ZN(n3025) );
  NAND2_X1 U2877 ( .A1(n2976), .A2(n2975), .ZN(n2247) );
  INV_X1 U2878 ( .A(n2668), .ZN(n2252) );
  NAND2_X1 U2879 ( .A1(n2255), .A2(n2886), .ZN(n2250) );
  NAND2_X1 U2880 ( .A1(n2252), .A2(n2715), .ZN(n2251) );
  NAND2_X1 U2881 ( .A1(n2886), .A2(n2715), .ZN(n2253) );
  OAI21_X1 U2882 ( .B1(n2150), .B2(n2262), .A(n2258), .ZN(n3669) );
  NAND2_X1 U2883 ( .A1(n3511), .A2(n2268), .ZN(n2266) );
  NAND2_X1 U2884 ( .A1(n3600), .A2(n2168), .ZN(n2278) );
  NAND2_X1 U2885 ( .A1(n2278), .A2(n2279), .ZN(n3591) );
  AND2_X1 U2886 ( .A1(n2520), .A2(n2291), .ZN(n2607) );
  NOR2_X1 U2887 ( .A1(n2520), .A2(n2291), .ZN(n2543) );
  NAND2_X1 U2888 ( .A1(n2291), .A2(STATE_REG_SCAN_IN), .ZN(n2388) );
  NAND2_X1 U2889 ( .A1(n4162), .A2(n2151), .ZN(n2292) );
  NAND2_X1 U2890 ( .A1(n2292), .A2(n2293), .ZN(n4105) );
  NAND2_X1 U2891 ( .A1(n4004), .A2(n3442), .ZN(n2312) );
  NAND2_X1 U2892 ( .A1(n2305), .A2(n2309), .ZN(n3969) );
  NAND2_X1 U2893 ( .A1(n4004), .A2(n2306), .ZN(n2305) );
  AND2_X1 U2894 ( .A1(n2312), .A2(n2172), .ZN(n3995) );
  AOI21_X2 U2895 ( .B1(n2315), .B2(n2164), .A(n2313), .ZN(n3232) );
  INV_X1 U2896 ( .A(n3104), .ZN(n2315) );
  NAND2_X1 U2897 ( .A1(n2318), .A2(n2316), .ZN(n3051) );
  NAND2_X1 U2898 ( .A1(n2862), .A2(n2861), .ZN(n2928) );
  INV_X1 U2899 ( .A(n2861), .ZN(n2320) );
  OR2_X1 U2900 ( .A1(n3883), .A2(n2926), .ZN(n2322) );
  AOI21_X2 U2901 ( .B1(n2324), .B2(n2323), .A(n3336), .ZN(n3342) );
  AND2_X1 U2903 ( .A1(n2354), .A2(n2332), .ZN(n2451) );
  NAND2_X1 U2904 ( .A1(n2354), .A2(n2329), .ZN(n2453) );
  NAND2_X1 U2905 ( .A1(n2354), .A2(n2152), .ZN(n2356) );
  OR2_X1 U2906 ( .A1(n2411), .A2(n3170), .ZN(n2413) );
  NAND2_X1 U2907 ( .A1(n2449), .A2(n2417), .ZN(n2416) );
  OAI22_X1 U2908 ( .A1(n2596), .A2(n3531), .B1(n2846), .B2(n3576), .ZN(n2643)
         );
  AND2_X1 U2909 ( .A1(n4862), .A2(DATAI_23_), .ZN(n4066) );
  NAND2_X1 U2910 ( .A1(n4862), .A2(DATAI_20_), .ZN(n4129) );
  OR2_X1 U2911 ( .A1(n3734), .A2(n4324), .ZN(n2603) );
  INV_X1 U2912 ( .A(n3734), .ZN(n2653) );
  AND2_X1 U2913 ( .A1(n2522), .A2(n2521), .ZN(n2334) );
  AND2_X1 U2914 ( .A1(n2374), .A2(n2372), .ZN(n2335) );
  AND2_X1 U2915 ( .A1(IR_REG_31__SCAN_IN), .A2(n2390), .ZN(n2336) );
  INV_X1 U2916 ( .A(n2757), .ZN(n2604) );
  AND2_X1 U2917 ( .A1(n4862), .A2(DATAI_27_), .ZN(n3996) );
  INV_X1 U2918 ( .A(n3996), .ZN(n3450) );
  NAND2_X1 U2919 ( .A1(n4862), .A2(DATAI_22_), .ZN(n4091) );
  INV_X1 U2920 ( .A(n3243), .ZN(n3230) );
  AND2_X1 U2921 ( .A1(n2581), .A2(n2580), .ZN(n2337) );
  AND2_X1 U2922 ( .A1(n3647), .A2(n3648), .ZN(n3516) );
  INV_X1 U2923 ( .A(n3876), .ZN(n3229) );
  NOR2_X1 U2924 ( .A1(n4013), .A2(n3450), .ZN(n3452) );
  INV_X1 U2925 ( .A(IR_REG_29__SCAN_IN), .ZN(n2390) );
  OR2_X1 U2926 ( .A1(n3577), .A2(n2803), .ZN(n2654) );
  NOR2_X1 U2927 ( .A1(n2560), .A2(n2408), .ZN(n2360) );
  AND2_X1 U2928 ( .A1(n3936), .A2(REG1_REG_15__SCAN_IN), .ZN(n3923) );
  INV_X1 U2929 ( .A(n4091), .ZN(n3408) );
  NAND2_X1 U2930 ( .A1(n3967), .A2(n3966), .ZN(n3968) );
  INV_X1 U2931 ( .A(n3778), .ZN(n3103) );
  NOR2_X1 U2932 ( .A1(n2890), .A2(n3012), .ZN(n3008) );
  INV_X1 U2933 ( .A(n2986), .ZN(n2984) );
  NAND2_X1 U2934 ( .A1(n3734), .A2(n2601), .ZN(n2602) );
  NAND2_X1 U2935 ( .A1(n2782), .A2(n2781), .ZN(n3007) );
  OR2_X1 U2936 ( .A1(n3427), .A2(n4576), .ZN(n3436) );
  INV_X1 U2937 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4831) );
  OR2_X1 U2938 ( .A1(n3954), .A2(n3461), .ZN(n3964) );
  NAND2_X1 U2939 ( .A1(n4067), .A2(n3408), .ZN(n3409) );
  AND2_X1 U2940 ( .A1(n3485), .A2(n4326), .ZN(n3385) );
  INV_X1 U2941 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2719) );
  INV_X1 U2942 ( .A(n2401), .ZN(n2561) );
  INV_X1 U2943 ( .A(n3004), .ZN(n2950) );
  INV_X1 U2944 ( .A(IR_REG_22__SCAN_IN), .ZN(n2412) );
  INV_X1 U2945 ( .A(n4068), .ZN(n3603) );
  NOR2_X1 U2946 ( .A1(n2937), .A2(n4831), .ZN(n3029) );
  NAND2_X1 U2947 ( .A1(n3734), .A2(DATAI_0_), .ZN(n2527) );
  OR2_X1 U2948 ( .A1(n3129), .A2(n3184), .ZN(n3208) );
  AND2_X1 U2949 ( .A1(n3029), .A2(REG3_REG_11__SCAN_IN), .ZN(n3087) );
  OR2_X1 U2950 ( .A1(n2585), .A2(n2577), .ZN(n3683) );
  INV_X1 U2951 ( .A(n3335), .ZN(n3707) );
  NOR2_X1 U2952 ( .A1(n2572), .A2(n2574), .ZN(n3866) );
  NOR2_X1 U2953 ( .A1(n3436), .A2(n3695), .ZN(n3443) );
  AOI21_X1 U2954 ( .B1(n4437), .B2(ADDR_REG_18__SCAN_IN), .A(n4436), .ZN(n4438) );
  MUX2_X1 U2955 ( .A(n4472), .B(n4471), .S(n4862), .Z(n3641) );
  INV_X1 U2956 ( .A(n4316), .ZN(n3950) );
  OR2_X1 U2957 ( .A1(n2564), .A2(D_REG_1__SCAN_IN), .ZN(n2735) );
  OR2_X1 U2958 ( .A1(n2564), .A2(D_REG_0__SCAN_IN), .ZN(n2563) );
  NOR2_X1 U2959 ( .A1(n3208), .A2(n3207), .ZN(n3247) );
  AND2_X1 U2960 ( .A1(n3387), .A2(REG3_REG_19__SCAN_IN), .ZN(n3393) );
  OR2_X1 U2961 ( .A1(n3398), .A2(n3621), .ZN(n3404) );
  OR2_X1 U2962 ( .A1(n3404), .A2(n4585), .ZN(n3410) );
  AND2_X1 U2963 ( .A1(n3417), .A2(n3416), .ZN(n4085) );
  AND2_X1 U2964 ( .A1(n3358), .A2(n3357), .ZN(n4173) );
  AND2_X1 U2965 ( .A1(n3090), .A2(n3089), .ZN(n3215) );
  INV_X1 U2966 ( .A(n4438), .ZN(n4439) );
  INV_X1 U2967 ( .A(n4190), .ZN(n4175) );
  NAND2_X1 U2968 ( .A1(n2759), .A2(n2758), .ZN(n2802) );
  AND2_X1 U2970 ( .A1(n4537), .A2(n4510), .ZN(n4215) );
  AND2_X1 U2971 ( .A1(n2563), .A2(n2562), .ZN(n2636) );
  AND2_X1 U2972 ( .A1(n4524), .A2(n4510), .ZN(n4276) );
  NAND2_X1 U2973 ( .A1(n2403), .A2(n2404), .ZN(n2564) );
  XNOR2_X1 U2974 ( .A(n2442), .B(n2441), .ZN(n2880) );
  AND2_X1 U2975 ( .A1(n2448), .A2(n2419), .ZN(n4437) );
  AND2_X1 U2976 ( .A1(n2675), .A2(n2674), .ZN(n4342) );
  OR2_X1 U2977 ( .A1(n2585), .A2(n2567), .ZN(n3712) );
  NAND2_X1 U2978 ( .A1(n3460), .A2(n3459), .ZN(n3967) );
  OAI211_X1 U2979 ( .C1(n2609), .C2(n4111), .A(n3402), .B(n3401), .ZN(n4123)
         );
  INV_X1 U2980 ( .A(n3215), .ZN(n3877) );
  OR2_X1 U2981 ( .A1(n3173), .A2(n3172), .ZN(n3199) );
  INV_X1 U2982 ( .A(n4107), .ZN(n4203) );
  AND2_X2 U2983 ( .A1(n2739), .A2(n4197), .ZN(n4465) );
  INV_X1 U2984 ( .A(n4215), .ZN(n4264) );
  INV_X1 U2985 ( .A(n4276), .ZN(n4310) );
  INV_X1 U2986 ( .A(n4524), .ZN(n4522) );
  INV_X1 U2987 ( .A(n4467), .ZN(n4466) );
  NOR2_X1 U2988 ( .A1(n2455), .A2(n2454), .ZN(n4314) );
  AND2_X1 U2989 ( .A1(n2671), .A2(STATE_REG_SCAN_IN), .ZN(n4468) );
  INV_X1 U2990 ( .A(n3199), .ZN(n4318) );
  INV_X1 U2991 ( .A(n3889), .ZN(U4043) );
  INV_X1 U2992 ( .A(n2370), .ZN(n2338) );
  NOR2_X1 U2993 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2342)
         );
  NAND2_X1 U2994 ( .A1(n3370), .A2(n2343), .ZN(n2379) );
  INV_X1 U2995 ( .A(n2379), .ZN(n2345) );
  NAND2_X1 U2996 ( .A1(n2345), .A2(n2344), .ZN(n2397) );
  INV_X1 U2997 ( .A(IR_REG_23__SCAN_IN), .ZN(n2346) );
  AND2_X1 U2998 ( .A1(n2412), .A2(n2346), .ZN(n2347) );
  NAND2_X1 U2999 ( .A1(n2411), .A2(n2347), .ZN(n2348) );
  OR2_X1 U3000 ( .A1(n2385), .A2(n3170), .ZN(n2355) );
  NAND2_X1 U3001 ( .A1(n2356), .A2(IR_REG_31__SCAN_IN), .ZN(n2357) );
  MUX2_X1 U3002 ( .A(IR_REG_31__SCAN_IN), .B(n2357), .S(IR_REG_25__SCAN_IN), 
        .Z(n2359) );
  INV_X1 U3003 ( .A(n2385), .ZN(n2358) );
  NAND2_X1 U3004 ( .A1(n2359), .A2(n2358), .ZN(n2408) );
  NAND2_X1 U3005 ( .A1(n2411), .A2(n2412), .ZN(n2361) );
  NAND2_X1 U3006 ( .A1(n2361), .A2(IR_REG_31__SCAN_IN), .ZN(n2362) );
  INV_X1 U3007 ( .A(n4468), .ZN(n2405) );
  OR2_X2 U3008 ( .A1(n2518), .A2(n2405), .ZN(n3889) );
  INV_X2 U3009 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND2_X1 U3010 ( .A1(n2363), .A2(IR_REG_31__SCAN_IN), .ZN(n2364) );
  MUX2_X1 U3011 ( .A(IR_REG_31__SCAN_IN), .B(n2364), .S(IR_REG_5__SCAN_IN), 
        .Z(n2367) );
  INV_X1 U3012 ( .A(n2365), .ZN(n2366) );
  NAND2_X1 U3013 ( .A1(n2367), .A2(n2366), .ZN(n2717) );
  INV_X1 U3014 ( .A(DATAI_5_), .ZN(n2368) );
  MUX2_X1 U3015 ( .A(n2717), .B(n2368), .S(U3149), .Z(n2369) );
  INV_X1 U3016 ( .A(n2369), .ZN(U3347) );
  INV_X1 U3017 ( .A(DATAI_4_), .ZN(n4729) );
  NAND2_X1 U3018 ( .A1(n2371), .A2(IR_REG_31__SCAN_IN), .ZN(n2432) );
  NAND2_X1 U3019 ( .A1(n2432), .A2(n2372), .ZN(n2373) );
  NAND2_X1 U3020 ( .A1(n2373), .A2(IR_REG_31__SCAN_IN), .ZN(n2375) );
  XNOR2_X1 U3021 ( .A(n2375), .B(n2374), .ZN(n4360) );
  MUX2_X1 U3022 ( .A(n4729), .B(n4360), .S(STATE_REG_SCAN_IN), .Z(n2376) );
  INV_X1 U3023 ( .A(n2376), .ZN(U3348) );
  NAND2_X1 U3024 ( .A1(U3149), .A2(DATAI_25_), .ZN(n2377) );
  OAI21_X1 U3025 ( .B1(n2408), .B2(U3149), .A(n2377), .ZN(U3327) );
  INV_X1 U3026 ( .A(DATAI_26_), .ZN(n4543) );
  NAND2_X1 U3027 ( .A1(n2404), .A2(STATE_REG_SCAN_IN), .ZN(n2378) );
  OAI21_X1 U3028 ( .B1(STATE_REG_SCAN_IN), .B2(n4543), .A(n2378), .ZN(U3326)
         );
  INV_X1 U3029 ( .A(DATAI_20_), .ZN(n4596) );
  NAND2_X1 U3030 ( .A1(n2379), .A2(IR_REG_31__SCAN_IN), .ZN(n2535) );
  INV_X1 U3031 ( .A(IR_REG_19__SCAN_IN), .ZN(n2380) );
  NAND2_X1 U3032 ( .A1(n2535), .A2(n2380), .ZN(n2381) );
  INV_X1 U3033 ( .A(IR_REG_20__SCAN_IN), .ZN(n2382) );
  INV_X1 U3034 ( .A(n3859), .ZN(n2618) );
  NAND2_X1 U3035 ( .A1(n2618), .A2(STATE_REG_SCAN_IN), .ZN(n2384) );
  OAI21_X1 U3036 ( .B1(STATE_REG_SCAN_IN), .B2(n4596), .A(n2384), .ZN(U3332)
         );
  INV_X1 U3037 ( .A(DATAI_30_), .ZN(n4829) );
  NOR2_X1 U3038 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_29__SCAN_IN), .ZN(n2386)
         );
  NAND2_X1 U3039 ( .A1(n2451), .A2(n2386), .ZN(n2391) );
  OAI21_X1 U3040 ( .B1(STATE_REG_SCAN_IN), .B2(n4829), .A(n2388), .ZN(U3322)
         );
  INV_X1 U3041 ( .A(DATAI_29_), .ZN(n2394) );
  NAND2_X1 U3042 ( .A1(n2453), .A2(IR_REG_31__SCAN_IN), .ZN(n2389) );
  NAND2_X1 U3043 ( .A1(n2520), .A2(STATE_REG_SCAN_IN), .ZN(n2393) );
  OAI21_X1 U3044 ( .B1(STATE_REG_SCAN_IN), .B2(n2394), .A(n2393), .ZN(U3323)
         );
  INV_X1 U3045 ( .A(DATAI_31_), .ZN(n2396) );
  OR4_X1 U3046 ( .A1(n2391), .A2(IR_REG_30__SCAN_IN), .A3(n3170), .A4(U3149), 
        .ZN(n2395) );
  OAI21_X1 U3047 ( .B1(STATE_REG_SCAN_IN), .B2(n2396), .A(n2395), .ZN(U3321)
         );
  INV_X1 U3048 ( .A(DATAI_21_), .ZN(n4540) );
  INV_X1 U3049 ( .A(IR_REG_21__SCAN_IN), .ZN(n2398) );
  NAND2_X1 U3050 ( .A1(n2517), .A2(STATE_REG_SCAN_IN), .ZN(n2400) );
  OAI21_X1 U3051 ( .B1(STATE_REG_SCAN_IN), .B2(n4540), .A(n2400), .ZN(U3331)
         );
  NAND2_X1 U3052 ( .A1(n2408), .A2(B_REG_SCAN_IN), .ZN(n2402) );
  MUX2_X1 U3053 ( .A(n2402), .B(B_REG_SCAN_IN), .S(n2401), .Z(n2403) );
  INV_X1 U3054 ( .A(n2734), .ZN(n2575) );
  INV_X1 U3055 ( .A(D_REG_0__SCAN_IN), .ZN(n2407) );
  NOR3_X1 U3056 ( .A1(n2405), .A2(n2404), .A3(n2401), .ZN(n2406) );
  AOI21_X1 U3057 ( .B1(n4467), .B2(n2407), .A(n2406), .ZN(U3458) );
  INV_X1 U3058 ( .A(D_REG_1__SCAN_IN), .ZN(n2410) );
  NAND2_X1 U3059 ( .A1(n2560), .A2(n2408), .ZN(n2627) );
  INV_X1 U3060 ( .A(n2627), .ZN(n2409) );
  AOI22_X1 U3061 ( .A1(n4467), .A2(n2410), .B1(n4468), .B2(n2409), .ZN(U3459)
         );
  OR2_X1 U3062 ( .A1(n2671), .A2(U3149), .ZN(n3870) );
  NAND2_X1 U3063 ( .A1(n2734), .A2(n3870), .ZN(n2448) );
  NAND2_X1 U3064 ( .A1(n4315), .A2(n2517), .ZN(n2614) );
  INV_X1 U3065 ( .A(n2614), .ZN(n2621) );
  NAND2_X1 U3066 ( .A1(n2385), .A2(n2414), .ZN(n2415) );
  NAND2_X1 U3067 ( .A1(n2417), .A2(IR_REG_27__SCAN_IN), .ZN(n2418) );
  AOI21_X1 U3068 ( .B1(n2621), .B2(n2671), .A(n2653), .ZN(n2447) );
  INV_X1 U3069 ( .A(n2447), .ZN(n2419) );
  NOR2_X1 U3070 ( .A1(n4437), .A2(U4043), .ZN(U3148) );
  INV_X1 U3071 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n2425) );
  INV_X1 U3072 ( .A(REG1_REG_30__SCAN_IN), .ZN(n2423) );
  NAND2_X1 U3073 ( .A1(n3725), .A2(REG2_REG_30__SCAN_IN), .ZN(n2422) );
  NAND2_X1 U3074 ( .A1(n3445), .A2(REG0_REG_30__SCAN_IN), .ZN(n2421) );
  OAI211_X1 U3075 ( .C1(n3729), .C2(n2423), .A(n2422), .B(n2421), .ZN(n3959)
         );
  NAND2_X1 U3076 ( .A1(U4043), .A2(n3959), .ZN(n2424) );
  OAI21_X1 U3077 ( .B1(U4043), .B2(n2425), .A(n2424), .ZN(U3580) );
  INV_X1 U3078 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2998) );
  INV_X1 U3079 ( .A(n2717), .ZN(n2500) );
  OR2_X1 U3080 ( .A1(n2426), .A2(n3170), .ZN(n2428) );
  XNOR2_X1 U3081 ( .A(n3902), .B(REG1_REG_2__SCAN_IN), .ZN(n3901) );
  INV_X1 U3082 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4527) );
  INV_X1 U3083 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4525) );
  NOR2_X1 U3084 ( .A1(n4547), .A2(n4525), .ZN(n3893) );
  INV_X1 U3085 ( .A(n3893), .ZN(n2429) );
  AOI21_X1 U3086 ( .B1(n3890), .B2(n4527), .A(n2429), .ZN(n2430) );
  NAND2_X1 U3087 ( .A1(n2430), .A2(n2431), .ZN(n3891) );
  NAND2_X1 U3088 ( .A1(n3891), .A2(n2431), .ZN(n3900) );
  INV_X1 U3089 ( .A(n3902), .ZN(n4324) );
  XNOR2_X1 U3090 ( .A(n2432), .B(IR_REG_3__SCAN_IN), .ZN(n4323) );
  XNOR2_X1 U3091 ( .A(n2433), .B(n2493), .ZN(n2487) );
  INV_X1 U3092 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2434) );
  OAI22_X1 U3093 ( .A1(n2487), .A2(n2434), .B1(n2433), .B2(n2493), .ZN(n2435)
         );
  XNOR2_X1 U3094 ( .A(n2435), .B(n4360), .ZN(n4359) );
  INV_X1 U3095 ( .A(n4360), .ZN(n2467) );
  INV_X1 U3096 ( .A(REG1_REG_5__SCAN_IN), .ZN(n4606) );
  MUX2_X1 U3097 ( .A(REG1_REG_5__SCAN_IN), .B(n4606), .S(n2717), .Z(n2497) );
  OR2_X1 U3098 ( .A1(n2365), .A2(n3170), .ZN(n2436) );
  XNOR2_X1 U3099 ( .A(n2436), .B(IR_REG_6__SCAN_IN), .ZN(n4322) );
  INV_X1 U3100 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2438) );
  OAI22_X1 U3101 ( .A1(n2480), .A2(n2438), .B1(n2437), .B2(n2482), .ZN(n2507)
         );
  OR2_X1 U3102 ( .A1(n2439), .A2(n3170), .ZN(n2442) );
  INV_X1 U3103 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4601) );
  NOR2_X1 U3104 ( .A1(n2880), .A2(n4601), .ZN(n2440) );
  INV_X1 U3105 ( .A(n2880), .ZN(n4321) );
  OAI22_X1 U3106 ( .A1(n2507), .A2(n2440), .B1(REG1_REG_7__SCAN_IN), .B2(n4321), .ZN(n2446) );
  NAND2_X1 U3107 ( .A1(n2442), .A2(n2441), .ZN(n2443) );
  NAND2_X1 U3108 ( .A1(n2443), .A2(IR_REG_31__SCAN_IN), .ZN(n2445) );
  INV_X1 U3109 ( .A(IR_REG_8__SCAN_IN), .ZN(n2444) );
  XNOR2_X1 U3110 ( .A(n2445), .B(n2444), .ZN(n2895) );
  NOR2_X1 U3111 ( .A1(n2446), .A2(n2895), .ZN(n2706) );
  NAND2_X1 U3112 ( .A1(n2448), .A2(n2447), .ZN(n4356) );
  XNOR2_X1 U3113 ( .A(n2449), .B(IR_REG_27__SCAN_IN), .ZN(n4353) );
  AOI211_X1 U3114 ( .C1(n2998), .C2(n2450), .A(n2705), .B(n4433), .ZN(n2459)
         );
  NOR2_X1 U3115 ( .A1(n2451), .A2(n3170), .ZN(n2452) );
  MUX2_X1 U3116 ( .A(n3170), .B(n2452), .S(IR_REG_28__SCAN_IN), .Z(n2455) );
  INV_X1 U3117 ( .A(n2453), .ZN(n2454) );
  NAND2_X1 U3118 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n2909) );
  INV_X1 U3119 ( .A(n2909), .ZN(n2456) );
  AOI21_X1 U3120 ( .B1(n4437), .B2(ADDR_REG_8__SCAN_IN), .A(n2456), .ZN(n2457)
         );
  OAI21_X1 U3121 ( .B1(n4449), .B2(n2895), .A(n2457), .ZN(n2458) );
  NOR2_X1 U3122 ( .A1(n2459), .A2(n2458), .ZN(n2478) );
  INV_X1 U3123 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2460) );
  MUX2_X1 U3124 ( .A(n2460), .B(REG2_REG_2__SCAN_IN), .S(n3902), .Z(n3907) );
  XNOR2_X1 U3125 ( .A(n3890), .B(REG2_REG_1__SCAN_IN), .ZN(n3894) );
  AND2_X1 U3126 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3911)
         );
  NAND2_X1 U3127 ( .A1(n3894), .A2(n3911), .ZN(n2462) );
  INV_X1 U3128 ( .A(n3890), .ZN(n4325) );
  NAND2_X1 U3129 ( .A1(n4325), .A2(REG2_REG_1__SCAN_IN), .ZN(n2461) );
  NAND2_X1 U3130 ( .A1(n2462), .A2(n2461), .ZN(n3906) );
  NAND2_X1 U3131 ( .A1(n3907), .A2(n3906), .ZN(n3905) );
  NAND2_X1 U3132 ( .A1(n4324), .A2(REG2_REG_2__SCAN_IN), .ZN(n2463) );
  NAND2_X1 U3133 ( .A1(n2488), .A2(REG2_REG_3__SCAN_IN), .ZN(n2466) );
  NAND2_X1 U3134 ( .A1(n2464), .A2(n4323), .ZN(n2465) );
  NAND2_X1 U3135 ( .A1(n2468), .A2(n2467), .ZN(n2469) );
  INV_X1 U3136 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2835) );
  MUX2_X1 U3137 ( .A(n2835), .B(REG2_REG_5__SCAN_IN), .S(n2717), .Z(n2503) );
  NAND2_X1 U3138 ( .A1(n2500), .A2(REG2_REG_5__SCAN_IN), .ZN(n2470) );
  NAND2_X1 U3139 ( .A1(n2471), .A2(n4322), .ZN(n2472) );
  INV_X1 U3140 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2473) );
  MUX2_X1 U3141 ( .A(n2473), .B(REG2_REG_7__SCAN_IN), .S(n2880), .Z(n2474) );
  OR2_X1 U3142 ( .A1(n2880), .A2(n2473), .ZN(n2475) );
  NAND2_X1 U3143 ( .A1(n4314), .A2(n4353), .ZN(n3909) );
  OR2_X1 U3144 ( .A1(n4356), .A2(n3909), .ZN(n4398) );
  OAI211_X1 U3145 ( .C1(n2476), .C2(REG2_REG_8__SCAN_IN), .A(n4445), .B(n2700), 
        .ZN(n2477) );
  NAND2_X1 U3146 ( .A1(n2478), .A2(n2477), .ZN(U3248) );
  XNOR2_X1 U3147 ( .A(n2479), .B(REG2_REG_6__SCAN_IN), .ZN(n2486) );
  XNOR2_X1 U31480 ( .A(n2480), .B(REG1_REG_6__SCAN_IN), .ZN(n2484) );
  INV_X1 U31490 ( .A(n4433), .ZN(n4429) );
  NOR2_X1 U3150 ( .A1(STATE_REG_SCAN_IN), .A2(n2719), .ZN(n2792) );
  AOI21_X1 U3151 ( .B1(n4437), .B2(ADDR_REG_6__SCAN_IN), .A(n2792), .ZN(n2481)
         );
  OAI21_X1 U3152 ( .B1(n4449), .B2(n2482), .A(n2481), .ZN(n2483) );
  AOI21_X1 U3153 ( .B1(n2484), .B2(n4429), .A(n2483), .ZN(n2485) );
  OAI21_X1 U3154 ( .B1(n2486), .B2(n4398), .A(n2485), .ZN(U3246) );
  XNOR2_X1 U3155 ( .A(n2487), .B(REG1_REG_3__SCAN_IN), .ZN(n2490) );
  INV_X1 U3156 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2768) );
  XNOR2_X1 U3157 ( .A(n2488), .B(n2768), .ZN(n2489) );
  AOI22_X1 U3158 ( .A1(n4429), .A2(n2490), .B1(n4445), .B2(n2489), .ZN(n2492)
         );
  INV_X1 U3159 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4549) );
  NOR2_X1 U3160 ( .A1(STATE_REG_SCAN_IN), .A2(n4549), .ZN(n2690) );
  AOI21_X1 U3161 ( .B1(n4437), .B2(ADDR_REG_3__SCAN_IN), .A(n2690), .ZN(n2491)
         );
  OAI211_X1 U3162 ( .C1(n2493), .C2(n4449), .A(n2492), .B(n2491), .ZN(U3243)
         );
  INV_X1 U3163 ( .A(n4449), .ZN(n4407) );
  INV_X1 U3164 ( .A(n4437), .ZN(n4410) );
  INV_X1 U3165 ( .A(ADDR_REG_5__SCAN_IN), .ZN(n2495) );
  AND2_X1 U3166 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n2726) );
  INV_X1 U3167 ( .A(n2726), .ZN(n2494) );
  OAI21_X1 U3168 ( .B1(n4410), .B2(n2495), .A(n2494), .ZN(n2499) );
  AOI211_X1 U3169 ( .C1(n2182), .C2(n2497), .A(n2496), .B(n4433), .ZN(n2498)
         );
  AOI211_X1 U3170 ( .C1(n4407), .C2(n2500), .A(n2499), .B(n2498), .ZN(n2505)
         );
  OAI211_X1 U3171 ( .C1(n2503), .C2(n2502), .A(n4445), .B(n2501), .ZN(n2504)
         );
  NAND2_X1 U3172 ( .A1(n2505), .A2(n2504), .ZN(U3245) );
  XOR2_X1 U3173 ( .A(n4601), .B(n2880), .Z(n2506) );
  XNOR2_X1 U3174 ( .A(n2507), .B(n2506), .ZN(n2516) );
  INV_X1 U3175 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2508) );
  NOR2_X1 U3176 ( .A1(STATE_REG_SCAN_IN), .A2(n2508), .ZN(n3001) );
  NOR2_X1 U3177 ( .A1(n4449), .A2(n2880), .ZN(n2509) );
  AOI211_X1 U3178 ( .C1(n4437), .C2(ADDR_REG_7__SCAN_IN), .A(n3001), .B(n2509), 
        .ZN(n2515) );
  MUX2_X1 U3179 ( .A(REG2_REG_7__SCAN_IN), .B(n2473), .S(n2880), .Z(n2510) );
  INV_X1 U3180 ( .A(n2510), .ZN(n2513) );
  OAI211_X1 U3181 ( .C1(n2513), .C2(n2512), .A(n4445), .B(n2511), .ZN(n2514)
         );
  OAI211_X1 U3182 ( .C1(n2516), .C2(n4433), .A(n2515), .B(n2514), .ZN(U3247)
         );
  OR2_X2 U3183 ( .A1(n3577), .A2(n4510), .ZN(n3531) );
  INV_X2 U3184 ( .A(n2542), .ZN(n2608) );
  NAND2_X1 U3185 ( .A1(n2608), .A2(REG1_REG_0__SCAN_IN), .ZN(n2524) );
  NAND2_X1 U3186 ( .A1(n2543), .A2(REG0_REG_0__SCAN_IN), .ZN(n2523) );
  NAND2_X1 U3187 ( .A1(n2159), .A2(REG2_REG_0__SCAN_IN), .ZN(n2522) );
  NAND2_X1 U3188 ( .A1(n2607), .A2(REG3_REG_0__SCAN_IN), .ZN(n2521) );
  NAND3_X1 U3189 ( .A1(n2524), .A2(n2523), .A3(n2334), .ZN(n2598) );
  INV_X1 U3190 ( .A(n2598), .ZN(n2525) );
  INV_X1 U3191 ( .A(n2740), .ZN(n2526) );
  INV_X1 U3192 ( .A(n2518), .ZN(n2529) );
  NAND2_X1 U3193 ( .A1(n2531), .A2(n2530), .ZN(n2591) );
  OR2_X1 U3194 ( .A1(n3577), .A2(n2841), .ZN(n2533) );
  NAND2_X1 U3195 ( .A1(n2598), .A2(n3561), .ZN(n2532) );
  AND2_X1 U3196 ( .A1(n2533), .A2(n2532), .ZN(n2538) );
  OR2_X1 U3197 ( .A1(n2518), .A2(n4525), .ZN(n2534) );
  NAND2_X1 U3198 ( .A1(n2538), .A2(n2534), .ZN(n2592) );
  NAND2_X1 U3199 ( .A1(n2591), .A2(n2592), .ZN(n2540) );
  NOR2_X1 U3200 ( .A1(n2536), .A2(n4316), .ZN(n2573) );
  INV_X1 U3201 ( .A(n2573), .ZN(n2537) );
  NAND2_X1 U3202 ( .A1(n2538), .A2(n3571), .ZN(n2539) );
  NAND2_X1 U3203 ( .A1(n2540), .A2(n2539), .ZN(n2641) );
  INV_X1 U3204 ( .A(DATAI_1_), .ZN(n2541) );
  NAND2_X1 U3205 ( .A1(n2608), .A2(REG1_REG_1__SCAN_IN), .ZN(n2547) );
  NAND2_X1 U3206 ( .A1(n2607), .A2(REG3_REG_1__SCAN_IN), .ZN(n2546) );
  NAND2_X1 U3207 ( .A1(n2159), .A2(REG2_REG_1__SCAN_IN), .ZN(n2545) );
  NAND2_X1 U3208 ( .A1(n2543), .A2(REG0_REG_1__SCAN_IN), .ZN(n2544) );
  XNOR2_X1 U3209 ( .A(n2642), .B(n2643), .ZN(n2640) );
  XNOR2_X1 U32100 ( .A(n2641), .B(n2640), .ZN(n2590) );
  NOR4_X1 U32110 ( .A1(D_REG_5__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_10__SCAN_IN), .ZN(n2552) );
  NOR4_X1 U32120 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_25__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_4__SCAN_IN), .ZN(n2551) );
  NOR4_X1 U32130 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2550) );
  NOR4_X1 U32140 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_13__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2549) );
  NAND4_X1 U32150 ( .A1(n2552), .A2(n2551), .A3(n2550), .A4(n2549), .ZN(n2558)
         );
  NOR2_X1 U32160 ( .A1(D_REG_30__SCAN_IN), .A2(D_REG_26__SCAN_IN), .ZN(n2556)
         );
  NOR4_X1 U32170 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n2555) );
  NOR4_X1 U32180 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_28__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_14__SCAN_IN), .ZN(n2554) );
  NOR4_X1 U32190 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_3__SCAN_IN), .ZN(n2553) );
  NAND4_X1 U32200 ( .A1(n2556), .A2(n2555), .A3(n2554), .A4(n2553), .ZN(n2557)
         );
  NOR2_X1 U32210 ( .A1(n2558), .A2(n2557), .ZN(n2559) );
  NAND2_X1 U32220 ( .A1(n2561), .A2(n2560), .ZN(n2562) );
  NAND3_X1 U32230 ( .A1(n2737), .A2(n2636), .A3(n2735), .ZN(n2585) );
  AND2_X1 U32240 ( .A1(n3859), .A2(n3950), .ZN(n2570) );
  INV_X1 U32250 ( .A(n2570), .ZN(n2565) );
  NAND2_X1 U32260 ( .A1(n2742), .A2(n2565), .ZN(n2566) );
  NAND2_X1 U32270 ( .A1(n2566), .A2(n2614), .ZN(n2568) );
  OR2_X1 U32280 ( .A1(n2734), .A2(n2568), .ZN(n2567) );
  NAND2_X1 U32290 ( .A1(n4207), .A2(n2568), .ZN(n2569) );
  NAND2_X1 U32300 ( .A1(n2585), .A2(n2569), .ZN(n2571) );
  OR2_X1 U32310 ( .A1(n2614), .A2(n2570), .ZN(n2732) );
  NAND2_X1 U32320 ( .A1(n2571), .A2(n2732), .ZN(n2673) );
  INV_X1 U32330 ( .A(n2673), .ZN(n2576) );
  NAND2_X1 U32340 ( .A1(n4468), .A2(n2573), .ZN(n2574) );
  NAND2_X1 U32350 ( .A1(n2585), .A2(n3866), .ZN(n2674) );
  NAND3_X1 U32360 ( .A1(n2576), .A2(n2575), .A3(n2674), .ZN(n2754) );
  NAND2_X1 U32370 ( .A1(n3866), .A2(n4314), .ZN(n2577) );
  INV_X1 U32380 ( .A(n4314), .ZN(n2578) );
  NAND2_X1 U32390 ( .A1(n3866), .A2(n2578), .ZN(n2579) );
  NAND2_X1 U32400 ( .A1(n2607), .A2(REG3_REG_2__SCAN_IN), .ZN(n2581) );
  NAND2_X1 U32410 ( .A1(n2159), .A2(REG2_REG_2__SCAN_IN), .ZN(n2580) );
  NAND2_X1 U32420 ( .A1(n2608), .A2(REG1_REG_2__SCAN_IN), .ZN(n2583) );
  NAND2_X1 U32430 ( .A1(n2543), .A2(REG0_REG_2__SCAN_IN), .ZN(n2582) );
  OAI22_X1 U32440 ( .A1(n2525), .A2(n3683), .B1(n4335), .B2(n2763), .ZN(n2588)
         );
  OR2_X1 U32450 ( .A1(n2734), .A2(n4207), .ZN(n2584) );
  OR2_X1 U32460 ( .A1(n2585), .A2(n2584), .ZN(n2586) );
  AND2_X1 U32470 ( .A1(n3859), .A2(n4316), .ZN(n2744) );
  NAND2_X1 U32480 ( .A1(n4521), .A2(n2519), .ZN(n2628) );
  AND2_X2 U32490 ( .A1(n2586), .A2(n4197), .ZN(n3684) );
  NOR2_X1 U32500 ( .A1(n3684), .A2(n2846), .ZN(n2587) );
  AOI211_X1 U32510 ( .C1(REG3_REG_1__SCAN_IN), .C2(n2754), .A(n2588), .B(n2587), .ZN(n2589) );
  OAI21_X1 U32520 ( .B1(n2590), .B2(n3712), .A(n2589), .ZN(U3219) );
  NAND2_X1 U32530 ( .A1(n2754), .A2(REG3_REG_0__SCAN_IN), .ZN(n2595) );
  XNOR2_X1 U32540 ( .A(n2592), .B(n2591), .ZN(n3908) );
  INV_X1 U32550 ( .A(n3908), .ZN(n2593) );
  AOI22_X1 U32560 ( .A1(n2593), .A2(n4337), .B1(n3704), .B2(n3888), .ZN(n2594)
         );
  OAI211_X1 U32570 ( .C1(n3684), .C2(n2841), .A(n2595), .B(n2594), .ZN(U3229)
         );
  INV_X1 U32580 ( .A(n2597), .ZN(n2596) );
  INV_X1 U32590 ( .A(n2846), .ZN(n2599) );
  NAND2_X1 U32600 ( .A1(n2596), .A2(n2599), .ZN(n3791) );
  NAND2_X1 U32610 ( .A1(n2597), .A2(n2846), .ZN(n3788) );
  NAND2_X1 U32620 ( .A1(n3791), .A2(n3788), .ZN(n2616) );
  NAND2_X1 U32630 ( .A1(n2616), .A2(n2843), .ZN(n2842) );
  NAND2_X1 U32640 ( .A1(n3888), .A2(n2599), .ZN(n2600) );
  INV_X1 U32650 ( .A(DATAI_2_), .ZN(n2601) );
  NAND2_X1 U32660 ( .A1(n3887), .A2(n2757), .ZN(n3795) );
  NAND2_X1 U32670 ( .A1(n2605), .A2(n2615), .ZN(n2759) );
  OAI21_X1 U32680 ( .B1(n2605), .B2(n2615), .A(n2759), .ZN(n4458) );
  XNOR2_X1 U32690 ( .A(n2740), .B(n4315), .ZN(n2606) );
  NAND2_X1 U32700 ( .A1(n2606), .A2(n3950), .ZN(n3219) );
  INV_X1 U32710 ( .A(n3219), .ZN(n2625) );
  NAND2_X1 U32720 ( .A1(n3412), .A2(n4549), .ZN(n2613) );
  NAND2_X1 U32730 ( .A1(n2608), .A2(REG1_REG_3__SCAN_IN), .ZN(n2612) );
  NAND2_X1 U32740 ( .A1(n2543), .A2(REG0_REG_3__SCAN_IN), .ZN(n2611) );
  NAND4_X1 U32750 ( .A1(n2613), .A2(n2612), .A3(n2611), .A4(n2610), .ZN(n3886)
         );
  INV_X1 U32760 ( .A(n2615), .ZN(n3775) );
  OR2_X1 U32770 ( .A1(n2598), .A2(n2841), .ZN(n3787) );
  OAI21_X1 U32780 ( .B1(n2616), .B2(n3787), .A(n3791), .ZN(n2617) );
  NAND2_X1 U32790 ( .A1(n2617), .A2(n3775), .ZN(n2760) );
  OAI21_X1 U32800 ( .B1(n3775), .B2(n2617), .A(n2760), .ZN(n2620) );
  NAND2_X1 U32810 ( .A1(n4315), .A2(n4316), .ZN(n2619) );
  NAND2_X1 U32820 ( .A1(n2618), .A2(n2517), .ZN(n3863) );
  NAND2_X1 U32830 ( .A1(n2620), .A2(n4175), .ZN(n2623) );
  AOI22_X1 U32840 ( .A1(n3888), .A2(n4188), .B1(n2604), .B2(n4217), .ZN(n2622)
         );
  OAI211_X1 U32850 ( .C1(n2804), .C2(n4185), .A(n2623), .B(n2622), .ZN(n2624)
         );
  AOI21_X1 U32860 ( .B1(n2625), .B2(n4458), .A(n2624), .ZN(n4464) );
  INV_X1 U32870 ( .A(n4464), .ZN(n2626) );
  AOI21_X1 U32880 ( .B1(n4521), .B2(n4458), .A(n2626), .ZN(n2639) );
  NAND2_X1 U32890 ( .A1(n2735), .A2(n2627), .ZN(n2632) );
  NAND2_X1 U32900 ( .A1(n2628), .A2(n2732), .ZN(n2629) );
  NOR2_X1 U32910 ( .A1(n2734), .A2(n2629), .ZN(n2631) );
  INV_X1 U32920 ( .A(n2633), .ZN(n2840) );
  NAND2_X1 U32930 ( .A1(n2840), .A2(n2604), .ZN(n2634) );
  NAND2_X1 U32940 ( .A1(n2633), .A2(n2757), .ZN(n2767) );
  AND2_X1 U32950 ( .A1(n2634), .A2(n2767), .ZN(n4460) );
  AOI22_X1 U32960 ( .A1(n4215), .A2(n4460), .B1(n4534), .B2(
        REG1_REG_2__SCAN_IN), .ZN(n2635) );
  OAI21_X1 U32970 ( .B1(n2639), .B2(n4534), .A(n2635), .ZN(U3520) );
  AOI22_X1 U32980 ( .A1(n4276), .A2(n4460), .B1(n4522), .B2(
        REG0_REG_2__SCAN_IN), .ZN(n2638) );
  OAI21_X1 U32990 ( .B1(n2639), .B2(n4522), .A(n2638), .ZN(U3471) );
  INV_X1 U33000 ( .A(n2642), .ZN(n2644) );
  NAND2_X1 U33010 ( .A1(n2644), .A2(n2643), .ZN(n2645) );
  NAND2_X1 U33020 ( .A1(n3887), .A2(n3561), .ZN(n2647) );
  OR2_X1 U33030 ( .A1(n3577), .A2(n2757), .ZN(n2646) );
  NAND2_X1 U33040 ( .A1(n2647), .A2(n2646), .ZN(n2648) );
  XNOR2_X1 U33050 ( .A(n2648), .B(n3571), .ZN(n2651) );
  NOR2_X1 U33060 ( .A1(n3576), .A2(n2757), .ZN(n2649) );
  NAND2_X1 U33070 ( .A1(n2651), .A2(n2650), .ZN(n2652) );
  NAND2_X1 U33080 ( .A1(n2749), .A2(n2652), .ZN(n2687) );
  NAND2_X1 U33090 ( .A1(n3886), .A2(n3561), .ZN(n2655) );
  MUX2_X1 U33100 ( .A(n4323), .B(DATAI_3_), .S(n3734), .Z(n2761) );
  NAND2_X1 U33110 ( .A1(n2655), .A2(n2654), .ZN(n2656) );
  XNOR2_X1 U33120 ( .A(n2656), .B(n3571), .ZN(n2667) );
  OAI22_X1 U33130 ( .A1(n2804), .A2(n3531), .B1(n2803), .B2(n3576), .ZN(n2665)
         );
  XNOR2_X1 U33140 ( .A(n2667), .B(n2665), .ZN(n2688) );
  NAND2_X1 U33150 ( .A1(n2687), .A2(n2688), .ZN(n2686) );
  NAND2_X1 U33160 ( .A1(n2608), .A2(REG1_REG_4__SCAN_IN), .ZN(n2661) );
  NAND2_X1 U33170 ( .A1(n3725), .A2(REG2_REG_4__SCAN_IN), .ZN(n2660) );
  NAND2_X1 U33180 ( .A1(n2543), .A2(REG0_REG_4__SCAN_IN), .ZN(n2659) );
  NOR2_X1 U33190 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2657) );
  NOR2_X1 U33200 ( .A1(n2676), .A2(n2657), .ZN(n2813) );
  NAND2_X1 U33210 ( .A1(n3412), .A2(n2813), .ZN(n2658) );
  NAND2_X1 U33220 ( .A1(n3885), .A2(n3561), .ZN(n2663) );
  MUX2_X1 U33230 ( .A(n4360), .B(n4729), .S(n3734), .Z(n2823) );
  OR2_X1 U33240 ( .A1(n3577), .A2(n2823), .ZN(n2662) );
  NAND2_X1 U33250 ( .A1(n2663), .A2(n2662), .ZN(n2664) );
  XNOR2_X1 U33260 ( .A(n2664), .B(n3571), .ZN(n2712) );
  INV_X1 U33270 ( .A(n3885), .ZN(n2832) );
  OAI22_X1 U33280 ( .A1(n2832), .A2(n3531), .B1(n2823), .B2(n3576), .ZN(n2713)
         );
  XNOR2_X1 U33290 ( .A(n2712), .B(n2713), .ZN(n2669) );
  INV_X1 U33300 ( .A(n2665), .ZN(n2666) );
  NAND2_X1 U33310 ( .A1(n2667), .A2(n2666), .ZN(n2670) );
  AND2_X1 U33320 ( .A1(n2669), .A2(n2670), .ZN(n2668) );
  NAND2_X1 U33330 ( .A1(n2716), .A2(n4337), .ZN(n2685) );
  AOI21_X1 U33340 ( .B1(n2686), .B2(n2670), .A(n2669), .ZN(n2684) );
  NAND2_X1 U33350 ( .A1(n2518), .A2(n2671), .ZN(n2672) );
  OAI21_X1 U33360 ( .B1(n2673), .B2(n2672), .A(STATE_REG_SCAN_IN), .ZN(n2675)
         );
  AOI22_X1 U33370 ( .A1(n2608), .A2(REG1_REG_5__SCAN_IN), .B1(n3445), .B2(
        REG0_REG_5__SCAN_IN), .ZN(n2679) );
  OAI21_X1 U33380 ( .B1(n2676), .B2(REG3_REG_5__SCAN_IN), .A(n2720), .ZN(n2677) );
  INV_X1 U33390 ( .A(n2677), .ZN(n2837) );
  AOI22_X1 U33400 ( .A1(n3412), .A2(n2837), .B1(n3725), .B2(
        REG2_REG_5__SCAN_IN), .ZN(n2678) );
  AND2_X1 U33410 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n4362) );
  AOI21_X1 U33420 ( .B1(n3704), .B2(n3884), .A(n4362), .ZN(n2681) );
  NAND2_X1 U33430 ( .A1(n4327), .A2(n3886), .ZN(n2680) );
  OAI211_X1 U33440 ( .C1(n3684), .C2(n2823), .A(n2681), .B(n2680), .ZN(n2682)
         );
  AOI21_X1 U33450 ( .B1(n3710), .B2(n2813), .A(n2682), .ZN(n2683) );
  OAI21_X1 U33460 ( .B1(n2685), .B2(n2684), .A(n2683), .ZN(U3227) );
  OAI21_X1 U33470 ( .B1(n2688), .B2(n2687), .A(n2686), .ZN(n2689) );
  NAND2_X1 U33480 ( .A1(n2689), .A2(n4337), .ZN(n2695) );
  OAI22_X1 U33490 ( .A1(n3684), .A2(n2803), .B1(n2763), .B2(n3683), .ZN(n2693)
         );
  INV_X1 U33500 ( .A(n2690), .ZN(n2691) );
  OAI21_X1 U33510 ( .B1(n4335), .B2(n2832), .A(n2691), .ZN(n2692) );
  NOR2_X1 U33520 ( .A1(n2693), .A2(n2692), .ZN(n2694) );
  OAI211_X1 U3353 ( .C1(REG3_REG_3__SCAN_IN), .C2(n4342), .A(n2695), .B(n2694), 
        .ZN(U3215) );
  OR2_X1 U33540 ( .A1(n2696), .A2(IR_REG_9__SCAN_IN), .ZN(n3168) );
  NAND2_X1 U3355 ( .A1(n3168), .A2(IR_REG_31__SCAN_IN), .ZN(n2697) );
  XNOR2_X1 U3356 ( .A(n2697), .B(IR_REG_10__SCAN_IN), .ZN(n4319) );
  INV_X1 U3357 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2948) );
  NAND2_X1 U3358 ( .A1(n2696), .A2(IR_REG_31__SCAN_IN), .ZN(n2698) );
  XNOR2_X1 U3359 ( .A(n2698), .B(IR_REG_9__SCAN_IN), .ZN(n2935) );
  INV_X1 U3360 ( .A(n2935), .ZN(n4476) );
  AOI22_X1 U3361 ( .A1(n2935), .A2(REG2_REG_9__SCAN_IN), .B1(n2948), .B2(n4476), .ZN(n4376) );
  INV_X1 U3362 ( .A(n2895), .ZN(n4320) );
  NAND2_X1 U3363 ( .A1(n2699), .A2(n4320), .ZN(n2701) );
  OAI211_X1 U3364 ( .C1(n2702), .C2(REG2_REG_10__SCAN_IN), .A(n4445), .B(n3176), .ZN(n2704) );
  NOR2_X1 U3365 ( .A1(STATE_REG_SCAN_IN), .A2(n4831), .ZN(n3028) );
  AOI21_X1 U3366 ( .B1(n4437), .B2(ADDR_REG_10__SCAN_IN), .A(n3028), .ZN(n2703) );
  OAI211_X1 U3367 ( .C1(n4449), .C2(n2209), .A(n2704), .B(n2703), .ZN(n2711)
         );
  INV_X1 U3368 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3124) );
  INV_X1 U3369 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4602) );
  AOI22_X1 U3370 ( .A1(n2935), .A2(n4602), .B1(REG1_REG_9__SCAN_IN), .B2(n4476), .ZN(n4370) );
  NOR2_X1 U3371 ( .A1(n4371), .A2(n4370), .ZN(n4369) );
  AND2_X1 U3372 ( .A1(n2935), .A2(REG1_REG_9__SCAN_IN), .ZN(n2707) );
  NAND2_X1 U3373 ( .A1(n2708), .A2(n4319), .ZN(n3185) );
  OAI21_X1 U3374 ( .B1(n2708), .B2(n4319), .A(n3185), .ZN(n2709) );
  AOI211_X1 U3375 ( .C1(n3124), .C2(n2709), .A(n3186), .B(n4433), .ZN(n2710)
         );
  OR2_X1 U3376 ( .A1(n2711), .A2(n2710), .ZN(U3250) );
  INV_X1 U3377 ( .A(n2712), .ZN(n2714) );
  NAND2_X1 U3378 ( .A1(n2714), .A2(n2713), .ZN(n2715) );
  MUX2_X1 U3379 ( .A(n2717), .B(n2368), .S(n3734), .Z(n2857) );
  OAI22_X1 U3380 ( .A1(n2867), .A2(n2572), .B1(n2857), .B2(n3577), .ZN(n2718)
         );
  XNOR2_X1 U3381 ( .A(n2718), .B(n3571), .ZN(n2774) );
  OAI22_X1 U3382 ( .A1(n2867), .A2(n3531), .B1(n2857), .B2(n3576), .ZN(n2775)
         );
  XNOR2_X1 U3383 ( .A(n2774), .B(n2775), .ZN(n2772) );
  XNOR2_X1 U3384 ( .A(n2773), .B(n2772), .ZN(n2731) );
  NAND2_X1 U3385 ( .A1(n2608), .A2(REG1_REG_6__SCAN_IN), .ZN(n2725) );
  AND2_X1 U3386 ( .A1(n2720), .A2(n2719), .ZN(n2721) );
  NOR2_X1 U3387 ( .A1(n2786), .A2(n2721), .ZN(n4450) );
  NAND2_X1 U3388 ( .A1(n3412), .A2(n4450), .ZN(n2724) );
  NAND2_X1 U3389 ( .A1(n3445), .A2(REG0_REG_6__SCAN_IN), .ZN(n2723) );
  NAND2_X1 U3390 ( .A1(n3725), .A2(REG2_REG_6__SCAN_IN), .ZN(n2722) );
  NAND4_X1 U3391 ( .A1(n2725), .A2(n2724), .A3(n2723), .A4(n2722), .ZN(n3883)
         );
  AOI21_X1 U3392 ( .B1(n3704), .B2(n3883), .A(n2726), .ZN(n2728) );
  NAND2_X1 U3393 ( .A1(n4327), .A2(n3885), .ZN(n2727) );
  OAI211_X1 U3394 ( .C1(n3684), .C2(n2857), .A(n2728), .B(n2727), .ZN(n2729)
         );
  AOI21_X1 U3395 ( .B1(n3710), .B2(n2837), .A(n2729), .ZN(n2730) );
  OAI21_X1 U3396 ( .B1(n2731), .B2(n3712), .A(n2730), .ZN(U3224) );
  NAND2_X1 U3397 ( .A1(n2598), .A2(n2841), .ZN(n3789) );
  AND2_X1 U3398 ( .A1(n3787), .A2(n3789), .ZN(n4480) );
  INV_X1 U3399 ( .A(n2732), .ZN(n2733) );
  NOR2_X1 U3400 ( .A1(n2734), .A2(n2733), .ZN(n2736) );
  NAND4_X1 U3401 ( .A1(n2738), .A2(n2737), .A3(n2736), .A4(n2735), .ZN(n2739)
         );
  OR2_X1 U3402 ( .A1(n2740), .A2(n3950), .ZN(n2817) );
  INV_X1 U3403 ( .A(n2817), .ZN(n2741) );
  INV_X1 U3404 ( .A(n4459), .ZN(n2853) );
  AOI21_X1 U3405 ( .B1(n4190), .B2(n3219), .A(n4480), .ZN(n2743) );
  AOI21_X1 U3406 ( .B1(n4169), .B2(n3888), .A(n2743), .ZN(n4479) );
  OAI21_X1 U3407 ( .B1(n2744), .B2(n4478), .A(n4479), .ZN(n2745) );
  AOI22_X1 U3408 ( .A1(n2745), .A2(n4350), .B1(REG3_REG_0__SCAN_IN), .B2(n4457), .ZN(n2747) );
  NAND2_X1 U3409 ( .A1(n4465), .A2(REG2_REG_0__SCAN_IN), .ZN(n2746) );
  OAI211_X1 U3410 ( .C1(n4480), .C2(n2853), .A(n2747), .B(n2746), .ZN(U3290)
         );
  INV_X1 U3411 ( .A(n2749), .ZN(n2750) );
  AOI21_X1 U3412 ( .B1(n2748), .B2(n2751), .A(n2750), .ZN(n2756) );
  OAI22_X1 U3413 ( .A1(n2804), .A2(n4335), .B1(n3683), .B2(n2596), .ZN(n2753)
         );
  NOR2_X1 U3414 ( .A1(n3684), .A2(n2757), .ZN(n2752) );
  AOI211_X1 U3415 ( .C1(REG3_REG_2__SCAN_IN), .C2(n2754), .A(n2753), .B(n2752), 
        .ZN(n2755) );
  OAI21_X1 U3416 ( .B1(n2756), .B2(n3712), .A(n2755), .ZN(U3234) );
  NAND2_X1 U3417 ( .A1(n2763), .A2(n2757), .ZN(n2758) );
  OR2_X1 U3418 ( .A1(n3886), .A2(n2803), .ZN(n3797) );
  NAND2_X1 U3419 ( .A1(n3886), .A2(n2803), .ZN(n3794) );
  XNOR2_X1 U3420 ( .A(n2802), .B(n2158), .ZN(n4488) );
  NAND2_X1 U3421 ( .A1(n2760), .A2(n3792), .ZN(n2799) );
  XNOR2_X1 U3422 ( .A(n2799), .B(n2158), .ZN(n2765) );
  AOI22_X1 U3423 ( .A1(n3885), .A2(n4169), .B1(n4217), .B2(n2761), .ZN(n2762)
         );
  OAI21_X1 U3424 ( .B1(n2763), .B2(n4172), .A(n2762), .ZN(n2764) );
  AOI21_X1 U3425 ( .B1(n2765), .B2(n4175), .A(n2764), .ZN(n2766) );
  OAI21_X1 U3426 ( .B1(n4488), .B2(n3219), .A(n2766), .ZN(n4489) );
  NAND2_X1 U3427 ( .A1(n4489), .A2(n4350), .ZN(n2771) );
  AOI21_X1 U3429 ( .B1(n2761), .B2(n2767), .A(n4858), .ZN(n4491) );
  OAI22_X1 U3430 ( .A1(n4350), .A2(n2768), .B1(n4197), .B2(REG3_REG_3__SCAN_IN), .ZN(n2769) );
  AOI21_X1 U3431 ( .B1(n4461), .B2(n4491), .A(n2769), .ZN(n2770) );
  OAI211_X1 U3432 ( .C1(n4488), .C2(n2853), .A(n2771), .B(n2770), .ZN(U3287)
         );
  INV_X1 U3433 ( .A(n2774), .ZN(n2776) );
  NAND2_X1 U3434 ( .A1(n2776), .A2(n2775), .ZN(n2884) );
  NAND2_X1 U3435 ( .A1(n2887), .A2(n2884), .ZN(n3006) );
  NAND2_X1 U3436 ( .A1(n3883), .A2(n3561), .ZN(n2778) );
  MUX2_X1 U3437 ( .A(n4322), .B(DATAI_6_), .S(n3734), .Z(n2926) );
  INV_X1 U3438 ( .A(n2926), .ZN(n2863) );
  OR2_X1 U3439 ( .A1(n3577), .A2(n2863), .ZN(n2777) );
  NAND2_X1 U3440 ( .A1(n2778), .A2(n2777), .ZN(n2779) );
  XNOR2_X1 U3441 ( .A(n2779), .B(n3578), .ZN(n2784) );
  INV_X1 U3442 ( .A(n2784), .ZN(n2782) );
  INV_X1 U3443 ( .A(n3883), .ZN(n2780) );
  OAI22_X1 U3444 ( .A1(n2780), .A2(n3531), .B1(n2863), .B2(n3576), .ZN(n2783)
         );
  INV_X1 U3445 ( .A(n2783), .ZN(n2781) );
  INV_X1 U3446 ( .A(n3007), .ZN(n2890) );
  AND2_X1 U3447 ( .A1(n2784), .A2(n2783), .ZN(n3005) );
  NOR2_X1 U3448 ( .A1(n2890), .A2(n3005), .ZN(n2785) );
  XNOR2_X1 U3449 ( .A(n3006), .B(n2785), .ZN(n2797) );
  NAND2_X1 U3450 ( .A1(n3400), .A2(REG1_REG_7__SCAN_IN), .ZN(n2791) );
  OR2_X1 U3451 ( .A1(n2786), .A2(REG3_REG_7__SCAN_IN), .ZN(n2787) );
  AND2_X1 U3452 ( .A1(n2903), .A2(n2787), .ZN(n3015) );
  NAND2_X1 U3453 ( .A1(n3412), .A2(n3015), .ZN(n2790) );
  NAND2_X1 U3454 ( .A1(n3445), .A2(REG0_REG_7__SCAN_IN), .ZN(n2789) );
  NAND2_X1 U3455 ( .A1(n3725), .A2(REG2_REG_7__SCAN_IN), .ZN(n2788) );
  AOI21_X1 U3456 ( .B1(n3704), .B2(n3882), .A(n2792), .ZN(n2794) );
  NAND2_X1 U3457 ( .A1(n4327), .A2(n3884), .ZN(n2793) );
  OAI211_X1 U34580 ( .C1(n3684), .C2(n2863), .A(n2794), .B(n2793), .ZN(n2795)
         );
  AOI21_X1 U34590 ( .B1(n3710), .B2(n4450), .A(n2795), .ZN(n2796) );
  OAI21_X1 U3460 ( .B1(n2797), .B2(n3712), .A(n2796), .ZN(U3236) );
  NAND2_X1 U3461 ( .A1(n2798), .A2(n2823), .ZN(n2836) );
  OAI211_X1 U3462 ( .C1(n4858), .C2(n2823), .A(n2836), .B(n4510), .ZN(n4493)
         );
  NOR2_X1 U3463 ( .A1(n4493), .A2(n4316), .ZN(n2812) );
  NAND2_X1 U3464 ( .A1(n3885), .A2(n2823), .ZN(n3800) );
  NAND2_X1 U3465 ( .A1(n3798), .A2(n3800), .ZN(n2820) );
  NAND2_X1 U3466 ( .A1(n2799), .A2(n2158), .ZN(n2800) );
  NAND2_X1 U34670 ( .A1(n2800), .A2(n3797), .ZN(n2829) );
  XNOR2_X1 U3468 ( .A(n2820), .B(n2829), .ZN(n2811) );
  OAI22_X1 U34690 ( .A1(n2804), .A2(n4172), .B1(n2823), .B2(n4207), .ZN(n2809)
         );
  NAND2_X1 U3470 ( .A1(n3886), .A2(n2761), .ZN(n2801) );
  NAND2_X1 U34710 ( .A1(n2802), .A2(n2801), .ZN(n2822) );
  NAND2_X1 U3472 ( .A1(n2804), .A2(n2803), .ZN(n2819) );
  NAND2_X1 U34730 ( .A1(n2822), .A2(n2819), .ZN(n2805) );
  INV_X1 U3474 ( .A(n2820), .ZN(n3776) );
  OR2_X1 U34750 ( .A1(n2805), .A2(n3776), .ZN(n2807) );
  NAND2_X1 U3476 ( .A1(n2805), .A2(n3776), .ZN(n2806) );
  NAND2_X1 U34770 ( .A1(n2807), .A2(n2806), .ZN(n2814) );
  NOR2_X1 U3478 ( .A1(n2814), .A2(n3219), .ZN(n2808) );
  AOI211_X1 U34790 ( .C1(n4169), .C2(n3884), .A(n2809), .B(n2808), .ZN(n2810)
         );
  OAI21_X1 U3480 ( .B1(n4190), .B2(n2811), .A(n2810), .ZN(n4494) );
  AOI211_X1 U34810 ( .C1(n4457), .C2(n2813), .A(n2812), .B(n4494), .ZN(n2816)
         );
  INV_X1 U3482 ( .A(n2814), .ZN(n4496) );
  AOI22_X1 U34830 ( .A1(n4496), .A2(n4459), .B1(REG2_REG_4__SCAN_IN), .B2(
        n4465), .ZN(n2815) );
  OAI21_X1 U3484 ( .B1(n2816), .B2(n4465), .A(n2815), .ZN(U3286) );
  NAND2_X1 U34850 ( .A1(n3219), .A2(n2817), .ZN(n2818) );
  AND2_X1 U3486 ( .A1(n2820), .A2(n2819), .ZN(n2821) );
  NAND2_X1 U34870 ( .A1(n2822), .A2(n2821), .ZN(n2826) );
  INV_X1 U3488 ( .A(n2823), .ZN(n2824) );
  NAND2_X1 U34890 ( .A1(n3885), .A2(n2824), .ZN(n2825) );
  NAND2_X1 U3490 ( .A1(n2826), .A2(n2825), .ZN(n2859) );
  AND2_X1 U34910 ( .A1(n3884), .A2(n2857), .ZN(n3801) );
  INV_X1 U3492 ( .A(n3801), .ZN(n2827) );
  OR2_X1 U34930 ( .A1(n3884), .A2(n2857), .ZN(n3814) );
  NAND2_X1 U3494 ( .A1(n2827), .A2(n3814), .ZN(n3772) );
  XNOR2_X1 U34950 ( .A(n2859), .B(n3772), .ZN(n4498) );
  INV_X1 U3496 ( .A(n3798), .ZN(n2828) );
  OR2_X1 U34970 ( .A1(n2829), .A2(n2828), .ZN(n2830) );
  NAND2_X1 U3498 ( .A1(n2830), .A2(n3800), .ZN(n2864) );
  XNOR2_X1 U34990 ( .A(n2864), .B(n3772), .ZN(n2834) );
  AOI22_X1 U3500 ( .A1(n3883), .A2(n4169), .B1(n4217), .B2(n2860), .ZN(n2831)
         );
  OAI21_X1 U35010 ( .B1(n2832), .B2(n4172), .A(n2831), .ZN(n2833) );
  AOI21_X1 U3502 ( .B1(n2834), .B2(n4175), .A(n2833), .ZN(n4499) );
  MUX2_X1 U35030 ( .A(n4499), .B(n2835), .S(n4465), .Z(n2839) );
  AOI21_X1 U3504 ( .B1(n2860), .B2(n2836), .A(n2189), .ZN(n4502) );
  AOI22_X1 U35050 ( .A1(n4461), .A2(n4502), .B1(n2837), .B2(n4457), .ZN(n2838)
         );
  OAI211_X1 U35060 ( .C1(n4203), .C2(n4498), .A(n2839), .B(n2838), .ZN(U3285)
         );
  OAI21_X1 U35070 ( .B1(n2841), .B2(n2846), .A(n2840), .ZN(n4482) );
  OAI21_X1 U35080 ( .B1(n2616), .B2(n2843), .A(n2842), .ZN(n4483) );
  NAND2_X1 U35090 ( .A1(n2598), .A2(n4188), .ZN(n2845) );
  NAND2_X1 U35100 ( .A1(n3887), .A2(n4169), .ZN(n2844) );
  OAI211_X1 U35110 ( .C1(n4207), .C2(n2846), .A(n2845), .B(n2844), .ZN(n2847)
         );
  INV_X1 U35120 ( .A(n2847), .ZN(n2850) );
  XNOR2_X1 U35130 ( .A(n2616), .B(n3787), .ZN(n2848) );
  NAND2_X1 U35140 ( .A1(n2848), .A2(n4175), .ZN(n2849) );
  OAI211_X1 U35150 ( .C1(n4483), .C2(n3219), .A(n2850), .B(n2849), .ZN(n4485)
         );
  INV_X1 U35160 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2852) );
  INV_X1 U35170 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2851) );
  OAI22_X1 U35180 ( .A1(n4350), .A2(n2852), .B1(n2851), .B2(n4197), .ZN(n2855)
         );
  NOR2_X1 U35190 ( .A1(n2853), .A2(n4483), .ZN(n2854) );
  AOI211_X1 U35200 ( .C1(n4350), .C2(n4485), .A(n2855), .B(n2854), .ZN(n2856)
         );
  OAI21_X1 U35210 ( .B1(n4195), .B2(n4482), .A(n2856), .ZN(U3289) );
  NAND2_X1 U35220 ( .A1(n2867), .A2(n2857), .ZN(n2858) );
  NAND2_X1 U35230 ( .A1(n2859), .A2(n2858), .ZN(n2862) );
  NAND2_X1 U35240 ( .A1(n3884), .A2(n2860), .ZN(n2861) );
  NAND2_X1 U35250 ( .A1(n3883), .A2(n2863), .ZN(n2915) );
  INV_X1 U35260 ( .A(n2915), .ZN(n3817) );
  NOR2_X1 U35270 ( .A1(n3883), .A2(n2863), .ZN(n3804) );
  OR2_X1 U35280 ( .A1(n3817), .A2(n3804), .ZN(n3769) );
  XNOR2_X1 U35290 ( .A(n2928), .B(n3769), .ZN(n4451) );
  OR2_X1 U35300 ( .A1(n2864), .A2(n3801), .ZN(n2865) );
  NAND2_X1 U35310 ( .A1(n2865), .A2(n3814), .ZN(n2916) );
  XOR2_X1 U35320 ( .A(n3769), .B(n2916), .Z(n2870) );
  AOI22_X1 U35330 ( .A1(n3882), .A2(n4169), .B1(n4217), .B2(n2926), .ZN(n2866)
         );
  OAI21_X1 U35340 ( .B1(n2867), .B2(n4172), .A(n2866), .ZN(n2869) );
  NOR2_X1 U35350 ( .A1(n4451), .A2(n3219), .ZN(n2868) );
  AOI211_X1 U35360 ( .C1(n2870), .C2(n4175), .A(n2869), .B(n2868), .ZN(n4456)
         );
  OAI21_X1 U35370 ( .B1(n4487), .B2(n4451), .A(n4456), .ZN(n2875) );
  NAND2_X1 U35380 ( .A1(n2875), .A2(n4537), .ZN(n2874) );
  NAND2_X1 U35390 ( .A1(n2871), .A2(n2926), .ZN(n2872) );
  AND2_X1 U35400 ( .A1(n2921), .A2(n2872), .ZN(n4452) );
  NAND2_X1 U35410 ( .A1(n4215), .A2(n4452), .ZN(n2873) );
  OAI211_X1 U35420 ( .C1(n4537), .C2(n2438), .A(n2874), .B(n2873), .ZN(U3524)
         );
  INV_X1 U35430 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2878) );
  NAND2_X1 U35440 ( .A1(n2875), .A2(n4524), .ZN(n2877) );
  NAND2_X1 U35450 ( .A1(n4276), .A2(n4452), .ZN(n2876) );
  OAI211_X1 U35460 ( .C1(n4524), .C2(n2878), .A(n2877), .B(n2876), .ZN(U3479)
         );
  XNOR2_X1 U35470 ( .A(n2903), .B(REG3_REG_8__SCAN_IN), .ZN(n2967) );
  INV_X1 U35480 ( .A(n2967), .ZN(n2914) );
  NAND2_X1 U35490 ( .A1(n3882), .A2(n3561), .ZN(n2882) );
  INV_X1 U35500 ( .A(DATAI_7_), .ZN(n2879) );
  MUX2_X1 U35510 ( .A(n2880), .B(n2879), .S(n3734), .Z(n3004) );
  OR2_X1 U35520 ( .A1(n3577), .A2(n3004), .ZN(n2881) );
  NAND2_X1 U35530 ( .A1(n2882), .A2(n2881), .ZN(n2883) );
  XNOR2_X1 U35540 ( .A(n2883), .B(n3578), .ZN(n2889) );
  INV_X1 U35550 ( .A(n3882), .ZN(n2899) );
  OAI22_X1 U35560 ( .A1(n2899), .A2(n3531), .B1(n3576), .B2(n3004), .ZN(n2888)
         );
  AND2_X1 U35570 ( .A1(n2889), .A2(n2888), .ZN(n2891) );
  NOR2_X1 U35580 ( .A1(n3005), .A2(n2891), .ZN(n2885) );
  AND2_X1 U35590 ( .A1(n2885), .A2(n2884), .ZN(n2886) );
  XNOR2_X1 U35600 ( .A(n2889), .B(n2888), .ZN(n3012) );
  NOR2_X1 U35610 ( .A1(n2891), .A2(n3008), .ZN(n2979) );
  NOR2_X1 U35620 ( .A1(n2981), .A2(n2979), .ZN(n2976) );
  AOI22_X1 U35630 ( .A1(n3400), .A2(REG1_REG_8__SCAN_IN), .B1(n3445), .B2(
        REG0_REG_8__SCAN_IN), .ZN(n2893) );
  AOI22_X1 U35640 ( .A1(n3412), .A2(n2967), .B1(n3725), .B2(
        REG2_REG_8__SCAN_IN), .ZN(n2892) );
  INV_X1 U35650 ( .A(DATAI_8_), .ZN(n2894) );
  MUX2_X1 U35660 ( .A(n2895), .B(n2894), .S(n3734), .Z(n2963) );
  OAI22_X1 U35670 ( .A1(n2951), .A2(n2572), .B1(n2963), .B2(n3577), .ZN(n2896)
         );
  XNOR2_X1 U35680 ( .A(n2896), .B(n3578), .ZN(n2975) );
  OAI22_X1 U35690 ( .A1(n2951), .A2(n3531), .B1(n2963), .B2(n3576), .ZN(n2977)
         );
  XNOR2_X1 U35700 ( .A(n2975), .B(n2977), .ZN(n2897) );
  XNOR2_X1 U35710 ( .A(n2976), .B(n2897), .ZN(n2898) );
  NAND2_X1 U35720 ( .A1(n2898), .A2(n4337), .ZN(n2913) );
  OAI22_X1 U35730 ( .A1(n3684), .A2(n2963), .B1(n2899), .B2(n3683), .ZN(n2911)
         );
  NAND2_X1 U35740 ( .A1(n2608), .A2(REG1_REG_9__SCAN_IN), .ZN(n2908) );
  INV_X1 U35750 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2901) );
  INV_X1 U35760 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2900) );
  OAI21_X1 U35770 ( .B1(n2903), .B2(n2901), .A(n2900), .ZN(n2904) );
  NAND2_X1 U35780 ( .A1(REG3_REG_8__SCAN_IN), .A2(REG3_REG_9__SCAN_IN), .ZN(
        n2902) );
  AND2_X1 U35790 ( .A1(n2904), .A2(n2937), .ZN(n2990) );
  NAND2_X1 U35800 ( .A1(n3412), .A2(n2990), .ZN(n2907) );
  NAND2_X1 U35810 ( .A1(n3445), .A2(REG0_REG_9__SCAN_IN), .ZN(n2906) );
  NAND2_X1 U3582 ( .A1(n3725), .A2(REG2_REG_9__SCAN_IN), .ZN(n2905) );
  NAND4_X1 U3583 ( .A1(n2908), .A2(n2907), .A3(n2906), .A4(n2905), .ZN(n3880)
         );
  INV_X1 U3584 ( .A(n3880), .ZN(n3056) );
  OAI21_X1 U3585 ( .B1(n4335), .B2(n3056), .A(n2909), .ZN(n2910) );
  NOR2_X1 U3586 ( .A1(n2911), .A2(n2910), .ZN(n2912) );
  OAI211_X1 U3587 ( .C1(n4342), .C2(n2914), .A(n2913), .B(n2912), .ZN(U3218)
         );
  OAI22_X1 U3588 ( .A1(n2951), .A2(n4185), .B1(n3004), .B2(n4207), .ZN(n2919)
         );
  OR2_X1 U3589 ( .A1(n3882), .A2(n3004), .ZN(n3803) );
  NAND2_X1 U3590 ( .A1(n3882), .A2(n3004), .ZN(n3809) );
  NAND2_X1 U3591 ( .A1(n3803), .A2(n3809), .ZN(n3773) );
  XNOR2_X1 U3592 ( .A(n2932), .B(n2321), .ZN(n2917) );
  NOR2_X1 U3593 ( .A1(n2917), .A2(n4190), .ZN(n2918) );
  AOI211_X1 U3594 ( .C1(n4188), .C2(n3883), .A(n2919), .B(n2918), .ZN(n4506)
         );
  NAND2_X1 U3595 ( .A1(n2921), .A2(n2950), .ZN(n2920) );
  NAND2_X1 U3596 ( .A1(n2920), .A2(n4510), .ZN(n2922) );
  OR2_X1 U3597 ( .A1(n2922), .A2(n2964), .ZN(n4505) );
  INV_X1 U3598 ( .A(n4505), .ZN(n2925) );
  INV_X1 U3599 ( .A(n3015), .ZN(n2923) );
  OAI22_X1 U3600 ( .A1(n4350), .A2(n2473), .B1(n2923), .B2(n4197), .ZN(n2924)
         );
  AOI21_X1 U3601 ( .B1(n2925), .B2(n4179), .A(n2924), .ZN(n2931) );
  AND2_X1 U3602 ( .A1(n3883), .A2(n2926), .ZN(n2927) );
  NAND2_X1 U3603 ( .A1(n2929), .A2(n2321), .ZN(n4503) );
  NAND3_X1 U3604 ( .A1(n3051), .A2(n4503), .A3(n4107), .ZN(n2930) );
  OAI211_X1 U3605 ( .C1(n4506), .C2(n4465), .A(n2931), .B(n2930), .ZN(U3283)
         );
  NAND2_X1 U3606 ( .A1(n2932), .A2(n3803), .ZN(n2933) );
  NAND2_X1 U3607 ( .A1(n2933), .A2(n3809), .ZN(n2958) );
  OR2_X1 U3608 ( .A1(n3881), .A2(n2963), .ZN(n3810) );
  NAND2_X1 U3609 ( .A1(n2958), .A2(n3810), .ZN(n2934) );
  NAND2_X1 U3610 ( .A1(n3881), .A2(n2963), .ZN(n3808) );
  NAND2_X1 U3611 ( .A1(n2934), .A2(n3808), .ZN(n3041) );
  MUX2_X1 U3612 ( .A(n2935), .B(DATAI_9_), .S(n3734), .Z(n3047) );
  AND2_X1 U3613 ( .A1(n3880), .A2(n3055), .ZN(n3815) );
  INV_X1 U3614 ( .A(n3815), .ZN(n2936) );
  OR2_X1 U3615 ( .A1(n3880), .A2(n3055), .ZN(n3811) );
  NAND2_X1 U3616 ( .A1(n2936), .A2(n3811), .ZN(n3768) );
  XNOR2_X1 U3617 ( .A(n3041), .B(n3768), .ZN(n2945) );
  NAND2_X1 U3618 ( .A1(n2608), .A2(REG1_REG_10__SCAN_IN), .ZN(n2942) );
  AND2_X1 U3619 ( .A1(n2937), .A2(n4831), .ZN(n2938) );
  NOR2_X1 U3620 ( .A1(n3029), .A2(n2938), .ZN(n3065) );
  NAND2_X1 U3621 ( .A1(n3412), .A2(n3065), .ZN(n2941) );
  NAND2_X1 U3622 ( .A1(n3445), .A2(REG0_REG_10__SCAN_IN), .ZN(n2940) );
  NAND2_X1 U3623 ( .A1(n3725), .A2(REG2_REG_10__SCAN_IN), .ZN(n2939) );
  NAND4_X1 U3624 ( .A1(n2942), .A2(n2941), .A3(n2940), .A4(n2939), .ZN(n3879)
         );
  AOI22_X1 U3625 ( .A1(n3879), .A2(n4169), .B1(n4217), .B2(n3047), .ZN(n2943)
         );
  OAI21_X1 U3626 ( .B1(n2951), .B2(n4172), .A(n2943), .ZN(n2944) );
  AOI21_X1 U3627 ( .B1(n2945), .B2(n4175), .A(n2944), .ZN(n4513) );
  NAND2_X1 U3628 ( .A1(n2966), .A2(n3047), .ZN(n2946) );
  AND2_X1 U3629 ( .A1(n3062), .A2(n2946), .ZN(n4511) );
  INV_X1 U3630 ( .A(n2990), .ZN(n2947) );
  OAI22_X1 U3631 ( .A1(n4350), .A2(n2948), .B1(n2947), .B2(n4197), .ZN(n2949)
         );
  AOI21_X1 U3632 ( .B1(n4511), .B2(n4461), .A(n2949), .ZN(n2957) );
  NAND2_X1 U3633 ( .A1(n3882), .A2(n2950), .ZN(n3049) );
  NAND2_X1 U3634 ( .A1(n3051), .A2(n3049), .ZN(n2962) );
  NAND2_X1 U3635 ( .A1(n2951), .A2(n2963), .ZN(n3053) );
  NAND2_X1 U3636 ( .A1(n2962), .A2(n3053), .ZN(n2953) );
  INV_X1 U3637 ( .A(n2963), .ZN(n2952) );
  NAND2_X1 U3638 ( .A1(n3881), .A2(n2952), .ZN(n3048) );
  NAND2_X1 U3639 ( .A1(n2953), .A2(n3048), .ZN(n2955) );
  INV_X1 U3640 ( .A(n3768), .ZN(n2954) );
  XNOR2_X1 U3641 ( .A(n2955), .B(n2954), .ZN(n4509) );
  NAND2_X1 U3642 ( .A1(n4509), .A2(n4107), .ZN(n2956) );
  OAI211_X1 U3643 ( .C1(n4513), .C2(n4465), .A(n2957), .B(n2956), .ZN(U3281)
         );
  NAND2_X1 U3644 ( .A1(n3810), .A2(n3808), .ZN(n3771) );
  XOR2_X1 U3645 ( .A(n3771), .B(n2958), .Z(n2961) );
  OAI22_X1 U3646 ( .A1(n3056), .A2(n4185), .B1(n4207), .B2(n2963), .ZN(n2959)
         );
  AOI21_X1 U3647 ( .B1(n4188), .B2(n3882), .A(n2959), .ZN(n2960) );
  OAI21_X1 U3648 ( .B1(n2961), .B2(n4190), .A(n2960), .ZN(n2993) );
  INV_X1 U3649 ( .A(n2993), .ZN(n2971) );
  XOR2_X1 U3650 ( .A(n3771), .B(n2962), .Z(n2994) );
  OR2_X1 U3651 ( .A1(n2964), .A2(n2963), .ZN(n2965) );
  NAND2_X1 U3652 ( .A1(n2966), .A2(n2965), .ZN(n3000) );
  AOI22_X1 U3653 ( .A1(n4465), .A2(REG2_REG_8__SCAN_IN), .B1(n2967), .B2(n4457), .ZN(n2968) );
  OAI21_X1 U3654 ( .B1(n4195), .B2(n3000), .A(n2968), .ZN(n2969) );
  AOI21_X1 U3655 ( .B1(n2994), .B2(n4107), .A(n2969), .ZN(n2970) );
  OAI21_X1 U3656 ( .B1(n2971), .B2(n4465), .A(n2970), .ZN(U3282) );
  NAND2_X1 U3657 ( .A1(n3880), .A2(n3561), .ZN(n2973) );
  OR2_X1 U3658 ( .A1(n3577), .A2(n3055), .ZN(n2972) );
  NAND2_X1 U3659 ( .A1(n2973), .A2(n2972), .ZN(n2974) );
  XNOR2_X1 U3660 ( .A(n2974), .B(n3578), .ZN(n3020) );
  OAI22_X1 U3661 ( .A1(n3056), .A2(n3531), .B1(n3055), .B2(n3576), .ZN(n3021)
         );
  XNOR2_X1 U3662 ( .A(n3020), .B(n3021), .ZN(n2986) );
  INV_X1 U3663 ( .A(n2977), .ZN(n2978) );
  OR2_X1 U3664 ( .A1(n2979), .A2(n2978), .ZN(n2980) );
  INV_X1 U3665 ( .A(n3025), .ZN(n2985) );
  AOI21_X1 U3666 ( .B1(n2986), .B2(n2983), .A(n2985), .ZN(n2992) );
  AND2_X1 U3667 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4372) );
  AOI21_X1 U3668 ( .B1(n3704), .B2(n3879), .A(n4372), .ZN(n2988) );
  NAND2_X1 U3669 ( .A1(n4327), .A2(n3881), .ZN(n2987) );
  OAI211_X1 U3670 ( .C1(n3684), .C2(n3055), .A(n2988), .B(n2987), .ZN(n2989)
         );
  AOI21_X1 U3671 ( .B1(n3710), .B2(n2990), .A(n2989), .ZN(n2991) );
  OAI21_X1 U3672 ( .B1(n2992), .B2(n3712), .A(n2991), .ZN(U3228) );
  INV_X1 U3673 ( .A(REG0_REG_8__SCAN_IN), .ZN(n2995) );
  AOI21_X1 U3674 ( .B1(n2994), .B2(n4508), .A(n2993), .ZN(n2997) );
  MUX2_X1 U3675 ( .A(n2995), .B(n2997), .S(n4524), .Z(n2996) );
  OAI21_X1 U3676 ( .B1(n3000), .B2(n4310), .A(n2996), .ZN(U3483) );
  MUX2_X1 U3677 ( .A(n2998), .B(n2997), .S(n4537), .Z(n2999) );
  OAI21_X1 U3678 ( .B1(n3000), .B2(n4264), .A(n2999), .ZN(U3526) );
  AOI21_X1 U3679 ( .B1(n4327), .B2(n3883), .A(n3001), .ZN(n3003) );
  NAND2_X1 U3680 ( .A1(n3704), .A2(n3881), .ZN(n3002) );
  OAI211_X1 U3681 ( .C1(n3684), .C2(n3004), .A(n3003), .B(n3002), .ZN(n3014)
         );
  OR2_X1 U3682 ( .A1(n3006), .A2(n3005), .ZN(n3009) );
  NAND2_X1 U3683 ( .A1(n3009), .A2(n3007), .ZN(n3011) );
  AND2_X1 U3684 ( .A1(n3009), .A2(n3008), .ZN(n3010) );
  AOI211_X1 U3685 ( .C1(n3012), .C2(n3011), .A(n3712), .B(n3010), .ZN(n3013)
         );
  AOI211_X1 U3686 ( .C1(n3015), .C2(n3710), .A(n3014), .B(n3013), .ZN(n3016)
         );
  INV_X1 U3687 ( .A(n3016), .ZN(U3210) );
  NAND2_X1 U3688 ( .A1(n3879), .A2(n3561), .ZN(n3018) );
  MUX2_X1 U3689 ( .A(n4319), .B(DATAI_10_), .S(n3734), .Z(n3098) );
  OR2_X1 U3690 ( .A1(n3577), .A2(n3099), .ZN(n3017) );
  NAND2_X1 U3691 ( .A1(n3018), .A2(n3017), .ZN(n3019) );
  XNOR2_X1 U3692 ( .A(n3019), .B(n3571), .ZN(n3080) );
  INV_X1 U3693 ( .A(n3879), .ZN(n3100) );
  OAI22_X1 U3694 ( .A1(n3100), .A2(n3531), .B1(n3576), .B2(n3099), .ZN(n3081)
         );
  XNOR2_X1 U3695 ( .A(n3080), .B(n3081), .ZN(n3026) );
  INV_X1 U3696 ( .A(n3020), .ZN(n3023) );
  INV_X1 U3697 ( .A(n3021), .ZN(n3022) );
  NAND2_X1 U3698 ( .A1(n3023), .A2(n3022), .ZN(n3027) );
  AND2_X1 U3699 ( .A1(n3026), .A2(n3027), .ZN(n3024) );
  NAND2_X1 U3700 ( .A1(n3025), .A2(n3024), .ZN(n3084) );
  NAND2_X1 U3701 ( .A1(n3084), .A2(n4337), .ZN(n3040) );
  AOI21_X1 U3702 ( .B1(n3025), .B2(n3027), .A(n3026), .ZN(n3039) );
  AOI21_X1 U3703 ( .B1(n4327), .B2(n3880), .A(n3028), .ZN(n3036) );
  NAND2_X1 U3704 ( .A1(n3400), .A2(REG1_REG_11__SCAN_IN), .ZN(n3034) );
  NOR2_X1 U3705 ( .A1(n3029), .A2(REG3_REG_11__SCAN_IN), .ZN(n3030) );
  NOR2_X1 U3706 ( .A1(n3087), .A2(n3030), .ZN(n3113) );
  NAND2_X1 U3707 ( .A1(n3412), .A2(n3113), .ZN(n3033) );
  NAND2_X1 U3708 ( .A1(n3445), .A2(REG0_REG_11__SCAN_IN), .ZN(n3032) );
  NAND2_X1 U3709 ( .A1(n3725), .A2(REG2_REG_11__SCAN_IN), .ZN(n3031) );
  NAND4_X1 U3710 ( .A1(n3034), .A2(n3033), .A3(n3032), .A4(n3031), .ZN(n3878)
         );
  NAND2_X1 U3711 ( .A1(n3704), .A2(n3878), .ZN(n3035) );
  OAI211_X1 U3712 ( .C1(n3684), .C2(n3099), .A(n3036), .B(n3035), .ZN(n3037)
         );
  AOI21_X1 U3713 ( .B1(n3710), .B2(n3065), .A(n3037), .ZN(n3038) );
  OAI21_X1 U3714 ( .B1(n3040), .B2(n3039), .A(n3038), .ZN(U3214) );
  NOR2_X1 U3715 ( .A1(n3879), .A2(n3099), .ZN(n3818) );
  NAND2_X1 U3716 ( .A1(n3879), .A2(n3099), .ZN(n3096) );
  INV_X1 U3717 ( .A(n3096), .ZN(n3824) );
  OR2_X1 U3718 ( .A1(n3818), .A2(n3824), .ZN(n3061) );
  INV_X1 U3719 ( .A(n3061), .ZN(n3763) );
  XNOR2_X1 U3720 ( .A(n3097), .B(n3763), .ZN(n3046) );
  NAND2_X1 U3721 ( .A1(n3880), .A2(n4188), .ZN(n3044) );
  NAND2_X1 U3722 ( .A1(n3878), .A2(n4169), .ZN(n3043) );
  OAI211_X1 U3723 ( .C1(n4207), .C2(n3099), .A(n3044), .B(n3043), .ZN(n3045)
         );
  AOI21_X1 U3724 ( .B1(n3046), .B2(n4175), .A(n3045), .ZN(n3119) );
  AND2_X1 U3725 ( .A1(n2169), .A2(n3048), .ZN(n3052) );
  AND2_X1 U3726 ( .A1(n3049), .A2(n3052), .ZN(n3050) );
  NAND2_X1 U3727 ( .A1(n3051), .A2(n3050), .ZN(n3060) );
  INV_X1 U3728 ( .A(n3052), .ZN(n3054) );
  OR2_X1 U3729 ( .A1(n3054), .A2(n3053), .ZN(n3058) );
  NAND2_X1 U3730 ( .A1(n3056), .A2(n3055), .ZN(n3057) );
  AND2_X1 U3731 ( .A1(n3058), .A2(n3057), .ZN(n3059) );
  NAND2_X1 U3732 ( .A1(n3060), .A2(n3059), .ZN(n3102) );
  XNOR2_X1 U3733 ( .A(n3102), .B(n3061), .ZN(n3118) );
  INV_X1 U3734 ( .A(n3062), .ZN(n3064) );
  INV_X1 U3735 ( .A(n3111), .ZN(n3063) );
  OAI21_X1 U3736 ( .B1(n3064), .B2(n3099), .A(n3063), .ZN(n3126) );
  AOI22_X1 U3737 ( .A1(n4465), .A2(REG2_REG_10__SCAN_IN), .B1(n3065), .B2(
        n4457), .ZN(n3066) );
  OAI21_X1 U3738 ( .B1(n3126), .B2(n4195), .A(n3066), .ZN(n3067) );
  AOI21_X1 U3739 ( .B1(n3118), .B2(n4107), .A(n3067), .ZN(n3068) );
  OAI21_X1 U3740 ( .B1(n3119), .B2(n4465), .A(n3068), .ZN(U3280) );
  NAND2_X1 U3741 ( .A1(n3878), .A2(n3561), .ZN(n3073) );
  OAI21_X1 U3742 ( .B1(n3168), .B2(IR_REG_10__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n3069) );
  OR2_X1 U3743 ( .A1(n3069), .A2(n4737), .ZN(n3070) );
  NAND2_X1 U3744 ( .A1(n3069), .A2(n4737), .ZN(n3127) );
  INV_X1 U3745 ( .A(DATAI_11_), .ZN(n3071) );
  MUX2_X1 U3746 ( .A(n4475), .B(n3071), .S(n3734), .Z(n3145) );
  OR2_X1 U3747 ( .A1(n3577), .A2(n3145), .ZN(n3072) );
  NAND2_X1 U3748 ( .A1(n3073), .A2(n3072), .ZN(n3074) );
  XNOR2_X1 U3749 ( .A(n3074), .B(n3571), .ZN(n3076) );
  NOR2_X1 U3750 ( .A1(n2572), .A2(n3145), .ZN(n3075) );
  AOI21_X1 U3751 ( .B1(n3566), .B2(n3878), .A(n3075), .ZN(n3077) );
  NAND2_X1 U3752 ( .A1(n3076), .A2(n3077), .ZN(n3151) );
  INV_X1 U3753 ( .A(n3076), .ZN(n3079) );
  INV_X1 U3754 ( .A(n3077), .ZN(n3078) );
  NAND2_X1 U3755 ( .A1(n3079), .A2(n3078), .ZN(n3153) );
  NAND2_X1 U3756 ( .A1(n3151), .A2(n3153), .ZN(n3085) );
  INV_X1 U3757 ( .A(n3080), .ZN(n3082) );
  NAND2_X1 U3758 ( .A1(n3082), .A2(n3081), .ZN(n3083) );
  NAND2_X1 U3759 ( .A1(n3084), .A2(n3083), .ZN(n3152) );
  XOR2_X1 U3760 ( .A(n3085), .B(n3152), .Z(n3095) );
  INV_X1 U3761 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3086) );
  NOR2_X1 U3762 ( .A1(STATE_REG_SCAN_IN), .A2(n3086), .ZN(n4382) );
  AOI21_X1 U3763 ( .B1(n4327), .B2(n3879), .A(n4382), .ZN(n3092) );
  AOI22_X1 U3764 ( .A1(n3400), .A2(REG1_REG_12__SCAN_IN), .B1(n3445), .B2(
        REG0_REG_12__SCAN_IN), .ZN(n3090) );
  OR2_X1 U3765 ( .A1(n3087), .A2(REG3_REG_12__SCAN_IN), .ZN(n3088) );
  AND2_X1 U3766 ( .A1(n3129), .A2(n3088), .ZN(n3141) );
  AOI22_X1 U3767 ( .A1(n3412), .A2(n3141), .B1(n3725), .B2(
        REG2_REG_12__SCAN_IN), .ZN(n3089) );
  NAND2_X1 U3768 ( .A1(n3704), .A2(n3877), .ZN(n3091) );
  OAI211_X1 U3769 ( .C1(n3684), .C2(n3145), .A(n3092), .B(n3091), .ZN(n3093)
         );
  AOI21_X1 U3770 ( .B1(n3710), .B2(n3113), .A(n3093), .ZN(n3094) );
  OAI21_X1 U3771 ( .B1(n3095), .B2(n3712), .A(n3094), .ZN(U3233) );
  OR2_X1 U3772 ( .A1(n3878), .A2(n3145), .ZN(n3241) );
  NAND2_X1 U3773 ( .A1(n3878), .A2(n3145), .ZN(n3238) );
  XNOR2_X1 U3774 ( .A(n3245), .B(n3778), .ZN(n3109) );
  OAI22_X1 U3775 ( .A1(n3215), .A2(n4185), .B1(n3145), .B2(n4207), .ZN(n3107)
         );
  NOR2_X1 U3776 ( .A1(n3879), .A2(n3098), .ZN(n3101) );
  OAI22_X1 U3777 ( .A1(n3102), .A2(n3101), .B1(n3100), .B2(n3099), .ZN(n3104)
         );
  NAND2_X1 U3778 ( .A1(n3104), .A2(n3778), .ZN(n3105) );
  AND2_X1 U3779 ( .A1(n3147), .A2(n3105), .ZN(n3110) );
  NOR2_X1 U3780 ( .A1(n3110), .A2(n3219), .ZN(n3106) );
  AOI211_X1 U3781 ( .C1(n4188), .C2(n3879), .A(n3107), .B(n3106), .ZN(n3108)
         );
  OAI21_X1 U3782 ( .B1(n4190), .B2(n3109), .A(n3108), .ZN(n4518) );
  INV_X1 U3783 ( .A(n4518), .ZN(n3117) );
  INV_X1 U3784 ( .A(n3110), .ZN(n4520) );
  NOR2_X1 U3785 ( .A1(n3111), .A2(n3145), .ZN(n3112) );
  OR2_X1 U3786 ( .A1(n3139), .A2(n3112), .ZN(n4517) );
  AOI22_X1 U3787 ( .A1(n4465), .A2(REG2_REG_11__SCAN_IN), .B1(n3113), .B2(
        n4457), .ZN(n3114) );
  OAI21_X1 U3788 ( .B1(n4517), .B2(n4195), .A(n3114), .ZN(n3115) );
  AOI21_X1 U3789 ( .B1(n4520), .B2(n4459), .A(n3115), .ZN(n3116) );
  OAI21_X1 U3790 ( .B1(n3117), .B2(n4465), .A(n3116), .ZN(U3279) );
  NAND2_X1 U3791 ( .A1(n3118), .A2(n4508), .ZN(n3120) );
  AND2_X1 U3792 ( .A1(n3120), .A2(n3119), .ZN(n3123) );
  INV_X1 U3793 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3121) );
  MUX2_X1 U3794 ( .A(n3123), .B(n3121), .S(n4522), .Z(n3122) );
  OAI21_X1 U3795 ( .B1(n3126), .B2(n4310), .A(n3122), .ZN(U3487) );
  MUX2_X1 U3796 ( .A(n3124), .B(n3123), .S(n4537), .Z(n3125) );
  OAI21_X1 U3797 ( .B1(n3126), .B2(n4264), .A(n3125), .ZN(U3528) );
  INV_X1 U3798 ( .A(n3238), .ZN(n3825) );
  AOI21_X1 U3799 ( .B1(n3245), .B2(n3241), .A(n3825), .ZN(n3205) );
  NAND2_X1 U3800 ( .A1(n3127), .A2(IR_REG_31__SCAN_IN), .ZN(n3128) );
  XNOR2_X1 U3801 ( .A(n3128), .B(IR_REG_12__SCAN_IN), .ZN(n3189) );
  MUX2_X1 U3802 ( .A(n3189), .B(DATAI_12_), .S(n3734), .Z(n3200) );
  OR2_X1 U3803 ( .A1(n3877), .A2(n3201), .ZN(n3240) );
  NAND2_X1 U3804 ( .A1(n3877), .A2(n3201), .ZN(n3237) );
  NAND2_X1 U3805 ( .A1(n3240), .A2(n3237), .ZN(n3148) );
  INV_X1 U3806 ( .A(n3148), .ZN(n3761) );
  XNOR2_X1 U3807 ( .A(n3205), .B(n3761), .ZN(n3138) );
  NAND2_X1 U3808 ( .A1(n3878), .A2(n4188), .ZN(n3136) );
  NAND2_X1 U3809 ( .A1(n3400), .A2(REG1_REG_13__SCAN_IN), .ZN(n3134) );
  NAND2_X1 U3810 ( .A1(n3129), .A2(n3184), .ZN(n3130) );
  AND2_X1 U3811 ( .A1(n3208), .A2(n3130), .ZN(n3279) );
  NAND2_X1 U3812 ( .A1(n3412), .A2(n3279), .ZN(n3133) );
  NAND2_X1 U3813 ( .A1(n3445), .A2(REG0_REG_13__SCAN_IN), .ZN(n3132) );
  NAND2_X1 U3814 ( .A1(n3725), .A2(REG2_REG_13__SCAN_IN), .ZN(n3131) );
  NAND4_X1 U3815 ( .A1(n3134), .A2(n3133), .A3(n3132), .A4(n3131), .ZN(n3876)
         );
  NAND2_X1 U3816 ( .A1(n3876), .A2(n4169), .ZN(n3135) );
  OAI211_X1 U3817 ( .C1(n4207), .C2(n3201), .A(n3136), .B(n3135), .ZN(n3137)
         );
  AOI21_X1 U3818 ( .B1(n3138), .B2(n4175), .A(n3137), .ZN(n3309) );
  OR2_X1 U3819 ( .A1(n3139), .A2(n3201), .ZN(n3140) );
  NAND2_X1 U3820 ( .A1(n3221), .A2(n3140), .ZN(n3315) );
  INV_X1 U3821 ( .A(n3315), .ZN(n3144) );
  INV_X1 U3822 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3142) );
  INV_X1 U3823 ( .A(n3141), .ZN(n3164) );
  OAI22_X1 U3824 ( .A1(n4350), .A2(n3142), .B1(n3164), .B2(n4197), .ZN(n3143)
         );
  AOI21_X1 U3825 ( .B1(n3144), .B2(n4461), .A(n3143), .ZN(n3150) );
  INV_X1 U3826 ( .A(n3878), .ZN(n3159) );
  NAND2_X1 U3827 ( .A1(n3159), .A2(n3145), .ZN(n3146) );
  XNOR2_X1 U3828 ( .A(n3203), .B(n3148), .ZN(n3307) );
  NAND2_X1 U3829 ( .A1(n3307), .A2(n4107), .ZN(n3149) );
  OAI211_X1 U3830 ( .C1(n3309), .C2(n4465), .A(n3150), .B(n3149), .ZN(U3278)
         );
  NAND2_X1 U3831 ( .A1(n3152), .A2(n3151), .ZN(n3154) );
  NAND2_X1 U3832 ( .A1(n3154), .A2(n3153), .ZN(n3296) );
  OAI22_X1 U3833 ( .A1(n3215), .A2(n2572), .B1(n3201), .B2(n3577), .ZN(n3155)
         );
  XNOR2_X1 U3834 ( .A(n3155), .B(n3571), .ZN(n3291) );
  NOR2_X1 U3835 ( .A1(n2572), .A2(n3201), .ZN(n3156) );
  AOI21_X1 U3836 ( .B1(n3877), .B2(n3566), .A(n3156), .ZN(n3290) );
  XNOR2_X1 U3837 ( .A(n3291), .B(n3290), .ZN(n3157) );
  XNOR2_X1 U3838 ( .A(n3296), .B(n3157), .ZN(n3158) );
  NAND2_X1 U3839 ( .A1(n3158), .A2(n4337), .ZN(n3163) );
  OAI22_X1 U3840 ( .A1(n3684), .A2(n3201), .B1(n3229), .B2(n4335), .ZN(n3161)
         );
  NAND2_X1 U3841 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4391) );
  OAI21_X1 U3842 ( .B1(n3683), .B2(n3159), .A(n4391), .ZN(n3160) );
  NOR2_X1 U3843 ( .A1(n3161), .A2(n3160), .ZN(n3162) );
  OAI211_X1 U3844 ( .C1(n4342), .C2(n3164), .A(n3163), .B(n3162), .ZN(U3221)
         );
  INV_X1 U3845 ( .A(IR_REG_10__SCAN_IN), .ZN(n3166) );
  INV_X1 U3846 ( .A(IR_REG_12__SCAN_IN), .ZN(n3165) );
  NAND3_X1 U3847 ( .A1(n3166), .A2(n4737), .A3(n3165), .ZN(n3167) );
  NOR2_X1 U3848 ( .A1(n3171), .A2(n3170), .ZN(n3169) );
  MUX2_X1 U3849 ( .A(n3170), .B(n3169), .S(IR_REG_13__SCAN_IN), .Z(n3173) );
  NAND2_X1 U3850 ( .A1(n3171), .A2(n4738), .ZN(n3318) );
  INV_X1 U3851 ( .A(n3318), .ZN(n3172) );
  NAND2_X1 U3852 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3188), .ZN(n3178) );
  INV_X1 U3853 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3174) );
  AOI22_X1 U3854 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3188), .B1(n4475), .B2(
        n3174), .ZN(n4386) );
  NAND2_X1 U3855 ( .A1(n3175), .A2(n4319), .ZN(n3177) );
  NAND2_X1 U3856 ( .A1(n3189), .A2(n3179), .ZN(n3180) );
  INV_X1 U3857 ( .A(n3189), .ZN(n4474) );
  XNOR2_X1 U3858 ( .A(n3179), .B(n4474), .ZN(n4395) );
  NAND2_X1 U3859 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4395), .ZN(n4394) );
  NAND2_X1 U3860 ( .A1(n3180), .A2(n4394), .ZN(n3932) );
  INV_X1 U3861 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3181) );
  NOR2_X1 U3862 ( .A1(n3199), .A2(n3181), .ZN(n3931) );
  AOI21_X1 U3863 ( .B1(n3181), .B2(n3199), .A(n3931), .ZN(n3183) );
  AOI21_X1 U3864 ( .B1(n3183), .B2(n3932), .A(n4398), .ZN(n3182) );
  OAI21_X1 U3865 ( .B1(n3932), .B2(n3183), .A(n3182), .ZN(n3198) );
  NOR2_X1 U3866 ( .A1(STATE_REG_SCAN_IN), .A2(n3184), .ZN(n3275) );
  INV_X1 U3867 ( .A(n3185), .ZN(n3187) );
  INV_X1 U3868 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4535) );
  AOI22_X1 U3869 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4475), .B1(n3188), .B2(
        n4535), .ZN(n4380) );
  NOR2_X1 U3870 ( .A1(n3190), .A2(n4474), .ZN(n3191) );
  INV_X1 U3871 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4633) );
  NOR2_X1 U3872 ( .A1(n3191), .A2(n4389), .ZN(n3195) );
  NAND2_X1 U3873 ( .A1(n4318), .A2(REG1_REG_13__SCAN_IN), .ZN(n3918) );
  INV_X1 U3874 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3365) );
  NAND2_X1 U3875 ( .A1(n3199), .A2(n3365), .ZN(n3192) );
  NAND2_X1 U3876 ( .A1(n3918), .A2(n3192), .ZN(n3194) );
  INV_X1 U3877 ( .A(n3919), .ZN(n3193) );
  AOI211_X1 U3878 ( .C1(n3195), .C2(n3194), .A(n3193), .B(n4433), .ZN(n3196)
         );
  AOI211_X1 U3879 ( .C1(n4437), .C2(ADDR_REG_13__SCAN_IN), .A(n3275), .B(n3196), .ZN(n3197) );
  OAI211_X1 U3880 ( .C1(n4449), .C2(n3199), .A(n3198), .B(n3197), .ZN(U3253)
         );
  NAND2_X1 U3881 ( .A1(n3877), .A2(n3200), .ZN(n3202) );
  MUX2_X1 U3882 ( .A(n4318), .B(DATAI_13_), .S(n3734), .Z(n3243) );
  XNOR2_X1 U3883 ( .A(n3876), .B(n3230), .ZN(n3764) );
  XNOR2_X1 U3884 ( .A(n3232), .B(n3764), .ZN(n3220) );
  INV_X1 U3885 ( .A(n3240), .ZN(n3204) );
  OAI21_X1 U3886 ( .B1(n3205), .B2(n3204), .A(n3237), .ZN(n3206) );
  XNOR2_X1 U3887 ( .A(n3206), .B(n3764), .ZN(n3217) );
  NAND2_X1 U3888 ( .A1(n3400), .A2(REG1_REG_14__SCAN_IN), .ZN(n3213) );
  INV_X1 U3889 ( .A(REG3_REG_14__SCAN_IN), .ZN(n3207) );
  AND2_X1 U3890 ( .A1(n3208), .A2(n3207), .ZN(n3209) );
  OR2_X1 U3891 ( .A1(n3247), .A2(n3209), .ZN(n3306) );
  INV_X1 U3892 ( .A(n3306), .ZN(n3259) );
  NAND2_X1 U3893 ( .A1(n3412), .A2(n3259), .ZN(n3212) );
  NAND2_X1 U3894 ( .A1(n3445), .A2(REG0_REG_14__SCAN_IN), .ZN(n3211) );
  NAND2_X1 U3895 ( .A1(n3725), .A2(REG2_REG_14__SCAN_IN), .ZN(n3210) );
  NAND4_X1 U3896 ( .A1(n3213), .A2(n3212), .A3(n3211), .A4(n3210), .ZN(n3875)
         );
  AOI22_X1 U3897 ( .A1(n3875), .A2(n4169), .B1(n4217), .B2(n3243), .ZN(n3214)
         );
  OAI21_X1 U3898 ( .B1(n3215), .B2(n4172), .A(n3214), .ZN(n3216) );
  AOI21_X1 U3899 ( .B1(n3217), .B2(n4175), .A(n3216), .ZN(n3218) );
  OAI21_X1 U3900 ( .B1(n3220), .B2(n3219), .A(n3218), .ZN(n3363) );
  INV_X1 U3901 ( .A(n3363), .ZN(n3226) );
  INV_X1 U3902 ( .A(n3220), .ZN(n3364) );
  NAND2_X1 U3903 ( .A1(n3221), .A2(n3243), .ZN(n3222) );
  NAND2_X1 U3904 ( .A1(n3257), .A2(n3222), .ZN(n3369) );
  AOI22_X1 U3905 ( .A1(n4465), .A2(REG2_REG_13__SCAN_IN), .B1(n3279), .B2(
        n4457), .ZN(n3223) );
  OAI21_X1 U3906 ( .B1(n3369), .B2(n4195), .A(n3223), .ZN(n3224) );
  AOI21_X1 U3907 ( .B1(n3364), .B2(n4459), .A(n3224), .ZN(n3225) );
  OAI21_X1 U3908 ( .B1(n3226), .B2(n4465), .A(n3225), .ZN(U3277) );
  NAND2_X1 U3909 ( .A1(n3318), .A2(IR_REG_31__SCAN_IN), .ZN(n3227) );
  INV_X1 U3910 ( .A(IR_REG_14__SCAN_IN), .ZN(n4750) );
  XNOR2_X1 U3911 ( .A(n3227), .B(n4750), .ZN(n3934) );
  INV_X1 U3912 ( .A(DATAI_14_), .ZN(n3228) );
  MUX2_X1 U3913 ( .A(n3934), .B(n3228), .S(n3734), .Z(n3317) );
  OR2_X1 U3914 ( .A1(n3875), .A2(n3317), .ZN(n3714) );
  NAND2_X1 U3915 ( .A1(n3875), .A2(n3317), .ZN(n3715) );
  NAND2_X1 U3916 ( .A1(n3714), .A2(n3715), .ZN(n3246) );
  NAND2_X1 U3917 ( .A1(n3232), .A2(n3231), .ZN(n3234) );
  NAND2_X1 U3918 ( .A1(n3876), .A2(n3243), .ZN(n3233) );
  NAND2_X1 U3919 ( .A1(n3234), .A2(n3233), .ZN(n3235) );
  AOI21_X1 U3920 ( .B1(n3779), .B2(n3235), .A(n3316), .ZN(n3282) );
  NAND2_X1 U3921 ( .A1(n3876), .A2(n3230), .ZN(n3236) );
  NAND2_X1 U3922 ( .A1(n3237), .A2(n3236), .ZN(n3823) );
  INV_X1 U3923 ( .A(n3823), .ZN(n3239) );
  NAND2_X1 U3924 ( .A1(n3239), .A2(n3238), .ZN(n3244) );
  AOI21_X1 U3925 ( .B1(n3241), .B2(n3240), .A(n3823), .ZN(n3242) );
  AOI21_X1 U3926 ( .B1(n3229), .B2(n3243), .A(n3242), .ZN(n3831) );
  OAI21_X2 U3927 ( .B1(n3245), .B2(n3244), .A(n3831), .ZN(n3718) );
  XNOR2_X1 U3928 ( .A(n3718), .B(n3246), .ZN(n3255) );
  NAND2_X1 U3929 ( .A1(n3400), .A2(REG1_REG_15__SCAN_IN), .ZN(n3252) );
  OR2_X1 U3930 ( .A1(n3247), .A2(REG3_REG_15__SCAN_IN), .ZN(n3248) );
  AND2_X1 U3931 ( .A1(n3355), .A2(n3248), .ZN(n3709) );
  NAND2_X1 U3932 ( .A1(n3412), .A2(n3709), .ZN(n3251) );
  NAND2_X1 U3933 ( .A1(n3445), .A2(REG0_REG_15__SCAN_IN), .ZN(n3250) );
  NAND2_X1 U3934 ( .A1(n3725), .A2(REG2_REG_15__SCAN_IN), .ZN(n3249) );
  NAND4_X1 U3935 ( .A1(n3252), .A2(n3251), .A3(n3250), .A4(n3249), .ZN(n3874)
         );
  INV_X1 U3936 ( .A(n3874), .ZN(n3640) );
  OAI22_X1 U3937 ( .A1(n3640), .A2(n4185), .B1(n3317), .B2(n4207), .ZN(n3253)
         );
  AOI21_X1 U3938 ( .B1(n4188), .B2(n3876), .A(n3253), .ZN(n3254) );
  OAI21_X1 U3939 ( .B1(n3255), .B2(n4190), .A(n3254), .ZN(n3283) );
  INV_X1 U3940 ( .A(n3317), .ZN(n3256) );
  INV_X1 U3941 ( .A(n4861), .ZN(n3258) );
  OAI21_X1 U3942 ( .B1(n2193), .B2(n3317), .A(n3258), .ZN(n3288) );
  AOI22_X1 U3943 ( .A1(n4465), .A2(REG2_REG_14__SCAN_IN), .B1(n3259), .B2(
        n4457), .ZN(n3260) );
  OAI21_X1 U3944 ( .B1(n3288), .B2(n4195), .A(n3260), .ZN(n3261) );
  AOI21_X1 U3945 ( .B1(n3283), .B2(n4350), .A(n3261), .ZN(n3262) );
  OAI21_X1 U3946 ( .B1(n3282), .B2(n4203), .A(n3262), .ZN(U3276) );
  NAND2_X1 U3947 ( .A1(n3876), .A2(n3561), .ZN(n3264) );
  OR2_X1 U3948 ( .A1(n3577), .A2(n3230), .ZN(n3263) );
  NAND2_X1 U3949 ( .A1(n3264), .A2(n3263), .ZN(n3265) );
  XNOR2_X1 U3950 ( .A(n3265), .B(n3578), .ZN(n3269) );
  INV_X1 U3951 ( .A(n3269), .ZN(n3267) );
  OAI22_X1 U3952 ( .A1(n3229), .A2(n3531), .B1(n3230), .B2(n3576), .ZN(n3268)
         );
  INV_X1 U3953 ( .A(n3268), .ZN(n3266) );
  NAND2_X1 U3954 ( .A1(n3267), .A2(n3266), .ZN(n3292) );
  NAND2_X1 U3955 ( .A1(n3269), .A2(n3268), .ZN(n3289) );
  NAND2_X1 U3956 ( .A1(n3292), .A2(n3289), .ZN(n3274) );
  INV_X1 U3957 ( .A(n3291), .ZN(n3270) );
  NOR2_X1 U3958 ( .A1(n3296), .A2(n3270), .ZN(n3272) );
  INV_X1 U3959 ( .A(n3296), .ZN(n3271) );
  OAI22_X1 U3960 ( .A1(n3272), .A2(n3290), .B1(n3271), .B2(n3291), .ZN(n3273)
         );
  XOR2_X1 U3961 ( .A(n3274), .B(n3273), .Z(n3281) );
  AOI21_X1 U3962 ( .B1(n4327), .B2(n3877), .A(n3275), .ZN(n3277) );
  NAND2_X1 U3963 ( .A1(n3704), .A2(n3875), .ZN(n3276) );
  OAI211_X1 U3964 ( .C1(n3684), .C2(n3230), .A(n3277), .B(n3276), .ZN(n3278)
         );
  AOI21_X1 U3965 ( .B1(n3710), .B2(n3279), .A(n3278), .ZN(n3280) );
  OAI21_X1 U3966 ( .B1(n3281), .B2(n3712), .A(n3280), .ZN(U3231) );
  INV_X1 U3967 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4402) );
  INV_X1 U3968 ( .A(n3282), .ZN(n3284) );
  AOI21_X1 U3969 ( .B1(n3284), .B2(n4508), .A(n3283), .ZN(n3286) );
  MUX2_X1 U3970 ( .A(n4402), .B(n3286), .S(n4537), .Z(n3285) );
  OAI21_X1 U3971 ( .B1(n4264), .B2(n3288), .A(n3285), .ZN(U3532) );
  INV_X1 U3972 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4723) );
  MUX2_X1 U3973 ( .A(n4723), .B(n3286), .S(n4524), .Z(n3287) );
  OAI21_X1 U3974 ( .B1(n3288), .B2(n4310), .A(n3287), .ZN(U3495) );
  OAI21_X1 U3975 ( .B1(n3291), .B2(n3290), .A(n3289), .ZN(n3295) );
  NAND3_X1 U3976 ( .A1(n3291), .A2(n3290), .A3(n3289), .ZN(n3293) );
  AND2_X1 U3977 ( .A1(n3293), .A2(n3292), .ZN(n3294) );
  NAND2_X1 U3978 ( .A1(n3875), .A2(n3561), .ZN(n3298) );
  OR2_X1 U3979 ( .A1(n3577), .A2(n3317), .ZN(n3297) );
  NAND2_X1 U3980 ( .A1(n3298), .A2(n3297), .ZN(n3299) );
  XNOR2_X1 U3981 ( .A(n3299), .B(n3571), .ZN(n3499) );
  INV_X1 U3982 ( .A(n3875), .ZN(n3329) );
  OAI22_X1 U3983 ( .A1(n3329), .A2(n3531), .B1(n3317), .B2(n3576), .ZN(n3496)
         );
  XNOR2_X1 U3984 ( .A(n3499), .B(n3496), .ZN(n3300) );
  XNOR2_X1 U3985 ( .A(n3498), .B(n3300), .ZN(n3301) );
  NAND2_X1 U3986 ( .A1(n3301), .A2(n4337), .ZN(n3305) );
  OAI22_X1 U3987 ( .A1(n3684), .A2(n3317), .B1(n3229), .B2(n3683), .ZN(n3303)
         );
  NAND2_X1 U3988 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4408) );
  OAI21_X1 U3989 ( .B1(n4335), .B2(n3640), .A(n4408), .ZN(n3302) );
  NOR2_X1 U3990 ( .A1(n3303), .A2(n3302), .ZN(n3304) );
  OAI211_X1 U3991 ( .C1(n4342), .C2(n3306), .A(n3305), .B(n3304), .ZN(U3212)
         );
  NAND2_X1 U3992 ( .A1(n3307), .A2(n4508), .ZN(n3308) );
  NAND2_X1 U3993 ( .A1(n3309), .A2(n3308), .ZN(n3312) );
  MUX2_X1 U3994 ( .A(REG1_REG_12__SCAN_IN), .B(n3312), .S(n4537), .Z(n3310) );
  INV_X1 U3995 ( .A(n3310), .ZN(n3311) );
  OAI21_X1 U3996 ( .B1(n4264), .B2(n3315), .A(n3311), .ZN(U3530) );
  MUX2_X1 U3997 ( .A(REG0_REG_12__SCAN_IN), .B(n3312), .S(n4524), .Z(n3313) );
  INV_X1 U3998 ( .A(n3313), .ZN(n3314) );
  OAI21_X1 U3999 ( .B1(n3315), .B2(n4310), .A(n3314), .ZN(U3491) );
  NAND2_X1 U4000 ( .A1(n3319), .A2(IR_REG_31__SCAN_IN), .ZN(n3338) );
  XNOR2_X1 U4001 ( .A(n3338), .B(IR_REG_15__SCAN_IN), .ZN(n3936) );
  MUX2_X1 U4002 ( .A(n3936), .B(DATAI_15_), .S(n4862), .Z(n3335) );
  OR2_X1 U4003 ( .A1(n3874), .A2(n3707), .ZN(n3717) );
  NAND2_X1 U4004 ( .A1(n3874), .A2(n3707), .ZN(n3716) );
  NAND2_X1 U4005 ( .A1(n3717), .A2(n3716), .ZN(n3321) );
  XNOR2_X1 U4006 ( .A(n3334), .B(n3321), .ZN(n4272) );
  INV_X1 U4007 ( .A(n3714), .ZN(n3320) );
  AOI21_X1 U4008 ( .B1(n3718), .B2(n3779), .A(n3320), .ZN(n3322) );
  INV_X1 U4009 ( .A(n3321), .ZN(n3777) );
  NAND2_X1 U4010 ( .A1(n3322), .A2(n3777), .ZN(n3350) );
  OAI211_X1 U4011 ( .C1(n3322), .C2(n3777), .A(n3350), .B(n4175), .ZN(n3328)
         );
  NAND2_X1 U4012 ( .A1(n2608), .A2(REG1_REG_16__SCAN_IN), .ZN(n3326) );
  XNOR2_X1 U4013 ( .A(n3355), .B(REG3_REG_16__SCAN_IN), .ZN(n3347) );
  NAND2_X1 U4014 ( .A1(n3412), .A2(n3347), .ZN(n3325) );
  NAND2_X1 U4015 ( .A1(n3445), .A2(REG0_REG_16__SCAN_IN), .ZN(n3324) );
  NAND2_X1 U4016 ( .A1(n3725), .A2(REG2_REG_16__SCAN_IN), .ZN(n3323) );
  NAND4_X1 U4017 ( .A1(n3326), .A2(n3325), .A3(n3324), .A4(n3323), .ZN(n4187)
         );
  AOI22_X1 U4018 ( .A1(n4187), .A2(n4169), .B1(n4217), .B2(n3335), .ZN(n3327)
         );
  OAI211_X1 U4019 ( .C1(n3329), .C2(n4172), .A(n3328), .B(n3327), .ZN(n4269)
         );
  XNOR2_X1 U4020 ( .A(n4861), .B(n3335), .ZN(n4270) );
  INV_X1 U4021 ( .A(n4270), .ZN(n3331) );
  AOI22_X1 U4022 ( .A1(n4465), .A2(REG2_REG_15__SCAN_IN), .B1(n3709), .B2(
        n4457), .ZN(n3330) );
  OAI21_X1 U4023 ( .B1(n3331), .B2(n4195), .A(n3330), .ZN(n3332) );
  AOI21_X1 U4024 ( .B1(n4269), .B2(n4350), .A(n3332), .ZN(n3333) );
  OAI21_X1 U4025 ( .B1(n4272), .B2(n4203), .A(n3333), .ZN(U3275) );
  INV_X1 U4026 ( .A(IR_REG_15__SCAN_IN), .ZN(n3337) );
  NAND2_X1 U4027 ( .A1(n3338), .A2(n3337), .ZN(n3339) );
  NAND2_X1 U4028 ( .A1(n3339), .A2(IR_REG_31__SCAN_IN), .ZN(n3341) );
  INV_X1 U4029 ( .A(IR_REG_16__SCAN_IN), .ZN(n3340) );
  INV_X1 U4030 ( .A(DATAI_16_), .ZN(n4471) );
  OR2_X1 U4031 ( .A1(n4187), .A2(n3641), .ZN(n3836) );
  NAND2_X1 U4032 ( .A1(n4187), .A2(n3641), .ZN(n3832) );
  NAND2_X1 U4033 ( .A1(n3836), .A2(n3832), .ZN(n3765) );
  NAND2_X1 U4034 ( .A1(n3342), .A2(n3765), .ZN(n3380) );
  OAI21_X1 U4035 ( .B1(n3342), .B2(n3765), .A(n3380), .ZN(n4268) );
  INV_X1 U4036 ( .A(n3641), .ZN(n3346) );
  INV_X1 U4037 ( .A(n3344), .ZN(n3345) );
  INV_X1 U4038 ( .A(n3486), .ZN(n4194) );
  AOI21_X1 U4039 ( .B1(n3346), .B2(n3345), .A(n4194), .ZN(n4266) );
  INV_X1 U4040 ( .A(REG2_REG_16__SCAN_IN), .ZN(n3348) );
  INV_X1 U4041 ( .A(n3347), .ZN(n3646) );
  OAI22_X1 U4042 ( .A1(n4350), .A2(n3348), .B1(n3646), .B2(n4197), .ZN(n3349)
         );
  AOI21_X1 U40430 ( .B1(n4266), .B2(n4461), .A(n3349), .ZN(n3362) );
  NAND2_X1 U4044 ( .A1(n3350), .A2(n3716), .ZN(n3352) );
  INV_X1 U4045 ( .A(n3765), .ZN(n3351) );
  NAND2_X1 U4046 ( .A1(n3352), .A2(n3351), .ZN(n3469) );
  OAI211_X1 U4047 ( .C1(n3352), .C2(n3351), .A(n3469), .B(n4175), .ZN(n3360)
         );
  INV_X1 U4048 ( .A(REG3_REG_16__SCAN_IN), .ZN(n3354) );
  INV_X1 U4049 ( .A(REG3_REG_17__SCAN_IN), .ZN(n3353) );
  OAI21_X1 U4050 ( .B1(n3355), .B2(n3354), .A(n3353), .ZN(n3356) );
  AND2_X1 U4051 ( .A1(n3356), .A2(n3373), .ZN(n4196) );
  AOI22_X1 U4052 ( .A1(n3412), .A2(n4196), .B1(n3445), .B2(
        REG0_REG_17__SCAN_IN), .ZN(n3358) );
  AOI22_X1 U4053 ( .A1(n3400), .A2(REG1_REG_17__SCAN_IN), .B1(n3725), .B2(
        REG2_REG_17__SCAN_IN), .ZN(n3357) );
  AOI22_X1 U4054 ( .A1(n4326), .A2(n4169), .B1(n4188), .B2(n3874), .ZN(n3359)
         );
  OAI211_X1 U4055 ( .C1(n4207), .C2(n3641), .A(n3360), .B(n3359), .ZN(n4265)
         );
  NAND2_X1 U4056 ( .A1(n4265), .A2(n4350), .ZN(n3361) );
  OAI211_X1 U4057 ( .C1(n4268), .C2(n4203), .A(n3362), .B(n3361), .ZN(U3274)
         );
  AOI21_X1 U4058 ( .B1(n4521), .B2(n3364), .A(n3363), .ZN(n3367) );
  MUX2_X1 U4059 ( .A(n3365), .B(n3367), .S(n4537), .Z(n3366) );
  OAI21_X1 U4060 ( .B1(n4264), .B2(n3369), .A(n3366), .ZN(U3531) );
  INV_X1 U4061 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4724) );
  MUX2_X1 U4062 ( .A(n4724), .B(n3367), .S(n4524), .Z(n3368) );
  OAI21_X1 U4063 ( .B1(n3369), .B2(n4310), .A(n3368), .ZN(U3493) );
  INV_X1 U4064 ( .A(REG1_REG_28__SCAN_IN), .ZN(n3484) );
  INV_X1 U4065 ( .A(n3370), .ZN(n3383) );
  NAND2_X1 U4066 ( .A1(n3383), .A2(IR_REG_31__SCAN_IN), .ZN(n3371) );
  XNOR2_X1 U4067 ( .A(n3371), .B(IR_REG_18__SCAN_IN), .ZN(n4469) );
  INV_X1 U4068 ( .A(n4469), .ZN(n4448) );
  INV_X1 U4069 ( .A(DATAI_18_), .ZN(n3372) );
  MUX2_X1 U4070 ( .A(n4448), .B(n3372), .S(n4862), .Z(n4164) );
  INV_X1 U4071 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4333) );
  AND2_X1 U4072 ( .A1(n3373), .A2(n4333), .ZN(n3374) );
  OR2_X1 U4073 ( .A1(n3374), .A2(n3387), .ZN(n4341) );
  INV_X1 U4074 ( .A(n4341), .ZN(n3375) );
  NAND2_X1 U4075 ( .A1(n3412), .A2(n3375), .ZN(n3379) );
  NAND2_X1 U4076 ( .A1(n2608), .A2(REG1_REG_18__SCAN_IN), .ZN(n3378) );
  NAND2_X1 U4077 ( .A1(n3445), .A2(REG0_REG_18__SCAN_IN), .ZN(n3377) );
  NAND2_X1 U4078 ( .A1(n3725), .A2(REG2_REG_18__SCAN_IN), .ZN(n3376) );
  NAND4_X1 U4079 ( .A1(n3379), .A2(n3378), .A3(n3377), .A4(n3376), .ZN(n4150)
         );
  INV_X1 U4080 ( .A(n4187), .ZN(n3508) );
  NAND2_X1 U4081 ( .A1(n3381), .A2(IR_REG_31__SCAN_IN), .ZN(n3382) );
  MUX2_X1 U4082 ( .A(IR_REG_31__SCAN_IN), .B(n3382), .S(IR_REG_17__SCAN_IN), 
        .Z(n3384) );
  NAND2_X1 U4083 ( .A1(n3384), .A2(n3383), .ZN(n3930) );
  INV_X1 U4084 ( .A(DATAI_17_), .ZN(n4550) );
  MUX2_X1 U4085 ( .A(n3930), .B(n4550), .S(n4862), .Z(n4193) );
  NAND2_X1 U4086 ( .A1(n4173), .A2(n4193), .ZN(n3386) );
  INV_X1 U4087 ( .A(n4193), .ZN(n3485) );
  OR2_X1 U4088 ( .A1(n4150), .A2(n4164), .ZN(n3472) );
  NAND2_X1 U4089 ( .A1(n4150), .A2(n4164), .ZN(n4143) );
  NAND2_X1 U4090 ( .A1(n3472), .A2(n4143), .ZN(n4168) );
  NOR2_X1 U4091 ( .A1(n3387), .A2(REG3_REG_19__SCAN_IN), .ZN(n3388) );
  OR2_X1 U4092 ( .A1(n3393), .A2(n3388), .ZN(n3615) );
  INV_X1 U4093 ( .A(n3615), .ZN(n4156) );
  NAND2_X1 U4094 ( .A1(n4156), .A2(n3412), .ZN(n3392) );
  NAND2_X1 U4095 ( .A1(n3400), .A2(REG1_REG_19__SCAN_IN), .ZN(n3391) );
  NAND2_X1 U4096 ( .A1(n3445), .A2(REG0_REG_19__SCAN_IN), .ZN(n3390) );
  NAND2_X1 U4097 ( .A1(n3725), .A2(REG2_REG_19__SCAN_IN), .ZN(n3389) );
  NAND4_X1 U4098 ( .A1(n3392), .A2(n3391), .A3(n3390), .A4(n3389), .ZN(n4170)
         );
  MUX2_X1 U4099 ( .A(n4316), .B(DATAI_19_), .S(n4862), .Z(n4152) );
  NOR2_X1 U4100 ( .A1(n4170), .A2(n4152), .ZN(n3750) );
  NAND2_X1 U4101 ( .A1(n4170), .A2(n4152), .ZN(n3748) );
  AOI22_X1 U4102 ( .A1(n2608), .A2(REG1_REG_20__SCAN_IN), .B1(n3445), .B2(
        REG0_REG_20__SCAN_IN), .ZN(n3397) );
  OR2_X1 U4103 ( .A1(n3393), .A2(REG3_REG_20__SCAN_IN), .ZN(n3394) );
  AND2_X1 U4104 ( .A1(n3398), .A2(n3394), .ZN(n3667) );
  NAND2_X1 U4105 ( .A1(n3667), .A2(n3412), .ZN(n3396) );
  NAND2_X1 U4106 ( .A1(n3725), .A2(REG2_REG_20__SCAN_IN), .ZN(n3395) );
  INV_X1 U4107 ( .A(n4129), .ZN(n4122) );
  NAND2_X1 U4108 ( .A1(n4139), .A2(n4129), .ZN(n3747) );
  INV_X1 U4109 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4111) );
  INV_X1 U4110 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3621) );
  NAND2_X1 U4111 ( .A1(n3398), .A2(n3621), .ZN(n3399) );
  NAND2_X1 U4112 ( .A1(n3404), .A2(n3399), .ZN(n4110) );
  OR2_X1 U4113 ( .A1(n4110), .A2(n3462), .ZN(n3402) );
  AOI22_X1 U4114 ( .A1(n3400), .A2(REG1_REG_21__SCAN_IN), .B1(n3445), .B2(
        REG0_REG_21__SCAN_IN), .ZN(n3401) );
  NAND2_X1 U4115 ( .A1(n4862), .A2(DATAI_21_), .ZN(n4109) );
  INV_X1 U4116 ( .A(n4109), .ZN(n4099) );
  NAND2_X1 U4117 ( .A1(n4123), .A2(n4099), .ZN(n3403) );
  INV_X1 U4118 ( .A(n4123), .ZN(n4086) );
  AOI22_X1 U4119 ( .A1(n4105), .A2(n3403), .B1(n4086), .B2(n4109), .ZN(n4082)
         );
  INV_X1 U4120 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4585) );
  NAND2_X1 U4121 ( .A1(n3404), .A2(n4585), .ZN(n3405) );
  NAND2_X1 U4122 ( .A1(n3410), .A2(n3405), .ZN(n4092) );
  AOI22_X1 U4123 ( .A1(n2608), .A2(REG1_REG_22__SCAN_IN), .B1(n3445), .B2(
        REG0_REG_22__SCAN_IN), .ZN(n3407) );
  NAND2_X1 U4124 ( .A1(n3725), .A2(REG2_REG_22__SCAN_IN), .ZN(n3406) );
  OAI211_X1 U4125 ( .C1(n4092), .C2(n3462), .A(n3407), .B(n3406), .ZN(n4067)
         );
  OR2_X1 U4126 ( .A1(n4067), .A2(n4091), .ZN(n4063) );
  NAND2_X1 U4127 ( .A1(n4067), .A2(n4091), .ZN(n3478) );
  NAND2_X1 U4128 ( .A1(n4063), .A2(n3478), .ZN(n4083) );
  NAND2_X1 U4129 ( .A1(n4082), .A2(n4083), .ZN(n4081) );
  INV_X1 U4130 ( .A(n4067), .ZN(n4102) );
  NAND2_X1 U4131 ( .A1(n4081), .A2(n3409), .ZN(n4058) );
  INV_X1 U4132 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4835) );
  AND2_X1 U4133 ( .A1(n3410), .A2(n4835), .ZN(n3411) );
  NOR2_X1 U4134 ( .A1(n3419), .A2(n3411), .ZN(n3598) );
  NAND2_X1 U4135 ( .A1(n3598), .A2(n3412), .ZN(n3417) );
  INV_X1 U4136 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4788) );
  NAND2_X1 U4137 ( .A1(n3725), .A2(REG2_REG_23__SCAN_IN), .ZN(n3414) );
  NAND2_X1 U4138 ( .A1(n3445), .A2(REG0_REG_23__SCAN_IN), .ZN(n3413) );
  OAI211_X1 U4139 ( .C1(n3729), .C2(n4788), .A(n3414), .B(n3413), .ZN(n3415)
         );
  INV_X1 U4140 ( .A(n3415), .ZN(n3416) );
  NAND2_X1 U4141 ( .A1(n4085), .A2(n4073), .ZN(n3418) );
  AOI22_X2 U4142 ( .A1(n4058), .A2(n3418), .B1(n4044), .B2(n4066), .ZN(n4038)
         );
  OR2_X1 U4143 ( .A1(n3419), .A2(REG3_REG_24__SCAN_IN), .ZN(n3420) );
  NAND2_X1 U4144 ( .A1(n3419), .A2(REG3_REG_24__SCAN_IN), .ZN(n3427) );
  AND2_X1 U4145 ( .A1(n3420), .A2(n3427), .ZN(n4053) );
  NAND2_X1 U4146 ( .A1(n4053), .A2(n3412), .ZN(n3425) );
  INV_X1 U4147 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4790) );
  NAND2_X1 U4148 ( .A1(n3725), .A2(REG2_REG_24__SCAN_IN), .ZN(n3422) );
  NAND2_X1 U4149 ( .A1(n3445), .A2(REG0_REG_24__SCAN_IN), .ZN(n3421) );
  OAI211_X1 U4150 ( .C1(n3729), .C2(n4790), .A(n3422), .B(n3421), .ZN(n3423)
         );
  INV_X1 U4151 ( .A(n3423), .ZN(n3424) );
  NAND2_X1 U4152 ( .A1(n4862), .A2(DATAI_24_), .ZN(n3551) );
  NAND2_X1 U4153 ( .A1(n4068), .A2(n4050), .ZN(n3426) );
  INV_X1 U4154 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4576) );
  NAND2_X1 U4155 ( .A1(n3427), .A2(n4576), .ZN(n3428) );
  NAND2_X1 U4156 ( .A1(n4033), .A2(n3412), .ZN(n3433) );
  INV_X1 U4157 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4235) );
  NAND2_X1 U4158 ( .A1(n3725), .A2(REG2_REG_25__SCAN_IN), .ZN(n3430) );
  NAND2_X1 U4159 ( .A1(n3445), .A2(REG0_REG_25__SCAN_IN), .ZN(n3429) );
  OAI211_X1 U4160 ( .C1(n3729), .C2(n4235), .A(n3430), .B(n3429), .ZN(n3431)
         );
  INV_X1 U4161 ( .A(n3431), .ZN(n3432) );
  INV_X1 U4162 ( .A(n4045), .ZN(n3434) );
  NAND2_X1 U4163 ( .A1(n4862), .A2(DATAI_25_), .ZN(n4032) );
  NAND2_X1 U4164 ( .A1(n3434), .A2(n4032), .ZN(n3435) );
  INV_X1 U4165 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3695) );
  AND2_X1 U4166 ( .A1(n3436), .A2(n3695), .ZN(n3437) );
  OR2_X1 U4167 ( .A1(n3437), .A2(n3443), .ZN(n3692) );
  INV_X1 U4168 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4231) );
  NAND2_X1 U4169 ( .A1(n3725), .A2(REG2_REG_26__SCAN_IN), .ZN(n3439) );
  NAND2_X1 U4170 ( .A1(n3445), .A2(REG0_REG_26__SCAN_IN), .ZN(n3438) );
  OAI211_X1 U4171 ( .C1(n3729), .C2(n4231), .A(n3439), .B(n3438), .ZN(n3440)
         );
  INV_X1 U4172 ( .A(n3440), .ZN(n3441) );
  NAND2_X1 U4173 ( .A1(n4862), .A2(DATAI_26_), .ZN(n4015) );
  INV_X1 U4174 ( .A(n4015), .ZN(n4010) );
  NAND2_X1 U4175 ( .A1(n4026), .A2(n4010), .ZN(n3442) );
  NOR2_X1 U4176 ( .A1(n3443), .A2(REG3_REG_27__SCAN_IN), .ZN(n3444) );
  INV_X1 U4177 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4800) );
  NAND2_X1 U4178 ( .A1(n3725), .A2(REG2_REG_27__SCAN_IN), .ZN(n3447) );
  NAND2_X1 U4179 ( .A1(n3445), .A2(REG0_REG_27__SCAN_IN), .ZN(n3446) );
  OAI211_X1 U4180 ( .C1(n3729), .C2(n4800), .A(n3447), .B(n3446), .ZN(n3448)
         );
  INV_X1 U4181 ( .A(n3448), .ZN(n3449) );
  INV_X1 U4182 ( .A(n3873), .ZN(n4013) );
  NAND2_X1 U4183 ( .A1(n3454), .A2(REG3_REG_28__SCAN_IN), .ZN(n3953) );
  OR2_X1 U4184 ( .A1(n3454), .A2(REG3_REG_28__SCAN_IN), .ZN(n3455) );
  NAND2_X1 U4185 ( .A1(n3980), .A2(n3412), .ZN(n3460) );
  NAND2_X1 U4186 ( .A1(n3725), .A2(REG2_REG_28__SCAN_IN), .ZN(n3457) );
  NAND2_X1 U4187 ( .A1(n3445), .A2(REG0_REG_28__SCAN_IN), .ZN(n3456) );
  OAI211_X1 U4188 ( .C1(n3729), .C2(n3484), .A(n3457), .B(n3456), .ZN(n3458)
         );
  INV_X1 U4189 ( .A(n3458), .ZN(n3459) );
  NAND2_X1 U4190 ( .A1(n4862), .A2(DATAI_28_), .ZN(n3585) );
  NOR2_X1 U4191 ( .A1(n3967), .A2(n3585), .ZN(n3954) );
  NAND2_X1 U4192 ( .A1(n3967), .A2(n3585), .ZN(n3955) );
  INV_X1 U4193 ( .A(n3955), .ZN(n3461) );
  INV_X1 U4194 ( .A(n3964), .ZN(n3786) );
  XNOR2_X1 U4195 ( .A(n3965), .B(n3786), .ZN(n3979) );
  OR2_X1 U4196 ( .A1(n3953), .A2(n3462), .ZN(n3468) );
  INV_X1 U4197 ( .A(REG1_REG_29__SCAN_IN), .ZN(n3465) );
  NAND2_X1 U4198 ( .A1(n3725), .A2(REG2_REG_29__SCAN_IN), .ZN(n3464) );
  NAND2_X1 U4199 ( .A1(n3445), .A2(REG0_REG_29__SCAN_IN), .ZN(n3463) );
  OAI211_X1 U4200 ( .C1(n3465), .C2(n3729), .A(n3464), .B(n3463), .ZN(n3466)
         );
  INV_X1 U4201 ( .A(n3466), .ZN(n3467) );
  OAI22_X1 U4202 ( .A1(n3737), .A2(n4185), .B1(n4207), .B2(n3585), .ZN(n3482)
         );
  NAND2_X1 U4203 ( .A1(n4100), .A2(n4129), .ZN(n3475) );
  NAND2_X1 U4204 ( .A1(n4326), .A2(n4193), .ZN(n3767) );
  AND2_X1 U4205 ( .A1(n3475), .A2(n3767), .ZN(n3471) );
  INV_X1 U4206 ( .A(n4152), .ZN(n4138) );
  NAND2_X1 U4207 ( .A1(n4170), .A2(n4138), .ZN(n3470) );
  AND2_X1 U4208 ( .A1(n4143), .A2(n3470), .ZN(n3473) );
  NAND2_X1 U4209 ( .A1(n3471), .A2(n3473), .ZN(n3835) );
  INV_X1 U4210 ( .A(n3472), .ZN(n4144) );
  NOR2_X1 U4211 ( .A1(n4326), .A2(n4193), .ZN(n4140) );
  NOR2_X1 U4212 ( .A1(n4144), .A2(n4140), .ZN(n3474) );
  INV_X1 U4213 ( .A(n3473), .ZN(n4117) );
  OAI22_X1 U4214 ( .A1(n3474), .A2(n4117), .B1(n4170), .B2(n4138), .ZN(n4118)
         );
  NOR2_X1 U4215 ( .A1(n4100), .A2(n4129), .ZN(n3476) );
  OAI21_X1 U4216 ( .B1(n4118), .B2(n3476), .A(n3475), .ZN(n4060) );
  INV_X1 U4217 ( .A(n4063), .ZN(n3477) );
  NOR2_X1 U4218 ( .A1(n4123), .A2(n4109), .ZN(n4062) );
  NOR2_X1 U4219 ( .A1(n3477), .A2(n4062), .ZN(n3844) );
  NAND2_X1 U4220 ( .A1(n4060), .A2(n3844), .ZN(n3722) );
  AND2_X1 U4221 ( .A1(n4123), .A2(n4109), .ZN(n3838) );
  OAI21_X1 U4222 ( .B1(n4085), .B2(n4066), .A(n3478), .ZN(n3842) );
  AOI21_X1 U4223 ( .B1(n3838), .B2(n4063), .A(n3842), .ZN(n3721) );
  OAI21_X1 U4224 ( .B1(n4059), .B2(n3722), .A(n3721), .ZN(n4041) );
  NOR2_X1 U4225 ( .A1(n4044), .A2(n4073), .ZN(n4039) );
  NOR2_X1 U4226 ( .A1(n4068), .A2(n3551), .ZN(n3751) );
  NOR2_X1 U4227 ( .A1(n4039), .A2(n3751), .ZN(n3845) );
  NAND2_X1 U4228 ( .A1(n4041), .A2(n3845), .ZN(n4023) );
  NAND2_X1 U4229 ( .A1(n4045), .A2(n4032), .ZN(n3756) );
  NAND2_X1 U4230 ( .A1(n4068), .A2(n3551), .ZN(n4022) );
  NAND2_X1 U4231 ( .A1(n4023), .A2(n3846), .ZN(n4006) );
  OR2_X1 U4232 ( .A1(n4026), .A2(n4015), .ZN(n3753) );
  OR2_X1 U4233 ( .A1(n4045), .A2(n4032), .ZN(n4005) );
  AND2_X1 U4234 ( .A1(n4026), .A2(n4015), .ZN(n3754) );
  AOI21_X1 U4235 ( .B1(n4006), .B2(n3853), .A(n3754), .ZN(n3989) );
  XNOR2_X1 U4236 ( .A(n3873), .B(n3996), .ZN(n3994) );
  NAND2_X1 U4237 ( .A1(n3989), .A2(n3994), .ZN(n3988) );
  NOR2_X1 U4238 ( .A1(n3873), .A2(n3450), .ZN(n3733) );
  INV_X1 U4239 ( .A(n3733), .ZN(n3479) );
  NAND2_X1 U4240 ( .A1(n3988), .A2(n3479), .ZN(n3956) );
  XNOR2_X1 U4241 ( .A(n3956), .B(n3964), .ZN(n3480) );
  NOR2_X1 U4242 ( .A1(n3480), .A2(n4190), .ZN(n3481) );
  AOI211_X1 U4243 ( .C1(n4188), .C2(n3873), .A(n3482), .B(n3481), .ZN(n3987)
         );
  INV_X1 U4244 ( .A(n3987), .ZN(n3483) );
  AOI21_X1 U4245 ( .B1(n3979), .B2(n4508), .A(n3483), .ZN(n3489) );
  INV_X1 U4246 ( .A(n3585), .ZN(n3966) );
  AOI21_X1 U4248 ( .B1(n3966), .B2(n2157), .A(n3974), .ZN(n3984) );
  NAND2_X1 U4249 ( .A1(n3984), .A2(n4215), .ZN(n3487) );
  NAND2_X1 U4250 ( .A1(n3488), .A2(n3487), .ZN(U3546) );
  INV_X1 U4251 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4804) );
  NAND2_X1 U4252 ( .A1(n3984), .A2(n4276), .ZN(n3490) );
  NAND2_X1 U4253 ( .A1(n3491), .A2(n3490), .ZN(U3514) );
  NAND2_X1 U4254 ( .A1(n4123), .A2(n3561), .ZN(n3493) );
  OR2_X1 U4255 ( .A1(n3577), .A2(n4109), .ZN(n3492) );
  NAND2_X1 U4256 ( .A1(n3493), .A2(n3492), .ZN(n3494) );
  XNOR2_X1 U4257 ( .A(n3494), .B(n3571), .ZN(n3617) );
  INV_X1 U4258 ( .A(n3617), .ZN(n3538) );
  NOR2_X1 U4259 ( .A1(n2572), .A2(n4109), .ZN(n3495) );
  AOI21_X1 U4260 ( .B1(n3566), .B2(n4123), .A(n3495), .ZN(n3536) );
  INV_X1 U4261 ( .A(n3536), .ZN(n3616) );
  NAND2_X1 U4262 ( .A1(n3498), .A2(n3499), .ZN(n3497) );
  NAND2_X1 U4263 ( .A1(n3497), .A2(n3496), .ZN(n3503) );
  INV_X1 U4264 ( .A(n3498), .ZN(n3501) );
  INV_X1 U4265 ( .A(n3499), .ZN(n3500) );
  NAND2_X1 U4266 ( .A1(n3501), .A2(n3500), .ZN(n3502) );
  NAND2_X1 U4267 ( .A1(n3874), .A2(n3561), .ZN(n3505) );
  OR2_X1 U4268 ( .A1(n3577), .A2(n3707), .ZN(n3504) );
  NAND2_X1 U4269 ( .A1(n3505), .A2(n3504), .ZN(n3506) );
  XNOR2_X1 U4270 ( .A(n3506), .B(n3578), .ZN(n3510) );
  NOR2_X1 U4271 ( .A1(n2572), .A2(n3707), .ZN(n3507) );
  AOI21_X1 U4272 ( .B1(n3566), .B2(n3874), .A(n3507), .ZN(n3701) );
  OAI22_X1 U4273 ( .A1(n3508), .A2(n3531), .B1(n3576), .B2(n3641), .ZN(n3512)
         );
  OAI22_X1 U4274 ( .A1(n3508), .A2(n2572), .B1(n3577), .B2(n3641), .ZN(n3509)
         );
  XNOR2_X1 U4275 ( .A(n3509), .B(n3578), .ZN(n3513) );
  XOR2_X1 U4276 ( .A(n3512), .B(n3513), .Z(n3638) );
  NOR2_X1 U4277 ( .A1(n3576), .A2(n4193), .ZN(n3514) );
  AOI21_X1 U4278 ( .B1(n4326), .B2(n3566), .A(n3514), .ZN(n3647) );
  OAI22_X1 U4279 ( .A1(n4173), .A2(n2572), .B1(n4193), .B2(n3577), .ZN(n3515)
         );
  XNOR2_X1 U4280 ( .A(n3515), .B(n3571), .ZN(n3648) );
  INV_X1 U4281 ( .A(n3647), .ZN(n3518) );
  INV_X1 U4282 ( .A(n3648), .ZN(n3517) );
  NAND2_X1 U4283 ( .A1(n4150), .A2(n3561), .ZN(n3520) );
  OR2_X1 U4284 ( .A1(n3577), .A2(n4164), .ZN(n3519) );
  NAND2_X1 U4285 ( .A1(n3520), .A2(n3519), .ZN(n3521) );
  XNOR2_X1 U4286 ( .A(n3521), .B(n3578), .ZN(n3523) );
  OAI22_X1 U4287 ( .A1(n2304), .A2(n3531), .B1(n3576), .B2(n4164), .ZN(n3522)
         );
  NAND2_X1 U4288 ( .A1(n3523), .A2(n3522), .ZN(n4330) );
  NOR2_X1 U4289 ( .A1(n3523), .A2(n3522), .ZN(n4331) );
  AOI22_X1 U4290 ( .A1(n3566), .A2(n4170), .B1(n3561), .B2(n4152), .ZN(n3527)
         );
  NAND2_X1 U4291 ( .A1(n4170), .A2(n3561), .ZN(n3525) );
  OR2_X1 U4292 ( .A1(n3577), .A2(n4138), .ZN(n3524) );
  NAND2_X1 U4293 ( .A1(n3525), .A2(n3524), .ZN(n3526) );
  XNOR2_X1 U4294 ( .A(n3526), .B(n3578), .ZN(n3529) );
  XOR2_X1 U4295 ( .A(n3527), .B(n3529), .Z(n3609) );
  INV_X1 U4296 ( .A(n3527), .ZN(n3528) );
  OAI22_X1 U4297 ( .A1(n4139), .A2(n2572), .B1(n3577), .B2(n4129), .ZN(n3530)
         );
  XNOR2_X1 U4298 ( .A(n3530), .B(n3578), .ZN(n3532) );
  OAI22_X1 U4299 ( .A1(n4139), .A2(n3531), .B1(n3576), .B2(n4129), .ZN(n3533)
         );
  NAND2_X1 U4300 ( .A1(n3532), .A2(n3533), .ZN(n3671) );
  INV_X1 U4301 ( .A(n3532), .ZN(n3535) );
  INV_X1 U4302 ( .A(n3533), .ZN(n3534) );
  NAND2_X1 U4303 ( .A1(n3535), .A2(n3534), .ZN(n3672) );
  AOI21_X1 U4304 ( .B1(n3617), .B2(n3536), .A(n3619), .ZN(n3537) );
  AOI21_X1 U4305 ( .B1(n3538), .B2(n3616), .A(n3537), .ZN(n3680) );
  OAI22_X1 U4306 ( .A1(n4102), .A2(n3531), .B1(n4091), .B2(n3576), .ZN(n3544)
         );
  NAND2_X1 U4307 ( .A1(n4067), .A2(n3561), .ZN(n3540) );
  OR2_X1 U4308 ( .A1(n3577), .A2(n4091), .ZN(n3539) );
  NAND2_X1 U4309 ( .A1(n3540), .A2(n3539), .ZN(n3541) );
  XNOR2_X1 U4310 ( .A(n3541), .B(n3578), .ZN(n3543) );
  XOR2_X1 U4311 ( .A(n3544), .B(n3543), .Z(n3681) );
  NAND2_X1 U4312 ( .A1(n3680), .A2(n3681), .ZN(n3679) );
  OAI22_X1 U4313 ( .A1(n4085), .A2(n3531), .B1(n4073), .B2(n3576), .ZN(n3549)
         );
  OAI22_X1 U4314 ( .A1(n4085), .A2(n2572), .B1(n4073), .B2(n3577), .ZN(n3542)
         );
  XNOR2_X1 U4315 ( .A(n3542), .B(n3578), .ZN(n3550) );
  XOR2_X1 U4316 ( .A(n3549), .B(n3550), .Z(n3601) );
  INV_X1 U4317 ( .A(n3543), .ZN(n3546) );
  INV_X1 U4318 ( .A(n3544), .ZN(n3545) );
  NAND2_X1 U4319 ( .A1(n3546), .A2(n3545), .ZN(n3599) );
  NOR2_X1 U4320 ( .A1(n3576), .A2(n3551), .ZN(n3548) );
  AOI21_X1 U4321 ( .B1(n4068), .B2(n3566), .A(n3548), .ZN(n3553) );
  NAND2_X1 U4322 ( .A1(n3550), .A2(n3549), .ZN(n3554) );
  OAI22_X1 U4323 ( .A1(n3603), .A2(n2572), .B1(n3551), .B2(n3577), .ZN(n3552)
         );
  XNOR2_X1 U4324 ( .A(n3552), .B(n3578), .ZN(n3657) );
  NAND2_X1 U4325 ( .A1(n4045), .A2(n3561), .ZN(n3556) );
  OR2_X1 U4326 ( .A1(n3577), .A2(n4032), .ZN(n3555) );
  NAND2_X1 U4327 ( .A1(n3556), .A2(n3555), .ZN(n3557) );
  XNOR2_X1 U4328 ( .A(n3557), .B(n3571), .ZN(n3560) );
  NOR2_X1 U4329 ( .A1(n3576), .A2(n4032), .ZN(n3558) );
  AOI21_X1 U4330 ( .B1(n4045), .B2(n3566), .A(n3558), .ZN(n3559) );
  AND2_X1 U4331 ( .A1(n3560), .A2(n3559), .ZN(n3626) );
  OR2_X1 U4332 ( .A1(n3560), .A2(n3559), .ZN(n3627) );
  NAND2_X1 U4333 ( .A1(n4026), .A2(n3561), .ZN(n3563) );
  OR2_X1 U4334 ( .A1(n3577), .A2(n4015), .ZN(n3562) );
  NAND2_X1 U4335 ( .A1(n3563), .A2(n3562), .ZN(n3564) );
  XNOR2_X1 U4336 ( .A(n3564), .B(n3571), .ZN(n3568) );
  NOR2_X1 U4337 ( .A1(n3576), .A2(n4015), .ZN(n3565) );
  AOI21_X1 U4338 ( .B1(n4026), .B2(n3566), .A(n3565), .ZN(n3567) );
  NOR2_X1 U4339 ( .A1(n3568), .A2(n3567), .ZN(n3689) );
  NAND2_X1 U4340 ( .A1(n3873), .A2(n3561), .ZN(n3570) );
  OR2_X1 U4341 ( .A1(n3577), .A2(n3450), .ZN(n3569) );
  NAND2_X1 U4342 ( .A1(n3570), .A2(n3569), .ZN(n3572) );
  XNOR2_X1 U4343 ( .A(n3572), .B(n3571), .ZN(n3574) );
  NOR2_X1 U4344 ( .A1(n3576), .A2(n3450), .ZN(n3573) );
  AOI21_X1 U4345 ( .B1(n3873), .B2(n3566), .A(n3573), .ZN(n3575) );
  XNOR2_X1 U4346 ( .A(n3574), .B(n3575), .ZN(n3590) );
  OAI22_X1 U4347 ( .A1(n3591), .A2(n3590), .B1(n3575), .B2(n3574), .ZN(n3583)
         );
  INV_X1 U4348 ( .A(n3967), .ZN(n3991) );
  OAI22_X1 U4349 ( .A1(n3991), .A2(n3531), .B1(n3585), .B2(n2572), .ZN(n3581)
         );
  OAI22_X1 U4350 ( .A1(n3991), .A2(n2572), .B1(n3585), .B2(n3577), .ZN(n3579)
         );
  XNOR2_X1 U4351 ( .A(n3579), .B(n3578), .ZN(n3580) );
  XOR2_X1 U4352 ( .A(n3581), .B(n3580), .Z(n3582) );
  XNOR2_X1 U4353 ( .A(n3583), .B(n3582), .ZN(n3589) );
  INV_X1 U4354 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3584) );
  OAI22_X1 U4355 ( .A1(n3737), .A2(n4335), .B1(STATE_REG_SCAN_IN), .B2(n3584), 
        .ZN(n3587) );
  OAI22_X1 U4356 ( .A1(n4013), .A2(n3683), .B1(n3684), .B2(n3585), .ZN(n3586)
         );
  AOI211_X1 U4357 ( .C1(n3980), .C2(n3710), .A(n3587), .B(n3586), .ZN(n3588)
         );
  OAI21_X1 U4358 ( .B1(n3589), .B2(n3712), .A(n3588), .ZN(U3217) );
  XNOR2_X1 U4359 ( .A(n3591), .B(n3590), .ZN(n3597) );
  INV_X1 U4360 ( .A(n3999), .ZN(n3595) );
  INV_X1 U4361 ( .A(n4026), .ZN(n3592) );
  INV_X1 U4362 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4808) );
  OAI22_X1 U4363 ( .A1(n3592), .A2(n3683), .B1(STATE_REG_SCAN_IN), .B2(n4808), 
        .ZN(n3594) );
  OAI22_X1 U4364 ( .A1(n3991), .A2(n4335), .B1(n3684), .B2(n3450), .ZN(n3593)
         );
  AOI211_X1 U4365 ( .C1(n3595), .C2(n3710), .A(n3594), .B(n3593), .ZN(n3596)
         );
  OAI21_X1 U4366 ( .B1(n3597), .B2(n3712), .A(n3596), .ZN(U3211) );
  INV_X1 U4367 ( .A(n3598), .ZN(n4075) );
  AND2_X1 U4368 ( .A1(n3679), .A2(n3599), .ZN(n3602) );
  OAI211_X1 U4369 ( .C1(n3602), .C2(n3601), .A(n4337), .B(n3600), .ZN(n3607)
         );
  OAI22_X1 U4370 ( .A1(n3684), .A2(n4073), .B1(n4102), .B2(n3683), .ZN(n3605)
         );
  OAI22_X1 U4371 ( .A1(n3603), .A2(n4335), .B1(STATE_REG_SCAN_IN), .B2(n4835), 
        .ZN(n3604) );
  NOR2_X1 U4372 ( .A1(n3605), .A2(n3604), .ZN(n3606) );
  OAI211_X1 U4373 ( .C1(n4342), .C2(n4075), .A(n3607), .B(n3606), .ZN(U3213)
         );
  XNOR2_X1 U4374 ( .A(n3608), .B(n3609), .ZN(n3610) );
  NAND2_X1 U4375 ( .A1(n3610), .A2(n4337), .ZN(n3614) );
  OAI22_X1 U4376 ( .A1(n3684), .A2(n4138), .B1(n4139), .B2(n4335), .ZN(n3612)
         );
  NAND2_X1 U4377 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3949) );
  OAI21_X1 U4378 ( .B1(n3683), .B2(n2304), .A(n3949), .ZN(n3611) );
  NOR2_X1 U4379 ( .A1(n3612), .A2(n3611), .ZN(n3613) );
  OAI211_X1 U4380 ( .C1(n4342), .C2(n3615), .A(n3614), .B(n3613), .ZN(U3216)
         );
  XNOR2_X1 U4381 ( .A(n3617), .B(n3616), .ZN(n3618) );
  XNOR2_X1 U4382 ( .A(n3619), .B(n3618), .ZN(n3620) );
  NAND2_X1 U4383 ( .A1(n3620), .A2(n4337), .ZN(n3625) );
  OAI22_X1 U4384 ( .A1(n3684), .A2(n4109), .B1(n4139), .B2(n3683), .ZN(n3623)
         );
  OAI22_X1 U4385 ( .A1(n4335), .A2(n4102), .B1(STATE_REG_SCAN_IN), .B2(n3621), 
        .ZN(n3622) );
  NOR2_X1 U4386 ( .A1(n3623), .A2(n3622), .ZN(n3624) );
  OAI211_X1 U4387 ( .C1(n4342), .C2(n4110), .A(n3625), .B(n3624), .ZN(U3220)
         );
  INV_X1 U4388 ( .A(n3626), .ZN(n3628) );
  NAND2_X1 U4389 ( .A1(n3628), .A2(n3627), .ZN(n3629) );
  XNOR2_X1 U4390 ( .A(n3630), .B(n3629), .ZN(n3636) );
  INV_X1 U4391 ( .A(n4033), .ZN(n3633) );
  INV_X1 U4392 ( .A(n3684), .ZN(n4329) );
  AOI22_X1 U4393 ( .A1(n4026), .A2(n3704), .B1(n4329), .B2(n2190), .ZN(n3632)
         );
  AOI22_X1 U4394 ( .A1(n4327), .A2(n4068), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n3631) );
  OAI211_X1 U4395 ( .C1(n4342), .C2(n3633), .A(n3632), .B(n3631), .ZN(n3634)
         );
  INV_X1 U4396 ( .A(n3634), .ZN(n3635) );
  OAI21_X1 U4397 ( .B1(n3636), .B2(n3712), .A(n3635), .ZN(U3222) );
  AOI21_X1 U4398 ( .B1(n3701), .B2(n3700), .A(n3699), .ZN(n3637) );
  XOR2_X1 U4399 ( .A(n3638), .B(n3637), .Z(n3639) );
  NAND2_X1 U4400 ( .A1(n3639), .A2(n4337), .ZN(n3645) );
  OAI22_X1 U4401 ( .A1(n3684), .A2(n3641), .B1(n3640), .B2(n3683), .ZN(n3643)
         );
  NAND2_X1 U4402 ( .A1(REG3_REG_16__SCAN_IN), .A2(U3149), .ZN(n4422) );
  OAI21_X1 U4403 ( .B1(n4335), .B2(n4173), .A(n4422), .ZN(n3642) );
  NOR2_X1 U4404 ( .A1(n3643), .A2(n3642), .ZN(n3644) );
  OAI211_X1 U4405 ( .C1(n4342), .C2(n3646), .A(n3645), .B(n3644), .ZN(U3223)
         );
  XNOR2_X1 U4406 ( .A(n3648), .B(n3647), .ZN(n3649) );
  XNOR2_X1 U4407 ( .A(n3650), .B(n3649), .ZN(n3655) );
  AND2_X1 U4408 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n3929) );
  AOI21_X1 U4409 ( .B1(n4327), .B2(n4187), .A(n3929), .ZN(n3652) );
  NAND2_X1 U4410 ( .A1(n3704), .A2(n4150), .ZN(n3651) );
  OAI211_X1 U4411 ( .C1(n3684), .C2(n4193), .A(n3652), .B(n3651), .ZN(n3653)
         );
  AOI21_X1 U4412 ( .B1(n3710), .B2(n4196), .A(n3653), .ZN(n3654) );
  OAI21_X1 U4413 ( .B1(n3655), .B2(n3712), .A(n3654), .ZN(U3225) );
  NOR2_X1 U4414 ( .A1(n3656), .A2(n2166), .ZN(n3658) );
  XNOR2_X1 U4415 ( .A(n3658), .B(n3657), .ZN(n3666) );
  INV_X1 U4416 ( .A(n4053), .ZN(n3663) );
  INV_X1 U4417 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3659) );
  OAI22_X1 U4418 ( .A1(n3683), .A2(n4085), .B1(STATE_REG_SCAN_IN), .B2(n3659), 
        .ZN(n3660) );
  INV_X1 U4419 ( .A(n3660), .ZN(n3662) );
  AOI22_X1 U4420 ( .A1(n4329), .A2(n4050), .B1(n3704), .B2(n4045), .ZN(n3661)
         );
  OAI211_X1 U4421 ( .C1(n4342), .C2(n3663), .A(n3662), .B(n3661), .ZN(n3664)
         );
  INV_X1 U4422 ( .A(n3664), .ZN(n3665) );
  OAI21_X1 U4423 ( .B1(n3666), .B2(n3712), .A(n3665), .ZN(U3226) );
  INV_X1 U4424 ( .A(n3667), .ZN(n4130) );
  INV_X1 U4425 ( .A(n3672), .ZN(n3668) );
  NOR2_X1 U4426 ( .A1(n3669), .A2(n3668), .ZN(n3674) );
  AOI21_X1 U4427 ( .B1(n3672), .B2(n3671), .A(n3670), .ZN(n3673) );
  OAI21_X1 U4428 ( .B1(n3674), .B2(n3673), .A(n4337), .ZN(n3678) );
  OAI22_X1 U4429 ( .A1(n3684), .A2(n4129), .B1(n4086), .B2(n4335), .ZN(n3676)
         );
  INV_X1 U4430 ( .A(n4170), .ZN(n4334) );
  INV_X1 U4431 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4586) );
  OAI22_X1 U4432 ( .A1(n3683), .A2(n4334), .B1(STATE_REG_SCAN_IN), .B2(n4586), 
        .ZN(n3675) );
  NOR2_X1 U4433 ( .A1(n3676), .A2(n3675), .ZN(n3677) );
  OAI211_X1 U4434 ( .C1(n4342), .C2(n4130), .A(n3678), .B(n3677), .ZN(U3230)
         );
  OAI21_X1 U4435 ( .B1(n3681), .B2(n3680), .A(n3679), .ZN(n3682) );
  NAND2_X1 U4436 ( .A1(n3682), .A2(n4337), .ZN(n3688) );
  OAI22_X1 U4437 ( .A1(n3684), .A2(n4091), .B1(n4086), .B2(n3683), .ZN(n3686)
         );
  OAI22_X1 U4438 ( .A1(n4335), .A2(n4085), .B1(STATE_REG_SCAN_IN), .B2(n4585), 
        .ZN(n3685) );
  NOR2_X1 U4439 ( .A1(n3686), .A2(n3685), .ZN(n3687) );
  OAI211_X1 U4440 ( .C1(n4342), .C2(n4092), .A(n3688), .B(n3687), .ZN(U3232)
         );
  NOR2_X1 U4441 ( .A1(n3689), .A2(n2173), .ZN(n3690) );
  XNOR2_X1 U4442 ( .A(n3691), .B(n3690), .ZN(n3698) );
  INV_X1 U4443 ( .A(n3692), .ZN(n4016) );
  NAND2_X1 U4444 ( .A1(n3873), .A2(n3704), .ZN(n3694) );
  AOI22_X1 U4445 ( .A1(n4329), .A2(n4010), .B1(n4327), .B2(n4045), .ZN(n3693)
         );
  OAI211_X1 U4446 ( .C1(STATE_REG_SCAN_IN), .C2(n3695), .A(n3694), .B(n3693), 
        .ZN(n3696) );
  AOI21_X1 U4447 ( .B1(n4016), .B2(n3710), .A(n3696), .ZN(n3697) );
  OAI21_X1 U4448 ( .B1(n3698), .B2(n3712), .A(n3697), .ZN(U3237) );
  NAND2_X1 U4449 ( .A1(n2277), .A2(n3700), .ZN(n3702) );
  XNOR2_X1 U4450 ( .A(n3702), .B(n3701), .ZN(n3713) );
  INV_X1 U4451 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3703) );
  NOR2_X1 U4452 ( .A1(STATE_REG_SCAN_IN), .A2(n3703), .ZN(n4415) );
  AOI21_X1 U4453 ( .B1(n3704), .B2(n4187), .A(n4415), .ZN(n3706) );
  NAND2_X1 U4454 ( .A1(n4327), .A2(n3875), .ZN(n3705) );
  OAI211_X1 U4455 ( .C1(n3684), .C2(n3707), .A(n3706), .B(n3705), .ZN(n3708)
         );
  AOI21_X1 U4456 ( .B1(n3710), .B2(n3709), .A(n3708), .ZN(n3711) );
  OAI21_X1 U4457 ( .B1(n3713), .B2(n3712), .A(n3711), .ZN(U3238) );
  NAND2_X1 U4458 ( .A1(n4862), .A2(DATAI_30_), .ZN(n4211) );
  INV_X1 U4459 ( .A(n4211), .ZN(n4216) );
  NAND2_X1 U4460 ( .A1(n4862), .A2(DATAI_31_), .ZN(n4208) );
  NAND2_X1 U4461 ( .A1(n3714), .A2(n3717), .ZN(n3827) );
  NAND2_X1 U4462 ( .A1(n3716), .A2(n3715), .ZN(n3813) );
  NAND2_X1 U4463 ( .A1(n3813), .A2(n3717), .ZN(n3828) );
  OAI21_X1 U4464 ( .B1(n3718), .B2(n3827), .A(n3828), .ZN(n3720) );
  INV_X1 U4465 ( .A(n3832), .ZN(n3719) );
  AOI211_X1 U4466 ( .C1(n3720), .C2(n3836), .A(n3719), .B(n3835), .ZN(n3723)
         );
  OAI21_X1 U4467 ( .B1(n3723), .B2(n3722), .A(n3721), .ZN(n3724) );
  NAND2_X1 U4468 ( .A1(n3724), .A2(n3845), .ZN(n3736) );
  INV_X1 U4469 ( .A(n3959), .ZN(n3732) );
  INV_X1 U4470 ( .A(REG1_REG_31__SCAN_IN), .ZN(n3728) );
  NAND2_X1 U4471 ( .A1(n3725), .A2(REG2_REG_31__SCAN_IN), .ZN(n3727) );
  NAND2_X1 U4472 ( .A1(n3445), .A2(REG0_REG_31__SCAN_IN), .ZN(n3726) );
  OAI211_X1 U4473 ( .C1(n3729), .C2(n3728), .A(n3727), .B(n3726), .ZN(n4206)
         );
  INV_X1 U4474 ( .A(n4206), .ZN(n3731) );
  INV_X1 U4475 ( .A(n4208), .ZN(n3730) );
  NOR2_X1 U4476 ( .A1(n3731), .A2(n3730), .ZN(n3856) );
  AOI21_X1 U4477 ( .B1(n3732), .B2(n4216), .A(n3856), .ZN(n3757) );
  NOR2_X1 U4478 ( .A1(n3954), .A2(n3733), .ZN(n3739) );
  AND2_X1 U4479 ( .A1(n4862), .A2(DATAI_29_), .ZN(n3975) );
  NAND2_X1 U4480 ( .A1(n3737), .A2(n3975), .ZN(n3744) );
  NAND4_X1 U4481 ( .A1(n3853), .A2(n3757), .A3(n3739), .A4(n3744), .ZN(n3735)
         );
  AOI21_X1 U4482 ( .B1(n3736), .B2(n3846), .A(n3735), .ZN(n3742) );
  INV_X1 U4483 ( .A(n3737), .ZN(n3872) );
  INV_X1 U4484 ( .A(n3975), .ZN(n3973) );
  NAND2_X1 U4485 ( .A1(n3872), .A2(n3973), .ZN(n3745) );
  NAND2_X1 U4486 ( .A1(n3745), .A2(n3955), .ZN(n3738) );
  NOR2_X1 U4487 ( .A1(n3754), .A2(n3738), .ZN(n3849) );
  OAI211_X1 U4488 ( .C1(n3739), .C2(n3738), .A(n3757), .B(n3744), .ZN(n3857)
         );
  AOI21_X1 U4489 ( .B1(n3994), .B2(n3849), .A(n3857), .ZN(n3741) );
  NAND2_X1 U4490 ( .A1(n3959), .A2(n4211), .ZN(n3746) );
  AOI21_X1 U4491 ( .B1(n3746), .B2(n4206), .A(n4208), .ZN(n3740) );
  NOR3_X1 U4492 ( .A1(n3742), .A2(n3741), .A3(n3740), .ZN(n3743) );
  AOI21_X1 U4493 ( .B1(n4216), .B2(n4208), .A(n3743), .ZN(n3864) );
  NAND2_X1 U4494 ( .A1(n3745), .A2(n3744), .ZN(n3970) );
  OAI21_X1 U4495 ( .B1(n4206), .B2(n4208), .A(n3746), .ZN(n3854) );
  AND2_X1 U4496 ( .A1(n2177), .A2(n3747), .ZN(n4121) );
  INV_X1 U4497 ( .A(n3748), .ZN(n3749) );
  OR2_X1 U4498 ( .A1(n3750), .A2(n3749), .ZN(n4145) );
  INV_X1 U4499 ( .A(n4145), .ZN(n4136) );
  XNOR2_X1 U4500 ( .A(n4085), .B(n4066), .ZN(n4064) );
  INV_X1 U4501 ( .A(n4022), .ZN(n3752) );
  OR2_X1 U4502 ( .A1(n3752), .A2(n3751), .ZN(n4042) );
  NOR4_X1 U4503 ( .A1(n4121), .A2(n4136), .A3(n4064), .A4(n4042), .ZN(n3759)
         );
  INV_X1 U4504 ( .A(n3753), .ZN(n3755) );
  NOR2_X1 U4505 ( .A1(n3755), .A2(n3754), .ZN(n4007) );
  AND2_X1 U4506 ( .A1(n4005), .A2(n3756), .ZN(n4024) );
  AND4_X1 U4507 ( .A1(n3994), .A2(n4007), .A3(n4024), .A4(n3757), .ZN(n3758)
         );
  NAND3_X1 U4508 ( .A1(n2519), .A2(n3759), .A3(n3758), .ZN(n3760) );
  NOR2_X1 U4509 ( .A1(n3854), .A2(n3760), .ZN(n3762) );
  NAND3_X1 U4510 ( .A1(n3763), .A2(n3762), .A3(n3761), .ZN(n3766) );
  NOR2_X1 U4511 ( .A1(n4062), .A2(n3838), .ZN(n4106) );
  INV_X1 U4512 ( .A(n4106), .ZN(n3770) );
  INV_X1 U4513 ( .A(n3767), .ZN(n4142) );
  OR2_X1 U4514 ( .A1(n4142), .A2(n4140), .ZN(n4184) );
  OR4_X1 U4515 ( .A1(n3770), .A2(n4184), .A3(n3769), .A4(n3768), .ZN(n3783) );
  OR4_X1 U4516 ( .A1(n4168), .A2(n3773), .A3(n3772), .A4(n3771), .ZN(n3782) );
  INV_X1 U4517 ( .A(n2616), .ZN(n3774) );
  NAND4_X1 U4518 ( .A1(n3776), .A2(n3775), .A3(n3774), .A4(n2158), .ZN(n3781)
         );
  NAND4_X1 U4519 ( .A1(n3779), .A2(n3778), .A3(n3777), .A4(n4480), .ZN(n3780)
         );
  NOR4_X1 U4520 ( .A1(n3783), .A2(n3782), .A3(n3781), .A4(n3780), .ZN(n3784)
         );
  NAND4_X1 U4521 ( .A1(n3786), .A2(n3971), .A3(n3785), .A4(n3784), .ZN(n3861)
         );
  INV_X1 U4522 ( .A(n3787), .ZN(n3790) );
  OAI211_X1 U4523 ( .C1(n3790), .C2(n2517), .A(n3789), .B(n3788), .ZN(n3793)
         );
  NAND3_X1 U4524 ( .A1(n3793), .A2(n3792), .A3(n3791), .ZN(n3796) );
  NAND3_X1 U4525 ( .A1(n3796), .A2(n3795), .A3(n3794), .ZN(n3799) );
  NAND3_X1 U4526 ( .A1(n3799), .A2(n3798), .A3(n3797), .ZN(n3807) );
  INV_X1 U4527 ( .A(n3800), .ZN(n3802) );
  NOR3_X1 U4528 ( .A1(n3817), .A2(n3802), .A3(n3801), .ZN(n3806) );
  INV_X1 U4529 ( .A(n3803), .ZN(n3805) );
  AOI211_X1 U4530 ( .C1(n3807), .C2(n3806), .A(n3805), .B(n3804), .ZN(n3812)
         );
  NAND2_X1 U4531 ( .A1(n3809), .A2(n3808), .ZN(n3816) );
  OAI211_X1 U4532 ( .C1(n3812), .C2(n3816), .A(n3811), .B(n3810), .ZN(n3822)
         );
  NOR2_X1 U4533 ( .A1(n3813), .A2(n3815), .ZN(n3821) );
  NOR4_X1 U4534 ( .A1(n3817), .A2(n3816), .A3(n3815), .A4(n3814), .ZN(n3819)
         );
  OR2_X1 U4535 ( .A1(n3819), .A2(n3818), .ZN(n3820) );
  AOI22_X1 U4536 ( .A1(n3822), .A2(n3821), .B1(n3828), .B2(n3820), .ZN(n3826)
         );
  NOR4_X1 U4537 ( .A1(n3826), .A2(n3825), .A3(n3824), .A4(n3823), .ZN(n3834)
         );
  INV_X1 U4538 ( .A(n3827), .ZN(n3830) );
  INV_X1 U4539 ( .A(n3828), .ZN(n3829) );
  AOI21_X1 U4540 ( .B1(n3831), .B2(n3830), .A(n3829), .ZN(n3833) );
  OAI21_X1 U4541 ( .B1(n3834), .B2(n3833), .A(n3832), .ZN(n3837) );
  AOI21_X1 U4542 ( .B1(n3837), .B2(n3836), .A(n3835), .ZN(n3841) );
  INV_X1 U4543 ( .A(n4060), .ZN(n3840) );
  INV_X1 U4544 ( .A(n3838), .ZN(n3839) );
  OAI21_X1 U4545 ( .B1(n3841), .B2(n3840), .A(n3839), .ZN(n3843) );
  AOI21_X1 U4546 ( .B1(n3844), .B2(n3843), .A(n3842), .ZN(n3848) );
  INV_X1 U4547 ( .A(n3845), .ZN(n3847) );
  OAI21_X1 U4548 ( .B1(n3848), .B2(n3847), .A(n3846), .ZN(n3852) );
  NOR2_X1 U4549 ( .A1(n4013), .A2(n3996), .ZN(n3851) );
  INV_X1 U4550 ( .A(n3849), .ZN(n3850) );
  AOI211_X1 U4551 ( .C1(n3853), .C2(n3852), .A(n3851), .B(n3850), .ZN(n3858)
         );
  INV_X1 U4552 ( .A(n3854), .ZN(n3855) );
  OAI22_X1 U4553 ( .A1(n3858), .A2(n3857), .B1(n3856), .B2(n3855), .ZN(n3860)
         );
  MUX2_X1 U4554 ( .A(n3861), .B(n3860), .S(n3859), .Z(n3862) );
  OAI21_X1 U4555 ( .B1(n3864), .B2(n3863), .A(n3862), .ZN(n3865) );
  XNOR2_X1 U4556 ( .A(n3865), .B(n4316), .ZN(n3871) );
  INV_X1 U4557 ( .A(n3866), .ZN(n3867) );
  NOR2_X1 U4558 ( .A1(n3867), .A2(n3909), .ZN(n3869) );
  OAI21_X1 U4559 ( .B1(n3870), .B2(n4315), .A(B_REG_SCAN_IN), .ZN(n3868) );
  OAI22_X1 U4560 ( .A1(n3871), .A2(n3870), .B1(n3869), .B2(n3868), .ZN(U3239)
         );
  MUX2_X1 U4561 ( .A(n4206), .B(DATAO_REG_31__SCAN_IN), .S(n3889), .Z(U3581)
         );
  MUX2_X1 U4562 ( .A(n3872), .B(DATAO_REG_29__SCAN_IN), .S(n3889), .Z(U3579)
         );
  MUX2_X1 U4563 ( .A(n3967), .B(DATAO_REG_28__SCAN_IN), .S(n3889), .Z(U3578)
         );
  MUX2_X1 U4564 ( .A(n3873), .B(DATAO_REG_27__SCAN_IN), .S(n3889), .Z(U3577)
         );
  MUX2_X1 U4565 ( .A(n4026), .B(DATAO_REG_26__SCAN_IN), .S(n3889), .Z(U3576)
         );
  MUX2_X1 U4566 ( .A(n4045), .B(DATAO_REG_25__SCAN_IN), .S(n3889), .Z(U3575)
         );
  MUX2_X1 U4567 ( .A(n4068), .B(DATAO_REG_24__SCAN_IN), .S(n3889), .Z(U3574)
         );
  MUX2_X1 U4568 ( .A(DATAO_REG_23__SCAN_IN), .B(n4044), .S(U4043), .Z(U3573)
         );
  MUX2_X1 U4569 ( .A(n4067), .B(DATAO_REG_22__SCAN_IN), .S(n3889), .Z(U3572)
         );
  MUX2_X1 U4570 ( .A(n4123), .B(DATAO_REG_21__SCAN_IN), .S(n3889), .Z(U3571)
         );
  MUX2_X1 U4571 ( .A(DATAO_REG_20__SCAN_IN), .B(n4100), .S(U4043), .Z(U3570)
         );
  MUX2_X1 U4572 ( .A(n4170), .B(DATAO_REG_19__SCAN_IN), .S(n3889), .Z(U3569)
         );
  MUX2_X1 U4573 ( .A(DATAO_REG_17__SCAN_IN), .B(n4326), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4574 ( .A(n4187), .B(DATAO_REG_16__SCAN_IN), .S(n3889), .Z(U3566)
         );
  MUX2_X1 U4575 ( .A(n3874), .B(DATAO_REG_15__SCAN_IN), .S(n3889), .Z(U3565)
         );
  MUX2_X1 U4576 ( .A(n3875), .B(DATAO_REG_14__SCAN_IN), .S(n3889), .Z(U3564)
         );
  MUX2_X1 U4577 ( .A(n3876), .B(DATAO_REG_13__SCAN_IN), .S(n3889), .Z(U3563)
         );
  MUX2_X1 U4578 ( .A(DATAO_REG_12__SCAN_IN), .B(n3877), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U4579 ( .A(n3878), .B(DATAO_REG_11__SCAN_IN), .S(n3889), .Z(U3561)
         );
  MUX2_X1 U4580 ( .A(n3879), .B(DATAO_REG_10__SCAN_IN), .S(n3889), .Z(U3560)
         );
  MUX2_X1 U4581 ( .A(n3880), .B(DATAO_REG_9__SCAN_IN), .S(n3889), .Z(U3559) );
  MUX2_X1 U4582 ( .A(DATAO_REG_8__SCAN_IN), .B(n3881), .S(U4043), .Z(U3558) );
  MUX2_X1 U4583 ( .A(n3882), .B(DATAO_REG_7__SCAN_IN), .S(n3889), .Z(U3557) );
  MUX2_X1 U4584 ( .A(n3883), .B(DATAO_REG_6__SCAN_IN), .S(n3889), .Z(U3556) );
  MUX2_X1 U4585 ( .A(DATAO_REG_5__SCAN_IN), .B(n3884), .S(U4043), .Z(U3555) );
  MUX2_X1 U4586 ( .A(n3885), .B(DATAO_REG_4__SCAN_IN), .S(n3889), .Z(U3554) );
  MUX2_X1 U4587 ( .A(n3886), .B(DATAO_REG_3__SCAN_IN), .S(n3889), .Z(U3553) );
  MUX2_X1 U4588 ( .A(n3887), .B(DATAO_REG_2__SCAN_IN), .S(n3889), .Z(U3552) );
  MUX2_X1 U4589 ( .A(n3888), .B(DATAO_REG_1__SCAN_IN), .S(n3889), .Z(U3551) );
  MUX2_X1 U4590 ( .A(n2598), .B(DATAO_REG_0__SCAN_IN), .S(n3889), .Z(U3550) );
  MUX2_X1 U4591 ( .A(n4527), .B(REG1_REG_1__SCAN_IN), .S(n3890), .Z(n3892) );
  OAI211_X1 U4592 ( .C1(n3893), .C2(n3892), .A(n4429), .B(n3891), .ZN(n3899)
         );
  NAND2_X1 U4593 ( .A1(n4407), .A2(n4325), .ZN(n3898) );
  XOR2_X1 U4594 ( .A(n3911), .B(n3894), .Z(n3895) );
  NAND2_X1 U4595 ( .A1(n4445), .A2(n3895), .ZN(n3897) );
  AOI22_X1 U4596 ( .A1(n4437), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3896) );
  NAND4_X1 U4597 ( .A1(n3899), .A2(n3898), .A3(n3897), .A4(n3896), .ZN(U3241)
         );
  AOI22_X1 U4598 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4437), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3917) );
  XNOR2_X1 U4599 ( .A(n3901), .B(n3900), .ZN(n3903) );
  OAI22_X1 U4600 ( .A1(n3903), .A2(n4433), .B1(n4449), .B2(n3902), .ZN(n3904)
         );
  INV_X1 U4601 ( .A(n3904), .ZN(n3916) );
  OAI211_X1 U4602 ( .C1(n3907), .C2(n3906), .A(n4445), .B(n3905), .ZN(n3915)
         );
  INV_X1 U4603 ( .A(n4353), .ZN(n3910) );
  NAND3_X1 U4604 ( .A1(n3908), .A2(n4314), .A3(n3910), .ZN(n3914) );
  INV_X1 U4605 ( .A(n3909), .ZN(n3912) );
  OAI21_X1 U4606 ( .B1(REG2_REG_0__SCAN_IN), .B2(n3910), .A(n4314), .ZN(n4351)
         );
  AOI22_X1 U4607 ( .A1(n3912), .A2(n3911), .B1(n4351), .B2(n4547), .ZN(n3913)
         );
  NAND3_X1 U4608 ( .A1(n3914), .A2(U4043), .A3(n3913), .ZN(n4367) );
  NAND4_X1 U4609 ( .A1(n3917), .A2(n3916), .A3(n3915), .A4(n4367), .ZN(U3242)
         );
  INV_X1 U4610 ( .A(n3930), .ZN(n4317) );
  XNOR2_X1 U4611 ( .A(n3930), .B(REG1_REG_17__SCAN_IN), .ZN(n3927) );
  INV_X1 U4612 ( .A(n3934), .ZN(n4406) );
  INV_X1 U4613 ( .A(n3936), .ZN(n4473) );
  INV_X1 U4614 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3922) );
  AOI22_X1 U4615 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4473), .B1(n3936), .B2(
        n3922), .ZN(n4412) );
  NAND2_X1 U4616 ( .A1(n3924), .A2(n4472), .ZN(n3925) );
  INV_X1 U4617 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4774) );
  NAND2_X1 U4618 ( .A1(n3926), .A2(n3927), .ZN(n3944) );
  OAI21_X1 U4619 ( .B1(n3927), .B2(n3926), .A(n3944), .ZN(n3928) );
  AOI22_X1 U4620 ( .A1(n4317), .A2(n4407), .B1(n4429), .B2(n3928), .ZN(n3943)
         );
  AOI21_X1 U4621 ( .B1(n4437), .B2(ADDR_REG_17__SCAN_IN), .A(n3929), .ZN(n3942) );
  XNOR2_X1 U4622 ( .A(n3930), .B(REG2_REG_17__SCAN_IN), .ZN(n3939) );
  INV_X1 U4623 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4641) );
  NOR2_X1 U4624 ( .A1(n3935), .A2(n4399), .ZN(n4417) );
  INV_X1 U4625 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4645) );
  AOI22_X1 U4626 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4473), .B1(n3936), .B2(
        n4645), .ZN(n4418) );
  NOR2_X1 U4627 ( .A1(n4417), .A2(n4418), .ZN(n4416) );
  NAND2_X1 U4628 ( .A1(n3937), .A2(n4424), .ZN(n3938) );
  NAND2_X1 U4629 ( .A1(n3938), .A2(n3939), .ZN(n3947) );
  OAI21_X1 U4630 ( .B1(n3939), .B2(n3938), .A(n3947), .ZN(n3940) );
  NAND2_X1 U4631 ( .A1(n4445), .A2(n3940), .ZN(n3941) );
  NAND3_X1 U4632 ( .A1(n3943), .A2(n3942), .A3(n3941), .ZN(U3257) );
  INV_X1 U4633 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4573) );
  AOI22_X1 U4634 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4448), .B1(n4469), .B2(
        n4573), .ZN(n4434) );
  OAI21_X1 U4635 ( .B1(n4317), .B2(REG1_REG_17__SCAN_IN), .A(n3944), .ZN(n4435) );
  XNOR2_X1 U4636 ( .A(n4316), .B(REG1_REG_19__SCAN_IN), .ZN(n3945) );
  NAND2_X1 U4637 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4469), .ZN(n3946) );
  OAI21_X1 U4638 ( .B1(REG2_REG_18__SCAN_IN), .B2(n4469), .A(n3946), .ZN(n4443) );
  OAI21_X1 U4639 ( .B1(n4317), .B2(REG2_REG_17__SCAN_IN), .A(n3947), .ZN(n4442) );
  NAND2_X1 U4640 ( .A1(n4437), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3948) );
  OAI211_X1 U4641 ( .C1(n4449), .C2(n3950), .A(n3949), .B(n3948), .ZN(n3951)
         );
  INV_X1 U4642 ( .A(n3953), .ZN(n3963) );
  AOI21_X1 U4643 ( .B1(n3956), .B2(n3955), .A(n3954), .ZN(n3957) );
  XOR2_X1 U4644 ( .A(n3970), .B(n3957), .Z(n3962) );
  AND2_X1 U4645 ( .A1(n4353), .A2(B_REG_SCAN_IN), .ZN(n3958) );
  NOR2_X1 U4646 ( .A1(n4185), .A2(n3958), .ZN(n4205) );
  AOI22_X1 U4647 ( .A1(n3959), .A2(n4205), .B1(n3975), .B2(n4217), .ZN(n3961)
         );
  NAND2_X1 U4648 ( .A1(n3967), .A2(n4188), .ZN(n3960) );
  OAI211_X1 U4649 ( .C1(n3962), .C2(n4190), .A(n3961), .B(n3960), .ZN(n4223)
         );
  AOI21_X1 U4650 ( .B1(n3963), .B2(n4457), .A(n4223), .ZN(n3978) );
  NAND2_X1 U4651 ( .A1(n3969), .A2(n3968), .ZN(n3972) );
  XNOR2_X1 U4652 ( .A(n3972), .B(n3971), .ZN(n4222) );
  NAND2_X1 U4653 ( .A1(n4222), .A2(n4107), .ZN(n3977) );
  AOI22_X1 U4654 ( .A1(n4224), .A2(n4461), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4465), .ZN(n3976) );
  OAI211_X1 U4655 ( .C1(n4465), .C2(n3978), .A(n3977), .B(n3976), .ZN(U3354)
         );
  NAND2_X1 U4656 ( .A1(n3979), .A2(n4107), .ZN(n3986) );
  INV_X1 U4657 ( .A(n3980), .ZN(n3982) );
  INV_X1 U4658 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3981) );
  OAI22_X1 U4659 ( .A1(n3982), .A2(n4197), .B1(n3981), .B2(n4350), .ZN(n3983)
         );
  AOI21_X1 U4660 ( .B1(n3984), .B2(n4461), .A(n3983), .ZN(n3985) );
  OAI211_X1 U4661 ( .C1(n3987), .C2(n4465), .A(n3986), .B(n3985), .ZN(U3262)
         );
  OAI21_X1 U4662 ( .B1(n3994), .B2(n3989), .A(n3988), .ZN(n3993) );
  AOI22_X1 U4663 ( .A1(n4026), .A2(n4188), .B1(n3996), .B2(n4217), .ZN(n3990)
         );
  OAI21_X1 U4664 ( .B1(n3991), .B2(n4185), .A(n3990), .ZN(n3992) );
  AOI21_X1 U4665 ( .B1(n3993), .B2(n4175), .A(n3992), .ZN(n4226) );
  XNOR2_X1 U4666 ( .A(n3995), .B(n3994), .ZN(n4225) );
  NAND2_X1 U4667 ( .A1(n4225), .A2(n4107), .ZN(n4003) );
  NAND2_X1 U4668 ( .A1(n4014), .A2(n3996), .ZN(n3997) );
  NAND2_X1 U4669 ( .A1(n2157), .A2(n3997), .ZN(n4228) );
  INV_X1 U4670 ( .A(n4228), .ZN(n4001) );
  INV_X1 U4671 ( .A(REG2_REG_27__SCAN_IN), .ZN(n3998) );
  OAI22_X1 U4672 ( .A1(n3999), .A2(n4197), .B1(n3998), .B2(n4350), .ZN(n4000)
         );
  AOI21_X1 U4673 ( .B1(n4001), .B2(n4461), .A(n4000), .ZN(n4002) );
  OAI211_X1 U4674 ( .C1(n4226), .C2(n4465), .A(n4003), .B(n4002), .ZN(U3263)
         );
  INV_X1 U4675 ( .A(n4230), .ZN(n4020) );
  NAND2_X1 U4676 ( .A1(n4006), .A2(n4005), .ZN(n4008) );
  XNOR2_X1 U4677 ( .A(n4008), .B(n4007), .ZN(n4009) );
  NAND2_X1 U4678 ( .A1(n4009), .A2(n4175), .ZN(n4012) );
  AOI22_X1 U4679 ( .A1(n4045), .A2(n4188), .B1(n4010), .B2(n4217), .ZN(n4011)
         );
  OAI211_X1 U4680 ( .C1(n4013), .C2(n4185), .A(n4012), .B(n4011), .ZN(n4229)
         );
  OAI21_X1 U4681 ( .B1(n4860), .B2(n4015), .A(n4014), .ZN(n4284) );
  AOI22_X1 U4682 ( .A1(n4016), .A2(n4457), .B1(n4465), .B2(
        REG2_REG_26__SCAN_IN), .ZN(n4017) );
  OAI21_X1 U4683 ( .B1(n4284), .B2(n4195), .A(n4017), .ZN(n4018) );
  AOI21_X1 U4684 ( .B1(n4229), .B2(n4350), .A(n4018), .ZN(n4019) );
  OAI21_X1 U4685 ( .B1(n4020), .B2(n4203), .A(n4019), .ZN(U3264) );
  XNOR2_X1 U4686 ( .A(n4021), .B(n4024), .ZN(n4234) );
  INV_X1 U4687 ( .A(n4234), .ZN(n4037) );
  NAND2_X1 U4688 ( .A1(n4023), .A2(n4022), .ZN(n4025) );
  XNOR2_X1 U4689 ( .A(n4025), .B(n4024), .ZN(n4029) );
  AOI22_X1 U4690 ( .A1(n4068), .A2(n4188), .B1(n2190), .B2(n4217), .ZN(n4028)
         );
  NAND2_X1 U4691 ( .A1(n4026), .A2(n4169), .ZN(n4027) );
  OAI211_X1 U4692 ( .C1(n4029), .C2(n4190), .A(n4028), .B(n4027), .ZN(n4233)
         );
  INV_X1 U4693 ( .A(n4860), .ZN(n4031) );
  OAI21_X1 U4694 ( .B1(n4049), .B2(n4032), .A(n4031), .ZN(n4288) );
  AOI22_X1 U4695 ( .A1(n4465), .A2(REG2_REG_25__SCAN_IN), .B1(n4033), .B2(
        n4457), .ZN(n4034) );
  OAI21_X1 U4696 ( .B1(n4288), .B2(n4195), .A(n4034), .ZN(n4035) );
  AOI21_X1 U4697 ( .B1(n4233), .B2(n4350), .A(n4035), .ZN(n4036) );
  OAI21_X1 U4698 ( .B1(n4037), .B2(n4203), .A(n4036), .ZN(U3265) );
  XNOR2_X1 U4699 ( .A(n4038), .B(n4042), .ZN(n4238) );
  INV_X1 U4700 ( .A(n4238), .ZN(n4057) );
  INV_X1 U4701 ( .A(n4039), .ZN(n4040) );
  NAND2_X1 U4702 ( .A1(n4041), .A2(n4040), .ZN(n4043) );
  XNOR2_X1 U4703 ( .A(n4043), .B(n4042), .ZN(n4048) );
  AOI22_X1 U4704 ( .A1(n4044), .A2(n4188), .B1(n4050), .B2(n4217), .ZN(n4047)
         );
  NAND2_X1 U4705 ( .A1(n4045), .A2(n4169), .ZN(n4046) );
  OAI211_X1 U4706 ( .C1(n4048), .C2(n4190), .A(n4047), .B(n4046), .ZN(n4237)
         );
  INV_X1 U4707 ( .A(n4049), .ZN(n4052) );
  NAND2_X1 U4708 ( .A1(n4072), .A2(n4050), .ZN(n4051) );
  NAND2_X1 U4709 ( .A1(n4052), .A2(n4051), .ZN(n4292) );
  AOI22_X1 U4710 ( .A1(n4465), .A2(REG2_REG_24__SCAN_IN), .B1(n4053), .B2(
        n4457), .ZN(n4054) );
  OAI21_X1 U4711 ( .B1(n4292), .B2(n4195), .A(n4054), .ZN(n4055) );
  AOI21_X1 U4712 ( .B1(n4237), .B2(n4350), .A(n4055), .ZN(n4056) );
  OAI21_X1 U4713 ( .B1(n4057), .B2(n4203), .A(n4056), .ZN(U3266) );
  XOR2_X1 U4714 ( .A(n4064), .B(n4058), .Z(n4241) );
  INV_X1 U4715 ( .A(n4241), .ZN(n4080) );
  INV_X1 U4716 ( .A(n4059), .ZN(n4061) );
  NAND2_X1 U4717 ( .A1(n4061), .A2(n4060), .ZN(n4098) );
  AOI21_X1 U4718 ( .B1(n4098), .B2(n4106), .A(n4062), .ZN(n4084) );
  OAI21_X1 U4719 ( .B1(n4084), .B2(n4083), .A(n4063), .ZN(n4065) );
  XNOR2_X1 U4720 ( .A(n4065), .B(n4064), .ZN(n4071) );
  AOI22_X1 U4721 ( .A1(n4067), .A2(n4188), .B1(n4217), .B2(n4066), .ZN(n4070)
         );
  NAND2_X1 U4722 ( .A1(n4068), .A2(n4169), .ZN(n4069) );
  OAI211_X1 U4723 ( .C1(n4071), .C2(n4190), .A(n4070), .B(n4069), .ZN(n4240)
         );
  INV_X1 U4724 ( .A(n4243), .ZN(n4074) );
  OAI21_X1 U4725 ( .B1(n4074), .B2(n4073), .A(n4072), .ZN(n4295) );
  NOR2_X1 U4726 ( .A1(n4295), .A2(n4195), .ZN(n4078) );
  INV_X1 U4727 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4076) );
  OAI22_X1 U4728 ( .A1(n4350), .A2(n4076), .B1(n4075), .B2(n4197), .ZN(n4077)
         );
  AOI211_X1 U4729 ( .C1(n4240), .C2(n4350), .A(n4078), .B(n4077), .ZN(n4079)
         );
  OAI21_X1 U4730 ( .B1(n4080), .B2(n4203), .A(n4079), .ZN(U3267) );
  OAI21_X1 U4731 ( .B1(n4082), .B2(n4083), .A(n4081), .ZN(n4247) );
  XNOR2_X1 U4732 ( .A(n4084), .B(n4083), .ZN(n4089) );
  NOR2_X1 U4733 ( .A1(n4085), .A2(n4185), .ZN(n4088) );
  OAI22_X1 U4734 ( .A1(n4086), .A2(n4172), .B1(n4091), .B2(n4207), .ZN(n4087)
         );
  AOI211_X1 U4735 ( .C1(n4089), .C2(n4175), .A(n4088), .B(n4087), .ZN(n4246)
         );
  INV_X1 U4736 ( .A(n4246), .ZN(n4096) );
  INV_X1 U4737 ( .A(n4090), .ZN(n4108) );
  NAND2_X1 U4738 ( .A1(n4108), .A2(n3408), .ZN(n4244) );
  AND3_X1 U4739 ( .A1(n4244), .A2(n4461), .A3(n4243), .ZN(n4095) );
  INV_X1 U4740 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4093) );
  OAI22_X1 U4741 ( .A1(n4350), .A2(n4093), .B1(n4092), .B2(n4197), .ZN(n4094)
         );
  AOI211_X1 U4742 ( .C1(n4096), .C2(n4350), .A(n4095), .B(n4094), .ZN(n4097)
         );
  OAI21_X1 U4743 ( .B1(n4247), .B2(n4203), .A(n4097), .ZN(U3268) );
  XNOR2_X1 U4744 ( .A(n4098), .B(n4106), .ZN(n4104) );
  AOI22_X1 U4745 ( .A1(n4100), .A2(n4188), .B1(n4217), .B2(n4099), .ZN(n4101)
         );
  OAI21_X1 U4746 ( .B1(n4102), .B2(n4185), .A(n4101), .ZN(n4103) );
  AOI21_X1 U4747 ( .B1(n4104), .B2(n4175), .A(n4103), .ZN(n4249) );
  XOR2_X1 U4748 ( .A(n4106), .B(n4105), .Z(n4248) );
  NAND2_X1 U4749 ( .A1(n4248), .A2(n4107), .ZN(n4115) );
  OAI21_X1 U4750 ( .B1(n4859), .B2(n4109), .A(n4108), .ZN(n4251) );
  INV_X1 U4751 ( .A(n4251), .ZN(n4113) );
  OAI22_X1 U4752 ( .A1(n4350), .A2(n4111), .B1(n4110), .B2(n4197), .ZN(n4112)
         );
  AOI21_X1 U4753 ( .B1(n4113), .B2(n4461), .A(n4112), .ZN(n4114) );
  OAI211_X1 U4754 ( .C1(n4465), .C2(n4249), .A(n4115), .B(n4114), .ZN(U3269)
         );
  XOR2_X1 U4755 ( .A(n4121), .B(n4116), .Z(n4253) );
  INV_X1 U4756 ( .A(n4253), .ZN(n4135) );
  NOR3_X1 U4757 ( .A1(n4183), .A2(n4142), .A3(n4117), .ZN(n4119) );
  NOR2_X1 U4758 ( .A1(n4119), .A2(n4118), .ZN(n4120) );
  XOR2_X1 U4759 ( .A(n4121), .B(n4120), .Z(n4126) );
  AOI22_X1 U4760 ( .A1(n4123), .A2(n4169), .B1(n4122), .B2(n4217), .ZN(n4125)
         );
  NAND2_X1 U4761 ( .A1(n4170), .A2(n4188), .ZN(n4124) );
  OAI211_X1 U4762 ( .C1(n4126), .C2(n4190), .A(n4125), .B(n4124), .ZN(n4252)
         );
  OAI21_X1 U4764 ( .B1(n4154), .B2(n4129), .A(n4857), .ZN(n4301) );
  NOR2_X1 U4765 ( .A1(n4301), .A2(n4195), .ZN(n4133) );
  INV_X1 U4766 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4131) );
  OAI22_X1 U4767 ( .A1(n4350), .A2(n4131), .B1(n4130), .B2(n4197), .ZN(n4132)
         );
  AOI211_X1 U4768 ( .C1(n4252), .C2(n4350), .A(n4133), .B(n4132), .ZN(n4134)
         );
  OAI21_X1 U4769 ( .B1(n4135), .B2(n4203), .A(n4134), .ZN(U3270) );
  XNOR2_X1 U4770 ( .A(n4137), .B(n4136), .ZN(n4256) );
  INV_X1 U4771 ( .A(n4256), .ZN(n4160) );
  OAI22_X1 U4772 ( .A1(n4139), .A2(n4185), .B1(n4207), .B2(n4138), .ZN(n4149)
         );
  INV_X1 U4773 ( .A(n4140), .ZN(n4141) );
  OAI21_X1 U4774 ( .B1(n4183), .B2(n4142), .A(n4141), .ZN(n4167) );
  OAI21_X1 U4775 ( .B1(n4167), .B2(n4144), .A(n4143), .ZN(n4146) );
  XNOR2_X1 U4776 ( .A(n4146), .B(n4145), .ZN(n4147) );
  NOR2_X1 U4777 ( .A1(n4147), .A2(n4190), .ZN(n4148) );
  AOI211_X1 U4778 ( .C1(n4188), .C2(n4150), .A(n4149), .B(n4148), .ZN(n4151)
         );
  INV_X1 U4779 ( .A(n4151), .ZN(n4255) );
  AND2_X1 U4780 ( .A1(n4153), .A2(n4152), .ZN(n4155) );
  OR2_X1 U4781 ( .A1(n4155), .A2(n4154), .ZN(n4305) );
  AOI22_X1 U4782 ( .A1(n4465), .A2(REG2_REG_19__SCAN_IN), .B1(n4156), .B2(
        n4457), .ZN(n4157) );
  OAI21_X1 U4783 ( .B1(n4305), .B2(n4195), .A(n4157), .ZN(n4158) );
  AOI21_X1 U4784 ( .B1(n4255), .B2(n4350), .A(n4158), .ZN(n4159) );
  OAI21_X1 U4785 ( .B1(n4160), .B2(n4203), .A(n4159), .ZN(U3271) );
  OAI21_X1 U4786 ( .B1(n4162), .B2(n4168), .A(n4161), .ZN(n4163) );
  INV_X1 U4787 ( .A(n4163), .ZN(n4260) );
  XNOR2_X1 U4788 ( .A(n4192), .B(n4164), .ZN(n4165) );
  NAND2_X1 U4789 ( .A1(n4165), .A2(n4510), .ZN(n4258) );
  INV_X1 U4790 ( .A(n4258), .ZN(n4180) );
  INV_X1 U4791 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4166) );
  OAI22_X1 U4792 ( .A1(n4350), .A2(n4166), .B1(n4341), .B2(n4197), .ZN(n4178)
         );
  XOR2_X1 U4793 ( .A(n4168), .B(n4167), .Z(n4176) );
  AOI22_X1 U4794 ( .A1(n4170), .A2(n4169), .B1(n4217), .B2(n4328), .ZN(n4171)
         );
  OAI21_X1 U4795 ( .B1(n4173), .B2(n4172), .A(n4171), .ZN(n4174) );
  AOI21_X1 U4796 ( .B1(n4176), .B2(n4175), .A(n4174), .ZN(n4259) );
  NOR2_X1 U4797 ( .A1(n4259), .A2(n4465), .ZN(n4177) );
  AOI211_X1 U4798 ( .C1(n4180), .C2(n4179), .A(n4178), .B(n4177), .ZN(n4181)
         );
  OAI21_X1 U4799 ( .B1(n4260), .B2(n4203), .A(n4181), .ZN(U3272) );
  XOR2_X1 U4800 ( .A(n4184), .B(n4182), .Z(n4262) );
  INV_X1 U4801 ( .A(n4262), .ZN(n4204) );
  XOR2_X1 U4802 ( .A(n4184), .B(n4183), .Z(n4191) );
  OAI22_X1 U4803 ( .A1(n2304), .A2(n4185), .B1(n4207), .B2(n4193), .ZN(n4186)
         );
  AOI21_X1 U4804 ( .B1(n4188), .B2(n4187), .A(n4186), .ZN(n4189) );
  OAI21_X1 U4805 ( .B1(n4191), .B2(n4190), .A(n4189), .ZN(n4261) );
  OAI21_X1 U4806 ( .B1(n4194), .B2(n4193), .A(n4192), .ZN(n4311) );
  NOR2_X1 U4807 ( .A1(n4311), .A2(n4195), .ZN(n4201) );
  INV_X1 U4808 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4199) );
  INV_X1 U4809 ( .A(n4196), .ZN(n4198) );
  OAI22_X1 U4810 ( .A1(n4350), .A2(n4199), .B1(n4198), .B2(n4197), .ZN(n4200)
         );
  AOI211_X1 U4811 ( .C1(n4261), .C2(n4350), .A(n4201), .B(n4200), .ZN(n4202)
         );
  OAI21_X1 U4812 ( .B1(n4204), .B2(n4203), .A(n4202), .ZN(U3273) );
  NAND2_X1 U4813 ( .A1(n4212), .A2(n4211), .ZN(n4214) );
  XNOR2_X1 U4814 ( .A(n4214), .B(n4208), .ZN(n4344) );
  NAND2_X1 U4815 ( .A1(n4344), .A2(n4215), .ZN(n4210) );
  NAND2_X1 U4816 ( .A1(n4206), .A2(n4205), .ZN(n4219) );
  OAI21_X1 U4817 ( .B1(n4208), .B2(n4207), .A(n4219), .ZN(n4343) );
  NAND2_X1 U4818 ( .A1(n4537), .A2(n4343), .ZN(n4209) );
  OAI211_X1 U4819 ( .C1(n4537), .C2(n3728), .A(n4210), .B(n4209), .ZN(U3549)
         );
  OR2_X1 U4820 ( .A1(n4212), .A2(n4211), .ZN(n4213) );
  NAND2_X1 U4821 ( .A1(n4348), .A2(n4215), .ZN(n4221) );
  NAND2_X1 U4822 ( .A1(n4217), .A2(n4216), .ZN(n4218) );
  NAND2_X1 U4823 ( .A1(n4219), .A2(n4218), .ZN(n4346) );
  NAND2_X1 U4824 ( .A1(n4537), .A2(n4346), .ZN(n4220) );
  OAI211_X1 U4825 ( .C1(n4537), .C2(n2423), .A(n4221), .B(n4220), .ZN(U3548)
         );
  MUX2_X1 U4826 ( .A(REG1_REG_29__SCAN_IN), .B(n4280), .S(n4537), .Z(U3547) );
  INV_X1 U4827 ( .A(n4510), .ZN(n4516) );
  NAND2_X1 U4828 ( .A1(n4225), .A2(n4508), .ZN(n4227) );
  OAI211_X1 U4829 ( .C1(n4516), .C2(n4228), .A(n4227), .B(n4226), .ZN(n4281)
         );
  MUX2_X1 U4830 ( .A(REG1_REG_27__SCAN_IN), .B(n4281), .S(n4537), .Z(U3545) );
  AOI21_X1 U4831 ( .B1(n4230), .B2(n4508), .A(n4229), .ZN(n4282) );
  MUX2_X1 U4832 ( .A(n4231), .B(n4282), .S(n4537), .Z(n4232) );
  OAI21_X1 U4833 ( .B1(n4264), .B2(n4284), .A(n4232), .ZN(U3544) );
  AOI21_X1 U4834 ( .B1(n4234), .B2(n4508), .A(n4233), .ZN(n4285) );
  MUX2_X1 U4835 ( .A(n4235), .B(n4285), .S(n4537), .Z(n4236) );
  OAI21_X1 U4836 ( .B1(n4264), .B2(n4288), .A(n4236), .ZN(U3543) );
  AOI21_X1 U4837 ( .B1(n4238), .B2(n4508), .A(n4237), .ZN(n4289) );
  MUX2_X1 U4838 ( .A(n4790), .B(n4289), .S(n4537), .Z(n4239) );
  OAI21_X1 U4839 ( .B1(n4264), .B2(n4292), .A(n4239), .ZN(U3542) );
  AOI21_X1 U4840 ( .B1(n4241), .B2(n4508), .A(n4240), .ZN(n4293) );
  MUX2_X1 U4841 ( .A(n4788), .B(n4293), .S(n4537), .Z(n4242) );
  OAI21_X1 U4842 ( .B1(n4264), .B2(n4295), .A(n4242), .ZN(U3541) );
  INV_X1 U4843 ( .A(n4508), .ZN(n4497) );
  NAND3_X1 U4844 ( .A1(n4244), .A2(n4510), .A3(n4243), .ZN(n4245) );
  OAI211_X1 U4845 ( .C1(n4247), .C2(n4497), .A(n4246), .B(n4245), .ZN(n4296)
         );
  MUX2_X1 U4846 ( .A(REG1_REG_22__SCAN_IN), .B(n4296), .S(n4537), .Z(U3540) );
  NAND2_X1 U4847 ( .A1(n4248), .A2(n4508), .ZN(n4250) );
  OAI211_X1 U4848 ( .C1(n4516), .C2(n4251), .A(n4250), .B(n4249), .ZN(n4297)
         );
  MUX2_X1 U4849 ( .A(REG1_REG_21__SCAN_IN), .B(n4297), .S(n4537), .Z(U3539) );
  INV_X1 U4850 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4786) );
  AOI21_X1 U4851 ( .B1(n4253), .B2(n4508), .A(n4252), .ZN(n4298) );
  MUX2_X1 U4852 ( .A(n4786), .B(n4298), .S(n4537), .Z(n4254) );
  OAI21_X1 U4853 ( .B1(n4264), .B2(n4301), .A(n4254), .ZN(U3538) );
  INV_X1 U4854 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4574) );
  AOI21_X1 U4855 ( .B1(n4256), .B2(n4508), .A(n4255), .ZN(n4302) );
  MUX2_X1 U4856 ( .A(n4574), .B(n4302), .S(n4537), .Z(n4257) );
  OAI21_X1 U4857 ( .B1(n4264), .B2(n4305), .A(n4257), .ZN(U3537) );
  OAI211_X1 U4858 ( .C1(n4260), .C2(n4497), .A(n4259), .B(n4258), .ZN(n4306)
         );
  MUX2_X1 U4859 ( .A(REG1_REG_18__SCAN_IN), .B(n4306), .S(n4537), .Z(U3536) );
  INV_X1 U4860 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4605) );
  AOI21_X1 U4861 ( .B1(n4262), .B2(n4508), .A(n4261), .ZN(n4307) );
  MUX2_X1 U4862 ( .A(n4605), .B(n4307), .S(n4537), .Z(n4263) );
  OAI21_X1 U4863 ( .B1(n4264), .B2(n4311), .A(n4263), .ZN(U3535) );
  AOI21_X1 U4864 ( .B1(n4510), .B2(n4266), .A(n4265), .ZN(n4267) );
  OAI21_X1 U4865 ( .B1(n4268), .B2(n4497), .A(n4267), .ZN(n4312) );
  MUX2_X1 U4866 ( .A(REG1_REG_16__SCAN_IN), .B(n4312), .S(n4537), .Z(U3534) );
  AOI21_X1 U4867 ( .B1(n4510), .B2(n4270), .A(n4269), .ZN(n4271) );
  OAI21_X1 U4868 ( .B1(n4272), .B2(n4497), .A(n4271), .ZN(n4313) );
  MUX2_X1 U4869 ( .A(REG1_REG_15__SCAN_IN), .B(n4313), .S(n4537), .Z(U3533) );
  INV_X1 U4870 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4275) );
  NAND2_X1 U4871 ( .A1(n4344), .A2(n4276), .ZN(n4274) );
  NAND2_X1 U4872 ( .A1(n4524), .A2(n4343), .ZN(n4273) );
  OAI211_X1 U4873 ( .C1(n4524), .C2(n4275), .A(n4274), .B(n4273), .ZN(U3517)
         );
  INV_X1 U4874 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4279) );
  NAND2_X1 U4875 ( .A1(n4348), .A2(n4276), .ZN(n4278) );
  NAND2_X1 U4876 ( .A1(n4524), .A2(n4346), .ZN(n4277) );
  OAI211_X1 U4877 ( .C1(n4524), .C2(n4279), .A(n4278), .B(n4277), .ZN(U3516)
         );
  MUX2_X1 U4878 ( .A(REG0_REG_29__SCAN_IN), .B(n4280), .S(n4524), .Z(U3515) );
  MUX2_X1 U4879 ( .A(REG0_REG_27__SCAN_IN), .B(n4281), .S(n4524), .Z(U3513) );
  INV_X1 U4880 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4801) );
  MUX2_X1 U4881 ( .A(n4801), .B(n4282), .S(n4524), .Z(n4283) );
  OAI21_X1 U4882 ( .B1(n4284), .B2(n4310), .A(n4283), .ZN(U3512) );
  INV_X1 U4883 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4286) );
  MUX2_X1 U4884 ( .A(n4286), .B(n4285), .S(n4524), .Z(n4287) );
  OAI21_X1 U4885 ( .B1(n4288), .B2(n4310), .A(n4287), .ZN(U3511) );
  INV_X1 U4886 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4290) );
  MUX2_X1 U4887 ( .A(n4290), .B(n4289), .S(n4524), .Z(n4291) );
  OAI21_X1 U4888 ( .B1(n4292), .B2(n4310), .A(n4291), .ZN(U3510) );
  INV_X1 U4889 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4791) );
  MUX2_X1 U4890 ( .A(n4791), .B(n4293), .S(n4524), .Z(n4294) );
  OAI21_X1 U4891 ( .B1(n4295), .B2(n4310), .A(n4294), .ZN(U3509) );
  MUX2_X1 U4892 ( .A(REG0_REG_22__SCAN_IN), .B(n4296), .S(n4524), .Z(U3508) );
  MUX2_X1 U4893 ( .A(REG0_REG_21__SCAN_IN), .B(n4297), .S(n4524), .Z(U3507) );
  INV_X1 U4894 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4299) );
  MUX2_X1 U4895 ( .A(n4299), .B(n4298), .S(n4524), .Z(n4300) );
  OAI21_X1 U4896 ( .B1(n4301), .B2(n4310), .A(n4300), .ZN(U3506) );
  INV_X1 U4897 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4303) );
  MUX2_X1 U4898 ( .A(n4303), .B(n4302), .S(n4524), .Z(n4304) );
  OAI21_X1 U4899 ( .B1(n4305), .B2(n4310), .A(n4304), .ZN(U3505) );
  MUX2_X1 U4900 ( .A(REG0_REG_18__SCAN_IN), .B(n4306), .S(n4524), .Z(U3503) );
  INV_X1 U4901 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4308) );
  MUX2_X1 U4902 ( .A(n4308), .B(n4307), .S(n4524), .Z(n4309) );
  OAI21_X1 U4903 ( .B1(n4311), .B2(n4310), .A(n4309), .ZN(U3501) );
  MUX2_X1 U4904 ( .A(REG0_REG_16__SCAN_IN), .B(n4312), .S(n4524), .Z(U3499) );
  MUX2_X1 U4905 ( .A(REG0_REG_15__SCAN_IN), .B(n4313), .S(n4524), .Z(U3497) );
  MUX2_X1 U4906 ( .A(n4314), .B(DATAI_28_), .S(U3149), .Z(U3324) );
  MUX2_X1 U4907 ( .A(n4353), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U4908 ( .A(DATAI_24_), .B(n2401), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U4909 ( .A(DATAI_22_), .B(n4315), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U4910 ( .A(DATAI_19_), .B(n4316), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U4911 ( .A(n4317), .B(DATAI_17_), .S(U3149), .Z(U3335) );
  MUX2_X1 U4912 ( .A(DATAI_14_), .B(n4406), .S(STATE_REG_SCAN_IN), .Z(U3338)
         );
  MUX2_X1 U4913 ( .A(n4318), .B(DATAI_13_), .S(U3149), .Z(U3339) );
  MUX2_X1 U4914 ( .A(n4319), .B(DATAI_10_), .S(U3149), .Z(U3342) );
  MUX2_X1 U4915 ( .A(DATAI_8_), .B(n4320), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U4916 ( .A(n4321), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U4917 ( .A(n4322), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U4918 ( .A(DATAI_3_), .B(n4323), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U4919 ( .A(n4324), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4920 ( .A(n4325), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  AOI22_X1 U4921 ( .A1(n4329), .A2(n4328), .B1(n4327), .B2(n4326), .ZN(n4340)
         );
  NOR2_X1 U4922 ( .A1(n4331), .A2(n2265), .ZN(n4332) );
  XNOR2_X1 U4923 ( .A(n2150), .B(n4332), .ZN(n4338) );
  NOR2_X1 U4924 ( .A1(STATE_REG_SCAN_IN), .A2(n4333), .ZN(n4436) );
  NOR2_X1 U4925 ( .A1(n4335), .A2(n4334), .ZN(n4336) );
  AOI211_X1 U4926 ( .C1(n4338), .C2(n4337), .A(n4436), .B(n4336), .ZN(n4339)
         );
  OAI211_X1 U4927 ( .C1(n4342), .C2(n4341), .A(n4340), .B(n4339), .ZN(U3235)
         );
  INV_X1 U4928 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4559) );
  AOI22_X1 U4929 ( .A1(n4344), .A2(n4461), .B1(n4350), .B2(n4343), .ZN(n4345)
         );
  OAI21_X1 U4930 ( .B1(n4350), .B2(n4559), .A(n4345), .ZN(U3260) );
  INV_X1 U4931 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4557) );
  AOI22_X1 U4932 ( .A1(n4348), .A2(n4461), .B1(n4350), .B2(n4346), .ZN(n4349)
         );
  OAI21_X1 U4933 ( .B1(n4557), .B2(n4350), .A(n4349), .ZN(U3261) );
  INV_X1 U4934 ( .A(n4351), .ZN(n4352) );
  OAI21_X1 U4935 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4353), .A(n4352), .ZN(n4354)
         );
  XNOR2_X1 U4936 ( .A(n4354), .B(n4547), .ZN(n4357) );
  AOI22_X1 U4937 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4437), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4355) );
  OAI21_X1 U4938 ( .B1(n4357), .B2(n4356), .A(n4355), .ZN(U3240) );
  XOR2_X1 U4939 ( .A(n4358), .B(REG2_REG_4__SCAN_IN), .Z(n4366) );
  XNOR2_X1 U4940 ( .A(n4359), .B(REG1_REG_4__SCAN_IN), .ZN(n4364) );
  NOR2_X1 U4941 ( .A1(n4449), .A2(n4360), .ZN(n4361) );
  AOI211_X1 U4942 ( .C1(n4437), .C2(ADDR_REG_4__SCAN_IN), .A(n4362), .B(n4361), 
        .ZN(n4363) );
  OAI21_X1 U4943 ( .B1(n4364), .B2(n4433), .A(n4363), .ZN(n4365) );
  AOI21_X1 U4944 ( .B1(n4445), .B2(n4366), .A(n4365), .ZN(n4368) );
  NAND2_X1 U4945 ( .A1(n4368), .A2(n4367), .ZN(U3244) );
  AOI211_X1 U4946 ( .C1(n4371), .C2(n4370), .A(n4369), .B(n4433), .ZN(n4373)
         );
  AOI211_X1 U4947 ( .C1(n4437), .C2(ADDR_REG_9__SCAN_IN), .A(n4373), .B(n4372), 
        .ZN(n4378) );
  OAI211_X1 U4948 ( .C1(n4376), .C2(n4375), .A(n4445), .B(n4374), .ZN(n4377)
         );
  OAI211_X1 U4949 ( .C1(n4449), .C2(n4476), .A(n4378), .B(n4377), .ZN(U3249)
         );
  AOI211_X1 U4950 ( .C1(n4381), .C2(n4380), .A(n4379), .B(n4433), .ZN(n4383)
         );
  AOI211_X1 U4951 ( .C1(n4437), .C2(ADDR_REG_11__SCAN_IN), .A(n4383), .B(n4382), .ZN(n4388) );
  OAI211_X1 U4952 ( .C1(n4386), .C2(n4385), .A(n4445), .B(n4384), .ZN(n4387)
         );
  OAI211_X1 U4953 ( .C1(n4449), .C2(n4475), .A(n4388), .B(n4387), .ZN(U3251)
         );
  AOI211_X1 U4954 ( .C1(n4633), .C2(n4390), .A(n4389), .B(n4433), .ZN(n4393)
         );
  INV_X1 U4955 ( .A(n4391), .ZN(n4392) );
  AOI211_X1 U4956 ( .C1(n4437), .C2(ADDR_REG_12__SCAN_IN), .A(n4393), .B(n4392), .ZN(n4397) );
  OAI211_X1 U4957 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4395), .A(n4445), .B(n4394), .ZN(n4396) );
  OAI211_X1 U4958 ( .C1(n4449), .C2(n4474), .A(n4397), .B(n4396), .ZN(U3252)
         );
  INV_X1 U4959 ( .A(ADDR_REG_14__SCAN_IN), .ZN(n4809) );
  AOI211_X1 U4960 ( .C1(n4400), .C2(n4641), .A(n4399), .B(n4398), .ZN(n4405)
         );
  AOI211_X1 U4961 ( .C1(n4403), .C2(n4402), .A(n4401), .B(n4433), .ZN(n4404)
         );
  AOI211_X1 U4962 ( .C1(n4407), .C2(n4406), .A(n4405), .B(n4404), .ZN(n4409)
         );
  OAI211_X1 U4963 ( .C1(n4410), .C2(n4809), .A(n4409), .B(n4408), .ZN(U3254)
         );
  AOI211_X1 U4964 ( .C1(n4413), .C2(n4412), .A(n4411), .B(n4433), .ZN(n4414)
         );
  AOI211_X1 U4965 ( .C1(n4437), .C2(ADDR_REG_15__SCAN_IN), .A(n4415), .B(n4414), .ZN(n4421) );
  AOI21_X1 U4966 ( .B1(n4418), .B2(n4417), .A(n4416), .ZN(n4419) );
  NAND2_X1 U4967 ( .A1(n4445), .A2(n4419), .ZN(n4420) );
  OAI211_X1 U4968 ( .C1(n4449), .C2(n4473), .A(n4421), .B(n4420), .ZN(U3255)
         );
  INV_X1 U4969 ( .A(n4422), .ZN(n4423) );
  AOI21_X1 U4970 ( .B1(n4437), .B2(ADDR_REG_16__SCAN_IN), .A(n4423), .ZN(n4432) );
  OAI21_X1 U4971 ( .B1(n4425), .B2(n3348), .A(n4424), .ZN(n4430) );
  OAI21_X1 U4972 ( .B1(n4427), .B2(n4774), .A(n4426), .ZN(n4428) );
  AOI22_X1 U4973 ( .A1(n4445), .A2(n4430), .B1(n4429), .B2(n4428), .ZN(n4431)
         );
  OAI211_X1 U4974 ( .C1(n4472), .C2(n4449), .A(n4432), .B(n4431), .ZN(U3256)
         );
  AOI21_X1 U4975 ( .B1(n4443), .B2(n4442), .A(n4441), .ZN(n4444) );
  NAND2_X1 U4976 ( .A1(n4445), .A2(n4444), .ZN(n4446) );
  OAI211_X1 U4977 ( .C1(n4449), .C2(n4448), .A(n4447), .B(n4446), .ZN(U3258)
         );
  AOI22_X1 U4978 ( .A1(n4465), .A2(REG2_REG_6__SCAN_IN), .B1(n4450), .B2(n4457), .ZN(n4455) );
  INV_X1 U4979 ( .A(n4451), .ZN(n4453) );
  AOI22_X1 U4980 ( .A1(n4453), .A2(n4459), .B1(n4461), .B2(n4452), .ZN(n4454)
         );
  OAI211_X1 U4981 ( .C1(n4465), .C2(n4456), .A(n4455), .B(n4454), .ZN(U3284)
         );
  AOI22_X1 U4982 ( .A1(REG2_REG_2__SCAN_IN), .A2(n4465), .B1(
        REG3_REG_2__SCAN_IN), .B2(n4457), .ZN(n4463) );
  AOI22_X1 U4983 ( .A1(n4461), .A2(n4460), .B1(n4459), .B2(n4458), .ZN(n4462)
         );
  OAI211_X1 U4984 ( .C1(n4465), .C2(n4464), .A(n4463), .B(n4462), .ZN(U3288)
         );
  AND2_X1 U4985 ( .A1(D_REG_31__SCAN_IN), .A2(n4467), .ZN(U3291) );
  INV_X1 U4986 ( .A(D_REG_30__SCAN_IN), .ZN(n4751) );
  NOR2_X1 U4987 ( .A1(n4466), .A2(n4751), .ZN(U3292) );
  AND2_X1 U4988 ( .A1(D_REG_29__SCAN_IN), .A2(n4467), .ZN(U3293) );
  INV_X1 U4989 ( .A(D_REG_28__SCAN_IN), .ZN(n4769) );
  NOR2_X1 U4990 ( .A1(n4466), .A2(n4769), .ZN(U3294) );
  AND2_X1 U4991 ( .A1(D_REG_27__SCAN_IN), .A2(n4467), .ZN(U3295) );
  INV_X1 U4992 ( .A(D_REG_26__SCAN_IN), .ZN(n4760) );
  NOR2_X1 U4993 ( .A1(n4466), .A2(n4760), .ZN(U3296) );
  INV_X1 U4994 ( .A(D_REG_25__SCAN_IN), .ZN(n4775) );
  NOR2_X1 U4995 ( .A1(n4466), .A2(n4775), .ZN(U3297) );
  AND2_X1 U4996 ( .A1(D_REG_24__SCAN_IN), .A2(n4467), .ZN(U3298) );
  AND2_X1 U4997 ( .A1(D_REG_23__SCAN_IN), .A2(n4467), .ZN(U3299) );
  AND2_X1 U4998 ( .A1(D_REG_22__SCAN_IN), .A2(n4467), .ZN(U3300) );
  INV_X1 U4999 ( .A(D_REG_21__SCAN_IN), .ZN(n4759) );
  NOR2_X1 U5000 ( .A1(n4466), .A2(n4759), .ZN(U3301) );
  INV_X1 U5001 ( .A(D_REG_20__SCAN_IN), .ZN(n4765) );
  NOR2_X1 U5002 ( .A1(n4466), .A2(n4765), .ZN(U3302) );
  INV_X1 U5003 ( .A(D_REG_19__SCAN_IN), .ZN(n4749) );
  NOR2_X1 U5004 ( .A1(n4466), .A2(n4749), .ZN(U3303) );
  INV_X1 U5005 ( .A(D_REG_18__SCAN_IN), .ZN(n4768) );
  NOR2_X1 U5006 ( .A1(n4466), .A2(n4768), .ZN(U3304) );
  AND2_X1 U5007 ( .A1(D_REG_17__SCAN_IN), .A2(n4467), .ZN(U3305) );
  INV_X1 U5008 ( .A(D_REG_16__SCAN_IN), .ZN(n4756) );
  NOR2_X1 U5009 ( .A1(n4466), .A2(n4756), .ZN(U3306) );
  AND2_X1 U5010 ( .A1(D_REG_15__SCAN_IN), .A2(n4467), .ZN(U3307) );
  INV_X1 U5011 ( .A(D_REG_14__SCAN_IN), .ZN(n4772) );
  NOR2_X1 U5012 ( .A1(n4466), .A2(n4772), .ZN(U3308) );
  AND2_X1 U5013 ( .A1(D_REG_13__SCAN_IN), .A2(n4467), .ZN(U3309) );
  INV_X1 U5014 ( .A(D_REG_12__SCAN_IN), .ZN(n4757) );
  NOR2_X1 U5015 ( .A1(n4466), .A2(n4757), .ZN(U3310) );
  AND2_X1 U5016 ( .A1(D_REG_11__SCAN_IN), .A2(n4467), .ZN(U3311) );
  AND2_X1 U5017 ( .A1(D_REG_10__SCAN_IN), .A2(n4467), .ZN(U3312) );
  AND2_X1 U5018 ( .A1(D_REG_9__SCAN_IN), .A2(n4467), .ZN(U3313) );
  INV_X1 U5019 ( .A(D_REG_8__SCAN_IN), .ZN(n4748) );
  NOR2_X1 U5020 ( .A1(n4466), .A2(n4748), .ZN(U3314) );
  INV_X1 U5021 ( .A(D_REG_7__SCAN_IN), .ZN(n4771) );
  NOR2_X1 U5022 ( .A1(n4466), .A2(n4771), .ZN(U3315) );
  AND2_X1 U5023 ( .A1(D_REG_6__SCAN_IN), .A2(n4467), .ZN(U3316) );
  AND2_X1 U5024 ( .A1(D_REG_5__SCAN_IN), .A2(n4467), .ZN(U3317) );
  AND2_X1 U5025 ( .A1(D_REG_4__SCAN_IN), .A2(n4467), .ZN(U3318) );
  INV_X1 U5026 ( .A(D_REG_3__SCAN_IN), .ZN(n4766) );
  NOR2_X1 U5027 ( .A1(n4466), .A2(n4766), .ZN(U3319) );
  AND2_X1 U5028 ( .A1(D_REG_2__SCAN_IN), .A2(n4467), .ZN(U3320) );
  INV_X1 U5029 ( .A(DATAI_23_), .ZN(n4541) );
  AOI21_X1 U5030 ( .B1(U3149), .B2(n4541), .A(n4468), .ZN(U3329) );
  OAI22_X1 U5031 ( .A1(U3149), .A2(n4469), .B1(DATAI_18_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4470) );
  INV_X1 U5032 ( .A(n4470), .ZN(U3334) );
  AOI22_X1 U5033 ( .A1(STATE_REG_SCAN_IN), .A2(n4472), .B1(n4471), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5034 ( .A(DATAI_15_), .ZN(n4642) );
  AOI22_X1 U5035 ( .A1(STATE_REG_SCAN_IN), .A2(n4473), .B1(n4642), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5036 ( .A(DATAI_12_), .ZN(n4736) );
  AOI22_X1 U5037 ( .A1(STATE_REG_SCAN_IN), .A2(n4474), .B1(n4736), .B2(U3149), 
        .ZN(U3340) );
  AOI22_X1 U5038 ( .A1(STATE_REG_SCAN_IN), .A2(n4475), .B1(n3071), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5039 ( .A(DATAI_9_), .ZN(n4818) );
  AOI22_X1 U5040 ( .A1(STATE_REG_SCAN_IN), .A2(n4476), .B1(n4818), .B2(U3149), 
        .ZN(U3343) );
  OAI22_X1 U5041 ( .A1(U3149), .A2(IR_REG_0__SCAN_IN), .B1(DATAI_0_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4477) );
  INV_X1 U5042 ( .A(n4477), .ZN(U3352) );
  OAI211_X1 U5043 ( .C1(n4480), .C2(n4487), .A(n4479), .B(n4478), .ZN(n4481)
         );
  INV_X1 U5044 ( .A(n4481), .ZN(n4526) );
  INV_X1 U5045 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4630) );
  AOI22_X1 U5046 ( .A1(n4524), .A2(n4526), .B1(n4630), .B2(n4522), .ZN(U3467)
         );
  OAI22_X1 U5047 ( .A1(n4483), .A2(n4487), .B1(n4516), .B2(n4482), .ZN(n4484)
         );
  NOR2_X1 U5048 ( .A1(n4485), .A2(n4484), .ZN(n4528) );
  INV_X1 U5049 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4486) );
  AOI22_X1 U5050 ( .A1(n4524), .A2(n4528), .B1(n4486), .B2(n4522), .ZN(U3469)
         );
  NOR2_X1 U5051 ( .A1(n4488), .A2(n4487), .ZN(n4490) );
  AOI211_X1 U5052 ( .C1(n4510), .C2(n4491), .A(n4490), .B(n4489), .ZN(n4529)
         );
  INV_X1 U5053 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4492) );
  AOI22_X1 U5054 ( .A1(n4524), .A2(n4529), .B1(n4492), .B2(n4522), .ZN(U3473)
         );
  INV_X1 U5055 ( .A(n4493), .ZN(n4495) );
  AOI211_X1 U5056 ( .C1(n4496), .C2(n4521), .A(n4495), .B(n4494), .ZN(n4530)
         );
  INV_X1 U5057 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4627) );
  AOI22_X1 U5058 ( .A1(n4524), .A2(n4530), .B1(n4627), .B2(n4522), .ZN(U3475)
         );
  NOR2_X1 U5059 ( .A1(n4498), .A2(n4497), .ZN(n4501) );
  INV_X1 U5060 ( .A(n4499), .ZN(n4500) );
  AOI211_X1 U5061 ( .C1(n4510), .C2(n4502), .A(n4501), .B(n4500), .ZN(n4531)
         );
  INV_X1 U5062 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4626) );
  AOI22_X1 U5063 ( .A1(n4524), .A2(n4531), .B1(n4626), .B2(n4522), .ZN(U3477)
         );
  NAND3_X1 U5064 ( .A1(n3051), .A2(n4503), .A3(n4508), .ZN(n4504) );
  AND3_X1 U5065 ( .A1(n4506), .A2(n4505), .A3(n4504), .ZN(n4532) );
  INV_X1 U5066 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4507) );
  AOI22_X1 U5067 ( .A1(n4524), .A2(n4532), .B1(n4507), .B2(n4522), .ZN(U3481)
         );
  NAND2_X1 U5068 ( .A1(n4509), .A2(n4508), .ZN(n4514) );
  NAND2_X1 U5069 ( .A1(n4511), .A2(n4510), .ZN(n4512) );
  AND3_X1 U5070 ( .A1(n4514), .A2(n4513), .A3(n4512), .ZN(n4533) );
  INV_X1 U5071 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4515) );
  AOI22_X1 U5072 ( .A1(n4524), .A2(n4533), .B1(n4515), .B2(n4522), .ZN(U3485)
         );
  NOR2_X1 U5073 ( .A1(n4517), .A2(n4516), .ZN(n4519) );
  AOI211_X1 U5074 ( .C1(n4521), .C2(n4520), .A(n4519), .B(n4518), .ZN(n4536)
         );
  INV_X1 U5075 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4523) );
  AOI22_X1 U5076 ( .A1(n4524), .A2(n4536), .B1(n4523), .B2(n4522), .ZN(U3489)
         );
  AOI22_X1 U5077 ( .A1(n4537), .A2(n4526), .B1(n4525), .B2(n4534), .ZN(U3518)
         );
  AOI22_X1 U5078 ( .A1(n4537), .A2(n4528), .B1(n4527), .B2(n4534), .ZN(U3519)
         );
  AOI22_X1 U5079 ( .A1(n4537), .A2(n4529), .B1(n2434), .B2(n4534), .ZN(U3521)
         );
  AOI22_X1 U5080 ( .A1(n4537), .A2(n4530), .B1(n2222), .B2(n4534), .ZN(U3522)
         );
  AOI22_X1 U5081 ( .A1(n4537), .A2(n4531), .B1(n4606), .B2(n4534), .ZN(U3523)
         );
  AOI22_X1 U5082 ( .A1(n4537), .A2(n4532), .B1(n4601), .B2(n4534), .ZN(U3525)
         );
  AOI22_X1 U5083 ( .A1(n4537), .A2(n4533), .B1(n4602), .B2(n4534), .ZN(U3527)
         );
  AOI22_X1 U5084 ( .A1(n4537), .A2(n4536), .B1(n4535), .B2(n4534), .ZN(U3529)
         );
  NAND2_X1 U5085 ( .A1(n2304), .A2(U4043), .ZN(n4538) );
  OAI21_X1 U5086 ( .B1(U4043), .B2(DATAO_REG_18__SCAN_IN), .A(n4538), .ZN(
        n4854) );
  AOI22_X1 U5087 ( .A1(n4541), .A2(keyinput40), .B1(keyinput82), .B2(n4540), 
        .ZN(n4539) );
  OAI221_X1 U5088 ( .B1(n4541), .B2(keyinput40), .C1(n4540), .C2(keyinput82), 
        .A(n4539), .ZN(n4554) );
  INV_X1 U5089 ( .A(DATAI_27_), .ZN(n4544) );
  AOI22_X1 U5090 ( .A1(n4544), .A2(keyinput114), .B1(keyinput2), .B2(n4543), 
        .ZN(n4542) );
  OAI221_X1 U5091 ( .B1(n4544), .B2(keyinput114), .C1(n4543), .C2(keyinput2), 
        .A(n4542), .ZN(n4553) );
  INV_X1 U5092 ( .A(keyinput20), .ZN(n4546) );
  AOI22_X1 U5093 ( .A1(n4547), .A2(keyinput72), .B1(ADDR_REG_0__SCAN_IN), .B2(
        n4546), .ZN(n4545) );
  OAI221_X1 U5094 ( .B1(n4547), .B2(keyinput72), .C1(n4546), .C2(
        ADDR_REG_0__SCAN_IN), .A(n4545), .ZN(n4552) );
  AOI22_X1 U5095 ( .A1(n4550), .A2(keyinput6), .B1(n4549), .B2(keyinput15), 
        .ZN(n4548) );
  OAI221_X1 U5096 ( .B1(n4550), .B2(keyinput6), .C1(n4549), .C2(keyinput15), 
        .A(n4548), .ZN(n4551) );
  NOR4_X1 U5097 ( .A1(n4554), .A2(n4553), .A3(n4552), .A4(n4551), .ZN(n4852)
         );
  INV_X1 U5098 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4556) );
  AOI22_X1 U5099 ( .A1(n4557), .A2(keyinput17), .B1(n4556), .B2(keyinput1), 
        .ZN(n4555) );
  OAI221_X1 U5100 ( .B1(n4557), .B2(keyinput17), .C1(n4556), .C2(keyinput1), 
        .A(n4555), .ZN(n4567) );
  INV_X1 U5101 ( .A(B_REG_SCAN_IN), .ZN(n4560) );
  AOI22_X1 U5102 ( .A1(n4560), .A2(keyinput93), .B1(keyinput83), .B2(n4559), 
        .ZN(n4558) );
  OAI221_X1 U5103 ( .B1(n4560), .B2(keyinput93), .C1(n4559), .C2(keyinput83), 
        .A(n4558), .ZN(n4566) );
  INV_X1 U5104 ( .A(DATAI_28_), .ZN(n4562) );
  AOI22_X1 U5105 ( .A1(n4111), .A2(keyinput102), .B1(n4562), .B2(keyinput81), 
        .ZN(n4561) );
  OAI221_X1 U5106 ( .B1(n4111), .B2(keyinput102), .C1(n4562), .C2(keyinput81), 
        .A(n4561), .ZN(n4565) );
  AOI22_X1 U5107 ( .A1(n4076), .A2(keyinput123), .B1(keyinput106), .B2(n4093), 
        .ZN(n4563) );
  OAI221_X1 U5108 ( .B1(n4076), .B2(keyinput123), .C1(n4093), .C2(keyinput106), 
        .A(n4563), .ZN(n4564) );
  NOR4_X1 U5109 ( .A1(n4567), .A2(n4566), .A3(n4565), .A4(n4564), .ZN(n4851)
         );
  INV_X1 U5110 ( .A(keyinput33), .ZN(n4569) );
  AOI22_X1 U5111 ( .A1(n2434), .A2(keyinput86), .B1(DATAO_REG_4__SCAN_IN), 
        .B2(n4569), .ZN(n4568) );
  OAI221_X1 U5112 ( .B1(n2434), .B2(keyinput86), .C1(n4569), .C2(
        DATAO_REG_4__SCAN_IN), .A(n4568), .ZN(n4660) );
  INV_X1 U5113 ( .A(DATAI_25_), .ZN(n4571) );
  AOI22_X1 U5114 ( .A1(U3149), .A2(keyinput113), .B1(keyinput66), .B2(n4571), 
        .ZN(n4570) );
  OAI221_X1 U5115 ( .B1(U3149), .B2(keyinput113), .C1(n4571), .C2(keyinput66), 
        .A(n4570), .ZN(n4659) );
  INV_X1 U5116 ( .A(keyinput90), .ZN(n4577) );
  AOI22_X1 U5117 ( .A1(n4574), .A2(keyinput5), .B1(keyinput47), .B2(n4573), 
        .ZN(n4572) );
  OAI221_X1 U5118 ( .B1(n4574), .B2(keyinput5), .C1(n4573), .C2(keyinput47), 
        .A(n4572), .ZN(n4575) );
  AOI221_X1 U5119 ( .B1(REG3_REG_25__SCAN_IN), .B2(n4577), .C1(n4576), .C2(
        keyinput90), .A(n4575), .ZN(n4595) );
  INV_X1 U5120 ( .A(keyinput56), .ZN(n4580) );
  INV_X1 U5121 ( .A(keyinput10), .ZN(n4579) );
  AOI22_X1 U5122 ( .A1(n4580), .A2(DATAO_REG_13__SCAN_IN), .B1(
        DATAO_REG_9__SCAN_IN), .B2(n4579), .ZN(n4578) );
  OAI221_X1 U5123 ( .B1(n4580), .B2(DATAO_REG_13__SCAN_IN), .C1(n4579), .C2(
        DATAO_REG_9__SCAN_IN), .A(n4578), .ZN(n4593) );
  INV_X1 U5124 ( .A(keyinput21), .ZN(n4583) );
  INV_X1 U5125 ( .A(keyinput43), .ZN(n4582) );
  AOI22_X1 U5126 ( .A1(n4583), .A2(DATAO_REG_6__SCAN_IN), .B1(
        DATAO_REG_11__SCAN_IN), .B2(n4582), .ZN(n4581) );
  OAI221_X1 U5127 ( .B1(n4583), .B2(DATAO_REG_6__SCAN_IN), .C1(n4582), .C2(
        DATAO_REG_11__SCAN_IN), .A(n4581), .ZN(n4592) );
  AOI22_X1 U5128 ( .A1(n4586), .A2(keyinput28), .B1(n4585), .B2(keyinput96), 
        .ZN(n4584) );
  OAI221_X1 U5129 ( .B1(n4586), .B2(keyinput28), .C1(n4585), .C2(keyinput96), 
        .A(n4584), .ZN(n4591) );
  INV_X1 U5130 ( .A(keyinput63), .ZN(n4589) );
  INV_X1 U5131 ( .A(keyinput92), .ZN(n4588) );
  AOI22_X1 U5132 ( .A1(n4589), .A2(DATAO_REG_15__SCAN_IN), .B1(
        DATAO_REG_14__SCAN_IN), .B2(n4588), .ZN(n4587) );
  OAI221_X1 U5133 ( .B1(n4589), .B2(DATAO_REG_15__SCAN_IN), .C1(n4588), .C2(
        DATAO_REG_14__SCAN_IN), .A(n4587), .ZN(n4590) );
  NOR4_X1 U5134 ( .A1(n4593), .A2(n4592), .A3(n4591), .A4(n4590), .ZN(n4594)
         );
  OAI211_X1 U5135 ( .C1(keyinput30), .C2(n4596), .A(n4595), .B(n4594), .ZN(
        n4658) );
  INV_X1 U5136 ( .A(ADDR_REG_13__SCAN_IN), .ZN(n4599) );
  INV_X1 U5137 ( .A(keyinput9), .ZN(n4598) );
  AOI22_X1 U5138 ( .A1(n4599), .A2(keyinput39), .B1(ADDR_REG_12__SCAN_IN), 
        .B2(n4598), .ZN(n4597) );
  OAI221_X1 U5139 ( .B1(n4599), .B2(keyinput39), .C1(n4598), .C2(
        ADDR_REG_12__SCAN_IN), .A(n4597), .ZN(n4612) );
  AOI22_X1 U5140 ( .A1(n4602), .A2(keyinput89), .B1(keyinput19), .B2(n4601), 
        .ZN(n4600) );
  OAI221_X1 U5141 ( .B1(n4602), .B2(keyinput89), .C1(n4601), .C2(keyinput19), 
        .A(n4600), .ZN(n4611) );
  INV_X1 U5142 ( .A(keyinput44), .ZN(n4604) );
  AOI22_X1 U5143 ( .A1(n4605), .A2(keyinput79), .B1(ADDR_REG_16__SCAN_IN), 
        .B2(n4604), .ZN(n4603) );
  OAI221_X1 U5144 ( .B1(n4605), .B2(keyinput79), .C1(n4604), .C2(
        ADDR_REG_16__SCAN_IN), .A(n4603), .ZN(n4610) );
  XOR2_X1 U5145 ( .A(n4606), .B(keyinput51), .Z(n4608) );
  XNOR2_X1 U5146 ( .A(REG1_REG_2__SCAN_IN), .B(keyinput24), .ZN(n4607) );
  NAND2_X1 U5147 ( .A1(n4608), .A2(n4607), .ZN(n4609) );
  NOR4_X1 U5148 ( .A1(n4612), .A2(n4611), .A3(n4610), .A4(n4609), .ZN(n4656)
         );
  INV_X1 U5149 ( .A(keyinput3), .ZN(n4614) );
  AOI22_X1 U5150 ( .A1(n2222), .A2(keyinput91), .B1(ADDR_REG_5__SCAN_IN), .B2(
        n4614), .ZN(n4613) );
  OAI221_X1 U5151 ( .B1(n2222), .B2(keyinput91), .C1(n4614), .C2(
        ADDR_REG_5__SCAN_IN), .A(n4613), .ZN(n4624) );
  INV_X1 U5152 ( .A(ADDR_REG_2__SCAN_IN), .ZN(n4617) );
  INV_X1 U5153 ( .A(ADDR_REG_4__SCAN_IN), .ZN(n4616) );
  AOI22_X1 U5154 ( .A1(n4617), .A2(keyinput14), .B1(keyinput4), .B2(n4616), 
        .ZN(n4615) );
  OAI221_X1 U5155 ( .B1(n4617), .B2(keyinput14), .C1(n4616), .C2(keyinput4), 
        .A(n4615), .ZN(n4623) );
  INV_X1 U5156 ( .A(keyinput16), .ZN(n4666) );
  AOI22_X1 U5157 ( .A1(n3142), .A2(keyinput31), .B1(ADDR_REG_9__SCAN_IN), .B2(
        n4666), .ZN(n4618) );
  OAI221_X1 U5158 ( .B1(n3142), .B2(keyinput31), .C1(n4666), .C2(
        ADDR_REG_9__SCAN_IN), .A(n4618), .ZN(n4622) );
  INV_X1 U5159 ( .A(keyinput125), .ZN(n4620) );
  AOI22_X1 U5160 ( .A1(n2197), .A2(keyinput95), .B1(ADDR_REG_7__SCAN_IN), .B2(
        n4620), .ZN(n4619) );
  OAI221_X1 U5161 ( .B1(n2197), .B2(keyinput95), .C1(n4620), .C2(
        ADDR_REG_7__SCAN_IN), .A(n4619), .ZN(n4621) );
  NOR4_X1 U5162 ( .A1(n4624), .A2(n4623), .A3(n4622), .A4(n4621), .ZN(n4655)
         );
  AOI22_X1 U5163 ( .A1(n4627), .A2(keyinput34), .B1(n4626), .B2(keyinput48), 
        .ZN(n4625) );
  OAI221_X1 U5164 ( .B1(n4627), .B2(keyinput34), .C1(n4626), .C2(keyinput48), 
        .A(n4625), .ZN(n4639) );
  INV_X1 U5165 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4629) );
  AOI22_X1 U5166 ( .A1(n4630), .A2(keyinput103), .B1(n4629), .B2(keyinput80), 
        .ZN(n4628) );
  OAI221_X1 U5167 ( .B1(n4630), .B2(keyinput103), .C1(n4629), .C2(keyinput80), 
        .A(n4628), .ZN(n4638) );
  INV_X1 U5168 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4632) );
  AOI22_X1 U5169 ( .A1(n4633), .A2(keyinput76), .B1(n4632), .B2(keyinput58), 
        .ZN(n4631) );
  OAI221_X1 U5170 ( .B1(n4633), .B2(keyinput76), .C1(n4632), .C2(keyinput58), 
        .A(n4631), .ZN(n4637) );
  XNOR2_X1 U5171 ( .A(REG3_REG_15__SCAN_IN), .B(keyinput46), .ZN(n4635) );
  XNOR2_X1 U5172 ( .A(IR_REG_28__SCAN_IN), .B(keyinput37), .ZN(n4634) );
  NAND2_X1 U5173 ( .A1(n4635), .A2(n4634), .ZN(n4636) );
  NOR4_X1 U5174 ( .A1(n4639), .A2(n4638), .A3(n4637), .A4(n4636), .ZN(n4654)
         );
  AOI22_X1 U5175 ( .A1(n4642), .A2(keyinput38), .B1(keyinput94), .B2(n4641), 
        .ZN(n4640) );
  OAI221_X1 U5176 ( .B1(n4642), .B2(keyinput38), .C1(n4641), .C2(keyinput94), 
        .A(n4640), .ZN(n4652) );
  INV_X1 U5177 ( .A(keyinput35), .ZN(n4644) );
  AOI22_X1 U5178 ( .A1(n4645), .A2(keyinput54), .B1(ADDR_REG_18__SCAN_IN), 
        .B2(n4644), .ZN(n4643) );
  OAI221_X1 U5179 ( .B1(n4645), .B2(keyinput54), .C1(n4644), .C2(
        ADDR_REG_18__SCAN_IN), .A(n4643), .ZN(n4651) );
  XNOR2_X1 U5180 ( .A(REG2_REG_1__SCAN_IN), .B(keyinput100), .ZN(n4649) );
  XNOR2_X1 U5181 ( .A(IR_REG_17__SCAN_IN), .B(keyinput122), .ZN(n4648) );
  XNOR2_X1 U5182 ( .A(REG0_REG_15__SCAN_IN), .B(keyinput18), .ZN(n4647) );
  XNOR2_X1 U5183 ( .A(keyinput112), .B(REG2_REG_7__SCAN_IN), .ZN(n4646) );
  NAND4_X1 U5184 ( .A1(n4649), .A2(n4648), .A3(n4647), .A4(n4646), .ZN(n4650)
         );
  NOR3_X1 U5185 ( .A1(n4652), .A2(n4651), .A3(n4650), .ZN(n4653) );
  NAND4_X1 U5186 ( .A1(n4656), .A2(n4655), .A3(n4654), .A4(n4653), .ZN(n4657)
         );
  NOR4_X1 U5187 ( .A1(n4660), .A2(n4659), .A3(n4658), .A4(n4657), .ZN(n4850)
         );
  NAND2_X1 U5188 ( .A1(keyinput19), .A2(keyinput89), .ZN(n4661) );
  NOR3_X1 U5189 ( .A1(keyinput79), .A2(keyinput24), .A3(n4661), .ZN(n4662) );
  NAND3_X1 U5190 ( .A1(keyinput39), .A2(keyinput44), .A3(n4662), .ZN(n4663) );
  NOR3_X1 U5191 ( .A1(keyinput31), .A2(keyinput9), .A3(n4663), .ZN(n4675) );
  INV_X1 U5192 ( .A(keyinput38), .ZN(n4664) );
  NOR4_X1 U5193 ( .A1(keyinput112), .A2(keyinput94), .A3(keyinput122), .A4(
        n4664), .ZN(n4674) );
  NAND2_X1 U5194 ( .A1(keyinput54), .A2(keyinput35), .ZN(n4665) );
  NOR3_X1 U5195 ( .A1(keyinput51), .A2(keyinput100), .A3(n4665), .ZN(n4673) );
  NAND4_X1 U5196 ( .A1(keyinput95), .A2(keyinput3), .A3(keyinput125), .A4(
        n4666), .ZN(n4671) );
  NAND4_X1 U5197 ( .A1(keyinput72), .A2(keyinput14), .A3(keyinput4), .A4(
        keyinput91), .ZN(n4670) );
  NOR3_X1 U5198 ( .A1(keyinput37), .A2(keyinput103), .A3(keyinput58), .ZN(
        n4667) );
  NAND2_X1 U5199 ( .A1(keyinput76), .A2(n4667), .ZN(n4669) );
  NAND4_X1 U5200 ( .A1(keyinput18), .A2(keyinput46), .A3(keyinput80), .A4(
        keyinput34), .ZN(n4668) );
  NOR4_X1 U5201 ( .A1(n4671), .A2(n4670), .A3(n4669), .A4(n4668), .ZN(n4672)
         );
  NAND4_X1 U5202 ( .A1(n4675), .A2(n4674), .A3(n4673), .A4(n4672), .ZN(n4721)
         );
  NAND2_X1 U5203 ( .A1(keyinput99), .A2(keyinput109), .ZN(n4676) );
  NOR3_X1 U5204 ( .A1(keyinput23), .A2(keyinput59), .A3(n4676), .ZN(n4719) );
  NOR4_X1 U5205 ( .A1(keyinput120), .A2(keyinput27), .A3(keyinput61), .A4(
        keyinput70), .ZN(n4718) );
  NAND2_X1 U5206 ( .A1(keyinput11), .A2(keyinput117), .ZN(n4677) );
  NOR3_X1 U5207 ( .A1(keyinput48), .A2(keyinput7), .A3(n4677), .ZN(n4678) );
  NAND3_X1 U5208 ( .A1(keyinput73), .A2(keyinput127), .A3(n4678), .ZN(n4686)
         );
  NAND3_X1 U5209 ( .A1(keyinput111), .A2(keyinput98), .A3(keyinput65), .ZN(
        n4679) );
  NOR2_X1 U5210 ( .A1(keyinput41), .A2(n4679), .ZN(n4684) );
  NOR4_X1 U5211 ( .A1(keyinput107), .A2(keyinput25), .A3(keyinput64), .A4(
        keyinput124), .ZN(n4683) );
  NOR4_X1 U5212 ( .A1(keyinput69), .A2(keyinput13), .A3(keyinput71), .A4(
        keyinput75), .ZN(n4682) );
  NAND2_X1 U5213 ( .A1(keyinput42), .A2(keyinput12), .ZN(n4680) );
  NOR3_X1 U5214 ( .A1(keyinput85), .A2(keyinput62), .A3(n4680), .ZN(n4681) );
  NAND4_X1 U5215 ( .A1(n4684), .A2(n4683), .A3(n4682), .A4(n4681), .ZN(n4685)
         );
  NOR4_X1 U5216 ( .A1(keyinput74), .A2(keyinput78), .A3(n4686), .A4(n4685), 
        .ZN(n4717) );
  NAND3_X1 U5217 ( .A1(keyinput86), .A2(keyinput66), .A3(keyinput47), .ZN(
        n4687) );
  NOR2_X1 U5218 ( .A1(keyinput113), .A2(n4687), .ZN(n4688) );
  NAND4_X1 U5219 ( .A1(keyinput55), .A2(keyinput90), .A3(keyinput5), .A4(n4688), .ZN(n4715) );
  INV_X1 U5220 ( .A(keyinput6), .ZN(n4689) );
  NOR4_X1 U5221 ( .A1(keyinput82), .A2(keyinput15), .A3(keyinput20), .A4(n4689), .ZN(n4699) );
  NAND2_X1 U5222 ( .A1(keyinput40), .A2(keyinput114), .ZN(n4690) );
  NOR3_X1 U5223 ( .A1(keyinput81), .A2(keyinput2), .A3(n4690), .ZN(n4698) );
  NAND4_X1 U5224 ( .A1(keyinput43), .A2(keyinput56), .A3(keyinput10), .A4(
        keyinput63), .ZN(n4696) );
  NOR2_X1 U5225 ( .A1(keyinput33), .A2(keyinput28), .ZN(n4691) );
  NAND3_X1 U5226 ( .A1(keyinput21), .A2(keyinput92), .A3(n4691), .ZN(n4695) );
  NAND4_X1 U5227 ( .A1(keyinput83), .A2(keyinput17), .A3(keyinput1), .A4(
        keyinput123), .ZN(n4694) );
  NOR3_X1 U5228 ( .A1(keyinput96), .A2(keyinput106), .A3(keyinput93), .ZN(
        n4692) );
  NAND2_X1 U5229 ( .A1(keyinput102), .A2(n4692), .ZN(n4693) );
  NOR4_X1 U5230 ( .A1(n4696), .A2(n4695), .A3(n4694), .A4(n4693), .ZN(n4697)
         );
  NAND3_X1 U5231 ( .A1(n4699), .A2(n4698), .A3(n4697), .ZN(n4714) );
  INV_X1 U5232 ( .A(keyinput101), .ZN(n4700) );
  NOR4_X1 U5233 ( .A1(keyinput68), .A2(keyinput52), .A3(keyinput105), .A4(
        n4700), .ZN(n4706) );
  AND4_X1 U5234 ( .A1(keyinput108), .A2(keyinput84), .A3(keyinput8), .A4(
        keyinput121), .ZN(n4705) );
  INV_X1 U5235 ( .A(keyinput110), .ZN(n4701) );
  NOR4_X1 U5236 ( .A1(keyinput118), .A2(keyinput67), .A3(keyinput119), .A4(
        n4701), .ZN(n4704) );
  NAND2_X1 U5237 ( .A1(keyinput87), .A2(keyinput53), .ZN(n4702) );
  NOR3_X1 U5238 ( .A1(keyinput49), .A2(keyinput29), .A3(n4702), .ZN(n4703) );
  NAND4_X1 U5239 ( .A1(n4706), .A2(n4705), .A3(n4704), .A4(n4703), .ZN(n4713)
         );
  NAND2_X1 U5240 ( .A1(keyinput57), .A2(keyinput50), .ZN(n4707) );
  NOR3_X1 U5241 ( .A1(keyinput32), .A2(keyinput26), .A3(n4707), .ZN(n4711) );
  NOR4_X1 U5242 ( .A1(keyinput77), .A2(keyinput22), .A3(keyinput126), .A4(
        keyinput104), .ZN(n4710) );
  AND4_X1 U5243 ( .A1(keyinput97), .A2(keyinput0), .A3(keyinput115), .A4(
        keyinput36), .ZN(n4709) );
  NOR4_X1 U5244 ( .A1(keyinput60), .A2(keyinput45), .A3(keyinput88), .A4(
        keyinput116), .ZN(n4708) );
  NAND4_X1 U5245 ( .A1(n4711), .A2(n4710), .A3(n4709), .A4(n4708), .ZN(n4712)
         );
  NOR4_X1 U5246 ( .A1(n4715), .A2(n4714), .A3(n4713), .A4(n4712), .ZN(n4716)
         );
  NAND4_X1 U5247 ( .A1(n4719), .A2(n4718), .A3(n4717), .A4(n4716), .ZN(n4720)
         );
  OAI21_X1 U5248 ( .B1(n4721), .B2(n4720), .A(DATAI_20_), .ZN(n4848) );
  AOI22_X1 U5249 ( .A1(n4724), .A2(keyinput117), .B1(n4723), .B2(keyinput74), 
        .ZN(n4722) );
  OAI221_X1 U5250 ( .B1(n4724), .B2(keyinput117), .C1(n4723), .C2(keyinput74), 
        .A(n4722), .ZN(n4734) );
  XNOR2_X1 U5251 ( .A(IR_REG_1__SCAN_IN), .B(keyinput11), .ZN(n4728) );
  XNOR2_X1 U5252 ( .A(DATAI_1_), .B(keyinput78), .ZN(n4727) );
  XNOR2_X1 U5253 ( .A(IR_REG_5__SCAN_IN), .B(keyinput127), .ZN(n4726) );
  XNOR2_X1 U5254 ( .A(IR_REG_4__SCAN_IN), .B(keyinput73), .ZN(n4725) );
  NAND4_X1 U5255 ( .A1(n4728), .A2(n4727), .A3(n4726), .A4(n4725), .ZN(n4733)
         );
  XNOR2_X1 U5256 ( .A(keyinput7), .B(n4729), .ZN(n4732) );
  INV_X1 U5257 ( .A(DATAI_6_), .ZN(n4730) );
  XNOR2_X1 U5258 ( .A(keyinput120), .B(n4730), .ZN(n4731) );
  NOR4_X1 U5259 ( .A1(n4734), .A2(n4733), .A3(n4732), .A4(n4731), .ZN(n4783)
         );
  AOI22_X1 U5260 ( .A1(n4737), .A2(keyinput70), .B1(keyinput99), .B2(n4736), 
        .ZN(n4735) );
  OAI221_X1 U5261 ( .B1(n4737), .B2(keyinput70), .C1(n4736), .C2(keyinput99), 
        .A(n4735), .ZN(n4746) );
  XNOR2_X1 U5262 ( .A(n4738), .B(keyinput59), .ZN(n4745) );
  XNOR2_X1 U5263 ( .A(keyinput61), .B(n3071), .ZN(n4744) );
  XNOR2_X1 U5264 ( .A(IR_REG_8__SCAN_IN), .B(keyinput27), .ZN(n4742) );
  XNOR2_X1 U5265 ( .A(DATAI_10_), .B(keyinput23), .ZN(n4741) );
  XNOR2_X1 U5266 ( .A(DATAI_14_), .B(keyinput107), .ZN(n4740) );
  XNOR2_X1 U5267 ( .A(IR_REG_10__SCAN_IN), .B(keyinput109), .ZN(n4739) );
  NAND4_X1 U5268 ( .A1(n4742), .A2(n4741), .A3(n4740), .A4(n4739), .ZN(n4743)
         );
  NOR4_X1 U5269 ( .A1(n4746), .A2(n4745), .A3(n4744), .A4(n4743), .ZN(n4782)
         );
  AOI22_X1 U5270 ( .A1(n4749), .A2(keyinput124), .B1(keyinput12), .B2(n4748), 
        .ZN(n4747) );
  OAI221_X1 U5271 ( .B1(n4749), .B2(keyinput124), .C1(n4748), .C2(keyinput12), 
        .A(n4747), .ZN(n4754) );
  XNOR2_X1 U5272 ( .A(n4750), .B(keyinput25), .ZN(n4753) );
  XNOR2_X1 U5273 ( .A(n4751), .B(keyinput65), .ZN(n4752) );
  OR3_X1 U5274 ( .A1(n4754), .A2(n4753), .A3(n4752), .ZN(n4763) );
  AOI22_X1 U5275 ( .A1(n4757), .A2(keyinput111), .B1(keyinput64), .B2(n4756), 
        .ZN(n4755) );
  OAI221_X1 U5276 ( .B1(n4757), .B2(keyinput111), .C1(n4756), .C2(keyinput64), 
        .A(n4755), .ZN(n4762) );
  AOI22_X1 U5277 ( .A1(n4760), .A2(keyinput41), .B1(keyinput98), .B2(n4759), 
        .ZN(n4758) );
  OAI221_X1 U5278 ( .B1(n4760), .B2(keyinput41), .C1(n4759), .C2(keyinput98), 
        .A(n4758), .ZN(n4761) );
  NOR3_X1 U5279 ( .A1(n4763), .A2(n4762), .A3(n4761), .ZN(n4781) );
  AOI22_X1 U5280 ( .A1(n4766), .A2(keyinput85), .B1(keyinput69), .B2(n4765), 
        .ZN(n4764) );
  OAI221_X1 U5281 ( .B1(n4766), .B2(keyinput85), .C1(n4765), .C2(keyinput69), 
        .A(n4764), .ZN(n4779) );
  AOI22_X1 U5282 ( .A1(n4769), .A2(keyinput13), .B1(keyinput42), .B2(n4768), 
        .ZN(n4767) );
  OAI221_X1 U5283 ( .B1(n4769), .B2(keyinput13), .C1(n4768), .C2(keyinput42), 
        .A(n4767), .ZN(n4778) );
  AOI22_X1 U5284 ( .A1(n4772), .A2(keyinput62), .B1(keyinput71), .B2(n4771), 
        .ZN(n4770) );
  OAI221_X1 U5285 ( .B1(n4772), .B2(keyinput62), .C1(n4771), .C2(keyinput71), 
        .A(n4770), .ZN(n4777) );
  AOI22_X1 U5286 ( .A1(n4775), .A2(keyinput75), .B1(keyinput77), .B2(n4774), 
        .ZN(n4773) );
  OAI221_X1 U5287 ( .B1(n4775), .B2(keyinput75), .C1(n4774), .C2(keyinput77), 
        .A(n4773), .ZN(n4776) );
  NOR4_X1 U5288 ( .A1(n4779), .A2(n4778), .A3(n4777), .A4(n4776), .ZN(n4780)
         );
  NAND4_X1 U5289 ( .A1(n4783), .A2(n4782), .A3(n4781), .A4(n4780), .ZN(n4847)
         );
  INV_X1 U5290 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4785) );
  AOI22_X1 U5291 ( .A1(n4786), .A2(keyinput22), .B1(n4785), .B2(keyinput32), 
        .ZN(n4784) );
  OAI221_X1 U5292 ( .B1(n4786), .B2(keyinput22), .C1(n4785), .C2(keyinput32), 
        .A(n4784), .ZN(n4798) );
  AOI22_X1 U5293 ( .A1(n3621), .A2(keyinput50), .B1(keyinput26), .B2(n4788), 
        .ZN(n4787) );
  OAI221_X1 U5294 ( .B1(n3621), .B2(keyinput50), .C1(n4788), .C2(keyinput26), 
        .A(n4787), .ZN(n4797) );
  AOI22_X1 U5295 ( .A1(n4791), .A2(keyinput57), .B1(keyinput126), .B2(n4790), 
        .ZN(n4789) );
  OAI221_X1 U5296 ( .B1(n4791), .B2(keyinput57), .C1(n4790), .C2(keyinput126), 
        .A(n4789), .ZN(n4796) );
  INV_X1 U5297 ( .A(keyinput104), .ZN(n4794) );
  INV_X1 U5298 ( .A(keyinput60), .ZN(n4793) );
  AOI22_X1 U5299 ( .A1(n4794), .A2(DATAO_REG_25__SCAN_IN), .B1(
        DATAO_REG_26__SCAN_IN), .B2(n4793), .ZN(n4792) );
  OAI221_X1 U5300 ( .B1(n4794), .B2(DATAO_REG_25__SCAN_IN), .C1(n4793), .C2(
        DATAO_REG_26__SCAN_IN), .A(n4792), .ZN(n4795) );
  NOR4_X1 U5301 ( .A1(n4798), .A2(n4797), .A3(n4796), .A4(n4795), .ZN(n4845)
         );
  AOI22_X1 U5302 ( .A1(n4801), .A2(keyinput45), .B1(n4800), .B2(keyinput97), 
        .ZN(n4799) );
  OAI221_X1 U5303 ( .B1(n4801), .B2(keyinput45), .C1(n4800), .C2(keyinput97), 
        .A(n4799), .ZN(n4813) );
  INV_X1 U5304 ( .A(keyinput115), .ZN(n4803) );
  AOI22_X1 U5305 ( .A1(n4804), .A2(keyinput0), .B1(DATAO_REG_29__SCAN_IN), 
        .B2(n4803), .ZN(n4802) );
  OAI221_X1 U5306 ( .B1(n4804), .B2(keyinput0), .C1(n4803), .C2(
        DATAO_REG_29__SCAN_IN), .A(n4802), .ZN(n4812) );
  INV_X1 U5307 ( .A(keyinput36), .ZN(n4806) );
  AOI22_X1 U5308 ( .A1(n2423), .A2(keyinput88), .B1(DATAO_REG_30__SCAN_IN), 
        .B2(n4806), .ZN(n4805) );
  OAI221_X1 U5309 ( .B1(n2423), .B2(keyinput88), .C1(n4806), .C2(
        DATAO_REG_30__SCAN_IN), .A(n4805), .ZN(n4811) );
  AOI22_X1 U5310 ( .A1(n4809), .A2(keyinput116), .B1(n4808), .B2(keyinput108), 
        .ZN(n4807) );
  OAI221_X1 U5311 ( .B1(n4809), .B2(keyinput116), .C1(n4808), .C2(keyinput108), 
        .A(n4807), .ZN(n4810) );
  NOR4_X1 U5312 ( .A1(n4813), .A2(n4812), .A3(n4811), .A4(n4810), .ZN(n4844)
         );
  INV_X1 U5313 ( .A(keyinput52), .ZN(n4816) );
  INV_X1 U5314 ( .A(keyinput8), .ZN(n4815) );
  AOI22_X1 U5315 ( .A1(n4816), .A2(DATAO_REG_1__SCAN_IN), .B1(
        DATAO_REG_22__SCAN_IN), .B2(n4815), .ZN(n4814) );
  OAI221_X1 U5316 ( .B1(n4816), .B2(DATAO_REG_1__SCAN_IN), .C1(n4815), .C2(
        DATAO_REG_22__SCAN_IN), .A(n4814), .ZN(n4827) );
  INV_X1 U5317 ( .A(REG0_REG_18__SCAN_IN), .ZN(n4819) );
  AOI22_X1 U5318 ( .A1(n4819), .A2(keyinput84), .B1(n4818), .B2(keyinput68), 
        .ZN(n4817) );
  OAI221_X1 U5319 ( .B1(n4819), .B2(keyinput84), .C1(n4818), .C2(keyinput68), 
        .A(n4817), .ZN(n4826) );
  INV_X1 U5320 ( .A(keyinput121), .ZN(n4820) );
  XOR2_X1 U5321 ( .A(DATAO_REG_10__SCAN_IN), .B(n4820), .Z(n4824) );
  XNOR2_X1 U5322 ( .A(IR_REG_25__SCAN_IN), .B(keyinput105), .ZN(n4823) );
  XNOR2_X1 U5323 ( .A(IR_REG_29__SCAN_IN), .B(keyinput101), .ZN(n4822) );
  XNOR2_X1 U5324 ( .A(IR_REG_26__SCAN_IN), .B(keyinput49), .ZN(n4821) );
  NAND4_X1 U5325 ( .A1(n4824), .A2(n4823), .A3(n4822), .A4(n4821), .ZN(n4825)
         );
  NOR3_X1 U5326 ( .A1(n4827), .A2(n4826), .A3(n4825), .ZN(n4843) );
  AOI22_X1 U5327 ( .A1(n2719), .A2(keyinput87), .B1(keyinput110), .B2(n4829), 
        .ZN(n4828) );
  OAI221_X1 U5328 ( .B1(n2719), .B2(keyinput87), .C1(n4829), .C2(keyinput110), 
        .A(n4828), .ZN(n4841) );
  INV_X1 U5329 ( .A(DATAI_13_), .ZN(n4832) );
  AOI22_X1 U5330 ( .A1(n4832), .A2(keyinput67), .B1(n4831), .B2(keyinput118), 
        .ZN(n4830) );
  OAI221_X1 U5331 ( .B1(n4832), .B2(keyinput67), .C1(n4831), .C2(keyinput118), 
        .A(n4830), .ZN(n4840) );
  INV_X1 U5332 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4834) );
  AOI22_X1 U5333 ( .A1(n4835), .A2(keyinput53), .B1(keyinput29), .B2(n4834), 
        .ZN(n4833) );
  OAI221_X1 U5334 ( .B1(n4835), .B2(keyinput53), .C1(n4834), .C2(keyinput29), 
        .A(n4833), .ZN(n4839) );
  XOR2_X1 U5335 ( .A(n2346), .B(keyinput119), .Z(n4837) );
  XNOR2_X1 U5336 ( .A(REG2_REG_0__SCAN_IN), .B(keyinput55), .ZN(n4836) );
  NAND2_X1 U5337 ( .A1(n4837), .A2(n4836), .ZN(n4838) );
  NOR4_X1 U5338 ( .A1(n4841), .A2(n4840), .A3(n4839), .A4(n4838), .ZN(n4842)
         );
  NAND4_X1 U5339 ( .A1(n4845), .A2(n4844), .A3(n4843), .A4(n4842), .ZN(n4846)
         );
  AOI211_X1 U5340 ( .C1(keyinput30), .C2(n4848), .A(n4847), .B(n4846), .ZN(
        n4849) );
  NAND4_X1 U5341 ( .A1(n4852), .A2(n4851), .A3(n4850), .A4(n4849), .ZN(n4853)
         );
  XOR2_X1 U5342 ( .A(n4854), .B(n4853), .Z(U3568) );
  NOR2_X1 U2415 ( .A1(n2162), .A2(n2328), .ZN(n2327) );
  NAND2_X1 U2416 ( .A1(n2338), .A2(n2335), .ZN(n2363) );
  CLKBUF_X1 U2417 ( .A(n2608), .Z(n3400) );
  OR2_X1 U2418 ( .A1(n4192), .A2(n4328), .ZN(n4153) );
  NOR2_X1 U2432 ( .A1(n3062), .A2(n3098), .ZN(n3111) );
  AND2_X1 U2631 ( .A1(n2354), .A2(n2330), .ZN(n2385) );
  MUX2_X1 U2633 ( .A(n3890), .B(n2541), .S(n3734), .Z(n2846) );
  OR2_X1 U2813 ( .A1(n3486), .A2(n3485), .ZN(n4192) );
  AND2_X1 U2834 ( .A1(n2528), .A2(n2527), .ZN(n2841) );
  OR3_X1 U2836 ( .A1(n4153), .A2(n4152), .A3(n4122), .ZN(n4857) );
  NOR2_X1 U2839 ( .A1(n2767), .A2(n2761), .ZN(n4858) );
  NOR3_X1 U2840 ( .A1(n4153), .A2(n4152), .A3(n4122), .ZN(n4859) );
  NOR3_X1 U2852 ( .A1(n4072), .A2(n4050), .A3(n2190), .ZN(n4860) );
  NOR3_X1 U2853 ( .A1(n3221), .A2(n3243), .A3(n3256), .ZN(n4861) );
  CLKBUF_X1 U2854 ( .A(n3734), .Z(n4862) );
  NOR2_X1 U2855 ( .A1(n2767), .A2(n2761), .ZN(n2798) );
  AND2_X1 U2902 ( .A1(n2846), .A2(n2841), .ZN(n2633) );
  NOR3_X1 U2969 ( .A1(n4153), .A2(n4152), .A3(n4122), .ZN(n4127) );
  NOR3_X1 U3428 ( .A1(n4072), .A2(n4050), .A3(n2190), .ZN(n4030) );
  OR2_X1 U4247 ( .A1(n4243), .A2(n4066), .ZN(n4072) );
  NOR3_X1 U4763 ( .A1(n3221), .A2(n3243), .A3(n3256), .ZN(n3343) );
  NAND2_X1 U5343 ( .A1(n3139), .A2(n3201), .ZN(n3221) );
  NOR2_X2 U5344 ( .A1(n2921), .A2(n2950), .ZN(n2964) );
  NAND2_X2 U5345 ( .A1(n2191), .A2(n2418), .ZN(n3734) );
  INV_X2 U5346 ( .A(n4465), .ZN(n4350) );
endmodule

