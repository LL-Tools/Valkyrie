

module b14_C_SARLock_k_64_7 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, U3352, U3351, U3350, U3349, U3348, U3347, 
        U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, 
        U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, 
        U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, 
        U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, 
        U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, 
        U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, 
        U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, 
        U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, 
        U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, 
        U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, 
        U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, 
        U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, 
        U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, 
        U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, 
        U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, 
        U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, 
        U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, 
        U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, 
        U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, 
        U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, 
        U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, 
        U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, 
        U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, 
        U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2037, n2038, n2039, n2040, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624;

  NAND4_X1 U2280 ( .A1(n2349), .A2(n2348), .A3(n2347), .A4(n2346), .ZN(n3582)
         );
  OR2_X2 U2281 ( .A1(n2259), .A2(n2812), .ZN(n2356) );
  AND2_X2 U2282 ( .A1(n2305), .A2(n2953), .ZN(n2645) );
  NAND2_X2 U2284 ( .A1(n2288), .A2(n2287), .ZN(n2363) );
  NAND2_X1 U2285 ( .A1(n2744), .A2(IR_REG_31__SCAN_IN), .ZN(n2266) );
  OR2_X1 U2286 ( .A1(n4507), .A2(n4271), .ZN(n4591) );
  AND2_X1 U2287 ( .A1(n2305), .A2(n2953), .ZN(n2037) );
  NAND2_X1 U2288 ( .A1(n4263), .A2(n2812), .ZN(n2354) );
  XNOR2_X2 U2289 ( .A(n2252), .B(IR_REG_29__SCAN_IN), .ZN(n2812) );
  NOR2_X2 U2290 ( .A1(n2725), .A2(n2742), .ZN(n2272) );
  XNOR2_X2 U2291 ( .A(n2266), .B(n2265), .ZN(n2725) );
  NAND4_X1 U2292 ( .A1(n2329), .A2(n2328), .A3(n2327), .A4(n2326), .ZN(n4480)
         );
  NAND4_X2 U2293 ( .A1(n2924), .A2(n2923), .A3(n2925), .A4(n2922), .ZN(n2304)
         );
  CLKBUF_X2 U2294 ( .A(n2543), .Z(n2042) );
  CLKBUF_X2 U2295 ( .A(n2543), .Z(n2043) );
  AND2_X1 U2296 ( .A1(n2259), .A2(n2812), .ZN(n2543) );
  OR2_X1 U2297 ( .A1(n2792), .A2(n2787), .ZN(n2807) );
  AND2_X1 U2298 ( .A1(n2133), .A2(n2132), .ZN(n3403) );
  NAND2_X1 U2299 ( .A1(n2124), .A2(n3361), .ZN(n3338) );
  NOR2_X1 U2300 ( .A1(n4291), .A2(n3345), .ZN(n2150) );
  AND2_X1 U2301 ( .A1(n2570), .A2(n2569), .ZN(n4291) );
  OAI21_X1 U2302 ( .B1(n3092), .B2(n3091), .A(n3448), .ZN(n3182) );
  AND2_X2 U2303 ( .A1(n2950), .A2(n4515), .ZN(n4296) );
  NAND4_X1 U2304 ( .A1(n2310), .A2(n2309), .A3(n2308), .A4(n2307), .ZN(n3584)
         );
  NAND4_X1 U2305 ( .A1(n2360), .A2(n2359), .A3(n2358), .A4(n2357), .ZN(n3581)
         );
  CLKBUF_X2 U2306 ( .A(n2354), .Z(n2039) );
  CLKBUF_X2 U2307 ( .A(n2354), .Z(n2040) );
  INV_X2 U2308 ( .A(n2080), .ZN(n2644) );
  NAND2_X1 U2309 ( .A1(n2299), .A2(n2300), .ZN(n4492) );
  INV_X4 U2310 ( .A(n2080), .ZN(n2038) );
  NAND2_X2 U2311 ( .A1(n2937), .A2(n2936), .ZN(n4502) );
  XNOR2_X1 U2312 ( .A(n2255), .B(n2808), .ZN(n2259) );
  NAND2_X1 U2313 ( .A1(n2811), .A2(IR_REG_31__SCAN_IN), .ZN(n2255) );
  NAND2_X1 U2314 ( .A1(n2752), .A2(n4270), .ZN(n2953) );
  XNOR2_X1 U2315 ( .A(n2271), .B(IR_REG_26__SCAN_IN), .ZN(n4266) );
  AND2_X1 U2316 ( .A1(n2282), .A2(n2232), .ZN(n2252) );
  XNOR2_X1 U2317 ( .A(n2277), .B(IR_REG_21__SCAN_IN), .ZN(n4270) );
  NOR2_X1 U2318 ( .A1(n2243), .A2(IR_REG_18__SCAN_IN), .ZN(n2177) );
  AND2_X1 U2319 ( .A1(n2050), .A2(n2235), .ZN(n2234) );
  NAND3_X1 U2320 ( .A1(n2157), .A2(n2156), .A3(n2155), .ZN(n4277) );
  NOR2_X1 U2321 ( .A1(n2386), .A2(n2061), .ZN(n2176) );
  AND2_X1 U2322 ( .A1(n2247), .A2(n2193), .ZN(n2192) );
  INV_X1 U2323 ( .A(IR_REG_2__SCAN_IN), .ZN(n2099) );
  INV_X1 U2324 ( .A(IR_REG_3__SCAN_IN), .ZN(n2340) );
  NOR2_X1 U2325 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2098)
         );
  NOR2_X1 U2326 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2240)
         );
  NOR2_X1 U2327 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2241)
         );
  NOR2_X1 U2328 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2242)
         );
  NOR2_X1 U2329 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2452)
         );
  AOI21_X2 U2330 ( .B1(n2957), .B2(n2958), .A(n2394), .ZN(n2965) );
  INV_X8 U2331 ( .A(n2658), .ZN(n2697) );
  AND2_X4 U2332 ( .A1(n2256), .A2(n2259), .ZN(n2353) );
  NAND2_X4 U2333 ( .A1(n2272), .A2(n4266), .ZN(n2305) );
  INV_X1 U2334 ( .A(n3901), .ZN(n2199) );
  NAND2_X1 U2335 ( .A1(n3893), .A2(n3916), .ZN(n2209) );
  AND2_X1 U2336 ( .A1(n2516), .A2(n3251), .ZN(n2538) );
  OR2_X1 U2337 ( .A1(n2282), .A2(n2283), .ZN(n2285) );
  AND4_X1 U2338 ( .A1(n2925), .A2(n2924), .A3(n2923), .A4(n2922), .ZN(n2926)
         );
  NAND2_X1 U2339 ( .A1(n2304), .A2(n2944), .ZN(n3426) );
  INV_X1 U2340 ( .A(n4492), .ZN(n2944) );
  NAND2_X1 U2341 ( .A1(n4345), .A2(n4346), .ZN(n4344) );
  XNOR2_X1 U2342 ( .A(n3140), .B(n4362), .ZN(n4357) );
  XNOR2_X1 U2343 ( .A(n3125), .B(n2166), .ZN(n4379) );
  XNOR2_X1 U2344 ( .A(n3618), .B(n3617), .ZN(n4412) );
  NAND2_X1 U2345 ( .A1(n2273), .A2(IR_REG_31__SCAN_IN), .ZN(n2294) );
  INV_X1 U2346 ( .A(n2386), .ZN(n2175) );
  NOR2_X1 U2347 ( .A1(n2215), .A2(n2058), .ZN(n2214) );
  INV_X1 U2348 ( .A(n2216), .ZN(n2215) );
  AND2_X1 U2349 ( .A1(n2114), .A2(n2113), .ZN(n3994) );
  INV_X1 U2350 ( .A(n3690), .ZN(n2113) );
  NAND2_X1 U2351 ( .A1(n4509), .A2(n2753), .ZN(n4596) );
  OAI21_X1 U2352 ( .B1(n2294), .B2(n2246), .A(n2293), .ZN(n3624) );
  INV_X1 U2353 ( .A(IR_REG_22__SCAN_IN), .ZN(n2193) );
  INV_X1 U2354 ( .A(n2143), .ZN(n2142) );
  OAI21_X1 U2355 ( .B1(n2541), .B2(n2144), .A(n2555), .ZN(n2143) );
  NAND2_X1 U2356 ( .A1(n4326), .A2(n4617), .ZN(n2091) );
  AND2_X1 U2357 ( .A1(n3774), .A2(n3502), .ZN(n3676) );
  NOR2_X1 U2358 ( .A1(n2673), .A2(n4037), .ZN(n2686) );
  OAI21_X1 U2359 ( .B1(n3832), .B2(n3675), .A(n3674), .ZN(n3775) );
  AND2_X1 U2360 ( .A1(n3540), .A2(n3539), .ZN(n3670) );
  AND2_X1 U2361 ( .A1(n3669), .A2(n2105), .ZN(n2103) );
  INV_X1 U2362 ( .A(n2103), .ZN(n2100) );
  NOR2_X1 U2363 ( .A1(n2202), .A2(n2198), .ZN(n2196) );
  AOI21_X1 U2364 ( .B1(n3935), .B2(n2106), .A(n3667), .ZN(n2105) );
  INV_X1 U2365 ( .A(n3666), .ZN(n2106) );
  NOR2_X1 U2366 ( .A1(n3945), .A2(n2107), .ZN(n2104) );
  NAND2_X1 U2367 ( .A1(n3944), .A2(n3935), .ZN(n2107) );
  NAND2_X1 U2368 ( .A1(n3201), .A2(n2118), .ZN(n3531) );
  NOR2_X1 U2369 ( .A1(n2119), .A2(n3422), .ZN(n2118) );
  NAND2_X1 U2370 ( .A1(n3182), .A2(n3442), .ZN(n2117) );
  NOR2_X1 U2371 ( .A1(n3431), .A2(n2977), .ZN(n2225) );
  NAND2_X1 U2372 ( .A1(n2935), .A2(n3523), .ZN(n2974) );
  AND2_X1 U2373 ( .A1(n4269), .A2(n4270), .ZN(n2938) );
  NOR2_X1 U2374 ( .A1(n2183), .A2(n3797), .ZN(n2182) );
  INV_X1 U2375 ( .A(n2184), .ZN(n2183) );
  NAND2_X1 U2376 ( .A1(n2204), .A2(n2209), .ZN(n2201) );
  NOR2_X1 U2377 ( .A1(n2208), .A2(n2203), .ZN(n2202) );
  INV_X1 U2378 ( .A(n2209), .ZN(n2203) );
  AND2_X1 U2379 ( .A1(n2047), .A2(n3220), .ZN(n2174) );
  INV_X1 U2380 ( .A(n4269), .ZN(n2753) );
  NAND2_X1 U2381 ( .A1(n3426), .A2(n3427), .ZN(n4486) );
  INV_X1 U2382 ( .A(IR_REG_17__SCAN_IN), .ZN(n2235) );
  INV_X1 U2383 ( .A(IR_REG_13__SCAN_IN), .ZN(n2244) );
  INV_X1 U2384 ( .A(IR_REG_4__SCAN_IN), .ZN(n2239) );
  NAND2_X1 U2385 ( .A1(n2572), .A2(n2571), .ZN(n2148) );
  NAND2_X1 U2386 ( .A1(n2151), .A2(n2150), .ZN(n2149) );
  NOR2_X1 U2387 ( .A1(n2518), .A2(n2257), .ZN(n2495) );
  AND2_X1 U2388 ( .A1(n2508), .A2(n2507), .ZN(n3249) );
  NAND2_X1 U2389 ( .A1(n2620), .A2(n2619), .ZN(n2621) );
  INV_X1 U2390 ( .A(n2617), .ZN(n2620) );
  INV_X1 U2391 ( .A(n2618), .ZN(n2619) );
  NOR2_X1 U2392 ( .A1(n2651), .A2(n2138), .ZN(n2137) );
  INV_X1 U2393 ( .A(n3374), .ZN(n2138) );
  INV_X1 U2394 ( .A(n3372), .ZN(n2135) );
  AOI22_X1 U2395 ( .A1(n2304), .A2(n2697), .B1(n2038), .B2(n4492), .ZN(n2322)
         );
  INV_X1 U2396 ( .A(n3336), .ZN(n2132) );
  INV_X1 U2397 ( .A(n2812), .ZN(n2256) );
  XNOR2_X1 U2398 ( .A(n3133), .B(n3113), .ZN(n2883) );
  NAND2_X1 U2399 ( .A1(n2887), .A2(n2888), .ZN(n3112) );
  XNOR2_X1 U2400 ( .A(n3112), .B(n3113), .ZN(n3111) );
  INV_X1 U2401 ( .A(n4274), .ZN(n3113) );
  NOR2_X1 U2402 ( .A1(n4303), .A2(n2094), .ZN(n3136) );
  AND2_X1 U2403 ( .A1(n3134), .A2(REG1_REG_5__SCAN_IN), .ZN(n2094) );
  OR2_X1 U2404 ( .A1(n4315), .A2(n4316), .ZN(n2189) );
  NAND2_X1 U2405 ( .A1(n2092), .A2(n2090), .ZN(n3137) );
  NAND2_X1 U2406 ( .A1(n2093), .A2(REG1_REG_7__SCAN_IN), .ZN(n2092) );
  NAND2_X1 U2407 ( .A1(n2091), .A2(n4323), .ZN(n2090) );
  INV_X1 U2408 ( .A(n4326), .ZN(n2093) );
  NAND2_X1 U2409 ( .A1(n4344), .A2(n3139), .ZN(n3140) );
  NAND2_X1 U2410 ( .A1(n4366), .A2(n2072), .ZN(n3125) );
  NAND2_X1 U2411 ( .A1(n4379), .A2(REG2_REG_12__SCAN_IN), .ZN(n4378) );
  OR2_X1 U2412 ( .A1(n2171), .A2(n4273), .ZN(n2170) );
  OAI21_X1 U2413 ( .B1(n4383), .B2(n2089), .A(n2087), .ZN(n3606) );
  INV_X1 U2414 ( .A(n2088), .ZN(n2087) );
  OAI21_X1 U2415 ( .B1(n3144), .B2(n2089), .A(n2085), .ZN(n2088) );
  NAND2_X1 U2416 ( .A1(n2170), .A2(REG2_REG_14__SCAN_IN), .ZN(n2169) );
  NOR2_X1 U2417 ( .A1(n4400), .A2(n2084), .ZN(n3618) );
  NAND2_X1 U2418 ( .A1(n4412), .A2(n2260), .ZN(n4411) );
  NAND2_X1 U2419 ( .A1(n4405), .A2(n2185), .ZN(n3609) );
  NAND2_X1 U2420 ( .A1(n3616), .A2(REG1_REG_15__SCAN_IN), .ZN(n2185) );
  OR2_X1 U2421 ( .A1(n4425), .A2(n4424), .ZN(n2188) );
  INV_X1 U2422 ( .A(n3806), .ZN(n3765) );
  OAI21_X1 U2423 ( .B1(n3831), .B2(n3649), .A(n3648), .ZN(n3792) );
  OAI22_X1 U2424 ( .A1(n3868), .A2(n3645), .B1(n3858), .B2(n3644), .ZN(n3847)
         );
  NAND2_X1 U2425 ( .A1(n2592), .A2(REG3_REG_18__SCAN_IN), .ZN(n2624) );
  AND2_X1 U2426 ( .A1(n3874), .A2(n3872), .ZN(n3901) );
  OAI22_X1 U2427 ( .A1(n3238), .A2(n3237), .B1(n3257), .B2(n3236), .ZN(n3951)
         );
  AOI21_X1 U2428 ( .B1(n2214), .B2(n3102), .A(n2045), .ZN(n2213) );
  OAI21_X1 U2429 ( .B1(n3041), .B2(n3040), .A(n3039), .ZN(n3097) );
  OAI21_X1 U2430 ( .B1(n3017), .B2(n3016), .A(n3445), .ZN(n3043) );
  NOR2_X1 U2431 ( .A1(n4564), .A2(n3432), .ZN(n2983) );
  OAI211_X1 U2432 ( .C1(n2191), .C2(n3426), .A(n2927), .B(n2190), .ZN(n3055)
         );
  NAND2_X1 U2433 ( .A1(n4485), .A2(n2122), .ZN(n2190) );
  OR2_X1 U2434 ( .A1(n2855), .A2(n2854), .ZN(n3075) );
  NAND2_X1 U2435 ( .A1(n2727), .A2(n4266), .ZN(n2814) );
  INV_X1 U2436 ( .A(n2250), .ZN(n2233) );
  AND2_X1 U2437 ( .A1(n2248), .A2(n2147), .ZN(n2146) );
  NAND2_X1 U2438 ( .A1(n2249), .A2(n2248), .ZN(n2270) );
  OR2_X1 U2439 ( .A1(n2039), .A2(n2947), .ZN(n2358) );
  OR2_X1 U2440 ( .A1(n2040), .A2(n3060), .ZN(n2327) );
  NAND2_X1 U2441 ( .A1(n2847), .A2(REG2_REG_3__SCAN_IN), .ZN(n2887) );
  NOR2_X1 U2442 ( .A1(n4305), .A2(n4304), .ZN(n4303) );
  XNOR2_X1 U2443 ( .A(n3136), .B(n2167), .ZN(n4315) );
  NAND2_X1 U2444 ( .A1(n4373), .A2(n4374), .ZN(n4372) );
  XNOR2_X1 U2445 ( .A(n3606), .B(n3128), .ZN(n3146) );
  NAND2_X1 U2446 ( .A1(n4406), .A2(n4407), .ZN(n4405) );
  XNOR2_X1 U2447 ( .A(n3609), .B(n3617), .ZN(n4415) );
  NOR2_X1 U2448 ( .A1(n4415), .A2(REG1_REG_16__SCAN_IN), .ZN(n4416) );
  NAND2_X1 U2449 ( .A1(n4439), .A2(n4440), .ZN(n4437) );
  INV_X1 U2450 ( .A(n3625), .ZN(n2161) );
  NAND2_X1 U2451 ( .A1(n3994), .A2(n2112), .ZN(n4214) );
  NOR2_X1 U2452 ( .A1(n2044), .A2(n2057), .ZN(n2112) );
  OAI21_X1 U2453 ( .B1(n3719), .B2(n3712), .A(n3711), .ZN(n4218) );
  OR2_X1 U2454 ( .A1(n2533), .A2(n2532), .ZN(n2535) );
  XNOR2_X1 U2455 ( .A(n2390), .B(n2722), .ZN(n2391) );
  INV_X1 U2456 ( .A(n4396), .ZN(n2089) );
  NOR2_X1 U2457 ( .A1(n3766), .A2(n3659), .ZN(n2173) );
  INV_X1 U2458 ( .A(n3746), .ZN(n3659) );
  AND2_X1 U2459 ( .A1(n3775), .A2(n3676), .ZN(n3755) );
  NOR2_X1 U2460 ( .A1(n2624), .A2(n2623), .ZN(n2637) );
  OR2_X1 U2461 ( .A1(n3631), .A2(n3630), .ZN(n3637) );
  NAND2_X1 U2462 ( .A1(n4475), .A2(n3427), .ZN(n2933) );
  AND2_X1 U2463 ( .A1(n2753), .A2(n2296), .ZN(n2769) );
  NAND2_X1 U2464 ( .A1(n2173), .A2(n3660), .ZN(n3709) );
  NOR2_X1 U2465 ( .A1(n3835), .A2(n3824), .ZN(n2184) );
  INV_X1 U2466 ( .A(n4493), .ZN(n4508) );
  INV_X1 U2467 ( .A(n2769), .ZN(n4507) );
  OR2_X1 U2468 ( .A1(n2054), .A2(n2597), .ZN(n2746) );
  INV_X1 U2469 ( .A(IR_REG_23__SCAN_IN), .ZN(n2745) );
  NAND2_X1 U2470 ( .A1(n2746), .A2(n2745), .ZN(n2744) );
  INV_X1 U2471 ( .A(n3836), .ZN(n3468) );
  AND2_X1 U2472 ( .A1(n2588), .A2(n2587), .ZN(n3352) );
  NAND2_X1 U2473 ( .A1(n2142), .A2(n2144), .ZN(n2139) );
  NOR2_X1 U2474 ( .A1(n2142), .A2(n2056), .ZN(n2140) );
  NOR2_X1 U2475 ( .A1(n2570), .A2(n2569), .ZN(n4288) );
  NAND2_X1 U2476 ( .A1(n2285), .A2(n2284), .ZN(n2288) );
  INV_X1 U2477 ( .A(n4527), .ZN(n2759) );
  OR2_X1 U2478 ( .A1(n2882), .A2(n2881), .ZN(n3133) );
  NAND2_X1 U2479 ( .A1(n4308), .A2(n2055), .ZN(n3117) );
  NAND2_X1 U2480 ( .A1(n4339), .A2(n3138), .ZN(n4345) );
  INV_X1 U2481 ( .A(REG3_REG_9__SCAN_IN), .ZN(n3156) );
  NAND2_X1 U2482 ( .A1(n4372), .A2(n2082), .ZN(n3143) );
  NOR2_X1 U2483 ( .A1(n3987), .A2(n3989), .ZN(n3986) );
  NAND2_X1 U2484 ( .A1(n3710), .A2(n3693), .ZN(n3987) );
  OAI22_X1 U2485 ( .A1(n3718), .A2(n3661), .B1(n3708), .B2(n3660), .ZN(n3700)
         );
  NAND2_X1 U2486 ( .A1(n3723), .A2(n3679), .ZN(n3702) );
  AND2_X1 U2487 ( .A1(n3680), .A2(n3682), .ZN(n3701) );
  INV_X1 U2488 ( .A(n3738), .ZN(n3708) );
  AOI21_X1 U2489 ( .B1(n3775), .B2(n2071), .A(n3677), .ZN(n3725) );
  NAND2_X1 U2490 ( .A1(n3725), .A2(n3724), .ZN(n3723) );
  INV_X1 U2491 ( .A(n2173), .ZN(n3745) );
  AND2_X1 U2492 ( .A1(n3679), .A2(n3489), .ZN(n3724) );
  NAND2_X1 U2493 ( .A1(n2230), .A2(n2048), .ZN(n2229) );
  NAND2_X1 U2494 ( .A1(n2231), .A2(n3657), .ZN(n2230) );
  AND2_X1 U2495 ( .A1(n2363), .A2(DATAI_24_), .ZN(n3779) );
  INV_X1 U2496 ( .A(n3737), .ZN(n3783) );
  OR3_X1 U2497 ( .A1(n2661), .A2(n3386), .A3(n3314), .ZN(n2673) );
  NAND2_X1 U2498 ( .A1(n2108), .A2(n3671), .ZN(n3832) );
  OR2_X1 U2499 ( .A1(n2104), .A2(n2101), .ZN(n2108) );
  NAND2_X1 U2500 ( .A1(n2103), .A2(n3539), .ZN(n2101) );
  OR2_X1 U2501 ( .A1(n2104), .A2(n2100), .ZN(n3850) );
  NAND2_X1 U2502 ( .A1(n2194), .A2(n2195), .ZN(n3868) );
  NOR2_X1 U2503 ( .A1(n2196), .A2(n2073), .ZN(n2195) );
  AND2_X1 U2504 ( .A1(REG3_REG_17__SCAN_IN), .A2(n2573), .ZN(n2592) );
  NOR2_X1 U2505 ( .A1(n2104), .A2(n2102), .ZN(n3908) );
  INV_X1 U2506 ( .A(n2105), .ZN(n2102) );
  OAI21_X1 U2507 ( .B1(n3945), .B2(n3957), .A(n3666), .ZN(n3923) );
  NOR2_X1 U2508 ( .A1(n2556), .A2(n4278), .ZN(n2557) );
  OR2_X1 U2509 ( .A1(n2545), .A2(n2544), .ZN(n2556) );
  NAND2_X1 U2510 ( .A1(n2120), .A2(n3532), .ZN(n3969) );
  INV_X1 U2511 ( .A(n3954), .ZN(n3973) );
  INV_X1 U2512 ( .A(n3627), .ZN(n3972) );
  NAND2_X1 U2513 ( .A1(n3201), .A2(n3421), .ZN(n3230) );
  AOI21_X1 U2514 ( .B1(n3181), .B2(n2052), .A(n2211), .ZN(n3238) );
  OAI21_X1 U2515 ( .B1(n2213), .B2(n2212), .A(n2060), .ZN(n2211) );
  INV_X1 U2516 ( .A(n3210), .ZN(n2212) );
  NAND2_X1 U2517 ( .A1(n2117), .A2(n2115), .ZN(n3199) );
  NOR2_X1 U2518 ( .A1(n3197), .A2(n2116), .ZN(n2115) );
  INV_X1 U2519 ( .A(n3447), .ZN(n2116) );
  NAND2_X1 U2520 ( .A1(n2219), .A2(n2214), .ZN(n3266) );
  NAND2_X1 U2521 ( .A1(n2117), .A2(n3447), .ZN(n3196) );
  NAND2_X1 U2522 ( .A1(n2218), .A2(n2217), .ZN(n2216) );
  OR2_X1 U2523 ( .A1(n3181), .A2(n3102), .ZN(n2219) );
  NOR2_X1 U2524 ( .A1(n2411), .A2(n2993), .ZN(n2432) );
  AND2_X1 U2525 ( .A1(n2222), .A2(n3005), .ZN(n2221) );
  OAI21_X1 U2526 ( .B1(n2998), .B2(n2997), .A(n3437), .ZN(n3017) );
  INV_X1 U2527 ( .A(n3018), .ZN(n3025) );
  AOI21_X1 U2528 ( .B1(n3002), .B2(n2225), .A(n2059), .ZN(n2224) );
  NAND2_X1 U2529 ( .A1(n3002), .A2(n2227), .ZN(n2226) );
  INV_X1 U2530 ( .A(n2931), .ZN(n2227) );
  INV_X1 U2531 ( .A(n2917), .ZN(n2946) );
  AND2_X1 U2532 ( .A1(n2983), .A2(n2946), .ZN(n3026) );
  NAND2_X1 U2533 ( .A1(n2974), .A2(n3433), .ZN(n2998) );
  OAI21_X1 U2534 ( .B1(n2971), .B2(n2931), .A(n2223), .ZN(n3003) );
  INV_X1 U2535 ( .A(n2225), .ZN(n2223) );
  AND2_X1 U2536 ( .A1(n2934), .A2(n3429), .ZN(n3519) );
  INV_X1 U2537 ( .A(n4478), .ZN(n3930) );
  NAND2_X1 U2538 ( .A1(n2121), .A2(n3426), .ZN(n4475) );
  NOR2_X1 U2539 ( .A1(n3518), .A2(n2122), .ZN(n2121) );
  NAND2_X1 U2540 ( .A1(n4264), .A2(n2938), .ZN(n4482) );
  NAND2_X1 U2541 ( .A1(n2944), .A2(n4508), .ZN(n4495) );
  OR2_X1 U2542 ( .A1(n4296), .A2(n2954), .ZN(n3007) );
  XNOR2_X1 U2543 ( .A(IR_REG_1__SCAN_IN), .B(keyinput41), .ZN(n4138) );
  NOR2_X1 U2544 ( .A1(n3709), .A2(n3704), .ZN(n3710) );
  AND2_X1 U2545 ( .A1(n3859), .A2(n2083), .ZN(n3784) );
  INV_X1 U2546 ( .A(n3809), .ZN(n3797) );
  AND2_X1 U2547 ( .A1(n3859), .A2(n2182), .ZN(n3796) );
  NAND2_X1 U2548 ( .A1(n3859), .A2(n2184), .ZN(n4168) );
  NAND2_X1 U2549 ( .A1(n3859), .A2(n3841), .ZN(n3840) );
  AND2_X1 U2550 ( .A1(n3883), .A2(n3861), .ZN(n3859) );
  INV_X1 U2551 ( .A(n3644), .ZN(n3882) );
  NOR2_X1 U2552 ( .A1(n3960), .A2(n2178), .ZN(n3883) );
  NAND2_X1 U2553 ( .A1(n2181), .A2(n2179), .ZN(n2178) );
  NOR2_X1 U2554 ( .A1(n3642), .A2(n3882), .ZN(n2179) );
  NAND2_X1 U2555 ( .A1(n2200), .A2(n2201), .ZN(n3900) );
  NAND2_X1 U2556 ( .A1(n2207), .A2(n2202), .ZN(n2200) );
  OR2_X1 U2557 ( .A1(n4203), .A2(n4285), .ZN(n3960) );
  OR2_X1 U2558 ( .A1(n3979), .A2(n3978), .ZN(n4203) );
  AND2_X1 U2559 ( .A1(n3178), .A2(n2078), .ZN(n3239) );
  NAND2_X1 U2560 ( .A1(n3178), .A2(n3103), .ZN(n3262) );
  NAND2_X1 U2561 ( .A1(n3178), .A2(n2047), .ZN(n4456) );
  NOR2_X1 U2562 ( .A1(n3049), .A2(n3098), .ZN(n3180) );
  AND2_X1 U2563 ( .A1(n3180), .A2(n2217), .ZN(n3178) );
  OR2_X1 U2564 ( .A1(n3024), .A2(n3038), .ZN(n3049) );
  NAND2_X1 U2565 ( .A1(n4487), .A2(n4596), .ZN(n4594) );
  NAND2_X1 U2566 ( .A1(n2172), .A2(n3066), .ZN(n4564) );
  INV_X1 U2567 ( .A(n4495), .ZN(n2172) );
  NAND2_X1 U2568 ( .A1(n4486), .A2(n4485), .ZN(n4484) );
  AND2_X1 U2569 ( .A1(n3079), .A2(n3078), .ZN(n3085) );
  INV_X1 U2570 ( .A(IR_REG_28__SCAN_IN), .ZN(n2286) );
  OAI21_X1 U2571 ( .B1(n2746), .B2(n2745), .A(n2744), .ZN(n2821) );
  XNOR2_X1 U2572 ( .A(n2274), .B(n2245), .ZN(n2752) );
  AND2_X1 U2573 ( .A1(n2234), .A2(n2487), .ZN(n2598) );
  INV_X1 U2574 ( .A(IR_REG_16__SCAN_IN), .ZN(n2154) );
  NOR2_X1 U2575 ( .A1(n2386), .A2(n2243), .ZN(n2487) );
  OR2_X1 U2576 ( .A1(n2502), .A2(IR_REG_10__SCAN_IN), .ZN(n2503) );
  OR2_X1 U2577 ( .A1(n2470), .A2(IR_REG_9__SCAN_IN), .ZN(n2502) );
  NAND2_X1 U2578 ( .A1(n2410), .A2(n2963), .ZN(n2990) );
  NAND2_X1 U2579 ( .A1(n2126), .A2(n2125), .ZN(n2780) );
  OR2_X1 U2580 ( .A1(n3400), .A2(n2130), .ZN(n2125) );
  NAND2_X1 U2581 ( .A1(n3338), .A2(n2127), .ZN(n2126) );
  NOR2_X1 U2582 ( .A1(n3400), .A2(n2129), .ZN(n2127) );
  NAND2_X1 U2583 ( .A1(n2542), .A2(n2541), .ZN(n3298) );
  INV_X1 U2584 ( .A(n3575), .ZN(n3207) );
  NAND2_X1 U2585 ( .A1(n2344), .A2(n2343), .ZN(n3432) );
  OR2_X1 U2586 ( .A1(n2363), .A2(n2165), .ZN(n2344) );
  NAND2_X1 U2587 ( .A1(n2123), .A2(n2049), .ZN(n2792) );
  NAND2_X1 U2588 ( .A1(n2130), .A2(n2129), .ZN(n2128) );
  OR2_X1 U2589 ( .A1(n2363), .A2(n2298), .ZN(n2299) );
  NAND2_X1 U2590 ( .A1(n2363), .A2(DATAI_1_), .ZN(n2300) );
  INV_X1 U2591 ( .A(n3779), .ZN(n3786) );
  NAND2_X1 U2592 ( .A1(n2312), .A2(n2311), .ZN(n4493) );
  NAND2_X1 U2593 ( .A1(n2363), .A2(DATAI_0_), .ZN(n2311) );
  OR2_X1 U2594 ( .A1(n2363), .A2(n2158), .ZN(n2312) );
  AOI21_X1 U2595 ( .B1(n2137), .B2(n2135), .A(n2075), .ZN(n2134) );
  INV_X1 U2596 ( .A(n2137), .ZN(n2136) );
  OR2_X1 U2597 ( .A1(n2334), .A2(n2333), .ZN(n2335) );
  INV_X1 U2598 ( .A(n3891), .ZN(n3858) );
  INV_X1 U2599 ( .A(n3580), .ZN(n3004) );
  NAND2_X1 U2600 ( .A1(n3338), .A2(n3335), .ZN(n2133) );
  INV_X1 U2601 ( .A(n4295), .ZN(n3408) );
  INV_X1 U2602 ( .A(n3574), .ZN(n4279) );
  INV_X1 U2603 ( .A(n3411), .ZN(n4290) );
  NAND4_X1 U2604 ( .A1(n2643), .A2(n2642), .A3(n2641), .A4(n2640), .ZN(n3855)
         );
  NAND4_X1 U2605 ( .A1(n2501), .A2(n2500), .A3(n2499), .A4(n2498), .ZN(n4445)
         );
  OAI21_X1 U2606 ( .B1(n4277), .B2(n2841), .A(n2160), .ZN(n3596) );
  NAND2_X1 U2607 ( .A1(n4277), .A2(n2841), .ZN(n2160) );
  XNOR2_X1 U2608 ( .A(n2886), .B(n2165), .ZN(n2847) );
  NOR2_X1 U2609 ( .A1(n2839), .A2(n4611), .ZN(n2882) );
  NAND2_X1 U2610 ( .A1(n2883), .A2(REG1_REG_4__SCAN_IN), .ZN(n3132) );
  OAI22_X1 U2611 ( .A1(n3115), .A2(n2355), .B1(n3114), .B2(n3113), .ZN(n4309)
         );
  NAND2_X1 U2612 ( .A1(n4309), .A2(n4310), .ZN(n4308) );
  AND2_X1 U2613 ( .A1(n3132), .A2(n2186), .ZN(n4305) );
  NAND2_X1 U2614 ( .A1(n3133), .A2(n4274), .ZN(n2186) );
  XNOR2_X1 U2615 ( .A(n3117), .B(n2167), .ZN(n4320) );
  INV_X1 U2616 ( .A(n2189), .ZN(n4314) );
  AND2_X1 U2617 ( .A1(n2189), .A2(n2063), .ZN(n4326) );
  XNOR2_X1 U2618 ( .A(n3137), .B(n4343), .ZN(n4340) );
  AND2_X1 U2619 ( .A1(n3588), .A2(n2846), .ZN(n4388) );
  INV_X1 U2620 ( .A(n4540), .ZN(n4377) );
  NAND2_X1 U2621 ( .A1(n4356), .A2(n3141), .ZN(n4373) );
  XNOR2_X1 U2622 ( .A(n3143), .B(n2166), .ZN(n4384) );
  NAND2_X1 U2623 ( .A1(n3126), .A2(n4378), .ZN(n4390) );
  NAND2_X1 U2624 ( .A1(n4383), .A2(n3144), .ZN(n4395) );
  NAND2_X1 U2625 ( .A1(n4395), .A2(n4396), .ZN(n4394) );
  NOR2_X1 U2626 ( .A1(n3615), .A2(n2169), .ZN(n3614) );
  NAND2_X1 U2627 ( .A1(n3607), .A2(n3608), .ZN(n4406) );
  AND2_X1 U2628 ( .A1(n2169), .A2(n2168), .ZN(n4402) );
  NAND2_X1 U2629 ( .A1(n4411), .A2(n3619), .ZN(n4419) );
  NOR2_X1 U2630 ( .A1(n4416), .A2(n3610), .ZN(n4425) );
  INV_X1 U2631 ( .A(n2188), .ZN(n4426) );
  AND2_X1 U2632 ( .A1(n2188), .A2(n2187), .ZN(n4439) );
  NAND2_X1 U2633 ( .A1(n4429), .A2(n4191), .ZN(n2187) );
  AND2_X1 U2634 ( .A1(n3588), .A2(n3585), .ZN(n4438) );
  OR2_X1 U2635 ( .A1(n2714), .A2(n2701), .ZN(n3748) );
  AOI21_X1 U2636 ( .B1(n3655), .B2(n2067), .A(n2236), .ZN(n3754) );
  NAND2_X1 U2637 ( .A1(n3655), .A2(n3654), .ZN(n3773) );
  NAND2_X1 U2638 ( .A1(n2207), .A2(n2206), .ZN(n2205) );
  NAND2_X1 U2639 ( .A1(n2210), .A2(n2213), .ZN(n4449) );
  NAND2_X1 U2640 ( .A1(n3181), .A2(n2214), .ZN(n2210) );
  INV_X1 U2641 ( .A(n4515), .ZN(n4491) );
  OR2_X1 U2642 ( .A1(n2855), .A2(n2771), .ZN(n4515) );
  INV_X1 U2643 ( .A(n3007), .ZN(n4501) );
  AND2_X2 U2644 ( .A1(n3085), .A2(n3080), .ZN(n4624) );
  AND2_X2 U2645 ( .A1(n3085), .A2(n3084), .ZN(n4605) );
  INV_X1 U2646 ( .A(IR_REG_30__SCAN_IN), .ZN(n2808) );
  INV_X1 U2647 ( .A(n2259), .ZN(n4263) );
  NOR2_X1 U2648 ( .A1(n2251), .A2(n2233), .ZN(n2232) );
  AND2_X1 U2649 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_28__SCAN_IN), .ZN(n2251)
         );
  NAND2_X1 U2650 ( .A1(n2270), .A2(IR_REG_31__SCAN_IN), .ZN(n2271) );
  NAND2_X1 U2651 ( .A1(n2821), .A2(STATE_REG_SCAN_IN), .ZN(n4527) );
  XNOR2_X1 U2652 ( .A(n2292), .B(IR_REG_22__SCAN_IN), .ZN(n4269) );
  NAND2_X1 U2653 ( .A1(n2291), .A2(IR_REG_31__SCAN_IN), .ZN(n2292) );
  INV_X1 U2654 ( .A(n2752), .ZN(n4271) );
  XNOR2_X1 U2655 ( .A(n2097), .B(IR_REG_2__SCAN_IN), .ZN(n4276) );
  OAI21_X1 U2656 ( .B1(IR_REG_1__SCAN_IN), .B2(IR_REG_0__SCAN_IN), .A(
        IR_REG_31__SCAN_IN), .ZN(n2097) );
  NAND3_X1 U2657 ( .A1(n2159), .A2(IR_REG_0__SCAN_IN), .A3(IR_REG_31__SCAN_IN), 
        .ZN(n2157) );
  NAND2_X1 U2658 ( .A1(n2158), .A2(IR_REG_1__SCAN_IN), .ZN(n2156) );
  NAND2_X1 U2659 ( .A1(n2597), .A2(IR_REG_1__SCAN_IN), .ZN(n2155) );
  OAI21_X1 U2660 ( .B1(n2096), .B2(n4313), .A(n2095), .ZN(U3259) );
  XNOR2_X1 U2661 ( .A(n3613), .B(n3612), .ZN(n2096) );
  AND2_X1 U2662 ( .A1(n2162), .A2(n2161), .ZN(n2095) );
  MUX2_X1 U2663 ( .A(n3997), .B(n4215), .S(n4624), .Z(n3998) );
  INV_X1 U2664 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2110) );
  MUX2_X1 U2665 ( .A(n4216), .B(n4215), .S(n4605), .Z(n4217) );
  INV_X1 U2666 ( .A(IR_REG_31__SCAN_IN), .ZN(n2597) );
  INV_X1 U2667 ( .A(n3578), .ZN(n2218) );
  NAND2_X1 U2668 ( .A1(n2201), .A2(n2199), .ZN(n2198) );
  AND2_X1 U2669 ( .A1(n3992), .A2(n4594), .ZN(n2044) );
  NAND2_X1 U2670 ( .A1(n2076), .A2(n3643), .ZN(n2204) );
  NAND2_X1 U2671 ( .A1(n2064), .A2(n3265), .ZN(n2045) );
  AND2_X1 U2672 ( .A1(n2426), .A2(n2963), .ZN(n2046) );
  INV_X1 U2673 ( .A(n4296), .ZN(n4511) );
  AND2_X1 U2674 ( .A1(n3103), .A2(n3263), .ZN(n2047) );
  NAND2_X1 U2675 ( .A1(n3737), .A2(n3656), .ZN(n2048) );
  AND3_X1 U2676 ( .A1(n2131), .A2(n2779), .A3(n2128), .ZN(n2049) );
  INV_X1 U2677 ( .A(n3400), .ZN(n2131) );
  AND4_X1 U2678 ( .A1(n2244), .A2(n2154), .A3(n2153), .A4(n2152), .ZN(n2050)
         );
  NAND2_X1 U2679 ( .A1(n2145), .A2(IR_REG_31__SCAN_IN), .ZN(n2282) );
  NAND2_X1 U2680 ( .A1(n3580), .A2(n3018), .ZN(n2051) );
  NAND4_X1 U2681 ( .A1(n2098), .A2(n2239), .A3(n2340), .A4(n2099), .ZN(n2386)
         );
  NAND2_X1 U2682 ( .A1(n2926), .A2(n4492), .ZN(n3427) );
  INV_X1 U2683 ( .A(n3427), .ZN(n2122) );
  AND2_X1 U2684 ( .A1(n2214), .A2(n3210), .ZN(n2052) );
  AND4_X1 U2685 ( .A1(n2147), .A2(n2286), .A3(n2283), .A4(n2253), .ZN(n2053)
         );
  AND2_X1 U2686 ( .A1(n2275), .A2(n2192), .ZN(n2054) );
  AND2_X1 U2687 ( .A1(n3537), .A2(n3536), .ZN(n3935) );
  OR2_X1 U2688 ( .A1(n4552), .A2(n3116), .ZN(n2055) );
  AND2_X1 U2689 ( .A1(n2541), .A2(n2144), .ZN(n2056) );
  NOR2_X1 U2690 ( .A1(n3993), .A2(n4591), .ZN(n2057) );
  NOR2_X1 U2691 ( .A1(n3577), .A2(n3206), .ZN(n2058) );
  INV_X1 U2692 ( .A(n2208), .ZN(n2206) );
  OR2_X1 U2693 ( .A1(n3640), .A2(n3935), .ZN(n2208) );
  AND2_X1 U2694 ( .A1(n3581), .A2(n2917), .ZN(n2059) );
  AND3_X1 U2695 ( .A1(n2177), .A2(n2176), .A3(n2234), .ZN(n2275) );
  OR2_X1 U2696 ( .A1(n3209), .A2(n3508), .ZN(n2060) );
  NAND2_X1 U2697 ( .A1(n2246), .A2(n2245), .ZN(n2061) );
  NOR2_X1 U2698 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2062)
         );
  OR2_X1 U2699 ( .A1(n3136), .A2(n2167), .ZN(n2063) );
  NAND2_X1 U2700 ( .A1(n3576), .A2(n3269), .ZN(n2064) );
  AND2_X1 U2701 ( .A1(n2051), .A2(n2224), .ZN(n2065) );
  XNOR2_X1 U2702 ( .A(n2303), .B(n2722), .ZN(n2321) );
  AND2_X1 U2703 ( .A1(n2062), .A2(n2192), .ZN(n2066) );
  INV_X1 U2704 ( .A(n2198), .ZN(n2197) );
  INV_X1 U2705 ( .A(IR_REG_0__SCAN_IN), .ZN(n2158) );
  INV_X1 U2706 ( .A(IR_REG_1__SCAN_IN), .ZN(n2159) );
  INV_X1 U2707 ( .A(n3642), .ZN(n3916) );
  INV_X1 U2708 ( .A(n3135), .ZN(n2167) );
  INV_X1 U2709 ( .A(IR_REG_20__SCAN_IN), .ZN(n2245) );
  INV_X1 U2710 ( .A(n3296), .ZN(n2144) );
  INV_X1 U2711 ( .A(n3183), .ZN(n2217) );
  INV_X1 U2712 ( .A(n4275), .ZN(n2165) );
  AND2_X1 U2713 ( .A1(n3654), .A2(n2238), .ZN(n2067) );
  AND2_X1 U2714 ( .A1(n2487), .A2(n2244), .ZN(n2279) );
  NAND2_X1 U2715 ( .A1(n3370), .A2(n3374), .ZN(n3326) );
  INV_X1 U2716 ( .A(IR_REG_19__SCAN_IN), .ZN(n2246) );
  INV_X1 U2717 ( .A(n3421), .ZN(n2119) );
  INV_X1 U2718 ( .A(n3335), .ZN(n2129) );
  INV_X1 U2719 ( .A(IR_REG_29__SCAN_IN), .ZN(n2253) );
  OR3_X1 U2720 ( .A1(n3960), .A2(n3642), .A3(n3936), .ZN(n2068) );
  AND3_X1 U2721 ( .A1(n2791), .A2(n2793), .A3(n4290), .ZN(n2069) );
  OR3_X1 U2722 ( .A1(n3960), .A2(n2180), .A3(n3642), .ZN(n2070) );
  NAND2_X1 U2723 ( .A1(n2487), .A2(n2050), .ZN(n2582) );
  AND2_X1 U2724 ( .A1(n3678), .A2(n3676), .ZN(n2071) );
  INV_X1 U2725 ( .A(IR_REG_14__SCAN_IN), .ZN(n2153) );
  NAND2_X1 U2726 ( .A1(n3371), .A2(n3372), .ZN(n3370) );
  OR2_X1 U2727 ( .A1(n4377), .A2(n2520), .ZN(n2072) );
  INV_X1 U2728 ( .A(n3235), .ZN(n3236) );
  AND2_X1 U2729 ( .A1(n3881), .A2(n3459), .ZN(n2073) );
  INV_X1 U2730 ( .A(n2151), .ZN(n4286) );
  OR2_X1 U2731 ( .A1(n4288), .A2(n4287), .ZN(n2151) );
  AND2_X1 U2732 ( .A1(n3533), .A2(n3666), .ZN(n3944) );
  AND2_X1 U2733 ( .A1(n2590), .A2(n2589), .ZN(n2074) );
  AND2_X1 U2734 ( .A1(n3328), .A2(n3327), .ZN(n2075) );
  INV_X1 U2735 ( .A(IR_REG_26__SCAN_IN), .ZN(n2147) );
  INV_X1 U2736 ( .A(n2181), .ZN(n2180) );
  NOR2_X1 U2737 ( .A1(n3936), .A2(n3896), .ZN(n2181) );
  NAND2_X1 U2738 ( .A1(n3947), .A2(n3936), .ZN(n2076) );
  AND2_X1 U2739 ( .A1(n2205), .A2(n2076), .ZN(n2077) );
  AND2_X1 U2740 ( .A1(n2174), .A2(n3236), .ZN(n2078) );
  AND2_X1 U2741 ( .A1(n2067), .A2(n2048), .ZN(n2079) );
  AND2_X1 U2742 ( .A1(n3401), .A2(n2132), .ZN(n2130) );
  NAND2_X2 U2743 ( .A1(n2305), .A2(n2278), .ZN(n2080) );
  INV_X1 U2744 ( .A(IR_REG_15__SCAN_IN), .ZN(n2152) );
  INV_X1 U2745 ( .A(n3142), .ZN(n2166) );
  NAND2_X1 U2746 ( .A1(n2991), .A2(n2431), .ZN(n3031) );
  AND2_X1 U2747 ( .A1(n3178), .A2(n2174), .ZN(n2081) );
  NAND2_X1 U2748 ( .A1(n2219), .A2(n2216), .ZN(n3205) );
  AND2_X1 U2749 ( .A1(n2377), .A2(n2376), .ZN(n2957) );
  INV_X1 U2750 ( .A(n2645), .ZN(n2692) );
  INV_X1 U2751 ( .A(n3835), .ZN(n3841) );
  AND2_X1 U2752 ( .A1(n2363), .A2(DATAI_21_), .ZN(n3835) );
  OR2_X1 U2753 ( .A1(n4377), .A2(n4622), .ZN(n2082) );
  AND2_X1 U2754 ( .A1(n2182), .A2(n3786), .ZN(n2083) );
  OAI21_X1 U2755 ( .B1(n2971), .B2(n2226), .A(n2224), .ZN(n3023) );
  AND2_X1 U2756 ( .A1(n2363), .A2(DATAI_27_), .ZN(n3727) );
  AND2_X1 U2757 ( .A1(n3616), .A2(REG2_REG_15__SCAN_IN), .ZN(n2084) );
  OR2_X1 U2758 ( .A1(n4399), .A2(n3145), .ZN(n2085) );
  AND2_X1 U2759 ( .A1(n3620), .A2(REG2_REG_18__SCAN_IN), .ZN(n2086) );
  NAND3_X1 U2760 ( .A1(n2159), .A2(n2099), .A3(n2158), .ZN(n2339) );
  NAND2_X1 U2761 ( .A1(n2111), .A2(n2109), .ZN(U3515) );
  OR2_X1 U2762 ( .A1(n4605), .A2(n2110), .ZN(n2109) );
  NAND2_X1 U2763 ( .A1(n4214), .A2(n4605), .ZN(n2111) );
  NAND2_X1 U2764 ( .A1(n3691), .A2(n4502), .ZN(n2114) );
  NAND2_X1 U2765 ( .A1(n3531), .A2(n3530), .ZN(n2120) );
  NAND3_X1 U2766 ( .A1(n2124), .A2(n3361), .A3(n2130), .ZN(n2123) );
  OR2_X2 U2767 ( .A1(n3360), .A2(n3363), .ZN(n2124) );
  OAI21_X2 U2768 ( .B1(n3371), .B2(n2136), .A(n2134), .ZN(n3383) );
  NOR2_X2 U2769 ( .A1(n3383), .A2(n3384), .ZN(n3382) );
  INV_X1 U2770 ( .A(n2542), .ZN(n2141) );
  OAI21_X2 U2771 ( .B1(n2141), .B2(n2140), .A(n2139), .ZN(n2570) );
  NAND2_X1 U2772 ( .A1(n2249), .A2(n2146), .ZN(n2145) );
  AOI21_X2 U2773 ( .B1(n3355), .B2(n2591), .A(n2074), .ZN(n3395) );
  AND2_X2 U2774 ( .A1(n2149), .A2(n2148), .ZN(n3355) );
  NAND2_X1 U2775 ( .A1(n2410), .A2(n2046), .ZN(n2991) );
  INV_X1 U2776 ( .A(n2899), .ZN(n2336) );
  NAND2_X1 U2777 ( .A1(n3044), .A2(n3439), .ZN(n3092) );
  NAND2_X1 U2778 ( .A1(n3968), .A2(n3665), .ZN(n3945) );
  NAND2_X1 U2779 ( .A1(n2275), .A2(n2247), .ZN(n2291) );
  NAND2_X1 U2780 ( .A1(n2163), .A2(n4388), .ZN(n2162) );
  XNOR2_X1 U2781 ( .A(n2164), .B(n3621), .ZN(n2163) );
  NOR2_X1 U2782 ( .A1(n4431), .A2(n2086), .ZN(n2164) );
  INV_X1 U2783 ( .A(n3615), .ZN(n2168) );
  NAND2_X1 U2784 ( .A1(n2168), .A2(n2170), .ZN(n3129) );
  INV_X1 U2785 ( .A(n3127), .ZN(n2171) );
  NAND3_X1 U2786 ( .A1(n2234), .A2(n2177), .A3(n2175), .ZN(n2273) );
  NAND4_X1 U2787 ( .A1(n2177), .A2(n2234), .A3(n2176), .A4(n2066), .ZN(n2267)
         );
  NOR2_X1 U2788 ( .A1(n3960), .A2(n3936), .ZN(n3937) );
  INV_X1 U2789 ( .A(n4485), .ZN(n2191) );
  INV_X1 U2790 ( .A(n2267), .ZN(n2249) );
  INV_X1 U2791 ( .A(n3641), .ZN(n2207) );
  NAND2_X1 U2792 ( .A1(n3641), .A2(n2197), .ZN(n2194) );
  NOR2_X1 U2793 ( .A1(n3641), .A2(n3640), .ZN(n3934) );
  NAND2_X1 U2794 ( .A1(n2971), .A2(n2065), .ZN(n2220) );
  NAND2_X1 U2795 ( .A1(n2221), .A2(n2220), .ZN(n3041) );
  NAND3_X1 U2796 ( .A1(n2051), .A2(n2224), .A3(n2226), .ZN(n2222) );
  NAND2_X1 U2797 ( .A1(n3655), .A2(n2079), .ZN(n2228) );
  NAND2_X1 U2798 ( .A1(n2228), .A2(n2229), .ZN(n3743) );
  INV_X1 U2799 ( .A(n2236), .ZN(n2231) );
  NAND2_X1 U2800 ( .A1(n2282), .A2(n2250), .ZN(n2760) );
  OR2_X1 U2801 ( .A1(n2375), .A2(n2912), .ZN(n2376) );
  AND2_X1 U2802 ( .A1(n2915), .A2(n2911), .ZN(n2912) );
  INV_X1 U2803 ( .A(n2322), .ZN(n2323) );
  CLKBUF_X1 U2804 ( .A(n2904), .Z(n2905) );
  NAND2_X1 U2805 ( .A1(n3239), .A2(n3636), .ZN(n3979) );
  NAND2_X1 U2806 ( .A1(n3784), .A2(n3767), .ZN(n3766) );
  OAI21_X2 U2807 ( .B1(n3319), .B2(n3320), .A(n2621), .ZN(n3371) );
  AOI21_X2 U2808 ( .B1(n3395), .B2(n3391), .A(n3392), .ZN(n3319) );
  NAND2_X1 U2809 ( .A1(n3987), .A2(n3694), .ZN(n3993) );
  NOR3_X4 U2810 ( .A1(n3382), .A2(n3311), .A3(n3310), .ZN(n3309) );
  AND2_X1 U2811 ( .A1(n3765), .A2(n3786), .ZN(n2236) );
  AND2_X1 U2812 ( .A1(n2805), .A2(n2804), .ZN(n2237) );
  NAND2_X1 U2813 ( .A1(n3806), .A2(n3779), .ZN(n2238) );
  OR2_X1 U2814 ( .A1(n3848), .A2(n3466), .ZN(n3540) );
  NAND2_X1 U2815 ( .A1(n3582), .A2(n2644), .ZN(n2350) );
  AND2_X1 U2816 ( .A1(n3803), .A2(n3801), .ZN(n3673) );
  INV_X1 U2817 ( .A(IR_REG_27__SCAN_IN), .ZN(n2283) );
  AND2_X1 U2818 ( .A1(n3545), .A2(n3544), .ZN(n3674) );
  INV_X1 U2819 ( .A(IR_REG_21__SCAN_IN), .ZN(n2247) );
  NAND2_X1 U2820 ( .A1(n2321), .A2(n2323), .ZN(n2324) );
  INV_X1 U2821 ( .A(n3295), .ZN(n2555) );
  OAI21_X1 U2822 ( .B1(n3652), .B2(n3793), .A(n3651), .ZN(n3653) );
  AOI21_X1 U2823 ( .B1(n3031), .B2(n3149), .A(n3155), .ZN(n2462) );
  INV_X1 U2824 ( .A(n4277), .ZN(n2298) );
  AND2_X1 U2825 ( .A1(n2686), .A2(REG3_REG_25__SCAN_IN), .ZN(n2700) );
  OR2_X1 U2826 ( .A1(n3710), .A2(n3693), .ZN(n3694) );
  AND2_X1 U2827 ( .A1(n2700), .A2(REG3_REG_26__SCAN_IN), .ZN(n2714) );
  INV_X1 U2828 ( .A(n3653), .ZN(n3654) );
  INV_X1 U2829 ( .A(n3935), .ZN(n3922) );
  OR2_X1 U2830 ( .A1(n2444), .A2(n3156), .ZN(n2463) );
  AND2_X1 U2831 ( .A1(n2363), .A2(DATAI_22_), .ZN(n3824) );
  INV_X1 U2832 ( .A(n3626), .ZN(n3636) );
  OR2_X1 U2833 ( .A1(n2540), .A2(n2539), .ZN(n2541) );
  NAND2_X1 U2834 ( .A1(n2363), .A2(DATAI_3_), .ZN(n2343) );
  INV_X1 U2835 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2993) );
  INV_X1 U2836 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3165) );
  INV_X1 U2837 ( .A(n3762), .ZN(n3731) );
  AND2_X1 U2838 ( .A1(n3490), .A2(n3526), .ZN(n3744) );
  INV_X1 U2839 ( .A(n3780), .ZN(n3823) );
  INV_X1 U2840 ( .A(n3926), .ZN(n3893) );
  INV_X1 U2841 ( .A(n3944), .ZN(n3957) );
  INV_X1 U2842 ( .A(n4445), .ZN(n3257) );
  OR2_X1 U2843 ( .A1(n2463), .A2(n3165), .ZN(n2518) );
  NAND2_X1 U2844 ( .A1(n3905), .A2(n4602), .ZN(n3961) );
  AND2_X1 U2845 ( .A1(n3436), .A2(n3445), .ZN(n3509) );
  AND3_X1 U2846 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2395) );
  INV_X1 U2847 ( .A(n3405), .ZN(n4284) );
  AND2_X1 U2848 ( .A1(n2838), .A2(n2837), .ZN(n3588) );
  AND2_X1 U2849 ( .A1(n2769), .A2(n4271), .ZN(n4478) );
  NOR2_X1 U2850 ( .A1(n4296), .A2(n4272), .ZN(n3905) );
  INV_X1 U2851 ( .A(n3902), .ZN(n3965) );
  INV_X1 U2852 ( .A(n3961), .ZN(n4498) );
  NAND2_X1 U2853 ( .A1(n2305), .A2(n2759), .ZN(n2855) );
  AND2_X1 U2854 ( .A1(n2731), .A2(n2730), .ZN(n3080) );
  INV_X1 U2855 ( .A(n4591), .ZN(n4602) );
  INV_X1 U2856 ( .A(n3080), .ZN(n3084) );
  AND2_X1 U2857 ( .A1(n2565), .A2(n2564), .ZN(n3616) );
  AND2_X1 U2858 ( .A1(n2440), .A2(n2422), .ZN(n4323) );
  AND2_X1 U2859 ( .A1(n2822), .A2(n2837), .ZN(n4436) );
  NAND2_X1 U2860 ( .A1(n2751), .A2(n2750), .ZN(n3411) );
  NAND2_X1 U2861 ( .A1(n2756), .A2(STATE_REG_SCAN_IN), .ZN(n4295) );
  NAND4_X1 U2862 ( .A1(n2705), .A2(n2704), .A3(n2703), .A4(n2702), .ZN(n3762)
         );
  NAND2_X1 U2863 ( .A1(n3588), .A2(n2939), .ZN(n4443) );
  AND2_X1 U2864 ( .A1(n3007), .A2(n3006), .ZN(n3902) );
  NAND2_X1 U2865 ( .A1(n4624), .A2(n4602), .ZN(n4201) );
  INV_X1 U2866 ( .A(n4624), .ZN(n4621) );
  NAND2_X1 U2867 ( .A1(n4605), .A2(n4602), .ZN(n4259) );
  INV_X1 U2868 ( .A(n4605), .ZN(n4603) );
  INV_X1 U2869 ( .A(n4526), .ZN(n4525) );
  NAND2_X1 U2870 ( .A1(n2815), .A2(n2814), .ZN(n4526) );
  INV_X1 U2871 ( .A(n4323), .ZN(n4549) );
  AND2_X1 U2872 ( .A1(n2361), .A2(n2342), .ZN(n4275) );
  INV_X1 U2873 ( .A(n3583), .ZN(U4043) );
  NAND4_X1 U2874 ( .A1(n2452), .A2(n2242), .A3(n2241), .A4(n2240), .ZN(n2243)
         );
  INV_X1 U2875 ( .A(IR_REG_25__SCAN_IN), .ZN(n2248) );
  NAND2_X1 U2876 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2250) );
  INV_X1 U2877 ( .A(n2270), .ZN(n2254) );
  NAND2_X1 U2878 ( .A1(n2254), .A2(n2053), .ZN(n2811) );
  NAND2_X1 U2879 ( .A1(n2043), .A2(REG1_REG_16__SCAN_IN), .ZN(n2264) );
  NAND2_X1 U2880 ( .A1(n2353), .A2(REG0_REG_16__SCAN_IN), .ZN(n2263) );
  NAND2_X1 U2881 ( .A1(n2395), .A2(REG3_REG_6__SCAN_IN), .ZN(n2411) );
  NAND2_X1 U2882 ( .A1(n2432), .A2(REG3_REG_8__SCAN_IN), .ZN(n2444) );
  NAND2_X1 U2883 ( .A1(REG3_REG_12__SCAN_IN), .A2(REG3_REG_11__SCAN_IN), .ZN(
        n2257) );
  NAND2_X1 U2884 ( .A1(n2495), .A2(REG3_REG_13__SCAN_IN), .ZN(n2545) );
  INV_X1 U2885 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2544) );
  INV_X1 U2886 ( .A(REG3_REG_15__SCAN_IN), .ZN(n4278) );
  OR2_X1 U2887 ( .A1(n2557), .A2(REG3_REG_16__SCAN_IN), .ZN(n2258) );
  NAND2_X1 U2888 ( .A1(n2557), .A2(REG3_REG_16__SCAN_IN), .ZN(n2574) );
  NAND2_X1 U2889 ( .A1(n2258), .A2(n2574), .ZN(n3347) );
  OR2_X1 U2890 ( .A1(n2040), .A2(n3347), .ZN(n2262) );
  INV_X1 U2891 ( .A(REG2_REG_16__SCAN_IN), .ZN(n2260) );
  OR2_X1 U2892 ( .A1(n2356), .A2(n2260), .ZN(n2261) );
  NAND4_X1 U2893 ( .A1(n2264), .A2(n2263), .A3(n2262), .A4(n2261), .ZN(n3947)
         );
  INV_X1 U2894 ( .A(IR_REG_24__SCAN_IN), .ZN(n2265) );
  NAND2_X1 U2895 ( .A1(n2267), .A2(IR_REG_31__SCAN_IN), .ZN(n2268) );
  MUX2_X1 U2896 ( .A(IR_REG_31__SCAN_IN), .B(n2268), .S(IR_REG_25__SCAN_IN), 
        .Z(n2269) );
  NAND2_X1 U2897 ( .A1(n2269), .A2(n2270), .ZN(n2742) );
  NAND2_X1 U2898 ( .A1(n2294), .A2(n2246), .ZN(n2293) );
  NAND2_X1 U2899 ( .A1(n2293), .A2(IR_REG_31__SCAN_IN), .ZN(n2274) );
  INV_X1 U2900 ( .A(n2275), .ZN(n2276) );
  NAND2_X1 U2901 ( .A1(n2276), .A2(IR_REG_31__SCAN_IN), .ZN(n2277) );
  INV_X1 U2902 ( .A(n2953), .ZN(n2278) );
  NAND2_X1 U2903 ( .A1(n3947), .A2(n2038), .ZN(n2290) );
  NAND2_X1 U2904 ( .A1(n2279), .A2(n2153), .ZN(n2280) );
  NAND2_X1 U2905 ( .A1(n2280), .A2(IR_REG_31__SCAN_IN), .ZN(n2563) );
  NAND2_X1 U2906 ( .A1(n2563), .A2(n2152), .ZN(n2565) );
  NAND2_X1 U2907 ( .A1(n2565), .A2(IR_REG_31__SCAN_IN), .ZN(n2281) );
  XNOR2_X1 U2908 ( .A(n2281), .B(IR_REG_16__SCAN_IN), .ZN(n3617) );
  NAND2_X1 U2909 ( .A1(n2282), .A2(n2286), .ZN(n2284) );
  NAND2_X1 U2910 ( .A1(n2286), .A2(IR_REG_27__SCAN_IN), .ZN(n2287) );
  MUX2_X1 U2911 ( .A(n3617), .B(DATAI_16_), .S(n2363), .Z(n3936) );
  NAND2_X1 U2912 ( .A1(n3936), .A2(n2645), .ZN(n2289) );
  NAND2_X1 U2913 ( .A1(n2290), .A2(n2289), .ZN(n2295) );
  NAND2_X1 U2914 ( .A1(n4269), .A2(n3624), .ZN(n2757) );
  NAND2_X2 U2915 ( .A1(n2757), .A2(n2953), .ZN(n2722) );
  INV_X2 U2916 ( .A(n2722), .ZN(n2783) );
  XNOR2_X1 U2917 ( .A(n2295), .B(n2783), .ZN(n2572) );
  INV_X1 U2918 ( .A(n4270), .ZN(n2296) );
  NAND2_X2 U2919 ( .A1(n2037), .A2(n4591), .ZN(n2658) );
  AOI22_X1 U2920 ( .A1(n3947), .A2(n2697), .B1(n2644), .B2(n3936), .ZN(n2571)
         );
  NAND2_X1 U2921 ( .A1(n2353), .A2(REG0_REG_1__SCAN_IN), .ZN(n2924) );
  INV_X1 U2922 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2297) );
  OR2_X1 U2923 ( .A1(n2354), .A2(n2297), .ZN(n2923) );
  NAND2_X1 U2924 ( .A1(n2543), .A2(REG1_REG_1__SCAN_IN), .ZN(n2925) );
  INV_X1 U2925 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2841) );
  OR2_X1 U2926 ( .A1(n2356), .A2(n2841), .ZN(n2922) );
  NAND2_X1 U2927 ( .A1(n2304), .A2(n2038), .ZN(n2302) );
  NAND2_X1 U2928 ( .A1(n4492), .A2(n2645), .ZN(n2301) );
  NAND2_X1 U2929 ( .A1(n2302), .A2(n2301), .ZN(n2303) );
  XNOR2_X1 U2930 ( .A(n2321), .B(n2322), .ZN(n2852) );
  INV_X1 U2931 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2314) );
  NAND2_X1 U2932 ( .A1(n2043), .A2(REG1_REG_0__SCAN_IN), .ZN(n2310) );
  NAND2_X1 U2933 ( .A1(n2353), .A2(REG0_REG_0__SCAN_IN), .ZN(n2309) );
  INV_X1 U2934 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2306) );
  OR2_X1 U2935 ( .A1(n2040), .A2(n2306), .ZN(n2308) );
  INV_X1 U2936 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2861) );
  OR2_X1 U2937 ( .A1(n2356), .A2(n2861), .ZN(n2307) );
  NAND2_X1 U2938 ( .A1(n3584), .A2(n2644), .ZN(n2313) );
  NAND2_X1 U2939 ( .A1(n4493), .A2(n2645), .ZN(n2318) );
  OAI211_X1 U2940 ( .C1(n2305), .C2(n2314), .A(n2313), .B(n2318), .ZN(n2864)
         );
  NAND2_X1 U2941 ( .A1(n3584), .A2(n2697), .ZN(n2317) );
  INV_X1 U2942 ( .A(n2305), .ZN(n2315) );
  AOI22_X1 U2943 ( .A1(n4493), .A2(n2644), .B1(n2315), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2316) );
  NAND2_X1 U2944 ( .A1(n2317), .A2(n2316), .ZN(n2863) );
  NAND2_X1 U2945 ( .A1(n2864), .A2(n2863), .ZN(n2320) );
  NAND2_X1 U2946 ( .A1(n2318), .A2(n2783), .ZN(n2319) );
  NAND2_X1 U2947 ( .A1(n2320), .A2(n2319), .ZN(n2853) );
  NAND2_X1 U2948 ( .A1(n2852), .A2(n2853), .ZN(n2325) );
  NAND2_X1 U2949 ( .A1(n2325), .A2(n2324), .ZN(n2896) );
  INV_X1 U2950 ( .A(n2896), .ZN(n2337) );
  NAND2_X1 U2951 ( .A1(n2353), .A2(REG0_REG_2__SCAN_IN), .ZN(n2329) );
  NAND2_X1 U2952 ( .A1(n2042), .A2(REG1_REG_2__SCAN_IN), .ZN(n2328) );
  INV_X1 U2953 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3060) );
  INV_X1 U2954 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2840) );
  OR2_X1 U2955 ( .A1(n2356), .A2(n2840), .ZN(n2326) );
  NAND2_X1 U2956 ( .A1(n4480), .A2(n2038), .ZN(n2331) );
  MUX2_X1 U2957 ( .A(n4276), .B(DATAI_2_), .S(n2363), .Z(n3058) );
  NAND2_X1 U2958 ( .A1(n3058), .A2(n2645), .ZN(n2330) );
  NAND2_X1 U2959 ( .A1(n2331), .A2(n2330), .ZN(n2332) );
  XNOR2_X1 U2960 ( .A(n2332), .B(n2783), .ZN(n2334) );
  AOI22_X1 U2961 ( .A1(n4480), .A2(n2697), .B1(n2644), .B2(n3058), .ZN(n2333)
         );
  NAND2_X1 U2962 ( .A1(n2334), .A2(n2333), .ZN(n2338) );
  NAND2_X1 U2963 ( .A1(n2335), .A2(n2338), .ZN(n2899) );
  NAND2_X1 U2964 ( .A1(n2337), .A2(n2336), .ZN(n2897) );
  NAND2_X1 U2965 ( .A1(n2897), .A2(n2338), .ZN(n2904) );
  NAND2_X1 U2966 ( .A1(n2339), .A2(IR_REG_31__SCAN_IN), .ZN(n2341) );
  NAND2_X1 U2967 ( .A1(n2341), .A2(n2340), .ZN(n2361) );
  OR2_X1 U2968 ( .A1(n2341), .A2(n2340), .ZN(n2342) );
  NAND2_X1 U2969 ( .A1(n3432), .A2(n2645), .ZN(n2351) );
  OR2_X1 U2970 ( .A1(n2039), .A2(REG3_REG_3__SCAN_IN), .ZN(n2349) );
  NAND2_X1 U2971 ( .A1(n2043), .A2(REG1_REG_3__SCAN_IN), .ZN(n2348) );
  NAND2_X1 U2972 ( .A1(n2353), .A2(REG0_REG_3__SCAN_IN), .ZN(n2347) );
  INV_X1 U2973 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2345) );
  OR2_X1 U2974 ( .A1(n2356), .A2(n2345), .ZN(n2346) );
  NAND2_X1 U2975 ( .A1(n2351), .A2(n2350), .ZN(n2352) );
  XNOR2_X1 U2976 ( .A(n2352), .B(n2722), .ZN(n2372) );
  AOI22_X1 U2977 ( .A1(n3582), .A2(n2697), .B1(n2644), .B2(n3432), .ZN(n2373)
         );
  XNOR2_X1 U2978 ( .A(n2372), .B(n2373), .ZN(n2903) );
  NAND2_X1 U2979 ( .A1(n2353), .A2(REG0_REG_4__SCAN_IN), .ZN(n2360) );
  NAND2_X1 U2980 ( .A1(n2042), .A2(REG1_REG_4__SCAN_IN), .ZN(n2359) );
  XNOR2_X1 U2981 ( .A(REG3_REG_4__SCAN_IN), .B(REG3_REG_3__SCAN_IN), .ZN(n2947) );
  INV_X1 U2982 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2355) );
  OR2_X1 U2983 ( .A1(n2356), .A2(n2355), .ZN(n2357) );
  NAND2_X1 U2984 ( .A1(n3581), .A2(n2644), .ZN(n2365) );
  NAND2_X1 U2985 ( .A1(n2361), .A2(IR_REG_31__SCAN_IN), .ZN(n2362) );
  XNOR2_X1 U2986 ( .A(n2362), .B(IR_REG_4__SCAN_IN), .ZN(n4274) );
  MUX2_X1 U2987 ( .A(n4274), .B(DATAI_4_), .S(n2363), .Z(n2917) );
  NAND2_X1 U2988 ( .A1(n2917), .A2(n2645), .ZN(n2364) );
  NAND2_X1 U2989 ( .A1(n2365), .A2(n2364), .ZN(n2366) );
  XNOR2_X1 U2990 ( .A(n2366), .B(n2722), .ZN(n2371) );
  AOI22_X1 U2991 ( .A1(n3581), .A2(n2697), .B1(n2038), .B2(n2917), .ZN(n2370)
         );
  INV_X1 U2992 ( .A(n2370), .ZN(n2367) );
  NAND2_X1 U2993 ( .A1(n2371), .A2(n2367), .ZN(n2369) );
  AND2_X1 U2994 ( .A1(n2903), .A2(n2369), .ZN(n2368) );
  NAND2_X1 U2995 ( .A1(n2904), .A2(n2368), .ZN(n2377) );
  INV_X1 U2996 ( .A(n2369), .ZN(n2375) );
  XNOR2_X1 U2997 ( .A(n2371), .B(n2370), .ZN(n2915) );
  INV_X1 U2998 ( .A(n2372), .ZN(n2374) );
  NAND2_X1 U2999 ( .A1(n2374), .A2(n2373), .ZN(n2911) );
  NAND2_X1 U3000 ( .A1(n2353), .A2(REG0_REG_5__SCAN_IN), .ZN(n2385) );
  NAND2_X1 U3001 ( .A1(n2042), .A2(REG1_REG_5__SCAN_IN), .ZN(n2384) );
  INV_X1 U3002 ( .A(n2395), .ZN(n2381) );
  INV_X1 U3003 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2379) );
  NAND2_X1 U3004 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2378) );
  NAND2_X1 U3005 ( .A1(n2379), .A2(n2378), .ZN(n2380) );
  NAND2_X1 U3006 ( .A1(n2381), .A2(n2380), .ZN(n3027) );
  OR2_X1 U3007 ( .A1(n2040), .A2(n3027), .ZN(n2383) );
  OR2_X1 U3008 ( .A1(n2356), .A2(n3116), .ZN(n2382) );
  NAND4_X1 U3009 ( .A1(n2385), .A2(n2384), .A3(n2383), .A4(n2382), .ZN(n3580)
         );
  NAND2_X1 U3010 ( .A1(n3580), .A2(n2644), .ZN(n2389) );
  NAND2_X1 U3011 ( .A1(n2386), .A2(IR_REG_31__SCAN_IN), .ZN(n2387) );
  XNOR2_X1 U3012 ( .A(n2387), .B(IR_REG_5__SCAN_IN), .ZN(n3134) );
  MUX2_X1 U3013 ( .A(n3134), .B(DATAI_5_), .S(n2363), .Z(n3018) );
  NAND2_X1 U3014 ( .A1(n3018), .A2(n2645), .ZN(n2388) );
  NAND2_X1 U3015 ( .A1(n2389), .A2(n2388), .ZN(n2390) );
  AOI22_X1 U3016 ( .A1(n3580), .A2(n2697), .B1(n2644), .B2(n3018), .ZN(n2392)
         );
  XNOR2_X1 U3017 ( .A(n2391), .B(n2392), .ZN(n2958) );
  INV_X1 U3018 ( .A(n2391), .ZN(n2393) );
  NOR2_X1 U3019 ( .A1(n2393), .A2(n2392), .ZN(n2394) );
  NAND2_X1 U3020 ( .A1(n2353), .A2(REG0_REG_6__SCAN_IN), .ZN(n2399) );
  NAND2_X1 U3021 ( .A1(n2043), .A2(REG1_REG_6__SCAN_IN), .ZN(n2398) );
  OAI21_X1 U3022 ( .B1(n2395), .B2(REG3_REG_6__SCAN_IN), .A(n2411), .ZN(n3010)
         );
  OR2_X1 U3023 ( .A1(n2040), .A2(n3010), .ZN(n2397) );
  INV_X1 U3024 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3011) );
  OR2_X1 U3025 ( .A1(n2832), .A2(n3011), .ZN(n2396) );
  NAND4_X1 U3026 ( .A1(n2399), .A2(n2398), .A3(n2397), .A4(n2396), .ZN(n3579)
         );
  NAND2_X1 U3027 ( .A1(n3579), .A2(n2644), .ZN(n2402) );
  NOR2_X1 U3028 ( .A1(n2386), .A2(IR_REG_5__SCAN_IN), .ZN(n2454) );
  OR2_X1 U3029 ( .A1(n2454), .A2(n2597), .ZN(n2400) );
  XNOR2_X1 U3030 ( .A(n2400), .B(IR_REG_6__SCAN_IN), .ZN(n3135) );
  MUX2_X1 U3031 ( .A(n3135), .B(DATAI_6_), .S(n2363), .Z(n3038) );
  NAND2_X1 U3032 ( .A1(n3038), .A2(n2645), .ZN(n2401) );
  NAND2_X1 U3033 ( .A1(n2402), .A2(n2401), .ZN(n2403) );
  XNOR2_X1 U3034 ( .A(n2403), .B(n2722), .ZN(n2406) );
  NAND2_X1 U3035 ( .A1(n3579), .A2(n2697), .ZN(n2405) );
  NAND2_X1 U3036 ( .A1(n3038), .A2(n2644), .ZN(n2404) );
  NAND2_X1 U3037 ( .A1(n2405), .A2(n2404), .ZN(n2407) );
  NAND2_X1 U3038 ( .A1(n2406), .A2(n2407), .ZN(n2964) );
  NAND2_X1 U3039 ( .A1(n2965), .A2(n2964), .ZN(n2410) );
  INV_X1 U3040 ( .A(n2406), .ZN(n2409) );
  INV_X1 U3041 ( .A(n2407), .ZN(n2408) );
  NAND2_X1 U3042 ( .A1(n2409), .A2(n2408), .ZN(n2963) );
  NAND2_X1 U3043 ( .A1(n2353), .A2(REG0_REG_7__SCAN_IN), .ZN(n2417) );
  NAND2_X1 U3044 ( .A1(n2042), .A2(REG1_REG_7__SCAN_IN), .ZN(n2416) );
  AND2_X1 U3045 ( .A1(n2411), .A2(n2993), .ZN(n2412) );
  OR2_X1 U3046 ( .A1(n2412), .A2(n2432), .ZN(n3050) );
  OR2_X1 U3047 ( .A1(n2039), .A2(n3050), .ZN(n2415) );
  INV_X1 U3048 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2413) );
  OR2_X1 U3049 ( .A1(n2356), .A2(n2413), .ZN(n2414) );
  NAND4_X1 U3050 ( .A1(n2417), .A2(n2416), .A3(n2415), .A4(n2414), .ZN(n3099)
         );
  NAND2_X1 U3051 ( .A1(n3099), .A2(n2038), .ZN(n2424) );
  INV_X1 U3052 ( .A(IR_REG_6__SCAN_IN), .ZN(n2418) );
  NAND2_X1 U3053 ( .A1(n2454), .A2(n2418), .ZN(n2419) );
  NAND2_X1 U3054 ( .A1(n2419), .A2(IR_REG_31__SCAN_IN), .ZN(n2421) );
  INV_X1 U3055 ( .A(IR_REG_7__SCAN_IN), .ZN(n2420) );
  NAND2_X1 U3056 ( .A1(n2421), .A2(n2420), .ZN(n2440) );
  OR2_X1 U3057 ( .A1(n2421), .A2(n2420), .ZN(n2422) );
  MUX2_X1 U3058 ( .A(n4323), .B(DATAI_7_), .S(n2363), .Z(n3098) );
  NAND2_X1 U3059 ( .A1(n3098), .A2(n2645), .ZN(n2423) );
  NAND2_X1 U3060 ( .A1(n2424), .A2(n2423), .ZN(n2425) );
  XNOR2_X1 U3061 ( .A(n2425), .B(n2783), .ZN(n2427) );
  AOI22_X1 U3062 ( .A1(n3099), .A2(n2697), .B1(n2644), .B2(n3098), .ZN(n2428)
         );
  XNOR2_X1 U3063 ( .A(n2427), .B(n2428), .ZN(n2989) );
  INV_X1 U3064 ( .A(n2989), .ZN(n2426) );
  INV_X1 U3065 ( .A(n2427), .ZN(n2430) );
  INV_X1 U3066 ( .A(n2428), .ZN(n2429) );
  NAND2_X1 U3067 ( .A1(n2430), .A2(n2429), .ZN(n2431) );
  NAND2_X1 U3068 ( .A1(n2353), .A2(REG0_REG_8__SCAN_IN), .ZN(n2439) );
  NAND2_X1 U3069 ( .A1(n2043), .A2(REG1_REG_8__SCAN_IN), .ZN(n2438) );
  OR2_X1 U3070 ( .A1(n2432), .A2(REG3_REG_8__SCAN_IN), .ZN(n2433) );
  AND2_X1 U3071 ( .A1(n2444), .A2(n2433), .ZN(n4468) );
  INV_X1 U3072 ( .A(n4468), .ZN(n2434) );
  OR2_X1 U3073 ( .A1(n2039), .A2(n2434), .ZN(n2437) );
  INV_X1 U3074 ( .A(REG2_REG_8__SCAN_IN), .ZN(n2435) );
  OR2_X1 U3075 ( .A1(n2832), .A2(n2435), .ZN(n2436) );
  NAND4_X1 U3076 ( .A1(n2439), .A2(n2438), .A3(n2437), .A4(n2436), .ZN(n3578)
         );
  NAND2_X1 U3077 ( .A1(n3578), .A2(n2697), .ZN(n2443) );
  NAND2_X1 U3078 ( .A1(n2440), .A2(IR_REG_31__SCAN_IN), .ZN(n2441) );
  XNOR2_X1 U3079 ( .A(n2441), .B(IR_REG_8__SCAN_IN), .ZN(n4546) );
  MUX2_X1 U3080 ( .A(n4546), .B(DATAI_8_), .S(n2363), .Z(n3183) );
  NAND2_X1 U3081 ( .A1(n3183), .A2(n2644), .ZN(n2442) );
  NAND2_X1 U3082 ( .A1(n2443), .A2(n2442), .ZN(n3149) );
  NAND2_X1 U3083 ( .A1(n2353), .A2(REG0_REG_9__SCAN_IN), .ZN(n2450) );
  NAND2_X1 U3084 ( .A1(n2042), .A2(REG1_REG_9__SCAN_IN), .ZN(n2449) );
  NAND2_X1 U3085 ( .A1(n2444), .A2(n3156), .ZN(n2445) );
  NAND2_X1 U3086 ( .A1(n2463), .A2(n2445), .ZN(n3105) );
  OR2_X1 U3087 ( .A1(n2040), .A2(n3105), .ZN(n2448) );
  INV_X1 U3088 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2446) );
  OR2_X1 U3089 ( .A1(n2832), .A2(n2446), .ZN(n2447) );
  NAND4_X1 U3090 ( .A1(n2450), .A2(n2449), .A3(n2448), .A4(n2447), .ZN(n3577)
         );
  NAND2_X1 U3091 ( .A1(n3577), .A2(n2644), .ZN(n2457) );
  INV_X1 U3092 ( .A(IR_REG_8__SCAN_IN), .ZN(n2451) );
  AND2_X1 U3093 ( .A1(n2452), .A2(n2451), .ZN(n2453) );
  NAND2_X1 U3094 ( .A1(n2454), .A2(n2453), .ZN(n2470) );
  NAND2_X1 U3095 ( .A1(n2470), .A2(IR_REG_31__SCAN_IN), .ZN(n2455) );
  XNOR2_X1 U3096 ( .A(n2455), .B(IR_REG_9__SCAN_IN), .ZN(n4544) );
  MUX2_X1 U3097 ( .A(n4544), .B(DATAI_9_), .S(n2363), .Z(n3206) );
  NAND2_X1 U3098 ( .A1(n3206), .A2(n2645), .ZN(n2456) );
  NAND2_X1 U3099 ( .A1(n2457), .A2(n2456), .ZN(n2458) );
  XNOR2_X1 U3100 ( .A(n2458), .B(n2783), .ZN(n2476) );
  AOI22_X1 U3101 ( .A1(n3577), .A2(n2697), .B1(n2038), .B2(n3206), .ZN(n2475)
         );
  XNOR2_X1 U3102 ( .A(n2476), .B(n2475), .ZN(n3155) );
  NAND2_X1 U3103 ( .A1(n3578), .A2(n2644), .ZN(n2460) );
  NAND2_X1 U3104 ( .A1(n3183), .A2(n2645), .ZN(n2459) );
  NAND2_X1 U3105 ( .A1(n2460), .A2(n2459), .ZN(n2461) );
  XNOR2_X1 U3106 ( .A(n2461), .B(n2722), .ZN(n3032) );
  OAI21_X2 U3107 ( .B1(n3031), .B2(n3149), .A(n3032), .ZN(n3151) );
  NAND2_X1 U3108 ( .A1(n2462), .A2(n3151), .ZN(n3152) );
  NAND2_X1 U3109 ( .A1(n2042), .A2(REG1_REG_10__SCAN_IN), .ZN(n2469) );
  NAND2_X1 U3110 ( .A1(n2353), .A2(REG0_REG_10__SCAN_IN), .ZN(n2468) );
  NAND2_X1 U3111 ( .A1(n2463), .A2(n3165), .ZN(n2464) );
  AND2_X1 U3112 ( .A1(n2518), .A2(n2464), .ZN(n4461) );
  INV_X1 U3113 ( .A(n4461), .ZN(n3169) );
  OR2_X1 U3114 ( .A1(n2039), .A2(n3169), .ZN(n2467) );
  INV_X1 U3115 ( .A(REG2_REG_10__SCAN_IN), .ZN(n2465) );
  OR2_X1 U3116 ( .A1(n2356), .A2(n2465), .ZN(n2466) );
  NAND4_X1 U3117 ( .A1(n2469), .A2(n2468), .A3(n2467), .A4(n2466), .ZN(n3576)
         );
  NAND2_X1 U3118 ( .A1(n3576), .A2(n2644), .ZN(n2473) );
  NAND2_X1 U3119 ( .A1(n2502), .A2(IR_REG_31__SCAN_IN), .ZN(n2471) );
  XNOR2_X1 U3120 ( .A(n2471), .B(IR_REG_10__SCAN_IN), .ZN(n4542) );
  MUX2_X1 U3121 ( .A(n4542), .B(DATAI_10_), .S(n2363), .Z(n3269) );
  NAND2_X1 U3122 ( .A1(n3269), .A2(n2645), .ZN(n2472) );
  NAND2_X1 U3123 ( .A1(n2473), .A2(n2472), .ZN(n2474) );
  XNOR2_X1 U3124 ( .A(n2474), .B(n2722), .ZN(n2480) );
  AOI22_X1 U3125 ( .A1(n3576), .A2(n2697), .B1(n2038), .B2(n3269), .ZN(n2478)
         );
  XNOR2_X1 U3126 ( .A(n2480), .B(n2478), .ZN(n3163) );
  NAND2_X1 U3127 ( .A1(n2476), .A2(n2475), .ZN(n3162) );
  AND2_X1 U3128 ( .A1(n3163), .A2(n3162), .ZN(n2477) );
  NAND2_X1 U3129 ( .A1(n3152), .A2(n2477), .ZN(n3171) );
  INV_X1 U3130 ( .A(n2478), .ZN(n2479) );
  NAND2_X1 U3131 ( .A1(n2480), .A2(n2479), .ZN(n3170) );
  NAND2_X1 U3132 ( .A1(n2353), .A2(REG0_REG_13__SCAN_IN), .ZN(n2486) );
  NAND2_X1 U3133 ( .A1(n2043), .A2(REG1_REG_13__SCAN_IN), .ZN(n2485) );
  OR2_X1 U3134 ( .A1(n2495), .A2(REG3_REG_13__SCAN_IN), .ZN(n2481) );
  NAND2_X1 U3135 ( .A1(n2545), .A2(n2481), .ZN(n3261) );
  OR2_X1 U3136 ( .A1(n2040), .A2(n3261), .ZN(n2484) );
  INV_X1 U3137 ( .A(REG2_REG_13__SCAN_IN), .ZN(n2482) );
  OR2_X1 U3138 ( .A1(n2356), .A2(n2482), .ZN(n2483) );
  NAND4_X1 U3139 ( .A1(n2486), .A2(n2485), .A3(n2484), .A4(n2483), .ZN(n3627)
         );
  NAND2_X1 U3140 ( .A1(n3627), .A2(n2644), .ZN(n2490) );
  OR2_X1 U3141 ( .A1(n2487), .A2(n2597), .ZN(n2488) );
  XNOR2_X1 U3142 ( .A(n2488), .B(IR_REG_13__SCAN_IN), .ZN(n4537) );
  MUX2_X1 U3143 ( .A(n4537), .B(DATAI_13_), .S(n2363), .Z(n3626) );
  NAND2_X1 U3144 ( .A1(n3626), .A2(n2645), .ZN(n2489) );
  NAND2_X1 U3145 ( .A1(n2490), .A2(n2489), .ZN(n2491) );
  XNOR2_X1 U3146 ( .A(n2491), .B(n2722), .ZN(n2512) );
  NAND2_X1 U3147 ( .A1(n3627), .A2(n2697), .ZN(n2493) );
  NAND2_X1 U31480 ( .A1(n3626), .A2(n2038), .ZN(n2492) );
  NAND2_X1 U31490 ( .A1(n2493), .A2(n2492), .ZN(n2513) );
  NAND2_X1 U3150 ( .A1(n2512), .A2(n2513), .ZN(n3252) );
  NAND2_X1 U3151 ( .A1(n2353), .A2(REG0_REG_12__SCAN_IN), .ZN(n2501) );
  NAND2_X1 U3152 ( .A1(n2043), .A2(REG1_REG_12__SCAN_IN), .ZN(n2500) );
  INV_X1 U3153 ( .A(n2518), .ZN(n2494) );
  AOI21_X1 U3154 ( .B1(n2494), .B2(REG3_REG_11__SCAN_IN), .A(
        REG3_REG_12__SCAN_IN), .ZN(n2496) );
  OR2_X1 U3155 ( .A1(n2496), .A2(n2495), .ZN(n3173) );
  OR2_X1 U3156 ( .A1(n2040), .A2(n3173), .ZN(n2499) );
  INV_X1 U3157 ( .A(REG2_REG_12__SCAN_IN), .ZN(n2497) );
  OR2_X1 U3158 ( .A1(n2832), .A2(n2497), .ZN(n2498) );
  NAND2_X1 U3159 ( .A1(n4445), .A2(n2697), .ZN(n2508) );
  NAND2_X1 U3160 ( .A1(n2503), .A2(IR_REG_31__SCAN_IN), .ZN(n2525) );
  INV_X1 U3161 ( .A(IR_REG_11__SCAN_IN), .ZN(n2504) );
  NAND2_X1 U3162 ( .A1(n2525), .A2(n2504), .ZN(n2505) );
  NAND2_X1 U3163 ( .A1(n2505), .A2(IR_REG_31__SCAN_IN), .ZN(n2506) );
  XNOR2_X1 U3164 ( .A(n2506), .B(IR_REG_12__SCAN_IN), .ZN(n3142) );
  MUX2_X1 U3165 ( .A(n3142), .B(DATAI_12_), .S(n2363), .Z(n3235) );
  NAND2_X1 U3166 ( .A1(n3235), .A2(n2644), .ZN(n2507) );
  NAND2_X1 U3167 ( .A1(n4445), .A2(n2038), .ZN(n2510) );
  NAND2_X1 U3168 ( .A1(n3235), .A2(n2645), .ZN(n2509) );
  NAND2_X1 U3169 ( .A1(n2510), .A2(n2509), .ZN(n2511) );
  XNOR2_X1 U3170 ( .A(n2511), .B(n2783), .ZN(n3247) );
  NAND3_X1 U3171 ( .A1(n3252), .A2(n3249), .A3(n3247), .ZN(n2516) );
  INV_X1 U3172 ( .A(n2512), .ZN(n2515) );
  INV_X1 U3173 ( .A(n2513), .ZN(n2514) );
  NAND2_X1 U3174 ( .A1(n2515), .A2(n2514), .ZN(n3251) );
  INV_X1 U3175 ( .A(n2538), .ZN(n2533) );
  OAI21_X1 U3176 ( .B1(n3247), .B2(n3249), .A(n3252), .ZN(n2517) );
  INV_X1 U3177 ( .A(n2517), .ZN(n2531) );
  NAND2_X1 U3178 ( .A1(n2353), .A2(REG0_REG_11__SCAN_IN), .ZN(n2524) );
  NAND2_X1 U3179 ( .A1(n2043), .A2(REG1_REG_11__SCAN_IN), .ZN(n2523) );
  XNOR2_X1 U3180 ( .A(n2518), .B(REG3_REG_11__SCAN_IN), .ZN(n4455) );
  INV_X1 U3181 ( .A(n4455), .ZN(n2519) );
  OR2_X1 U3182 ( .A1(n2039), .A2(n2519), .ZN(n2522) );
  INV_X1 U3183 ( .A(REG2_REG_11__SCAN_IN), .ZN(n2520) );
  OR2_X1 U3184 ( .A1(n2832), .A2(n2520), .ZN(n2521) );
  NAND4_X1 U3185 ( .A1(n2524), .A2(n2523), .A3(n2522), .A4(n2521), .ZN(n3575)
         );
  NAND2_X1 U3186 ( .A1(n3575), .A2(n2038), .ZN(n2527) );
  XNOR2_X1 U3187 ( .A(n2525), .B(IR_REG_11__SCAN_IN), .ZN(n4540) );
  MUX2_X1 U3188 ( .A(n4540), .B(DATAI_11_), .S(n2363), .Z(n4457) );
  NAND2_X1 U3189 ( .A1(n4457), .A2(n2645), .ZN(n2526) );
  NAND2_X1 U3190 ( .A1(n2527), .A2(n2526), .ZN(n2528) );
  XNOR2_X1 U3191 ( .A(n2528), .B(n2783), .ZN(n2537) );
  INV_X1 U3192 ( .A(n2537), .ZN(n2530) );
  AOI22_X1 U3193 ( .A1(n3575), .A2(n2697), .B1(n2644), .B2(n4457), .ZN(n2536)
         );
  INV_X1 U3194 ( .A(n2536), .ZN(n2529) );
  NAND2_X1 U3195 ( .A1(n2530), .A2(n2529), .ZN(n3225) );
  AND2_X1 U3196 ( .A1(n2531), .A2(n3225), .ZN(n2532) );
  AND2_X1 U3197 ( .A1(n3170), .A2(n2535), .ZN(n2534) );
  NAND2_X1 U3198 ( .A1(n3171), .A2(n2534), .ZN(n2542) );
  INV_X1 U3199 ( .A(n2535), .ZN(n2540) );
  NAND2_X1 U3200 ( .A1(n2537), .A2(n2536), .ZN(n3223) );
  AND2_X1 U3201 ( .A1(n3223), .A2(n2538), .ZN(n2539) );
  NAND2_X1 U3202 ( .A1(n2353), .A2(REG0_REG_14__SCAN_IN), .ZN(n2550) );
  NAND2_X1 U3203 ( .A1(n2042), .A2(REG1_REG_14__SCAN_IN), .ZN(n2549) );
  NAND2_X1 U3204 ( .A1(n2545), .A2(n2544), .ZN(n2546) );
  NAND2_X1 U3205 ( .A1(n2556), .A2(n2546), .ZN(n3980) );
  OR2_X1 U3206 ( .A1(n2039), .A2(n3980), .ZN(n2548) );
  INV_X1 U3207 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3981) );
  OR2_X1 U3208 ( .A1(n2356), .A2(n3981), .ZN(n2547) );
  NAND4_X1 U3209 ( .A1(n2550), .A2(n2549), .A3(n2548), .A4(n2547), .ZN(n3574)
         );
  NAND2_X1 U32100 ( .A1(n3574), .A2(n2038), .ZN(n2553) );
  OR2_X1 U32110 ( .A1(n2279), .A2(n2597), .ZN(n2551) );
  XNOR2_X1 U32120 ( .A(n2551), .B(IR_REG_14__SCAN_IN), .ZN(n4273) );
  MUX2_X1 U32130 ( .A(n4273), .B(DATAI_14_), .S(n2363), .Z(n3978) );
  NAND2_X1 U32140 ( .A1(n3978), .A2(n2645), .ZN(n2552) );
  NAND2_X1 U32150 ( .A1(n2553), .A2(n2552), .ZN(n2554) );
  XNOR2_X1 U32160 ( .A(n2554), .B(n2783), .ZN(n3296) );
  AOI22_X1 U32170 ( .A1(n3574), .A2(n2697), .B1(n2038), .B2(n3978), .ZN(n3295)
         );
  NAND2_X1 U32180 ( .A1(n2042), .A2(REG1_REG_15__SCAN_IN), .ZN(n2562) );
  NAND2_X1 U32190 ( .A1(n2353), .A2(REG0_REG_15__SCAN_IN), .ZN(n2561) );
  AND2_X1 U32200 ( .A1(n2556), .A2(n4278), .ZN(n2558) );
  OR2_X1 U32210 ( .A1(n2558), .A2(n2557), .ZN(n4294) );
  OR2_X1 U32220 ( .A1(n2039), .A2(n4294), .ZN(n2560) );
  INV_X1 U32230 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3962) );
  OR2_X1 U32240 ( .A1(n2832), .A2(n3962), .ZN(n2559) );
  NAND4_X1 U32250 ( .A1(n2562), .A2(n2561), .A3(n2560), .A4(n2559), .ZN(n3970)
         );
  NAND2_X1 U32260 ( .A1(n3970), .A2(n2644), .ZN(n2567) );
  OR2_X1 U32270 ( .A1(n2563), .A2(n2152), .ZN(n2564) );
  MUX2_X1 U32280 ( .A(n3616), .B(DATAI_15_), .S(n2363), .Z(n4285) );
  NAND2_X1 U32290 ( .A1(n4285), .A2(n2645), .ZN(n2566) );
  NAND2_X1 U32300 ( .A1(n2567), .A2(n2566), .ZN(n2568) );
  XNOR2_X1 U32310 ( .A(n2568), .B(n2722), .ZN(n2569) );
  AOI22_X1 U32320 ( .A1(n3970), .A2(n2697), .B1(n2644), .B2(n4285), .ZN(n4287)
         );
  XNOR2_X1 U32330 ( .A(n2572), .B(n2571), .ZN(n3345) );
  NAND2_X1 U32340 ( .A1(n2353), .A2(REG0_REG_17__SCAN_IN), .ZN(n2581) );
  NAND2_X1 U32350 ( .A1(n2043), .A2(REG1_REG_17__SCAN_IN), .ZN(n2580) );
  INV_X1 U32360 ( .A(n2574), .ZN(n2573) );
  INV_X1 U32370 ( .A(n2592), .ZN(n2577) );
  INV_X1 U32380 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2575) );
  NAND2_X1 U32390 ( .A1(n2575), .A2(n2574), .ZN(n2576) );
  NAND2_X1 U32400 ( .A1(n2577), .A2(n2576), .ZN(n3917) );
  OR2_X1 U32410 ( .A1(n2040), .A2(n3917), .ZN(n2579) );
  INV_X1 U32420 ( .A(REG2_REG_17__SCAN_IN), .ZN(n3918) );
  OR2_X1 U32430 ( .A1(n2356), .A2(n3918), .ZN(n2578) );
  NAND4_X1 U32440 ( .A1(n2581), .A2(n2580), .A3(n2579), .A4(n2578), .ZN(n3926)
         );
  NAND2_X1 U32450 ( .A1(n3926), .A2(n2038), .ZN(n2585) );
  NAND2_X1 U32460 ( .A1(n2582), .A2(IR_REG_31__SCAN_IN), .ZN(n2583) );
  XNOR2_X1 U32470 ( .A(n2583), .B(IR_REG_17__SCAN_IN), .ZN(n4531) );
  MUX2_X1 U32480 ( .A(n4531), .B(DATAI_17_), .S(n2363), .Z(n3642) );
  NAND2_X1 U32490 ( .A1(n3642), .A2(n2645), .ZN(n2584) );
  NAND2_X1 U32500 ( .A1(n2585), .A2(n2584), .ZN(n2586) );
  XNOR2_X1 U32510 ( .A(n2586), .B(n2783), .ZN(n3353) );
  NAND2_X1 U32520 ( .A1(n3926), .A2(n2697), .ZN(n2588) );
  NAND2_X1 U32530 ( .A1(n3642), .A2(n2644), .ZN(n2587) );
  NAND2_X1 U32540 ( .A1(n3353), .A2(n3352), .ZN(n2591) );
  INV_X1 U32550 ( .A(n3353), .ZN(n2590) );
  INV_X1 U32560 ( .A(n3352), .ZN(n2589) );
  NAND2_X1 U32570 ( .A1(n2353), .A2(REG0_REG_18__SCAN_IN), .ZN(n2596) );
  NAND2_X1 U32580 ( .A1(n2042), .A2(REG1_REG_18__SCAN_IN), .ZN(n2595) );
  OAI21_X1 U32590 ( .B1(n2592), .B2(REG3_REG_18__SCAN_IN), .A(n2624), .ZN(
        n3898) );
  OR2_X1 U32600 ( .A1(n2039), .A2(n3898), .ZN(n2594) );
  INV_X1 U32610 ( .A(REG2_REG_18__SCAN_IN), .ZN(n3899) );
  OR2_X1 U32620 ( .A1(n2356), .A2(n3899), .ZN(n2593) );
  NAND4_X1 U32630 ( .A1(n2596), .A2(n2595), .A3(n2594), .A4(n2593), .ZN(n3909)
         );
  NAND2_X1 U32640 ( .A1(n3909), .A2(n2038), .ZN(n2601) );
  OR2_X1 U32650 ( .A1(n2598), .A2(n2597), .ZN(n2599) );
  XNOR2_X1 U32660 ( .A(n2599), .B(IR_REG_18__SCAN_IN), .ZN(n3620) );
  MUX2_X1 U32670 ( .A(n3620), .B(DATAI_18_), .S(n2363), .Z(n3896) );
  NAND2_X1 U32680 ( .A1(n3896), .A2(n2645), .ZN(n2600) );
  NAND2_X1 U32690 ( .A1(n2601), .A2(n2600), .ZN(n2602) );
  XNOR2_X1 U32700 ( .A(n2602), .B(n2783), .ZN(n2606) );
  INV_X1 U32710 ( .A(n2606), .ZN(n2604) );
  AOI22_X1 U32720 ( .A1(n3909), .A2(n2697), .B1(n2038), .B2(n3896), .ZN(n2605)
         );
  INV_X1 U32730 ( .A(n2605), .ZN(n2603) );
  NAND2_X1 U32740 ( .A1(n2604), .A2(n2603), .ZN(n3391) );
  AND2_X1 U32750 ( .A1(n2606), .A2(n2605), .ZN(n3392) );
  NAND2_X1 U32760 ( .A1(n2353), .A2(REG0_REG_19__SCAN_IN), .ZN(n2612) );
  NAND2_X1 U32770 ( .A1(n2042), .A2(REG1_REG_19__SCAN_IN), .ZN(n2611) );
  INV_X1 U32780 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2607) );
  XNOR2_X1 U32790 ( .A(n2624), .B(n2607), .ZN(n3321) );
  OR2_X1 U32800 ( .A1(n2039), .A2(n3321), .ZN(n2610) );
  INV_X1 U32810 ( .A(REG2_REG_19__SCAN_IN), .ZN(n2608) );
  OR2_X1 U32820 ( .A1(n2832), .A2(n2608), .ZN(n2609) );
  NAND4_X1 U32830 ( .A1(n2612), .A2(n2611), .A3(n2610), .A4(n2609), .ZN(n3891)
         );
  NAND2_X1 U32840 ( .A1(n3891), .A2(n2038), .ZN(n2615) );
  INV_X1 U32850 ( .A(DATAI_19_), .ZN(n2613) );
  MUX2_X1 U32860 ( .A(n3624), .B(n2613), .S(n2363), .Z(n3644) );
  OR2_X1 U32870 ( .A1(n3644), .A2(n2692), .ZN(n2614) );
  NAND2_X1 U32880 ( .A1(n2615), .A2(n2614), .ZN(n2616) );
  XNOR2_X1 U32890 ( .A(n2616), .B(n2722), .ZN(n2617) );
  OAI22_X1 U32900 ( .A1(n3858), .A2(n2658), .B1(n2080), .B2(n3644), .ZN(n2618)
         );
  XNOR2_X1 U32910 ( .A(n2617), .B(n2618), .ZN(n3320) );
  NAND2_X1 U32920 ( .A1(n2353), .A2(REG0_REG_20__SCAN_IN), .ZN(n2630) );
  NAND2_X1 U32930 ( .A1(n2043), .A2(REG1_REG_20__SCAN_IN), .ZN(n2629) );
  INV_X1 U32940 ( .A(n2624), .ZN(n2622) );
  AOI21_X1 U32950 ( .B1(n2622), .B2(REG3_REG_19__SCAN_IN), .A(
        REG3_REG_20__SCAN_IN), .ZN(n2625) );
  NAND2_X1 U32960 ( .A1(REG3_REG_19__SCAN_IN), .A2(REG3_REG_20__SCAN_IN), .ZN(
        n2623) );
  OR2_X1 U32970 ( .A1(n2625), .A2(n2637), .ZN(n3376) );
  OR2_X1 U32980 ( .A1(n2040), .A2(n3376), .ZN(n2628) );
  INV_X1 U32990 ( .A(REG2_REG_20__SCAN_IN), .ZN(n2626) );
  OR2_X1 U33000 ( .A1(n2832), .A2(n2626), .ZN(n2627) );
  NAND4_X1 U33010 ( .A1(n2630), .A2(n2629), .A3(n2628), .A4(n2627), .ZN(n3878)
         );
  NAND2_X1 U33020 ( .A1(n3878), .A2(n2644), .ZN(n2632) );
  NAND2_X1 U33030 ( .A1(n2363), .A2(DATAI_20_), .ZN(n3861) );
  OR2_X1 U33040 ( .A1(n3861), .A2(n2692), .ZN(n2631) );
  NAND2_X1 U33050 ( .A1(n2632), .A2(n2631), .ZN(n2633) );
  XNOR2_X1 U33060 ( .A(n2633), .B(n2783), .ZN(n2636) );
  NOR2_X1 U33070 ( .A1(n3861), .A2(n2080), .ZN(n2634) );
  AOI21_X1 U33080 ( .B1(n3878), .B2(n2697), .A(n2634), .ZN(n2635) );
  OR2_X1 U33090 ( .A1(n2636), .A2(n2635), .ZN(n3372) );
  NAND2_X1 U33100 ( .A1(n2636), .A2(n2635), .ZN(n3374) );
  NAND2_X1 U33110 ( .A1(n2353), .A2(REG0_REG_21__SCAN_IN), .ZN(n2643) );
  NAND2_X1 U33120 ( .A1(n2043), .A2(REG1_REG_21__SCAN_IN), .ZN(n2642) );
  NAND2_X1 U33130 ( .A1(n2637), .A2(REG3_REG_21__SCAN_IN), .ZN(n2661) );
  OR2_X1 U33140 ( .A1(n2637), .A2(REG3_REG_21__SCAN_IN), .ZN(n2638) );
  NAND2_X1 U33150 ( .A1(n2661), .A2(n2638), .ZN(n3330) );
  OR2_X1 U33160 ( .A1(n2040), .A2(n3330), .ZN(n2641) );
  INV_X1 U33170 ( .A(REG2_REG_21__SCAN_IN), .ZN(n2639) );
  OR2_X1 U33180 ( .A1(n2356), .A2(n2639), .ZN(n2640) );
  NAND2_X1 U33190 ( .A1(n3855), .A2(n2038), .ZN(n2647) );
  NAND2_X1 U33200 ( .A1(n3835), .A2(n2645), .ZN(n2646) );
  NAND2_X1 U33210 ( .A1(n2647), .A2(n2646), .ZN(n2648) );
  XNOR2_X1 U33220 ( .A(n2648), .B(n2722), .ZN(n3328) );
  NAND2_X1 U33230 ( .A1(n3855), .A2(n2697), .ZN(n2650) );
  NAND2_X1 U33240 ( .A1(n3835), .A2(n2038), .ZN(n2649) );
  NAND2_X1 U33250 ( .A1(n2650), .A2(n2649), .ZN(n3327) );
  NOR2_X1 U33260 ( .A1(n3328), .A2(n3327), .ZN(n2651) );
  NAND2_X1 U33270 ( .A1(n2353), .A2(REG0_REG_22__SCAN_IN), .ZN(n2656) );
  NAND2_X1 U33280 ( .A1(n2042), .A2(REG1_REG_22__SCAN_IN), .ZN(n2655) );
  INV_X1 U33290 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3386) );
  XNOR2_X1 U33300 ( .A(n2661), .B(n3386), .ZN(n3385) );
  OR2_X1 U33310 ( .A1(n2040), .A2(n3385), .ZN(n2654) );
  INV_X1 U33320 ( .A(REG2_REG_22__SCAN_IN), .ZN(n2652) );
  OR2_X1 U33330 ( .A1(n2832), .A2(n2652), .ZN(n2653) );
  NAND4_X1 U33340 ( .A1(n2656), .A2(n2655), .A3(n2654), .A4(n2653), .ZN(n3836)
         );
  INV_X1 U33350 ( .A(n3824), .ZN(n3471) );
  OAI22_X1 U33360 ( .A1(n3468), .A2(n2080), .B1(n2692), .B2(n3471), .ZN(n2657)
         );
  XNOR2_X1 U33370 ( .A(n2657), .B(n2722), .ZN(n2660) );
  OAI22_X1 U33380 ( .A1(n3468), .A2(n2658), .B1(n2080), .B2(n3471), .ZN(n2659)
         );
  XNOR2_X1 U33390 ( .A(n2660), .B(n2659), .ZN(n3384) );
  NOR2_X1 U33400 ( .A1(n2660), .A2(n2659), .ZN(n3311) );
  NAND2_X1 U33410 ( .A1(n2353), .A2(REG0_REG_23__SCAN_IN), .ZN(n2666) );
  NAND2_X1 U33420 ( .A1(n2042), .A2(REG1_REG_23__SCAN_IN), .ZN(n2665) );
  INV_X1 U33430 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3314) );
  OAI21_X1 U33440 ( .B1(n2661), .B2(n3386), .A(n3314), .ZN(n2662) );
  NAND2_X1 U33450 ( .A1(n2662), .A2(n2673), .ZN(n3798) );
  OR2_X1 U33460 ( .A1(n2039), .A2(n3798), .ZN(n2664) );
  INV_X1 U33470 ( .A(REG2_REG_23__SCAN_IN), .ZN(n3799) );
  OR2_X1 U33480 ( .A1(n2356), .A2(n3799), .ZN(n2663) );
  NAND4_X1 U33490 ( .A1(n2666), .A2(n2665), .A3(n2664), .A4(n2663), .ZN(n3780)
         );
  NAND2_X1 U33500 ( .A1(n3780), .A2(n2644), .ZN(n2668) );
  NAND2_X1 U33510 ( .A1(n2363), .A2(DATAI_23_), .ZN(n3809) );
  OR2_X1 U33520 ( .A1(n3809), .A2(n2692), .ZN(n2667) );
  NAND2_X1 U3353 ( .A1(n2668), .A2(n2667), .ZN(n2669) );
  XNOR2_X1 U33540 ( .A(n2669), .B(n2783), .ZN(n2672) );
  NOR2_X1 U3355 ( .A1(n3809), .A2(n2080), .ZN(n2670) );
  AOI21_X1 U3356 ( .B1(n3780), .B2(n2697), .A(n2670), .ZN(n2671) );
  XNOR2_X1 U3357 ( .A(n2672), .B(n2671), .ZN(n3310) );
  NOR2_X1 U3358 ( .A1(n2672), .A2(n2671), .ZN(n2684) );
  NAND2_X1 U3359 ( .A1(n2353), .A2(REG0_REG_24__SCAN_IN), .ZN(n2679) );
  NAND2_X1 U3360 ( .A1(n2042), .A2(REG1_REG_24__SCAN_IN), .ZN(n2678) );
  INV_X1 U3361 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4037) );
  AND2_X1 U3362 ( .A1(n2673), .A2(n4037), .ZN(n2674) );
  OR2_X1 U3363 ( .A1(n2674), .A2(n2686), .ZN(n3365) );
  OR2_X1 U3364 ( .A1(n2039), .A2(n3365), .ZN(n2677) );
  INV_X1 U3365 ( .A(REG2_REG_24__SCAN_IN), .ZN(n2675) );
  OR2_X1 U3366 ( .A1(n2832), .A2(n2675), .ZN(n2676) );
  NAND4_X1 U3367 ( .A1(n2679), .A2(n2678), .A3(n2677), .A4(n2676), .ZN(n3806)
         );
  NAND2_X1 U3368 ( .A1(n3806), .A2(n2697), .ZN(n2681) );
  NAND2_X1 U3369 ( .A1(n3779), .A2(n2038), .ZN(n2680) );
  NAND2_X1 U3370 ( .A1(n2681), .A2(n2680), .ZN(n2683) );
  NOR3_X2 U3371 ( .A1(n3309), .A2(n2684), .A3(n2683), .ZN(n3360) );
  OAI22_X1 U3372 ( .A1(n3765), .A2(n2080), .B1(n2692), .B2(n3786), .ZN(n2682)
         );
  XOR2_X1 U3373 ( .A(n2722), .B(n2682), .Z(n3363) );
  OAI21_X1 U3374 ( .B1(n3309), .B2(n2684), .A(n2683), .ZN(n3361) );
  NAND2_X1 U3375 ( .A1(n2042), .A2(REG1_REG_25__SCAN_IN), .ZN(n2691) );
  NAND2_X1 U3376 ( .A1(n2353), .A2(REG0_REG_25__SCAN_IN), .ZN(n2690) );
  INV_X1 U3377 ( .A(REG2_REG_25__SCAN_IN), .ZN(n2685) );
  OR2_X1 U3378 ( .A1(n2832), .A2(n2685), .ZN(n2689) );
  NOR2_X1 U3379 ( .A1(n2686), .A2(REG3_REG_25__SCAN_IN), .ZN(n2687) );
  OR2_X1 U3380 ( .A1(n2700), .A2(n2687), .ZN(n3339) );
  OR2_X1 U3381 ( .A1(n2039), .A2(n3339), .ZN(n2688) );
  NAND4_X1 U3382 ( .A1(n2691), .A2(n2690), .A3(n2689), .A4(n2688), .ZN(n3737)
         );
  NAND2_X1 U3383 ( .A1(n3737), .A2(n2038), .ZN(n2694) );
  NAND2_X1 U3384 ( .A1(n2363), .A2(DATAI_25_), .ZN(n3767) );
  OR2_X1 U3385 ( .A1(n3767), .A2(n2692), .ZN(n2693) );
  NAND2_X1 U3386 ( .A1(n2694), .A2(n2693), .ZN(n2695) );
  XNOR2_X1 U3387 ( .A(n2695), .B(n2783), .ZN(n2699) );
  NOR2_X1 U3388 ( .A1(n3767), .A2(n2080), .ZN(n2696) );
  AOI21_X1 U3389 ( .B1(n3737), .B2(n2697), .A(n2696), .ZN(n2698) );
  NAND2_X1 U3390 ( .A1(n2699), .A2(n2698), .ZN(n3335) );
  NOR2_X1 U3391 ( .A1(n2699), .A2(n2698), .ZN(n3336) );
  NAND2_X1 U3392 ( .A1(n2353), .A2(REG0_REG_26__SCAN_IN), .ZN(n2705) );
  NAND2_X1 U3393 ( .A1(n2043), .A2(REG1_REG_26__SCAN_IN), .ZN(n2704) );
  NOR2_X1 U3394 ( .A1(n2700), .A2(REG3_REG_26__SCAN_IN), .ZN(n2701) );
  OR2_X1 U3395 ( .A1(n2040), .A2(n3748), .ZN(n2703) );
  INV_X1 U3396 ( .A(REG2_REG_26__SCAN_IN), .ZN(n3749) );
  OR2_X1 U3397 ( .A1(n2356), .A2(n3749), .ZN(n2702) );
  NAND2_X1 U3398 ( .A1(n3762), .A2(n2038), .ZN(n2707) );
  NAND2_X1 U3399 ( .A1(n2363), .A2(DATAI_26_), .ZN(n3746) );
  OR2_X1 U3400 ( .A1(n3746), .A2(n2692), .ZN(n2706) );
  NAND2_X1 U3401 ( .A1(n2707), .A2(n2706), .ZN(n2708) );
  XNOR2_X1 U3402 ( .A(n2708), .B(n2783), .ZN(n2713) );
  INV_X1 U3403 ( .A(n2713), .ZN(n2711) );
  NOR2_X1 U3404 ( .A1(n3746), .A2(n2080), .ZN(n2709) );
  AOI21_X1 U3405 ( .B1(n3762), .B2(n2697), .A(n2709), .ZN(n2712) );
  INV_X1 U3406 ( .A(n2712), .ZN(n2710) );
  NAND2_X1 U3407 ( .A1(n2711), .A2(n2710), .ZN(n3401) );
  AND2_X1 U3408 ( .A1(n2713), .A2(n2712), .ZN(n3400) );
  NAND2_X1 U3409 ( .A1(n2353), .A2(REG0_REG_27__SCAN_IN), .ZN(n2719) );
  NAND2_X1 U3410 ( .A1(n2043), .A2(REG1_REG_27__SCAN_IN), .ZN(n2718) );
  NAND2_X1 U3411 ( .A1(n2714), .A2(REG3_REG_27__SCAN_IN), .ZN(n2762) );
  OR2_X1 U3412 ( .A1(n2714), .A2(REG3_REG_27__SCAN_IN), .ZN(n2715) );
  NAND2_X1 U3413 ( .A1(n2762), .A2(n2715), .ZN(n3720) );
  OR2_X1 U3414 ( .A1(n2039), .A2(n3720), .ZN(n2717) );
  INV_X1 U3415 ( .A(REG2_REG_27__SCAN_IN), .ZN(n3721) );
  OR2_X1 U3416 ( .A1(n2832), .A2(n3721), .ZN(n2716) );
  NAND4_X1 U3417 ( .A1(n2719), .A2(n2718), .A3(n2717), .A4(n2716), .ZN(n3738)
         );
  NAND2_X1 U3418 ( .A1(n3738), .A2(n2644), .ZN(n2721) );
  NAND2_X1 U3419 ( .A1(n3727), .A2(n2645), .ZN(n2720) );
  NAND2_X1 U3420 ( .A1(n2721), .A2(n2720), .ZN(n2723) );
  XNOR2_X1 U3421 ( .A(n2723), .B(n2722), .ZN(n2790) );
  AND2_X1 U3422 ( .A1(n3727), .A2(n2644), .ZN(n2724) );
  AOI21_X1 U3423 ( .B1(n3738), .B2(n2697), .A(n2724), .ZN(n2788) );
  XNOR2_X1 U3424 ( .A(n2790), .B(n2788), .ZN(n2779) );
  XNOR2_X1 U3425 ( .A(n2780), .B(n2779), .ZN(n2778) );
  NAND2_X1 U3426 ( .A1(n2725), .A2(n2742), .ZN(n2726) );
  MUX2_X1 U3427 ( .A(n2725), .B(n2726), .S(B_REG_SCAN_IN), .Z(n2727) );
  INV_X1 U3428 ( .A(n2814), .ZN(n2728) );
  INV_X1 U3429 ( .A(D_REG_0__SCAN_IN), .ZN(n2817) );
  NAND2_X1 U3430 ( .A1(n2728), .A2(n2817), .ZN(n2731) );
  INV_X1 U3431 ( .A(n4266), .ZN(n2729) );
  NAND2_X1 U3432 ( .A1(n2729), .A2(n2725), .ZN(n2730) );
  NOR4_X1 U3433 ( .A1(D_REG_9__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_28__SCAN_IN), .ZN(n2740) );
  NOR4_X1 U3434 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_2__SCAN_IN), .A3(
        D_REG_3__SCAN_IN), .A4(D_REG_4__SCAN_IN), .ZN(n2739) );
  INV_X1 U3435 ( .A(D_REG_12__SCAN_IN), .ZN(n4522) );
  INV_X1 U3436 ( .A(D_REG_16__SCAN_IN), .ZN(n4520) );
  INV_X1 U3437 ( .A(D_REG_21__SCAN_IN), .ZN(n4517) );
  INV_X1 U3438 ( .A(D_REG_18__SCAN_IN), .ZN(n4519) );
  NAND4_X1 U3439 ( .A1(n4522), .A2(n4520), .A3(n4517), .A4(n4519), .ZN(n2737)
         );
  NOR4_X1 U3440 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2735) );
  NOR4_X1 U3441 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_5__SCAN_IN), .A3(
        D_REG_6__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2734) );
  NOR4_X1 U3442 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2733) );
  NOR4_X1 U3443 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_22__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2732) );
  NAND4_X1 U3444 ( .A1(n2735), .A2(n2734), .A3(n2733), .A4(n2732), .ZN(n2736)
         );
  NOR4_X1 U3445 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(n2737), 
        .A4(n2736), .ZN(n2738) );
  AND3_X1 U3446 ( .A1(n2740), .A2(n2739), .A3(n2738), .ZN(n2741) );
  NOR2_X1 U3447 ( .A1(n2814), .A2(n2741), .ZN(n3077) );
  INV_X1 U3448 ( .A(n2742), .ZN(n4267) );
  OAI22_X1 U3449 ( .A1(n2814), .A2(D_REG_1__SCAN_IN), .B1(n4266), .B2(n4267), 
        .ZN(n3078) );
  NOR2_X1 U3450 ( .A1(n3077), .A2(n3078), .ZN(n2743) );
  NAND2_X1 U3451 ( .A1(n3080), .A2(n2743), .ZN(n2770) );
  INV_X1 U3452 ( .A(n2770), .ZN(n2751) );
  INV_X1 U3453 ( .A(n2938), .ZN(n2748) );
  NAND2_X1 U3454 ( .A1(n2752), .A2(n3624), .ZN(n2754) );
  NAND2_X1 U3455 ( .A1(n2769), .A2(n2754), .ZN(n2747) );
  NAND2_X1 U3456 ( .A1(n2748), .A2(n2747), .ZN(n2749) );
  NOR2_X1 U3457 ( .A1(n2855), .A2(n2749), .ZN(n2750) );
  INV_X1 U34580 ( .A(n3720), .ZN(n2776) );
  INV_X1 U34590 ( .A(n3624), .ZN(n4272) );
  AND2_X1 U3460 ( .A1(n2752), .A2(n4272), .ZN(n4509) );
  NOR2_X1 U3461 ( .A1(n4596), .A2(n4270), .ZN(n3074) );
  INV_X1 U3462 ( .A(n3074), .ZN(n2771) );
  NAND2_X1 U3463 ( .A1(n2770), .A2(n2771), .ZN(n2857) );
  AND2_X1 U3464 ( .A1(n2938), .A2(n2754), .ZN(n2854) );
  INV_X1 U3465 ( .A(n2854), .ZN(n2755) );
  NAND4_X1 U3466 ( .A1(n2857), .A2(n2821), .A3(n2305), .A4(n2755), .ZN(n2756)
         );
  INV_X1 U34670 ( .A(n2757), .ZN(n2758) );
  NAND3_X1 U3468 ( .A1(n2038), .A2(n2759), .A3(n2758), .ZN(n3569) );
  NOR2_X1 U34690 ( .A1(n2770), .A2(n3569), .ZN(n2761) );
  XNOR2_X1 U3470 ( .A(n2760), .B(IR_REG_28__SCAN_IN), .ZN(n2939) );
  INV_X1 U34710 ( .A(n2939), .ZN(n4264) );
  NAND2_X2 U3472 ( .A1(n2761), .A2(n4264), .ZN(n4280) );
  NAND2_X2 U34730 ( .A1(n2761), .A2(n2939), .ZN(n4281) );
  NAND2_X1 U3474 ( .A1(n2353), .A2(REG0_REG_28__SCAN_IN), .ZN(n2768) );
  NAND2_X1 U34750 ( .A1(n2043), .A2(REG1_REG_28__SCAN_IN), .ZN(n2767) );
  INV_X1 U3476 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2801) );
  OR2_X1 U34770 ( .A1(n2762), .A2(n2801), .ZN(n3692) );
  NAND2_X1 U3478 ( .A1(n2762), .A2(n2801), .ZN(n2763) );
  NAND2_X1 U34790 ( .A1(n3692), .A2(n2763), .ZN(n2796) );
  OR2_X1 U3480 ( .A1(n2039), .A2(n2796), .ZN(n2766) );
  INV_X1 U34810 ( .A(REG2_REG_28__SCAN_IN), .ZN(n2764) );
  OR2_X1 U3482 ( .A1(n2832), .A2(n2764), .ZN(n2765) );
  NAND4_X1 U34830 ( .A1(n2768), .A2(n2767), .A3(n2766), .A4(n2765), .ZN(n3728)
         );
  INV_X1 U3484 ( .A(n3728), .ZN(n3689) );
  OAI22_X1 U34850 ( .A1(n3731), .A2(n4280), .B1(n4281), .B2(n3689), .ZN(n2775)
         );
  NOR3_X1 U3486 ( .A1(n2770), .A2(n2855), .A3(n3930), .ZN(n2772) );
  NOR2_X2 U34870 ( .A1(n2772), .A2(n4491), .ZN(n3405) );
  INV_X1 U3488 ( .A(n3727), .ZN(n3660) );
  INV_X1 U34890 ( .A(REG3_REG_27__SCAN_IN), .ZN(n2773) );
  OAI22_X1 U3490 ( .A1(n3405), .A2(n3660), .B1(STATE_REG_SCAN_IN), .B2(n2773), 
        .ZN(n2774) );
  AOI211_X1 U34910 ( .C1(n2776), .C2(n3408), .A(n2775), .B(n2774), .ZN(n2777)
         );
  OAI21_X1 U3492 ( .B1(n2778), .B2(n3411), .A(n2777), .ZN(U3211) );
  NAND2_X1 U34930 ( .A1(n3728), .A2(n2644), .ZN(n2782) );
  AND2_X1 U3494 ( .A1(n2363), .A2(DATAI_28_), .ZN(n3704) );
  NAND2_X1 U34950 ( .A1(n3704), .A2(n2645), .ZN(n2781) );
  NAND2_X1 U3496 ( .A1(n2782), .A2(n2781), .ZN(n2784) );
  XNOR2_X1 U34970 ( .A(n2784), .B(n2783), .ZN(n2786) );
  AOI22_X1 U3498 ( .A1(n3728), .A2(n2697), .B1(n2038), .B2(n3704), .ZN(n2785)
         );
  XNOR2_X1 U34990 ( .A(n2786), .B(n2785), .ZN(n2794) );
  NAND2_X1 U3500 ( .A1(n2794), .A2(n4290), .ZN(n2787) );
  INV_X1 U35010 ( .A(n2794), .ZN(n2791) );
  INV_X1 U3502 ( .A(n2788), .ZN(n2789) );
  NAND2_X1 U35030 ( .A1(n2790), .A2(n2789), .ZN(n2793) );
  NAND2_X1 U3504 ( .A1(n2792), .A2(n2069), .ZN(n2806) );
  INV_X1 U35050 ( .A(n2793), .ZN(n2795) );
  NAND3_X1 U35060 ( .A1(n2795), .A2(n4290), .A3(n2794), .ZN(n2805) );
  INV_X1 U35070 ( .A(n2796), .ZN(n3713) );
  NAND2_X1 U35080 ( .A1(n2043), .A2(REG1_REG_29__SCAN_IN), .ZN(n2800) );
  NAND2_X1 U35090 ( .A1(n2353), .A2(REG0_REG_29__SCAN_IN), .ZN(n2799) );
  OR2_X1 U35100 ( .A1(n2040), .A2(n3692), .ZN(n2798) );
  INV_X1 U35110 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3695) );
  OR2_X1 U35120 ( .A1(n2832), .A2(n3695), .ZN(n2797) );
  NAND4_X1 U35130 ( .A1(n2800), .A2(n2799), .A3(n2798), .A4(n2797), .ZN(n3705)
         );
  INV_X1 U35140 ( .A(n3705), .ZN(n3477) );
  OAI22_X1 U35150 ( .A1(n3708), .A2(n4280), .B1(n4281), .B2(n3477), .ZN(n2803)
         );
  INV_X1 U35160 ( .A(n3704), .ZN(n3712) );
  OAI22_X1 U35170 ( .A1(n3405), .A2(n3712), .B1(STATE_REG_SCAN_IN), .B2(n2801), 
        .ZN(n2802) );
  AOI211_X1 U35180 ( .C1(n3408), .C2(n3713), .A(n2803), .B(n2802), .ZN(n2804)
         );
  NAND3_X1 U35190 ( .A1(n2807), .A2(n2806), .A3(n2237), .ZN(U3217) );
  OR2_X2 U35200 ( .A1(n2305), .A2(n4527), .ZN(n3583) );
  INV_X2 U35210 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND3_X1 U35220 ( .A1(n2808), .A2(STATE_REG_SCAN_IN), .A3(IR_REG_31__SCAN_IN), .ZN(n2810) );
  INV_X1 U35230 ( .A(DATAI_31_), .ZN(n2809) );
  OAI22_X1 U35240 ( .A1(n2811), .A2(n2810), .B1(STATE_REG_SCAN_IN), .B2(n2809), 
        .ZN(U3321) );
  INV_X1 U35250 ( .A(DATAI_29_), .ZN(n4040) );
  NAND2_X1 U35260 ( .A1(n2812), .A2(STATE_REG_SCAN_IN), .ZN(n2813) );
  OAI21_X1 U35270 ( .B1(STATE_REG_SCAN_IN), .B2(n4040), .A(n2813), .ZN(U3323)
         );
  INV_X1 U35280 ( .A(n2855), .ZN(n2815) );
  INV_X1 U35290 ( .A(n2725), .ZN(n4268) );
  NOR3_X1 U35300 ( .A1(n4268), .A2(n4266), .A3(n4527), .ZN(n2816) );
  AOI21_X1 U35310 ( .B1(n4526), .B2(n2817), .A(n2816), .ZN(U3458) );
  INV_X1 U35320 ( .A(D_REG_1__SCAN_IN), .ZN(n2819) );
  NOR3_X1 U35330 ( .A1(n4266), .A2(n4267), .A3(n4527), .ZN(n2818) );
  AOI21_X1 U35340 ( .B1(n4526), .B2(n2819), .A(n2818), .ZN(U3459) );
  NAND2_X1 U35350 ( .A1(n2821), .A2(n2938), .ZN(n2820) );
  AND2_X1 U35360 ( .A1(n2363), .A2(n2820), .ZN(n2838) );
  INV_X1 U35370 ( .A(n2838), .ZN(n2822) );
  OR2_X1 U35380 ( .A1(n2821), .A2(U3149), .ZN(n3572) );
  NAND2_X1 U35390 ( .A1(n2855), .A2(n3572), .ZN(n2837) );
  NOR2_X1 U35400 ( .A1(n4436), .A2(U4043), .ZN(U3148) );
  INV_X1 U35410 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n4080) );
  NAND2_X1 U35420 ( .A1(n3099), .A2(U4043), .ZN(n2823) );
  OAI21_X1 U35430 ( .B1(U4043), .B2(n4080), .A(n2823), .ZN(U3557) );
  INV_X1 U35440 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n2828) );
  INV_X1 U35450 ( .A(REG2_REG_30__SCAN_IN), .ZN(n2826) );
  NAND2_X1 U35460 ( .A1(n2042), .A2(REG1_REG_30__SCAN_IN), .ZN(n2825) );
  NAND2_X1 U35470 ( .A1(n2353), .A2(REG0_REG_30__SCAN_IN), .ZN(n2824) );
  OAI211_X1 U35480 ( .C1(n2832), .C2(n2826), .A(n2825), .B(n2824), .ZN(n3687)
         );
  NAND2_X1 U35490 ( .A1(n3687), .A2(U4043), .ZN(n2827) );
  OAI21_X1 U35500 ( .B1(U4043), .B2(n2828), .A(n2827), .ZN(U3580) );
  INV_X1 U35510 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n2834) );
  INV_X1 U35520 ( .A(REG2_REG_31__SCAN_IN), .ZN(n2831) );
  NAND2_X1 U35530 ( .A1(n2042), .A2(REG1_REG_31__SCAN_IN), .ZN(n2830) );
  NAND2_X1 U35540 ( .A1(n2353), .A2(REG0_REG_31__SCAN_IN), .ZN(n2829) );
  OAI211_X1 U35550 ( .C1(n2832), .C2(n2831), .A(n2830), .B(n2829), .ZN(n3556)
         );
  NAND2_X1 U35560 ( .A1(n3556), .A2(U4043), .ZN(n2833) );
  OAI21_X1 U35570 ( .B1(U4043), .B2(n2834), .A(n2833), .ZN(U3581) );
  INV_X1 U35580 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4611) );
  INV_X1 U35590 ( .A(REG1_REG_2__SCAN_IN), .ZN(n4609) );
  MUX2_X1 U35600 ( .A(REG1_REG_2__SCAN_IN), .B(n4609), .S(n4276), .Z(n2869) );
  INV_X1 U35610 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4607) );
  MUX2_X1 U35620 ( .A(REG1_REG_1__SCAN_IN), .B(n4607), .S(n4277), .Z(n3600) );
  AND2_X1 U35630 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3599) );
  NAND2_X1 U35640 ( .A1(n3600), .A2(n3599), .ZN(n3598) );
  NAND2_X1 U35650 ( .A1(n4277), .A2(REG1_REG_1__SCAN_IN), .ZN(n2835) );
  NAND2_X1 U35660 ( .A1(n3598), .A2(n2835), .ZN(n2868) );
  NAND2_X1 U35670 ( .A1(n2869), .A2(n2868), .ZN(n2867) );
  NAND2_X1 U35680 ( .A1(n4276), .A2(REG1_REG_2__SCAN_IN), .ZN(n2836) );
  NAND2_X1 U35690 ( .A1(n2867), .A2(n2836), .ZN(n2880) );
  XNOR2_X1 U35700 ( .A(n2880), .B(n4275), .ZN(n2839) );
  XNOR2_X1 U35710 ( .A(n2282), .B(IR_REG_27__SCAN_IN), .ZN(n4265) );
  INV_X1 U35720 ( .A(n4265), .ZN(n3585) );
  INV_X1 U35730 ( .A(n4438), .ZN(n4313) );
  AOI211_X1 U35740 ( .C1(n4611), .C2(n2839), .A(n2882), .B(n4313), .ZN(n2851)
         );
  MUX2_X1 U35750 ( .A(REG2_REG_2__SCAN_IN), .B(n2840), .S(n4276), .Z(n2844) );
  AND2_X1 U35760 ( .A1(REG2_REG_0__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2842) );
  NAND2_X1 U35770 ( .A1(n3596), .A2(n2842), .ZN(n3595) );
  NAND2_X1 U35780 ( .A1(n4277), .A2(REG2_REG_1__SCAN_IN), .ZN(n2870) );
  NAND2_X1 U35790 ( .A1(n3595), .A2(n2870), .ZN(n2843) );
  NAND2_X1 U35800 ( .A1(n2844), .A2(n2843), .ZN(n2873) );
  NAND2_X1 U35810 ( .A1(n4276), .A2(REG2_REG_2__SCAN_IN), .ZN(n2845) );
  NAND2_X1 U3582 ( .A1(n2873), .A2(n2845), .ZN(n2886) );
  OR2_X1 U3583 ( .A1(n3585), .A2(n2939), .ZN(n3568) );
  INV_X1 U3584 ( .A(n3568), .ZN(n2846) );
  OAI211_X1 U3585 ( .C1(REG2_REG_3__SCAN_IN), .C2(n2847), .A(n4388), .B(n2887), 
        .ZN(n2849) );
  INV_X1 U3586 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2984) );
  NOR2_X1 U3587 ( .A1(STATE_REG_SCAN_IN), .A2(n2984), .ZN(n2908) );
  AOI21_X1 U3588 ( .B1(n4436), .B2(ADDR_REG_3__SCAN_IN), .A(n2908), .ZN(n2848)
         );
  OAI211_X1 U3589 ( .C1(n4443), .C2(n2165), .A(n2849), .B(n2848), .ZN(n2850)
         );
  OR2_X1 U3590 ( .A1(n2851), .A2(n2850), .ZN(U3243) );
  XNOR2_X1 U3591 ( .A(n2853), .B(n2852), .ZN(n2860) );
  INV_X1 U3592 ( .A(n3075), .ZN(n2856) );
  NAND2_X1 U3593 ( .A1(n2857), .A2(n2856), .ZN(n3305) );
  AOI22_X1 U3594 ( .A1(n4284), .A2(n4492), .B1(REG3_REG_1__SCAN_IN), .B2(n3305), .ZN(n2859) );
  INV_X1 U3595 ( .A(n4280), .ZN(n3217) );
  INV_X1 U3596 ( .A(n4281), .ZN(n3218) );
  AOI22_X1 U3597 ( .A1(n3217), .A2(n3584), .B1(n3218), .B2(n4480), .ZN(n2858)
         );
  OAI211_X1 U3598 ( .C1(n2860), .C2(n3411), .A(n2859), .B(n2858), .ZN(U3219)
         );
  AND2_X1 U3599 ( .A1(n4265), .A2(n2861), .ZN(n2862) );
  OR2_X1 U3600 ( .A1(n2862), .A2(n2939), .ZN(n3587) );
  NAND2_X1 U3601 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3594) );
  OAI21_X1 U3602 ( .B1(n3568), .B2(n3594), .A(U4043), .ZN(n2866) );
  XOR2_X1 U3603 ( .A(n2864), .B(n2863), .Z(n3306) );
  NOR3_X1 U3604 ( .A1(n3306), .A2(n2939), .A3(n4265), .ZN(n2865) );
  AOI211_X1 U3605 ( .C1(n2158), .C2(n3587), .A(n2866), .B(n2865), .ZN(n2895)
         );
  AOI22_X1 U3606 ( .A1(n4436), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n2878) );
  OAI211_X1 U3607 ( .C1(n2869), .C2(n2868), .A(n4438), .B(n2867), .ZN(n2877)
         );
  MUX2_X1 U3608 ( .A(n2840), .B(REG2_REG_2__SCAN_IN), .S(n4276), .Z(n2871) );
  NAND3_X1 U3609 ( .A1(n2871), .A2(n3595), .A3(n2870), .ZN(n2872) );
  NAND3_X1 U3610 ( .A1(n4388), .A2(n2873), .A3(n2872), .ZN(n2876) );
  INV_X1 U3611 ( .A(n4276), .ZN(n2874) );
  OR2_X1 U3612 ( .A1(n4443), .A2(n2874), .ZN(n2875) );
  NAND4_X1 U3613 ( .A1(n2878), .A2(n2877), .A3(n2876), .A4(n2875), .ZN(n2879)
         );
  OR2_X1 U3614 ( .A1(n2895), .A2(n2879), .ZN(U3242) );
  AND2_X1 U3615 ( .A1(n2880), .A2(n4275), .ZN(n2881) );
  INV_X1 U3616 ( .A(n2883), .ZN(n2884) );
  INV_X1 U3617 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4613) );
  NAND2_X1 U3618 ( .A1(n2884), .A2(n4613), .ZN(n2885) );
  NAND3_X1 U3619 ( .A1(n4438), .A2(n3132), .A3(n2885), .ZN(n2893) );
  NAND2_X1 U3620 ( .A1(n2886), .A2(n4275), .ZN(n2888) );
  XNOR2_X1 U3621 ( .A(n3111), .B(n2355), .ZN(n2889) );
  NAND2_X1 U3622 ( .A1(n4388), .A2(n2889), .ZN(n2892) );
  AND2_X1 U3623 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n2919) );
  AOI21_X1 U3624 ( .B1(n4436), .B2(ADDR_REG_4__SCAN_IN), .A(n2919), .ZN(n2891)
         );
  OR2_X1 U3625 ( .A1(n4443), .A2(n3113), .ZN(n2890) );
  NAND4_X1 U3626 ( .A1(n2893), .A2(n2892), .A3(n2891), .A4(n2890), .ZN(n2894)
         );
  OR2_X1 U3627 ( .A1(n2895), .A2(n2894), .ZN(U3244) );
  INV_X1 U3628 ( .A(n2897), .ZN(n2898) );
  AOI21_X1 U3629 ( .B1(n2896), .B2(n2899), .A(n2898), .ZN(n2902) );
  AOI22_X1 U3630 ( .A1(n4284), .A2(n3058), .B1(REG3_REG_2__SCAN_IN), .B2(n3305), .ZN(n2901) );
  INV_X1 U3631 ( .A(n2304), .ZN(n4506) );
  AOI22_X1 U3632 ( .A1(n3218), .A2(n3582), .B1(n3217), .B2(n2304), .ZN(n2900)
         );
  OAI211_X1 U3633 ( .C1(n2902), .C2(n3411), .A(n2901), .B(n2900), .ZN(U3234)
         );
  NAND2_X1 U3634 ( .A1(n2905), .A2(n2903), .ZN(n2913) );
  OAI21_X1 U3635 ( .B1(n2903), .B2(n2905), .A(n2913), .ZN(n2906) );
  NAND2_X1 U3636 ( .A1(n2906), .A2(n4290), .ZN(n2910) );
  INV_X1 U3637 ( .A(n4480), .ZN(n2929) );
  INV_X1 U3638 ( .A(n3581), .ZN(n3020) );
  OAI22_X1 U3639 ( .A1(n2929), .A2(n4280), .B1(n4281), .B2(n3020), .ZN(n2907)
         );
  AOI211_X1 U3640 ( .C1(n3432), .C2(n4284), .A(n2908), .B(n2907), .ZN(n2909)
         );
  OAI211_X1 U3641 ( .C1(REG3_REG_3__SCAN_IN), .C2(n4295), .A(n2910), .B(n2909), 
        .ZN(U3215) );
  AND2_X1 U3642 ( .A1(n2913), .A2(n2911), .ZN(n2916) );
  NAND2_X1 U3643 ( .A1(n2913), .A2(n2912), .ZN(n2914) );
  OAI211_X1 U3644 ( .C1(n2916), .C2(n2915), .A(n4290), .B(n2914), .ZN(n2921)
         );
  INV_X1 U3645 ( .A(n3582), .ZN(n3431) );
  OAI22_X1 U3646 ( .A1(n3004), .A2(n4281), .B1(n4280), .B2(n3431), .ZN(n2918)
         );
  AOI211_X1 U3647 ( .C1(n2917), .C2(n4284), .A(n2919), .B(n2918), .ZN(n2920)
         );
  OAI211_X1 U3648 ( .C1(n4295), .C2(n2947), .A(n2921), .B(n2920), .ZN(U3227)
         );
  AND2_X1 U3649 ( .A1(n3584), .A2(n4493), .ZN(n4485) );
  NAND2_X1 U3650 ( .A1(n2304), .A2(n4492), .ZN(n2927) );
  INV_X1 U3651 ( .A(n3055), .ZN(n2928) );
  NAND2_X1 U3652 ( .A1(n2929), .A2(n3058), .ZN(n2934) );
  INV_X1 U3653 ( .A(n3058), .ZN(n3066) );
  NAND2_X1 U3654 ( .A1(n4480), .A2(n3066), .ZN(n3429) );
  NAND2_X1 U3655 ( .A1(n2928), .A2(n3061), .ZN(n3057) );
  NAND2_X1 U3656 ( .A1(n2929), .A2(n3066), .ZN(n2930) );
  NAND2_X1 U3657 ( .A1(n3057), .A2(n2930), .ZN(n2971) );
  NOR2_X1 U3658 ( .A1(n3582), .A2(n3432), .ZN(n2931) );
  INV_X1 U3659 ( .A(n3432), .ZN(n2977) );
  NAND2_X1 U3660 ( .A1(n3020), .A2(n2917), .ZN(n3434) );
  NAND2_X1 U3661 ( .A1(n3581), .A2(n2946), .ZN(n3437) );
  NAND2_X1 U3662 ( .A1(n3434), .A2(n3437), .ZN(n3002) );
  XNOR2_X1 U3663 ( .A(n3003), .B(n3002), .ZN(n2952) );
  XNOR2_X1 U3664 ( .A(n4269), .B(n2953), .ZN(n2932) );
  NAND2_X1 U3665 ( .A1(n2932), .A2(n3624), .ZN(n4487) );
  INV_X1 U3666 ( .A(n3584), .ZN(n4483) );
  NAND2_X1 U3667 ( .A1(n4483), .A2(n4493), .ZN(n3518) );
  NAND2_X1 U3668 ( .A1(n2933), .A2(n3519), .ZN(n3063) );
  NAND2_X1 U3669 ( .A1(n3063), .A2(n2934), .ZN(n2935) );
  XNOR2_X1 U3670 ( .A(n3582), .B(n3432), .ZN(n3523) );
  NAND2_X1 U3671 ( .A1(n3431), .A2(n3432), .ZN(n3433) );
  INV_X1 U3672 ( .A(n3002), .ZN(n3510) );
  XNOR2_X1 U3673 ( .A(n2998), .B(n3510), .ZN(n2942) );
  NAND2_X1 U3674 ( .A1(n4269), .A2(n4272), .ZN(n2937) );
  NAND2_X1 U3675 ( .A1(n4271), .A2(n4270), .ZN(n2936) );
  NAND2_X1 U3676 ( .A1(n2939), .A2(n2938), .ZN(n4505) );
  INV_X2 U3677 ( .A(n4505), .ZN(n4479) );
  AOI22_X1 U3678 ( .A1(n3580), .A2(n4479), .B1(n2917), .B2(n4478), .ZN(n2940)
         );
  OAI21_X1 U3679 ( .B1(n3431), .B2(n4482), .A(n2940), .ZN(n2941) );
  AOI21_X1 U3680 ( .B1(n2942), .B2(n4502), .A(n2941), .ZN(n2943) );
  OAI21_X1 U3681 ( .B1(n2952), .B2(n4487), .A(n2943), .ZN(n4575) );
  INV_X1 U3682 ( .A(n3026), .ZN(n2945) );
  OAI211_X1 U3683 ( .C1(n2983), .C2(n2946), .A(n2945), .B(n4602), .ZN(n4574)
         );
  OAI22_X1 U3684 ( .A1(n4574), .A2(n4272), .B1(n4515), .B2(n2947), .ZN(n2951)
         );
  INV_X1 U3685 ( .A(n3078), .ZN(n2949) );
  NOR2_X1 U3686 ( .A1(n3077), .A2(n3075), .ZN(n2948) );
  NAND3_X1 U3687 ( .A1(n3084), .A2(n2949), .A3(n2948), .ZN(n2950) );
  OAI21_X1 U3688 ( .B1(n4575), .B2(n2951), .A(n4511), .ZN(n2956) );
  INV_X1 U3689 ( .A(n2952), .ZN(n4578) );
  OR2_X1 U3690 ( .A1(n2953), .A2(n3624), .ZN(n2954) );
  AOI22_X1 U3691 ( .A1(n4578), .A2(n4501), .B1(REG2_REG_4__SCAN_IN), .B2(n4296), .ZN(n2955) );
  NAND2_X1 U3692 ( .A1(n2956), .A2(n2955), .ZN(U3286) );
  XOR2_X1 U3693 ( .A(n2957), .B(n2958), .Z(n2959) );
  NAND2_X1 U3694 ( .A1(n2959), .A2(n4290), .ZN(n2962) );
  AND2_X1 U3695 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n4306) );
  INV_X1 U3696 ( .A(n3579), .ZN(n3048) );
  OAI22_X1 U3697 ( .A1(n3020), .A2(n4280), .B1(n4281), .B2(n3048), .ZN(n2960)
         );
  AOI211_X1 U3698 ( .C1(n3018), .C2(n4284), .A(n4306), .B(n2960), .ZN(n2961)
         );
  OAI211_X1 U3699 ( .C1(n4295), .C2(n3027), .A(n2962), .B(n2961), .ZN(U3224)
         );
  NAND2_X1 U3700 ( .A1(n2964), .A2(n2963), .ZN(n2966) );
  XOR2_X1 U3701 ( .A(n2966), .B(n2965), .Z(n2967) );
  NAND2_X1 U3702 ( .A1(n2967), .A2(n4290), .ZN(n2970) );
  INV_X1 U3703 ( .A(REG3_REG_6__SCAN_IN), .ZN(n4110) );
  NOR2_X1 U3704 ( .A1(STATE_REG_SCAN_IN), .A2(n4110), .ZN(n4318) );
  INV_X1 U3705 ( .A(n3099), .ZN(n3185) );
  OAI22_X1 U3706 ( .A1(n3004), .A2(n4280), .B1(n4281), .B2(n3185), .ZN(n2968)
         );
  AOI211_X1 U3707 ( .C1(n3038), .C2(n4284), .A(n4318), .B(n2968), .ZN(n2969)
         );
  OAI211_X1 U3708 ( .C1(n4295), .C2(n3010), .A(n2970), .B(n2969), .ZN(U3236)
         );
  INV_X1 U3709 ( .A(n3523), .ZN(n2972) );
  XNOR2_X1 U3710 ( .A(n2971), .B(n2972), .ZN(n4570) );
  INV_X1 U3711 ( .A(n4487), .ZN(n4503) );
  NAND2_X1 U3712 ( .A1(n4570), .A2(n4503), .ZN(n2981) );
  NAND3_X1 U3713 ( .A1(n3063), .A2(n2934), .A3(n2972), .ZN(n2973) );
  NAND2_X1 U3714 ( .A1(n2974), .A2(n2973), .ZN(n2979) );
  INV_X1 U3715 ( .A(n4482), .ZN(n3925) );
  NAND2_X1 U3716 ( .A1(n4480), .A2(n3925), .ZN(n2976) );
  NAND2_X1 U3717 ( .A1(n3581), .A2(n4479), .ZN(n2975) );
  OAI211_X1 U3718 ( .C1(n3930), .C2(n2977), .A(n2976), .B(n2975), .ZN(n2978)
         );
  AOI21_X1 U3719 ( .B1(n2979), .B2(n4502), .A(n2978), .ZN(n2980) );
  AND2_X1 U3720 ( .A1(n2981), .A2(n2980), .ZN(n4572) );
  AND2_X1 U3721 ( .A1(n4564), .A2(n3432), .ZN(n2982) );
  NOR2_X1 U3722 ( .A1(n2983), .A2(n2982), .ZN(n4569) );
  INV_X1 U3723 ( .A(n4569), .ZN(n2986) );
  AOI22_X1 U3724 ( .A1(n4296), .A2(REG2_REG_3__SCAN_IN), .B1(n4491), .B2(n2984), .ZN(n2985) );
  OAI21_X1 U3725 ( .B1(n2986), .B2(n3961), .A(n2985), .ZN(n2987) );
  AOI21_X1 U3726 ( .B1(n4570), .B2(n4501), .A(n2987), .ZN(n2988) );
  OAI21_X1 U3727 ( .B1(n4572), .B2(n4296), .A(n2988), .ZN(U3287) );
  AOI21_X1 U3728 ( .B1(n2990), .B2(n2989), .A(n3411), .ZN(n2992) );
  NAND2_X1 U3729 ( .A1(n2992), .A2(n2991), .ZN(n2996) );
  NOR2_X1 U3730 ( .A1(STATE_REG_SCAN_IN), .A2(n2993), .ZN(n4327) );
  OAI22_X1 U3731 ( .A1(n3048), .A2(n4280), .B1(n4281), .B2(n2218), .ZN(n2994)
         );
  AOI211_X1 U3732 ( .C1(n3098), .C2(n4284), .A(n4327), .B(n2994), .ZN(n2995)
         );
  OAI211_X1 U3733 ( .C1(n4295), .C2(n3050), .A(n2996), .B(n2995), .ZN(U3210)
         );
  INV_X1 U3734 ( .A(n3434), .ZN(n2997) );
  AND2_X1 U3735 ( .A1(n3580), .A2(n3025), .ZN(n3016) );
  NAND2_X1 U3736 ( .A1(n3004), .A2(n3018), .ZN(n3445) );
  NAND2_X1 U3737 ( .A1(n3048), .A2(n3038), .ZN(n3439) );
  INV_X1 U3738 ( .A(n3038), .ZN(n3008) );
  NAND2_X1 U3739 ( .A1(n3579), .A2(n3008), .ZN(n3446) );
  AND2_X1 U3740 ( .A1(n3439), .A2(n3446), .ZN(n3514) );
  XNOR2_X1 U3741 ( .A(n3043), .B(n3514), .ZN(n2999) );
  NAND2_X1 U3742 ( .A1(n2999), .A2(n4502), .ZN(n3001) );
  AOI22_X1 U3743 ( .A1(n3099), .A2(n4479), .B1(n4478), .B2(n3038), .ZN(n3000)
         );
  OAI211_X1 U3744 ( .C1(n3004), .C2(n4482), .A(n3001), .B(n3000), .ZN(n3081)
         );
  INV_X1 U3745 ( .A(n3081), .ZN(n3015) );
  NAND2_X1 U3746 ( .A1(n3004), .A2(n3025), .ZN(n3005) );
  XOR2_X1 U3747 ( .A(n3514), .B(n3041), .Z(n3082) );
  OR2_X1 U3748 ( .A1(n4296), .A2(n4487), .ZN(n3006) );
  NAND2_X1 U3749 ( .A1(n3026), .A2(n3025), .ZN(n3024) );
  INV_X1 U3750 ( .A(n3024), .ZN(n3009) );
  OAI21_X1 U3751 ( .B1(n3009), .B2(n3008), .A(n3049), .ZN(n3089) );
  NOR2_X1 U3752 ( .A1(n3089), .A2(n3961), .ZN(n3013) );
  OAI22_X1 U3753 ( .A1(n4511), .A2(n3011), .B1(n3010), .B2(n4515), .ZN(n3012)
         );
  AOI211_X1 U3754 ( .C1(n3082), .C2(n3965), .A(n3013), .B(n3012), .ZN(n3014)
         );
  OAI21_X1 U3755 ( .B1(n4296), .B2(n3015), .A(n3014), .ZN(U3284) );
  INV_X1 U3756 ( .A(n3016), .ZN(n3436) );
  XOR2_X1 U3757 ( .A(n3509), .B(n3017), .Z(n3022) );
  AOI22_X1 U3758 ( .A1(n3579), .A2(n4479), .B1(n4478), .B2(n3018), .ZN(n3019)
         );
  OAI21_X1 U3759 ( .B1(n3020), .B2(n4482), .A(n3019), .ZN(n3021) );
  AOI21_X1 U3760 ( .B1(n3022), .B2(n4502), .A(n3021), .ZN(n4580) );
  XNOR2_X1 U3761 ( .A(n3023), .B(n3509), .ZN(n4583) );
  OAI21_X1 U3762 ( .B1(n3026), .B2(n3025), .A(n3024), .ZN(n4581) );
  NOR2_X1 U3763 ( .A1(n4581), .A2(n3961), .ZN(n3029) );
  INV_X1 U3764 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3116) );
  OAI22_X1 U3765 ( .A1(n4511), .A2(n3116), .B1(n3027), .B2(n4515), .ZN(n3028)
         );
  AOI211_X1 U3766 ( .C1(n4583), .C2(n3965), .A(n3029), .B(n3028), .ZN(n3030)
         );
  OAI21_X1 U3767 ( .B1(n4580), .B2(n4296), .A(n3030), .ZN(U3285) );
  XOR2_X1 U3768 ( .A(n3149), .B(n3032), .Z(n3033) );
  XNOR2_X1 U3769 ( .A(n3031), .B(n3033), .ZN(n3037) );
  AOI22_X1 U3770 ( .A1(n3217), .A2(n3099), .B1(n3218), .B2(n3577), .ZN(n3034)
         );
  NAND2_X1 U3771 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n4336) );
  OAI211_X1 U3772 ( .C1(n3405), .C2(n2217), .A(n3034), .B(n4336), .ZN(n3035)
         );
  AOI21_X1 U3773 ( .B1(n4468), .B2(n3408), .A(n3035), .ZN(n3036) );
  OAI21_X1 U3774 ( .B1(n3037), .B2(n3411), .A(n3036), .ZN(U3218) );
  NOR2_X1 U3775 ( .A1(n3579), .A2(n3038), .ZN(n3040) );
  NAND2_X1 U3776 ( .A1(n3579), .A2(n3038), .ZN(n3039) );
  NAND2_X1 U3777 ( .A1(n3185), .A2(n3098), .ZN(n3090) );
  INV_X1 U3778 ( .A(n3098), .ZN(n3042) );
  NAND2_X1 U3779 ( .A1(n3099), .A2(n3042), .ZN(n3448) );
  NAND2_X1 U3780 ( .A1(n3090), .A2(n3448), .ZN(n3096) );
  INV_X1 U3781 ( .A(n3096), .ZN(n3520) );
  XNOR2_X1 U3782 ( .A(n3097), .B(n3520), .ZN(n4587) );
  INV_X1 U3783 ( .A(n4587), .ZN(n3054) );
  NAND2_X1 U3784 ( .A1(n3043), .A2(n3446), .ZN(n3044) );
  XNOR2_X1 U3785 ( .A(n3092), .B(n3520), .ZN(n3045) );
  NAND2_X1 U3786 ( .A1(n3045), .A2(n4502), .ZN(n3047) );
  AOI22_X1 U3787 ( .A1(n3578), .A2(n4479), .B1(n4478), .B2(n3098), .ZN(n3046)
         );
  OAI211_X1 U3788 ( .C1(n3048), .C2(n4482), .A(n3047), .B(n3046), .ZN(n4585)
         );
  NAND2_X1 U3789 ( .A1(n4585), .A2(n4511), .ZN(n3053) );
  AOI211_X1 U3790 ( .C1(n3098), .C2(n3049), .A(n4591), .B(n3180), .ZN(n4586)
         );
  OAI22_X1 U3791 ( .A1(n4511), .A2(n2413), .B1(n3050), .B2(n4515), .ZN(n3051)
         );
  AOI21_X1 U3792 ( .B1(n4586), .B2(n3905), .A(n3051), .ZN(n3052) );
  OAI211_X1 U3793 ( .C1(n3054), .C2(n3902), .A(n3053), .B(n3052), .ZN(U3283)
         );
  NAND2_X1 U3794 ( .A1(n3055), .A2(n3519), .ZN(n3056) );
  NAND2_X1 U3795 ( .A1(n3057), .A2(n3056), .ZN(n4567) );
  NAND2_X1 U3796 ( .A1(n4495), .A2(n3058), .ZN(n4563) );
  NAND3_X1 U3797 ( .A1(n4498), .A2(n4564), .A3(n4563), .ZN(n3059) );
  OAI21_X1 U3798 ( .B1(n4515), .B2(n3060), .A(n3059), .ZN(n3072) );
  INV_X1 U3799 ( .A(n3519), .ZN(n3061) );
  NAND3_X1 U3800 ( .A1(n3061), .A2(n3427), .A3(n4475), .ZN(n3062) );
  NAND2_X1 U3801 ( .A1(n3063), .A2(n3062), .ZN(n3068) );
  NAND2_X1 U3802 ( .A1(n2304), .A2(n3925), .ZN(n3065) );
  NAND2_X1 U3803 ( .A1(n3582), .A2(n4479), .ZN(n3064) );
  OAI211_X1 U3804 ( .C1(n3930), .C2(n3066), .A(n3065), .B(n3064), .ZN(n3067)
         );
  AOI21_X1 U3805 ( .B1(n3068), .B2(n4502), .A(n3067), .ZN(n3070) );
  NAND2_X1 U3806 ( .A1(n4567), .A2(n4503), .ZN(n3069) );
  NAND2_X1 U3807 ( .A1(n3070), .A2(n3069), .ZN(n4565) );
  MUX2_X1 U3808 ( .A(n4565), .B(REG2_REG_2__SCAN_IN), .S(n4296), .Z(n3071) );
  AOI211_X1 U3809 ( .C1(n4501), .C2(n4567), .A(n3072), .B(n3071), .ZN(n3073)
         );
  INV_X1 U3810 ( .A(n3073), .ZN(U3288) );
  OR2_X1 U3811 ( .A1(n3075), .A2(n3074), .ZN(n3076) );
  NOR2_X1 U3812 ( .A1(n3077), .A2(n3076), .ZN(n3079) );
  INV_X1 U3813 ( .A(REG1_REG_6__SCAN_IN), .ZN(n4316) );
  AOI21_X1 U3814 ( .B1(n3082), .B2(n4594), .A(n3081), .ZN(n3086) );
  MUX2_X1 U3815 ( .A(n4316), .B(n3086), .S(n4624), .Z(n3083) );
  OAI21_X1 U3816 ( .B1(n3089), .B2(n4201), .A(n3083), .ZN(U3524) );
  INV_X1 U3817 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3087) );
  MUX2_X1 U3818 ( .A(n3087), .B(n3086), .S(n4605), .Z(n3088) );
  OAI21_X1 U3819 ( .B1(n3089), .B2(n4259), .A(n3088), .ZN(U3479) );
  INV_X1 U3820 ( .A(n3206), .ZN(n3103) );
  AND2_X1 U3821 ( .A1(n3577), .A2(n3103), .ZN(n3197) );
  INV_X1 U3822 ( .A(n3577), .ZN(n3271) );
  NAND2_X1 U3823 ( .A1(n3271), .A2(n3206), .ZN(n3443) );
  AND2_X1 U3824 ( .A1(n3198), .A2(n3443), .ZN(n3504) );
  INV_X1 U3825 ( .A(n3090), .ZN(n3091) );
  NAND2_X1 U3826 ( .A1(n2218), .A2(n3183), .ZN(n3442) );
  NAND2_X1 U3827 ( .A1(n3578), .A2(n2217), .ZN(n3447) );
  XOR2_X1 U3828 ( .A(n3504), .B(n3196), .Z(n3095) );
  AOI22_X1 U3829 ( .A1(n3576), .A2(n4479), .B1(n4478), .B2(n3206), .ZN(n3093)
         );
  OAI21_X1 U3830 ( .B1(n2218), .B2(n4482), .A(n3093), .ZN(n3094) );
  AOI21_X1 U3831 ( .B1(n3095), .B2(n4502), .A(n3094), .ZN(n4589) );
  NAND2_X1 U3832 ( .A1(n3097), .A2(n3096), .ZN(n3101) );
  NAND2_X1 U3833 ( .A1(n3099), .A2(n3098), .ZN(n3100) );
  NAND2_X1 U3834 ( .A1(n3101), .A2(n3100), .ZN(n3181) );
  AND2_X1 U3835 ( .A1(n3578), .A2(n3183), .ZN(n3102) );
  XOR2_X1 U3836 ( .A(n3504), .B(n3205), .Z(n4593) );
  OR2_X1 U3837 ( .A1(n3178), .A2(n3103), .ZN(n3104) );
  NAND2_X1 U3838 ( .A1(n3262), .A2(n3104), .ZN(n4590) );
  INV_X1 U3839 ( .A(n3105), .ZN(n3158) );
  AOI22_X1 U3840 ( .A1(n4296), .A2(REG2_REG_9__SCAN_IN), .B1(n3158), .B2(n4491), .ZN(n3106) );
  OAI21_X1 U3841 ( .B1(n4590), .B2(n3961), .A(n3106), .ZN(n3107) );
  AOI21_X1 U3842 ( .B1(n4593), .B2(n3965), .A(n3107), .ZN(n3108) );
  OAI21_X1 U3843 ( .B1(n4296), .B2(n4589), .A(n3108), .ZN(U3281) );
  INV_X1 U3844 ( .A(n4443), .ZN(n3593) );
  NAND2_X1 U3845 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n3299) );
  INV_X1 U3846 ( .A(n3299), .ZN(n3109) );
  AOI21_X1 U3847 ( .B1(n4436), .B2(ADDR_REG_14__SCAN_IN), .A(n3109), .ZN(n3110) );
  INV_X1 U3848 ( .A(n3110), .ZN(n3131) );
  INV_X1 U3849 ( .A(n4273), .ZN(n3128) );
  AOI22_X1 U3850 ( .A1(n4540), .A2(REG2_REG_11__SCAN_IN), .B1(n2520), .B2(
        n4377), .ZN(n4368) );
  NAND2_X1 U3851 ( .A1(REG2_REG_9__SCAN_IN), .A2(n4544), .ZN(n3122) );
  INV_X1 U3852 ( .A(n4544), .ZN(n4352) );
  AOI22_X1 U3853 ( .A1(REG2_REG_9__SCAN_IN), .A2(n4544), .B1(n4352), .B2(n2446), .ZN(n4349) );
  NAND2_X1 U3854 ( .A1(n4323), .A2(REG2_REG_7__SCAN_IN), .ZN(n3119) );
  AOI22_X1 U3855 ( .A1(n4323), .A2(REG2_REG_7__SCAN_IN), .B1(n2413), .B2(n4549), .ZN(n4331) );
  INV_X1 U3856 ( .A(n3134), .ZN(n4552) );
  AOI22_X1 U3857 ( .A1(REG2_REG_5__SCAN_IN), .A2(n3134), .B1(n4552), .B2(n3116), .ZN(n4310) );
  INV_X1 U3858 ( .A(n3111), .ZN(n3115) );
  INV_X1 U3859 ( .A(n3112), .ZN(n3114) );
  NAND2_X1 U3860 ( .A1(n3135), .A2(n3117), .ZN(n3118) );
  NAND2_X1 U3861 ( .A1(REG2_REG_6__SCAN_IN), .A2(n4320), .ZN(n4319) );
  NAND2_X1 U3862 ( .A1(n3118), .A2(n4319), .ZN(n4330) );
  NAND2_X1 U3863 ( .A1(n4331), .A2(n4330), .ZN(n4329) );
  NAND2_X1 U3864 ( .A1(n3119), .A2(n4329), .ZN(n3120) );
  NAND2_X1 U3865 ( .A1(n4546), .A2(n3120), .ZN(n3121) );
  INV_X1 U3866 ( .A(n4546), .ZN(n4343) );
  XNOR2_X1 U3867 ( .A(n3120), .B(n4343), .ZN(n4335) );
  NAND2_X1 U3868 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4335), .ZN(n4334) );
  NAND2_X1 U3869 ( .A1(n3121), .A2(n4334), .ZN(n4348) );
  NAND2_X1 U3870 ( .A1(n4349), .A2(n4348), .ZN(n4347) );
  NAND2_X1 U3871 ( .A1(n3122), .A2(n4347), .ZN(n3123) );
  NAND2_X1 U3872 ( .A1(n4542), .A2(n3123), .ZN(n3124) );
  INV_X1 U3873 ( .A(n4542), .ZN(n4362) );
  XNOR2_X1 U3874 ( .A(n3123), .B(n4362), .ZN(n4359) );
  NAND2_X1 U3875 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4359), .ZN(n4358) );
  NAND2_X1 U3876 ( .A1(n3124), .A2(n4358), .ZN(n4367) );
  NAND2_X1 U3877 ( .A1(n4368), .A2(n4367), .ZN(n4366) );
  NAND2_X1 U3878 ( .A1(n3142), .A2(n3125), .ZN(n3126) );
  INV_X1 U3879 ( .A(n4537), .ZN(n4399) );
  NOR2_X1 U3880 ( .A1(n4399), .A2(n2482), .ZN(n4387) );
  OAI22_X1 U3881 ( .A1(n4390), .A2(n4387), .B1(n4537), .B2(
        REG2_REG_13__SCAN_IN), .ZN(n3127) );
  NOR2_X1 U3882 ( .A1(n3127), .A2(n3128), .ZN(n3615) );
  INV_X1 U3883 ( .A(n4388), .ZN(n4430) );
  AOI211_X1 U3884 ( .C1(n3981), .C2(n3129), .A(n3614), .B(n4430), .ZN(n3130)
         );
  AOI211_X1 U3885 ( .C1(n3593), .C2(n4273), .A(n3131), .B(n3130), .ZN(n3148)
         );
  INV_X1 U3886 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3145) );
  AOI22_X1 U3887 ( .A1(n4537), .A2(REG1_REG_13__SCAN_IN), .B1(n3145), .B2(
        n4399), .ZN(n4396) );
  INV_X1 U3888 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4622) );
  AOI22_X1 U3889 ( .A1(n4540), .A2(REG1_REG_11__SCAN_IN), .B1(n4622), .B2(
        n4377), .ZN(n4374) );
  NAND2_X1 U3890 ( .A1(REG1_REG_9__SCAN_IN), .A2(n4544), .ZN(n3139) );
  INV_X1 U3891 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4619) );
  AOI22_X1 U3892 ( .A1(REG1_REG_9__SCAN_IN), .A2(n4544), .B1(n4352), .B2(n4619), .ZN(n4346) );
  INV_X1 U3893 ( .A(REG1_REG_5__SCAN_IN), .ZN(n4615) );
  AOI22_X1 U3894 ( .A1(REG1_REG_5__SCAN_IN), .A2(n4552), .B1(n3134), .B2(n4615), .ZN(n4304) );
  INV_X1 U3895 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4617) );
  NAND2_X1 U3896 ( .A1(n4546), .A2(n3137), .ZN(n3138) );
  NAND2_X1 U3897 ( .A1(REG1_REG_8__SCAN_IN), .A2(n4340), .ZN(n4339) );
  NAND2_X1 U3898 ( .A1(n4542), .A2(n3140), .ZN(n3141) );
  NAND2_X1 U3899 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4357), .ZN(n4356) );
  NAND2_X1 U3900 ( .A1(n3142), .A2(n3143), .ZN(n3144) );
  NAND2_X1 U3901 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4384), .ZN(n4383) );
  NAND2_X1 U3902 ( .A1(REG1_REG_14__SCAN_IN), .A2(n3146), .ZN(n3607) );
  OAI211_X1 U3903 ( .C1(n3146), .C2(REG1_REG_14__SCAN_IN), .A(n4438), .B(n3607), .ZN(n3147) );
  NAND2_X1 U3904 ( .A1(n3148), .A2(n3147), .ZN(U3254) );
  NAND2_X1 U3905 ( .A1(n3031), .A2(n3149), .ZN(n3150) );
  NAND2_X1 U3906 ( .A1(n3151), .A2(n3150), .ZN(n3154) );
  INV_X1 U3907 ( .A(n3152), .ZN(n3153) );
  AOI21_X1 U3908 ( .B1(n3155), .B2(n3154), .A(n3153), .ZN(n3161) );
  NOR2_X1 U3909 ( .A1(STATE_REG_SCAN_IN), .A2(n3156), .ZN(n4354) );
  INV_X1 U3910 ( .A(n3576), .ZN(n4447) );
  OAI22_X1 U3911 ( .A1(n2218), .A2(n4280), .B1(n4281), .B2(n4447), .ZN(n3157)
         );
  AOI211_X1 U3912 ( .C1(n3206), .C2(n4284), .A(n4354), .B(n3157), .ZN(n3160)
         );
  NAND2_X1 U3913 ( .A1(n3408), .A2(n3158), .ZN(n3159) );
  OAI211_X1 U3914 ( .C1(n3161), .C2(n3411), .A(n3160), .B(n3159), .ZN(U3228)
         );
  AND2_X1 U3915 ( .A1(n3152), .A2(n3162), .ZN(n3164) );
  OAI211_X1 U3916 ( .C1(n3164), .C2(n3163), .A(n4290), .B(n3171), .ZN(n3168)
         );
  NOR2_X1 U3917 ( .A1(STATE_REG_SCAN_IN), .A2(n3165), .ZN(n4364) );
  OAI22_X1 U3918 ( .A1(n3271), .A2(n4280), .B1(n4281), .B2(n3207), .ZN(n3166)
         );
  AOI211_X1 U3919 ( .C1(n3269), .C2(n4284), .A(n4364), .B(n3166), .ZN(n3167)
         );
  OAI211_X1 U3920 ( .C1(n4295), .C2(n3169), .A(n3168), .B(n3167), .ZN(U3214)
         );
  NAND2_X1 U3921 ( .A1(n3171), .A2(n3170), .ZN(n3222) );
  NAND2_X1 U3922 ( .A1(n3222), .A2(n3223), .ZN(n3221) );
  NAND2_X1 U3923 ( .A1(n3221), .A2(n3225), .ZN(n3246) );
  INV_X1 U3924 ( .A(n3247), .ZN(n3245) );
  XNOR2_X1 U3925 ( .A(n3245), .B(n3249), .ZN(n3172) );
  XNOR2_X1 U3926 ( .A(n3246), .B(n3172), .ZN(n3177) );
  INV_X1 U3927 ( .A(n3173), .ZN(n3212) );
  OAI22_X1 U3928 ( .A1(n3972), .A2(n4281), .B1(n4280), .B2(n3207), .ZN(n3175)
         );
  NAND2_X1 U3929 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4381) );
  OAI21_X1 U3930 ( .B1(n3405), .B2(n3236), .A(n4381), .ZN(n3174) );
  AOI211_X1 U3931 ( .C1(n3212), .C2(n3408), .A(n3175), .B(n3174), .ZN(n3176)
         );
  OAI21_X1 U3932 ( .B1(n3177), .B2(n3411), .A(n3176), .ZN(U3221) );
  INV_X1 U3933 ( .A(n3178), .ZN(n3179) );
  OAI21_X1 U3934 ( .B1(n3180), .B2(n2217), .A(n3179), .ZN(n4469) );
  INV_X1 U3935 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3191) );
  INV_X1 U3936 ( .A(n4596), .ZN(n4577) );
  AND2_X1 U3937 ( .A1(n3442), .A2(n3447), .ZN(n3513) );
  XOR2_X1 U3938 ( .A(n3513), .B(n3181), .Z(n3186) );
  INV_X1 U3939 ( .A(n3186), .ZN(n4471) );
  XOR2_X1 U3940 ( .A(n3182), .B(n3513), .Z(n3189) );
  AOI22_X1 U3941 ( .A1(n3577), .A2(n4479), .B1(n4478), .B2(n3183), .ZN(n3184)
         );
  OAI21_X1 U3942 ( .B1(n3185), .B2(n4482), .A(n3184), .ZN(n3188) );
  NOR2_X1 U3943 ( .A1(n3186), .A2(n4487), .ZN(n3187) );
  AOI211_X1 U3944 ( .C1(n4502), .C2(n3189), .A(n3188), .B(n3187), .ZN(n4474)
         );
  INV_X1 U3945 ( .A(n4474), .ZN(n3190) );
  AOI21_X1 U3946 ( .B1(n4577), .B2(n4471), .A(n3190), .ZN(n3193) );
  MUX2_X1 U3947 ( .A(n3191), .B(n3193), .S(n4624), .Z(n3192) );
  OAI21_X1 U3948 ( .B1(n4469), .B2(n4201), .A(n3192), .ZN(U3526) );
  INV_X1 U3949 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3194) );
  MUX2_X1 U3950 ( .A(n3194), .B(n3193), .S(n4605), .Z(n3195) );
  OAI21_X1 U3951 ( .B1(n4469), .B2(n4259), .A(n3195), .ZN(U3483) );
  INV_X1 U3952 ( .A(n3197), .ZN(n3198) );
  NAND2_X1 U3953 ( .A1(n3199), .A2(n3443), .ZN(n3268) );
  INV_X1 U3954 ( .A(n3269), .ZN(n3263) );
  NAND2_X1 U3955 ( .A1(n3576), .A2(n3263), .ZN(n3418) );
  NAND2_X1 U3956 ( .A1(n3268), .A2(n3418), .ZN(n3200) );
  NAND2_X1 U3957 ( .A1(n4447), .A2(n3269), .ZN(n3415) );
  NAND2_X1 U3958 ( .A1(n3200), .A2(n3415), .ZN(n4444) );
  INV_X1 U3959 ( .A(n4457), .ZN(n3220) );
  NAND2_X1 U3960 ( .A1(n3575), .A2(n3220), .ZN(n3419) );
  NAND2_X1 U3961 ( .A1(n4444), .A2(n3419), .ZN(n3201) );
  NAND2_X1 U3962 ( .A1(n3207), .A2(n4457), .ZN(n3421) );
  XNOR2_X1 U3963 ( .A(n4445), .B(n3235), .ZN(n3487) );
  XNOR2_X1 U3964 ( .A(n3230), .B(n3487), .ZN(n3202) );
  NAND2_X1 U3965 ( .A1(n3202), .A2(n4502), .ZN(n3204) );
  AOI22_X1 U3966 ( .A1(n3627), .A2(n4479), .B1(n4478), .B2(n3235), .ZN(n3203)
         );
  OAI211_X1 U3967 ( .C1(n3207), .C2(n4482), .A(n3204), .B(n3203), .ZN(n3282)
         );
  INV_X1 U3968 ( .A(n3282), .ZN(n3216) );
  NAND2_X1 U3969 ( .A1(n3577), .A2(n3206), .ZN(n3265) );
  NAND2_X1 U3970 ( .A1(n4447), .A2(n3263), .ZN(n4448) );
  NAND2_X1 U3971 ( .A1(n3207), .A2(n3220), .ZN(n3208) );
  AND2_X1 U3972 ( .A1(n4448), .A2(n3208), .ZN(n3210) );
  INV_X1 U3973 ( .A(n3208), .ZN(n3209) );
  NAND2_X1 U3974 ( .A1(n3421), .A2(n3419), .ZN(n3508) );
  XOR2_X1 U3975 ( .A(n3487), .B(n3238), .Z(n3283) );
  INV_X1 U3976 ( .A(n3239), .ZN(n3211) );
  OAI21_X1 U3977 ( .B1(n2081), .B2(n3236), .A(n3211), .ZN(n3289) );
  AOI22_X1 U3978 ( .A1(n4296), .A2(REG2_REG_12__SCAN_IN), .B1(n3212), .B2(
        n4491), .ZN(n3213) );
  OAI21_X1 U3979 ( .B1(n3289), .B2(n3961), .A(n3213), .ZN(n3214) );
  AOI21_X1 U3980 ( .B1(n3283), .B2(n3965), .A(n3214), .ZN(n3215) );
  OAI21_X1 U3981 ( .B1(n4296), .B2(n3216), .A(n3215), .ZN(U3278) );
  AOI22_X1 U3982 ( .A1(n3218), .A2(n4445), .B1(n3217), .B2(n3576), .ZN(n3219)
         );
  NAND2_X1 U3983 ( .A1(REG3_REG_11__SCAN_IN), .A2(U3149), .ZN(n4369) );
  OAI211_X1 U3984 ( .C1(n3405), .C2(n3220), .A(n3219), .B(n4369), .ZN(n3228)
         );
  INV_X1 U3985 ( .A(n3221), .ZN(n3226) );
  AOI21_X1 U3986 ( .B1(n3225), .B2(n3223), .A(n3222), .ZN(n3224) );
  AOI211_X1 U3987 ( .C1(n3226), .C2(n3225), .A(n3411), .B(n3224), .ZN(n3227)
         );
  AOI211_X1 U3988 ( .C1(n3408), .C2(n4455), .A(n3228), .B(n3227), .ZN(n3229)
         );
  INV_X1 U3989 ( .A(n3229), .ZN(U3233) );
  NOR2_X1 U3990 ( .A1(n4445), .A2(n3236), .ZN(n3422) );
  NAND2_X1 U3991 ( .A1(n4445), .A2(n3236), .ZN(n3416) );
  NAND2_X1 U3992 ( .A1(n3531), .A2(n3416), .ZN(n3231) );
  NAND2_X1 U3993 ( .A1(n3972), .A2(n3626), .ZN(n3532) );
  NAND2_X1 U3994 ( .A1(n3627), .A2(n3636), .ZN(n3417) );
  AND2_X1 U3995 ( .A1(n3532), .A2(n3417), .ZN(n3488) );
  XOR2_X1 U3996 ( .A(n3231), .B(n3488), .Z(n3234) );
  AOI22_X1 U3997 ( .A1(n3574), .A2(n4479), .B1(n4478), .B2(n3626), .ZN(n3232)
         );
  OAI21_X1 U3998 ( .B1(n3257), .B2(n4482), .A(n3232), .ZN(n3233) );
  AOI21_X1 U3999 ( .B1(n3234), .B2(n4502), .A(n3233), .ZN(n4209) );
  NOR2_X1 U4000 ( .A1(n4445), .A2(n3235), .ZN(n3237) );
  XNOR2_X1 U4001 ( .A(n3951), .B(n3488), .ZN(n4207) );
  OR2_X1 U4002 ( .A1(n3239), .A2(n3636), .ZN(n3240) );
  NAND2_X1 U4003 ( .A1(n3979), .A2(n3240), .ZN(n4210) );
  NOR2_X1 U4004 ( .A1(n4515), .A2(n3261), .ZN(n3241) );
  AOI21_X1 U4005 ( .B1(n4296), .B2(REG2_REG_13__SCAN_IN), .A(n3241), .ZN(n3242) );
  OAI21_X1 U4006 ( .B1(n4210), .B2(n3961), .A(n3242), .ZN(n3243) );
  AOI21_X1 U4007 ( .B1(n4207), .B2(n3965), .A(n3243), .ZN(n3244) );
  OAI21_X1 U4008 ( .B1(n4209), .B2(n4296), .A(n3244), .ZN(U3277) );
  NOR2_X1 U4009 ( .A1(n3246), .A2(n3245), .ZN(n3250) );
  INV_X1 U4010 ( .A(n3246), .ZN(n3248) );
  OAI22_X1 U4011 ( .A1(n3250), .A2(n3249), .B1(n3248), .B2(n3247), .ZN(n3254)
         );
  NAND2_X1 U4012 ( .A1(n3252), .A2(n3251), .ZN(n3253) );
  XNOR2_X1 U4013 ( .A(n3254), .B(n3253), .ZN(n3255) );
  NAND2_X1 U4014 ( .A1(n3255), .A2(n4290), .ZN(n3260) );
  INV_X1 U4015 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3256) );
  NOR2_X1 U4016 ( .A1(STATE_REG_SCAN_IN), .A2(n3256), .ZN(n4392) );
  OAI22_X1 U4017 ( .A1(n3257), .A2(n4280), .B1(n4281), .B2(n4279), .ZN(n3258)
         );
  AOI211_X1 U4018 ( .C1(n3626), .C2(n4284), .A(n4392), .B(n3258), .ZN(n3259)
         );
  OAI211_X1 U4019 ( .C1(n4295), .C2(n3261), .A(n3260), .B(n3259), .ZN(U3231)
         );
  INV_X1 U4020 ( .A(n3262), .ZN(n3264) );
  OAI21_X1 U4021 ( .B1(n3264), .B2(n3263), .A(n4456), .ZN(n4462) );
  INV_X1 U4022 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3277) );
  AND2_X1 U4023 ( .A1(n3415), .A2(n3418), .ZN(n3486) );
  NAND2_X1 U4024 ( .A1(n3266), .A2(n3265), .ZN(n3267) );
  XOR2_X1 U4025 ( .A(n3486), .B(n3267), .Z(n3272) );
  INV_X1 U4026 ( .A(n3272), .ZN(n4464) );
  XNOR2_X1 U4027 ( .A(n3268), .B(n3486), .ZN(n3275) );
  AOI22_X1 U4028 ( .A1(n3575), .A2(n4479), .B1(n4478), .B2(n3269), .ZN(n3270)
         );
  OAI21_X1 U4029 ( .B1(n3271), .B2(n4482), .A(n3270), .ZN(n3274) );
  NOR2_X1 U4030 ( .A1(n3272), .A2(n4487), .ZN(n3273) );
  AOI211_X1 U4031 ( .C1(n3275), .C2(n4502), .A(n3274), .B(n3273), .ZN(n4467)
         );
  INV_X1 U4032 ( .A(n4467), .ZN(n3276) );
  AOI21_X1 U4033 ( .B1(n4577), .B2(n4464), .A(n3276), .ZN(n3279) );
  MUX2_X1 U4034 ( .A(n3277), .B(n3279), .S(n4605), .Z(n3278) );
  OAI21_X1 U4035 ( .B1(n4462), .B2(n4259), .A(n3278), .ZN(U3487) );
  INV_X1 U4036 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3280) );
  MUX2_X1 U4037 ( .A(n3280), .B(n3279), .S(n4624), .Z(n3281) );
  OAI21_X1 U4038 ( .B1(n4462), .B2(n4201), .A(n3281), .ZN(U3528) );
  AOI21_X1 U4039 ( .B1(n3283), .B2(n4594), .A(n3282), .ZN(n3287) );
  INV_X1 U4040 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3284) );
  MUX2_X1 U4041 ( .A(n3287), .B(n3284), .S(n4603), .Z(n3285) );
  OAI21_X1 U4042 ( .B1(n3289), .B2(n4259), .A(n3285), .ZN(U3491) );
  INV_X1 U40430 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3286) );
  MUX2_X1 U4044 ( .A(n3287), .B(n3286), .S(n4621), .Z(n3288) );
  OAI21_X1 U4045 ( .B1(n3289), .B2(n4201), .A(n3288), .ZN(U3530) );
  NAND2_X1 U4046 ( .A1(n2363), .A2(DATAI_31_), .ZN(n3475) );
  NAND2_X1 U4047 ( .A1(n2363), .A2(DATAI_29_), .ZN(n3693) );
  AND2_X1 U4048 ( .A1(n2363), .A2(DATAI_30_), .ZN(n3989) );
  XOR2_X1 U4049 ( .A(n3475), .B(n3986), .Z(n4297) );
  INV_X1 U4050 ( .A(n4297), .ZN(n3294) );
  INV_X1 U4051 ( .A(REG0_REG_31__SCAN_IN), .ZN(n3290) );
  INV_X1 U4052 ( .A(n3475), .ZN(n3558) );
  AOI21_X1 U4053 ( .B1(B_REG_SCAN_IN), .B2(n4265), .A(n4505), .ZN(n3686) );
  AND2_X1 U4054 ( .A1(n3556), .A2(n3686), .ZN(n3988) );
  AOI21_X1 U4055 ( .B1(n3558), .B2(n4478), .A(n3988), .ZN(n4299) );
  MUX2_X1 U4056 ( .A(n3290), .B(n4299), .S(n4605), .Z(n3291) );
  OAI21_X1 U4057 ( .B1(n3294), .B2(n4259), .A(n3291), .ZN(U3517) );
  INV_X1 U4058 ( .A(REG1_REG_31__SCAN_IN), .ZN(n3292) );
  MUX2_X1 U4059 ( .A(n3292), .B(n4299), .S(n4624), .Z(n3293) );
  OAI21_X1 U4060 ( .B1(n3294), .B2(n4201), .A(n3293), .ZN(U3549) );
  XNOR2_X1 U4061 ( .A(n3296), .B(n3295), .ZN(n3297) );
  XNOR2_X1 U4062 ( .A(n3298), .B(n3297), .ZN(n3304) );
  INV_X1 U4063 ( .A(n3980), .ZN(n3302) );
  INV_X1 U4064 ( .A(n3970), .ZN(n3414) );
  OAI22_X1 U4065 ( .A1(n3972), .A2(n4280), .B1(n4281), .B2(n3414), .ZN(n3301)
         );
  INV_X1 U4066 ( .A(n3978), .ZN(n3628) );
  OAI21_X1 U4067 ( .B1(n3405), .B2(n3628), .A(n3299), .ZN(n3300) );
  AOI211_X1 U4068 ( .C1(n3302), .C2(n3408), .A(n3301), .B(n3300), .ZN(n3303)
         );
  OAI21_X1 U4069 ( .B1(n3304), .B2(n3411), .A(n3303), .ZN(U3212) );
  AOI22_X1 U4070 ( .A1(n4284), .A2(n4493), .B1(REG3_REG_0__SCAN_IN), .B2(n3305), .ZN(n3308) );
  NAND2_X1 U4071 ( .A1(n3306), .A2(n4290), .ZN(n3307) );
  OAI211_X1 U4072 ( .C1(n4506), .C2(n4281), .A(n3308), .B(n3307), .ZN(U3229)
         );
  INV_X1 U4073 ( .A(n3309), .ZN(n3313) );
  OAI21_X1 U4074 ( .B1(n3382), .B2(n3311), .A(n3310), .ZN(n3312) );
  NAND3_X1 U4075 ( .A1(n3313), .A2(n4290), .A3(n3312), .ZN(n3318) );
  OAI22_X1 U4076 ( .A1(n3405), .A2(n3809), .B1(STATE_REG_SCAN_IN), .B2(n3314), 
        .ZN(n3316) );
  OAI22_X1 U4077 ( .A1(n3765), .A2(n4281), .B1(n4280), .B2(n3468), .ZN(n3315)
         );
  NOR2_X1 U4078 ( .A1(n3316), .A2(n3315), .ZN(n3317) );
  OAI211_X1 U4079 ( .C1(n4295), .C2(n3798), .A(n3318), .B(n3317), .ZN(U3213)
         );
  XOR2_X1 U4080 ( .A(n3320), .B(n3319), .Z(n3325) );
  INV_X1 U4081 ( .A(n3321), .ZN(n3885) );
  INV_X1 U4082 ( .A(n3909), .ZN(n3881) );
  INV_X1 U4083 ( .A(n3878), .ZN(n3839) );
  OAI22_X1 U4084 ( .A1(n3881), .A2(n4280), .B1(n4281), .B2(n3839), .ZN(n3323)
         );
  NAND2_X1 U4085 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3623) );
  OAI21_X1 U4086 ( .B1(n3405), .B2(n3644), .A(n3623), .ZN(n3322) );
  AOI211_X1 U4087 ( .C1(n3885), .C2(n3408), .A(n3323), .B(n3322), .ZN(n3324)
         );
  OAI21_X1 U4088 ( .B1(n3325), .B2(n3411), .A(n3324), .ZN(U3216) );
  XNOR2_X1 U4089 ( .A(n3328), .B(n3327), .ZN(n3329) );
  XNOR2_X1 U4090 ( .A(n3326), .B(n3329), .ZN(n3334) );
  INV_X1 U4091 ( .A(n3330), .ZN(n3842) );
  OAI22_X1 U4092 ( .A1(n3839), .A2(n4280), .B1(n4281), .B2(n3468), .ZN(n3332)
         );
  INV_X1 U4093 ( .A(REG3_REG_21__SCAN_IN), .ZN(n4089) );
  OAI22_X1 U4094 ( .A1(n3405), .A2(n3841), .B1(STATE_REG_SCAN_IN), .B2(n4089), 
        .ZN(n3331) );
  AOI211_X1 U4095 ( .C1(n3842), .C2(n3408), .A(n3332), .B(n3331), .ZN(n3333)
         );
  OAI21_X1 U4096 ( .B1(n3334), .B2(n3411), .A(n3333), .ZN(U3220) );
  NOR2_X1 U4097 ( .A1(n3336), .A2(n2129), .ZN(n3337) );
  XNOR2_X1 U4098 ( .A(n3338), .B(n3337), .ZN(n3344) );
  INV_X1 U4099 ( .A(n3339), .ZN(n3768) );
  OAI22_X1 U4100 ( .A1(n3765), .A2(n4280), .B1(n4281), .B2(n3731), .ZN(n3342)
         );
  INV_X1 U4101 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3340) );
  OAI22_X1 U4102 ( .A1(n3405), .A2(n3767), .B1(STATE_REG_SCAN_IN), .B2(n3340), 
        .ZN(n3341) );
  AOI211_X1 U4103 ( .C1(n3768), .C2(n3408), .A(n3342), .B(n3341), .ZN(n3343)
         );
  OAI21_X1 U4104 ( .B1(n3344), .B2(n3411), .A(n3343), .ZN(U3222) );
  NOR2_X1 U4105 ( .A1(n4286), .A2(n4291), .ZN(n3346) );
  XNOR2_X1 U4106 ( .A(n3346), .B(n3345), .ZN(n3351) );
  INV_X1 U4107 ( .A(n3347), .ZN(n3939) );
  OAI22_X1 U4108 ( .A1(n3414), .A2(n4280), .B1(n4281), .B2(n3893), .ZN(n3349)
         );
  INV_X1 U4109 ( .A(n3936), .ZN(n3929) );
  NAND2_X1 U4110 ( .A1(REG3_REG_16__SCAN_IN), .A2(U3149), .ZN(n4410) );
  OAI21_X1 U4111 ( .B1(n3405), .B2(n3929), .A(n4410), .ZN(n3348) );
  AOI211_X1 U4112 ( .C1(n3939), .C2(n3408), .A(n3349), .B(n3348), .ZN(n3350)
         );
  OAI21_X1 U4113 ( .B1(n3351), .B2(n3411), .A(n3350), .ZN(U3223) );
  XNOR2_X1 U4114 ( .A(n3353), .B(n3352), .ZN(n3354) );
  XNOR2_X1 U4115 ( .A(n3355), .B(n3354), .ZN(n3356) );
  NAND2_X1 U4116 ( .A1(n3356), .A2(n4290), .ZN(n3359) );
  AND2_X1 U4117 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4423) );
  INV_X1 U4118 ( .A(n3947), .ZN(n4282) );
  OAI22_X1 U4119 ( .A1(n4282), .A2(n4280), .B1(n4281), .B2(n3881), .ZN(n3357)
         );
  AOI211_X1 U4120 ( .C1(n3642), .C2(n4284), .A(n4423), .B(n3357), .ZN(n3358)
         );
  OAI211_X1 U4121 ( .C1(n4295), .C2(n3917), .A(n3359), .B(n3358), .ZN(U3225)
         );
  INV_X1 U4122 ( .A(n3360), .ZN(n3362) );
  NAND2_X1 U4123 ( .A1(n3362), .A2(n3361), .ZN(n3364) );
  XNOR2_X1 U4124 ( .A(n3364), .B(n3363), .ZN(n3369) );
  INV_X1 U4125 ( .A(n3365), .ZN(n3787) );
  OAI22_X1 U4126 ( .A1(n3823), .A2(n4280), .B1(n4281), .B2(n3783), .ZN(n3367)
         );
  OAI22_X1 U4127 ( .A1(n3405), .A2(n3786), .B1(STATE_REG_SCAN_IN), .B2(n4037), 
        .ZN(n3366) );
  AOI211_X1 U4128 ( .C1(n3787), .C2(n3408), .A(n3367), .B(n3366), .ZN(n3368)
         );
  OAI21_X1 U4129 ( .B1(n3369), .B2(n3411), .A(n3368), .ZN(U3226) );
  INV_X1 U4130 ( .A(n3370), .ZN(n3375) );
  AOI21_X1 U4131 ( .B1(n3374), .B2(n3372), .A(n3371), .ZN(n3373) );
  AOI21_X1 U4132 ( .B1(n3375), .B2(n3374), .A(n3373), .ZN(n3381) );
  INV_X1 U4133 ( .A(n3376), .ZN(n3862) );
  INV_X1 U4134 ( .A(n3855), .ZN(n3469) );
  OAI22_X1 U4135 ( .A1(n3858), .A2(n4280), .B1(n4281), .B2(n3469), .ZN(n3379)
         );
  INV_X1 U4136 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3377) );
  OAI22_X1 U4137 ( .A1(n3405), .A2(n3861), .B1(STATE_REG_SCAN_IN), .B2(n3377), 
        .ZN(n3378) );
  AOI211_X1 U4138 ( .C1(n3862), .C2(n3408), .A(n3379), .B(n3378), .ZN(n3380)
         );
  OAI21_X1 U4139 ( .B1(n3381), .B2(n3411), .A(n3380), .ZN(U3230) );
  AOI21_X1 U4140 ( .B1(n3384), .B2(n3383), .A(n3382), .ZN(n3390) );
  INV_X1 U4141 ( .A(n3385), .ZN(n3826) );
  OAI22_X1 U4142 ( .A1(n3823), .A2(n4281), .B1(n4280), .B2(n3469), .ZN(n3388)
         );
  OAI22_X1 U4143 ( .A1(n3405), .A2(n3471), .B1(STATE_REG_SCAN_IN), .B2(n3386), 
        .ZN(n3387) );
  AOI211_X1 U4144 ( .C1(n3826), .C2(n3408), .A(n3388), .B(n3387), .ZN(n3389)
         );
  OAI21_X1 U4145 ( .B1(n3390), .B2(n3411), .A(n3389), .ZN(U3232) );
  INV_X1 U4146 ( .A(n3391), .ZN(n3393) );
  NOR2_X1 U4147 ( .A1(n3393), .A2(n3392), .ZN(n3394) );
  XNOR2_X1 U4148 ( .A(n3395), .B(n3394), .ZN(n3396) );
  NAND2_X1 U4149 ( .A1(n3396), .A2(n4290), .ZN(n3399) );
  INV_X1 U4150 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4112) );
  NOR2_X1 U4151 ( .A1(STATE_REG_SCAN_IN), .A2(n4112), .ZN(n4435) );
  OAI22_X1 U4152 ( .A1(n3858), .A2(n4281), .B1(n4280), .B2(n3893), .ZN(n3397)
         );
  AOI211_X1 U4153 ( .C1(n3896), .C2(n4284), .A(n4435), .B(n3397), .ZN(n3398)
         );
  OAI211_X1 U4154 ( .C1(n4295), .C2(n3898), .A(n3399), .B(n3398), .ZN(U3235)
         );
  NAND2_X1 U4155 ( .A1(n2131), .A2(n3401), .ZN(n3402) );
  XNOR2_X1 U4156 ( .A(n3403), .B(n3402), .ZN(n3412) );
  INV_X1 U4157 ( .A(n3748), .ZN(n3409) );
  OAI22_X1 U4158 ( .A1(n3783), .A2(n4280), .B1(n4281), .B2(n3708), .ZN(n3407)
         );
  INV_X1 U4159 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3404) );
  OAI22_X1 U4160 ( .A1(n3405), .A2(n3746), .B1(STATE_REG_SCAN_IN), .B2(n3404), 
        .ZN(n3406) );
  AOI211_X1 U4161 ( .C1(n3409), .C2(n3408), .A(n3407), .B(n3406), .ZN(n3410)
         );
  OAI21_X1 U4162 ( .B1(n3412), .B2(n3411), .A(n3410), .ZN(U3237) );
  AND2_X1 U4163 ( .A1(n3855), .A2(n3841), .ZN(n3543) );
  NAND2_X1 U4164 ( .A1(n4282), .A2(n3936), .ZN(n3537) );
  NAND2_X1 U4165 ( .A1(n3947), .A2(n3929), .ZN(n3536) );
  INV_X1 U4166 ( .A(n4285), .ZN(n3413) );
  NAND2_X1 U4167 ( .A1(n3970), .A2(n3413), .ZN(n3666) );
  NAND2_X1 U4168 ( .A1(n3574), .A2(n3628), .ZN(n3511) );
  NAND2_X1 U4169 ( .A1(n3666), .A2(n3511), .ZN(n3451) );
  NAND2_X1 U4170 ( .A1(n3414), .A2(n4285), .ZN(n3533) );
  NAND2_X1 U4171 ( .A1(n3451), .A2(n3533), .ZN(n3534) );
  INV_X1 U4172 ( .A(n3534), .ZN(n3457) );
  INV_X1 U4173 ( .A(n3415), .ZN(n3425) );
  AND2_X1 U4174 ( .A1(n3417), .A2(n3416), .ZN(n3530) );
  AND2_X1 U4175 ( .A1(n3419), .A2(n3418), .ZN(n3420) );
  AND2_X1 U4176 ( .A1(n3530), .A2(n3420), .ZN(n3453) );
  OAI21_X1 U4177 ( .B1(n2119), .B2(n3422), .A(n3530), .ZN(n3423) );
  NAND2_X1 U4178 ( .A1(n4279), .A2(n3978), .ZN(n3665) );
  NAND4_X1 U4179 ( .A1(n3423), .A2(n3665), .A3(n3532), .A4(n3533), .ZN(n3424)
         );
  AOI21_X1 U4180 ( .B1(n3425), .B2(n3453), .A(n3424), .ZN(n3456) );
  INV_X1 U4181 ( .A(n3518), .ZN(n4476) );
  NAND2_X1 U4182 ( .A1(n3584), .A2(n4508), .ZN(n3517) );
  OAI211_X1 U4183 ( .C1(n4476), .C2(n4270), .A(n3517), .B(n3426), .ZN(n3428)
         );
  NAND3_X1 U4184 ( .A1(n3428), .A2(n2934), .A3(n3427), .ZN(n3430) );
  OAI211_X1 U4185 ( .C1(n3432), .C2(n3431), .A(n3430), .B(n3429), .ZN(n3435)
         );
  NAND3_X1 U4186 ( .A1(n3435), .A2(n3434), .A3(n3433), .ZN(n3438) );
  NAND4_X1 U4187 ( .A1(n3438), .A2(n3437), .A3(n3436), .A4(n3446), .ZN(n3440)
         );
  NAND3_X1 U4188 ( .A1(n3440), .A2(n3520), .A3(n3439), .ZN(n3441) );
  NAND3_X1 U4189 ( .A1(n3441), .A2(n3448), .A3(n3447), .ZN(n3444) );
  AND3_X1 U4190 ( .A1(n3444), .A2(n3443), .A3(n3442), .ZN(n3452) );
  INV_X1 U4191 ( .A(n3445), .ZN(n3449) );
  NAND4_X1 U4192 ( .A1(n3449), .A2(n3448), .A3(n3447), .A4(n3446), .ZN(n3450)
         );
  OAI22_X1 U4193 ( .A1(n3452), .A2(n3451), .B1(n3457), .B2(n3450), .ZN(n3454)
         );
  NAND3_X1 U4194 ( .A1(n3454), .A2(n3453), .A3(n3198), .ZN(n3455) );
  OAI21_X1 U4195 ( .B1(n3457), .B2(n3456), .A(n3455), .ZN(n3458) );
  NAND2_X1 U4196 ( .A1(n3536), .A2(n3458), .ZN(n3461) );
  AND2_X1 U4197 ( .A1(n3878), .A2(n3861), .ZN(n3672) );
  INV_X1 U4198 ( .A(n3896), .ZN(n3459) );
  NAND2_X1 U4199 ( .A1(n3909), .A2(n3459), .ZN(n3872) );
  NAND2_X1 U4200 ( .A1(n3891), .A2(n3644), .ZN(n3460) );
  AND2_X1 U4201 ( .A1(n3872), .A2(n3460), .ZN(n3462) );
  NAND2_X1 U4202 ( .A1(n3926), .A2(n3916), .ZN(n3871) );
  NAND2_X1 U4203 ( .A1(n3462), .A2(n3871), .ZN(n3668) );
  AOI211_X1 U4204 ( .C1(n3537), .C2(n3461), .A(n3672), .B(n3668), .ZN(n3467)
         );
  NAND2_X1 U4205 ( .A1(n3881), .A2(n3896), .ZN(n3874) );
  NAND2_X1 U4206 ( .A1(n3893), .A2(n3642), .ZN(n3869) );
  NAND2_X1 U4207 ( .A1(n3874), .A2(n3869), .ZN(n3463) );
  NAND2_X1 U4208 ( .A1(n3463), .A2(n3462), .ZN(n3465) );
  NAND2_X1 U4209 ( .A1(n3858), .A2(n3882), .ZN(n3464) );
  NAND2_X1 U4210 ( .A1(n3465), .A2(n3464), .ZN(n3848) );
  NOR2_X1 U4211 ( .A1(n3878), .A2(n3861), .ZN(n3466) );
  INV_X1 U4212 ( .A(n3672), .ZN(n3539) );
  NOR2_X1 U4213 ( .A1(n3467), .A2(n3670), .ZN(n3470) );
  NAND2_X1 U4214 ( .A1(n3468), .A2(n3824), .ZN(n3803) );
  NAND2_X1 U4215 ( .A1(n3469), .A2(n3835), .ZN(n3801) );
  OAI21_X1 U4216 ( .B1(n3543), .B2(n3470), .A(n3673), .ZN(n3472) );
  NAND2_X1 U4217 ( .A1(n3836), .A2(n3471), .ZN(n3512) );
  NAND2_X1 U4218 ( .A1(n3780), .A2(n3809), .ZN(n3501) );
  AND2_X1 U4219 ( .A1(n3512), .A2(n3501), .ZN(n3544) );
  INV_X1 U4220 ( .A(n3767), .ZN(n3656) );
  NAND2_X1 U4221 ( .A1(n3783), .A2(n3656), .ZN(n3734) );
  NAND2_X1 U4222 ( .A1(n3731), .A2(n3659), .ZN(n3490) );
  NAND2_X1 U4223 ( .A1(n3734), .A2(n3490), .ZN(n3549) );
  NAND2_X1 U4224 ( .A1(n3823), .A2(n3797), .ZN(n3774) );
  NAND2_X1 U4225 ( .A1(n3765), .A2(n3779), .ZN(n3502) );
  INV_X1 U4226 ( .A(n3676), .ZN(n3546) );
  AOI211_X1 U4227 ( .C1(n3472), .C2(n3544), .A(n3549), .B(n3546), .ZN(n3474)
         );
  NAND2_X1 U4228 ( .A1(n3738), .A2(n3660), .ZN(n3489) );
  INV_X1 U4229 ( .A(n3489), .ZN(n3473) );
  NAND2_X1 U4230 ( .A1(n3806), .A2(n3786), .ZN(n3756) );
  NAND2_X1 U4231 ( .A1(n3737), .A2(n3767), .ZN(n3500) );
  AND2_X1 U4232 ( .A1(n3756), .A2(n3500), .ZN(n3548) );
  NAND2_X1 U4233 ( .A1(n3762), .A2(n3746), .ZN(n3526) );
  OAI21_X1 U4234 ( .B1(n3549), .B2(n3548), .A(n3526), .ZN(n3677) );
  INV_X1 U4235 ( .A(n3693), .ZN(n3685) );
  NAND2_X1 U4236 ( .A1(n3728), .A2(n3712), .ZN(n3682) );
  OAI21_X1 U4237 ( .B1(n3477), .B2(n3685), .A(n3682), .ZN(n3527) );
  NOR4_X1 U4238 ( .A1(n3474), .A2(n3473), .A3(n3677), .A4(n3527), .ZN(n3485)
         );
  NAND2_X1 U4239 ( .A1(n3556), .A2(n3475), .ZN(n3482) );
  INV_X1 U4240 ( .A(n3989), .ZN(n3557) );
  OR2_X1 U4241 ( .A1(n3687), .A2(n3557), .ZN(n3476) );
  AND2_X1 U4242 ( .A1(n3482), .A2(n3476), .ZN(n3492) );
  NAND2_X1 U4243 ( .A1(n3477), .A2(n3685), .ZN(n3478) );
  NAND2_X1 U4244 ( .A1(n3492), .A2(n3478), .ZN(n3480) );
  INV_X1 U4245 ( .A(n3480), .ZN(n3481) );
  NAND2_X1 U4246 ( .A1(n3689), .A2(n3704), .ZN(n3680) );
  NAND2_X1 U4247 ( .A1(n3708), .A2(n3727), .ZN(n3679) );
  NAND2_X1 U4248 ( .A1(n3680), .A2(n3679), .ZN(n3479) );
  NOR2_X1 U4249 ( .A1(n3480), .A2(n3479), .ZN(n3550) );
  AOI21_X1 U4250 ( .B1(n3481), .B2(n3527), .A(n3550), .ZN(n3554) );
  INV_X1 U4251 ( .A(n3482), .ZN(n3484) );
  INV_X1 U4252 ( .A(n3556), .ZN(n3559) );
  INV_X1 U4253 ( .A(n3687), .ZN(n3483) );
  NOR2_X1 U4254 ( .A1(n3483), .A2(n3989), .ZN(n3560) );
  AOI21_X1 U4255 ( .B1(n3558), .B2(n3559), .A(n3560), .ZN(n3491) );
  OAI22_X1 U4256 ( .A1(n3485), .A2(n3554), .B1(n3484), .B2(n3491), .ZN(n3566)
         );
  INV_X1 U4257 ( .A(n3543), .ZN(n3800) );
  NAND2_X1 U4258 ( .A1(n3800), .A2(n3801), .ZN(n3833) );
  INV_X1 U4259 ( .A(n3833), .ZN(n3499) );
  NAND4_X1 U4260 ( .A1(n3944), .A2(n3488), .A3(n3487), .A4(n3486), .ZN(n3495)
         );
  XOR2_X1 U4261 ( .A(n3693), .B(n3705), .Z(n3684) );
  NAND4_X1 U4262 ( .A1(n3684), .A2(n3701), .A3(n3901), .A4(n3935), .ZN(n3494)
         );
  NAND4_X1 U4263 ( .A1(n3724), .A2(n3744), .A3(n3492), .A4(n3491), .ZN(n3493)
         );
  NOR3_X1 U4264 ( .A1(n3495), .A2(n3494), .A3(n3493), .ZN(n3498) );
  INV_X1 U4265 ( .A(n3861), .ZN(n3496) );
  AND2_X1 U4266 ( .A1(n3878), .A2(n3496), .ZN(n3647) );
  INV_X1 U4267 ( .A(n3647), .ZN(n3497) );
  NAND2_X1 U4268 ( .A1(n3839), .A2(n3861), .ZN(n3646) );
  NAND2_X1 U4269 ( .A1(n3497), .A2(n3646), .ZN(n3851) );
  NAND3_X1 U4270 ( .A1(n3499), .A2(n3498), .A3(n3851), .ZN(n3507) );
  NAND2_X1 U4271 ( .A1(n3734), .A2(n3500), .ZN(n3758) );
  INV_X1 U4272 ( .A(n3758), .ZN(n3505) );
  NAND2_X1 U4273 ( .A1(n3774), .A2(n3501), .ZN(n3794) );
  INV_X1 U4274 ( .A(n3794), .ZN(n3804) );
  NAND2_X1 U4275 ( .A1(n3502), .A2(n3756), .ZN(n3777) );
  INV_X1 U4276 ( .A(n3777), .ZN(n3503) );
  NAND4_X1 U4277 ( .A1(n3505), .A2(n3804), .A3(n3504), .A4(n3503), .ZN(n3506)
         );
  NOR2_X1 U4278 ( .A1(n3507), .A2(n3506), .ZN(n3525) );
  INV_X1 U4279 ( .A(n3508), .ZN(n4450) );
  AND2_X1 U4280 ( .A1(n3869), .A2(n3871), .ZN(n3914) );
  NAND4_X1 U4281 ( .A1(n4450), .A2(n3510), .A3(n3509), .A4(n3914), .ZN(n3516)
         );
  NAND2_X1 U4282 ( .A1(n3665), .A2(n3511), .ZN(n3954) );
  NAND2_X1 U4283 ( .A1(n3803), .A2(n3512), .ZN(n3816) );
  INV_X1 U4284 ( .A(n3816), .ZN(n3819) );
  NAND4_X1 U4285 ( .A1(n3973), .A2(n3819), .A3(n3514), .A4(n3513), .ZN(n3515)
         );
  NOR2_X1 U4286 ( .A1(n3516), .A2(n3515), .ZN(n3524) );
  NAND2_X1 U4287 ( .A1(n3518), .A2(n3517), .ZN(n4555) );
  NOR2_X1 U4288 ( .A1(n4486), .A2(n4555), .ZN(n3521) );
  XNOR2_X1 U4289 ( .A(n3891), .B(n3644), .ZN(n3867) );
  INV_X1 U4290 ( .A(n3867), .ZN(n3875) );
  AND4_X1 U4291 ( .A1(n3521), .A2(n3520), .A3(n3519), .A4(n3875), .ZN(n3522)
         );
  NAND4_X1 U4292 ( .A1(n3525), .A2(n3524), .A3(n3523), .A4(n3522), .ZN(n3564)
         );
  INV_X1 U4293 ( .A(n3724), .ZN(n3529) );
  INV_X1 U4294 ( .A(n3526), .ZN(n3528) );
  NOR3_X1 U4295 ( .A1(n3529), .A2(n3528), .A3(n3527), .ZN(n3553) );
  NAND2_X1 U4296 ( .A1(n3665), .A2(n3533), .ZN(n3535) );
  OAI21_X1 U4297 ( .B1(n3969), .B2(n3535), .A(n3534), .ZN(n3538) );
  INV_X1 U4298 ( .A(n3536), .ZN(n3667) );
  AOI211_X1 U4299 ( .C1(n3538), .C2(n3537), .A(n3667), .B(n3668), .ZN(n3541)
         );
  OAI21_X1 U4300 ( .B1(n3541), .B2(n3540), .A(n3539), .ZN(n3542) );
  NAND2_X1 U4301 ( .A1(n3542), .A2(n3673), .ZN(n3547) );
  NAND2_X1 U4302 ( .A1(n3803), .A2(n3543), .ZN(n3545) );
  AOI21_X1 U4303 ( .B1(n3547), .B2(n3674), .A(n3546), .ZN(n3551) );
  INV_X1 U4304 ( .A(n3548), .ZN(n3735) );
  INV_X1 U4305 ( .A(n3549), .ZN(n3678) );
  OAI211_X1 U4306 ( .C1(n3551), .C2(n3735), .A(n3678), .B(n3550), .ZN(n3552)
         );
  OAI21_X1 U4307 ( .B1(n3554), .B2(n3553), .A(n3552), .ZN(n3555) );
  OAI21_X1 U4308 ( .B1(n3557), .B2(n3556), .A(n3555), .ZN(n3562) );
  OAI21_X1 U4309 ( .B1(n3560), .B2(n3559), .A(n3558), .ZN(n3561) );
  NAND2_X1 U4310 ( .A1(n3562), .A2(n3561), .ZN(n3563) );
  MUX2_X1 U4311 ( .A(n3564), .B(n3563), .S(n4270), .Z(n3565) );
  MUX2_X1 U4312 ( .A(n3566), .B(n3565), .S(n4271), .Z(n3567) );
  XNOR2_X1 U4313 ( .A(n3567), .B(n3624), .ZN(n3573) );
  NOR2_X1 U4314 ( .A1(n3569), .A2(n3568), .ZN(n3571) );
  OAI21_X1 U4315 ( .B1(n3572), .B2(n4269), .A(B_REG_SCAN_IN), .ZN(n3570) );
  OAI22_X1 U4316 ( .A1(n3573), .A2(n3572), .B1(n3571), .B2(n3570), .ZN(U3239)
         );
  MUX2_X1 U4317 ( .A(n3705), .B(DATAO_REG_29__SCAN_IN), .S(n3583), .Z(U3579)
         );
  MUX2_X1 U4318 ( .A(n3728), .B(DATAO_REG_28__SCAN_IN), .S(n3583), .Z(U3578)
         );
  MUX2_X1 U4319 ( .A(n3738), .B(DATAO_REG_27__SCAN_IN), .S(n3583), .Z(U3577)
         );
  MUX2_X1 U4320 ( .A(n3762), .B(DATAO_REG_26__SCAN_IN), .S(n3583), .Z(U3576)
         );
  MUX2_X1 U4321 ( .A(n3737), .B(DATAO_REG_25__SCAN_IN), .S(n3583), .Z(U3575)
         );
  MUX2_X1 U4322 ( .A(n3806), .B(DATAO_REG_24__SCAN_IN), .S(n3583), .Z(U3574)
         );
  MUX2_X1 U4323 ( .A(n3780), .B(DATAO_REG_23__SCAN_IN), .S(n3583), .Z(U3573)
         );
  MUX2_X1 U4324 ( .A(n3836), .B(DATAO_REG_22__SCAN_IN), .S(n3583), .Z(U3572)
         );
  MUX2_X1 U4325 ( .A(n3855), .B(DATAO_REG_21__SCAN_IN), .S(n3583), .Z(U3571)
         );
  MUX2_X1 U4326 ( .A(n3878), .B(DATAO_REG_20__SCAN_IN), .S(n3583), .Z(U3570)
         );
  MUX2_X1 U4327 ( .A(n3891), .B(DATAO_REG_19__SCAN_IN), .S(n3583), .Z(U3569)
         );
  MUX2_X1 U4328 ( .A(n3909), .B(DATAO_REG_18__SCAN_IN), .S(n3583), .Z(U3568)
         );
  MUX2_X1 U4329 ( .A(n3926), .B(DATAO_REG_17__SCAN_IN), .S(n3583), .Z(U3567)
         );
  MUX2_X1 U4330 ( .A(n3947), .B(DATAO_REG_16__SCAN_IN), .S(n3583), .Z(U3566)
         );
  MUX2_X1 U4331 ( .A(n3970), .B(DATAO_REG_15__SCAN_IN), .S(n3583), .Z(U3565)
         );
  MUX2_X1 U4332 ( .A(n3574), .B(DATAO_REG_14__SCAN_IN), .S(n3583), .Z(U3564)
         );
  MUX2_X1 U4333 ( .A(n3627), .B(DATAO_REG_13__SCAN_IN), .S(n3583), .Z(U3563)
         );
  MUX2_X1 U4334 ( .A(n4445), .B(DATAO_REG_12__SCAN_IN), .S(n3583), .Z(U3562)
         );
  MUX2_X1 U4335 ( .A(n3575), .B(DATAO_REG_11__SCAN_IN), .S(n3583), .Z(U3561)
         );
  MUX2_X1 U4336 ( .A(n3576), .B(DATAO_REG_10__SCAN_IN), .S(n3583), .Z(U3560)
         );
  MUX2_X1 U4337 ( .A(n3577), .B(DATAO_REG_9__SCAN_IN), .S(n3583), .Z(U3559) );
  MUX2_X1 U4338 ( .A(n3578), .B(DATAO_REG_8__SCAN_IN), .S(n3583), .Z(U3558) );
  MUX2_X1 U4339 ( .A(n3579), .B(DATAO_REG_6__SCAN_IN), .S(n3583), .Z(U3556) );
  MUX2_X1 U4340 ( .A(n3580), .B(DATAO_REG_5__SCAN_IN), .S(n3583), .Z(U3555) );
  MUX2_X1 U4341 ( .A(n3581), .B(DATAO_REG_4__SCAN_IN), .S(n3583), .Z(U3554) );
  MUX2_X1 U4342 ( .A(n3582), .B(DATAO_REG_3__SCAN_IN), .S(n3583), .Z(U3553) );
  MUX2_X1 U4343 ( .A(n4480), .B(DATAO_REG_2__SCAN_IN), .S(n3583), .Z(U3552) );
  MUX2_X1 U4344 ( .A(n2304), .B(DATAO_REG_1__SCAN_IN), .S(n3583), .Z(U3551) );
  MUX2_X1 U4345 ( .A(n3584), .B(DATAO_REG_0__SCAN_IN), .S(n3583), .Z(U3550) );
  AOI22_X1 U4346 ( .A1(n4436), .A2(ADDR_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n3592) );
  AOI21_X1 U4347 ( .B1(n2314), .B2(n3585), .A(n3587), .ZN(n3586) );
  MUX2_X1 U4348 ( .A(n3587), .B(n3586), .S(n2158), .Z(n3589) );
  NAND2_X1 U4349 ( .A1(n3589), .A2(n3588), .ZN(n3591) );
  NAND3_X1 U4350 ( .A1(n4438), .A2(IR_REG_0__SCAN_IN), .A3(n2314), .ZN(n3590)
         );
  NAND3_X1 U4351 ( .A1(n3592), .A2(n3591), .A3(n3590), .ZN(U3240) );
  NAND2_X1 U4352 ( .A1(n3593), .A2(n4277), .ZN(n3605) );
  INV_X1 U4353 ( .A(n3594), .ZN(n3597) );
  OAI211_X1 U4354 ( .C1(n3597), .C2(n3596), .A(n4388), .B(n3595), .ZN(n3604)
         );
  OAI211_X1 U4355 ( .C1(n3600), .C2(n3599), .A(n4438), .B(n3598), .ZN(n3603)
         );
  NOR2_X1 U4356 ( .A1(STATE_REG_SCAN_IN), .A2(n2297), .ZN(n3601) );
  AOI21_X1 U4357 ( .B1(n4436), .B2(ADDR_REG_1__SCAN_IN), .A(n3601), .ZN(n3602)
         );
  NAND4_X1 U4358 ( .A1(n3605), .A2(n3604), .A3(n3603), .A4(n3602), .ZN(U3241)
         );
  INV_X1 U4359 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3611) );
  INV_X1 U4360 ( .A(n3620), .ZN(n4530) );
  AOI22_X1 U4361 ( .A1(n3620), .A2(REG1_REG_18__SCAN_IN), .B1(n3611), .B2(
        n4530), .ZN(n4440) );
  INV_X1 U4362 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4191) );
  INV_X1 U4363 ( .A(n4531), .ZN(n4429) );
  INV_X1 U4364 ( .A(n3616), .ZN(n4536) );
  INV_X1 U4365 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4199) );
  AOI22_X1 U4366 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3616), .B1(n4536), .B2(
        n4199), .ZN(n4407) );
  NAND2_X1 U4367 ( .A1(n3606), .A2(n4273), .ZN(n3608) );
  NOR2_X1 U4368 ( .A1(n3617), .A2(n3609), .ZN(n3610) );
  AOI22_X1 U4369 ( .A1(REG1_REG_17__SCAN_IN), .A2(n4429), .B1(n4531), .B2(
        n4191), .ZN(n4424) );
  OAI21_X1 U4370 ( .B1(n3611), .B2(n4530), .A(n4437), .ZN(n3613) );
  XNOR2_X1 U4371 ( .A(n3624), .B(REG1_REG_19__SCAN_IN), .ZN(n3612) );
  AOI22_X1 U4372 ( .A1(n3620), .A2(n3899), .B1(REG2_REG_18__SCAN_IN), .B2(
        n4530), .ZN(n4433) );
  AOI22_X1 U4373 ( .A1(REG2_REG_17__SCAN_IN), .A2(n4531), .B1(n4429), .B2(
        n3918), .ZN(n4421) );
  AOI22_X1 U4374 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4536), .B1(n3616), .B2(
        n3962), .ZN(n4401) );
  NOR2_X1 U4375 ( .A1(n4402), .A2(n4401), .ZN(n4400) );
  INV_X1 U4376 ( .A(n3617), .ZN(n4534) );
  NAND2_X1 U4377 ( .A1(n3618), .A2(n4534), .ZN(n3619) );
  NAND2_X1 U4378 ( .A1(n4421), .A2(n4419), .ZN(n4420) );
  OAI21_X1 U4379 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4531), .A(n4420), .ZN(n4432) );
  NOR2_X1 U4380 ( .A1(n4433), .A2(n4432), .ZN(n4431) );
  XNOR2_X1 U4381 ( .A(n3624), .B(REG2_REG_19__SCAN_IN), .ZN(n3621) );
  NAND2_X1 U4382 ( .A1(n4436), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3622) );
  OAI211_X1 U4383 ( .C1(n4443), .C2(n3624), .A(n3623), .B(n3622), .ZN(n3625)
         );
  AND2_X1 U4384 ( .A1(n3627), .A2(n3626), .ZN(n3950) );
  NAND2_X1 U4385 ( .A1(n3970), .A2(n4285), .ZN(n3632) );
  INV_X1 U4386 ( .A(n3632), .ZN(n3631) );
  OR2_X1 U4387 ( .A1(n3970), .A2(n4285), .ZN(n3629) );
  NAND2_X1 U4388 ( .A1(n4279), .A2(n3628), .ZN(n3955) );
  AND2_X1 U4389 ( .A1(n3629), .A2(n3955), .ZN(n3630) );
  INV_X1 U4390 ( .A(n3637), .ZN(n3634) );
  AND2_X1 U4391 ( .A1(n3954), .A2(n3632), .ZN(n3633) );
  NOR2_X1 U4392 ( .A1(n3634), .A2(n3633), .ZN(n3639) );
  OR2_X1 U4393 ( .A1(n3950), .A2(n3639), .ZN(n3635) );
  NOR2_X1 U4394 ( .A1(n3951), .A2(n3635), .ZN(n3641) );
  NAND2_X1 U4395 ( .A1(n3972), .A2(n3636), .ZN(n3952) );
  AND2_X1 U4396 ( .A1(n3952), .A2(n3637), .ZN(n3638) );
  NOR2_X1 U4397 ( .A1(n3639), .A2(n3638), .ZN(n3640) );
  NAND2_X1 U4398 ( .A1(n3926), .A2(n3642), .ZN(n3643) );
  NOR2_X1 U4399 ( .A1(n3891), .A2(n3882), .ZN(n3645) );
  OAI21_X1 U4400 ( .B1(n3847), .B2(n3647), .A(n3646), .ZN(n3831) );
  NOR2_X1 U4401 ( .A1(n3855), .A2(n3835), .ZN(n3649) );
  NAND2_X1 U4402 ( .A1(n3855), .A2(n3835), .ZN(n3648) );
  NAND2_X1 U4403 ( .A1(n3823), .A2(n3809), .ZN(n3650) );
  NAND3_X1 U4404 ( .A1(n3792), .A2(n3650), .A3(n3816), .ZN(n3655) );
  INV_X1 U4405 ( .A(n3650), .ZN(n3652) );
  NAND2_X1 U4406 ( .A1(n3836), .A2(n3824), .ZN(n3793) );
  NAND2_X1 U4407 ( .A1(n3780), .A2(n3797), .ZN(n3651) );
  NAND2_X1 U4408 ( .A1(n3783), .A2(n3767), .ZN(n3657) );
  OAI21_X1 U4409 ( .B1(n3731), .B2(n3746), .A(n3743), .ZN(n3658) );
  OAI21_X1 U4410 ( .B1(n3659), .B2(n3762), .A(n3658), .ZN(n3718) );
  NOR2_X1 U4411 ( .A1(n3738), .A2(n3727), .ZN(n3661) );
  INV_X1 U4412 ( .A(n3701), .ZN(n3662) );
  AOI22_X1 U4413 ( .A1(n3700), .A2(n3662), .B1(n3728), .B2(n3704), .ZN(n3664)
         );
  INV_X1 U4414 ( .A(n3684), .ZN(n3663) );
  XNOR2_X1 U4415 ( .A(n3664), .B(n3663), .ZN(n3992) );
  INV_X1 U4416 ( .A(n3992), .ZN(n3699) );
  NAND2_X1 U4417 ( .A1(n3969), .A2(n3973), .ZN(n3968) );
  INV_X1 U4418 ( .A(n3668), .ZN(n3669) );
  INV_X1 U4419 ( .A(n3670), .ZN(n3671) );
  INV_X1 U4420 ( .A(n3673), .ZN(n3675) );
  INV_X1 U4421 ( .A(n3680), .ZN(n3681) );
  AOI21_X1 U4422 ( .B1(n3702), .B2(n3682), .A(n3681), .ZN(n3683) );
  XOR2_X1 U4423 ( .A(n3684), .B(n3683), .Z(n3691) );
  AOI22_X1 U4424 ( .A1(n3687), .A2(n3686), .B1(n4478), .B2(n3685), .ZN(n3688)
         );
  OAI21_X1 U4425 ( .B1(n3689), .B2(n4482), .A(n3688), .ZN(n3690) );
  OAI21_X1 U4426 ( .B1(n4515), .B2(n3692), .A(n3994), .ZN(n3697) );
  OAI22_X1 U4427 ( .A1(n3993), .A2(n3961), .B1(n3695), .B2(n4511), .ZN(n3696)
         );
  AOI21_X1 U4428 ( .B1(n3697), .B2(n4511), .A(n3696), .ZN(n3698) );
  OAI21_X1 U4429 ( .B1(n3699), .B2(n3902), .A(n3698), .ZN(U3354) );
  XNOR2_X1 U4430 ( .A(n3700), .B(n3701), .ZN(n3996) );
  INV_X1 U4431 ( .A(n3996), .ZN(n3717) );
  XNOR2_X1 U4432 ( .A(n3702), .B(n3701), .ZN(n3703) );
  NAND2_X1 U4433 ( .A1(n3703), .A2(n4502), .ZN(n3707) );
  AOI22_X1 U4434 ( .A1(n3705), .A2(n4479), .B1(n4478), .B2(n3704), .ZN(n3706)
         );
  OAI211_X1 U4435 ( .C1(n3708), .C2(n4482), .A(n3707), .B(n3706), .ZN(n3995)
         );
  INV_X1 U4436 ( .A(n3709), .ZN(n3719) );
  INV_X1 U4437 ( .A(n3710), .ZN(n3711) );
  AOI22_X1 U4438 ( .A1(n4296), .A2(REG2_REG_28__SCAN_IN), .B1(n4491), .B2(
        n3713), .ZN(n3714) );
  OAI21_X1 U4439 ( .B1(n4218), .B2(n3961), .A(n3714), .ZN(n3715) );
  AOI21_X1 U4440 ( .B1(n3995), .B2(n4511), .A(n3715), .ZN(n3716) );
  OAI21_X1 U4441 ( .B1(n3717), .B2(n3902), .A(n3716), .ZN(U3262) );
  XNOR2_X1 U4442 ( .A(n3718), .B(n3724), .ZN(n4002) );
  AOI21_X1 U4443 ( .B1(n3727), .B2(n3745), .A(n3719), .ZN(n4000) );
  OAI22_X1 U4444 ( .A1(n4511), .A2(n3721), .B1(n3720), .B2(n4515), .ZN(n3722)
         );
  AOI21_X1 U4445 ( .B1(n4000), .B2(n4498), .A(n3722), .ZN(n3733) );
  OAI21_X1 U4446 ( .B1(n3725), .B2(n3724), .A(n3723), .ZN(n3726) );
  NAND2_X1 U4447 ( .A1(n3726), .A2(n4502), .ZN(n3730) );
  AOI22_X1 U4448 ( .A1(n3728), .A2(n4479), .B1(n3727), .B2(n4478), .ZN(n3729)
         );
  OAI211_X1 U4449 ( .C1(n3731), .C2(n4482), .A(n3730), .B(n3729), .ZN(n3999)
         );
  NAND2_X1 U4450 ( .A1(n3999), .A2(n4511), .ZN(n3732) );
  OAI211_X1 U4451 ( .C1(n4002), .C2(n3902), .A(n3733), .B(n3732), .ZN(U3263)
         );
  OAI21_X1 U4452 ( .B1(n3755), .B2(n3735), .A(n3734), .ZN(n3736) );
  XNOR2_X1 U4453 ( .A(n3736), .B(n3744), .ZN(n3742) );
  NAND2_X1 U4454 ( .A1(n3737), .A2(n3925), .ZN(n3740) );
  NAND2_X1 U4455 ( .A1(n3738), .A2(n4479), .ZN(n3739) );
  OAI211_X1 U4456 ( .C1(n3930), .C2(n3746), .A(n3740), .B(n3739), .ZN(n3741)
         );
  AOI21_X1 U4457 ( .B1(n3742), .B2(n4502), .A(n3741), .ZN(n4004) );
  XOR2_X1 U4458 ( .A(n3744), .B(n3743), .Z(n4003) );
  NAND2_X1 U4459 ( .A1(n4003), .A2(n3965), .ZN(n3753) );
  INV_X1 U4460 ( .A(n3766), .ZN(n3747) );
  OAI21_X1 U4461 ( .B1(n3747), .B2(n3746), .A(n3745), .ZN(n4006) );
  INV_X1 U4462 ( .A(n4006), .ZN(n3751) );
  OAI22_X1 U4463 ( .A1(n4511), .A2(n3749), .B1(n3748), .B2(n4515), .ZN(n3750)
         );
  AOI21_X1 U4464 ( .B1(n3751), .B2(n4498), .A(n3750), .ZN(n3752) );
  OAI211_X1 U4465 ( .C1(n4296), .C2(n4004), .A(n3753), .B(n3752), .ZN(U3264)
         );
  XOR2_X1 U4466 ( .A(n3758), .B(n3754), .Z(n4154) );
  INV_X1 U4467 ( .A(n4154), .ZN(n3772) );
  INV_X1 U4468 ( .A(n3755), .ZN(n3757) );
  NAND2_X1 U4469 ( .A1(n3757), .A2(n3756), .ZN(n3759) );
  XNOR2_X1 U4470 ( .A(n3759), .B(n3758), .ZN(n3760) );
  NAND2_X1 U4471 ( .A1(n3760), .A2(n4502), .ZN(n3764) );
  NOR2_X1 U4472 ( .A1(n3767), .A2(n3930), .ZN(n3761) );
  AOI21_X1 U4473 ( .B1(n3762), .B2(n4479), .A(n3761), .ZN(n3763) );
  OAI211_X1 U4474 ( .C1(n3765), .C2(n4482), .A(n3764), .B(n3763), .ZN(n4153)
         );
  OAI21_X1 U4475 ( .B1(n3784), .B2(n3767), .A(n3766), .ZN(n4224) );
  AOI22_X1 U4476 ( .A1(n4296), .A2(REG2_REG_25__SCAN_IN), .B1(n3768), .B2(
        n4491), .ZN(n3769) );
  OAI21_X1 U4477 ( .B1(n4224), .B2(n3961), .A(n3769), .ZN(n3770) );
  AOI21_X1 U4478 ( .B1(n4153), .B2(n4511), .A(n3770), .ZN(n3771) );
  OAI21_X1 U4479 ( .B1(n3772), .B2(n3902), .A(n3771), .ZN(U3265) );
  XOR2_X1 U4480 ( .A(n3777), .B(n3773), .Z(n4158) );
  INV_X1 U4481 ( .A(n4158), .ZN(n3791) );
  NAND2_X1 U4482 ( .A1(n3775), .A2(n3774), .ZN(n3776) );
  XOR2_X1 U4483 ( .A(n3777), .B(n3776), .Z(n3778) );
  NAND2_X1 U4484 ( .A1(n3778), .A2(n4502), .ZN(n3782) );
  AOI22_X1 U4485 ( .A1(n3780), .A2(n3925), .B1(n4478), .B2(n3779), .ZN(n3781)
         );
  OAI211_X1 U4486 ( .C1(n3783), .C2(n4505), .A(n3782), .B(n3781), .ZN(n4157)
         );
  INV_X1 U4487 ( .A(n3784), .ZN(n3785) );
  OAI21_X1 U4488 ( .B1(n3796), .B2(n3786), .A(n3785), .ZN(n4228) );
  AOI22_X1 U4489 ( .A1(n4296), .A2(REG2_REG_24__SCAN_IN), .B1(n3787), .B2(
        n4491), .ZN(n3788) );
  OAI21_X1 U4490 ( .B1(n4228), .B2(n3961), .A(n3788), .ZN(n3789) );
  AOI21_X1 U4491 ( .B1(n4157), .B2(n4511), .A(n3789), .ZN(n3790) );
  OAI21_X1 U4492 ( .B1(n3791), .B2(n3902), .A(n3790), .ZN(U3266) );
  NAND2_X1 U4493 ( .A1(n3792), .A2(n3816), .ZN(n3815) );
  NAND2_X1 U4494 ( .A1(n3815), .A2(n3793), .ZN(n3795) );
  XNOR2_X1 U4495 ( .A(n3795), .B(n3794), .ZN(n4162) );
  AOI21_X1 U4496 ( .B1(n3797), .B2(n4168), .A(n3796), .ZN(n4232) );
  OAI22_X1 U4497 ( .A1(n4511), .A2(n3799), .B1(n3798), .B2(n4515), .ZN(n3813)
         );
  NAND2_X1 U4498 ( .A1(n3832), .A2(n3800), .ZN(n3802) );
  NAND2_X1 U4499 ( .A1(n3802), .A2(n3801), .ZN(n3818) );
  NAND2_X1 U4500 ( .A1(n3818), .A2(n3819), .ZN(n3817) );
  NAND2_X1 U4501 ( .A1(n3817), .A2(n3803), .ZN(n3805) );
  XNOR2_X1 U4502 ( .A(n3805), .B(n3804), .ZN(n3811) );
  NAND2_X1 U4503 ( .A1(n3806), .A2(n4479), .ZN(n3808) );
  NAND2_X1 U4504 ( .A1(n3836), .A2(n3925), .ZN(n3807) );
  OAI211_X1 U4505 ( .C1(n3930), .C2(n3809), .A(n3808), .B(n3807), .ZN(n3810)
         );
  AOI21_X1 U4506 ( .B1(n3811), .B2(n4502), .A(n3810), .ZN(n4161) );
  NOR2_X1 U4507 ( .A1(n4161), .A2(n4296), .ZN(n3812) );
  AOI211_X1 U4508 ( .C1(n4232), .C2(n4498), .A(n3813), .B(n3812), .ZN(n3814)
         );
  OAI21_X1 U4509 ( .B1(n4162), .B2(n3902), .A(n3814), .ZN(U3267) );
  OAI21_X1 U4510 ( .B1(n3792), .B2(n3816), .A(n3815), .ZN(n4171) );
  OAI21_X1 U4511 ( .B1(n3819), .B2(n3818), .A(n3817), .ZN(n3820) );
  NAND2_X1 U4512 ( .A1(n3820), .A2(n4502), .ZN(n3822) );
  AOI22_X1 U4513 ( .A1(n3855), .A2(n3925), .B1(n3824), .B2(n4478), .ZN(n3821)
         );
  OAI211_X1 U4514 ( .C1(n3823), .C2(n4505), .A(n3822), .B(n3821), .ZN(n4167)
         );
  AND2_X1 U4515 ( .A1(n3840), .A2(n3824), .ZN(n4166) );
  INV_X1 U4516 ( .A(n4166), .ZN(n3825) );
  NAND3_X1 U4517 ( .A1(n3825), .A2(n4498), .A3(n4168), .ZN(n3828) );
  AOI22_X1 U4518 ( .A1(n4296), .A2(REG2_REG_22__SCAN_IN), .B1(n3826), .B2(
        n4491), .ZN(n3827) );
  NAND2_X1 U4519 ( .A1(n3828), .A2(n3827), .ZN(n3829) );
  AOI21_X1 U4520 ( .B1(n4167), .B2(n4511), .A(n3829), .ZN(n3830) );
  OAI21_X1 U4521 ( .B1(n4171), .B2(n3902), .A(n3830), .ZN(U3268) );
  XNOR2_X1 U4522 ( .A(n3831), .B(n3833), .ZN(n4173) );
  INV_X1 U4523 ( .A(n4173), .ZN(n3846) );
  XOR2_X1 U4524 ( .A(n3833), .B(n3832), .Z(n3834) );
  NAND2_X1 U4525 ( .A1(n3834), .A2(n4502), .ZN(n3838) );
  AOI22_X1 U4526 ( .A1(n3836), .A2(n4479), .B1(n4478), .B2(n3835), .ZN(n3837)
         );
  OAI211_X1 U4527 ( .C1(n3839), .C2(n4482), .A(n3838), .B(n3837), .ZN(n4172)
         );
  OAI21_X1 U4528 ( .B1(n3859), .B2(n3841), .A(n3840), .ZN(n4238) );
  AOI22_X1 U4529 ( .A1(n4296), .A2(REG2_REG_21__SCAN_IN), .B1(n3842), .B2(
        n4491), .ZN(n3843) );
  OAI21_X1 U4530 ( .B1(n4238), .B2(n3961), .A(n3843), .ZN(n3844) );
  AOI21_X1 U4531 ( .B1(n4172), .B2(n4511), .A(n3844), .ZN(n3845) );
  OAI21_X1 U4532 ( .B1(n3846), .B2(n3902), .A(n3845), .ZN(U3269) );
  XNOR2_X1 U4533 ( .A(n3847), .B(n3851), .ZN(n4177) );
  INV_X1 U4534 ( .A(n4177), .ZN(n3866) );
  INV_X1 U4535 ( .A(n3848), .ZN(n3849) );
  NAND2_X1 U4536 ( .A1(n3850), .A2(n3849), .ZN(n3852) );
  XNOR2_X1 U4537 ( .A(n3852), .B(n3851), .ZN(n3853) );
  NAND2_X1 U4538 ( .A1(n3853), .A2(n4502), .ZN(n3857) );
  NOR2_X1 U4539 ( .A1(n3861), .A2(n3930), .ZN(n3854) );
  AOI21_X1 U4540 ( .B1(n3855), .B2(n4479), .A(n3854), .ZN(n3856) );
  OAI211_X1 U4541 ( .C1(n3858), .C2(n4482), .A(n3857), .B(n3856), .ZN(n4176)
         );
  INV_X1 U4542 ( .A(n3859), .ZN(n3860) );
  OAI21_X1 U4543 ( .B1(n3883), .B2(n3861), .A(n3860), .ZN(n4242) );
  AOI22_X1 U4544 ( .A1(n4296), .A2(REG2_REG_20__SCAN_IN), .B1(n3862), .B2(
        n4491), .ZN(n3863) );
  OAI21_X1 U4545 ( .B1(n4242), .B2(n3961), .A(n3863), .ZN(n3864) );
  AOI21_X1 U4546 ( .B1(n4176), .B2(n4511), .A(n3864), .ZN(n3865) );
  OAI21_X1 U4547 ( .B1(n3866), .B2(n3902), .A(n3865), .ZN(U3270) );
  XNOR2_X1 U4548 ( .A(n3868), .B(n3867), .ZN(n4181) );
  INV_X1 U4549 ( .A(n4181), .ZN(n3889) );
  INV_X1 U4550 ( .A(n3869), .ZN(n3870) );
  AOI21_X1 U4551 ( .B1(n3908), .B2(n3871), .A(n3870), .ZN(n3890) );
  INV_X1 U4552 ( .A(n3872), .ZN(n3873) );
  AOI21_X1 U4553 ( .B1(n3890), .B2(n3874), .A(n3873), .ZN(n3876) );
  XNOR2_X1 U4554 ( .A(n3876), .B(n3875), .ZN(n3877) );
  NAND2_X1 U4555 ( .A1(n3877), .A2(n4502), .ZN(n3880) );
  AOI22_X1 U4556 ( .A1(n3878), .A2(n4479), .B1(n3882), .B2(n4478), .ZN(n3879)
         );
  OAI211_X1 U4557 ( .C1(n3881), .C2(n4482), .A(n3880), .B(n3879), .ZN(n4180)
         );
  AND2_X1 U4558 ( .A1(n2070), .A2(n3882), .ZN(n3884) );
  OR2_X1 U4559 ( .A1(n3884), .A2(n3883), .ZN(n4246) );
  AOI22_X1 U4560 ( .A1(n4296), .A2(REG2_REG_19__SCAN_IN), .B1(n3885), .B2(
        n4491), .ZN(n3886) );
  OAI21_X1 U4561 ( .B1(n4246), .B2(n3961), .A(n3886), .ZN(n3887) );
  AOI21_X1 U4562 ( .B1(n4180), .B2(n4511), .A(n3887), .ZN(n3888) );
  OAI21_X1 U4563 ( .B1(n3889), .B2(n3902), .A(n3888), .ZN(U3271) );
  XOR2_X1 U4564 ( .A(n3901), .B(n3890), .Z(n3895) );
  AOI22_X1 U4565 ( .A1(n3891), .A2(n4479), .B1(n3896), .B2(n4478), .ZN(n3892)
         );
  OAI21_X1 U4566 ( .B1(n3893), .B2(n4482), .A(n3892), .ZN(n3894) );
  AOI21_X1 U4567 ( .B1(n3895), .B2(n4502), .A(n3894), .ZN(n4185) );
  AOI21_X1 U4568 ( .B1(n2068), .B2(n3896), .A(n4591), .ZN(n3897) );
  NAND2_X1 U4569 ( .A1(n3897), .A2(n2070), .ZN(n4184) );
  INV_X1 U4570 ( .A(n4184), .ZN(n3906) );
  OAI22_X1 U4571 ( .A1(n4511), .A2(n3899), .B1(n3898), .B2(n4515), .ZN(n3904)
         );
  XOR2_X1 U4572 ( .A(n3901), .B(n3900), .Z(n4187) );
  NOR2_X1 U4573 ( .A1(n4187), .A2(n3902), .ZN(n3903) );
  AOI211_X1 U4574 ( .C1(n3906), .C2(n3905), .A(n3904), .B(n3903), .ZN(n3907)
         );
  OAI21_X1 U4575 ( .B1(n4296), .B2(n4185), .A(n3907), .ZN(U3272) );
  XNOR2_X1 U4576 ( .A(n3908), .B(n3914), .ZN(n3913) );
  NAND2_X1 U4577 ( .A1(n3947), .A2(n3925), .ZN(n3911) );
  NAND2_X1 U4578 ( .A1(n3909), .A2(n4479), .ZN(n3910) );
  OAI211_X1 U4579 ( .C1(n3930), .C2(n3916), .A(n3911), .B(n3910), .ZN(n3912)
         );
  AOI21_X1 U4580 ( .B1(n3913), .B2(n4502), .A(n3912), .ZN(n4189) );
  INV_X1 U4581 ( .A(n3914), .ZN(n3915) );
  XNOR2_X1 U4582 ( .A(n2077), .B(n3915), .ZN(n4188) );
  OAI21_X1 U4583 ( .B1(n3937), .B2(n3916), .A(n2068), .ZN(n4251) );
  NOR2_X1 U4584 ( .A1(n4251), .A2(n3961), .ZN(n3920) );
  OAI22_X1 U4585 ( .A1(n4511), .A2(n3918), .B1(n3917), .B2(n4515), .ZN(n3919)
         );
  AOI211_X1 U4586 ( .C1(n4188), .C2(n3965), .A(n3920), .B(n3919), .ZN(n3921)
         );
  OAI21_X1 U4587 ( .B1(n4296), .B2(n4189), .A(n3921), .ZN(U3273) );
  XNOR2_X1 U4588 ( .A(n3923), .B(n3922), .ZN(n3924) );
  NAND2_X1 U4589 ( .A1(n3924), .A2(n4502), .ZN(n3933) );
  NAND2_X1 U4590 ( .A1(n3970), .A2(n3925), .ZN(n3928) );
  NAND2_X1 U4591 ( .A1(n3926), .A2(n4479), .ZN(n3927) );
  OAI211_X1 U4592 ( .C1(n3930), .C2(n3929), .A(n3928), .B(n3927), .ZN(n3931)
         );
  INV_X1 U4593 ( .A(n3931), .ZN(n3932) );
  NAND2_X1 U4594 ( .A1(n3933), .A2(n3932), .ZN(n4193) );
  INV_X1 U4595 ( .A(n4193), .ZN(n3943) );
  XNOR2_X1 U4596 ( .A(n3934), .B(n3935), .ZN(n4194) );
  AND2_X1 U4597 ( .A1(n3960), .A2(n3936), .ZN(n3938) );
  OR2_X1 U4598 ( .A1(n3938), .A2(n3937), .ZN(n4255) );
  AOI22_X1 U4599 ( .A1(n4296), .A2(REG2_REG_16__SCAN_IN), .B1(n3939), .B2(
        n4491), .ZN(n3940) );
  OAI21_X1 U4600 ( .B1(n4255), .B2(n3961), .A(n3940), .ZN(n3941) );
  AOI21_X1 U4601 ( .B1(n4194), .B2(n3965), .A(n3941), .ZN(n3942) );
  OAI21_X1 U4602 ( .B1(n4296), .B2(n3943), .A(n3942), .ZN(U3274) );
  XNOR2_X1 U4603 ( .A(n3945), .B(n3944), .ZN(n3946) );
  NAND2_X1 U4604 ( .A1(n3946), .A2(n4502), .ZN(n3949) );
  AOI22_X1 U4605 ( .A1(n3947), .A2(n4479), .B1(n4285), .B2(n4478), .ZN(n3948)
         );
  OAI211_X1 U4606 ( .C1(n4279), .C2(n4482), .A(n3949), .B(n3948), .ZN(n4197)
         );
  INV_X1 U4607 ( .A(n4197), .ZN(n3967) );
  OR2_X1 U4608 ( .A1(n3951), .A2(n3950), .ZN(n3953) );
  NAND2_X1 U4609 ( .A1(n3953), .A2(n3952), .ZN(n3974) );
  NAND2_X1 U4610 ( .A1(n3974), .A2(n3954), .ZN(n3956) );
  NAND2_X1 U4611 ( .A1(n3956), .A2(n3955), .ZN(n3958) );
  XNOR2_X1 U4612 ( .A(n3958), .B(n3957), .ZN(n4198) );
  NAND2_X1 U4613 ( .A1(n4203), .A2(n4285), .ZN(n3959) );
  NAND2_X1 U4614 ( .A1(n3960), .A2(n3959), .ZN(n4260) );
  NOR2_X1 U4615 ( .A1(n4260), .A2(n3961), .ZN(n3964) );
  OAI22_X1 U4616 ( .A1(n4511), .A2(n3962), .B1(n4294), .B2(n4515), .ZN(n3963)
         );
  AOI211_X1 U4617 ( .C1(n4198), .C2(n3965), .A(n3964), .B(n3963), .ZN(n3966)
         );
  OAI21_X1 U4618 ( .B1(n4296), .B2(n3967), .A(n3966), .ZN(U3275) );
  OAI21_X1 U4619 ( .B1(n3973), .B2(n3969), .A(n3968), .ZN(n3977) );
  AOI22_X1 U4620 ( .A1(n3970), .A2(n4479), .B1(n4478), .B2(n3978), .ZN(n3971)
         );
  OAI21_X1 U4621 ( .B1(n3972), .B2(n4482), .A(n3971), .ZN(n3976) );
  XNOR2_X1 U4622 ( .A(n3974), .B(n3973), .ZN(n4206) );
  NOR2_X1 U4623 ( .A1(n4206), .A2(n4487), .ZN(n3975) );
  AOI211_X1 U4624 ( .C1(n4502), .C2(n3977), .A(n3976), .B(n3975), .ZN(n4205)
         );
  INV_X1 U4625 ( .A(n4206), .ZN(n3984) );
  NAND2_X1 U4626 ( .A1(n3979), .A2(n3978), .ZN(n4202) );
  AND3_X1 U4627 ( .A1(n4203), .A2(n4498), .A3(n4202), .ZN(n3983) );
  OAI22_X1 U4628 ( .A1(n4511), .A2(n3981), .B1(n3980), .B2(n4515), .ZN(n3982)
         );
  AOI211_X1 U4629 ( .C1(n3984), .C2(n4501), .A(n3983), .B(n3982), .ZN(n3985)
         );
  OAI21_X1 U4630 ( .B1(n4205), .B2(n4296), .A(n3985), .ZN(U3276) );
  AOI21_X1 U4631 ( .B1(n3989), .B2(n3987), .A(n3986), .ZN(n4300) );
  INV_X1 U4632 ( .A(n4300), .ZN(n4213) );
  INV_X1 U4633 ( .A(REG1_REG_30__SCAN_IN), .ZN(n3990) );
  AOI21_X1 U4634 ( .B1(n3989), .B2(n4478), .A(n3988), .ZN(n4302) );
  MUX2_X1 U4635 ( .A(n3990), .B(n4302), .S(n4624), .Z(n3991) );
  OAI21_X1 U4636 ( .B1(n4213), .B2(n4201), .A(n3991), .ZN(U3548) );
  MUX2_X1 U4637 ( .A(REG1_REG_29__SCAN_IN), .B(n4214), .S(n4624), .Z(U3547) );
  INV_X1 U4638 ( .A(REG1_REG_28__SCAN_IN), .ZN(n3997) );
  AOI21_X1 U4639 ( .B1(n3996), .B2(n4594), .A(n3995), .ZN(n4215) );
  OAI21_X1 U4640 ( .B1(n4218), .B2(n4201), .A(n3998), .ZN(U3546) );
  INV_X1 U4641 ( .A(n4594), .ZN(n4186) );
  AOI21_X1 U4642 ( .B1(n4602), .B2(n4000), .A(n3999), .ZN(n4001) );
  OAI21_X1 U4643 ( .B1(n4002), .B2(n4186), .A(n4001), .ZN(n4219) );
  MUX2_X1 U4644 ( .A(REG1_REG_27__SCAN_IN), .B(n4219), .S(n4624), .Z(U3545) );
  NAND2_X1 U4645 ( .A1(n4003), .A2(n4594), .ZN(n4005) );
  OAI211_X1 U4646 ( .C1(n4591), .C2(n4006), .A(n4005), .B(n4004), .ZN(n4220)
         );
  MUX2_X1 U4647 ( .A(REG1_REG_26__SCAN_IN), .B(n4220), .S(n4624), .Z(n4152) );
  NAND3_X1 U4648 ( .A1(keyinput5), .A2(keyinput8), .A3(keyinput17), .ZN(n4011)
         );
  INV_X1 U4649 ( .A(keyinput9), .ZN(n4007) );
  NAND4_X1 U4650 ( .A1(keyinput30), .A2(keyinput23), .A3(keyinput52), .A4(
        n4007), .ZN(n4010) );
  NOR4_X1 U4651 ( .A1(keyinput10), .A2(keyinput2), .A3(keyinput7), .A4(
        keyinput60), .ZN(n4008) );
  INV_X1 U4652 ( .A(keyinput55), .ZN(n4083) );
  NAND4_X1 U4653 ( .A1(keyinput25), .A2(keyinput59), .A3(n4008), .A4(n4083), 
        .ZN(n4009) );
  NOR4_X1 U4654 ( .A1(keyinput26), .A2(n4011), .A3(n4010), .A4(n4009), .ZN(
        n4026) );
  NAND2_X1 U4655 ( .A1(keyinput41), .A2(keyinput61), .ZN(n4014) );
  INV_X1 U4656 ( .A(keyinput45), .ZN(n4012) );
  NAND4_X1 U4657 ( .A1(keyinput4), .A2(keyinput3), .A3(keyinput42), .A4(n4012), 
        .ZN(n4013) );
  NOR4_X1 U4658 ( .A1(keyinput54), .A2(keyinput38), .A3(n4014), .A4(n4013), 
        .ZN(n4025) );
  NAND2_X1 U4659 ( .A1(keyinput57), .A2(keyinput37), .ZN(n4017) );
  NOR2_X1 U4660 ( .A1(keyinput21), .A2(keyinput48), .ZN(n4015) );
  NAND3_X1 U4661 ( .A1(keyinput1), .A2(keyinput39), .A3(n4015), .ZN(n4016) );
  NOR4_X1 U4662 ( .A1(keyinput36), .A2(keyinput14), .A3(n4017), .A4(n4016), 
        .ZN(n4024) );
  NAND3_X1 U4663 ( .A1(keyinput53), .A2(keyinput6), .A3(keyinput19), .ZN(n4022) );
  NAND4_X1 U4664 ( .A1(keyinput0), .A2(keyinput33), .A3(keyinput51), .A4(
        keyinput58), .ZN(n4021) );
  NOR3_X1 U4665 ( .A1(keyinput20), .A2(keyinput22), .A3(keyinput16), .ZN(n4019) );
  NOR3_X1 U4666 ( .A1(keyinput35), .A2(keyinput50), .A3(keyinput29), .ZN(n4018) );
  NAND4_X1 U4667 ( .A1(keyinput47), .A2(n4019), .A3(keyinput46), .A4(n4018), 
        .ZN(n4020) );
  NOR4_X1 U4668 ( .A1(keyinput31), .A2(n4022), .A3(n4021), .A4(n4020), .ZN(
        n4023) );
  NAND4_X1 U4669 ( .A1(n4026), .A2(n4025), .A3(n4024), .A4(n4023), .ZN(n4034)
         );
  NOR3_X1 U4670 ( .A1(keyinput32), .A2(keyinput49), .A3(keyinput12), .ZN(n4032) );
  NAND2_X1 U4671 ( .A1(keyinput11), .A2(keyinput56), .ZN(n4027) );
  NOR3_X1 U4672 ( .A1(keyinput28), .A2(keyinput44), .A3(n4027), .ZN(n4031) );
  NAND3_X1 U4673 ( .A1(keyinput18), .A2(keyinput40), .A3(keyinput34), .ZN(
        n4029) );
  NAND3_X1 U4674 ( .A1(keyinput13), .A2(keyinput24), .A3(keyinput43), .ZN(
        n4028) );
  NOR4_X1 U4675 ( .A1(keyinput27), .A2(keyinput15), .A3(n4029), .A4(n4028), 
        .ZN(n4030) );
  NAND4_X1 U4676 ( .A1(keyinput62), .A2(n4032), .A3(n4031), .A4(n4030), .ZN(
        n4033) );
  OAI21_X1 U4677 ( .B1(n4034), .B2(n4033), .A(keyinput63), .ZN(n4067) );
  INV_X1 U4678 ( .A(B_REG_SCAN_IN), .ZN(n4036) );
  AOI22_X1 U4679 ( .A1(n4037), .A2(keyinput9), .B1(n4036), .B2(keyinput23), 
        .ZN(n4035) );
  OAI221_X1 U4680 ( .B1(n4037), .B2(keyinput9), .C1(n4036), .C2(keyinput23), 
        .A(n4035), .ZN(n4048) );
  INV_X1 U4681 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4039) );
  AOI22_X1 U4682 ( .A1(n4040), .A2(keyinput52), .B1(keyinput10), .B2(n4039), 
        .ZN(n4038) );
  OAI221_X1 U4683 ( .B1(n4040), .B2(keyinput52), .C1(n4039), .C2(keyinput10), 
        .A(n4038), .ZN(n4047) );
  AOI22_X1 U4684 ( .A1(n2297), .A2(keyinput2), .B1(keyinput7), .B2(n2314), 
        .ZN(n4041) );
  OAI221_X1 U4685 ( .B1(n2297), .B2(keyinput2), .C1(n2314), .C2(keyinput7), 
        .A(n4041), .ZN(n4046) );
  INV_X1 U4686 ( .A(keyinput60), .ZN(n4044) );
  INV_X1 U4687 ( .A(keyinput32), .ZN(n4043) );
  AOI22_X1 U4688 ( .A1(n4044), .A2(ADDR_REG_2__SCAN_IN), .B1(
        ADDR_REG_4__SCAN_IN), .B2(n4043), .ZN(n4042) );
  OAI221_X1 U4689 ( .B1(n4044), .B2(ADDR_REG_2__SCAN_IN), .C1(n4043), .C2(
        ADDR_REG_4__SCAN_IN), .A(n4042), .ZN(n4045) );
  NOR4_X1 U4690 ( .A1(n4048), .A2(n4047), .A3(n4046), .A4(n4045), .ZN(n4065)
         );
  INV_X1 U4691 ( .A(keyinput24), .ZN(n4051) );
  INV_X1 U4692 ( .A(keyinput43), .ZN(n4050) );
  AOI22_X1 U4693 ( .A1(n4051), .A2(DATAO_REG_18__SCAN_IN), .B1(
        DATAO_REG_20__SCAN_IN), .B2(n4050), .ZN(n4049) );
  OAI221_X1 U4694 ( .B1(n4051), .B2(DATAO_REG_18__SCAN_IN), .C1(n4050), .C2(
        DATAO_REG_20__SCAN_IN), .A(n4049), .ZN(n4063) );
  INV_X1 U4695 ( .A(keyinput15), .ZN(n4054) );
  INV_X1 U4696 ( .A(keyinput28), .ZN(n4053) );
  AOI22_X1 U4697 ( .A1(n4054), .A2(DATAO_REG_25__SCAN_IN), .B1(
        DATAO_REG_28__SCAN_IN), .B2(n4053), .ZN(n4052) );
  OAI221_X1 U4698 ( .B1(n4054), .B2(DATAO_REG_25__SCAN_IN), .C1(n4053), .C2(
        DATAO_REG_28__SCAN_IN), .A(n4052), .ZN(n4062) );
  INV_X1 U4699 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4216) );
  INV_X1 U4700 ( .A(keyinput11), .ZN(n4056) );
  AOI22_X1 U4701 ( .A1(n4216), .A2(keyinput56), .B1(DATAO_REG_30__SCAN_IN), 
        .B2(n4056), .ZN(n4055) );
  OAI221_X1 U4702 ( .B1(n4216), .B2(keyinput56), .C1(n4056), .C2(
        DATAO_REG_30__SCAN_IN), .A(n4055), .ZN(n4061) );
  INV_X1 U4703 ( .A(keyinput44), .ZN(n4059) );
  INV_X1 U4704 ( .A(keyinput57), .ZN(n4058) );
  AOI22_X1 U4705 ( .A1(n4059), .A2(DATAO_REG_31__SCAN_IN), .B1(
        REG0_REG_31__SCAN_IN), .B2(n4058), .ZN(n4057) );
  OAI221_X1 U4706 ( .B1(n4059), .B2(DATAO_REG_31__SCAN_IN), .C1(n4058), .C2(
        REG0_REG_31__SCAN_IN), .A(n4057), .ZN(n4060) );
  NOR4_X1 U4707 ( .A1(n4063), .A2(n4062), .A3(n4061), .A4(n4060), .ZN(n4064)
         );
  NAND2_X1 U4708 ( .A1(n4065), .A2(n4064), .ZN(n4066) );
  AOI21_X1 U4709 ( .B1(DATAO_REG_7__SCAN_IN), .B2(n4067), .A(n4066), .ZN(n4150) );
  INV_X1 U4710 ( .A(keyinput49), .ZN(n4069) );
  AOI22_X1 U4711 ( .A1(n3011), .A2(keyinput62), .B1(ADDR_REG_6__SCAN_IN), .B2(
        n4069), .ZN(n4068) );
  OAI221_X1 U4712 ( .B1(n3011), .B2(keyinput62), .C1(n4069), .C2(
        ADDR_REG_6__SCAN_IN), .A(n4068), .ZN(n4079) );
  INV_X1 U4713 ( .A(keyinput27), .ZN(n4071) );
  AOI22_X1 U4714 ( .A1(n2435), .A2(keyinput12), .B1(ADDR_REG_12__SCAN_IN), 
        .B2(n4071), .ZN(n4070) );
  OAI221_X1 U4715 ( .B1(n2435), .B2(keyinput12), .C1(n4071), .C2(
        ADDR_REG_12__SCAN_IN), .A(n4070), .ZN(n4078) );
  INV_X1 U4716 ( .A(keyinput18), .ZN(n4074) );
  INV_X1 U4717 ( .A(keyinput40), .ZN(n4073) );
  AOI22_X1 U4718 ( .A1(n4074), .A2(ADDR_REG_14__SCAN_IN), .B1(
        ADDR_REG_17__SCAN_IN), .B2(n4073), .ZN(n4072) );
  OAI221_X1 U4719 ( .B1(n4074), .B2(ADDR_REG_14__SCAN_IN), .C1(n4073), .C2(
        ADDR_REG_17__SCAN_IN), .A(n4072), .ZN(n4077) );
  AOI22_X1 U4720 ( .A1(n3962), .A2(keyinput34), .B1(keyinput13), .B2(n2840), 
        .ZN(n4075) );
  OAI221_X1 U4721 ( .B1(n3962), .B2(keyinput34), .C1(n2840), .C2(keyinput13), 
        .A(n4075), .ZN(n4076) );
  NOR4_X1 U4722 ( .A1(n4079), .A2(n4078), .A3(n4077), .A4(n4076), .ZN(n4149)
         );
  AOI22_X1 U4723 ( .A1(keyinput25), .A2(U3149), .B1(keyinput63), .B2(n4080), 
        .ZN(n4081) );
  OAI21_X1 U4724 ( .B1(U3149), .B2(keyinput25), .A(n4081), .ZN(n4093) );
  AOI22_X1 U4725 ( .A1(n4611), .A2(keyinput5), .B1(DATAI_30_), .B2(n4083), 
        .ZN(n4082) );
  OAI221_X1 U4726 ( .B1(n4611), .B2(keyinput5), .C1(n4083), .C2(DATAI_30_), 
        .A(n4082), .ZN(n4092) );
  INV_X1 U4727 ( .A(keyinput26), .ZN(n4086) );
  INV_X1 U4728 ( .A(keyinput8), .ZN(n4085) );
  AOI22_X1 U4729 ( .A1(n4086), .A2(DATAO_REG_6__SCAN_IN), .B1(
        DATAO_REG_11__SCAN_IN), .B2(n4085), .ZN(n4084) );
  OAI221_X1 U4730 ( .B1(n4086), .B2(DATAO_REG_6__SCAN_IN), .C1(n4085), .C2(
        DATAO_REG_11__SCAN_IN), .A(n4084), .ZN(n4091) );
  INV_X1 U4731 ( .A(keyinput17), .ZN(n4088) );
  AOI22_X1 U4732 ( .A1(n4089), .A2(keyinput30), .B1(DATAO_REG_14__SCAN_IN), 
        .B2(n4088), .ZN(n4087) );
  OAI221_X1 U4733 ( .B1(n4089), .B2(keyinput30), .C1(n4088), .C2(
        DATAO_REG_14__SCAN_IN), .A(n4087), .ZN(n4090) );
  NOR4_X1 U4734 ( .A1(n4093), .A2(n4092), .A3(n4091), .A4(n4090), .ZN(n4148)
         );
  INV_X1 U4735 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4096) );
  INV_X1 U4736 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4095) );
  AOI22_X1 U4737 ( .A1(n4096), .A2(keyinput54), .B1(n4095), .B2(keyinput38), 
        .ZN(n4094) );
  OAI221_X1 U4738 ( .B1(n4096), .B2(keyinput54), .C1(n4095), .C2(keyinput38), 
        .A(n4094), .ZN(n4099) );
  INV_X1 U4739 ( .A(DATAI_15_), .ZN(n4535) );
  AOI22_X1 U4740 ( .A1(n4535), .A2(keyinput61), .B1(n2152), .B2(keyinput3), 
        .ZN(n4097) );
  OAI221_X1 U4741 ( .B1(n4535), .B2(keyinput61), .C1(n2152), .C2(keyinput3), 
        .A(n4097), .ZN(n4098) );
  NOR2_X1 U4742 ( .A1(n4099), .A2(n4098), .ZN(n4107) );
  INV_X1 U4743 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4101) );
  INV_X1 U4744 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4244) );
  AOI22_X1 U4745 ( .A1(n4101), .A2(keyinput37), .B1(n4244), .B2(keyinput36), 
        .ZN(n4100) );
  OAI221_X1 U4746 ( .B1(n4101), .B2(keyinput37), .C1(n4244), .C2(keyinput36), 
        .A(n4100), .ZN(n4105) );
  XNOR2_X1 U4747 ( .A(REG2_REG_26__SCAN_IN), .B(keyinput20), .ZN(n4103) );
  XNOR2_X1 U4748 ( .A(REG0_REG_27__SCAN_IN), .B(keyinput47), .ZN(n4102) );
  NAND2_X1 U4749 ( .A1(n4103), .A2(n4102), .ZN(n4104) );
  NOR2_X1 U4750 ( .A1(n4105), .A2(n4104), .ZN(n4106) );
  AND2_X1 U4751 ( .A1(n4107), .A2(n4106), .ZN(n4122) );
  INV_X1 U4752 ( .A(D_REG_11__SCAN_IN), .ZN(n4523) );
  INV_X1 U4753 ( .A(keyinput29), .ZN(n4108) );
  XNOR2_X1 U4754 ( .A(n4523), .B(n4108), .ZN(n4121) );
  INV_X1 U4755 ( .A(DATAI_5_), .ZN(n4551) );
  AOI22_X1 U4756 ( .A1(n4110), .A2(keyinput1), .B1(keyinput48), .B2(n4551), 
        .ZN(n4109) );
  OAI221_X1 U4757 ( .B1(n4110), .B2(keyinput1), .C1(n4551), .C2(keyinput48), 
        .A(n4109), .ZN(n4114) );
  INV_X1 U4758 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4595) );
  AOI22_X1 U4759 ( .A1(n4112), .A2(keyinput14), .B1(keyinput21), .B2(n4595), 
        .ZN(n4111) );
  OAI221_X1 U4760 ( .B1(n4112), .B2(keyinput14), .C1(n4595), .C2(keyinput21), 
        .A(n4111), .ZN(n4113) );
  NOR2_X1 U4761 ( .A1(n4114), .A2(n4113), .ZN(n4120) );
  INV_X1 U4762 ( .A(D_REG_9__SCAN_IN), .ZN(n4524) );
  INV_X1 U4763 ( .A(D_REG_19__SCAN_IN), .ZN(n4518) );
  AOI22_X1 U4764 ( .A1(n4524), .A2(keyinput31), .B1(keyinput35), .B2(n4518), 
        .ZN(n4115) );
  OAI221_X1 U4765 ( .B1(n4524), .B2(keyinput31), .C1(n4518), .C2(keyinput35), 
        .A(n4115), .ZN(n4118) );
  INV_X1 U4766 ( .A(D_REG_13__SCAN_IN), .ZN(n4521) );
  INV_X1 U4767 ( .A(D_REG_28__SCAN_IN), .ZN(n4516) );
  AOI22_X1 U4768 ( .A1(n4521), .A2(keyinput46), .B1(keyinput50), .B2(n4516), 
        .ZN(n4116) );
  OAI221_X1 U4769 ( .B1(n4521), .B2(keyinput46), .C1(n4516), .C2(keyinput50), 
        .A(n4116), .ZN(n4117) );
  NOR2_X1 U4770 ( .A1(n4118), .A2(n4117), .ZN(n4119) );
  NAND4_X1 U4771 ( .A1(n4122), .A2(n4121), .A3(n4120), .A4(n4119), .ZN(n4146)
         );
  INV_X1 U4772 ( .A(DATAI_0_), .ZN(n4124) );
  AOI22_X1 U4773 ( .A1(n4124), .A2(keyinput59), .B1(n2248), .B2(keyinput58), 
        .ZN(n4123) );
  OAI221_X1 U4774 ( .B1(n4124), .B2(keyinput59), .C1(n2248), .C2(keyinput58), 
        .A(n4123), .ZN(n4127) );
  INV_X1 U4775 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4178) );
  INV_X1 U4776 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4155) );
  AOI22_X1 U4777 ( .A1(n4178), .A2(keyinput4), .B1(keyinput42), .B2(n4155), 
        .ZN(n4125) );
  OAI221_X1 U4778 ( .B1(n4178), .B2(keyinput4), .C1(n4155), .C2(keyinput42), 
        .A(n4125), .ZN(n4126) );
  NOR2_X1 U4779 ( .A1(n4127), .A2(n4126), .ZN(n4144) );
  AOI22_X1 U4780 ( .A1(n4517), .A2(keyinput6), .B1(keyinput19), .B2(n4519), 
        .ZN(n4128) );
  OAI221_X1 U4781 ( .B1(n4517), .B2(keyinput6), .C1(n4519), .C2(keyinput19), 
        .A(n4128), .ZN(n4129) );
  INV_X1 U4782 ( .A(n4129), .ZN(n4143) );
  AOI22_X1 U4783 ( .A1(n4522), .A2(keyinput16), .B1(keyinput53), .B2(n4520), 
        .ZN(n4130) );
  OAI221_X1 U4784 ( .B1(n4522), .B2(keyinput16), .C1(n4520), .C2(keyinput53), 
        .A(n4130), .ZN(n4131) );
  INV_X1 U4785 ( .A(n4131), .ZN(n4142) );
  XNOR2_X1 U4786 ( .A(IR_REG_14__SCAN_IN), .B(keyinput33), .ZN(n4135) );
  XNOR2_X1 U4787 ( .A(IR_REG_23__SCAN_IN), .B(keyinput0), .ZN(n4134) );
  XNOR2_X1 U4788 ( .A(IR_REG_19__SCAN_IN), .B(keyinput22), .ZN(n4133) );
  XNOR2_X1 U4789 ( .A(IR_REG_28__SCAN_IN), .B(keyinput45), .ZN(n4132) );
  NAND4_X1 U4790 ( .A1(n4135), .A2(n4134), .A3(n4133), .A4(n4132), .ZN(n4140)
         );
  XNOR2_X1 U4791 ( .A(DATAI_16_), .B(keyinput51), .ZN(n4137) );
  XNOR2_X1 U4792 ( .A(keyinput39), .B(REG0_REG_0__SCAN_IN), .ZN(n4136) );
  NAND3_X1 U4793 ( .A1(n4138), .A2(n4137), .A3(n4136), .ZN(n4139) );
  NOR2_X1 U4794 ( .A1(n4140), .A2(n4139), .ZN(n4141) );
  NAND4_X1 U4795 ( .A1(n4144), .A2(n4143), .A3(n4142), .A4(n4141), .ZN(n4145)
         );
  NOR2_X1 U4796 ( .A1(n4146), .A2(n4145), .ZN(n4147) );
  NAND4_X1 U4797 ( .A1(n4150), .A2(n4149), .A3(n4148), .A4(n4147), .ZN(n4151)
         );
  XNOR2_X1 U4798 ( .A(n4152), .B(n4151), .ZN(U3544) );
  AOI21_X1 U4799 ( .B1(n4154), .B2(n4594), .A(n4153), .ZN(n4221) );
  MUX2_X1 U4800 ( .A(n4155), .B(n4221), .S(n4624), .Z(n4156) );
  OAI21_X1 U4801 ( .B1(n4201), .B2(n4224), .A(n4156), .ZN(U3543) );
  INV_X1 U4802 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4159) );
  AOI21_X1 U4803 ( .B1(n4158), .B2(n4594), .A(n4157), .ZN(n4225) );
  MUX2_X1 U4804 ( .A(n4159), .B(n4225), .S(n4624), .Z(n4160) );
  OAI21_X1 U4805 ( .B1(n4201), .B2(n4228), .A(n4160), .ZN(U3542) );
  INV_X1 U4806 ( .A(n4201), .ZN(n4164) );
  OAI21_X1 U4807 ( .B1(n4162), .B2(n4186), .A(n4161), .ZN(n4229) );
  MUX2_X1 U4808 ( .A(REG1_REG_23__SCAN_IN), .B(n4229), .S(n4624), .Z(n4163) );
  AOI21_X1 U4809 ( .B1(n4164), .B2(n4232), .A(n4163), .ZN(n4165) );
  INV_X1 U4810 ( .A(n4165), .ZN(U3541) );
  NOR2_X1 U4811 ( .A1(n4166), .A2(n4591), .ZN(n4169) );
  AOI21_X1 U4812 ( .B1(n4169), .B2(n4168), .A(n4167), .ZN(n4170) );
  OAI21_X1 U4813 ( .B1(n4171), .B2(n4186), .A(n4170), .ZN(n4234) );
  MUX2_X1 U4814 ( .A(REG1_REG_22__SCAN_IN), .B(n4234), .S(n4624), .Z(U3540) );
  INV_X1 U4815 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4174) );
  AOI21_X1 U4816 ( .B1(n4173), .B2(n4594), .A(n4172), .ZN(n4235) );
  MUX2_X1 U4817 ( .A(n4174), .B(n4235), .S(n4624), .Z(n4175) );
  OAI21_X1 U4818 ( .B1(n4201), .B2(n4238), .A(n4175), .ZN(U3539) );
  AOI21_X1 U4819 ( .B1(n4177), .B2(n4594), .A(n4176), .ZN(n4239) );
  MUX2_X1 U4820 ( .A(n4178), .B(n4239), .S(n4624), .Z(n4179) );
  OAI21_X1 U4821 ( .B1(n4201), .B2(n4242), .A(n4179), .ZN(U3538) );
  INV_X1 U4822 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4182) );
  AOI21_X1 U4823 ( .B1(n4181), .B2(n4594), .A(n4180), .ZN(n4243) );
  MUX2_X1 U4824 ( .A(n4182), .B(n4243), .S(n4624), .Z(n4183) );
  OAI21_X1 U4825 ( .B1(n4201), .B2(n4246), .A(n4183), .ZN(U3537) );
  OAI211_X1 U4826 ( .C1(n4187), .C2(n4186), .A(n4185), .B(n4184), .ZN(n4247)
         );
  MUX2_X1 U4827 ( .A(REG1_REG_18__SCAN_IN), .B(n4247), .S(n4624), .Z(U3536) );
  NAND2_X1 U4828 ( .A1(n4188), .A2(n4594), .ZN(n4190) );
  AND2_X1 U4829 ( .A1(n4190), .A2(n4189), .ZN(n4248) );
  MUX2_X1 U4830 ( .A(n4191), .B(n4248), .S(n4624), .Z(n4192) );
  OAI21_X1 U4831 ( .B1(n4201), .B2(n4251), .A(n4192), .ZN(U3535) );
  INV_X1 U4832 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4195) );
  AOI21_X1 U4833 ( .B1(n4194), .B2(n4594), .A(n4193), .ZN(n4252) );
  MUX2_X1 U4834 ( .A(n4195), .B(n4252), .S(n4624), .Z(n4196) );
  OAI21_X1 U4835 ( .B1(n4201), .B2(n4255), .A(n4196), .ZN(U3534) );
  AOI21_X1 U4836 ( .B1(n4594), .B2(n4198), .A(n4197), .ZN(n4256) );
  MUX2_X1 U4837 ( .A(n4199), .B(n4256), .S(n4624), .Z(n4200) );
  OAI21_X1 U4838 ( .B1(n4201), .B2(n4260), .A(n4200), .ZN(U3533) );
  NAND3_X1 U4839 ( .A1(n4203), .A2(n4602), .A3(n4202), .ZN(n4204) );
  OAI211_X1 U4840 ( .C1(n4206), .C2(n4596), .A(n4205), .B(n4204), .ZN(n4261)
         );
  MUX2_X1 U4841 ( .A(REG1_REG_14__SCAN_IN), .B(n4261), .S(n4624), .Z(U3532) );
  NAND2_X1 U4842 ( .A1(n4207), .A2(n4594), .ZN(n4208) );
  OAI211_X1 U4843 ( .C1(n4591), .C2(n4210), .A(n4209), .B(n4208), .ZN(n4262)
         );
  MUX2_X1 U4844 ( .A(REG1_REG_13__SCAN_IN), .B(n4262), .S(n4624), .Z(U3531) );
  INV_X1 U4845 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4211) );
  MUX2_X1 U4846 ( .A(n4211), .B(n4302), .S(n4605), .Z(n4212) );
  OAI21_X1 U4847 ( .B1(n4213), .B2(n4259), .A(n4212), .ZN(U3516) );
  OAI21_X1 U4848 ( .B1(n4218), .B2(n4259), .A(n4217), .ZN(U3514) );
  MUX2_X1 U4849 ( .A(REG0_REG_27__SCAN_IN), .B(n4219), .S(n4605), .Z(U3513) );
  MUX2_X1 U4850 ( .A(REG0_REG_26__SCAN_IN), .B(n4220), .S(n4605), .Z(U3512) );
  INV_X1 U4851 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4222) );
  MUX2_X1 U4852 ( .A(n4222), .B(n4221), .S(n4605), .Z(n4223) );
  OAI21_X1 U4853 ( .B1(n4224), .B2(n4259), .A(n4223), .ZN(U3511) );
  INV_X1 U4854 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4226) );
  MUX2_X1 U4855 ( .A(n4226), .B(n4225), .S(n4605), .Z(n4227) );
  OAI21_X1 U4856 ( .B1(n4228), .B2(n4259), .A(n4227), .ZN(U3510) );
  INV_X1 U4857 ( .A(n4259), .ZN(n4231) );
  MUX2_X1 U4858 ( .A(REG0_REG_23__SCAN_IN), .B(n4229), .S(n4605), .Z(n4230) );
  AOI21_X1 U4859 ( .B1(n4232), .B2(n4231), .A(n4230), .ZN(n4233) );
  INV_X1 U4860 ( .A(n4233), .ZN(U3509) );
  MUX2_X1 U4861 ( .A(REG0_REG_22__SCAN_IN), .B(n4234), .S(n4605), .Z(U3508) );
  INV_X1 U4862 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4236) );
  MUX2_X1 U4863 ( .A(n4236), .B(n4235), .S(n4605), .Z(n4237) );
  OAI21_X1 U4864 ( .B1(n4238), .B2(n4259), .A(n4237), .ZN(U3507) );
  INV_X1 U4865 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4240) );
  MUX2_X1 U4866 ( .A(n4240), .B(n4239), .S(n4605), .Z(n4241) );
  OAI21_X1 U4867 ( .B1(n4242), .B2(n4259), .A(n4241), .ZN(U3506) );
  MUX2_X1 U4868 ( .A(n4244), .B(n4243), .S(n4605), .Z(n4245) );
  OAI21_X1 U4869 ( .B1(n4246), .B2(n4259), .A(n4245), .ZN(U3505) );
  MUX2_X1 U4870 ( .A(REG0_REG_18__SCAN_IN), .B(n4247), .S(n4605), .Z(U3503) );
  INV_X1 U4871 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4249) );
  MUX2_X1 U4872 ( .A(n4249), .B(n4248), .S(n4605), .Z(n4250) );
  OAI21_X1 U4873 ( .B1(n4251), .B2(n4259), .A(n4250), .ZN(U3501) );
  INV_X1 U4874 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4253) );
  MUX2_X1 U4875 ( .A(n4253), .B(n4252), .S(n4605), .Z(n4254) );
  OAI21_X1 U4876 ( .B1(n4255), .B2(n4259), .A(n4254), .ZN(U3499) );
  INV_X1 U4877 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4257) );
  MUX2_X1 U4878 ( .A(n4257), .B(n4256), .S(n4605), .Z(n4258) );
  OAI21_X1 U4879 ( .B1(n4260), .B2(n4259), .A(n4258), .ZN(U3497) );
  MUX2_X1 U4880 ( .A(REG0_REG_14__SCAN_IN), .B(n4261), .S(n4605), .Z(U3495) );
  MUX2_X1 U4881 ( .A(REG0_REG_13__SCAN_IN), .B(n4262), .S(n4605), .Z(U3493) );
  MUX2_X1 U4882 ( .A(DATAI_30_), .B(n4263), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U4883 ( .A(DATAI_28_), .B(n4264), .S(STATE_REG_SCAN_IN), .Z(U3324)
         );
  MUX2_X1 U4884 ( .A(n4265), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U4885 ( .A(n4266), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U4886 ( .A(DATAI_25_), .B(n4267), .S(STATE_REG_SCAN_IN), .Z(U3327)
         );
  MUX2_X1 U4887 ( .A(n4268), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U4888 ( .A(n4269), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U4889 ( .A(DATAI_21_), .B(n4270), .S(STATE_REG_SCAN_IN), .Z(U3331)
         );
  MUX2_X1 U4890 ( .A(DATAI_20_), .B(n4271), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4891 ( .A(n4272), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U4892 ( .A(n4273), .B(DATAI_14_), .S(U3149), .Z(U3338) );
  MUX2_X1 U4893 ( .A(DATAI_4_), .B(n4274), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4894 ( .A(n4275), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U4895 ( .A(n4276), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4896 ( .A(n4277), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  MUX2_X1 U4897 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(STATE_REG_SCAN_IN), 
        .Z(U3352) );
  NOR2_X1 U4898 ( .A1(STATE_REG_SCAN_IN), .A2(n4278), .ZN(n4404) );
  OAI22_X1 U4899 ( .A1(n4282), .A2(n4281), .B1(n4280), .B2(n4279), .ZN(n4283)
         );
  AOI211_X1 U4900 ( .C1(n4285), .C2(n4284), .A(n4404), .B(n4283), .ZN(n4293)
         );
  OAI21_X1 U4901 ( .B1(n4288), .B2(n4291), .A(n4287), .ZN(n4289) );
  OAI211_X1 U4902 ( .C1(n2151), .C2(n4291), .A(n4290), .B(n4289), .ZN(n4292)
         );
  OAI211_X1 U4903 ( .C1(n4295), .C2(n4294), .A(n4293), .B(n4292), .ZN(U3238)
         );
  AOI22_X1 U4904 ( .A1(n4297), .A2(n4498), .B1(n4296), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n4298) );
  OAI21_X1 U4905 ( .B1(n4296), .B2(n4299), .A(n4298), .ZN(U3260) );
  AOI22_X1 U4906 ( .A1(n4300), .A2(n4498), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4296), .ZN(n4301) );
  OAI21_X1 U4907 ( .B1(n4296), .B2(n4302), .A(n4301), .ZN(U3261) );
  AOI211_X1 U4908 ( .C1(n4305), .C2(n4304), .A(n4303), .B(n4313), .ZN(n4307)
         );
  AOI211_X1 U4909 ( .C1(n4436), .C2(ADDR_REG_5__SCAN_IN), .A(n4307), .B(n4306), 
        .ZN(n4312) );
  OAI211_X1 U4910 ( .C1(n4310), .C2(n4309), .A(n4388), .B(n4308), .ZN(n4311)
         );
  OAI211_X1 U4911 ( .C1(n4443), .C2(n4552), .A(n4312), .B(n4311), .ZN(U3245)
         );
  AOI211_X1 U4912 ( .C1(n4316), .C2(n4315), .A(n4314), .B(n4313), .ZN(n4317)
         );
  AOI211_X1 U4913 ( .C1(n4436), .C2(ADDR_REG_6__SCAN_IN), .A(n4318), .B(n4317), 
        .ZN(n4322) );
  OAI211_X1 U4914 ( .C1(REG2_REG_6__SCAN_IN), .C2(n4320), .A(n4388), .B(n4319), 
        .ZN(n4321) );
  OAI211_X1 U4915 ( .C1(n4443), .C2(n2167), .A(n4322), .B(n4321), .ZN(U3246)
         );
  AOI22_X1 U4916 ( .A1(n4323), .A2(n4617), .B1(REG1_REG_7__SCAN_IN), .B2(n4549), .ZN(n4325) );
  OAI21_X1 U4917 ( .B1(n4326), .B2(n4325), .A(n4438), .ZN(n4324) );
  AOI21_X1 U4918 ( .B1(n4326), .B2(n4325), .A(n4324), .ZN(n4328) );
  AOI211_X1 U4919 ( .C1(n4436), .C2(ADDR_REG_7__SCAN_IN), .A(n4328), .B(n4327), 
        .ZN(n4333) );
  OAI211_X1 U4920 ( .C1(n4331), .C2(n4330), .A(n4388), .B(n4329), .ZN(n4332)
         );
  OAI211_X1 U4921 ( .C1(n4443), .C2(n4549), .A(n4333), .B(n4332), .ZN(U3247)
         );
  OAI211_X1 U4922 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4335), .A(n4388), .B(n4334), 
        .ZN(n4337) );
  NAND2_X1 U4923 ( .A1(n4337), .A2(n4336), .ZN(n4338) );
  AOI21_X1 U4924 ( .B1(n4436), .B2(ADDR_REG_8__SCAN_IN), .A(n4338), .ZN(n4342)
         );
  OAI211_X1 U4925 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4340), .A(n4438), .B(n4339), 
        .ZN(n4341) );
  OAI211_X1 U4926 ( .C1(n4443), .C2(n4343), .A(n4342), .B(n4341), .ZN(U3248)
         );
  OAI211_X1 U4927 ( .C1(n4346), .C2(n4345), .A(n4438), .B(n4344), .ZN(n4351)
         );
  OAI211_X1 U4928 ( .C1(n4349), .C2(n4348), .A(n4388), .B(n4347), .ZN(n4350)
         );
  OAI211_X1 U4929 ( .C1(n4443), .C2(n4352), .A(n4351), .B(n4350), .ZN(n4353)
         );
  AOI211_X1 U4930 ( .C1(n4436), .C2(ADDR_REG_9__SCAN_IN), .A(n4354), .B(n4353), 
        .ZN(n4355) );
  INV_X1 U4931 ( .A(n4355), .ZN(U3249) );
  OAI211_X1 U4932 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4357), .A(n4438), .B(n4356), .ZN(n4361) );
  OAI211_X1 U4933 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4359), .A(n4388), .B(n4358), .ZN(n4360) );
  OAI211_X1 U4934 ( .C1(n4443), .C2(n4362), .A(n4361), .B(n4360), .ZN(n4363)
         );
  AOI211_X1 U4935 ( .C1(n4436), .C2(ADDR_REG_10__SCAN_IN), .A(n4364), .B(n4363), .ZN(n4365) );
  INV_X1 U4936 ( .A(n4365), .ZN(U3250) );
  OAI211_X1 U4937 ( .C1(n4368), .C2(n4367), .A(n4388), .B(n4366), .ZN(n4370)
         );
  NAND2_X1 U4938 ( .A1(n4370), .A2(n4369), .ZN(n4371) );
  AOI21_X1 U4939 ( .B1(n4436), .B2(ADDR_REG_11__SCAN_IN), .A(n4371), .ZN(n4376) );
  OAI211_X1 U4940 ( .C1(n4374), .C2(n4373), .A(n4438), .B(n4372), .ZN(n4375)
         );
  OAI211_X1 U4941 ( .C1(n4443), .C2(n4377), .A(n4376), .B(n4375), .ZN(U3251)
         );
  OAI211_X1 U4942 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4379), .A(n4388), .B(n4378), .ZN(n4380) );
  NAND2_X1 U4943 ( .A1(n4381), .A2(n4380), .ZN(n4382) );
  AOI21_X1 U4944 ( .B1(n4436), .B2(ADDR_REG_12__SCAN_IN), .A(n4382), .ZN(n4386) );
  OAI211_X1 U4945 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4384), .A(n4438), .B(n4383), .ZN(n4385) );
  OAI211_X1 U4946 ( .C1(n4443), .C2(n2166), .A(n4386), .B(n4385), .ZN(U3252)
         );
  AOI21_X1 U4947 ( .B1(n4399), .B2(n2482), .A(n4387), .ZN(n4391) );
  OAI21_X1 U4948 ( .B1(n4391), .B2(n4390), .A(n4388), .ZN(n4389) );
  AOI21_X1 U4949 ( .B1(n4391), .B2(n4390), .A(n4389), .ZN(n4393) );
  AOI211_X1 U4950 ( .C1(n4436), .C2(ADDR_REG_13__SCAN_IN), .A(n4393), .B(n4392), .ZN(n4398) );
  OAI211_X1 U4951 ( .C1(n4396), .C2(n4395), .A(n4438), .B(n4394), .ZN(n4397)
         );
  OAI211_X1 U4952 ( .C1(n4443), .C2(n4399), .A(n4398), .B(n4397), .ZN(U3253)
         );
  AOI211_X1 U4953 ( .C1(n4402), .C2(n4401), .A(n4400), .B(n4430), .ZN(n4403)
         );
  AOI211_X1 U4954 ( .C1(n4436), .C2(ADDR_REG_15__SCAN_IN), .A(n4404), .B(n4403), .ZN(n4409) );
  OAI211_X1 U4955 ( .C1(n4407), .C2(n4406), .A(n4438), .B(n4405), .ZN(n4408)
         );
  OAI211_X1 U4956 ( .C1(n4443), .C2(n4536), .A(n4409), .B(n4408), .ZN(U3255)
         );
  INV_X1 U4957 ( .A(n4410), .ZN(n4414) );
  AOI221_X1 U4958 ( .B1(n4412), .B2(n4411), .C1(n2260), .C2(n4411), .A(n4430), 
        .ZN(n4413) );
  AOI211_X1 U4959 ( .C1(n4436), .C2(ADDR_REG_16__SCAN_IN), .A(n4414), .B(n4413), .ZN(n4418) );
  OAI221_X1 U4960 ( .B1(n4416), .B2(REG1_REG_16__SCAN_IN), .C1(n4416), .C2(
        n4415), .A(n4438), .ZN(n4417) );
  OAI211_X1 U4961 ( .C1(n4443), .C2(n4534), .A(n4418), .B(n4417), .ZN(U3256)
         );
  AOI221_X1 U4962 ( .B1(n4421), .B2(n4420), .C1(n4419), .C2(n4420), .A(n4430), 
        .ZN(n4422) );
  AOI211_X1 U4963 ( .C1(ADDR_REG_17__SCAN_IN), .C2(n4436), .A(n4423), .B(n4422), .ZN(n4428) );
  OAI221_X1 U4964 ( .B1(n4426), .B2(n4425), .C1(n4426), .C2(n4424), .A(n4438), 
        .ZN(n4427) );
  OAI211_X1 U4965 ( .C1(n4443), .C2(n4429), .A(n4428), .B(n4427), .ZN(U3257)
         );
  AOI211_X1 U4966 ( .C1(n4433), .C2(n4432), .A(n4431), .B(n4430), .ZN(n4434)
         );
  AOI211_X1 U4967 ( .C1(n4436), .C2(ADDR_REG_18__SCAN_IN), .A(n4435), .B(n4434), .ZN(n4442) );
  OAI211_X1 U4968 ( .C1(n4440), .C2(n4439), .A(n4438), .B(n4437), .ZN(n4441)
         );
  OAI211_X1 U4969 ( .C1(n4443), .C2(n4530), .A(n4442), .B(n4441), .ZN(U3258)
         );
  XNOR2_X1 U4970 ( .A(n4444), .B(n4450), .ZN(n4454) );
  AOI22_X1 U4971 ( .A1(n4445), .A2(n4479), .B1(n4457), .B2(n4478), .ZN(n4446)
         );
  OAI21_X1 U4972 ( .B1(n4447), .B2(n4482), .A(n4446), .ZN(n4453) );
  NAND2_X1 U4973 ( .A1(n4449), .A2(n4448), .ZN(n4451) );
  XNOR2_X1 U4974 ( .A(n4451), .B(n4450), .ZN(n4597) );
  NOR2_X1 U4975 ( .A1(n4597), .A2(n4487), .ZN(n4452) );
  AOI211_X1 U4976 ( .C1(n4454), .C2(n4502), .A(n4453), .B(n4452), .ZN(n4598)
         );
  AOI22_X1 U4977 ( .A1(n4455), .A2(n4491), .B1(REG2_REG_11__SCAN_IN), .B2(
        n4296), .ZN(n4460) );
  INV_X1 U4978 ( .A(n4597), .ZN(n4458) );
  AOI21_X1 U4979 ( .B1(n4457), .B2(n4456), .A(n2081), .ZN(n4601) );
  AOI22_X1 U4980 ( .A1(n4458), .A2(n4501), .B1(n4498), .B2(n4601), .ZN(n4459)
         );
  OAI211_X1 U4981 ( .C1(n4296), .C2(n4598), .A(n4460), .B(n4459), .ZN(U3279)
         );
  AOI22_X1 U4982 ( .A1(n4461), .A2(n4491), .B1(REG2_REG_10__SCAN_IN), .B2(
        n4296), .ZN(n4466) );
  INV_X1 U4983 ( .A(n4462), .ZN(n4463) );
  AOI22_X1 U4984 ( .A1(n4464), .A2(n4501), .B1(n4498), .B2(n4463), .ZN(n4465)
         );
  OAI211_X1 U4985 ( .C1(n4296), .C2(n4467), .A(n4466), .B(n4465), .ZN(U3280)
         );
  AOI22_X1 U4986 ( .A1(n4468), .A2(n4491), .B1(REG2_REG_8__SCAN_IN), .B2(n4296), .ZN(n4473) );
  INV_X1 U4987 ( .A(n4469), .ZN(n4470) );
  AOI22_X1 U4988 ( .A1(n4471), .A2(n4501), .B1(n4498), .B2(n4470), .ZN(n4472)
         );
  OAI211_X1 U4989 ( .C1(n4296), .C2(n4474), .A(n4473), .B(n4472), .ZN(U3282)
         );
  INV_X1 U4990 ( .A(n4486), .ZN(n4477) );
  OAI21_X1 U4991 ( .B1(n4477), .B2(n4476), .A(n4475), .ZN(n4490) );
  AOI22_X1 U4992 ( .A1(n4480), .A2(n4479), .B1(n4478), .B2(n4492), .ZN(n4481)
         );
  OAI21_X1 U4993 ( .B1(n4483), .B2(n4482), .A(n4481), .ZN(n4489) );
  OAI21_X1 U4994 ( .B1(n4486), .B2(n4485), .A(n4484), .ZN(n4559) );
  NOR2_X1 U4995 ( .A1(n4559), .A2(n4487), .ZN(n4488) );
  AOI211_X1 U4996 ( .C1(n4502), .C2(n4490), .A(n4489), .B(n4488), .ZN(n4557)
         );
  AOI22_X1 U4997 ( .A1(REG3_REG_1__SCAN_IN), .A2(n4491), .B1(
        REG2_REG_1__SCAN_IN), .B2(n4296), .ZN(n4500) );
  NAND2_X1 U4998 ( .A1(n4493), .A2(n4492), .ZN(n4494) );
  NAND2_X1 U4999 ( .A1(n4495), .A2(n4494), .ZN(n4558) );
  INV_X1 U5000 ( .A(n4558), .ZN(n4497) );
  INV_X1 U5001 ( .A(n4559), .ZN(n4496) );
  AOI22_X1 U5002 ( .A1(n4498), .A2(n4497), .B1(n4496), .B2(n4501), .ZN(n4499)
         );
  OAI211_X1 U5003 ( .C1(n4296), .C2(n4557), .A(n4500), .B(n4499), .ZN(U3289)
         );
  AOI22_X1 U5004 ( .A1(n4501), .A2(n4555), .B1(REG2_REG_0__SCAN_IN), .B2(n4296), .ZN(n4514) );
  OAI21_X1 U5005 ( .B1(n4503), .B2(n4502), .A(n4555), .ZN(n4504) );
  OAI21_X1 U5006 ( .B1(n4506), .B2(n4505), .A(n4504), .ZN(n4553) );
  NOR2_X1 U5007 ( .A1(n4508), .A2(n4507), .ZN(n4554) );
  INV_X1 U5008 ( .A(n4554), .ZN(n4510) );
  NOR2_X1 U5009 ( .A1(n4510), .A2(n4509), .ZN(n4512) );
  OAI21_X1 U5010 ( .B1(n4553), .B2(n4512), .A(n4511), .ZN(n4513) );
  OAI211_X1 U5011 ( .C1(n4515), .C2(n2306), .A(n4514), .B(n4513), .ZN(U3290)
         );
  AND2_X1 U5012 ( .A1(D_REG_31__SCAN_IN), .A2(n4526), .ZN(U3291) );
  AND2_X1 U5013 ( .A1(D_REG_30__SCAN_IN), .A2(n4526), .ZN(U3292) );
  AND2_X1 U5014 ( .A1(D_REG_29__SCAN_IN), .A2(n4526), .ZN(U3293) );
  NOR2_X1 U5015 ( .A1(n4525), .A2(n4516), .ZN(U3294) );
  AND2_X1 U5016 ( .A1(D_REG_27__SCAN_IN), .A2(n4526), .ZN(U3295) );
  AND2_X1 U5017 ( .A1(D_REG_26__SCAN_IN), .A2(n4526), .ZN(U3296) );
  AND2_X1 U5018 ( .A1(D_REG_25__SCAN_IN), .A2(n4526), .ZN(U3297) );
  AND2_X1 U5019 ( .A1(D_REG_24__SCAN_IN), .A2(n4526), .ZN(U3298) );
  AND2_X1 U5020 ( .A1(D_REG_23__SCAN_IN), .A2(n4526), .ZN(U3299) );
  AND2_X1 U5021 ( .A1(D_REG_22__SCAN_IN), .A2(n4526), .ZN(U3300) );
  NOR2_X1 U5022 ( .A1(n4525), .A2(n4517), .ZN(U3301) );
  AND2_X1 U5023 ( .A1(D_REG_20__SCAN_IN), .A2(n4526), .ZN(U3302) );
  NOR2_X1 U5024 ( .A1(n4525), .A2(n4518), .ZN(U3303) );
  NOR2_X1 U5025 ( .A1(n4525), .A2(n4519), .ZN(U3304) );
  AND2_X1 U5026 ( .A1(D_REG_17__SCAN_IN), .A2(n4526), .ZN(U3305) );
  NOR2_X1 U5027 ( .A1(n4525), .A2(n4520), .ZN(U3306) );
  AND2_X1 U5028 ( .A1(D_REG_15__SCAN_IN), .A2(n4526), .ZN(U3307) );
  AND2_X1 U5029 ( .A1(D_REG_14__SCAN_IN), .A2(n4526), .ZN(U3308) );
  NOR2_X1 U5030 ( .A1(n4525), .A2(n4521), .ZN(U3309) );
  NOR2_X1 U5031 ( .A1(n4525), .A2(n4522), .ZN(U3310) );
  NOR2_X1 U5032 ( .A1(n4525), .A2(n4523), .ZN(U3311) );
  AND2_X1 U5033 ( .A1(D_REG_10__SCAN_IN), .A2(n4526), .ZN(U3312) );
  NOR2_X1 U5034 ( .A1(n4525), .A2(n4524), .ZN(U3313) );
  AND2_X1 U5035 ( .A1(D_REG_8__SCAN_IN), .A2(n4526), .ZN(U3314) );
  AND2_X1 U5036 ( .A1(D_REG_7__SCAN_IN), .A2(n4526), .ZN(U3315) );
  AND2_X1 U5037 ( .A1(D_REG_6__SCAN_IN), .A2(n4526), .ZN(U3316) );
  AND2_X1 U5038 ( .A1(D_REG_5__SCAN_IN), .A2(n4526), .ZN(U3317) );
  AND2_X1 U5039 ( .A1(D_REG_4__SCAN_IN), .A2(n4526), .ZN(U3318) );
  AND2_X1 U5040 ( .A1(D_REG_3__SCAN_IN), .A2(n4526), .ZN(U3319) );
  AND2_X1 U5041 ( .A1(D_REG_2__SCAN_IN), .A2(n4526), .ZN(U3320) );
  OAI21_X1 U5042 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4527), .ZN(
        n4528) );
  INV_X1 U5043 ( .A(n4528), .ZN(U3329) );
  INV_X1 U5044 ( .A(DATAI_18_), .ZN(n4529) );
  AOI22_X1 U5045 ( .A1(STATE_REG_SCAN_IN), .A2(n4530), .B1(n4529), .B2(U3149), 
        .ZN(U3334) );
  OAI22_X1 U5046 ( .A1(U3149), .A2(n4531), .B1(DATAI_17_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4532) );
  INV_X1 U5047 ( .A(n4532), .ZN(U3335) );
  INV_X1 U5048 ( .A(DATAI_16_), .ZN(n4533) );
  AOI22_X1 U5049 ( .A1(STATE_REG_SCAN_IN), .A2(n4534), .B1(n4533), .B2(U3149), 
        .ZN(U3336) );
  AOI22_X1 U5050 ( .A1(STATE_REG_SCAN_IN), .A2(n4536), .B1(n4535), .B2(U3149), 
        .ZN(U3337) );
  OAI22_X1 U5051 ( .A1(U3149), .A2(n4537), .B1(DATAI_13_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4538) );
  INV_X1 U5052 ( .A(n4538), .ZN(U3339) );
  INV_X1 U5053 ( .A(DATAI_12_), .ZN(n4539) );
  AOI22_X1 U5054 ( .A1(STATE_REG_SCAN_IN), .A2(n2166), .B1(n4539), .B2(U3149), 
        .ZN(U3340) );
  OAI22_X1 U5055 ( .A1(U3149), .A2(n4540), .B1(DATAI_11_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4541) );
  INV_X1 U5056 ( .A(n4541), .ZN(U3341) );
  OAI22_X1 U5057 ( .A1(U3149), .A2(n4542), .B1(DATAI_10_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4543) );
  INV_X1 U5058 ( .A(n4543), .ZN(U3342) );
  OAI22_X1 U5059 ( .A1(U3149), .A2(n4544), .B1(DATAI_9_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4545) );
  INV_X1 U5060 ( .A(n4545), .ZN(U3343) );
  OAI22_X1 U5061 ( .A1(U3149), .A2(n4546), .B1(DATAI_8_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4547) );
  INV_X1 U5062 ( .A(n4547), .ZN(U3344) );
  INV_X1 U5063 ( .A(DATAI_7_), .ZN(n4548) );
  AOI22_X1 U5064 ( .A1(STATE_REG_SCAN_IN), .A2(n4549), .B1(n4548), .B2(U3149), 
        .ZN(U3345) );
  INV_X1 U5065 ( .A(DATAI_6_), .ZN(n4550) );
  AOI22_X1 U5066 ( .A1(STATE_REG_SCAN_IN), .A2(n2167), .B1(n4550), .B2(U3149), 
        .ZN(U3346) );
  AOI22_X1 U5067 ( .A1(STATE_REG_SCAN_IN), .A2(n4552), .B1(n4551), .B2(U3149), 
        .ZN(U3347) );
  AOI211_X1 U5068 ( .C1(n4577), .C2(n4555), .A(n4554), .B(n4553), .ZN(n4606)
         );
  INV_X1 U5069 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4556) );
  AOI22_X1 U5070 ( .A1(n4605), .A2(n4606), .B1(n4556), .B2(n4603), .ZN(U3467)
         );
  INV_X1 U5071 ( .A(n4557), .ZN(n4561) );
  OAI22_X1 U5072 ( .A1(n4559), .A2(n4596), .B1(n4591), .B2(n4558), .ZN(n4560)
         );
  NOR2_X1 U5073 ( .A1(n4561), .A2(n4560), .ZN(n4608) );
  INV_X1 U5074 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4562) );
  AOI22_X1 U5075 ( .A1(n4605), .A2(n4608), .B1(n4562), .B2(n4603), .ZN(U3469)
         );
  AND3_X1 U5076 ( .A1(n4564), .A2(n4602), .A3(n4563), .ZN(n4566) );
  AOI211_X1 U5077 ( .C1(n4577), .C2(n4567), .A(n4566), .B(n4565), .ZN(n4610)
         );
  INV_X1 U5078 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4568) );
  AOI22_X1 U5079 ( .A1(n4605), .A2(n4610), .B1(n4568), .B2(n4603), .ZN(U3471)
         );
  AOI22_X1 U5080 ( .A1(n4570), .A2(n4577), .B1(n4602), .B2(n4569), .ZN(n4571)
         );
  AND2_X1 U5081 ( .A1(n4572), .A2(n4571), .ZN(n4612) );
  INV_X1 U5082 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4573) );
  AOI22_X1 U5083 ( .A1(n4605), .A2(n4612), .B1(n4573), .B2(n4603), .ZN(U3473)
         );
  INV_X1 U5084 ( .A(n4574), .ZN(n4576) );
  AOI211_X1 U5085 ( .C1(n4578), .C2(n4577), .A(n4576), .B(n4575), .ZN(n4614)
         );
  INV_X1 U5086 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4579) );
  AOI22_X1 U5087 ( .A1(n4605), .A2(n4614), .B1(n4579), .B2(n4603), .ZN(U3475)
         );
  OAI21_X1 U5088 ( .B1(n4591), .B2(n4581), .A(n4580), .ZN(n4582) );
  AOI21_X1 U5089 ( .B1(n4583), .B2(n4594), .A(n4582), .ZN(n4616) );
  INV_X1 U5090 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4584) );
  AOI22_X1 U5091 ( .A1(n4605), .A2(n4616), .B1(n4584), .B2(n4603), .ZN(U3477)
         );
  AOI211_X1 U5092 ( .C1(n4587), .C2(n4594), .A(n4586), .B(n4585), .ZN(n4618)
         );
  INV_X1 U5093 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4588) );
  AOI22_X1 U5094 ( .A1(n4605), .A2(n4618), .B1(n4588), .B2(n4603), .ZN(U3481)
         );
  OAI21_X1 U5095 ( .B1(n4591), .B2(n4590), .A(n4589), .ZN(n4592) );
  AOI21_X1 U5096 ( .B1(n4594), .B2(n4593), .A(n4592), .ZN(n4620) );
  AOI22_X1 U5097 ( .A1(n4605), .A2(n4620), .B1(n4595), .B2(n4603), .ZN(U3485)
         );
  NOR2_X1 U5098 ( .A1(n4597), .A2(n4596), .ZN(n4600) );
  INV_X1 U5099 ( .A(n4598), .ZN(n4599) );
  AOI211_X1 U5100 ( .C1(n4602), .C2(n4601), .A(n4600), .B(n4599), .ZN(n4623)
         );
  INV_X1 U5101 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4604) );
  AOI22_X1 U5102 ( .A1(n4605), .A2(n4623), .B1(n4604), .B2(n4603), .ZN(U3489)
         );
  AOI22_X1 U5103 ( .A1(n4624), .A2(n4606), .B1(n2314), .B2(n4621), .ZN(U3518)
         );
  AOI22_X1 U5104 ( .A1(n4624), .A2(n4608), .B1(n4607), .B2(n4621), .ZN(U3519)
         );
  AOI22_X1 U5105 ( .A1(n4624), .A2(n4610), .B1(n4609), .B2(n4621), .ZN(U3520)
         );
  AOI22_X1 U5106 ( .A1(n4624), .A2(n4612), .B1(n4611), .B2(n4621), .ZN(U3521)
         );
  AOI22_X1 U5107 ( .A1(n4624), .A2(n4614), .B1(n4613), .B2(n4621), .ZN(U3522)
         );
  AOI22_X1 U5108 ( .A1(n4624), .A2(n4616), .B1(n4615), .B2(n4621), .ZN(U3523)
         );
  AOI22_X1 U5109 ( .A1(n4624), .A2(n4618), .B1(n4617), .B2(n4621), .ZN(U3525)
         );
  AOI22_X1 U5110 ( .A1(n4624), .A2(n4620), .B1(n4619), .B2(n4621), .ZN(U3527)
         );
  AOI22_X1 U5111 ( .A1(n4624), .A2(n4623), .B1(n4622), .B2(n4621), .ZN(U3529)
         );
  CLKBUF_X1 U2283 ( .A(n2356), .Z(n2832) );
endmodule

