

module b21_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898;

  NAND2_X1 U5108 ( .A1(n5256), .A2(n5088), .ZN(n8242) );
  CLKBUF_X2 U5109 ( .A(n6552), .Z(n9423) );
  CLKBUF_X1 U5110 ( .A(n6576), .Z(n6931) );
  INV_X1 U5111 ( .A(n8242), .ZN(n5255) );
  INV_X1 U5112 ( .A(n9287), .ZN(n9198) );
  INV_X1 U5113 ( .A(n6231), .ZN(n9427) );
  INV_X1 U5114 ( .A(n8531), .ZN(n6757) );
  AND3_X1 U5115 ( .A1(n7094), .A2(n7093), .A3(n7092), .ZN(n10677) );
  INV_X1 U5116 ( .A(n9287), .ZN(n9235) );
  INV_X1 U5117 ( .A(n6813), .ZN(n10662) );
  NAND2_X1 U5118 ( .A1(n8877), .A2(n8878), .ZN(n8876) );
  INV_X1 U5119 ( .A(n8047), .ZN(n8263) );
  OR2_X1 U5120 ( .A1(n5698), .A2(n9146), .ZN(n5706) );
  NAND2_X1 U5121 ( .A1(n7182), .A2(n7181), .ZN(n7393) );
  NAND2_X1 U5122 ( .A1(n5635), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5634) );
  XNOR2_X1 U5123 ( .A(n5645), .B(P1_IR_REG_22__SCAN_IN), .ZN(n9661) );
  AND2_X1 U5124 ( .A1(n5312), .A2(n5048), .ZN(n5044) );
  OAI21_X2 U5125 ( .B1(n9303), .B2(n9301), .A(n9299), .ZN(n9362) );
  AOI22_X2 U5126 ( .A1(n8894), .A2(n8902), .B1(n8901), .B2(n8772), .ZN(n8877)
         );
  INV_X4 U5127 ( .A(n5712), .ZN(n5713) );
  NAND2_X2 U5128 ( .A1(n5456), .A2(n5455), .ZN(n5712) );
  XNOR2_X2 U5129 ( .A(n8704), .B(n7142), .ZN(n8047) );
  XNOR2_X2 U5130 ( .A(n5634), .B(n5651), .ZN(n5750) );
  OAI22_X2 U5131 ( .A1(n9002), .A2(n8763), .B1(n8762), .B2(n9123), .ZN(n8989)
         );
  XNOR2_X2 U5132 ( .A(n5697), .B(P2_IR_REG_1__SCAN_IN), .ZN(n10600) );
  XNOR2_X2 U5133 ( .A(n5706), .B(n5705), .ZN(n6701) );
  AOI211_X1 U5134 ( .C1(n10877), .C2(n9958), .A(n9957), .B(n9956), .ZN(n9959)
         );
  AND2_X1 U5135 ( .A1(n8059), .A2(n8058), .ZN(n9031) );
  NAND2_X1 U5136 ( .A1(n7269), .A2(n7268), .ZN(n7400) );
  NAND2_X1 U5137 ( .A1(n6964), .A2(n8038), .ZN(n8259) );
  INV_X1 U5138 ( .A(n6914), .ZN(n5317) );
  INV_X1 U5139 ( .A(n6860), .ZN(n7003) );
  NAND2_X1 U5140 ( .A1(n6870), .A2(n6732), .ZN(n6871) );
  NAND2_X2 U5141 ( .A1(n8028), .A2(n8027), .ZN(n6732) );
  INV_X1 U5142 ( .A(n6849), .ZN(n5046) );
  AND2_X1 U5143 ( .A1(n6514), .A2(n6756), .ZN(n6698) );
  INV_X2 U5144 ( .A(n10648), .ZN(n9444) );
  INV_X1 U5145 ( .A(n6220), .ZN(n6160) );
  OR2_X1 U5147 ( .A1(n9653), .A2(n9657), .ZN(n6626) );
  NAND2_X1 U5148 ( .A1(n7966), .A2(P1_U3084), .ZN(n10455) );
  OR2_X1 U5149 ( .A1(n5643), .A2(n5884), .ZN(n6018) );
  NAND2_X1 U5150 ( .A1(n5688), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5455) );
  AND3_X2 U5151 ( .A1(n5052), .A2(n5051), .A3(n5050), .ZN(n5746) );
  AND2_X1 U5152 ( .A1(n5395), .A2(n5142), .ZN(n5394) );
  MUX2_X1 U5153 ( .A(n5077), .B(n8281), .S(n8242), .Z(n8245) );
  NAND2_X1 U5154 ( .A1(n5053), .A2(n8780), .ZN(n8800) );
  NAND2_X1 U5155 ( .A1(n5054), .A2(n8778), .ZN(n8815) );
  NAND2_X1 U5156 ( .A1(n9267), .A2(n5589), .ZN(n5588) );
  AOI21_X1 U5157 ( .B1(n9265), .B2(n5586), .A(n5585), .ZN(n5584) );
  NAND2_X1 U5158 ( .A1(n7972), .A2(n7971), .ZN(n8746) );
  NAND2_X1 U5159 ( .A1(n7979), .A2(n7978), .ZN(n8757) );
  NAND2_X1 U5160 ( .A1(n8845), .A2(n8844), .ZN(n8777) );
  XNOR2_X1 U5161 ( .A(n7969), .B(n7968), .ZN(n9419) );
  NAND2_X1 U5162 ( .A1(n8858), .A2(n5147), .ZN(n8845) );
  XNOR2_X1 U5163 ( .A(n7977), .B(n7976), .ZN(n9412) );
  NAND2_X1 U5164 ( .A1(n8876), .A2(n5117), .ZN(n8858) );
  AOI21_X1 U5165 ( .B1(n9377), .B2(n5609), .A(n5603), .ZN(n5602) );
  OAI21_X1 U5166 ( .B1(n7981), .B2(n10229), .A(n7961), .ZN(n7977) );
  NAND2_X1 U5167 ( .A1(n8371), .A2(n8370), .ZN(n9803) );
  NAND2_X1 U5168 ( .A1(n8934), .A2(n8933), .ZN(n8932) );
  NAND2_X1 U5169 ( .A1(n9101), .A2(n5096), .ZN(n8926) );
  NAND2_X1 U5170 ( .A1(n8941), .A2(n8943), .ZN(n9101) );
  AND2_X1 U5171 ( .A1(n5365), .A2(n5364), .ZN(n9794) );
  NAND2_X1 U5172 ( .A1(n8428), .A2(n8427), .ZN(n9951) );
  AOI21_X1 U5173 ( .B1(n8956), .B2(n8768), .A(n5047), .ZN(n8941) );
  NAND2_X1 U5174 ( .A1(n5409), .A2(n5410), .ZN(n8956) );
  NAND2_X1 U5175 ( .A1(n9893), .A2(n9892), .ZN(n9891) );
  NAND2_X1 U5176 ( .A1(n8001), .A2(n8000), .ZN(n9081) );
  NAND2_X1 U5177 ( .A1(n8013), .A2(n8012), .ZN(n9086) );
  NOR2_X1 U5178 ( .A1(n7868), .A2(n8084), .ZN(n8760) );
  NAND2_X1 U5179 ( .A1(n7867), .A2(n5094), .ZN(n7868) );
  NAND2_X1 U5180 ( .A1(n7823), .A2(n5425), .ZN(n7867) );
  NAND2_X1 U5181 ( .A1(n7659), .A2(n7658), .ZN(n7691) );
  NAND2_X1 U5182 ( .A1(n10787), .A2(n5098), .ZN(n7823) );
  NOR2_X1 U5183 ( .A1(n9108), .A2(n8695), .ZN(n5047) );
  NOR2_X2 U5184 ( .A1(n9998), .A2(n5075), .ZN(n9871) );
  OAI21_X1 U5185 ( .B1(n7864), .B2(P2_REG2_REG_14__SCAN_IN), .A(n7552), .ZN(
        n7836) );
  AOI21_X1 U5186 ( .B1(n5572), .B2(n7488), .A(n5569), .ZN(n5568) );
  NAND2_X1 U5187 ( .A1(n5146), .A2(n7415), .ZN(n5055) );
  NAND2_X1 U5188 ( .A1(n7758), .A2(n7757), .ZN(n10876) );
  AND2_X1 U5189 ( .A1(n8286), .A2(n8090), .ZN(n8084) );
  NAND2_X1 U5190 ( .A1(n7208), .A2(n7207), .ZN(n7209) );
  NAND2_X1 U5191 ( .A1(n7809), .A2(n8076), .ZN(n8255) );
  NAND2_X1 U5192 ( .A1(n7519), .A2(n7518), .ZN(n10815) );
  AOI21_X1 U5193 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n7574), .A(n7155), .ZN(
        n7158) );
  NAND2_X1 U5194 ( .A1(n7576), .A2(n7575), .ZN(n7821) );
  NAND2_X1 U5195 ( .A1(n6410), .A2(n6409), .ZN(n6442) );
  NAND2_X1 U5196 ( .A1(n7368), .A2(n7367), .ZN(n9032) );
  AOI21_X1 U5197 ( .B1(n5060), .B2(n9031), .A(n5105), .ZN(n5426) );
  OAI21_X1 U5198 ( .B1(n7535), .B2(P2_REG2_REG_11__SCAN_IN), .A(n7064), .ZN(
        n7066) );
  NAND2_X1 U5199 ( .A1(n6944), .A2(n6943), .ZN(n7141) );
  NAND2_X1 U5200 ( .A1(n6730), .A2(n8259), .ZN(n6944) );
  NAND2_X1 U5201 ( .A1(n6785), .A2(n8030), .ZN(n6730) );
  XNOR2_X1 U5202 ( .A(n5194), .B(n5867), .ZN(n7370) );
  NAND2_X1 U5203 ( .A1(n5819), .A2(n5818), .ZN(n5194) );
  INV_X1 U5204 ( .A(n10677), .ZN(n8049) );
  INV_X2 U5205 ( .A(n10783), .ZN(n10778) );
  INV_X2 U5206 ( .A(n10896), .ZN(n5045) );
  AND3_X2 U5207 ( .A1(n6951), .A2(n6950), .A3(n6949), .ZN(n7142) );
  CLKBUF_X3 U5208 ( .A(n6651), .Z(n9243) );
  INV_X1 U5209 ( .A(n6759), .ZN(n6832) );
  AND3_X1 U5210 ( .A1(n6717), .A2(n6716), .A3(n6715), .ZN(n6795) );
  AND2_X2 U5211 ( .A1(n6755), .A2(n6754), .ZN(n6764) );
  NOR2_X2 U5212 ( .A1(n9289), .A2(n6038), .ZN(n9239) );
  OR2_X2 U5213 ( .A1(n6615), .A2(n10640), .ZN(n8531) );
  OR2_X1 U5214 ( .A1(n6946), .A2(n5702), .ZN(n5057) );
  AND3_X2 U5215 ( .A1(n6079), .A2(n6078), .A3(n6077), .ZN(n10648) );
  INV_X2 U5216 ( .A(n6702), .ZN(n8211) );
  OAI211_X1 U5217 ( .C1(n6149), .C2(n6148), .A(n5559), .B(n5558), .ZN(n6220)
         );
  NAND2_X2 U5218 ( .A1(n6039), .A2(n6626), .ZN(n9289) );
  OR2_X1 U5219 ( .A1(n6729), .A2(n6701), .ZN(n5056) );
  CLKBUF_X3 U5220 ( .A(n6707), .Z(n8169) );
  OAI21_X1 U5221 ( .B1(n5430), .B2(n5432), .A(n5722), .ZN(n5728) );
  INV_X2 U5222 ( .A(n6537), .ZN(n8352) );
  OR2_X1 U5223 ( .A1(n5721), .A2(n5720), .ZN(n5722) );
  INV_X1 U5224 ( .A(n6382), .ZN(n9154) );
  NAND2_X1 U5225 ( .A1(n5648), .A2(n5647), .ZN(n9653) );
  NAND2_X4 U5226 ( .A1(n10503), .A2(n10452), .ZN(n6537) );
  AND2_X1 U5227 ( .A1(n5946), .A2(n9147), .ZN(n6382) );
  AND2_X1 U5228 ( .A1(n5313), .A2(n5044), .ZN(n5809) );
  NAND2_X1 U5229 ( .A1(n5657), .A2(n5656), .ZN(n10503) );
  OR2_X1 U5230 ( .A1(n5941), .A2(n9146), .ZN(n5813) );
  XNOR2_X1 U5231 ( .A(n6020), .B(n6019), .ZN(n9812) );
  MUX2_X1 U5232 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5653), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5654) );
  AND4_X1 U5233 ( .A1(n5453), .A2(SI_0_), .A3(n5451), .A4(n5450), .ZN(n5690)
         );
  NAND2_X2 U5234 ( .A1(n7958), .A2(P1_U3084), .ZN(n10451) );
  AND3_X1 U5235 ( .A1(n5070), .A2(n5667), .A3(n5940), .ZN(n5227) );
  AND2_X1 U5236 ( .A1(n5391), .A2(n5518), .ZN(n5643) );
  AND2_X1 U5237 ( .A1(n5676), .A2(n5360), .ZN(n5671) );
  AND2_X1 U5238 ( .A1(n5059), .A2(n5521), .ZN(n5391) );
  AND3_X1 U5239 ( .A1(n5363), .A2(n5362), .A3(n5361), .ZN(n5676) );
  AND3_X1 U5240 ( .A1(n10196), .A2(n5632), .A3(n6017), .ZN(n5633) );
  INV_X1 U5241 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5048) );
  INV_X1 U5242 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n10204) );
  INV_X1 U5243 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n10390) );
  NOR2_X1 U5244 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5730) );
  NOR2_X1 U5245 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n6057) );
  INV_X1 U5246 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5658) );
  INV_X1 U5247 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6598) );
  NOR2_X1 U5248 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5517) );
  NOR2_X1 U5249 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5050) );
  NOR2_X1 U5250 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5051) );
  NOR2_X1 U5251 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5052) );
  INV_X1 U5252 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n5421) );
  INV_X1 U5253 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10396) );
  INV_X1 U5254 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7684) );
  INV_X4 U5255 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NAND2_X1 U5256 ( .A1(n5313), .A2(n5312), .ZN(n5049) );
  NAND2_X1 U5257 ( .A1(n5049), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5673) );
  NAND2_X1 U5258 ( .A1(n7141), .A2(n8047), .ZN(n7144) );
  NAND2_X1 U5259 ( .A1(n8815), .A2(n8824), .ZN(n5053) );
  NAND2_X1 U5260 ( .A1(n8832), .A2(n8834), .ZN(n5054) );
  NAND2_X1 U5261 ( .A1(n5055), .A2(n7580), .ZN(n10789) );
  NAND2_X1 U5262 ( .A1(n5055), .A2(n7417), .ZN(n10741) );
  OAI211_X2 U5263 ( .C1(n6702), .C2(n6703), .A(n5057), .B(n5056), .ZN(n6888)
         );
  NAND2_X2 U5264 ( .A1(n6729), .A2(n7958), .ZN(n6946) );
  NAND2_X2 U5265 ( .A1(n6729), .A2(n7966), .ZN(n6702) );
  NAND2_X2 U5266 ( .A1(n6279), .A2(n6278), .ZN(n6729) );
  NAND2_X1 U5267 ( .A1(n6537), .A2(n5713), .ZN(n5058) );
  NAND2_X1 U5268 ( .A1(n6537), .A2(n5713), .ZN(n6231) );
  NAND2_X1 U5269 ( .A1(n6672), .A2(n9446), .ZN(n6805) );
  INV_X4 U5270 ( .A(n5370), .ZN(n6031) );
  INV_X1 U5271 ( .A(n8169), .ZN(n8219) );
  AND2_X1 U5272 ( .A1(n7130), .A2(n7129), .ZN(n8045) );
  AND2_X1 U5273 ( .A1(n6039), .A2(n6034), .ZN(n6147) );
  OR2_X1 U5274 ( .A1(n9936), .A2(n9484), .ZN(n9624) );
  OR2_X1 U5275 ( .A1(n9958), .A2(n9754), .ZN(n9498) );
  OR2_X1 U5276 ( .A1(n10886), .A2(n9336), .ZN(n9544) );
  OR2_X1 U5277 ( .A1(n7400), .A2(n9670), .ZN(n5540) );
  NAND2_X1 U5278 ( .A1(n10749), .A2(n10750), .ZN(n5543) );
  BUF_X1 U5280 ( .A(n6946), .Z(n5137) );
  INV_X1 U5281 ( .A(n9289), .ZN(n5169) );
  NAND2_X1 U5282 ( .A1(n9936), .A2(n9484), .ZN(n9623) );
  INV_X1 U5283 ( .A(n6931), .ZN(n8400) );
  NAND2_X1 U5284 ( .A1(n8474), .A2(n5886), .ZN(n5370) );
  INV_X1 U5285 ( .A(n5369), .ZN(n6552) );
  AOI21_X1 U5286 ( .B1(n5236), .B2(n8178), .A(n5235), .ZN(n8183) );
  AND2_X1 U5287 ( .A1(n9091), .A2(n8177), .ZN(n5235) );
  NAND2_X1 U5288 ( .A1(n8163), .A2(n5237), .ZN(n5236) );
  INV_X1 U5289 ( .A(n6888), .ZN(n5318) );
  AND2_X1 U5290 ( .A1(n9593), .A2(n9489), .ZN(n9493) );
  NOR2_X1 U5291 ( .A1(n6198), .A2(n5449), .ZN(n5448) );
  INV_X1 U5292 ( .A(n6127), .ZN(n5449) );
  INV_X1 U5293 ( .A(SI_10_), .ZN(n10047) );
  NAND2_X2 U5294 ( .A1(n5686), .A2(n5685), .ZN(n5456) );
  INV_X1 U5295 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5685) );
  INV_X1 U5296 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5684) );
  INV_X1 U5297 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5687) );
  AND2_X1 U5298 ( .A1(n8313), .A2(n8312), .ZN(n8785) );
  NAND2_X1 U5299 ( .A1(n8848), .A2(n8310), .ZN(n5216) );
  OR2_X1 U5300 ( .A1(n9076), .A2(n8601), .ZN(n8307) );
  OR2_X1 U5301 ( .A1(n9091), .A2(n8935), .ZN(n8771) );
  OR2_X1 U5302 ( .A1(n9114), .A2(n8764), .ZN(n8295) );
  AND2_X1 U5303 ( .A1(n8289), .A2(n8288), .ZN(n8763) );
  AND2_X1 U5304 ( .A1(n8084), .A2(n8082), .ZN(n5338) );
  AOI21_X1 U5305 ( .B1(n10461), .B2(n10463), .A(n10464), .ZN(n6609) );
  INV_X1 U5306 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5360) );
  OAI21_X1 U5307 ( .B1(n6482), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7037) );
  NAND2_X1 U5308 ( .A1(n10876), .A2(n5169), .ZN(n9174) );
  NAND2_X1 U5309 ( .A1(n7780), .A2(n5169), .ZN(n7732) );
  NAND2_X1 U5310 ( .A1(n9736), .A2(n9750), .ZN(n5375) );
  NOR2_X1 U5311 ( .A1(n5095), .A2(n5377), .ZN(n5376) );
  NOR2_X1 U5312 ( .A1(n9738), .A2(n5379), .ZN(n5377) );
  OR2_X1 U5313 ( .A1(n9998), .A2(n9890), .ZN(n9548) );
  OR2_X1 U5314 ( .A1(n9755), .A2(n9958), .ZN(n9743) );
  NOR2_X1 U5315 ( .A1(n9636), .A2(n5542), .ZN(n5541) );
  INV_X1 U5316 ( .A(n7638), .ZN(n5542) );
  AND3_X1 U5317 ( .A1(n5521), .A2(n5633), .A3(n10200), .ZN(n5171) );
  INV_X1 U5318 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n10174) );
  AND2_X1 U5319 ( .A1(n5445), .A2(n5127), .ZN(n5444) );
  INV_X1 U5320 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n10397) );
  NAND2_X1 U5321 ( .A1(n5871), .A2(n5870), .ZN(n5988) );
  OR2_X1 U5322 ( .A1(n8015), .A2(n10291), .ZN(n8005) );
  AOI21_X1 U5323 ( .B1(n5487), .B2(n5183), .A(n5486), .ZN(n5485) );
  INV_X1 U5324 ( .A(n8538), .ZN(n5486) );
  NAND2_X1 U5325 ( .A1(n8607), .A2(n8608), .ZN(n8606) );
  AND2_X1 U5326 ( .A1(n8550), .A2(n6382), .ZN(n6719) );
  NAND2_X1 U5327 ( .A1(n8550), .A2(n9154), .ZN(n6707) );
  NAND2_X1 U5328 ( .A1(n6383), .A2(n9154), .ZN(n6718) );
  NAND2_X1 U5329 ( .A1(n5515), .A2(n5620), .ZN(n5514) );
  AOI21_X1 U5330 ( .B1(n8801), .B2(n8191), .A(n7991), .ZN(n8787) );
  NAND2_X1 U5331 ( .A1(n5332), .A2(n8302), .ZN(n8903) );
  OAI21_X1 U5332 ( .B1(n8926), .B2(n5419), .A(n5417), .ZN(n8894) );
  INV_X1 U5333 ( .A(n5420), .ZN(n5419) );
  AOI21_X1 U5334 ( .B1(n5420), .B2(n8933), .A(n5418), .ZN(n5417) );
  INV_X1 U5335 ( .A(n8771), .ZN(n5418) );
  OR2_X1 U5336 ( .A1(n8251), .A2(n10640), .ZN(n6690) );
  INV_X1 U5337 ( .A(n6946), .ZN(n8135) );
  OAI22_X1 U5338 ( .A1(n7344), .A2(n7343), .B1(n10677), .B2(n8703), .ZN(n7380)
         );
  INV_X1 U5339 ( .A(n8806), .ZN(n9012) );
  AND2_X1 U5340 ( .A1(n6278), .A2(n6522), .ZN(n9014) );
  INV_X1 U5341 ( .A(n10797), .ZN(n9017) );
  NAND2_X1 U5342 ( .A1(n8213), .A2(n8212), .ZN(n9059) );
  NAND2_X1 U5343 ( .A1(n8252), .A2(n8314), .ZN(n10640) );
  NOR2_X1 U5344 ( .A1(n5666), .A2(n5665), .ZN(n5667) );
  INV_X1 U5345 ( .A(n5820), .ZN(n5314) );
  XNOR2_X1 U5346 ( .A(n5811), .B(n5810), .ZN(n6279) );
  OR2_X1 U5347 ( .A1(n5809), .A2(n9146), .ZN(n5811) );
  XNOR2_X1 U5348 ( .A(n5808), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8284) );
  XNOR2_X1 U5349 ( .A(n5513), .B(n6486), .ZN(n6513) );
  INV_X1 U5350 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6486) );
  OAI21_X1 U5351 ( .B1(n6484), .B2(P2_IR_REG_19__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5513) );
  OR2_X1 U5352 ( .A1(n9166), .A2(n9165), .ZN(n9255) );
  NAND2_X1 U5353 ( .A1(n9958), .A2(n5169), .ZN(n9229) );
  NAND2_X1 U5354 ( .A1(n10886), .A2(n5169), .ZN(n9169) );
  INV_X1 U5355 ( .A(n7265), .ZN(n5164) );
  NOR2_X1 U5356 ( .A1(n5165), .A2(n5158), .ZN(n5157) );
  NOR2_X1 U5357 ( .A1(n7265), .A2(n7184), .ZN(n5165) );
  INV_X1 U5358 ( .A(n7174), .ZN(n5158) );
  NAND2_X1 U5359 ( .A1(n6152), .A2(n6151), .ZN(n6154) );
  AND2_X1 U5360 ( .A1(n5304), .A2(n5303), .ZN(n9600) );
  INV_X1 U5361 ( .A(n9595), .ZN(n5303) );
  INV_X1 U5362 ( .A(n9653), .ZN(n9597) );
  AND2_X1 U5363 ( .A1(n9684), .A2(n9583), .ZN(n9686) );
  NOR2_X1 U5364 ( .A1(n9714), .A2(n5555), .ZN(n5554) );
  INV_X1 U5365 ( .A(n8435), .ZN(n5555) );
  AND4_X1 U5366 ( .A1(n6606), .A2(n6605), .A3(n6604), .A4(n6603), .ZN(n9723)
         );
  AOI21_X1 U5367 ( .B1(n9738), .B2(n5526), .A(n5106), .ZN(n5525) );
  OR2_X1 U5368 ( .A1(n5072), .A2(n8456), .ZN(n5380) );
  AOI21_X1 U5369 ( .B1(n9914), .B2(n9915), .A(n7783), .ZN(n7784) );
  OAI21_X1 U5370 ( .B1(n7750), .B2(n7749), .A(n9530), .ZN(n7788) );
  AOI21_X1 U5371 ( .B1(n5534), .B2(n5536), .A(n5067), .ZN(n5533) );
  NAND2_X1 U5372 ( .A1(n5403), .A2(n5401), .ZN(n7398) );
  AOI21_X1 U5373 ( .B1(n5404), .B2(n5407), .A(n5402), .ZN(n5401) );
  NOR2_X1 U5374 ( .A1(n9513), .A2(n5405), .ZN(n5404) );
  NAND2_X1 U5375 ( .A1(n7011), .A2(n9634), .ZN(n7208) );
  NAND2_X1 U5376 ( .A1(n6666), .A2(n6665), .ZN(n6804) );
  NAND2_X1 U5377 ( .A1(n9430), .A2(n9429), .ZN(n9936) );
  NAND2_X1 U5378 ( .A1(n8444), .A2(n8443), .ZN(n9941) );
  XNOR2_X1 U5379 ( .A(n5564), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5888) );
  OR2_X1 U5380 ( .A1(n5885), .A2(n5884), .ZN(n5564) );
  INV_X1 U5381 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5651) );
  AOI21_X1 U5382 ( .B1(n5638), .B2(n10204), .A(n5884), .ZN(n5148) );
  NAND2_X1 U5383 ( .A1(n7887), .A2(n7886), .ZN(n7923) );
  NAND2_X1 U5384 ( .A1(n7691), .A2(n7690), .ZN(n7695) );
  NAND2_X1 U5385 ( .A1(n6052), .A2(n6051), .ZN(n6128) );
  BUF_X1 U5386 ( .A(n5712), .Z(n7966) );
  NAND2_X1 U5387 ( .A1(n9993), .A2(n5169), .ZN(n9192) );
  NAND2_X1 U5388 ( .A1(n8029), .A2(n5251), .ZN(n8035) );
  NAND2_X1 U5389 ( .A1(n5254), .A2(n5252), .ZN(n5251) );
  AOI21_X1 U5390 ( .B1(n5253), .B2(n8242), .A(n6732), .ZN(n5252) );
  AND2_X1 U5391 ( .A1(n5241), .A2(n5242), .ZN(n5246) );
  AOI21_X1 U5392 ( .B1(n5250), .B2(n5092), .A(n5243), .ZN(n5242) );
  NAND2_X1 U5393 ( .A1(n5240), .A2(n5245), .ZN(n5241) );
  NAND2_X1 U5394 ( .A1(n5244), .A2(n5066), .ZN(n5247) );
  NAND2_X1 U5395 ( .A1(n8046), .A2(n8047), .ZN(n5244) );
  AND2_X1 U5396 ( .A1(n8083), .A2(n8084), .ZN(n5277) );
  OAI21_X1 U5397 ( .B1(n9533), .B2(n9590), .A(n9907), .ZN(n5289) );
  NOR2_X1 U5398 ( .A1(n9532), .A2(n9558), .ZN(n5290) );
  NAND2_X1 U5399 ( .A1(n8148), .A2(n8147), .ZN(n8162) );
  NAND2_X1 U5400 ( .A1(n5239), .A2(n5238), .ZN(n5237) );
  NOR2_X1 U5401 ( .A1(n9096), .A2(n8920), .ZN(n5238) );
  INV_X1 U5402 ( .A(n8162), .ZN(n5239) );
  NOR2_X1 U5403 ( .A1(n5220), .A2(n5209), .ZN(n5208) );
  INV_X1 U5404 ( .A(n8310), .ZN(n5209) );
  AOI21_X1 U5405 ( .B1(n5219), .B2(n5214), .A(n5218), .ZN(n5213) );
  NOR2_X1 U5406 ( .A1(n5286), .A2(n5285), .ZN(n5284) );
  NAND2_X1 U5407 ( .A1(n9736), .A2(n9577), .ZN(n5285) );
  AOI21_X1 U5408 ( .B1(n9572), .B2(n5085), .A(n9578), .ZN(n5286) );
  INV_X1 U5409 ( .A(n8064), .ZN(n5341) );
  INV_X1 U5410 ( .A(n9493), .ZN(n9491) );
  OR2_X1 U5411 ( .A1(n9948), .A2(n9723), .ZN(n9495) );
  INV_X1 U5412 ( .A(n5456), .ZN(n5454) );
  NOR2_X1 U5413 ( .A1(n8483), .A2(n8617), .ZN(n5192) );
  NOR2_X1 U5414 ( .A1(n5266), .A2(n5265), .ZN(n5264) );
  INV_X1 U5415 ( .A(n8238), .ZN(n5266) );
  NAND2_X1 U5416 ( .A1(n8316), .A2(n8239), .ZN(n5265) );
  INV_X1 U5417 ( .A(n5264), .ZN(n5259) );
  INV_X1 U5418 ( .A(n8245), .ZN(n5261) );
  NOR2_X1 U5419 ( .A1(n5217), .A2(n8824), .ZN(n5215) );
  OR2_X1 U5420 ( .A1(n9065), .A2(n8602), .ZN(n8253) );
  NOR2_X1 U5421 ( .A1(n9076), .A2(n5329), .ZN(n5328) );
  INV_X1 U5422 ( .A(n5330), .ZN(n5329) );
  OR2_X1 U5423 ( .A1(n9103), .A2(n8769), .ZN(n8299) );
  AND2_X1 U5424 ( .A1(n8064), .A2(n9031), .ZN(n5222) );
  OAI21_X1 U5425 ( .B1(n5342), .B2(n5341), .A(n8067), .ZN(n5340) );
  AND2_X1 U5426 ( .A1(n7383), .A2(n8058), .ZN(n5342) );
  INV_X1 U5427 ( .A(n9103), .ZN(n8949) );
  AOI221_X1 U5428 ( .B1(P2_B_REG_SCAN_IN), .B2(n6479), .C1(n6478), .C2(n7702), 
        .A(n6492), .ZN(n6494) );
  INV_X1 U5429 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5273) );
  INV_X1 U5430 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6443) );
  INV_X1 U5431 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6445) );
  AND2_X1 U5432 ( .A1(n5517), .A2(n5516), .ZN(n5515) );
  INV_X1 U5433 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U5434 ( .A1(n9921), .A2(n5169), .ZN(n9161) );
  INV_X1 U5435 ( .A(n7728), .ZN(n5600) );
  INV_X1 U5436 ( .A(n7324), .ZN(n5570) );
  NAND2_X1 U5437 ( .A1(n7164), .A2(n5169), .ZN(n6650) );
  NAND2_X1 U5438 ( .A1(n9361), .A2(n9365), .ZN(n9224) );
  INV_X1 U5439 ( .A(n10449), .ZN(n5886) );
  NOR2_X1 U5440 ( .A1(n9948), .A2(n9941), .ZN(n5359) );
  NOR2_X1 U5441 ( .A1(n9709), .A2(n5375), .ZN(n5374) );
  AND2_X1 U5442 ( .A1(n9495), .A2(n9586), .ZN(n9714) );
  INV_X1 U5443 ( .A(n6602), .ZN(n8445) );
  OR2_X1 U5444 ( .A1(n9971), .A2(n9808), .ZN(n9791) );
  OR2_X1 U5445 ( .A1(n9978), .A2(n9820), .ZN(n8459) );
  INV_X1 U5446 ( .A(n9855), .ZN(n5551) );
  NOR2_X1 U5447 ( .A1(n9876), .A2(n5550), .ZN(n5549) );
  INV_X1 U5448 ( .A(n8333), .ZN(n5550) );
  OR2_X1 U5449 ( .A1(n9921), .A2(n9403), .ZN(n9534) );
  OR2_X1 U5450 ( .A1(n10815), .A2(n10754), .ZN(n9524) );
  OR2_X1 U5451 ( .A1(n7275), .A2(n7274), .ZN(n7277) );
  NAND2_X1 U5452 ( .A1(n6160), .A2(n5046), .ZN(n9448) );
  NAND2_X1 U5453 ( .A1(n6208), .A2(n9444), .ZN(n6212) );
  NOR2_X1 U5454 ( .A1(n5334), .A2(n5767), .ZN(n5518) );
  NOR2_X1 U5455 ( .A1(n5460), .A2(n5458), .ZN(n5457) );
  INV_X1 U5456 ( .A(n7934), .ZN(n5458) );
  INV_X1 U5457 ( .A(n7654), .ZN(n5472) );
  INV_X1 U5458 ( .A(SI_20_), .ZN(n10039) );
  NOR2_X1 U5459 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5628) );
  NOR2_X1 U5460 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5627) );
  INV_X1 U5461 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5631) );
  OAI21_X1 U5462 ( .B1(n6442), .B2(n5463), .A(n5461), .ZN(n7083) );
  INV_X1 U5463 ( .A(n5462), .ZN(n5461) );
  OAI21_X1 U5464 ( .B1(n5468), .B2(n5463), .A(n6984), .ZN(n5462) );
  INV_X1 U5465 ( .A(n5464), .ZN(n5463) );
  NOR2_X1 U5466 ( .A1(n6590), .A2(n5469), .ZN(n5468) );
  INV_X1 U5467 ( .A(n6441), .ZN(n5469) );
  INV_X1 U5468 ( .A(SI_15_), .ZN(n10252) );
  INV_X1 U5469 ( .A(n5448), .ZN(n5447) );
  AOI21_X1 U5470 ( .B1(n5446), .B2(n5448), .A(n5112), .ZN(n5445) );
  INV_X1 U5471 ( .A(n6051), .ZN(n5446) );
  NAND2_X1 U5472 ( .A1(n5452), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5198) );
  OAI21_X1 U5473 ( .B1(n7958), .B2(n5702), .A(n5701), .ZN(n5703) );
  NAND2_X1 U5474 ( .A1(n5713), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5701) );
  INV_X1 U5475 ( .A(n9195), .ZN(n5576) );
  OAI22_X1 U5476 ( .A1(n8566), .A2(n8527), .B1(n5183), .B2(n5103), .ZN(n5182)
         );
  NAND2_X1 U5477 ( .A1(n8591), .A2(n5176), .ZN(n5178) );
  NOR2_X1 U5478 ( .A1(n8516), .A2(n5177), .ZN(n5176) );
  INV_X1 U5479 ( .A(n8592), .ZN(n5177) );
  INV_X1 U5480 ( .A(n7439), .ZN(n5492) );
  NAND2_X1 U5481 ( .A1(n5485), .A2(n5481), .ZN(n5484) );
  AND2_X1 U5482 ( .A1(n8498), .A2(n8497), .ZN(n8504) );
  AND2_X1 U5483 ( .A1(n5175), .A2(n5174), .ZN(n7711) );
  NAND2_X1 U5484 ( .A1(n7708), .A2(n7707), .ZN(n5174) );
  NAND2_X1 U5485 ( .A1(n7710), .A2(n7709), .ZN(n5175) );
  NAND2_X1 U5486 ( .A1(n7711), .A2(n7712), .ZN(n7852) );
  NAND2_X1 U5487 ( .A1(n8572), .A2(n5079), .ZN(n8519) );
  INV_X1 U5488 ( .A(n8656), .ZN(n5511) );
  NAND2_X1 U5489 ( .A1(n6377), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8151) );
  OR2_X1 U5490 ( .A1(n8151), .A2(n10320), .ZN(n8167) );
  INV_X1 U5491 ( .A(n5494), .ZN(n5493) );
  AND2_X1 U5492 ( .A1(n5196), .A2(n5195), .ZN(n5490) );
  NOR2_X1 U5493 ( .A1(n7532), .A2(n7461), .ZN(n5195) );
  NAND2_X1 U5494 ( .A1(n5496), .A2(n5499), .ZN(n8607) );
  AOI21_X1 U5495 ( .B1(n8682), .B2(n8475), .A(n8480), .ZN(n5499) );
  NOR2_X1 U5496 ( .A1(n5500), .A2(n5498), .ZN(n5497) );
  NAND2_X1 U5497 ( .A1(n5505), .A2(n5507), .ZN(n7225) );
  INV_X1 U5498 ( .A(n5508), .ZN(n5507) );
  OAI21_X1 U5499 ( .B1(n6977), .B2(n7097), .A(n7101), .ZN(n5508) );
  NAND2_X1 U5500 ( .A1(n6976), .A2(n6977), .ZN(n7099) );
  AND2_X1 U5501 ( .A1(n6687), .A2(n6610), .ZN(n6613) );
  NAND2_X1 U5502 ( .A1(n7898), .A2(n7899), .ZN(n8477) );
  NAND2_X1 U5503 ( .A1(n5228), .A2(n5143), .ZN(n5437) );
  NAND2_X1 U5504 ( .A1(n8317), .A2(n8316), .ZN(n5232) );
  NAND2_X1 U5505 ( .A1(n5231), .A2(n5230), .ZN(n5229) );
  AND3_X1 U5506 ( .A1(n7998), .A2(n7997), .A3(n7996), .ZN(n8601) );
  AND4_X1 U5507 ( .A1(n8022), .A2(n8021), .A3(n8020), .A4(n8019), .ZN(n8772)
         );
  AND2_X1 U5508 ( .A1(n6520), .A2(n6519), .ZN(n5428) );
  OR2_X1 U5509 ( .A1(n6718), .A2(n6264), .ZN(n6520) );
  OR2_X1 U5510 ( .A1(n6707), .A2(n5200), .ZN(n6505) );
  INV_X1 U5511 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6444) );
  NAND2_X1 U5512 ( .A1(n8232), .A2(n8311), .ZN(n8781) );
  INV_X1 U5513 ( .A(n8311), .ZN(n5218) );
  NAND2_X1 U5514 ( .A1(n5216), .A2(n5212), .ZN(n5211) );
  NOR2_X1 U5515 ( .A1(n5218), .A2(n5214), .ZN(n5212) );
  INV_X1 U5516 ( .A(n8785), .ZN(n8783) );
  NAND2_X1 U5517 ( .A1(n5216), .A2(n5215), .ZN(n5221) );
  NOR2_X1 U5518 ( .A1(n9065), .A2(n8846), .ZN(n8838) );
  NAND2_X1 U5519 ( .A1(n8307), .A2(n8254), .ZN(n8870) );
  NAND2_X1 U5520 ( .A1(n8903), .A2(n8893), .ZN(n5225) );
  NAND2_X1 U5521 ( .A1(n8932), .A2(n8300), .ZN(n8917) );
  AND2_X1 U5522 ( .A1(n8916), .A2(n8770), .ZN(n5420) );
  NAND2_X1 U5523 ( .A1(n8946), .A2(n8299), .ZN(n8934) );
  INV_X1 U5524 ( .A(n5411), .ZN(n5410) );
  OAI21_X1 U5525 ( .B1(n5414), .B2(n5412), .A(n8766), .ZN(n5411) );
  NAND2_X1 U5526 ( .A1(n8973), .A2(n5415), .ZN(n5414) );
  INV_X1 U5527 ( .A(n5416), .ZN(n5415) );
  INV_X1 U5528 ( .A(n5336), .ZN(n5335) );
  OAI21_X1 U5529 ( .B1(n5338), .B2(n5337), .A(n8288), .ZN(n5336) );
  AND2_X1 U5530 ( .A1(n8292), .A2(n8291), .ZN(n8993) );
  NOR2_X1 U5531 ( .A1(n8989), .A2(n8993), .ZN(n8988) );
  OR2_X1 U5532 ( .A1(n9005), .A2(n9123), .ZN(n9003) );
  NAND2_X1 U5533 ( .A1(n7871), .A2(n5338), .ZN(n8287) );
  OAI21_X1 U5534 ( .B1(n7811), .B2(n8077), .A(n8079), .ZN(n7870) );
  CLKBUF_X1 U5535 ( .A(n7823), .Z(n7582) );
  AND2_X1 U5536 ( .A1(n6755), .A2(n8246), .ZN(n10797) );
  NAND2_X1 U5537 ( .A1(n8263), .A2(n6965), .ZN(n7130) );
  NAND2_X1 U5538 ( .A1(n5429), .A2(n7985), .ZN(n9054) );
  NAND2_X1 U5539 ( .A1(n8441), .A2(n8211), .ZN(n5429) );
  NAND2_X1 U5540 ( .A1(n8166), .A2(n8165), .ZN(n9091) );
  NAND2_X1 U5541 ( .A1(n8094), .A2(n8093), .ZN(n9119) );
  OR2_X1 U5542 ( .A1(n7089), .A2(n6702), .ZN(n7094) );
  INV_X1 U5543 ( .A(n6888), .ZN(n10656) );
  NAND2_X1 U5544 ( .A1(n6615), .A2(n6526), .ZN(n10860) );
  NOR2_X1 U5545 ( .A1(n6493), .A2(n6609), .ZN(n6530) );
  NOR2_X1 U5546 ( .A1(n7929), .A2(n6494), .ZN(n10461) );
  OR2_X1 U5547 ( .A1(n5945), .A2(n9146), .ZN(n5942) );
  NOR2_X1 U5548 ( .A1(n5812), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n5424) );
  OR2_X1 U5549 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n5812) );
  NOR2_X1 U5550 ( .A1(n5423), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n5312) );
  INV_X1 U5551 ( .A(n5807), .ZN(n5313) );
  INV_X1 U5552 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6483) );
  INV_X1 U5553 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6450) );
  NAND2_X1 U5554 ( .A1(n7634), .A2(n5169), .ZN(n7329) );
  NAND2_X1 U5555 ( .A1(n7175), .A2(n7174), .ZN(n5166) );
  AOI21_X1 U5556 ( .B1(n7325), .B2(n5568), .A(n5566), .ZN(n5565) );
  NAND2_X1 U5557 ( .A1(n5567), .A2(n7510), .ZN(n5566) );
  NAND2_X1 U5558 ( .A1(n5568), .A2(n5571), .ZN(n5567) );
  NAND2_X1 U5559 ( .A1(n10815), .A2(n5169), .ZN(n7521) );
  OR2_X1 U5560 ( .A1(n9226), .A2(n9227), .ZN(n5595) );
  NAND2_X1 U5561 ( .A1(n9265), .A2(n9268), .ZN(n5594) );
  NAND2_X1 U5562 ( .A1(n6545), .A2(n5574), .ZN(n6566) );
  AND2_X1 U5563 ( .A1(n6546), .A2(n6544), .ZN(n5574) );
  NAND2_X1 U5564 ( .A1(n5163), .A2(n7184), .ZN(n5162) );
  INV_X1 U5565 ( .A(n7179), .ZN(n5163) );
  AND2_X1 U5566 ( .A1(n7179), .A2(n5583), .ZN(n5582) );
  INV_X1 U5567 ( .A(n7184), .ZN(n5583) );
  AND2_X1 U5568 ( .A1(n6042), .A2(n6041), .ZN(n6082) );
  INV_X1 U5569 ( .A(n5167), .ZN(n6036) );
  OAI21_X1 U5570 ( .B1(n6855), .B2(n9289), .A(n5168), .ZN(n5167) );
  NAND2_X1 U5571 ( .A1(n7723), .A2(n7722), .ZN(n7780) );
  OR2_X1 U5572 ( .A1(n7730), .A2(n7729), .ZN(n5601) );
  NAND2_X1 U5573 ( .A1(n9971), .A2(n5169), .ZN(n9214) );
  NAND2_X1 U5574 ( .A1(n7641), .A2(n5169), .ZN(n7495) );
  AND4_X1 U5575 ( .A1(n5912), .A2(n5911), .A3(n5910), .A4(n5909), .ZN(n7198)
         );
  NAND2_X1 U5576 ( .A1(n9422), .A2(n9421), .ZN(n9593) );
  NOR2_X1 U5577 ( .A1(n9936), .A2(n5358), .ZN(n5357) );
  INV_X1 U5578 ( .A(n5359), .ZN(n5358) );
  OR2_X1 U5579 ( .A1(n9948), .A2(n8440), .ZN(n5556) );
  NAND2_X1 U5580 ( .A1(n9729), .A2(n9717), .ZN(n9706) );
  XOR2_X1 U5581 ( .A(n9714), .B(n9713), .Z(n9949) );
  NAND2_X1 U5582 ( .A1(n8436), .A2(n8435), .ZN(n9713) );
  AND2_X1 U5583 ( .A1(n5372), .A2(n5376), .ZN(n9724) );
  INV_X1 U5584 ( .A(n5375), .ZN(n5373) );
  NOR2_X1 U5585 ( .A1(n8416), .A2(n5529), .ZN(n5528) );
  INV_X1 U5586 ( .A(n8402), .ZN(n5529) );
  NAND2_X1 U5587 ( .A1(n9350), .A2(n9741), .ZN(n5530) );
  OAI21_X1 U5588 ( .B1(n9794), .B2(n9792), .A(n9791), .ZN(n9774) );
  OAI21_X1 U5589 ( .B1(n9782), .B2(n8388), .A(n8389), .ZN(n9765) );
  NAND2_X1 U5590 ( .A1(n9891), .A2(n5549), .ZN(n5548) );
  AND2_X1 U5591 ( .A1(n9553), .A2(n9554), .ZN(n9855) );
  AND4_X1 U5592 ( .A1(n7764), .A2(n7763), .A3(n7762), .A4(n7761), .ZN(n9887)
         );
  NAND2_X1 U5593 ( .A1(n7755), .A2(n5081), .ZN(n8455) );
  NAND2_X1 U5594 ( .A1(n7779), .A2(n7778), .ZN(n7787) );
  OAI21_X1 U5595 ( .B1(n10752), .B2(n7649), .A(n9526), .ZN(n7750) );
  OR2_X1 U5596 ( .A1(n7396), .A2(n5537), .ZN(n5536) );
  INV_X1 U5597 ( .A(n7394), .ZN(n5537) );
  NAND2_X1 U5598 ( .A1(n5406), .A2(n9462), .ZN(n10713) );
  NAND2_X1 U5599 ( .A1(n5281), .A2(n9505), .ZN(n7204) );
  OAI211_X1 U5600 ( .C1(n7001), .C2(n5282), .A(n5383), .B(n9457), .ZN(n5281)
         );
  NAND3_X1 U5601 ( .A1(n5384), .A2(n5385), .A3(n9459), .ZN(n5383) );
  AND2_X1 U5602 ( .A1(n7009), .A2(n7008), .ZN(n5552) );
  AND2_X1 U5603 ( .A1(n9505), .A2(n9507), .ZN(n9632) );
  NAND2_X1 U5604 ( .A1(n6846), .A2(n6214), .ZN(n9450) );
  NAND2_X1 U5605 ( .A1(n6212), .A2(n6213), .ZN(n6847) );
  NAND2_X1 U5606 ( .A1(n6847), .A2(n6848), .ZN(n6846) );
  NAND2_X1 U5607 ( .A1(n10452), .A2(n9598), .ZN(n10753) );
  OR2_X1 U5608 ( .A1(n10452), .A2(n6091), .ZN(n10755) );
  OR2_X1 U5609 ( .A1(n10817), .A2(n9597), .ZN(n6061) );
  OR2_X1 U5610 ( .A1(n9949), .A2(n10831), .ZN(n5395) );
  INV_X1 U5611 ( .A(n9743), .ZN(n8467) );
  OR2_X1 U5612 ( .A1(n6537), .A2(n10627), .ZN(n5558) );
  OR2_X1 U5613 ( .A1(n5058), .A2(n6703), .ZN(n5559) );
  AND4_X1 U5614 ( .A1(n5614), .A2(n5391), .A3(n5387), .A4(n5518), .ZN(n5885)
         );
  AND2_X1 U5615 ( .A1(n5389), .A2(n5390), .ZN(n5387) );
  INV_X1 U5616 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5389) );
  NAND2_X1 U5617 ( .A1(n5639), .A2(n5615), .ZN(n5560) );
  INV_X1 U5618 ( .A(n5148), .ZN(n5636) );
  AND2_X1 U5619 ( .A1(n5476), .A2(n7694), .ZN(n5475) );
  INV_X1 U5620 ( .A(n7697), .ZN(n5476) );
  NAND2_X1 U5621 ( .A1(n7472), .A2(n7471), .ZN(n7655) );
  NAND2_X1 U5622 ( .A1(n7313), .A2(n5470), .ZN(n7472) );
  NOR2_X1 U5623 ( .A1(n7315), .A2(n5471), .ZN(n5470) );
  INV_X1 U5624 ( .A(n7312), .ZN(n5471) );
  INV_X1 U5625 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5626) );
  NAND2_X1 U5626 ( .A1(n5172), .A2(n5059), .ZN(n5520) );
  NOR2_X1 U5627 ( .A1(n6593), .A2(n5467), .ZN(n5464) );
  NAND2_X1 U5628 ( .A1(n6442), .A2(n5468), .ZN(n5465) );
  NAND2_X1 U5629 ( .A1(n6047), .A2(n6046), .ZN(n6052) );
  NAND2_X1 U5630 ( .A1(n5798), .A2(n5797), .ZN(n5819) );
  OAI21_X1 U5631 ( .B1(n5709), .B2(n5433), .A(n5737), .ZN(n5430) );
  OAI21_X1 U5632 ( .B1(n5710), .B2(n5433), .A(n5740), .ZN(n5432) );
  NAND2_X1 U5633 ( .A1(n5579), .A2(n5083), .ZN(n5578) );
  INV_X1 U5634 ( .A(n9333), .ZN(n5579) );
  INV_X1 U5635 ( .A(n9320), .ZN(n9178) );
  NAND2_X1 U5636 ( .A1(n6479), .A2(n5679), .ZN(n6490) );
  NAND2_X1 U5637 ( .A1(n8574), .A2(n8573), .ZN(n8572) );
  OR2_X1 U5638 ( .A1(n7440), .A2(n5493), .ZN(n5491) );
  NAND2_X1 U5639 ( .A1(n5502), .A2(n5501), .ZN(n6903) );
  NAND2_X1 U5640 ( .A1(n5503), .A2(n5504), .ZN(n5502) );
  NAND2_X1 U5641 ( .A1(n6837), .A2(n6768), .ZN(n5501) );
  NOR2_X1 U5642 ( .A1(n6769), .A2(n6763), .ZN(n5503) );
  INV_X1 U5643 ( .A(n8705), .ZN(n6961) );
  AND2_X1 U5644 ( .A1(n7987), .A2(n7986), .ZN(n8801) );
  OR2_X1 U5645 ( .A1(n6778), .A2(n6779), .ZN(n5504) );
  AND3_X1 U5646 ( .A1(n8008), .A2(n8007), .A3(n8006), .ZN(n8773) );
  INV_X1 U5647 ( .A(n8707), .ZN(n6839) );
  AND2_X1 U5648 ( .A1(n5504), .A2(n6762), .ZN(n6838) );
  INV_X1 U5649 ( .A(n9013), .ZN(n8761) );
  NAND2_X1 U5650 ( .A1(n8322), .A2(n8323), .ZN(n5267) );
  NOR3_X1 U5651 ( .A1(n8285), .A2(n8284), .A3(n8283), .ZN(n8321) );
  NAND2_X1 U5652 ( .A1(n6490), .A2(n10583), .ZN(n10462) );
  NAND2_X1 U5653 ( .A1(n6523), .A2(n6522), .ZN(n8806) );
  XNOR2_X1 U5654 ( .A(n5806), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8324) );
  INV_X1 U5655 ( .A(n6514), .ZN(n6780) );
  AND2_X1 U5656 ( .A1(n5139), .A2(n5138), .ZN(n9062) );
  AOI22_X1 U5657 ( .A1(n8827), .A2(n9014), .B1(n9012), .B2(n8826), .ZN(n5138)
         );
  NAND2_X1 U5658 ( .A1(n8828), .A2(n9017), .ZN(n5139) );
  NAND2_X1 U5659 ( .A1(n8107), .A2(n8106), .ZN(n9114) );
  NAND2_X1 U5660 ( .A1(n10811), .A2(n10803), .ZN(n9008) );
  INV_X1 U5661 ( .A(n8793), .ZN(n9020) );
  NAND2_X2 U5662 ( .A1(n6695), .A2(n8981), .ZN(n10811) );
  NAND2_X1 U5663 ( .A1(n8392), .A2(n8391), .ZN(n9966) );
  OAI21_X1 U5664 ( .B1(n9292), .B2(n5151), .A(n9298), .ZN(n5150) );
  NAND2_X1 U5665 ( .A1(n9283), .A2(n9376), .ZN(n5151) );
  NAND2_X1 U5666 ( .A1(n7393), .A2(n5169), .ZN(n7186) );
  INV_X1 U5667 ( .A(n5605), .ZN(n5603) );
  AND4_X1 U5668 ( .A1(n8345), .A2(n8344), .A3(n8343), .A4(n8342), .ZN(n9890)
         );
  NAND2_X1 U5669 ( .A1(n8332), .A2(n8331), .ZN(n10886) );
  NAND2_X1 U5670 ( .A1(n8337), .A2(n8336), .ZN(n9998) );
  INV_X1 U5671 ( .A(n6208), .ZN(n9445) );
  AND4_X1 U5672 ( .A1(n8425), .A2(n8424), .A3(n8423), .A4(n8422), .ZN(n9754)
         );
  OR2_X1 U5673 ( .A1(n8085), .A2(n6231), .ZN(n7758) );
  INV_X1 U5674 ( .A(n10755), .ZN(n9912) );
  OAI21_X1 U5675 ( .B1(n9603), .B2(n9604), .A(n5295), .ZN(n5294) );
  NAND2_X1 U5676 ( .A1(n9602), .A2(n9601), .ZN(n9603) );
  NOR2_X1 U5677 ( .A1(n9656), .A2(n7264), .ZN(n5295) );
  AOI21_X1 U5678 ( .B1(n9658), .B2(n7264), .A(n9663), .ZN(n5293) );
  INV_X1 U5679 ( .A(n9593), .ZN(n9930) );
  AOI21_X1 U5680 ( .B1(n9695), .B2(n10758), .A(n9694), .ZN(n9940) );
  NAND2_X1 U5681 ( .A1(n9693), .A2(n9692), .ZN(n9694) );
  XNOR2_X1 U5682 ( .A(n9688), .B(n9648), .ZN(n9695) );
  XNOR2_X1 U5683 ( .A(n9704), .B(n9703), .ZN(n9935) );
  OR2_X1 U5684 ( .A1(n9701), .A2(n9712), .ZN(n5622) );
  NAND2_X1 U5685 ( .A1(n5400), .A2(n5397), .ZN(n9946) );
  INV_X1 U5686 ( .A(n5398), .ZN(n5397) );
  OR2_X1 U5687 ( .A1(n9711), .A2(n9888), .ZN(n5400) );
  OAI21_X1 U5688 ( .B1(n9712), .B2(n10753), .A(n5399), .ZN(n5398) );
  NAND2_X1 U5689 ( .A1(n10783), .A2(n6629), .ZN(n10780) );
  AND2_X1 U5690 ( .A1(n10783), .A2(n6627), .ZN(n10773) );
  INV_X1 U5691 ( .A(n9812), .ZN(n9760) );
  AND2_X1 U5692 ( .A1(n10783), .A2(n6631), .ZN(n10772) );
  AND2_X1 U5693 ( .A1(n6016), .A2(n6015), .ZN(n10442) );
  NAND2_X1 U5694 ( .A1(n6039), .A2(n5756), .ZN(n10441) );
  OAI21_X1 U5695 ( .B1(n8256), .B2(n8314), .A(n6879), .ZN(n5253) );
  NAND2_X1 U5696 ( .A1(n8026), .A2(n5255), .ZN(n5254) );
  INV_X1 U5697 ( .A(n8046), .ZN(n5240) );
  NOR2_X1 U5698 ( .A1(n5248), .A2(n8268), .ZN(n5245) );
  INV_X1 U5699 ( .A(n8057), .ZN(n5243) );
  AOI21_X1 U5700 ( .B1(n8035), .B2(n8032), .A(n8031), .ZN(n8037) );
  NAND2_X1 U5701 ( .A1(n5302), .A2(n5300), .ZN(n5299) );
  NOR2_X1 U5702 ( .A1(n10712), .A2(n5301), .ZN(n5300) );
  NAND2_X1 U5703 ( .A1(n10713), .A2(n9558), .ZN(n5302) );
  AND2_X1 U5704 ( .A1(n5408), .A2(n9590), .ZN(n5301) );
  OAI21_X1 U5705 ( .B1(n8048), .B2(n5247), .A(n5246), .ZN(n5249) );
  NAND2_X1 U5706 ( .A1(n5279), .A2(n5277), .ZN(n5276) );
  AOI21_X1 U5707 ( .B1(n5275), .B2(n5277), .A(n5278), .ZN(n5274) );
  NAND2_X1 U5708 ( .A1(n8763), .A2(n8091), .ZN(n5278) );
  NAND2_X1 U5709 ( .A1(n8080), .A2(n8270), .ZN(n5275) );
  NAND2_X1 U5710 ( .A1(n5297), .A2(n5296), .ZN(n9514) );
  OAI21_X1 U5711 ( .B1(n5299), .B2(n5090), .A(n5298), .ZN(n5297) );
  NAND2_X1 U5712 ( .A1(n5299), .A2(n5093), .ZN(n5296) );
  NOR2_X1 U5713 ( .A1(n9513), .A2(n9558), .ZN(n5298) );
  NAND2_X1 U5714 ( .A1(n5288), .A2(n5287), .ZN(n9547) );
  AND2_X1 U5715 ( .A1(n9641), .A2(n9543), .ZN(n5287) );
  OAI21_X1 U5716 ( .B1(n5290), .B2(n5289), .A(n5111), .ZN(n5288) );
  NAND2_X1 U5717 ( .A1(n5207), .A2(n5065), .ZN(n5434) );
  OR2_X1 U5718 ( .A1(n9108), .A2(n8767), .ZN(n8297) );
  OAI21_X1 U5719 ( .B1(n5284), .B2(n5283), .A(n5109), .ZN(n9582) );
  NAND2_X1 U5720 ( .A1(n9580), .A2(n9579), .ZN(n5283) );
  INV_X1 U5721 ( .A(n9498), .ZN(n5378) );
  NOR2_X1 U5722 ( .A1(n7922), .A2(n5474), .ZN(n5473) );
  INV_X1 U5723 ( .A(n7886), .ZN(n5474) );
  INV_X1 U5724 ( .A(n5334), .ZN(n5333) );
  INV_X1 U5725 ( .A(SI_19_), .ZN(n10244) );
  INV_X1 U5726 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n10391) );
  INV_X1 U5727 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n10192) );
  INV_X1 U5728 ( .A(SI_13_), .ZN(n10255) );
  INV_X1 U5729 ( .A(SI_9_), .ZN(n10263) );
  NOR2_X1 U5730 ( .A1(n5867), .A2(n5440), .ZN(n5439) );
  INV_X1 U5731 ( .A(n5818), .ZN(n5440) );
  INV_X1 U5732 ( .A(n8682), .ZN(n5500) );
  INV_X1 U5733 ( .A(n7899), .ZN(n5498) );
  NOR2_X1 U5734 ( .A1(n7097), .A2(n6973), .ZN(n5506) );
  INV_X1 U5735 ( .A(n8084), .ZN(n8273) );
  NAND2_X1 U5736 ( .A1(n8315), .A2(n9046), .ZN(n5231) );
  NOR2_X1 U5737 ( .A1(n8694), .A2(n8314), .ZN(n5230) );
  OR2_X1 U5738 ( .A1(n9054), .A2(n8787), .ZN(n8232) );
  INV_X1 U5739 ( .A(n5215), .ZN(n5214) );
  NOR2_X1 U5740 ( .A1(n9081), .A2(n9086), .ZN(n5330) );
  NOR2_X1 U5741 ( .A1(n9003), .A2(n5323), .ZN(n8927) );
  NAND2_X1 U5742 ( .A1(n5324), .A2(n8949), .ZN(n5323) );
  NOR2_X1 U5743 ( .A1(n5325), .A2(n9108), .ZN(n5324) );
  INV_X1 U5744 ( .A(n8993), .ZN(n5412) );
  INV_X1 U5745 ( .A(n5414), .ZN(n5413) );
  INV_X1 U5746 ( .A(n8286), .ZN(n5337) );
  NOR2_X1 U5747 ( .A1(n7821), .A2(n10804), .ZN(n5320) );
  OR2_X1 U5748 ( .A1(n6962), .A2(n8042), .ZN(n7135) );
  OR2_X1 U5749 ( .A1(n6879), .A2(n6732), .ZN(n6881) );
  NAND2_X1 U5750 ( .A1(n8911), .A2(n5063), .ZN(n8846) );
  AND2_X1 U5751 ( .A1(n7869), .A2(n7822), .ZN(n5425) );
  NAND4_X1 U5752 ( .A1(n10639), .A2(n6832), .A3(n10656), .A4(n5316), .ZN(n6962) );
  AND2_X1 U5753 ( .A1(n6795), .A2(n5317), .ZN(n5316) );
  INV_X1 U5754 ( .A(n10640), .ZN(n6526) );
  AND2_X1 U5755 ( .A1(n5319), .A2(n6832), .ZN(n6875) );
  NOR2_X1 U5756 ( .A1(n6756), .A2(n6888), .ZN(n5319) );
  NAND2_X1 U5757 ( .A1(n6832), .A2(n10639), .ZN(n6873) );
  NAND2_X1 U5758 ( .A1(n5314), .A2(n5227), .ZN(n5943) );
  NAND2_X1 U5759 ( .A1(n5669), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5680) );
  INV_X1 U5760 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5422) );
  NAND2_X1 U5761 ( .A1(n7206), .A2(n5169), .ZN(n6925) );
  NAND2_X1 U5762 ( .A1(n9978), .A2(n5169), .ZN(n9207) );
  NAND2_X1 U5763 ( .A1(n6035), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5168) );
  INV_X1 U5764 ( .A(n9275), .ZN(n5613) );
  NAND2_X1 U5765 ( .A1(n9981), .A2(n5169), .ZN(n9200) );
  MUX2_X1 U5766 ( .A(n9605), .B(n9494), .S(n9590), .Z(n9595) );
  NAND2_X1 U5767 ( .A1(n5309), .A2(n5307), .ZN(n5306) );
  NOR2_X1 U5768 ( .A1(n5308), .A2(n9558), .ZN(n5307) );
  OR2_X1 U5769 ( .A1(n9589), .A2(n9618), .ZN(n5309) );
  INV_X1 U5770 ( .A(n9623), .ZN(n5308) );
  OR2_X1 U5771 ( .A1(n9941), .A2(n9712), .ZN(n9684) );
  NOR2_X1 U5772 ( .A1(n9736), .A2(n5524), .ZN(n5523) );
  INV_X1 U5773 ( .A(n5528), .ZN(n5524) );
  INV_X1 U5774 ( .A(n5530), .ZN(n5526) );
  INV_X1 U5775 ( .A(n9566), .ZN(n5364) );
  NOR2_X1 U5776 ( .A1(n9993), .A2(n9987), .ZN(n5348) );
  AND2_X1 U5777 ( .A1(n7759), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7767) );
  NOR2_X1 U5778 ( .A1(n9921), .A2(n7780), .ZN(n5354) );
  INV_X1 U5779 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5958) );
  INV_X1 U5780 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5980) );
  INV_X1 U5781 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7274) );
  INV_X1 U5782 ( .A(n9462), .ZN(n5405) );
  INV_X1 U5783 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7189) );
  OR2_X1 U5784 ( .A1(n7190), .A2(n7189), .ZN(n7275) );
  OR2_X1 U5785 ( .A1(n5408), .A2(n7205), .ZN(n5407) );
  INV_X1 U5786 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5906) );
  INV_X1 U5787 ( .A(n9456), .ZN(n5385) );
  NAND2_X1 U5788 ( .A1(n6667), .A2(n10662), .ZN(n9453) );
  NAND2_X1 U5789 ( .A1(n9766), .A2(n9350), .ZN(n9755) );
  AND2_X1 U5790 ( .A1(n9871), .A2(n9862), .ZN(n9863) );
  XNOR2_X1 U5791 ( .A(n7960), .B(n7959), .ZN(n7981) );
  AND2_X1 U5792 ( .A1(n5616), .A2(n5633), .ZN(n5614) );
  NOR2_X1 U5793 ( .A1(n5617), .A2(n5621), .ZN(n5616) );
  NAND2_X1 U5794 ( .A1(n10208), .A2(n10200), .ZN(n5617) );
  INV_X1 U5795 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5390) );
  NOR2_X1 U5796 ( .A1(n5621), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n5615) );
  AND2_X1 U5797 ( .A1(n7947), .A2(n7938), .ZN(n7946) );
  NAND2_X1 U5798 ( .A1(n7931), .A2(n7930), .ZN(n5459) );
  INV_X1 U5799 ( .A(SI_23_), .ZN(n10236) );
  INV_X1 U5800 ( .A(SI_12_), .ZN(n10254) );
  NAND2_X1 U5801 ( .A1(n5454), .A2(n5689), .ZN(n5453) );
  NAND2_X1 U5802 ( .A1(n5452), .A2(n5689), .ZN(n5451) );
  OR2_X1 U5803 ( .A1(n8214), .A2(n8567), .ZN(n8216) );
  OR2_X1 U5804 ( .A1(n8216), .A2(n10292), .ZN(n7987) );
  NAND2_X1 U5805 ( .A1(n6975), .A2(n6974), .ZN(n6976) );
  NAND2_X1 U5806 ( .A1(n7440), .A2(n7439), .ZN(n5495) );
  NAND2_X1 U5807 ( .A1(n7852), .A2(n7851), .ZN(n7853) );
  NAND2_X1 U5808 ( .A1(n6379), .A2(n6378), .ZN(n8015) );
  NAND2_X1 U5809 ( .A1(n5187), .A2(n5185), .ZN(n8655) );
  AOI21_X1 U5810 ( .B1(n5188), .B2(n5191), .A(n5186), .ZN(n5185) );
  INV_X1 U5811 ( .A(n8660), .ZN(n5186) );
  AOI21_X1 U5812 ( .B1(n5190), .B2(n5192), .A(n5189), .ZN(n5188) );
  INV_X1 U5813 ( .A(n8618), .ZN(n5189) );
  INV_X1 U5814 ( .A(n8608), .ZN(n5190) );
  INV_X1 U5815 ( .A(n5192), .ZN(n5191) );
  OR2_X1 U5816 ( .A1(n8120), .A2(n10117), .ZN(n8138) );
  AOI21_X1 U5817 ( .B1(n6615), .B2(n6522), .A(n6491), .ZN(n6771) );
  OR2_X1 U5818 ( .A1(n7873), .A2(n6374), .ZN(n8095) );
  AOI21_X1 U5819 ( .B1(n8245), .B2(n5263), .A(n8244), .ZN(n8249) );
  NAND2_X1 U5820 ( .A1(n8547), .A2(n5256), .ZN(n8251) );
  NAND2_X1 U5821 ( .A1(n5258), .A2(n5260), .ZN(n8250) );
  NOR2_X1 U5822 ( .A1(n8244), .A2(n5259), .ZN(n5257) );
  NAND2_X1 U5823 ( .A1(n5668), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5806) );
  INV_X1 U5824 ( .A(n5672), .ZN(n5668) );
  AND2_X1 U5825 ( .A1(n8209), .A2(n8208), .ZN(n8602) );
  NOR2_X1 U5826 ( .A1(n5514), .A2(n5270), .ZN(n6447) );
  AOI21_X1 U5827 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n8720), .A(n8719), .ZN(
        n8723) );
  NAND2_X1 U5828 ( .A1(n5315), .A2(n9048), .ZN(n8792) );
  NOR2_X1 U5829 ( .A1(n8792), .A2(n8757), .ZN(n8753) );
  OR2_X1 U5830 ( .A1(n9071), .A2(n8672), .ZN(n8833) );
  OR2_X1 U5831 ( .A1(n8189), .A2(n10309), .ZN(n8202) );
  NAND2_X1 U5832 ( .A1(n8253), .A2(n8309), .ZN(n8834) );
  OR2_X1 U5833 ( .A1(n9076), .A2(n8775), .ZN(n5147) );
  NAND2_X1 U5834 ( .A1(n8911), .A2(n5328), .ZN(n8862) );
  NAND2_X1 U5835 ( .A1(n8911), .A2(n8901), .ZN(n8895) );
  AND2_X1 U5836 ( .A1(n8928), .A2(n8915), .ZN(n8911) );
  AND2_X1 U5837 ( .A1(n8771), .A2(n8176), .ZN(n8916) );
  AND2_X1 U5838 ( .A1(n8927), .A2(n8931), .ZN(n8928) );
  NAND2_X1 U5839 ( .A1(n8926), .A2(n8925), .ZN(n8924) );
  OR2_X1 U5840 ( .A1(n9114), .A2(n9119), .ZN(n5325) );
  NOR2_X1 U5841 ( .A1(n9003), .A2(n5322), .ZN(n8957) );
  INV_X1 U5842 ( .A(n5324), .ZN(n5322) );
  OR2_X1 U5843 ( .A1(n7564), .A2(n10319), .ZN(n7873) );
  NAND2_X1 U5844 ( .A1(n10793), .A2(n5320), .ZN(n7817) );
  NAND2_X1 U5845 ( .A1(n10793), .A2(n10794), .ZN(n10791) );
  OR2_X1 U5846 ( .A1(n7373), .A2(n10080), .ZN(n7539) );
  INV_X1 U5847 ( .A(n5340), .ZN(n5339) );
  NOR2_X1 U5848 ( .A1(n9027), .A2(n7441), .ZN(n7429) );
  AND2_X1 U5849 ( .A1(n7429), .A2(n10742), .ZN(n10793) );
  NAND2_X1 U5850 ( .A1(n7418), .A2(n8064), .ZN(n7571) );
  OR2_X1 U5851 ( .A1(n9026), .A2(n9034), .ZN(n9027) );
  NAND2_X1 U5852 ( .A1(n9023), .A2(n9031), .ZN(n7382) );
  NAND2_X1 U5853 ( .A1(n7382), .A2(n5342), .ZN(n7418) );
  NOR2_X1 U5854 ( .A1(n7135), .A2(n8049), .ZN(n7340) );
  NAND2_X1 U5855 ( .A1(n5206), .A2(n8045), .ZN(n7344) );
  NAND2_X1 U5856 ( .A1(n6788), .A2(n6735), .ZN(n7131) );
  NAND2_X1 U5857 ( .A1(n6790), .A2(n6789), .ZN(n6788) );
  NAND2_X1 U5858 ( .A1(n6500), .A2(n10640), .ZN(n8979) );
  OR3_X1 U5859 ( .A1(n6689), .A2(n6688), .A3(n6687), .ZN(n6695) );
  INV_X1 U5860 ( .A(n8757), .ZN(n9046) );
  NAND2_X1 U5861 ( .A1(n8150), .A2(n8149), .ZN(n9096) );
  NAND2_X1 U5862 ( .A1(n8088), .A2(n8087), .ZN(n9123) );
  NAND2_X1 U5863 ( .A1(n5624), .A2(n5060), .ZN(n7409) );
  OR2_X1 U5864 ( .A1(n9032), .A2(n9031), .ZN(n5624) );
  INV_X1 U5865 ( .A(n8560), .ZN(n10692) );
  CLKBUF_X1 U5866 ( .A(n7338), .Z(n10681) );
  NAND2_X1 U5867 ( .A1(n8547), .A2(n6526), .ZN(n10862) );
  NAND2_X1 U5868 ( .A1(n8979), .A2(n10653), .ZN(n10866) );
  OR2_X1 U5869 ( .A1(n8251), .A2(n8324), .ZN(n10653) );
  OR2_X1 U5870 ( .A1(n6946), .A2(n5145), .ZN(n5311) );
  INV_X1 U5871 ( .A(n10862), .ZN(n10792) );
  XNOR2_X1 U5872 ( .A(n5678), .B(P2_IR_REG_25__SCAN_IN), .ZN(n6492) );
  NAND2_X1 U5873 ( .A1(n5680), .A2(n5361), .ZN(n5682) );
  AND2_X1 U5874 ( .A1(n6446), .A2(n5273), .ZN(n5271) );
  AND3_X1 U5875 ( .A1(n6445), .A2(n6444), .A3(n6443), .ZN(n6446) );
  AND2_X1 U5876 ( .A1(n5746), .A2(n5659), .ZN(n5787) );
  INV_X1 U5877 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5659) );
  NOR2_X1 U5878 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5509) );
  NOR2_X1 U5879 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5698) );
  AND2_X1 U5880 ( .A1(n5598), .A2(n9165), .ZN(n5597) );
  OR2_X1 U5881 ( .A1(n7730), .A2(n5073), .ZN(n5596) );
  OR2_X1 U5882 ( .A1(n5061), .A2(n5599), .ZN(n5598) );
  AOI21_X1 U5883 ( .B1(n5609), .B2(n5607), .A(n5606), .ZN(n5605) );
  INV_X1 U5884 ( .A(n9352), .ZN(n5606) );
  INV_X1 U5885 ( .A(n5612), .ZN(n5607) );
  NAND2_X1 U5886 ( .A1(n9998), .A2(n5169), .ZN(n9185) );
  NAND2_X1 U5887 ( .A1(n5591), .A2(n5592), .ZN(n9340) );
  AND2_X1 U5888 ( .A1(n5594), .A2(n9342), .ZN(n5591) );
  NAND2_X1 U5889 ( .A1(n7400), .A2(n5169), .ZN(n7271) );
  NAND2_X1 U5890 ( .A1(n9197), .A2(n5613), .ZN(n5612) );
  NOR2_X1 U5891 ( .A1(n9197), .A2(n5613), .ZN(n5610) );
  NOR2_X1 U5892 ( .A1(n7489), .A2(n7488), .ZN(n5571) );
  AND2_X1 U5893 ( .A1(n5570), .A2(n7489), .ZN(n5569) );
  NOR2_X1 U5894 ( .A1(n8341), .A2(n5895), .ZN(n8355) );
  OR2_X1 U5895 ( .A1(n8339), .A2(n8338), .ZN(n8341) );
  NAND2_X1 U5896 ( .A1(n7077), .A2(n5169), .ZN(n6570) );
  OAI21_X1 U5897 ( .B1(n5590), .B2(n9342), .A(n5113), .ZN(n5585) );
  NOR2_X1 U5898 ( .A1(n5590), .A2(n5587), .ZN(n5586) );
  INV_X1 U5899 ( .A(n9268), .ZN(n5587) );
  NAND2_X1 U5900 ( .A1(n9951), .A2(n5169), .ZN(n9237) );
  NAND2_X1 U5901 ( .A1(n9600), .A2(n9599), .ZN(n9602) );
  AND2_X1 U5902 ( .A1(n9930), .A2(n9677), .ZN(n9651) );
  NOR2_X1 U5903 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5629) );
  NOR2_X1 U5904 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5630) );
  NAND2_X1 U5905 ( .A1(n5553), .A2(n5097), .ZN(n9702) );
  AND2_X1 U5906 ( .A1(n8448), .A2(n8447), .ZN(n9294) );
  OR2_X1 U5907 ( .A1(n9742), .A2(n10755), .ZN(n5399) );
  NAND2_X1 U5908 ( .A1(n9751), .A2(n5374), .ZN(n5371) );
  AND2_X1 U5909 ( .A1(n9783), .A2(n9771), .ZN(n9766) );
  NAND2_X1 U5910 ( .A1(n9871), .A2(n5344), .ZN(n9810) );
  NOR2_X1 U5911 ( .A1(n9978), .A2(n5346), .ZN(n5344) );
  NAND2_X1 U5912 ( .A1(n5557), .A2(n8384), .ZN(n9782) );
  NAND2_X1 U5913 ( .A1(n9871), .A2(n5348), .ZN(n9839) );
  NOR2_X1 U5914 ( .A1(n9834), .A2(n9835), .ZN(n9833) );
  OAI21_X1 U5915 ( .B1(n9891), .B2(n5547), .A(n5544), .ZN(n9832) );
  AOI21_X1 U5916 ( .B1(n5546), .B2(n5545), .A(n5084), .ZN(n5544) );
  INV_X1 U5917 ( .A(n5549), .ZN(n5545) );
  NAND2_X1 U5918 ( .A1(n5354), .A2(n8466), .ZN(n5353) );
  NAND2_X1 U5919 ( .A1(n7755), .A2(n9534), .ZN(n7765) );
  OR2_X1 U5920 ( .A1(n7499), .A2(n5958), .ZN(n5960) );
  INV_X1 U5921 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6429) );
  NOR2_X1 U5922 ( .A1(n5960), .A2(n6429), .ZN(n7759) );
  NOR2_X1 U5923 ( .A1(n7793), .A2(n5352), .ZN(n9916) );
  INV_X1 U5924 ( .A(n5354), .ZN(n5352) );
  NOR2_X1 U5925 ( .A1(n7793), .A2(n7780), .ZN(n9918) );
  AND4_X1 U5926 ( .A1(n5956), .A2(n5955), .A3(n5954), .A4(n5953), .ZN(n9403)
         );
  AND2_X1 U5927 ( .A1(n9528), .A2(n9905), .ZN(n7789) );
  NOR2_X1 U5928 ( .A1(n10708), .A2(n7400), .ZN(n10709) );
  NAND2_X1 U5929 ( .A1(n7395), .A2(n7394), .ZN(n10707) );
  OR2_X1 U5930 ( .A1(n7215), .A2(n7393), .ZN(n10708) );
  NAND2_X1 U5931 ( .A1(n5539), .A2(n5538), .ZN(n7395) );
  INV_X1 U5932 ( .A(n7209), .ZN(n5539) );
  NOR2_X1 U5933 ( .A1(n7204), .A2(n7203), .ZN(n9607) );
  NAND2_X1 U5934 ( .A1(n7030), .A2(n10685), .ZN(n7215) );
  AND4_X1 U5935 ( .A1(n6937), .A2(n6936), .A3(n6935), .A4(n6934), .ZN(n10714)
         );
  NOR2_X1 U5936 ( .A1(n7048), .A2(n7164), .ZN(n7030) );
  NAND2_X1 U5937 ( .A1(n5351), .A2(n5291), .ZN(n7048) );
  NAND2_X1 U5938 ( .A1(n6670), .A2(n6674), .ZN(n7005) );
  AND4_X1 U5939 ( .A1(n5892), .A2(n5891), .A3(n5890), .A4(n5889), .ZN(n7046)
         );
  AND2_X1 U5940 ( .A1(n6209), .A2(n6212), .ZN(n6210) );
  NAND2_X1 U5941 ( .A1(n9627), .A2(n6210), .ZN(n6666) );
  AND2_X1 U5942 ( .A1(n9697), .A2(n8468), .ZN(n9942) );
  NAND2_X1 U5943 ( .A1(n5543), .A2(n7638), .ZN(n7640) );
  INV_X1 U5944 ( .A(n10878), .ZN(n10833) );
  AND2_X1 U5945 ( .A1(n6630), .A2(n7264), .ZN(n10878) );
  AND3_X1 U5946 ( .A1(n6624), .A2(n6064), .A3(n6063), .ZN(n6072) );
  XNOR2_X1 U5947 ( .A(n7945), .B(n7946), .ZN(n8437) );
  NAND2_X1 U5948 ( .A1(n5459), .A2(n7934), .ZN(n7945) );
  NAND2_X1 U5949 ( .A1(n7472), .A2(n5129), .ZN(n7659) );
  INV_X1 U5950 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n10196) );
  INV_X1 U5951 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U5952 ( .A1(n6442), .A2(n6441), .ZN(n6591) );
  NAND2_X1 U5953 ( .A1(n5443), .A2(n5441), .ZN(n6410) );
  AOI21_X1 U5954 ( .B1(n5445), .B2(n5064), .A(n5442), .ZN(n5441) );
  INV_X1 U5955 ( .A(n6404), .ZN(n5442) );
  AND2_X1 U5956 ( .A1(n6441), .A2(n6408), .ZN(n6409) );
  OAI21_X1 U5957 ( .B1(n6052), .B2(n5447), .A(n5445), .ZN(n6405) );
  NAND2_X1 U5958 ( .A1(n6128), .A2(n6127), .ZN(n6199) );
  NAND2_X1 U5959 ( .A1(n5438), .A2(n5991), .ZN(n6045) );
  AND2_X1 U5960 ( .A1(n5873), .A2(n5872), .ZN(n5875) );
  AND2_X1 U5961 ( .A1(n5802), .A2(n5822), .ZN(n7180) );
  AND2_X1 U5962 ( .A1(n5716), .A2(n5738), .ZN(n5737) );
  OR2_X1 U5963 ( .A1(n5703), .A2(SI_2_), .ZN(n5704) );
  OAI21_X1 U5964 ( .B1(n5713), .B2(n5145), .A(n5144), .ZN(n5693) );
  NAND2_X1 U5965 ( .A1(n5713), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5144) );
  AOI21_X1 U5966 ( .B1(n9320), .B2(n5580), .A(n5069), .ZN(n9374) );
  NAND2_X1 U5967 ( .A1(n5580), .A2(n9176), .ZN(n5575) );
  INV_X1 U5968 ( .A(n8670), .ZN(n5181) );
  NAND2_X1 U5969 ( .A1(n5182), .A2(n5104), .ZN(n5180) );
  AND2_X1 U5970 ( .A1(n8512), .A2(n8511), .ZN(n8574) );
  AND2_X1 U5971 ( .A1(n5178), .A2(n8507), .ZN(n8512) );
  INV_X1 U5972 ( .A(n6704), .ZN(n6791) );
  NAND2_X1 U5973 ( .A1(n8655), .A2(n8656), .ZN(n8654) );
  NOR2_X1 U5974 ( .A1(n8540), .A2(n5481), .ZN(n5478) );
  NOR2_X1 U5975 ( .A1(n5483), .A2(n5480), .ZN(n5479) );
  NAND2_X1 U5976 ( .A1(n5484), .A2(n8539), .ZN(n5483) );
  NOR3_X1 U5977 ( .A1(n8540), .A2(n5481), .A3(n8566), .ZN(n5480) );
  INV_X1 U5978 ( .A(n5485), .ZN(n5482) );
  AND2_X1 U5979 ( .A1(n7235), .A2(n7234), .ZN(n10702) );
  NAND2_X1 U5980 ( .A1(n8637), .A2(n8496), .ZN(n8591) );
  NAND2_X1 U5981 ( .A1(n8591), .A2(n8592), .ZN(n8590) );
  INV_X1 U5982 ( .A(n8698), .ZN(n7716) );
  NAND2_X1 U5983 ( .A1(n8606), .A2(n8484), .ZN(n8621) );
  XNOR2_X1 U5984 ( .A(n8519), .B(n8517), .ZN(n8631) );
  AOI22_X1 U5985 ( .A1(n6903), .A2(n6902), .B1(n6901), .B2(n6900), .ZN(n6904)
         );
  AND2_X1 U5986 ( .A1(n5495), .A2(n5080), .ZN(n7445) );
  NAND2_X1 U5987 ( .A1(n5495), .A2(n5494), .ZN(n7463) );
  NAND2_X1 U5988 ( .A1(n5512), .A2(n5510), .ZN(n8637) );
  AND2_X1 U5989 ( .A1(n8638), .A2(n5062), .ZN(n5510) );
  AND2_X1 U5990 ( .A1(n5512), .A2(n5062), .ZN(n8639) );
  AOI21_X1 U5991 ( .B1(n5490), .B2(n5493), .A(n5110), .ZN(n5488) );
  NAND2_X1 U5992 ( .A1(n5184), .A2(n5188), .ZN(n8658) );
  OR2_X1 U5993 ( .A1(n8607), .A2(n5191), .ZN(n5184) );
  NAND2_X1 U5994 ( .A1(n7099), .A2(n7098), .ZN(n7100) );
  NOR2_X1 U5995 ( .A1(n6615), .A2(n6612), .ZN(n8676) );
  OR3_X1 U5996 ( .A1(n6614), .A2(n10860), .A3(n10462), .ZN(n8693) );
  NAND2_X1 U5997 ( .A1(n8681), .A2(n8682), .ZN(n8680) );
  NAND2_X1 U5998 ( .A1(n8477), .A2(n8476), .ZN(n8681) );
  INV_X1 U5999 ( .A(n8667), .ZN(n8683) );
  OR2_X1 U6000 ( .A1(n5437), .A2(n5436), .ZN(n5343) );
  INV_X1 U6001 ( .A(n8319), .ZN(n5436) );
  INV_X1 U6002 ( .A(n8602), .ZN(n8826) );
  NAND2_X1 U6003 ( .A1(n6724), .A2(n6723), .ZN(n8705) );
  OR2_X1 U6004 ( .A1(n8217), .A2(n6911), .ZN(n6723) );
  OR2_X1 U6005 ( .A1(n6718), .A2(n6826), .ZN(n6509) );
  INV_X2 U6006 ( .A(P2_U3966), .ZN(n8708) );
  AOI21_X1 U6007 ( .B1(n10612), .B2(P2_REG2_REG_2__SCAN_IN), .A(n10608), .ZN(
        n6335) );
  AOI21_X1 U6008 ( .B1(n6268), .B2(P2_REG2_REG_4__SCAN_IN), .A(n6310), .ZN(
        n6301) );
  AOI21_X1 U6009 ( .B1(n7090), .B2(P2_REG2_REG_6__SCAN_IN), .A(n6345), .ZN(
        n6323) );
  AOI21_X1 U6010 ( .B1(n7371), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6389), .ZN(
        n6393) );
  NAND2_X1 U6011 ( .A1(n5272), .A2(n5746), .ZN(n6126) );
  INV_X1 U6012 ( .A(n5514), .ZN(n5272) );
  AOI21_X1 U6013 ( .B1(n8092), .B2(P2_REG2_REG_16__SCAN_IN), .A(n7908), .ZN(
        n7911) );
  AND2_X1 U6014 ( .A1(n5817), .A2(n5816), .ZN(n10606) );
  NAND3_X1 U6015 ( .A1(n6283), .A2(n6523), .A3(n8747), .ZN(n10607) );
  XNOR2_X1 U6016 ( .A(n8753), .B(n8745), .ZN(n9041) );
  INV_X1 U6017 ( .A(n8746), .ZN(n8745) );
  NAND2_X1 U6018 ( .A1(n5211), .A2(n5210), .ZN(n8786) );
  OR2_X1 U6019 ( .A1(n5219), .A2(n5218), .ZN(n5210) );
  AND2_X1 U6020 ( .A1(n5221), .A2(n5082), .ZN(n8805) );
  INV_X1 U6021 ( .A(n9054), .ZN(n8803) );
  NAND2_X1 U6022 ( .A1(n8201), .A2(n8200), .ZN(n9065) );
  NAND2_X1 U6023 ( .A1(n8876), .A2(n5076), .ZN(n8860) );
  NAND2_X1 U6024 ( .A1(n5225), .A2(n8303), .ZN(n8879) );
  NAND2_X1 U6025 ( .A1(n8137), .A2(n8136), .ZN(n9103) );
  OR2_X1 U6026 ( .A1(n8988), .A2(n5414), .ZN(n8971) );
  NAND2_X1 U6027 ( .A1(n6692), .A2(n6691), .ZN(n8981) );
  NAND2_X1 U6028 ( .A1(n8287), .A2(n8286), .ZN(n9011) );
  AND2_X1 U6029 ( .A1(n7582), .A2(n7822), .ZN(n7824) );
  INV_X1 U6030 ( .A(n10702), .ZN(n9034) );
  INV_X1 U6031 ( .A(n8981), .ZN(n10801) );
  OR2_X1 U6032 ( .A1(n6695), .A2(n8531), .ZN(n8793) );
  NAND2_X1 U6033 ( .A1(n7144), .A2(n7143), .ZN(n7146) );
  INV_X1 U6034 ( .A(n7142), .ZN(n8042) );
  AOI21_X1 U6035 ( .B1(n6524), .B2(n9017), .A(n5203), .ZN(n6835) );
  NAND2_X1 U6036 ( .A1(n5205), .A2(n5204), .ZN(n5203) );
  INV_X1 U6037 ( .A(n9008), .ZN(n9035) );
  AND2_X2 U6038 ( .A1(n6530), .A2(n6498), .ZN(n10873) );
  AND2_X1 U6039 ( .A1(n6489), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10583) );
  OR2_X1 U6040 ( .A1(n10462), .A2(n10461), .ZN(n10580) );
  AND2_X1 U6041 ( .A1(n5314), .A2(n5226), .ZN(n5941) );
  CLKBUF_X1 U6042 ( .A(n6279), .Z(n6280) );
  NAND2_X1 U6043 ( .A1(n5675), .A2(n5674), .ZN(n7929) );
  XNOR2_X1 U6044 ( .A(n5670), .B(n5362), .ZN(n7702) );
  NAND2_X1 U6045 ( .A1(n5682), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5670) );
  INV_X1 U6046 ( .A(n8324), .ZN(n8252) );
  INV_X1 U6047 ( .A(n8284), .ZN(n8314) );
  NAND2_X1 U6048 ( .A1(n6487), .A2(n6485), .ZN(n5280) );
  OR2_X1 U6049 ( .A1(n6487), .A2(n6485), .ZN(n6488) );
  NAND2_X1 U6050 ( .A1(n6484), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6487) );
  AND4_X1 U6051 ( .A1(n6583), .A2(n6582), .A3(n6581), .A4(n6580), .ZN(n7047)
         );
  AND4_X1 U6052 ( .A1(n5985), .A2(n5984), .A3(n5983), .A4(n5982), .ZN(n7651)
         );
  NAND2_X1 U6053 ( .A1(n7325), .A2(n7324), .ZN(n7490) );
  AND4_X2 U6054 ( .A1(n5933), .A2(n5932), .A3(n5931), .A4(n5930), .ZN(n6849)
         );
  AND2_X1 U6055 ( .A1(n9292), .A2(n5154), .ZN(n5153) );
  AND2_X1 U6056 ( .A1(n9284), .A2(n9376), .ZN(n5154) );
  NAND2_X1 U6057 ( .A1(n5166), .A2(n5582), .ZN(n7266) );
  NAND2_X1 U6058 ( .A1(n5159), .A2(n7184), .ZN(n7267) );
  NAND2_X1 U6059 ( .A1(n5166), .A2(n7179), .ZN(n5159) );
  AND3_X1 U6060 ( .A1(n8369), .A2(n8368), .A3(n8367), .ZN(n9838) );
  AND4_X1 U6061 ( .A1(n5965), .A2(n5964), .A3(n5963), .A4(n5962), .ZN(n9260)
         );
  NAND2_X1 U6062 ( .A1(n9340), .A2(n5595), .ZN(n9313) );
  NAND2_X1 U6063 ( .A1(n6566), .A2(n6565), .ZN(n6646) );
  AND4_X1 U6064 ( .A1(n7772), .A2(n7771), .A3(n7770), .A4(n7769), .ZN(n9336)
         );
  NAND2_X1 U6065 ( .A1(n5581), .A2(n9183), .ZN(n9332) );
  NAND2_X1 U6066 ( .A1(n6545), .A2(n6544), .ZN(n6548) );
  AND4_X1 U6067 ( .A1(n7281), .A2(n7280), .A3(n7279), .A4(n7278), .ZN(n10756)
         );
  INV_X1 U6068 ( .A(n5161), .ZN(n5160) );
  OAI21_X1 U6069 ( .B1(n5582), .B2(n5164), .A(n5162), .ZN(n5161) );
  INV_X1 U6070 ( .A(n10456), .ZN(n5350) );
  NAND2_X1 U6071 ( .A1(n5611), .A2(n5608), .ZN(n9355) );
  INV_X1 U6072 ( .A(n5610), .ZN(n5608) );
  NAND2_X1 U6073 ( .A1(n5125), .A2(n5612), .ZN(n5611) );
  NAND2_X1 U6074 ( .A1(n5601), .A2(n7728), .ZN(n7740) );
  NAND2_X1 U6075 ( .A1(n8387), .A2(n8386), .ZN(n9971) );
  AND4_X1 U6076 ( .A1(n7504), .A2(n7503), .A3(n7502), .A4(n7501), .ZN(n10754)
         );
  OAI21_X1 U6077 ( .B1(n7325), .B2(n5571), .A(n5568), .ZN(n7511) );
  NAND2_X1 U6078 ( .A1(n6153), .A2(n6154), .ZN(n6157) );
  AND4_X1 U6079 ( .A1(n5904), .A2(n5903), .A3(n5902), .A4(n5901), .ZN(n6671)
         );
  OR2_X1 U6080 ( .A1(n6094), .A2(n6093), .ZN(n9402) );
  NAND2_X1 U6081 ( .A1(n6021), .A2(n9897), .ZN(n9407) );
  AND4_X1 U6082 ( .A1(n6439), .A2(n6438), .A3(n6437), .A4(n6436), .ZN(n9484)
         );
  INV_X1 U6083 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5702) );
  NAND2_X1 U6084 ( .A1(n5366), .A2(n6032), .ZN(n6208) );
  NOR2_X1 U6085 ( .A1(n5100), .A2(n5367), .ZN(n5366) );
  OAI22_X1 U6086 ( .A1(n5370), .A2(n5849), .B1(n5369), .B2(n5368), .ZN(n5367)
         );
  OR2_X1 U6087 ( .A1(n6117), .A2(n10452), .ZN(n7688) );
  NOR2_X1 U6088 ( .A1(n9680), .A2(n5356), .ZN(n5355) );
  INV_X1 U6089 ( .A(n5357), .ZN(n5356) );
  INV_X1 U6090 ( .A(n5140), .ZN(n9954) );
  OAI21_X1 U6091 ( .B1(n9727), .B2(n9888), .A(n5141), .ZN(n5140) );
  AOI21_X1 U6092 ( .B1(n9950), .B2(n10822), .A(n9728), .ZN(n5141) );
  NAND2_X1 U6093 ( .A1(n8419), .A2(n8418), .ZN(n9958) );
  NAND2_X1 U6094 ( .A1(n5527), .A2(n5530), .ZN(n9737) );
  NAND2_X1 U6095 ( .A1(n8403), .A2(n5528), .ZN(n5527) );
  NAND2_X1 U6096 ( .A1(n8403), .A2(n8402), .ZN(n9749) );
  NAND2_X1 U6097 ( .A1(n5548), .A2(n5546), .ZN(n9851) );
  NAND2_X1 U6098 ( .A1(n5548), .A2(n8346), .ZN(n9849) );
  NAND2_X1 U6099 ( .A1(n9891), .A2(n8333), .ZN(n9870) );
  NAND2_X1 U6100 ( .A1(n8455), .A2(n9542), .ZN(n9886) );
  NAND2_X1 U6101 ( .A1(n7209), .A2(n5532), .ZN(n5531) );
  INV_X1 U6102 ( .A(n5536), .ZN(n5532) );
  NAND2_X1 U6103 ( .A1(n7042), .A2(n7008), .ZN(n7026) );
  INV_X1 U6104 ( .A(n9946), .ZN(n5396) );
  NOR2_X1 U6105 ( .A1(n9947), .A2(n5126), .ZN(n5142) );
  NAND2_X1 U6106 ( .A1(n6072), .A2(n6623), .ZN(n10896) );
  NAND2_X1 U6107 ( .A1(n5883), .A2(n10443), .ZN(n10449) );
  MUX2_X1 U6108 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5882), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5883) );
  NAND2_X1 U6109 ( .A1(n5635), .A2(n5637), .ZN(n7888) );
  INV_X1 U6110 ( .A(n9661), .ZN(n9596) );
  NAND2_X1 U6111 ( .A1(n7313), .A2(n7312), .ZN(n7316) );
  NAND2_X1 U6112 ( .A1(n5521), .A2(n5089), .ZN(n5519) );
  AND2_X1 U6113 ( .A1(n6987), .A2(n6600), .ZN(n8335) );
  NAND2_X1 U6114 ( .A1(n5465), .A2(n5464), .ZN(n6985) );
  NAND2_X1 U6115 ( .A1(n5465), .A2(n5466), .ZN(n6594) );
  OR2_X1 U6116 ( .A1(n6052), .A2(n6051), .ZN(n6053) );
  OR2_X1 U6117 ( .A1(n5765), .A2(n5764), .ZN(n5766) );
  NOR2_X1 U6118 ( .A1(n7619), .A2(n7618), .ZN(n10491) );
  NOR2_X1 U6119 ( .A1(n10489), .A2(n10488), .ZN(n7618) );
  NAND2_X1 U6120 ( .A1(n5581), .A2(n5580), .ZN(n5577) );
  NAND2_X1 U6121 ( .A1(n5491), .A2(n5074), .ZN(n7533) );
  NOR2_X1 U6122 ( .A1(n6838), .A2(n6837), .ZN(n6836) );
  INV_X1 U6123 ( .A(n5201), .ZN(P2_U3552) );
  AOI21_X1 U6124 ( .B1(n8708), .B2(P2_DATAO_REG_0__SCAN_IN), .A(n5202), .ZN(
        n5201) );
  NOR2_X1 U6125 ( .A1(n9062), .A2(n10813), .ZN(n8829) );
  OAI211_X1 U6126 ( .C1(n9285), .C2(n5155), .A(n5152), .B(n5149), .ZN(P1_U3218) );
  OR2_X1 U6127 ( .A1(n9292), .A2(n9410), .ZN(n5155) );
  INV_X1 U6128 ( .A(n5150), .ZN(n5149) );
  NAND2_X1 U6129 ( .A1(n9285), .A2(n5153), .ZN(n5152) );
  NAND2_X1 U6130 ( .A1(n5292), .A2(n9662), .ZN(P1_U3240) );
  NAND2_X1 U6131 ( .A1(n5294), .A2(n5293), .ZN(n5292) );
  INV_X1 U6132 ( .A(n5562), .ZN(n5561) );
  OAI21_X1 U6133 ( .B1(n9940), .B2(n10778), .A(n5563), .ZN(n5562) );
  AOI21_X1 U6134 ( .B1(n9937), .B2(n10772), .A(n9705), .ZN(n5563) );
  NAND2_X1 U6135 ( .A1(n5393), .A2(n5392), .ZN(P1_U3550) );
  NAND2_X1 U6136 ( .A1(n10894), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5392) );
  NAND2_X1 U6137 ( .A1(n10007), .A2(n10722), .ZN(n5393) );
  AND4_X2 U6138 ( .A1(n10391), .A2(n10192), .A3(n10390), .A4(n6598), .ZN(n5059) );
  INV_X1 U6139 ( .A(n8566), .ZN(n5183) );
  AND2_X1 U6140 ( .A1(n8266), .A2(n7369), .ZN(n5060) );
  INV_X1 U6141 ( .A(n5590), .ZN(n5589) );
  NAND2_X1 U6142 ( .A1(n5102), .A2(n5595), .ZN(n5590) );
  AOI21_X1 U6143 ( .B1(n8566), .B2(n8527), .A(n8530), .ZN(n5487) );
  INV_X1 U6144 ( .A(n5487), .ZN(n5481) );
  INV_X1 U6145 ( .A(n9511), .ZN(n5538) );
  NAND2_X1 U6146 ( .A1(n6568), .A2(n6569), .ZN(n7077) );
  INV_X1 U6147 ( .A(n7077), .ZN(n5291) );
  NAND2_X1 U6148 ( .A1(n8406), .A2(n8405), .ZN(n9963) );
  NOR2_X1 U6149 ( .A1(n7741), .A2(n5600), .ZN(n5061) );
  NAND2_X1 U6150 ( .A1(n8492), .A2(n8491), .ZN(n5062) );
  NAND2_X1 U6151 ( .A1(n8924), .A2(n5420), .ZN(n8909) );
  NAND2_X1 U6152 ( .A1(n8350), .A2(n8349), .ZN(n9993) );
  AND2_X1 U6153 ( .A1(n5328), .A2(n5327), .ZN(n5063) );
  AND2_X1 U6154 ( .A1(n5447), .A2(n5127), .ZN(n5064) );
  NAND2_X1 U6155 ( .A1(n8374), .A2(n8373), .ZN(n9978) );
  NAND2_X1 U6156 ( .A1(n7983), .A2(n7982), .ZN(n8791) );
  AND2_X1 U6157 ( .A1(n5213), .A2(n8312), .ZN(n5065) );
  AND2_X1 U6158 ( .A1(n8054), .A2(n5250), .ZN(n5066) );
  AND2_X1 U6159 ( .A1(n9515), .A2(n9516), .ZN(n5067) );
  AND2_X1 U6160 ( .A1(n5320), .A2(n10843), .ZN(n5068) );
  NAND2_X1 U6161 ( .A1(n5122), .A2(n5575), .ZN(n5069) );
  AND2_X1 U6162 ( .A1(n5671), .A2(n5424), .ZN(n5070) );
  NOR2_X1 U6163 ( .A1(n8582), .A2(n5511), .ZN(n5071) );
  AND2_X1 U6164 ( .A1(n9544), .A2(n5381), .ZN(n5072) );
  OR2_X1 U6165 ( .A1(n5599), .A2(n7729), .ZN(n5073) );
  INV_X2 U6166 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U6167 ( .A(n6499), .ZN(n5256) );
  NAND2_X1 U6168 ( .A1(n9871), .A2(n5345), .ZN(n5349) );
  AND2_X1 U6169 ( .A1(n5196), .A2(n7462), .ZN(n5074) );
  OR3_X1 U6170 ( .A1(n7793), .A2(n10886), .A3(n5353), .ZN(n5075) );
  OR2_X1 U6171 ( .A1(n8774), .A2(n8773), .ZN(n5076) );
  AND2_X1 U6172 ( .A1(n8241), .A2(n8239), .ZN(n5077) );
  NOR2_X1 U6173 ( .A1(n5807), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n5672) );
  NAND2_X1 U6174 ( .A1(n5643), .A2(n5388), .ZN(n5078) );
  NAND2_X1 U6175 ( .A1(n5172), .A2(n5631), .ZN(n5769) );
  NAND2_X1 U6176 ( .A1(n9054), .A2(n8787), .ZN(n8311) );
  INV_X1 U6177 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9146) );
  INV_X2 U6178 ( .A(n5908), .ZN(n6933) );
  INV_X1 U6179 ( .A(n5143), .ZN(n8318) );
  NAND2_X1 U6180 ( .A1(n8746), .A2(n8749), .ZN(n5143) );
  OR2_X1 U6181 ( .A1(n8644), .A2(n8516), .ZN(n5079) );
  NAND2_X1 U6182 ( .A1(n7437), .A2(n7438), .ZN(n5080) );
  AND2_X1 U6183 ( .A1(n5382), .A2(n9534), .ZN(n5081) );
  NAND2_X1 U6184 ( .A1(n5636), .A2(n5650), .ZN(n5635) );
  OR2_X1 U6185 ( .A1(n9059), .A2(n8807), .ZN(n5082) );
  NOR2_X1 U6186 ( .A1(n5610), .A2(n9351), .ZN(n5609) );
  NAND2_X1 U6187 ( .A1(n9190), .A2(n9189), .ZN(n5083) );
  INV_X1 U6188 ( .A(n8268), .ZN(n5250) );
  XNOR2_X1 U6189 ( .A(n5942), .B(P2_IR_REG_30__SCAN_IN), .ZN(n6383) );
  INV_X1 U6190 ( .A(n6383), .ZN(n8550) );
  INV_X2 U6191 ( .A(n6764), .ZN(n6765) );
  AND2_X1 U6192 ( .A1(n9993), .A2(n9878), .ZN(n5084) );
  AND2_X1 U6193 ( .A1(n9571), .A2(n9773), .ZN(n5085) );
  AND4_X1 U6194 ( .A1(n5343), .A2(n5268), .A3(n5435), .A4(n5267), .ZN(n5086)
         );
  OR2_X1 U6195 ( .A1(n5520), .A2(n5519), .ZN(n5087) );
  AND2_X1 U6196 ( .A1(n10640), .A2(n8252), .ZN(n5088) );
  AND3_X1 U6197 ( .A1(n5628), .A2(n5627), .A3(n5631), .ZN(n5089) );
  AND3_X1 U6198 ( .A1(n9512), .A2(n9511), .A3(n9510), .ZN(n5090) );
  AND3_X1 U6199 ( .A1(n5422), .A2(n5421), .A3(n5658), .ZN(n5091) );
  NAND2_X1 U6200 ( .A1(n5509), .A2(n5091), .ZN(n5744) );
  NAND2_X1 U6201 ( .A1(n5698), .A2(n5509), .ZN(n5735) );
  NAND2_X1 U6202 ( .A1(n7753), .A2(n7752), .ZN(n9921) );
  INV_X1 U6203 ( .A(n9948), .ZN(n9717) );
  NAND2_X1 U6204 ( .A1(n8439), .A2(n8438), .ZN(n9948) );
  NAND2_X1 U6205 ( .A1(n7994), .A2(n7993), .ZN(n9076) );
  AND2_X1 U6206 ( .A1(n8053), .A2(n8052), .ZN(n5092) );
  INV_X1 U6207 ( .A(n8824), .ZN(n8816) );
  XNOR2_X1 U6208 ( .A(n9059), .B(n8807), .ZN(n8824) );
  NOR2_X1 U6209 ( .A1(n5402), .A2(n9590), .ZN(n5093) );
  OR2_X1 U6210 ( .A1(n10843), .A2(n7903), .ZN(n5094) );
  OR2_X1 U6211 ( .A1(n9726), .A2(n5378), .ZN(n5095) );
  OR2_X1 U6212 ( .A1(n8949), .A2(n8769), .ZN(n5096) );
  AND2_X1 U6213 ( .A1(n9645), .A2(n5556), .ZN(n5097) );
  AND2_X1 U6214 ( .A1(n8255), .A2(n7581), .ZN(n5098) );
  INV_X1 U6215 ( .A(n9504), .ZN(n5402) );
  AND2_X1 U6216 ( .A1(n5081), .A2(n9544), .ZN(n5099) );
  NAND2_X1 U6217 ( .A1(n8354), .A2(n8353), .ZN(n9987) );
  AND2_X1 U6218 ( .A1(n6932), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5100) );
  AND2_X1 U6219 ( .A1(n7145), .A2(n7143), .ZN(n5101) );
  NAND2_X1 U6220 ( .A1(n8119), .A2(n8118), .ZN(n9108) );
  AND2_X1 U6221 ( .A1(n5083), .A2(n9183), .ZN(n5580) );
  INV_X1 U6222 ( .A(n6855), .ZN(n6820) );
  OR2_X1 U6223 ( .A1(n9311), .A2(n9310), .ZN(n5102) );
  INV_X1 U6224 ( .A(n9680), .ZN(n9934) );
  NAND2_X1 U6225 ( .A1(n9415), .A2(n9414), .ZN(n9680) );
  NOR2_X1 U6226 ( .A1(n8670), .A2(n8527), .ZN(n5103) );
  INV_X1 U6227 ( .A(n9503), .ZN(n5408) );
  INV_X1 U6228 ( .A(n5365), .ZN(n9818) );
  OR2_X1 U6229 ( .A1(n9833), .A2(n9473), .ZN(n5365) );
  OR2_X1 U6230 ( .A1(n5183), .A2(n8527), .ZN(n5104) );
  AND2_X1 U6231 ( .A1(n9524), .A2(n9530), .ZN(n9636) );
  INV_X1 U6232 ( .A(n5455), .ZN(n5452) );
  NOR2_X1 U6233 ( .A1(n7441), .A2(n8700), .ZN(n5105) );
  NOR2_X1 U6234 ( .A1(n9958), .A2(n9665), .ZN(n5106) );
  OR2_X1 U6235 ( .A1(n8566), .A2(n5181), .ZN(n5107) );
  INV_X1 U6236 ( .A(n5220), .ZN(n5219) );
  NAND2_X1 U6237 ( .A1(n8804), .A2(n5082), .ZN(n5220) );
  NAND2_X1 U6238 ( .A1(n5746), .A2(n5515), .ZN(n5108) );
  INV_X1 U6239 ( .A(n5535), .ZN(n5534) );
  OAI21_X1 U6240 ( .B1(n5538), .B2(n5536), .A(n5540), .ZN(n5535) );
  AND2_X1 U6241 ( .A1(n9581), .A2(n9714), .ZN(n5109) );
  XNOR2_X1 U6242 ( .A(n7981), .B(SI_29_), .ZN(n9428) );
  NOR2_X1 U6243 ( .A1(n7531), .A2(n7530), .ZN(n5110) );
  NOR2_X1 U6244 ( .A1(n8817), .A2(n9054), .ZN(n5315) );
  INV_X1 U6245 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n10200) );
  INV_X1 U6246 ( .A(n5346), .ZN(n5345) );
  NAND2_X1 U6247 ( .A1(n5348), .A2(n5347), .ZN(n5346) );
  AND2_X1 U6248 ( .A1(n9540), .A2(n5382), .ZN(n5111) );
  INV_X1 U6249 ( .A(n5547), .ZN(n5546) );
  NAND2_X1 U6250 ( .A1(n5551), .A2(n8346), .ZN(n5547) );
  AND2_X1 U6251 ( .A1(n6197), .A2(n10255), .ZN(n5112) );
  INV_X1 U6252 ( .A(n8244), .ZN(n5262) );
  OR2_X1 U6253 ( .A1(n9234), .A2(n9233), .ZN(n5113) );
  OR2_X1 U6254 ( .A1(n9739), .A2(n9738), .ZN(n5114) );
  INV_X1 U6255 ( .A(n8054), .ZN(n5248) );
  INV_X1 U6256 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n10208) );
  AND2_X1 U6257 ( .A1(n6735), .A2(n8263), .ZN(n5115) );
  AND2_X1 U6258 ( .A1(n5182), .A2(n5107), .ZN(n5116) );
  NAND2_X1 U6259 ( .A1(n5652), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5638) );
  AND2_X1 U6260 ( .A1(n8870), .A2(n5076), .ZN(n5117) );
  AND2_X1 U6261 ( .A1(n5623), .A2(n5991), .ZN(n5118) );
  AND2_X1 U6262 ( .A1(n8924), .A2(n8770), .ZN(n5119) );
  AND2_X1 U6263 ( .A1(n8304), .A2(n8303), .ZN(n5120) );
  OR2_X1 U6264 ( .A1(n5376), .A2(n9709), .ZN(n5121) );
  AND2_X1 U6265 ( .A1(n5578), .A2(n5576), .ZN(n5122) );
  AND2_X1 U6266 ( .A1(n5068), .A2(n10861), .ZN(n5123) );
  NAND2_X1 U6267 ( .A1(n9255), .A2(n9167), .ZN(n9320) );
  INV_X1 U6268 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5940) );
  AND2_X1 U6269 ( .A1(n5492), .A2(n5080), .ZN(n5124) );
  INV_X1 U6270 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5650) );
  INV_X1 U6271 ( .A(n8309), .ZN(n5217) );
  INV_X2 U6272 ( .A(n10811), .ZN(n10813) );
  NAND2_X1 U6273 ( .A1(n7381), .A2(n8055), .ZN(n9023) );
  NAND2_X1 U6274 ( .A1(n8188), .A2(n8187), .ZN(n9071) );
  INV_X1 U6275 ( .A(n9071), .ZN(n5327) );
  INV_X1 U6276 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5199) );
  NOR2_X1 U6277 ( .A1(n9372), .A2(n9377), .ZN(n5125) );
  INV_X1 U6278 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5145) );
  AND2_X1 U6279 ( .A1(n9948), .A2(n10877), .ZN(n5126) );
  AND2_X1 U6280 ( .A1(n6404), .A2(n6203), .ZN(n5127) );
  INV_X1 U6281 ( .A(n9542), .ZN(n5381) );
  NOR2_X1 U6282 ( .A1(n5269), .A2(n5514), .ZN(n6451) );
  NAND3_X1 U6283 ( .A1(n5730), .A2(n5629), .A3(n5630), .ZN(n5767) );
  INV_X1 U6284 ( .A(n5767), .ZN(n5172) );
  OR2_X1 U6285 ( .A1(n9003), .A2(n5325), .ZN(n5128) );
  INV_X1 U6286 ( .A(n8807), .ZN(n8779) );
  AND2_X1 U6287 ( .A1(n8226), .A2(n8225), .ZN(n8807) );
  AND2_X1 U6288 ( .A1(n5472), .A2(n7471), .ZN(n5129) );
  NAND2_X1 U6289 ( .A1(n8911), .A2(n5330), .ZN(n5331) );
  INV_X1 U6290 ( .A(n5326), .ZN(n8996) );
  NOR2_X1 U6291 ( .A1(n9003), .A2(n9119), .ZN(n5326) );
  INV_X1 U6292 ( .A(n5467), .ZN(n5466) );
  NOR2_X1 U6293 ( .A1(n6589), .A2(SI_16_), .ZN(n5467) );
  INV_X1 U6294 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6485) );
  OR2_X1 U6295 ( .A1(n7793), .A2(n5353), .ZN(n5130) );
  NOR2_X1 U6296 ( .A1(n8988), .A2(n5416), .ZN(n5131) );
  AND2_X1 U6297 ( .A1(n7871), .A2(n8082), .ZN(n5132) );
  INV_X1 U6298 ( .A(n9158), .ZN(n5599) );
  OAI21_X1 U6299 ( .B1(n6805), .B2(n6673), .A(n9453), .ZN(n7001) );
  NAND2_X1 U6300 ( .A1(n5531), .A2(n5534), .ZN(n7633) );
  NOR2_X1 U6301 ( .A1(n9607), .A2(n7205), .ZN(n5133) );
  NAND2_X1 U6302 ( .A1(n8364), .A2(n8363), .ZN(n9981) );
  INV_X1 U6303 ( .A(n9981), .ZN(n5347) );
  NAND2_X1 U6304 ( .A1(n5291), .A2(n9673), .ZN(n9459) );
  INV_X1 U6305 ( .A(n9459), .ZN(n5386) );
  NAND2_X1 U6306 ( .A1(n10793), .A2(n5068), .ZN(n5321) );
  AND3_X1 U6307 ( .A1(n5333), .A2(n5170), .A3(n5172), .ZN(n5639) );
  AND2_X1 U6308 ( .A1(n5624), .A2(n7369), .ZN(n5134) );
  AND2_X1 U6309 ( .A1(n10787), .A2(n7581), .ZN(n5135) );
  AND2_X1 U6310 ( .A1(n7382), .A2(n8058), .ZN(n5136) );
  INV_X1 U6311 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5363) );
  NAND2_X1 U6312 ( .A1(n8248), .A2(n8284), .ZN(n6755) );
  NAND2_X1 U6313 ( .A1(n9596), .A2(n9760), .ZN(n9590) );
  INV_X1 U6314 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5362) );
  INV_X1 U6315 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5361) );
  OR2_X1 U6316 ( .A1(n6810), .A2(n6860), .ZN(n7043) );
  INV_X1 U6317 ( .A(n7043), .ZN(n5351) );
  XNOR2_X1 U6318 ( .A(n6018), .B(n6017), .ZN(n7264) );
  INV_X1 U6319 ( .A(n5888), .ZN(n8474) );
  INV_X1 U6320 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5200) );
  INV_X1 U6321 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5368) );
  AOI21_X1 U6322 ( .B1(n10861), .B2(n8761), .A(n8760), .ZN(n9002) );
  NAND2_X1 U6323 ( .A1(n10789), .A2(n10788), .ZN(n10787) );
  NAND2_X1 U6324 ( .A1(n8942), .A2(n8298), .ZN(n8946) );
  INV_X1 U6325 ( .A(n9639), .ZN(n5382) );
  NAND2_X1 U6326 ( .A1(n6788), .A2(n5115), .ZN(n5206) );
  NAND2_X1 U6327 ( .A1(n7007), .A2(n7006), .ZN(n7042) );
  NAND2_X1 U6328 ( .A1(n7928), .A2(n7927), .ZN(n7931) );
  NAND2_X1 U6329 ( .A1(n7957), .A2(n7956), .ZN(n7960) );
  AOI21_X1 U6330 ( .B1(n5261), .B2(n5262), .A(n8248), .ZN(n5260) );
  OAI21_X1 U6331 ( .B1(n7262), .B2(n7261), .A(n7260), .ZN(n7309) );
  NAND2_X1 U6332 ( .A1(n9159), .A2(n9158), .ZN(n9166) );
  NAND2_X1 U6333 ( .A1(n5577), .A2(n5578), .ZN(n9196) );
  NAND2_X1 U6334 ( .A1(n9248), .A2(n9247), .ZN(n9285) );
  NAND2_X1 U6335 ( .A1(n5588), .A2(n5584), .ZN(n9386) );
  NAND2_X1 U6336 ( .A1(n5604), .A2(n5602), .ZN(n9303) );
  NAND2_X1 U6337 ( .A1(n9362), .A2(n9363), .ZN(n9361) );
  NAND2_X1 U6338 ( .A1(n7370), .A2(n8211), .ZN(n5193) );
  INV_X1 U6339 ( .A(n7416), .ZN(n5146) );
  NAND2_X1 U6340 ( .A1(n5427), .A2(n5426), .ZN(n7416) );
  NAND2_X1 U6341 ( .A1(n9607), .A2(n5404), .ZN(n5403) );
  NAND2_X1 U6342 ( .A1(n5114), .A2(n9498), .ZN(n9725) );
  AOI21_X1 U6343 ( .B1(n7755), .B2(n5099), .A(n5380), .ZN(n9877) );
  NAND2_X1 U6344 ( .A1(n9459), .A2(n5384), .ZN(n5282) );
  NAND2_X1 U6345 ( .A1(n7338), .A2(n7337), .ZN(n7368) );
  NAND2_X1 U6346 ( .A1(n5543), .A2(n5541), .ZN(n7779) );
  NAND2_X1 U6347 ( .A1(n9803), .A2(n9806), .ZN(n5557) );
  OAI21_X1 U6348 ( .B1(n7787), .B2(n7789), .A(n7781), .ZN(n9914) );
  NAND2_X1 U6349 ( .A1(n5522), .A2(n5525), .ZN(n9722) );
  NAND2_X1 U6350 ( .A1(n5396), .A2(n5394), .ZN(n10007) );
  NAND2_X1 U6351 ( .A1(n5173), .A2(n5793), .ZN(n5798) );
  NAND2_X1 U6352 ( .A1(n5783), .A2(n5782), .ZN(n5792) );
  NAND2_X1 U6353 ( .A1(n7965), .A2(n7964), .ZN(n7969) );
  NAND2_X1 U6354 ( .A1(n5988), .A2(n5987), .ZN(n5438) );
  NAND2_X1 U6355 ( .A1(n7950), .A2(n7949), .ZN(n7957) );
  NAND2_X1 U6356 ( .A1(n7085), .A2(n7084), .ZN(n7262) );
  INV_X1 U6357 ( .A(n8250), .ZN(n8285) );
  NAND2_X1 U6358 ( .A1(n7887), .A2(n5473), .ZN(n7928) );
  INV_X1 U6359 ( .A(n8321), .ZN(n5268) );
  NOR2_X2 U6360 ( .A1(n9224), .A2(n9223), .ZN(n9267) );
  NAND2_X1 U6361 ( .A1(n5148), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n5637) );
  NAND2_X1 U6362 ( .A1(n7175), .A2(n5157), .ZN(n5156) );
  NAND2_X1 U6363 ( .A1(n5156), .A2(n5160), .ZN(n7320) );
  AND3_X1 U6364 ( .A1(n5059), .A2(n5521), .A3(n5633), .ZN(n5170) );
  NAND4_X1 U6365 ( .A1(n5333), .A2(n5172), .A3(n5059), .A4(n5171), .ZN(n5652)
         );
  AND4_X2 U6366 ( .A1(n10396), .A2(n10397), .A3(n10174), .A4(n5626), .ZN(n5521) );
  NAND2_X1 U6367 ( .A1(n5792), .A2(n5791), .ZN(n5173) );
  NAND2_X1 U6368 ( .A1(n5765), .A2(n5764), .ZN(n5783) );
  NAND2_X1 U6369 ( .A1(n5488), .A2(n5489), .ZN(n7710) );
  NAND2_X1 U6370 ( .A1(n8671), .A2(n5116), .ZN(n5179) );
  OAI211_X1 U6371 ( .C1(n8671), .C2(n5180), .A(n8683), .B(n5179), .ZN(n8571)
         );
  NAND2_X1 U6372 ( .A1(n8671), .A2(n8670), .ZN(n8669) );
  NAND2_X1 U6373 ( .A1(n8607), .A2(n5188), .ZN(n5187) );
  NAND2_X2 U6374 ( .A1(n5193), .A2(n7372), .ZN(n7441) );
  AND2_X1 U6375 ( .A1(n7444), .A2(n5080), .ZN(n5494) );
  NAND2_X1 U6376 ( .A1(n5124), .A2(n7444), .ZN(n5196) );
  OAI211_X1 U6377 ( .C1(n5456), .C2(n5199), .A(n5198), .B(n5197), .ZN(n5714)
         );
  NAND3_X1 U6378 ( .A1(n5456), .A2(n5455), .A3(P2_DATAO_REG_3__SCAN_IN), .ZN(
        n5197) );
  NAND2_X1 U6379 ( .A1(n6514), .A2(n10639), .ZN(n8023) );
  NOR2_X1 U6380 ( .A1(n8708), .A2(n6780), .ZN(n5202) );
  NAND2_X1 U6381 ( .A1(n9012), .A2(n6514), .ZN(n5204) );
  NAND2_X1 U6382 ( .A1(n6704), .A2(n9014), .ZN(n5205) );
  NAND2_X1 U6383 ( .A1(n8848), .A2(n5208), .ZN(n5207) );
  AND2_X1 U6384 ( .A1(n5216), .A2(n8309), .ZN(n8825) );
  NAND2_X1 U6385 ( .A1(n9023), .A2(n5222), .ZN(n5224) );
  NAND2_X1 U6386 ( .A1(n5223), .A2(n8070), .ZN(n7811) );
  NAND2_X1 U6387 ( .A1(n5339), .A2(n5224), .ZN(n5223) );
  NAND2_X1 U6388 ( .A1(n5225), .A2(n5120), .ZN(n8867) );
  NAND2_X1 U6389 ( .A1(n5314), .A2(n5667), .ZN(n5807) );
  AND2_X1 U6390 ( .A1(n5070), .A2(n5667), .ZN(n5226) );
  NOR2_X2 U6391 ( .A1(n5943), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n5945) );
  NAND3_X1 U6392 ( .A1(n5232), .A2(n5077), .A3(n5229), .ZN(n5228) );
  NAND2_X1 U6393 ( .A1(n5233), .A2(n5255), .ZN(n8198) );
  NAND2_X1 U6394 ( .A1(n5234), .A2(n8833), .ZN(n5233) );
  NAND2_X1 U6395 ( .A1(n8196), .A2(n8866), .ZN(n5234) );
  NAND2_X1 U6396 ( .A1(n8184), .A2(n8185), .ZN(n8196) );
  NAND2_X1 U6397 ( .A1(n5249), .A2(n9031), .ZN(n8061) );
  NAND2_X1 U6398 ( .A1(n8240), .A2(n5264), .ZN(n5263) );
  NAND2_X1 U6399 ( .A1(n8240), .A2(n5257), .ZN(n5258) );
  NAND2_X1 U6400 ( .A1(n5271), .A2(n5746), .ZN(n5269) );
  NAND2_X1 U6401 ( .A1(n5746), .A2(n5273), .ZN(n5270) );
  OAI21_X1 U6402 ( .B1(n8075), .B2(n5276), .A(n5274), .ZN(n8105) );
  NOR2_X1 U6403 ( .A1(n8074), .A2(n8255), .ZN(n5279) );
  NAND2_X2 U6404 ( .A1(n6488), .A2(n5280), .ZN(n6499) );
  NAND3_X1 U6405 ( .A1(n5306), .A2(n5305), .A3(n9594), .ZN(n5304) );
  NAND3_X1 U6406 ( .A1(n9585), .A2(n9624), .A3(n9558), .ZN(n5305) );
  OAI211_X2 U6407 ( .C1(n6702), .C2(n6511), .A(n5311), .B(n5310), .ZN(n6759)
         );
  OR2_X1 U6408 ( .A1(n6729), .A2(n6512), .ZN(n5310) );
  NAND4_X1 U6409 ( .A1(n10639), .A2(n6832), .A3(n10656), .A4(n6795), .ZN(n6797) );
  NAND2_X1 U6410 ( .A1(n10793), .A2(n5123), .ZN(n9005) );
  INV_X1 U6411 ( .A(n5321), .ZN(n8744) );
  INV_X1 U6412 ( .A(n5331), .ZN(n8888) );
  NAND2_X1 U6413 ( .A1(n5318), .A2(n6704), .ZN(n8027) );
  NAND2_X1 U6414 ( .A1(n8917), .A2(n8301), .ZN(n5332) );
  NAND4_X1 U6415 ( .A1(n5627), .A2(n5628), .A3(n5631), .A4(n6019), .ZN(n5334)
         );
  OAI21_X1 U6416 ( .B1(n7871), .B2(n5337), .A(n5335), .ZN(n8290) );
  INV_X1 U6417 ( .A(n5349), .ZN(n9809) );
  MUX2_X1 U6418 ( .A(n6166), .B(n5350), .S(n6537), .Z(n6855) );
  AND2_X1 U6419 ( .A1(n9729), .A2(n5357), .ZN(n9696) );
  NAND2_X1 U6420 ( .A1(n9729), .A2(n5355), .ZN(n9675) );
  NAND2_X1 U6421 ( .A1(n9729), .A2(n5359), .ZN(n9697) );
  NAND2_X1 U6422 ( .A1(n9450), .A2(n6215), .ZN(n6672) );
  NAND2_X1 U6423 ( .A1(n8474), .A2(n10449), .ZN(n5369) );
  NAND2_X1 U6424 ( .A1(n9751), .A2(n5373), .ZN(n5372) );
  AOI21_X1 U6425 ( .B1(n9751), .B2(n9750), .A(n9574), .ZN(n9739) );
  NAND2_X1 U6426 ( .A1(n5371), .A2(n5121), .ZN(n9710) );
  INV_X1 U6427 ( .A(n9574), .ZN(n5379) );
  NAND2_X1 U6428 ( .A1(n7000), .A2(n9456), .ZN(n5384) );
  OAI21_X1 U6429 ( .B1(n7001), .B2(n7000), .A(n9456), .ZN(n7044) );
  AND2_X1 U6430 ( .A1(n5614), .A2(n5390), .ZN(n5388) );
  NAND2_X1 U6431 ( .A1(n5643), .A2(n5614), .ZN(n5656) );
  OR2_X1 U6432 ( .A1(n9607), .A2(n5407), .ZN(n5406) );
  NAND2_X1 U6433 ( .A1(n7788), .A2(n7789), .ZN(n9906) );
  NAND2_X1 U6434 ( .A1(n9856), .A2(n9855), .ZN(n9854) );
  NAND2_X1 U6435 ( .A1(n7398), .A2(n5067), .ZN(n7648) );
  NAND2_X1 U6436 ( .A1(n5434), .A2(n8313), .ZN(n8315) );
  NAND2_X1 U6437 ( .A1(n8290), .A2(n8289), .ZN(n8992) );
  NAND2_X1 U6438 ( .A1(n8961), .A2(n8297), .ZN(n8942) );
  NAND2_X1 U6439 ( .A1(n5437), .A2(n8320), .ZN(n5435) );
  NAND2_X1 U6440 ( .A1(n9877), .A2(n9876), .ZN(n9875) );
  XNOR2_X1 U6441 ( .A(n9710), .B(n9714), .ZN(n9711) );
  NAND2_X1 U6442 ( .A1(n5560), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5655) );
  NAND2_X2 U6443 ( .A1(n8850), .A2(n8849), .ZN(n8848) );
  NAND2_X1 U6444 ( .A1(n8989), .A2(n5413), .ZN(n5409) );
  AND2_X1 U6445 ( .A1(n9119), .A2(n9015), .ZN(n5416) );
  NAND2_X1 U6446 ( .A1(n7144), .A2(n5101), .ZN(n7338) );
  INV_X1 U6447 ( .A(n5671), .ZN(n5423) );
  NAND2_X1 U6448 ( .A1(n9032), .A2(n5060), .ZN(n5427) );
  NAND3_X1 U6449 ( .A1(n5428), .A2(n6888), .A3(n6521), .ZN(n8028) );
  NAND2_X1 U6450 ( .A1(n5428), .A2(n6521), .ZN(n6704) );
  NAND2_X1 U6451 ( .A1(n5431), .A2(n5711), .ZN(n5718) );
  NAND2_X1 U6452 ( .A1(n5709), .A2(n5710), .ZN(n5431) );
  INV_X1 U6453 ( .A(n5711), .ZN(n5433) );
  INV_X1 U6454 ( .A(n8315), .ZN(n8317) );
  NAND2_X1 U6455 ( .A1(n5438), .A2(n5118), .ZN(n6047) );
  NAND2_X1 U6456 ( .A1(n5819), .A2(n5439), .ZN(n5871) );
  NAND2_X1 U6457 ( .A1(n6052), .A2(n5444), .ZN(n5443) );
  NAND3_X1 U6458 ( .A1(n5456), .A2(n5455), .A3(n6023), .ZN(n5450) );
  NAND2_X1 U6459 ( .A1(n5459), .A2(n5457), .ZN(n7948) );
  INV_X1 U6460 ( .A(n7946), .ZN(n5460) );
  NAND2_X1 U6461 ( .A1(n7695), .A2(n5475), .ZN(n7887) );
  NAND2_X1 U6462 ( .A1(n7695), .A2(n7694), .ZN(n7698) );
  NAND2_X1 U6463 ( .A1(n8669), .A2(n5478), .ZN(n5477) );
  OAI211_X1 U6464 ( .C1(n8669), .C2(n5482), .A(n5479), .B(n5477), .ZN(n8544)
         );
  NAND2_X1 U6465 ( .A1(n7440), .A2(n5490), .ZN(n5489) );
  NAND2_X1 U6466 ( .A1(n7898), .A2(n5497), .ZN(n5496) );
  INV_X1 U6467 ( .A(n5504), .ZN(n6777) );
  NAND2_X1 U6468 ( .A1(n6975), .A2(n5506), .ZN(n5505) );
  NAND2_X1 U6469 ( .A1(n8655), .A2(n5071), .ZN(n5512) );
  INV_X1 U6470 ( .A(n5512), .ZN(n8581) );
  NAND2_X1 U6471 ( .A1(n5746), .A2(n5517), .ZN(n5820) );
  NAND2_X1 U6472 ( .A1(n9448), .A2(n9446), .ZN(n9627) );
  NAND2_X1 U6473 ( .A1(n8403), .A2(n5523), .ZN(n5522) );
  OAI21_X1 U6474 ( .B1(n7209), .B2(n5535), .A(n5533), .ZN(n7636) );
  NAND2_X1 U6475 ( .A1(n7042), .A2(n5552), .ZN(n7024) );
  NAND2_X1 U6476 ( .A1(n8436), .A2(n5554), .ZN(n5553) );
  NAND2_X1 U6477 ( .A1(n5553), .A2(n5556), .ZN(n8453) );
  NAND2_X2 U6478 ( .A1(n6537), .A2(n7966), .ZN(n6149) );
  OAI21_X1 U6479 ( .B1(n9935), .B2(n9885), .A(n5561), .ZN(P1_U3355) );
  INV_X1 U6480 ( .A(n5565), .ZN(n7516) );
  NAND2_X1 U6481 ( .A1(n5573), .A2(n7324), .ZN(n5572) );
  INV_X1 U6482 ( .A(n7489), .ZN(n5573) );
  NAND2_X1 U6483 ( .A1(n9178), .A2(n9177), .ZN(n5581) );
  INV_X1 U6484 ( .A(n9267), .ZN(n5592) );
  NOR2_X1 U6485 ( .A1(n9267), .A2(n5593), .ZN(n9341) );
  INV_X1 U6486 ( .A(n5594), .ZN(n5593) );
  NAND2_X1 U6487 ( .A1(n5596), .A2(n5597), .ZN(n9254) );
  NAND2_X1 U6488 ( .A1(n5601), .A2(n5061), .ZN(n9159) );
  NAND2_X1 U6489 ( .A1(n9372), .A2(n5609), .ZN(n5604) );
  OR2_X1 U6490 ( .A1(n8820), .A2(n8217), .ZN(n8226) );
  OR2_X1 U6491 ( .A1(n8840), .A2(n8217), .ZN(n8209) );
  INV_X1 U6492 ( .A(n6516), .ZN(n8217) );
  OR2_X1 U6493 ( .A1(n6707), .A2(n6529), .ZN(n6510) );
  AND2_X1 U6494 ( .A1(n6722), .A2(n6721), .ZN(n6724) );
  AND2_X1 U6495 ( .A1(n6516), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6517) );
  CLKBUF_X1 U6496 ( .A(n7867), .Z(n10847) );
  INV_X1 U6497 ( .A(n8465), .ZN(n9944) );
  OAI21_X1 U6498 ( .B1(n9945), .B2(n10718), .A(n8464), .ZN(n8465) );
  NAND2_X1 U6499 ( .A1(n8631), .A2(n8630), .ZN(n8629) );
  CLKBUF_X1 U6500 ( .A(n6513), .Z(n8547) );
  AOI21_X1 U6501 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n6719), .A(n5618), .ZN(
        n6722) );
  BUF_X4 U6502 ( .A(n6719), .Z(n8192) );
  NAND2_X1 U6503 ( .A1(n9702), .A2(n5622), .ZN(n9704) );
  XNOR2_X1 U6504 ( .A(n6832), .B(n6764), .ZN(n6760) );
  OR2_X1 U6505 ( .A1(n9935), .A2(n10831), .ZN(n9939) );
  AND2_X1 U6506 ( .A1(n6207), .A2(n6820), .ZN(n6845) );
  OAI22_X2 U6507 ( .A1(n8551), .A2(n8552), .B1(n7231), .B2(n7230), .ZN(n7440)
         );
  NOR2_X1 U6508 ( .A1(n6718), .A2(n6266), .ZN(n5618) );
  NAND2_X1 U6509 ( .A1(n10811), .A2(n10809), .ZN(n9022) );
  OR2_X1 U6510 ( .A1(n9966), .A2(n9799), .ZN(n5619) );
  INV_X1 U6511 ( .A(n8878), .ZN(n8304) );
  AND2_X1 U6512 ( .A1(n6057), .A2(n6056), .ZN(n5620) );
  NAND2_X1 U6513 ( .A1(n6072), .A2(n10442), .ZN(n10894) );
  INV_X2 U6514 ( .A(n10894), .ZN(n10722) );
  NAND2_X2 U6515 ( .A1(n7015), .A2(n9897), .ZN(n10783) );
  NAND3_X1 U6516 ( .A1(n5651), .A2(n5650), .A3(n10204), .ZN(n5621) );
  NAND2_X1 U6517 ( .A1(n6761), .A2(n6760), .ZN(n6762) );
  AND2_X1 U6518 ( .A1(n6046), .A2(n5995), .ZN(n5623) );
  AND3_X1 U6519 ( .A1(n8195), .A2(n8194), .A3(n8193), .ZN(n8672) );
  INV_X1 U6520 ( .A(n8965), .ZN(n8764) );
  INV_X4 U6521 ( .A(n5712), .ZN(n7958) );
  OR2_X1 U6522 ( .A1(n9054), .A2(n8827), .ZN(n5625) );
  INV_X1 U6523 ( .A(n9607), .ZN(n9610) );
  INV_X1 U6524 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5663) );
  INV_X1 U6525 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5632) );
  NAND2_X1 U6526 ( .A1(n5046), .A2(n9239), .ZN(n6152) );
  INV_X1 U6527 ( .A(n8167), .ZN(n6379) );
  INV_X1 U6528 ( .A(n8138), .ZN(n6377) );
  NAND2_X1 U6529 ( .A1(n5327), .A2(n8672), .ZN(n8776) );
  NAND2_X1 U6530 ( .A1(n8261), .A2(n8024), .ZN(n6879) );
  INV_X1 U6531 ( .A(n8266), .ZN(n7383) );
  NAND2_X1 U6532 ( .A1(n5806), .A2(n5363), .ZN(n5669) );
  INV_X1 U6533 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6056) );
  INV_X1 U6534 ( .A(n9651), .ZN(n9601) );
  NAND2_X1 U6535 ( .A1(n7767), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8339) );
  OR2_X1 U6536 ( .A1(n8375), .A2(n9304), .ZN(n8377) );
  NOR2_X1 U6537 ( .A1(n7277), .A2(n5980), .ZN(n7498) );
  INV_X1 U6538 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5884) );
  INV_X1 U6539 ( .A(n8095), .ZN(n6375) );
  INV_X1 U6540 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n10319) );
  INV_X1 U6541 ( .A(n8171), .ZN(n8218) );
  INV_X1 U6542 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10080) );
  OR2_X1 U6543 ( .A1(n9065), .A2(n8826), .ZN(n8778) );
  INV_X1 U6544 ( .A(n9114), .ZN(n8765) );
  INV_X1 U6545 ( .A(n8264), .ZN(n7145) );
  INV_X1 U6546 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5810) );
  INV_X1 U6547 ( .A(n6549), .ZN(n6546) );
  OR2_X1 U6548 ( .A1(n8365), .A2(n9356), .ZN(n8375) );
  NOR2_X1 U6549 ( .A1(n8377), .A2(n9367), .ZN(n8393) );
  AND2_X1 U6550 ( .A1(n9462), .A2(n9503), .ZN(n9511) );
  OR2_X1 U6551 ( .A1(n9513), .A2(n5402), .ZN(n10712) );
  AND2_X1 U6552 ( .A1(n9596), .A2(n9653), .ZN(n6630) );
  OR2_X1 U6553 ( .A1(n7960), .A2(n7959), .ZN(n7961) );
  INV_X1 U6554 ( .A(SI_26_), .ZN(n10027) );
  OR2_X1 U6555 ( .A1(n6413), .A2(n6412), .ZN(n6454) );
  INV_X1 U6556 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10291) );
  INV_X1 U6557 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10293) );
  INV_X1 U6558 ( .A(n8964), .ZN(n8769) );
  INV_X1 U6559 ( .A(n8508), .ZN(n8514) );
  NAND2_X1 U6560 ( .A1(n6767), .A2(n6766), .ZN(n6768) );
  NAND2_X1 U6561 ( .A1(n8676), .A2(n9012), .ZN(n8688) );
  INV_X1 U6562 ( .A(n8192), .ZN(n8223) );
  INV_X1 U6563 ( .A(n9108), .ZN(n8960) );
  AND2_X1 U6564 ( .A1(n8070), .A2(n8067), .ZN(n7419) );
  OR2_X1 U6565 ( .A1(n7236), .A2(n10293), .ZN(n7244) );
  AND2_X1 U6566 ( .A1(n8324), .A2(n8284), .ZN(n6522) );
  INV_X1 U6567 ( .A(n10860), .ZN(n9124) );
  INV_X1 U6568 ( .A(n8696), .ZN(n7903) );
  INV_X2 U6569 ( .A(n6651), .ZN(n9208) );
  AND3_X1 U6570 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6578) );
  AND2_X1 U6571 ( .A1(n6157), .A2(n6239), .ZN(n6158) );
  OR2_X1 U6572 ( .A1(n6094), .A2(n6030), .ZN(n9388) );
  INV_X1 U6573 ( .A(n6091), .ZN(n9598) );
  AND2_X1 U6574 ( .A1(n8393), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8407) );
  AOI21_X1 U6575 ( .B1(n8463), .B2(n10758), .A(n8462), .ZN(n8464) );
  INV_X1 U6576 ( .A(n9799), .ZN(n9752) );
  INV_X1 U6577 ( .A(n9966), .ZN(n9771) );
  OR2_X1 U6578 ( .A1(n10441), .A2(n6061), .ZN(n9897) );
  AND2_X1 U6579 ( .A1(n6630), .A2(n6092), .ZN(n10877) );
  INV_X1 U6580 ( .A(n10758), .ZN(n9888) );
  AND2_X1 U6581 ( .A1(n5752), .A2(n5751), .ZN(n10018) );
  XNOR2_X1 U6582 ( .A(n6589), .B(SI_16_), .ZN(n6590) );
  AND2_X1 U6583 ( .A1(n6127), .A2(n6050), .ZN(n6051) );
  AND2_X1 U6584 ( .A1(n5818), .A2(n5796), .ZN(n5797) );
  INV_X1 U6585 ( .A(n7702), .ZN(n6479) );
  INV_X1 U6586 ( .A(n8555), .ZN(n8685) );
  AND2_X1 U6587 ( .A1(n6772), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8690) );
  NAND2_X1 U6588 ( .A1(n6719), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6508) );
  INV_X1 U6589 ( .A(n10586), .ZN(n10615) );
  INV_X1 U6590 ( .A(n10607), .ZN(n10584) );
  INV_X1 U6591 ( .A(n8781), .ZN(n8804) );
  INV_X1 U6592 ( .A(n8768), .ZN(n8962) );
  INV_X1 U6593 ( .A(n8763), .ZN(n9010) );
  INV_X1 U6594 ( .A(n9022), .ZN(n9033) );
  AND2_X1 U6595 ( .A1(n10579), .A2(n6497), .ZN(n6687) );
  INV_X1 U6596 ( .A(n10866), .ZN(n10841) );
  INV_X1 U6597 ( .A(n7929), .ZN(n6496) );
  AND2_X1 U6598 ( .A1(n5748), .A2(n5747), .ZN(n6948) );
  NAND2_X1 U6599 ( .A1(n6243), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9401) );
  INV_X1 U6600 ( .A(n9410), .ZN(n9376) );
  INV_X1 U6601 ( .A(n9401), .ZN(n9347) );
  INV_X1 U6602 ( .A(n7264), .ZN(n9657) );
  AND4_X1 U6603 ( .A1(n8452), .A2(n8451), .A3(n8450), .A4(n8449), .ZN(n9712)
         );
  AND2_X1 U6604 ( .A1(n8383), .A2(n8382), .ZN(n9820) );
  INV_X1 U6605 ( .A(n7688), .ZN(n10633) );
  INV_X1 U6606 ( .A(n10566), .ZN(n10628) );
  INV_X1 U6607 ( .A(n10626), .ZN(n10550) );
  AND2_X1 U6608 ( .A1(n5863), .A2(n10452), .ZN(n10566) );
  AND2_X1 U6609 ( .A1(n9791), .A2(n9570), .ZN(n9788) );
  AND2_X1 U6610 ( .A1(n9548), .A2(n9549), .ZN(n9876) );
  NAND2_X1 U6611 ( .A1(n6067), .A2(n6066), .ZN(n10758) );
  INV_X1 U6612 ( .A(n10877), .ZN(n10888) );
  OR2_X1 U6613 ( .A1(n9590), .A2(n9657), .ZN(n10817) );
  AND2_X1 U6614 ( .A1(n10718), .A2(n10817), .ZN(n10831) );
  INV_X1 U6615 ( .A(n10718), .ZN(n10822) );
  INV_X1 U6616 ( .A(n10442), .ZN(n6623) );
  INV_X1 U6617 ( .A(n10441), .ZN(n10020) );
  INV_X1 U6618 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6019) );
  AND2_X1 U6619 ( .A1(n6204), .A2(n6133), .ZN(n7721) );
  NOR2_X1 U6620 ( .A1(n10476), .A2(n7598), .ZN(n7599) );
  NOR2_X1 U6621 ( .A1(n10487), .A2(n10486), .ZN(n7615) );
  INV_X1 U6622 ( .A(n10583), .ZN(n5683) );
  INV_X1 U6623 ( .A(n7892), .ZN(n10861) );
  INV_X1 U6624 ( .A(n9076), .ZN(n8866) );
  NAND2_X1 U6625 ( .A1(n10860), .A2(n6618), .ZN(n8667) );
  INV_X1 U6626 ( .A(n8672), .ZN(n8872) );
  INV_X1 U6627 ( .A(n10613), .ZN(n10585) );
  OR2_X1 U6628 ( .A1(n10813), .A2(n6872), .ZN(n8987) );
  INV_X1 U6629 ( .A(n10870), .ZN(n10868) );
  AND2_X2 U6630 ( .A1(n6530), .A2(n6687), .ZN(n10870) );
  INV_X1 U6631 ( .A(n10873), .ZN(n10871) );
  NOR2_X1 U6632 ( .A1(n6492), .A2(n6496), .ZN(n10464) );
  INV_X1 U6633 ( .A(n9921), .ZN(n10853) );
  INV_X1 U6634 ( .A(n9407), .ZN(n9384) );
  OR2_X1 U6635 ( .A1(n6094), .A2(n6033), .ZN(n9410) );
  OAI21_X1 U6636 ( .B1(n9768), .B2(n8400), .A(n8399), .ZN(n9799) );
  OR2_X1 U6637 ( .A1(n6039), .A2(n5755), .ZN(n9674) );
  OR2_X1 U6638 ( .A1(P1_U3083), .A2(n5861), .ZN(n10626) );
  INV_X1 U6639 ( .A(n9926), .ZN(n9885) );
  AND3_X1 U6640 ( .A1(n10882), .A2(n10881), .A3(n10880), .ZN(n10885) );
  AND2_X1 U6641 ( .A1(n10775), .A2(n10767), .ZN(n10769) );
  NAND2_X1 U6642 ( .A1(n10020), .A2(n10019), .ZN(n10460) );
  XNOR2_X1 U6643 ( .A(n5638), .B(n10204), .ZN(n7701) );
  NOR2_X1 U6644 ( .A1(n7616), .A2(n7615), .ZN(n10489) );
  NOR2_X1 U6645 ( .A1(n6490), .A2(n5683), .ZN(P2_U3966) );
  INV_X2 U6646 ( .A(n9674), .ZN(P1_U4006) );
  OR3_X4 U6647 ( .A1(n5750), .A2(n7888), .A3(n7701), .ZN(n6039) );
  INV_X1 U6648 ( .A(n5639), .ZN(n5640) );
  NAND2_X1 U6649 ( .A1(n5640), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5641) );
  MUX2_X1 U6650 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5641), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n5642) );
  NAND2_X1 U6651 ( .A1(n5642), .A2(n5652), .ZN(n5860) );
  NAND2_X1 U6652 ( .A1(n5860), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5755) );
  NAND2_X1 U6653 ( .A1(n6018), .A2(n6017), .ZN(n5644) );
  NAND2_X1 U6654 ( .A1(n5644), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5646) );
  NAND2_X1 U6655 ( .A1(n5646), .A2(n10196), .ZN(n5647) );
  NAND2_X1 U6656 ( .A1(n5647), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5645) );
  OR2_X1 U6657 ( .A1(n5646), .A2(n10196), .ZN(n5648) );
  NAND2_X1 U6658 ( .A1(n9661), .A2(n9597), .ZN(n6091) );
  NAND2_X1 U6659 ( .A1(n6039), .A2(n6091), .ZN(n5649) );
  NAND2_X1 U6660 ( .A1(n5649), .A2(n5860), .ZN(n5844) );
  NAND2_X1 U6661 ( .A1(n5656), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5653) );
  NAND2_X2 U6662 ( .A1(n5654), .A2(n5078), .ZN(n10452) );
  MUX2_X1 U6663 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5655), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n5657) );
  NAND2_X1 U6664 ( .A1(n5844), .A2(n6537), .ZN(n5845) );
  NAND2_X1 U6665 ( .A1(n5845), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  NOR2_X1 U6666 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5662) );
  NOR2_X1 U6667 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5661) );
  NOR2_X1 U6668 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5660) );
  NAND4_X1 U6669 ( .A1(n6057), .A2(n5662), .A3(n5661), .A4(n5660), .ZN(n5666)
         );
  NOR2_X1 U6670 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5664) );
  NAND4_X1 U6671 ( .A1(n5664), .A2(n6485), .A3(n5663), .A4(n6445), .ZN(n5665)
         );
  MUX2_X1 U6672 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5673), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5675) );
  INV_X1 U6673 ( .A(n5809), .ZN(n5674) );
  NAND2_X1 U6674 ( .A1(n5672), .A2(n5676), .ZN(n5677) );
  NAND2_X1 U6675 ( .A1(n5677), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5678) );
  INV_X1 U6676 ( .A(n6492), .ZN(n7891) );
  NOR2_X1 U6677 ( .A1(n7929), .A2(n7891), .ZN(n5679) );
  OR2_X1 U6678 ( .A1(n5680), .A2(n5361), .ZN(n5681) );
  NAND2_X1 U6679 ( .A1(n5682), .A2(n5681), .ZN(n6489) );
  NAND2_X1 U6680 ( .A1(n7684), .A2(n5684), .ZN(n5686) );
  NAND2_X1 U6681 ( .A1(n5687), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n5688) );
  NOR2_X1 U6682 ( .A1(n7966), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9149) );
  INV_X2 U6683 ( .A(n9149), .ZN(n9151) );
  AND2_X1 U6684 ( .A1(n7966), .A2(P2_U3152), .ZN(n7663) );
  INV_X2 U6685 ( .A(n7663), .ZN(n9153) );
  INV_X1 U6686 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6023) );
  INV_X1 U6687 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5689) );
  INV_X1 U6688 ( .A(SI_0_), .ZN(n6022) );
  NAND2_X1 U6689 ( .A1(n5690), .A2(SI_1_), .ZN(n5699) );
  OR2_X1 U6690 ( .A1(n5690), .A2(SI_1_), .ZN(n5691) );
  AND2_X1 U6691 ( .A1(n5699), .A2(n5691), .ZN(n5692) );
  NAND2_X1 U6692 ( .A1(n5692), .A2(n5693), .ZN(n5700) );
  INV_X1 U6693 ( .A(n5692), .ZN(n5695) );
  INV_X1 U6694 ( .A(n5693), .ZN(n5694) );
  NAND2_X1 U6695 ( .A1(n5695), .A2(n5694), .ZN(n5696) );
  NAND2_X1 U6696 ( .A1(n5700), .A2(n5696), .ZN(n6511) );
  NAND2_X1 U6697 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5697) );
  INV_X1 U6698 ( .A(n10600), .ZN(n6512) );
  OAI222_X1 U6699 ( .A1(n9151), .A2(n5145), .B1(n9153), .B2(n6511), .C1(
        P2_U3152), .C2(n6512), .ZN(P2_U3357) );
  INV_X1 U6700 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5705) );
  NAND2_X1 U6701 ( .A1(n5700), .A2(n5699), .ZN(n5709) );
  INV_X1 U6702 ( .A(SI_2_), .ZN(n10276) );
  NAND2_X1 U6703 ( .A1(n5703), .A2(SI_2_), .ZN(n5711) );
  AND2_X2 U6704 ( .A1(n5704), .A2(n5711), .ZN(n5710) );
  XNOR2_X1 U6705 ( .A(n5709), .B(n5710), .ZN(n6703) );
  OAI222_X1 U6706 ( .A1(n6701), .A2(P2_U3152), .B1(n9153), .B2(n6703), .C1(
        n9151), .C2(n5702), .ZN(P2_U3356) );
  NAND2_X1 U6707 ( .A1(n5706), .A2(n5705), .ZN(n5707) );
  NAND2_X1 U6708 ( .A1(n5707), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5708) );
  XNOR2_X1 U6709 ( .A(n5708), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6714) );
  INV_X1 U6710 ( .A(n6714), .ZN(n6342) );
  NAND2_X1 U6711 ( .A1(n5714), .A2(SI_3_), .ZN(n5738) );
  INV_X1 U6712 ( .A(n5714), .ZN(n5715) );
  INV_X1 U6713 ( .A(SI_3_), .ZN(n10063) );
  NAND2_X1 U6714 ( .A1(n5715), .A2(n10063), .ZN(n5716) );
  XNOR2_X1 U6715 ( .A(n5718), .B(n5737), .ZN(n6713) );
  OAI222_X1 U6716 ( .A1(n6342), .A2(P2_U3152), .B1(n9153), .B2(n6713), .C1(
        n9151), .C2(n5199), .ZN(P2_U3355) );
  MUX2_X1 U6717 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5713), .Z(n5719) );
  INV_X1 U6718 ( .A(n5719), .ZN(n5717) );
  INV_X1 U6719 ( .A(SI_4_), .ZN(n10271) );
  NAND2_X1 U6720 ( .A1(n5717), .A2(n10271), .ZN(n5740) );
  INV_X1 U6721 ( .A(n5740), .ZN(n5721) );
  NAND2_X1 U6722 ( .A1(n5719), .A2(SI_4_), .ZN(n5741) );
  AND2_X1 U6723 ( .A1(n5738), .A2(n5741), .ZN(n5720) );
  MUX2_X1 U6724 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n7958), .Z(n5723) );
  NAND2_X1 U6725 ( .A1(n5723), .A2(SI_5_), .ZN(n5758) );
  INV_X1 U6726 ( .A(n5723), .ZN(n5725) );
  INV_X1 U6727 ( .A(SI_5_), .ZN(n5724) );
  NAND2_X1 U6728 ( .A1(n5725), .A2(n5724), .ZN(n5726) );
  AND2_X1 U6729 ( .A1(n5758), .A2(n5726), .ZN(n5727) );
  NAND2_X1 U6730 ( .A1(n5728), .A2(n5727), .ZN(n5759) );
  OR2_X1 U6731 ( .A1(n5728), .A2(n5727), .ZN(n5729) );
  NAND2_X1 U6732 ( .A1(n5759), .A2(n5729), .ZN(n6945) );
  OR2_X1 U6733 ( .A1(n5730), .A2(n5884), .ZN(n5731) );
  OAI21_X1 U6734 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(P1_IR_REG_0__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5773) );
  AND2_X1 U6735 ( .A1(n5731), .A2(n5773), .ZN(n5776) );
  INV_X1 U6736 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5732) );
  NAND2_X1 U6737 ( .A1(n5776), .A2(n5732), .ZN(n5779) );
  NAND2_X1 U6738 ( .A1(n5779), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5733) );
  XNOR2_X1 U6739 ( .A(n5733), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6567) );
  INV_X1 U6740 ( .A(n6567), .ZN(n5970) );
  INV_X1 U6741 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n5734) );
  OAI222_X1 U6742 ( .A1(n10451), .A2(n6945), .B1(n5970), .B2(P1_U3084), .C1(
        n5734), .C2(n10455), .ZN(P1_U3348) );
  NAND2_X1 U6743 ( .A1(n5735), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5736) );
  XNOR2_X1 U6744 ( .A(n5736), .B(n5658), .ZN(n6728) );
  NAND2_X1 U6745 ( .A1(n5718), .A2(n5737), .ZN(n5739) );
  NAND2_X1 U6746 ( .A1(n5739), .A2(n5738), .ZN(n5743) );
  AND2_X1 U6747 ( .A1(n5741), .A2(n5740), .ZN(n5742) );
  XNOR2_X1 U6748 ( .A(n5743), .B(n5742), .ZN(n6725) );
  INV_X1 U6749 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5894) );
  OAI222_X1 U6750 ( .A1(n6728), .A2(P2_U3152), .B1(n9153), .B2(n6725), .C1(
        n9151), .C2(n5894), .ZN(P2_U3354) );
  NAND2_X1 U6751 ( .A1(n5744), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5745) );
  MUX2_X1 U6752 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5745), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n5748) );
  INV_X1 U6753 ( .A(n5746), .ZN(n5747) );
  INV_X1 U6754 ( .A(n6948), .ZN(n6307) );
  INV_X1 U6755 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6947) );
  OAI222_X1 U6756 ( .A1(P2_U3152), .A2(n6307), .B1(n9153), .B2(n6945), .C1(
        n6947), .C2(n9151), .ZN(P2_U3353) );
  NAND2_X1 U6757 ( .A1(n7888), .A2(P1_B_REG_SCAN_IN), .ZN(n5749) );
  MUX2_X1 U6758 ( .A(P1_B_REG_SCAN_IN), .B(n5749), .S(n7701), .Z(n5752) );
  INV_X1 U6759 ( .A(n5750), .ZN(n5751) );
  INV_X1 U6760 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10214) );
  NAND2_X1 U6761 ( .A1(n10018), .A2(n10214), .ZN(n5754) );
  NAND2_X1 U6762 ( .A1(n5750), .A2(n7888), .ZN(n5753) );
  NAND2_X1 U6763 ( .A1(n5754), .A2(n5753), .ZN(n6063) );
  INV_X1 U6764 ( .A(n5755), .ZN(n5756) );
  NAND2_X1 U6765 ( .A1(n10441), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5757) );
  OAI21_X1 U6766 ( .B1(n6063), .B2(n10441), .A(n5757), .ZN(P1_U3441) );
  NAND2_X1 U6767 ( .A1(n5759), .A2(n5758), .ZN(n5765) );
  MUX2_X1 U6768 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7958), .Z(n5760) );
  NAND2_X1 U6769 ( .A1(n5760), .A2(SI_6_), .ZN(n5782) );
  INV_X1 U6770 ( .A(n5760), .ZN(n5762) );
  INV_X1 U6771 ( .A(SI_6_), .ZN(n5761) );
  NAND2_X1 U6772 ( .A1(n5762), .A2(n5761), .ZN(n5763) );
  AND2_X1 U6773 ( .A1(n5782), .A2(n5763), .ZN(n5764) );
  NAND2_X1 U6774 ( .A1(n5783), .A2(n5766), .ZN(n7089) );
  NAND2_X1 U6775 ( .A1(n5767), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5768) );
  MUX2_X1 U6776 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5768), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n5770) );
  AND2_X1 U6777 ( .A1(n5770), .A2(n5769), .ZN(n10513) );
  INV_X1 U6778 ( .A(n10513), .ZN(n5839) );
  INV_X1 U6779 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n5771) );
  OAI222_X1 U6780 ( .A1(n10451), .A2(n7089), .B1(n5839), .B2(P1_U3084), .C1(
        n5771), .C2(n10455), .ZN(P1_U3347) );
  OR2_X1 U6781 ( .A1(n5746), .A2(n9146), .ZN(n5772) );
  XNOR2_X1 U6782 ( .A(n5772), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7090) );
  INV_X1 U6783 ( .A(n7090), .ZN(n6353) );
  INV_X1 U6784 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7091) );
  OAI222_X1 U6785 ( .A1(P2_U3152), .A2(n6353), .B1(n9153), .B2(n7089), .C1(
        n7091), .C2(n9151), .ZN(P2_U3352) );
  INV_X1 U6786 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6148) );
  INV_X1 U6787 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n10167) );
  XNOR2_X1 U6788 ( .A(n5773), .B(n10167), .ZN(n10627) );
  OAI222_X1 U6789 ( .A1(n10455), .A2(n6148), .B1(n10451), .B2(n6703), .C1(
        P1_U3084), .C2(n10627), .ZN(P1_U3351) );
  INV_X1 U6790 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U6791 ( .A1(n5773), .A2(n10167), .ZN(n5774) );
  NAND2_X1 U6792 ( .A1(n5774), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5775) );
  XNOR2_X1 U6793 ( .A(n5775), .B(P1_IR_REG_3__SCAN_IN), .ZN(n10549) );
  INV_X1 U6794 ( .A(n10549), .ZN(n6235) );
  OAI222_X1 U6795 ( .A1(n10455), .A2(n6232), .B1(n10451), .B2(n6713), .C1(
        P1_U3084), .C2(n6235), .ZN(P1_U3350) );
  INV_X1 U6796 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n5780) );
  INV_X1 U6797 ( .A(n5776), .ZN(n5777) );
  NAND2_X1 U6798 ( .A1(n5777), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5778) );
  NAND2_X1 U6799 ( .A1(n5779), .A2(n5778), .ZN(n6536) );
  OAI222_X1 U6800 ( .A1(n10455), .A2(n5780), .B1(n10451), .B2(n6725), .C1(
        P1_U3084), .C2(n6536), .ZN(P1_U3349) );
  INV_X1 U6801 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U6802 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5781) );
  XNOR2_X1 U6803 ( .A(n5781), .B(P1_IR_REG_1__SCAN_IN), .ZN(n10565) );
  INV_X1 U6804 ( .A(n10565), .ZN(n5830) );
  OAI222_X1 U6805 ( .A1(n10455), .A2(n6076), .B1(n5830), .B2(P1_U3084), .C1(
        n10451), .C2(n6511), .ZN(P1_U3352) );
  INV_X1 U6806 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n5786) );
  MUX2_X1 U6807 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7958), .Z(n5784) );
  NAND2_X1 U6808 ( .A1(n5784), .A2(SI_7_), .ZN(n5793) );
  OAI21_X1 U6809 ( .B1(n5784), .B2(SI_7_), .A(n5793), .ZN(n5790) );
  XNOR2_X1 U6810 ( .A(n5792), .B(n5790), .ZN(n7226) );
  INV_X1 U6811 ( .A(n7226), .ZN(n5789) );
  NAND2_X1 U6812 ( .A1(n5769), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5785) );
  XNOR2_X1 U6813 ( .A(n5785), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6917) );
  INV_X1 U6814 ( .A(n6917), .ZN(n5827) );
  OAI222_X1 U6815 ( .A1(n10455), .A2(n5786), .B1(n10451), .B2(n5789), .C1(
        P1_U3084), .C2(n5827), .ZN(P1_U3346) );
  OR2_X1 U6816 ( .A1(n5787), .A2(n9146), .ZN(n5788) );
  XNOR2_X1 U6817 ( .A(n5788), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7227) );
  INV_X1 U6818 ( .A(n7227), .ZN(n6330) );
  INV_X1 U6819 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n5914) );
  OAI222_X1 U6820 ( .A1(n6330), .A2(P2_U3152), .B1(n9153), .B2(n5789), .C1(
        n9151), .C2(n5914), .ZN(P2_U3351) );
  INV_X1 U6821 ( .A(n5790), .ZN(n5791) );
  MUX2_X1 U6822 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n7958), .Z(n5794) );
  NAND2_X1 U6823 ( .A1(n5794), .A2(SI_8_), .ZN(n5818) );
  INV_X1 U6824 ( .A(n5794), .ZN(n5795) );
  INV_X1 U6825 ( .A(SI_8_), .ZN(n10264) );
  NAND2_X1 U6826 ( .A1(n5795), .A2(n10264), .ZN(n5796) );
  OR2_X1 U6827 ( .A1(n5798), .A2(n5797), .ZN(n5799) );
  NAND2_X1 U6828 ( .A1(n5819), .A2(n5799), .ZN(n7232) );
  NOR2_X1 U6829 ( .A1(n5769), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5873) );
  OR2_X1 U6830 ( .A1(n5873), .A2(n5884), .ZN(n5801) );
  INV_X1 U6831 ( .A(n5801), .ZN(n5800) );
  NAND2_X1 U6832 ( .A1(n5800), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5802) );
  NAND2_X1 U6833 ( .A1(n5801), .A2(n10174), .ZN(n5822) );
  INV_X1 U6834 ( .A(n7180), .ZN(n5925) );
  INV_X1 U6835 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5803) );
  OAI222_X1 U6836 ( .A1(n10451), .A2(n7232), .B1(n5925), .B2(P1_U3084), .C1(
        n5803), .C2(n10455), .ZN(P1_U3345) );
  NAND2_X1 U6837 ( .A1(n5820), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5804) );
  XNOR2_X1 U6838 ( .A(n5804), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7233) );
  INV_X1 U6839 ( .A(n7233), .ZN(n6365) );
  INV_X1 U6840 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n5805) );
  OAI222_X1 U6841 ( .A1(P2_U3152), .A2(n6365), .B1(n9153), .B2(n7232), .C1(
        n5805), .C2(n9151), .ZN(P2_U3350) );
  NAND2_X1 U6842 ( .A1(n5807), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5808) );
  INV_X1 U6843 ( .A(n6522), .ZN(n5814) );
  XNOR2_X2 U6844 ( .A(n5813), .B(n5940), .ZN(n6278) );
  OAI21_X1 U6845 ( .B1(n10462), .B2(n5814), .A(n6729), .ZN(n5817) );
  INV_X1 U6846 ( .A(n6489), .ZN(n5815) );
  NAND2_X1 U6847 ( .A1(n5815), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8327) );
  NAND2_X1 U6848 ( .A1(n10462), .A2(n8327), .ZN(n5816) );
  NOR2_X1 U6849 ( .A1(n10606), .A2(P2_U3966), .ZN(P2_U3151) );
  MUX2_X1 U6850 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n7958), .Z(n5868) );
  XNOR2_X1 U6851 ( .A(n5868), .B(SI_9_), .ZN(n5867) );
  INV_X1 U6852 ( .A(n7370), .ZN(n5824) );
  NAND2_X1 U6853 ( .A1(n5108), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5878) );
  XNOR2_X1 U6854 ( .A(n5878), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7371) );
  AOI22_X1 U6855 ( .A1(n7371), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n9149), .ZN(n5821) );
  OAI21_X1 U6856 ( .B1(n5824), .B2(n9153), .A(n5821), .ZN(P2_U3349) );
  INV_X1 U6857 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5825) );
  NAND2_X1 U6858 ( .A1(n5822), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5823) );
  XNOR2_X1 U6859 ( .A(n5823), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10525) );
  INV_X1 U6860 ( .A(n10525), .ZN(n6101) );
  OAI222_X1 U6861 ( .A1(n10455), .A2(n5825), .B1(n10451), .B2(n5824), .C1(
        P1_U3084), .C2(n6101), .ZN(P1_U3344) );
  INV_X1 U6862 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n5828) );
  NOR2_X1 U6863 ( .A1(n6917), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5916) );
  INV_X1 U6864 ( .A(n5916), .ZN(n5826) );
  OAI21_X1 U6865 ( .B1(n5828), .B2(n5827), .A(n5826), .ZN(n5843) );
  NAND2_X1 U6866 ( .A1(n10513), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5841) );
  INV_X1 U6867 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5837) );
  MUX2_X1 U6868 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n5837), .S(n6567), .Z(n5969)
         );
  NAND2_X1 U6869 ( .A1(n6536), .A2(n6680), .ZN(n5835) );
  NAND2_X1 U6870 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(n10549), .ZN(n5833) );
  INV_X1 U6871 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5831) );
  MUX2_X1 U6872 ( .A(n5831), .B(P1_REG2_REG_2__SCAN_IN), .S(n10627), .Z(n10634) );
  INV_X1 U6873 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5829) );
  MUX2_X1 U6874 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n5829), .S(n10565), .Z(n10575) );
  NAND3_X1 U6875 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .A3(n10575), .ZN(n10574) );
  OAI21_X1 U6876 ( .B1(n5830), .B2(n5829), .A(n10574), .ZN(n10635) );
  NAND2_X1 U6877 ( .A1(n10634), .A2(n10635), .ZN(n10632) );
  OAI21_X1 U6878 ( .B1(n5831), .B2(n10627), .A(n10632), .ZN(n10557) );
  INV_X1 U6879 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5832) );
  MUX2_X1 U6880 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n5832), .S(n10549), .Z(n10556) );
  NAND2_X1 U6881 ( .A1(n10557), .A2(n10556), .ZN(n10555) );
  NAND2_X1 U6882 ( .A1(n5833), .A2(n10555), .ZN(n6174) );
  INV_X1 U6883 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6680) );
  OAI21_X1 U6884 ( .B1(n6536), .B2(n6680), .A(n5835), .ZN(n6173) );
  NOR2_X1 U6885 ( .A1(n6174), .A2(n6173), .ZN(n6172) );
  INV_X1 U6886 ( .A(n6172), .ZN(n5834) );
  NAND2_X1 U6887 ( .A1(n5835), .A2(n5834), .ZN(n5968) );
  NAND2_X1 U6888 ( .A1(n5969), .A2(n5968), .ZN(n5967) );
  INV_X1 U6889 ( .A(n5967), .ZN(n5836) );
  AOI21_X1 U6890 ( .B1(n5837), .B2(n5970), .A(n5836), .ZN(n10519) );
  INV_X1 U6891 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5840) );
  INV_X1 U6892 ( .A(n5841), .ZN(n5838) );
  AOI21_X1 U6893 ( .B1(n5840), .B2(n5839), .A(n5838), .ZN(n10520) );
  NAND2_X1 U6894 ( .A1(n10519), .A2(n10520), .ZN(n10518) );
  NAND2_X1 U6895 ( .A1(n5841), .A2(n10518), .ZN(n5842) );
  NOR2_X1 U6896 ( .A1(n5842), .A2(n5843), .ZN(n5915) );
  AOI21_X1 U6897 ( .B1(n5843), .B2(n5842), .A(n5915), .ZN(n5866) );
  NOR2_X1 U6898 ( .A1(n10503), .A2(P1_U3084), .ZN(n7939) );
  NAND2_X1 U6899 ( .A1(n5844), .A2(n7939), .ZN(n6117) );
  OR2_X1 U6900 ( .A1(n5845), .A2(P1_U3084), .ZN(n10512) );
  INV_X1 U6901 ( .A(n10512), .ZN(n5846) );
  NAND2_X1 U6902 ( .A1(n5846), .A2(n10503), .ZN(n10621) );
  INV_X1 U6903 ( .A(n10621), .ZN(n10573) );
  XOR2_X1 U6904 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n6917), .Z(n5859) );
  NAND2_X1 U6905 ( .A1(n6567), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5856) );
  OAI21_X1 U6906 ( .B1(n6567), .B2(P1_REG1_REG_5__SCAN_IN), .A(n5856), .ZN(
        n5974) );
  INV_X1 U6907 ( .A(n6536), .ZN(n5855) );
  XNOR2_X1 U6908 ( .A(n6536), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n6176) );
  INV_X1 U6909 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n5847) );
  OR2_X1 U6910 ( .A1(n10627), .A2(n5847), .ZN(n5850) );
  NAND2_X1 U6911 ( .A1(n10627), .A2(n5847), .ZN(n5848) );
  NAND2_X1 U6912 ( .A1(n5850), .A2(n5848), .ZN(n10623) );
  INV_X1 U6913 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6166) );
  INV_X1 U6914 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10502) );
  INV_X1 U6915 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n5849) );
  MUX2_X1 U6916 ( .A(n5849), .B(P1_REG1_REG_1__SCAN_IN), .S(n10565), .Z(n10564) );
  NOR3_X1 U6917 ( .A1(n6166), .A2(n10502), .A3(n10564), .ZN(n10562) );
  AOI21_X1 U6918 ( .B1(n10565), .B2(P1_REG1_REG_1__SCAN_IN), .A(n10562), .ZN(
        n10624) );
  NOR2_X1 U6919 ( .A1(n10623), .A2(n10624), .ZN(n10622) );
  INV_X1 U6920 ( .A(n5850), .ZN(n5851) );
  OR2_X1 U6921 ( .A1(n10622), .A2(n5851), .ZN(n10553) );
  OR2_X1 U6922 ( .A1(n10549), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5853) );
  NAND2_X1 U6923 ( .A1(P1_REG1_REG_3__SCAN_IN), .A2(n10549), .ZN(n5852) );
  AND2_X1 U6924 ( .A1(n5853), .A2(n5852), .ZN(n10554) );
  AND2_X1 U6925 ( .A1(n10553), .A2(n10554), .ZN(n10551) );
  AOI21_X1 U6926 ( .B1(n10549), .B2(P1_REG1_REG_3__SCAN_IN), .A(n10551), .ZN(
        n6177) );
  NAND2_X1 U6927 ( .A1(n6176), .A2(n6177), .ZN(n5854) );
  OAI21_X1 U6928 ( .B1(n5855), .B2(P1_REG1_REG_4__SCAN_IN), .A(n5854), .ZN(
        n5975) );
  NOR2_X1 U6929 ( .A1(n5974), .A2(n5975), .ZN(n5973) );
  INV_X1 U6930 ( .A(n5856), .ZN(n5857) );
  NOR2_X1 U6931 ( .A1(n5973), .A2(n5857), .ZN(n10516) );
  XNOR2_X1 U6932 ( .A(n10513), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n10515) );
  NOR2_X1 U6933 ( .A1(n10516), .A2(n10515), .ZN(n10514) );
  AOI21_X1 U6934 ( .B1(n10513), .B2(P1_REG1_REG_6__SCAN_IN), .A(n10514), .ZN(
        n5858) );
  NAND2_X1 U6935 ( .A1(n5858), .A2(n5859), .ZN(n5920) );
  OAI21_X1 U6936 ( .B1(n5859), .B2(n5858), .A(n5920), .ZN(n5862) );
  INV_X1 U6937 ( .A(n5860), .ZN(n7660) );
  NOR2_X1 U6938 ( .A1(n6039), .A2(n7660), .ZN(n5861) );
  AOI22_X1 U6939 ( .A1(n10573), .A2(n5862), .B1(n10550), .B2(
        P1_ADDR_REG_7__SCAN_IN), .ZN(n5865) );
  INV_X1 U6940 ( .A(n6117), .ZN(n5863) );
  AND2_X1 U6941 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6940) );
  AOI21_X1 U6942 ( .B1(n10566), .B2(n6917), .A(n6940), .ZN(n5864) );
  OAI211_X1 U6943 ( .C1(n5866), .C2(n7688), .A(n5865), .B(n5864), .ZN(P1_U3248) );
  INV_X1 U6944 ( .A(n5868), .ZN(n5869) );
  NAND2_X1 U6945 ( .A1(n5869), .A2(n10263), .ZN(n5870) );
  MUX2_X1 U6946 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n7958), .Z(n5989) );
  XNOR2_X1 U6947 ( .A(n5989), .B(n10047), .ZN(n5987) );
  XNOR2_X1 U6948 ( .A(n5988), .B(n5987), .ZN(n7410) );
  INV_X1 U6949 ( .A(n7410), .ZN(n5881) );
  NOR2_X1 U6950 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5872) );
  NOR2_X1 U6951 ( .A1(n5875), .A2(n5884), .ZN(n5874) );
  MUX2_X1 U6952 ( .A(n5884), .B(n5874), .S(P1_IR_REG_10__SCAN_IN), .Z(n5876)
         );
  AND2_X1 U6953 ( .A1(n5875), .A2(n10390), .ZN(n6054) );
  NOR2_X1 U6954 ( .A1(n5876), .A2(n6054), .ZN(n10544) );
  INV_X1 U6955 ( .A(n10455), .ZN(n10445) );
  AOI22_X1 U6956 ( .A1(n10544), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10445), .ZN(n5877) );
  OAI21_X1 U6957 ( .B1(n5881), .B2(n10451), .A(n5877), .ZN(P1_U3343) );
  NAND2_X1 U6958 ( .A1(n5878), .A2(n6056), .ZN(n5879) );
  NAND2_X1 U6959 ( .A1(n5879), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5999) );
  XNOR2_X1 U6960 ( .A(n5999), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7411) );
  AOI22_X1 U6961 ( .A1(n7411), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n9149), .ZN(n5880) );
  OAI21_X1 U6962 ( .B1(n5881), .B2(n9153), .A(n5880), .ZN(P2_U3348) );
  NAND2_X1 U6963 ( .A1(n5078), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5882) );
  INV_X1 U6964 ( .A(n5885), .ZN(n10443) );
  NAND2_X1 U6965 ( .A1(n6031), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5892) );
  AND2_X2 U6966 ( .A1(n5886), .A2(n5888), .ZN(n6576) );
  INV_X1 U6967 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5887) );
  XNOR2_X1 U6968 ( .A(n5887), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n6550) );
  NAND2_X1 U6969 ( .A1(n6931), .A2(n6550), .ZN(n5891) );
  AND2_X2 U6970 ( .A1(n5888), .A2(n10449), .ZN(n6932) );
  INV_X1 U6971 ( .A(n6932), .ZN(n5908) );
  NAND2_X1 U6972 ( .A1(n6932), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5890) );
  NAND2_X1 U6973 ( .A1(n6552), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5889) );
  INV_X1 U6974 ( .A(n7046), .ZN(n6669) );
  NAND2_X1 U6975 ( .A1(n6669), .A2(P1_U4006), .ZN(n5893) );
  OAI21_X1 U6976 ( .B1(P1_U4006), .B2(n5894), .A(n5893), .ZN(P1_U3559) );
  INV_X1 U6977 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7038) );
  NAND2_X1 U6978 ( .A1(n6578), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6577) );
  NOR2_X1 U6979 ( .A1(n6577), .A2(n5906), .ZN(n6929) );
  NAND2_X1 U6980 ( .A1(n6929), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7190) );
  NAND2_X1 U6981 ( .A1(n7498), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7499) );
  INV_X1 U6982 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8338) );
  INV_X1 U6983 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5895) );
  AND2_X1 U6984 ( .A1(n8341), .A2(n5895), .ZN(n5896) );
  OR2_X1 U6985 ( .A1(n5896), .A2(n8355), .ZN(n9859) );
  AOI22_X1 U6986 ( .A1(n6031), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n6933), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n5898) );
  NAND2_X1 U6987 ( .A1(n9423), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5897) );
  OAI211_X1 U6988 ( .C1(n9859), .C2(n8400), .A(n5898), .B(n5897), .ZN(n9878)
         );
  NAND2_X1 U6989 ( .A1(n9878), .A2(P1_U4006), .ZN(n5899) );
  OAI21_X1 U6990 ( .B1(n7038), .B2(P1_U4006), .A(n5899), .ZN(P1_U3573) );
  NAND2_X1 U6991 ( .A1(n6031), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5904) );
  INV_X1 U6992 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5900) );
  NAND2_X1 U6993 ( .A1(n6576), .A2(n5900), .ZN(n5903) );
  NAND2_X1 U6994 ( .A1(n6932), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5902) );
  NAND2_X1 U6995 ( .A1(n6552), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5901) );
  INV_X1 U6996 ( .A(n6671), .ZN(n6667) );
  NAND2_X1 U6997 ( .A1(n6667), .A2(P1_U4006), .ZN(n5905) );
  OAI21_X1 U6998 ( .B1(P1_U4006), .B2(n5199), .A(n5905), .ZN(P1_U3558) );
  NAND2_X1 U6999 ( .A1(n6031), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5912) );
  AND2_X1 U7000 ( .A1(n6577), .A2(n5906), .ZN(n5907) );
  NOR2_X1 U7001 ( .A1(n6929), .A2(n5907), .ZN(n7016) );
  NAND2_X1 U7002 ( .A1(n6931), .A2(n7016), .ZN(n5911) );
  NAND2_X1 U7003 ( .A1(n6933), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5910) );
  NAND2_X1 U7004 ( .A1(n9423), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5909) );
  INV_X1 U7005 ( .A(n7198), .ZN(n7211) );
  NAND2_X1 U7006 ( .A1(n7211), .A2(P1_U4006), .ZN(n5913) );
  OAI21_X1 U7007 ( .B1(P1_U4006), .B2(n5914), .A(n5913), .ZN(P1_U3562) );
  NOR2_X1 U7008 ( .A1(n5916), .A2(n5915), .ZN(n5919) );
  INV_X1 U7009 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5917) );
  AOI22_X1 U7010 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n5925), .B1(n7180), .B2(
        n5917), .ZN(n5918) );
  NOR2_X1 U7011 ( .A1(n5919), .A2(n5918), .ZN(n6108) );
  AOI21_X1 U7012 ( .B1(n5919), .B2(n5918), .A(n6108), .ZN(n5929) );
  OAI21_X1 U7013 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n6917), .A(n5920), .ZN(
        n5922) );
  INV_X1 U7014 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7304) );
  AOI22_X1 U7015 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n7180), .B1(n5925), .B2(
        n7304), .ZN(n5921) );
  NAND2_X1 U7016 ( .A1(n5921), .A2(n5922), .ZN(n6102) );
  OAI21_X1 U7017 ( .B1(n5922), .B2(n5921), .A(n6102), .ZN(n5927) );
  NAND2_X1 U7018 ( .A1(n10550), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U7019 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3084), .ZN(n5923) );
  OAI211_X1 U7020 ( .C1(n10628), .C2(n5925), .A(n5924), .B(n5923), .ZN(n5926)
         );
  AOI21_X1 U7021 ( .B1(n10573), .B2(n5927), .A(n5926), .ZN(n5928) );
  OAI21_X1 U7022 ( .B1(n5929), .B2(n7688), .A(n5928), .ZN(P1_U3249) );
  NAND2_X1 U7023 ( .A1(n6576), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5933) );
  NAND2_X1 U7024 ( .A1(n6031), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5932) );
  NAND2_X1 U7025 ( .A1(n6932), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U7026 ( .A1(n6552), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5930) );
  NAND2_X1 U7027 ( .A1(n5046), .A2(P1_U4006), .ZN(n5934) );
  OAI21_X1 U7028 ( .B1(P1_U4006), .B2(n5702), .A(n5934), .ZN(P1_U3557) );
  NAND2_X1 U7029 ( .A1(n6031), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5938) );
  NAND2_X1 U7030 ( .A1(n6552), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5937) );
  NAND2_X1 U7031 ( .A1(n6932), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5936) );
  NAND2_X1 U7032 ( .A1(n6576), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5935) );
  NAND4_X2 U7033 ( .A1(n5938), .A2(n5937), .A3(n5936), .A4(n5935), .ZN(n6207)
         );
  NAND2_X1 U7034 ( .A1(n6207), .A2(P1_U4006), .ZN(n5939) );
  OAI21_X1 U7035 ( .B1(P1_U4006), .B2(n5689), .A(n5939), .ZN(P1_U3555) );
  NAND2_X1 U7036 ( .A1(n5943), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5944) );
  MUX2_X1 U7037 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5944), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5946) );
  INV_X1 U7038 ( .A(n5945), .ZN(n9147) );
  NAND2_X1 U7039 ( .A1(n8192), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5950) );
  INV_X1 U7040 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8755) );
  OR2_X1 U7041 ( .A1(n8171), .A2(n8755), .ZN(n5949) );
  INV_X1 U7042 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n5947) );
  OR2_X1 U7043 ( .A1(n8169), .A2(n5947), .ZN(n5948) );
  AND3_X1 U7044 ( .A1(n5950), .A2(n5949), .A3(n5948), .ZN(n8789) );
  NAND2_X1 U7045 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n8708), .ZN(n5951) );
  OAI21_X1 U7046 ( .B1(n8789), .B2(n8708), .A(n5951), .ZN(P2_U3582) );
  INV_X1 U7047 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6230) );
  NAND2_X1 U7048 ( .A1(n6031), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5956) );
  AND2_X1 U7049 ( .A1(n5960), .A2(n6429), .ZN(n5952) );
  NOR2_X1 U7050 ( .A1(n7759), .A2(n5952), .ZN(n9919) );
  NAND2_X1 U7051 ( .A1(n6576), .A2(n9919), .ZN(n5955) );
  NAND2_X1 U7052 ( .A1(n6933), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5954) );
  NAND2_X1 U7053 ( .A1(n9423), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5953) );
  INV_X1 U7054 ( .A(n9403), .ZN(n7782) );
  NAND2_X1 U7055 ( .A1(n7782), .A2(P1_U4006), .ZN(n5957) );
  OAI21_X1 U7056 ( .B1(n6230), .B2(P1_U4006), .A(n5957), .ZN(P1_U3569) );
  INV_X1 U7057 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6129) );
  NAND2_X1 U7058 ( .A1(n7499), .A2(n5958), .ZN(n5959) );
  NAND2_X1 U7059 ( .A1(n5960), .A2(n5959), .ZN(n7796) );
  INV_X1 U7060 ( .A(n7796), .ZN(n5961) );
  NAND2_X1 U7061 ( .A1(n6576), .A2(n5961), .ZN(n5965) );
  NAND2_X1 U7062 ( .A1(n6031), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U7063 ( .A1(n6933), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5963) );
  NAND2_X1 U7064 ( .A1(n9423), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5962) );
  INV_X1 U7065 ( .A(n9260), .ZN(n9913) );
  NAND2_X1 U7066 ( .A1(n9913), .A2(P1_U4006), .ZN(n5966) );
  OAI21_X1 U7067 ( .B1(n6129), .B2(P1_U4006), .A(n5966), .ZN(P1_U3568) );
  INV_X1 U7068 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n5979) );
  OAI21_X1 U7069 ( .B1(n5969), .B2(n5968), .A(n5967), .ZN(n5972) );
  AND2_X1 U7070 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6585) );
  NOR2_X1 U7071 ( .A1(n10628), .A2(n5970), .ZN(n5971) );
  AOI211_X1 U7072 ( .C1(n10633), .C2(n5972), .A(n6585), .B(n5971), .ZN(n5978)
         );
  AOI211_X1 U7073 ( .C1(n5975), .C2(n5974), .A(n5973), .B(n10621), .ZN(n5976)
         );
  INV_X1 U7074 ( .A(n5976), .ZN(n5977) );
  OAI211_X1 U7075 ( .C1(n5979), .C2(n10626), .A(n5978), .B(n5977), .ZN(
        P1_U3246) );
  INV_X1 U7076 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6003) );
  NAND2_X1 U7077 ( .A1(n6031), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5985) );
  AND2_X1 U7078 ( .A1(n7277), .A2(n5980), .ZN(n5981) );
  NOR2_X1 U7079 ( .A1(n7498), .A2(n5981), .ZN(n10777) );
  NAND2_X1 U7080 ( .A1(n6931), .A2(n10777), .ZN(n5984) );
  NAND2_X1 U7081 ( .A1(n6933), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5983) );
  NAND2_X1 U7082 ( .A1(n9423), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5982) );
  INV_X1 U7083 ( .A(n7651), .ZN(n7637) );
  NAND2_X1 U7084 ( .A1(n7637), .A2(P1_U4006), .ZN(n5986) );
  OAI21_X1 U7085 ( .B1(n6003), .B2(P1_U4006), .A(n5986), .ZN(P1_U3566) );
  INV_X1 U7086 ( .A(n5989), .ZN(n5990) );
  NAND2_X1 U7087 ( .A1(n5990), .A2(n10047), .ZN(n5991) );
  MUX2_X1 U7088 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n5713), .Z(n5992) );
  NAND2_X1 U7089 ( .A1(n5992), .A2(SI_11_), .ZN(n6046) );
  INV_X1 U7090 ( .A(n5992), .ZN(n5994) );
  INV_X1 U7091 ( .A(SI_11_), .ZN(n5993) );
  NAND2_X1 U7092 ( .A1(n5994), .A2(n5993), .ZN(n5995) );
  XNOR2_X1 U7093 ( .A(n6045), .B(n5623), .ZN(n7534) );
  INV_X1 U7094 ( .A(n7534), .ZN(n6002) );
  OR2_X1 U7095 ( .A1(n6054), .A2(n5884), .ZN(n5996) );
  XNOR2_X1 U7096 ( .A(n5996), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7491) );
  INV_X1 U7097 ( .A(n7491), .ZN(n6112) );
  INV_X1 U7098 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5997) );
  OAI222_X1 U7099 ( .A1(n10451), .A2(n6002), .B1(n6112), .B2(P1_U3084), .C1(
        n5997), .C2(n10455), .ZN(P1_U3342) );
  INV_X1 U7100 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5998) );
  NAND2_X1 U7101 ( .A1(n5999), .A2(n5998), .ZN(n6000) );
  NAND2_X1 U7102 ( .A1(n6000), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6001) );
  XNOR2_X1 U7103 ( .A(n6001), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7535) );
  INV_X1 U7104 ( .A(n7535), .ZN(n7057) );
  OAI222_X1 U7105 ( .A1(n7057), .A2(P2_U3152), .B1(n9151), .B2(n6003), .C1(
        n6002), .C2(n9153), .ZN(P2_U3347) );
  NOR4_X1 U7106 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_27__SCAN_IN), .ZN(n6012) );
  NOR4_X1 U7107 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n6011) );
  OR4_X1 U7108 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6009) );
  NOR4_X1 U7109 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n6007) );
  NOR4_X1 U7110 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n6006) );
  NOR4_X1 U7111 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n6005) );
  NOR4_X1 U7112 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n6004) );
  NAND4_X1 U7113 ( .A1(n6007), .A2(n6006), .A3(n6005), .A4(n6004), .ZN(n6008)
         );
  NOR4_X1 U7114 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        n6009), .A4(n6008), .ZN(n6010) );
  NAND3_X1 U7115 ( .A1(n6012), .A2(n6011), .A3(n6010), .ZN(n6013) );
  NAND2_X1 U7116 ( .A1(n10018), .A2(n6013), .ZN(n6062) );
  INV_X1 U7117 ( .A(n6062), .ZN(n6014) );
  NOR2_X1 U7118 ( .A1(n6014), .A2(n6063), .ZN(n6625) );
  INV_X1 U7119 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10213) );
  NAND2_X1 U7120 ( .A1(n10018), .A2(n10213), .ZN(n6016) );
  NAND2_X1 U7121 ( .A1(n5750), .A2(n7701), .ZN(n6015) );
  AND2_X1 U7122 ( .A1(n6625), .A2(n10442), .ZN(n6025) );
  NAND2_X1 U7123 ( .A1(n6025), .A2(n10020), .ZN(n6094) );
  NAND2_X1 U7124 ( .A1(n6630), .A2(n9657), .ZN(n6628) );
  OR2_X1 U7125 ( .A1(n6094), .A2(n6628), .ZN(n6021) );
  NAND2_X1 U7126 ( .A1(n5087), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6020) );
  NOR2_X1 U7127 ( .A1(n7966), .A2(n6022), .ZN(n6024) );
  XNOR2_X1 U7128 ( .A(n6024), .B(n6023), .ZN(n10456) );
  INV_X1 U7129 ( .A(n6025), .ZN(n6026) );
  NAND2_X1 U7130 ( .A1(n6026), .A2(n6061), .ZN(n6029) );
  NAND2_X1 U7131 ( .A1(n7264), .A2(n9812), .ZN(n6092) );
  AND2_X1 U7132 ( .A1(n9598), .A2(n6092), .ZN(n6060) );
  NOR2_X1 U7133 ( .A1(n6060), .A2(n7660), .ZN(n6027) );
  AND2_X1 U7134 ( .A1(n6027), .A2(n6039), .ZN(n6028) );
  NAND2_X1 U7135 ( .A1(n6029), .A2(n6028), .ZN(n6243) );
  NOR2_X1 U7136 ( .A1(n6243), .A2(P1_U3084), .ZN(n6161) );
  INV_X1 U7137 ( .A(n6161), .ZN(n6097) );
  OR2_X1 U7138 ( .A1(n10753), .A2(n6092), .ZN(n6030) );
  INV_X1 U7139 ( .A(n9388), .ZN(n9406) );
  NAND2_X1 U7140 ( .A1(n6576), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6032) );
  AOI22_X1 U7141 ( .A1(n6097), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n9406), .B2(
        n6208), .ZN(n6044) );
  OR2_X1 U7142 ( .A1(n10877), .A2(n9598), .ZN(n6033) );
  INV_X1 U7143 ( .A(n6626), .ZN(n6034) );
  NAND2_X1 U7144 ( .A1(n6207), .A2(n6147), .ZN(n6037) );
  INV_X1 U7145 ( .A(n6039), .ZN(n6035) );
  NAND2_X1 U7146 ( .A1(n6037), .A2(n6036), .ZN(n6084) );
  NOR2_X1 U7147 ( .A1(n9661), .A2(n6092), .ZN(n6038) );
  NAND2_X1 U7148 ( .A1(n6207), .A2(n9239), .ZN(n6042) );
  NOR2_X1 U7149 ( .A1(n6039), .A2(n6166), .ZN(n6040) );
  AOI21_X1 U7150 ( .B1(n6820), .B2(n6147), .A(n6040), .ZN(n6041) );
  XNOR2_X1 U7151 ( .A(n6084), .B(n6082), .ZN(n6168) );
  NAND2_X1 U7152 ( .A1(n9376), .A2(n6168), .ZN(n6043) );
  OAI211_X1 U7153 ( .C1(n9384), .C2(n6855), .A(n6044), .B(n6043), .ZN(P1_U3230) );
  MUX2_X1 U7154 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n7958), .Z(n6048) );
  NAND2_X1 U7155 ( .A1(n6048), .A2(SI_12_), .ZN(n6127) );
  INV_X1 U7156 ( .A(n6048), .ZN(n6049) );
  NAND2_X1 U7157 ( .A1(n6049), .A2(n10254), .ZN(n6050) );
  NAND2_X1 U7158 ( .A1(n6128), .A2(n6053), .ZN(n7573) );
  NAND2_X1 U7159 ( .A1(n6054), .A2(n10391), .ZN(n6413) );
  NAND2_X1 U7160 ( .A1(n6413), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6130) );
  XNOR2_X1 U7161 ( .A(n6130), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7517) );
  INV_X1 U7162 ( .A(n7517), .ZN(n6188) );
  INV_X1 U7163 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6055) );
  OAI222_X1 U7164 ( .A1(n10451), .A2(n7573), .B1(n6188), .B2(P1_U3084), .C1(
        n6055), .C2(n10455), .ZN(P1_U3341) );
  NAND2_X1 U7165 ( .A1(n6126), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6058) );
  XNOR2_X1 U7166 ( .A(n6058), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7574) );
  INV_X1 U7167 ( .A(n7574), .ZN(n7152) );
  INV_X1 U7168 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6059) );
  OAI222_X1 U7169 ( .A1(P2_U3152), .A2(n7152), .B1(n9153), .B2(n7573), .C1(
        n6059), .C2(n9151), .ZN(P2_U3346) );
  NOR2_X1 U7170 ( .A1(n10441), .A2(n6060), .ZN(n6624) );
  AND2_X1 U7171 ( .A1(n6062), .A2(n6061), .ZN(n6064) );
  INV_X1 U7172 ( .A(n6630), .ZN(n6070) );
  NOR2_X1 U7173 ( .A1(n6207), .A2(n6855), .ZN(n6848) );
  INV_X1 U7174 ( .A(n6848), .ZN(n6065) );
  NAND2_X1 U7175 ( .A1(n6207), .A2(n6855), .ZN(n9443) );
  NAND2_X1 U7176 ( .A1(n6065), .A2(n9443), .ZN(n9626) );
  NAND2_X1 U7177 ( .A1(n9661), .A2(n9760), .ZN(n6067) );
  OR2_X1 U7178 ( .A1(n9653), .A2(n7264), .ZN(n6066) );
  NAND2_X1 U7179 ( .A1(n9596), .A2(n6626), .ZN(n6068) );
  NAND2_X1 U7180 ( .A1(n6091), .A2(n6068), .ZN(n7071) );
  NAND2_X1 U7181 ( .A1(n9888), .A2(n7071), .ZN(n6069) );
  INV_X1 U7182 ( .A(n10753), .ZN(n9910) );
  AOI22_X1 U7183 ( .A1(n9626), .A2(n6069), .B1(n9910), .B2(n6208), .ZN(n6817)
         );
  OAI21_X1 U7184 ( .B1(n6855), .B2(n6070), .A(n6817), .ZN(n6073) );
  NAND2_X1 U7185 ( .A1(n6073), .A2(n10722), .ZN(n6071) );
  OAI21_X1 U7186 ( .B1(n10722), .B2(n10502), .A(n6071), .ZN(P1_U3523) );
  INV_X1 U7187 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U7188 ( .A1(n6073), .A2(n5045), .ZN(n6074) );
  OAI21_X1 U7189 ( .B1(n5045), .B2(n6075), .A(n6074), .ZN(P1_U3454) );
  INV_X2 U7190 ( .A(n9239), .ZN(n9286) );
  OR2_X1 U7191 ( .A1(n9445), .A2(n9286), .ZN(n6081) );
  OR2_X1 U7192 ( .A1(n6149), .A2(n6076), .ZN(n6079) );
  OR2_X1 U7193 ( .A1(n5058), .A2(n6511), .ZN(n6078) );
  NAND2_X1 U7194 ( .A1(n8352), .A2(n10565), .ZN(n6077) );
  NAND2_X1 U7195 ( .A1(n9444), .A2(n9198), .ZN(n6080) );
  NAND2_X1 U7196 ( .A1(n6081), .A2(n6080), .ZN(n6143) );
  OR2_X2 U7197 ( .A1(n7071), .A2(n9760), .ZN(n10718) );
  NAND2_X1 U7198 ( .A1(n10718), .A2(n6626), .ZN(n6651) );
  NAND2_X1 U7199 ( .A1(n6082), .A2(n6084), .ZN(n6083) );
  OAI21_X1 U7200 ( .B1(n6084), .B2(n9208), .A(n6083), .ZN(n6087) );
  INV_X2 U7201 ( .A(n6147), .ZN(n9287) );
  OAI22_X1 U7202 ( .A1(n9445), .A2(n9287), .B1(n10648), .B2(n9289), .ZN(n6085)
         );
  XNOR2_X1 U7203 ( .A(n6085), .B(n9208), .ZN(n6086) );
  NAND2_X1 U7204 ( .A1(n6087), .A2(n6086), .ZN(n6144) );
  INV_X1 U7205 ( .A(n6086), .ZN(n6089) );
  INV_X1 U7206 ( .A(n6087), .ZN(n6088) );
  NAND2_X1 U7207 ( .A1(n6089), .A2(n6088), .ZN(n6145) );
  NAND2_X1 U7208 ( .A1(n6144), .A2(n6145), .ZN(n6090) );
  XOR2_X1 U7209 ( .A(n6143), .B(n6090), .Z(n6099) );
  INV_X1 U7210 ( .A(n6207), .ZN(n6850) );
  INV_X1 U7211 ( .A(n6092), .ZN(n9659) );
  NAND2_X1 U7212 ( .A1(n9912), .A2(n9659), .ZN(n6093) );
  OAI22_X1 U7213 ( .A1(n6850), .A2(n9402), .B1(n9388), .B2(n6849), .ZN(n6096)
         );
  NOR2_X1 U7214 ( .A1(n9384), .A2(n10648), .ZN(n6095) );
  AOI211_X1 U7215 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n6097), .A(n6096), .B(
        n6095), .ZN(n6098) );
  OAI21_X1 U7216 ( .B1(n6099), .B2(n9410), .A(n6098), .ZN(P1_U3220) );
  INV_X1 U7217 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6100) );
  MUX2_X1 U7218 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n6100), .S(n7491), .Z(n6105)
         );
  INV_X1 U7219 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10721) );
  AOI22_X1 U7220 ( .A1(n10525), .A2(P1_REG1_REG_9__SCAN_IN), .B1(n10721), .B2(
        n6101), .ZN(n10527) );
  OAI21_X1 U7221 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n7180), .A(n6102), .ZN(
        n10528) );
  NAND2_X1 U7222 ( .A1(n10527), .A2(n10528), .ZN(n10526) );
  OAI21_X1 U7223 ( .B1(n10525), .B2(P1_REG1_REG_9__SCAN_IN), .A(n10526), .ZN(
        n10539) );
  INV_X1 U7224 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6103) );
  MUX2_X1 U7225 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6103), .S(n10544), .Z(
        n10538) );
  NAND2_X1 U7226 ( .A1(n10539), .A2(n10538), .ZN(n10537) );
  OAI21_X1 U7227 ( .B1(n10544), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10537), .ZN(
        n6104) );
  NAND2_X1 U7228 ( .A1(n6104), .A2(n6105), .ZN(n6184) );
  OAI21_X1 U7229 ( .B1(n6105), .B2(n6104), .A(n6184), .ZN(n6124) );
  NAND2_X1 U7230 ( .A1(n10525), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6109) );
  INV_X1 U7231 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6106) );
  MUX2_X1 U7232 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n6106), .S(n10525), .Z(n10531) );
  NOR2_X1 U7233 ( .A1(n7180), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6107) );
  NOR2_X1 U7234 ( .A1(n6108), .A2(n6107), .ZN(n10532) );
  NAND2_X1 U7235 ( .A1(n10531), .A2(n10532), .ZN(n10530) );
  NAND2_X1 U7236 ( .A1(n6109), .A2(n10530), .ZN(n10543) );
  INV_X1 U7237 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6110) );
  MUX2_X1 U7238 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n6110), .S(n10544), .Z(
        n10542) );
  NAND2_X1 U7239 ( .A1(n10543), .A2(n10542), .ZN(n10541) );
  NAND2_X1 U7240 ( .A1(n10544), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6111) );
  NAND2_X1 U7241 ( .A1(n10541), .A2(n6111), .ZN(n6116) );
  INV_X1 U7242 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6118) );
  NOR2_X1 U7243 ( .A1(n6112), .A2(n6118), .ZN(n6113) );
  OAI22_X1 U7244 ( .A1(n6116), .A2(n6113), .B1(P1_REG2_REG_11__SCAN_IN), .B2(
        n7491), .ZN(n6191) );
  INV_X1 U7245 ( .A(n6191), .ZN(n6115) );
  NOR3_X1 U7246 ( .A1(n6116), .A2(n7491), .A3(P1_REG2_REG_11__SCAN_IN), .ZN(
        n6114) );
  NOR3_X1 U7247 ( .A1(n6115), .A2(n6114), .A3(n7688), .ZN(n6123) );
  INV_X1 U7248 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7590) );
  INV_X1 U7249 ( .A(n6116), .ZN(n6119) );
  NOR3_X1 U7250 ( .A1(n6119), .A2(n6118), .A3(n6117), .ZN(n6120) );
  OAI21_X1 U7251 ( .B1(n6120), .B2(n10566), .A(n7491), .ZN(n6121) );
  NAND2_X1 U7252 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3084), .ZN(n7505) );
  OAI211_X1 U7253 ( .C1(n7590), .C2(n10626), .A(n6121), .B(n7505), .ZN(n6122)
         );
  AOI211_X1 U7254 ( .C1(n10573), .C2(n6124), .A(n6123), .B(n6122), .ZN(n6125)
         );
  INV_X1 U7255 ( .A(n6125), .ZN(P1_U3252) );
  OR2_X1 U7256 ( .A1(n6447), .A2(n9146), .ZN(n6227) );
  XNOR2_X1 U7257 ( .A(n6227), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7813) );
  INV_X1 U7258 ( .A(n7813), .ZN(n7287) );
  MUX2_X1 U7259 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n5713), .Z(n6196) );
  XNOR2_X1 U7260 ( .A(n6196), .B(SI_13_), .ZN(n6198) );
  XNOR2_X1 U7261 ( .A(n6199), .B(n6198), .ZN(n7812) );
  INV_X1 U7262 ( .A(n7812), .ZN(n6134) );
  OAI222_X1 U7263 ( .A1(n7287), .A2(P2_U3152), .B1(n9153), .B2(n6134), .C1(
        n9151), .C2(n6129), .ZN(P2_U3345) );
  INV_X1 U7264 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7265 ( .A1(n6130), .A2(n10396), .ZN(n6131) );
  NAND2_X1 U7266 ( .A1(n6131), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6132) );
  NAND2_X1 U7267 ( .A1(n6132), .A2(n10397), .ZN(n6204) );
  OR2_X1 U7268 ( .A1(n6132), .A2(n10397), .ZN(n6133) );
  INV_X1 U7269 ( .A(n7721), .ZN(n6254) );
  OAI222_X1 U7270 ( .A1(n10455), .A2(n6135), .B1(n10451), .B2(n6134), .C1(
        P1_U3084), .C2(n6254), .ZN(P1_U3340) );
  INV_X1 U7271 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7473) );
  NAND2_X1 U7272 ( .A1(n8355), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8365) );
  INV_X1 U7273 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9356) );
  INV_X1 U7274 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9304) );
  INV_X1 U7275 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9367) );
  AND2_X1 U7276 ( .A1(n8377), .A2(n9367), .ZN(n6136) );
  OR2_X1 U7277 ( .A1(n6136), .A2(n8393), .ZN(n9784) );
  INV_X1 U7278 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n6139) );
  INV_X1 U7279 ( .A(n6031), .ZN(n8412) );
  NAND2_X1 U7280 ( .A1(n6933), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U7281 ( .A1(n9423), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6137) );
  OAI211_X1 U7282 ( .C1(n6139), .C2(n8412), .A(n6138), .B(n6137), .ZN(n6140)
         );
  INV_X1 U7283 ( .A(n6140), .ZN(n6141) );
  OAI21_X1 U7284 ( .B1(n9784), .B2(n8400), .A(n6141), .ZN(n9775) );
  NAND2_X1 U7285 ( .A1(n9775), .A2(P1_U4006), .ZN(n6142) );
  OAI21_X1 U7286 ( .B1(n7473), .B2(P1_U4006), .A(n6142), .ZN(P1_U3577) );
  NAND2_X1 U7287 ( .A1(n6144), .A2(n6143), .ZN(n6146) );
  AND2_X1 U7288 ( .A1(n6146), .A2(n6145), .ZN(n6159) );
  OAI22_X1 U7289 ( .A1(n6849), .A2(n9287), .B1(n6160), .B2(n9289), .ZN(n6150)
         );
  XNOR2_X1 U7290 ( .A(n6150), .B(n9208), .ZN(n6156) );
  INV_X1 U7291 ( .A(n6156), .ZN(n6153) );
  NAND2_X1 U7292 ( .A1(n6220), .A2(n9198), .ZN(n6151) );
  INV_X1 U7293 ( .A(n6154), .ZN(n6155) );
  NAND2_X1 U7294 ( .A1(n6156), .A2(n6155), .ZN(n6239) );
  NAND2_X1 U7295 ( .A1(n6159), .A2(n6158), .ZN(n6240) );
  OAI21_X1 U7296 ( .B1(n6159), .B2(n6158), .A(n6240), .ZN(n6164) );
  OAI22_X1 U7297 ( .A1(n9445), .A2(n9402), .B1(n9388), .B2(n6671), .ZN(n6163)
         );
  INV_X1 U7298 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10638) );
  OAI22_X1 U7299 ( .A1(n9384), .A2(n6160), .B1(n6161), .B2(n10638), .ZN(n6162)
         );
  AOI211_X1 U7300 ( .C1(n6164), .C2(n9376), .A(n6163), .B(n6162), .ZN(n6165)
         );
  INV_X1 U7301 ( .A(n6165), .ZN(P1_U3235) );
  INV_X1 U7302 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6823) );
  NOR2_X1 U7303 ( .A1(n6166), .A2(n6823), .ZN(n10576) );
  INV_X1 U7304 ( .A(n10576), .ZN(n6167) );
  INV_X1 U7305 ( .A(n10503), .ZN(n9676) );
  MUX2_X1 U7306 ( .A(n6168), .B(n6167), .S(n9676), .Z(n6169) );
  NOR2_X1 U7307 ( .A1(n6169), .A2(n10452), .ZN(n6171) );
  NOR2_X1 U7308 ( .A1(n10503), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6170) );
  NOR2_X1 U7309 ( .A1(n10452), .A2(n6170), .ZN(n10504) );
  NOR2_X1 U7310 ( .A1(n10504), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n10501) );
  NOR3_X1 U7311 ( .A1(n6171), .A2(n10501), .A3(n9674), .ZN(n10631) );
  AOI21_X1 U7312 ( .B1(n6174), .B2(n6173), .A(n6172), .ZN(n6175) );
  NOR2_X1 U7313 ( .A1(n7688), .A2(n6175), .ZN(n6182) );
  NAND2_X1 U7314 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n6557) );
  OAI21_X1 U7315 ( .B1(n10628), .B2(n6536), .A(n6557), .ZN(n6181) );
  XOR2_X1 U7316 ( .A(n6177), .B(n6176), .Z(n6179) );
  INV_X1 U7317 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n6178) );
  OAI22_X1 U7318 ( .A1(n10621), .A2(n6179), .B1(n10626), .B2(n6178), .ZN(n6180) );
  OR4_X1 U7319 ( .A1(n10631), .A2(n6182), .A3(n6181), .A4(n6180), .ZN(P1_U3245) );
  INV_X1 U7320 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6183) );
  MUX2_X1 U7321 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6183), .S(n7517), .Z(n6186)
         );
  OAI21_X1 U7322 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n7491), .A(n6184), .ZN(
        n6185) );
  NAND2_X1 U7323 ( .A1(n6185), .A2(n6186), .ZN(n6250) );
  OAI21_X1 U7324 ( .B1(n6186), .B2(n6185), .A(n6250), .ZN(n6194) );
  NAND2_X1 U7325 ( .A1(n10550), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6187) );
  NAND2_X1 U7326 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n7525) );
  OAI211_X1 U7327 ( .C1(n10628), .C2(n6188), .A(n6187), .B(n7525), .ZN(n6193)
         );
  NAND2_X1 U7328 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7517), .ZN(n6189) );
  OAI21_X1 U7329 ( .B1(n7517), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6189), .ZN(
        n6190) );
  NOR2_X1 U7330 ( .A1(n6191), .A2(n6190), .ZN(n6255) );
  AOI211_X1 U7331 ( .C1(n6191), .C2(n6190), .A(n7688), .B(n6255), .ZN(n6192)
         );
  AOI211_X1 U7332 ( .C1(n10573), .C2(n6194), .A(n6193), .B(n6192), .ZN(n6195)
         );
  INV_X1 U7333 ( .A(n6195), .ZN(P1_U3253) );
  INV_X1 U7334 ( .A(n6196), .ZN(n6197) );
  MUX2_X1 U7335 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n7958), .Z(n6200) );
  NAND2_X1 U7336 ( .A1(n6200), .A2(SI_14_), .ZN(n6404) );
  INV_X1 U7337 ( .A(n6200), .ZN(n6202) );
  INV_X1 U7338 ( .A(SI_14_), .ZN(n6201) );
  NAND2_X1 U7339 ( .A1(n6202), .A2(n6201), .ZN(n6203) );
  XNOR2_X1 U7340 ( .A(n6405), .B(n5127), .ZN(n7863) );
  INV_X1 U7341 ( .A(n7863), .ZN(n6229) );
  NAND2_X1 U7342 ( .A1(n6204), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6205) );
  XNOR2_X1 U7343 ( .A(n6205), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7751) );
  INV_X1 U7344 ( .A(n7751), .ZN(n6425) );
  INV_X1 U7345 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6206) );
  OAI222_X1 U7346 ( .A1(n10451), .A2(n6229), .B1(n6425), .B2(P1_U3084), .C1(
        n6206), .C2(n10455), .ZN(P1_U3339) );
  NAND2_X1 U7347 ( .A1(n9445), .A2(n10648), .ZN(n6213) );
  NAND2_X1 U7348 ( .A1(n6213), .A2(n6845), .ZN(n6209) );
  NAND2_X1 U7349 ( .A1(n6849), .A2(n6220), .ZN(n9446) );
  OR2_X1 U7350 ( .A1(n6210), .A2(n9627), .ZN(n6211) );
  NAND2_X1 U7351 ( .A1(n6211), .A2(n6666), .ZN(n6637) );
  INV_X1 U7352 ( .A(n6637), .ZN(n6222) );
  INV_X1 U7353 ( .A(n9627), .ZN(n6215) );
  NAND2_X1 U7354 ( .A1(n9445), .A2(n9444), .ZN(n6214) );
  OAI21_X1 U7355 ( .B1(n6215), .B2(n9450), .A(n6672), .ZN(n6218) );
  AOI22_X1 U7356 ( .A1(n9912), .A2(n6208), .B1(n6667), .B2(n9910), .ZN(n6216)
         );
  OAI21_X1 U7357 ( .B1(n6222), .B2(n10718), .A(n6216), .ZN(n6217) );
  AOI21_X1 U7358 ( .B1(n10758), .B2(n6218), .A(n6217), .ZN(n6639) );
  NAND2_X1 U7359 ( .A1(n10648), .A2(n6855), .ZN(n6854) );
  NOR2_X1 U7360 ( .A1(n6854), .A2(n6220), .ZN(n6678) );
  AND2_X1 U7361 ( .A1(n6854), .A2(n6220), .ZN(n6219) );
  NOR2_X1 U7362 ( .A1(n6678), .A2(n6219), .ZN(n6632) );
  AOI22_X1 U7363 ( .A1(n6632), .A2(n10878), .B1(n10877), .B2(n6220), .ZN(n6221) );
  OAI211_X1 U7364 ( .C1(n6222), .C2(n10817), .A(n6639), .B(n6221), .ZN(n6224)
         );
  NAND2_X1 U7365 ( .A1(n6224), .A2(n10722), .ZN(n6223) );
  OAI21_X1 U7366 ( .B1(n10722), .B2(n5847), .A(n6223), .ZN(P1_U3525) );
  INV_X1 U7367 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6226) );
  NAND2_X1 U7368 ( .A1(n6224), .A2(n5045), .ZN(n6225) );
  OAI21_X1 U7369 ( .B1(n5045), .B2(n6226), .A(n6225), .ZN(P1_U3460) );
  NAND2_X1 U7370 ( .A1(n6227), .A2(n6445), .ZN(n6228) );
  NAND2_X1 U7371 ( .A1(n6228), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6416) );
  XNOR2_X1 U7372 ( .A(n6416), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7864) );
  INV_X1 U7373 ( .A(n7864), .ZN(n7559) );
  OAI222_X1 U7374 ( .A1(n7559), .A2(P2_U3152), .B1(n9151), .B2(n6230), .C1(
        n6229), .C2(n9153), .ZN(P2_U3344) );
  OR2_X1 U7375 ( .A1(n6231), .A2(n6713), .ZN(n6234) );
  OR2_X1 U7376 ( .A1(n6149), .A2(n6232), .ZN(n6233) );
  OAI211_X1 U7377 ( .C1(n6537), .C2(n6235), .A(n6234), .B(n6233), .ZN(n6813)
         );
  OAI22_X1 U7378 ( .A1(n6671), .A2(n9287), .B1(n10662), .B2(n9289), .ZN(n6236)
         );
  XNOR2_X1 U7379 ( .A(n6236), .B(n9208), .ZN(n6543) );
  OR2_X1 U7380 ( .A1(n6671), .A2(n9286), .ZN(n6238) );
  NAND2_X1 U7381 ( .A1(n6813), .A2(n9198), .ZN(n6237) );
  NAND2_X1 U7382 ( .A1(n6238), .A2(n6237), .ZN(n6541) );
  XNOR2_X1 U7383 ( .A(n6543), .B(n6541), .ZN(n6242) );
  NAND2_X1 U7384 ( .A1(n6240), .A2(n6239), .ZN(n6241) );
  NAND2_X1 U7385 ( .A1(n6241), .A2(n6242), .ZN(n6545) );
  OAI21_X1 U7386 ( .B1(n6242), .B2(n6241), .A(n6545), .ZN(n6248) );
  OAI22_X1 U7387 ( .A1(n6849), .A2(n9402), .B1(n9401), .B2(
        P1_REG3_REG_3__SCAN_IN), .ZN(n6247) );
  NAND2_X1 U7388 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n10560) );
  INV_X1 U7389 ( .A(n10560), .ZN(n6244) );
  AOI21_X1 U7390 ( .B1(n9406), .B2(n6669), .A(n6244), .ZN(n6245) );
  OAI21_X1 U7391 ( .B1(n9384), .B2(n10662), .A(n6245), .ZN(n6246) );
  AOI211_X1 U7392 ( .C1(n6248), .C2(n9376), .A(n6247), .B(n6246), .ZN(n6249)
         );
  INV_X1 U7393 ( .A(n6249), .ZN(P1_U3216) );
  OAI21_X1 U7394 ( .B1(n7517), .B2(P1_REG1_REG_12__SCAN_IN), .A(n6250), .ZN(
        n6252) );
  MUX2_X1 U7395 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10838), .S(n7721), .Z(n6251) );
  NAND2_X1 U7396 ( .A1(n6251), .A2(n6252), .ZN(n6426) );
  OAI21_X1 U7397 ( .B1(n6252), .B2(n6251), .A(n6426), .ZN(n6261) );
  NAND2_X1 U7398 ( .A1(n10550), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n6253) );
  NAND2_X1 U7399 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7744) );
  OAI211_X1 U7400 ( .C1(n10628), .C2(n6254), .A(n6253), .B(n7744), .ZN(n6260)
         );
  AOI21_X1 U7401 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7517), .A(n6255), .ZN(
        n6258) );
  NAND2_X1 U7402 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7721), .ZN(n6256) );
  OAI21_X1 U7403 ( .B1(n7721), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6256), .ZN(
        n6257) );
  NOR2_X1 U7404 ( .A1(n6258), .A2(n6257), .ZN(n6421) );
  AOI211_X1 U7405 ( .C1(n6258), .C2(n6257), .A(n6421), .B(n7688), .ZN(n6259)
         );
  AOI211_X1 U7406 ( .C1(n10573), .C2(n6261), .A(n6260), .B(n6259), .ZN(n6262)
         );
  INV_X1 U7407 ( .A(n6262), .ZN(P1_U3254) );
  INV_X1 U7408 ( .A(n6728), .ZN(n6268) );
  INV_X1 U7409 ( .A(n6701), .ZN(n10612) );
  NAND2_X1 U7410 ( .A1(n10600), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6263) );
  OAI21_X1 U7411 ( .B1(n10600), .B2(P2_REG2_REG_1__SCAN_IN), .A(n6263), .ZN(
        n10596) );
  NAND2_X1 U7412 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n10597) );
  NOR2_X1 U7413 ( .A1(n10596), .A2(n10597), .ZN(n10595) );
  AOI21_X1 U7414 ( .B1(n10600), .B2(P2_REG2_REG_1__SCAN_IN), .A(n10595), .ZN(
        n10610) );
  INV_X1 U7415 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6264) );
  MUX2_X1 U7416 ( .A(n6264), .B(P2_REG2_REG_2__SCAN_IN), .S(n6701), .Z(n6265)
         );
  INV_X1 U7417 ( .A(n6265), .ZN(n10609) );
  NOR2_X1 U7418 ( .A1(n10610), .A2(n10609), .ZN(n10608) );
  INV_X1 U7419 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6708) );
  MUX2_X1 U7420 ( .A(n6708), .B(P2_REG2_REG_3__SCAN_IN), .S(n6714), .Z(n6334)
         );
  NOR2_X1 U7421 ( .A1(n6335), .A2(n6334), .ZN(n6333) );
  AOI21_X1 U7422 ( .B1(n6714), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6333), .ZN(
        n6312) );
  INV_X1 U7423 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6266) );
  MUX2_X1 U7424 ( .A(n6266), .B(P2_REG2_REG_4__SCAN_IN), .S(n6728), .Z(n6267)
         );
  INV_X1 U7425 ( .A(n6267), .ZN(n6311) );
  NOR2_X1 U7426 ( .A1(n6312), .A2(n6311), .ZN(n6310) );
  NAND2_X1 U7427 ( .A1(n6948), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6269) );
  OAI21_X1 U7428 ( .B1(n6948), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6269), .ZN(
        n6300) );
  NOR2_X1 U7429 ( .A1(n6301), .A2(n6300), .ZN(n6299) );
  AOI21_X1 U7430 ( .B1(n6948), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6299), .ZN(
        n6347) );
  NAND2_X1 U7431 ( .A1(n7090), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6270) );
  OAI21_X1 U7432 ( .B1(n7090), .B2(P2_REG2_REG_6__SCAN_IN), .A(n6270), .ZN(
        n6346) );
  NOR2_X1 U7433 ( .A1(n6347), .A2(n6346), .ZN(n6345) );
  INV_X1 U7434 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6271) );
  MUX2_X1 U7435 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n6271), .S(n7227), .Z(n6272)
         );
  INV_X1 U7436 ( .A(n6272), .ZN(n6322) );
  NOR2_X1 U7437 ( .A1(n6323), .A2(n6322), .ZN(n6321) );
  AOI21_X1 U7438 ( .B1(n7227), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6321), .ZN(
        n6358) );
  NAND2_X1 U7439 ( .A1(n7233), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6273) );
  OAI21_X1 U7440 ( .B1(n7233), .B2(P2_REG2_REG_8__SCAN_IN), .A(n6273), .ZN(
        n6357) );
  NOR2_X1 U7441 ( .A1(n6358), .A2(n6357), .ZN(n6356) );
  AOI21_X1 U7442 ( .B1(n7233), .B2(P2_REG2_REG_8__SCAN_IN), .A(n6356), .ZN(
        n6282) );
  MUX2_X1 U7443 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n7247), .S(n7371), .Z(n6274)
         );
  INV_X1 U7444 ( .A(n6274), .ZN(n6281) );
  NOR2_X1 U7445 ( .A1(n6282), .A2(n6281), .ZN(n6389) );
  OR2_X1 U7446 ( .A1(n10462), .A2(n6522), .ZN(n6617) );
  INV_X1 U7447 ( .A(n6490), .ZN(n6275) );
  NAND2_X1 U7448 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6275), .ZN(n6276) );
  NAND3_X1 U7449 ( .A1(n6617), .A2(n8327), .A3(n6276), .ZN(n6277) );
  NAND2_X1 U7450 ( .A1(n6277), .A2(n6729), .ZN(n6291) );
  NAND2_X1 U7451 ( .A1(n6291), .A2(n8708), .ZN(n6283) );
  INV_X1 U7452 ( .A(n6278), .ZN(n6523) );
  INV_X1 U7453 ( .A(n6280), .ZN(n8747) );
  AOI211_X1 U7454 ( .C1(n6282), .C2(n6281), .A(n6389), .B(n10607), .ZN(n6298)
         );
  AND2_X1 U7455 ( .A1(n6283), .A2(n6278), .ZN(n10613) );
  INV_X1 U7456 ( .A(n7371), .ZN(n6396) );
  NAND2_X1 U7457 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7447) );
  INV_X1 U7458 ( .A(n7447), .ZN(n6284) );
  AOI21_X1 U7459 ( .B1(n10606), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n6284), .ZN(
        n6296) );
  INV_X1 U7460 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10705) );
  MUX2_X1 U7461 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n10705), .S(n7233), .Z(n6361)
         );
  INV_X1 U7462 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10697) );
  MUX2_X1 U7463 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10697), .S(n7227), .Z(n6326)
         );
  NAND2_X1 U7464 ( .A1(n7090), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6289) );
  INV_X1 U7465 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6285) );
  MUX2_X1 U7466 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6285), .S(n7090), .Z(n6349)
         );
  NAND2_X1 U7467 ( .A1(n6948), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6288) );
  INV_X1 U7468 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6286) );
  MUX2_X1 U7469 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6286), .S(n6948), .Z(n6304)
         );
  INV_X1 U7470 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10674) );
  MUX2_X1 U7471 ( .A(n10674), .B(P2_REG1_REG_4__SCAN_IN), .S(n6728), .Z(n6315)
         );
  INV_X1 U7472 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6802) );
  MUX2_X1 U7473 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6802), .S(n6714), .Z(n6338)
         );
  INV_X1 U7474 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10660) );
  MUX2_X1 U7475 ( .A(n10660), .B(P2_REG1_REG_2__SCAN_IN), .S(n6701), .Z(n10616) );
  NAND2_X1 U7476 ( .A1(n10600), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6287) );
  MUX2_X1 U7477 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6533), .S(n10600), .Z(n10602) );
  NAND3_X1 U7478 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .A3(n10602), .ZN(n10601) );
  NAND2_X1 U7479 ( .A1(n6287), .A2(n10601), .ZN(n10617) );
  NAND2_X1 U7480 ( .A1(n10616), .A2(n10617), .ZN(n10614) );
  OAI21_X1 U7481 ( .B1(n6701), .B2(n10660), .A(n10614), .ZN(n6339) );
  NAND2_X1 U7482 ( .A1(n6338), .A2(n6339), .ZN(n6337) );
  OAI21_X1 U7483 ( .B1(n6342), .B2(n6802), .A(n6337), .ZN(n6316) );
  NAND2_X1 U7484 ( .A1(n6315), .A2(n6316), .ZN(n6314) );
  OAI21_X1 U7485 ( .B1(n6728), .B2(n10674), .A(n6314), .ZN(n6303) );
  NAND2_X1 U7486 ( .A1(n6304), .A2(n6303), .ZN(n6302) );
  NAND2_X1 U7487 ( .A1(n6288), .A2(n6302), .ZN(n6350) );
  NAND2_X1 U7488 ( .A1(n6349), .A2(n6350), .ZN(n6348) );
  NAND2_X1 U7489 ( .A1(n6289), .A2(n6348), .ZN(n6327) );
  NAND2_X1 U7490 ( .A1(n6326), .A2(n6327), .ZN(n6325) );
  OAI21_X1 U7491 ( .B1(n6330), .B2(n10697), .A(n6325), .ZN(n6362) );
  NAND2_X1 U7492 ( .A1(n6361), .A2(n6362), .ZN(n6360) );
  OAI21_X1 U7493 ( .B1(n6365), .B2(n10705), .A(n6360), .ZN(n6294) );
  INV_X1 U7494 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6290) );
  MUX2_X1 U7495 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n6290), .S(n7371), .Z(n6293)
         );
  INV_X1 U7496 ( .A(n6291), .ZN(n6292) );
  NAND2_X1 U7497 ( .A1(n6292), .A2(n6280), .ZN(n10586) );
  NAND2_X1 U7498 ( .A1(n6293), .A2(n6294), .ZN(n6395) );
  OAI211_X1 U7499 ( .C1(n6294), .C2(n6293), .A(n10615), .B(n6395), .ZN(n6295)
         );
  OAI211_X1 U7500 ( .C1(n10585), .C2(n6396), .A(n6296), .B(n6295), .ZN(n6297)
         );
  OR2_X1 U7501 ( .A1(n6298), .A2(n6297), .ZN(P2_U3254) );
  AOI211_X1 U7502 ( .C1(n6301), .C2(n6300), .A(n6299), .B(n10607), .ZN(n6309)
         );
  INV_X1 U7503 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10096) );
  NOR2_X1 U7504 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10096), .ZN(n6979) );
  AOI21_X1 U7505 ( .B1(n10606), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6979), .ZN(
        n6306) );
  OAI211_X1 U7506 ( .C1(n6304), .C2(n6303), .A(n10615), .B(n6302), .ZN(n6305)
         );
  OAI211_X1 U7507 ( .C1(n10585), .C2(n6307), .A(n6306), .B(n6305), .ZN(n6308)
         );
  OR2_X1 U7508 ( .A1(n6309), .A2(n6308), .ZN(P2_U3250) );
  AOI211_X1 U7509 ( .C1(n6312), .C2(n6311), .A(n6310), .B(n10607), .ZN(n6320)
         );
  INV_X1 U7510 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6313) );
  NOR2_X1 U7511 ( .A1(n6313), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6907) );
  AOI21_X1 U7512 ( .B1(n10606), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n6907), .ZN(
        n6318) );
  OAI211_X1 U7513 ( .C1(n6316), .C2(n6315), .A(n10615), .B(n6314), .ZN(n6317)
         );
  OAI211_X1 U7514 ( .C1(n10585), .C2(n6728), .A(n6318), .B(n6317), .ZN(n6319)
         );
  OR2_X1 U7515 ( .A1(n6320), .A2(n6319), .ZN(P2_U3249) );
  AOI211_X1 U7516 ( .C1(n6323), .C2(n6322), .A(n6321), .B(n10607), .ZN(n6332)
         );
  INV_X1 U7517 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8554) );
  NOR2_X1 U7518 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8554), .ZN(n6324) );
  AOI21_X1 U7519 ( .B1(n10606), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n6324), .ZN(
        n6329) );
  OAI211_X1 U7520 ( .C1(n6327), .C2(n6326), .A(n10615), .B(n6325), .ZN(n6328)
         );
  OAI211_X1 U7521 ( .C1(n10585), .C2(n6330), .A(n6329), .B(n6328), .ZN(n6331)
         );
  OR2_X1 U7522 ( .A1(n6332), .A2(n6331), .ZN(P2_U3252) );
  AOI211_X1 U7523 ( .C1(n6335), .C2(n6334), .A(n6333), .B(n10607), .ZN(n6344)
         );
  INV_X1 U7524 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10082) );
  NOR2_X1 U7525 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10082), .ZN(n6336) );
  AOI21_X1 U7526 ( .B1(n10606), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n6336), .ZN(
        n6341) );
  OAI211_X1 U7527 ( .C1(n6339), .C2(n6338), .A(n10615), .B(n6337), .ZN(n6340)
         );
  OAI211_X1 U7528 ( .C1(n10585), .C2(n6342), .A(n6341), .B(n6340), .ZN(n6343)
         );
  OR2_X1 U7529 ( .A1(n6344), .A2(n6343), .ZN(P2_U3248) );
  AOI211_X1 U7530 ( .C1(n6347), .C2(n6346), .A(n6345), .B(n10607), .ZN(n6355)
         );
  INV_X1 U7531 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10331) );
  NOR2_X1 U7532 ( .A1(n10331), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7110) );
  AOI21_X1 U7533 ( .B1(n10606), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n7110), .ZN(
        n6352) );
  OAI211_X1 U7534 ( .C1(n6350), .C2(n6349), .A(n10615), .B(n6348), .ZN(n6351)
         );
  OAI211_X1 U7535 ( .C1(n10585), .C2(n6353), .A(n6352), .B(n6351), .ZN(n6354)
         );
  OR2_X1 U7536 ( .A1(n6355), .A2(n6354), .ZN(P2_U3251) );
  AOI211_X1 U7537 ( .C1(n6358), .C2(n6357), .A(n6356), .B(n10607), .ZN(n6367)
         );
  NOR2_X1 U7538 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10293), .ZN(n6359) );
  AOI21_X1 U7539 ( .B1(n10606), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6359), .ZN(
        n6364) );
  OAI211_X1 U7540 ( .C1(n6362), .C2(n6361), .A(n10615), .B(n6360), .ZN(n6363)
         );
  OAI211_X1 U7541 ( .C1(n10585), .C2(n6365), .A(n6364), .B(n6363), .ZN(n6366)
         );
  OR2_X1 U7542 ( .A1(n6367), .A2(n6366), .ZN(P2_U3253) );
  NAND2_X1 U7543 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6737) );
  INV_X1 U7544 ( .A(n6737), .ZN(n6368) );
  NAND2_X1 U7545 ( .A1(n6368), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6952) );
  INV_X1 U7546 ( .A(n6952), .ZN(n6369) );
  NAND2_X1 U7547 ( .A1(n6369), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7103) );
  INV_X1 U7548 ( .A(n7103), .ZN(n6370) );
  NAND2_X1 U7549 ( .A1(n6370), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7236) );
  INV_X1 U7550 ( .A(n7244), .ZN(n6371) );
  NAND2_X1 U7551 ( .A1(n6371), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7373) );
  INV_X1 U7552 ( .A(n7539), .ZN(n6373) );
  AND2_X1 U7553 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n6372) );
  NAND2_X1 U7554 ( .A1(n6373), .A2(n6372), .ZN(n7564) );
  NAND2_X1 U7555 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_REG3_REG_15__SCAN_IN), 
        .ZN(n6374) );
  NAND2_X1 U7556 ( .A1(n6375), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8109) );
  INV_X1 U7557 ( .A(n8109), .ZN(n6376) );
  NAND2_X1 U7558 ( .A1(n6376), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8120) );
  INV_X1 U7559 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10117) );
  INV_X1 U7560 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10320) );
  AND2_X1 U7561 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n6378) );
  INV_X1 U7562 ( .A(n8005), .ZN(n6380) );
  NAND2_X1 U7563 ( .A1(n6380), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8189) );
  INV_X1 U7564 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10309) );
  INV_X1 U7565 ( .A(n8202), .ZN(n6381) );
  NAND2_X1 U7566 ( .A1(n6381), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n8214) );
  INV_X1 U7567 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8567) );
  INV_X1 U7568 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n10292) );
  INV_X1 U7569 ( .A(n7987), .ZN(n8794) );
  AND2_X2 U7570 ( .A1(n6383), .A2(n6382), .ZN(n6516) );
  INV_X1 U7571 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6386) );
  NAND2_X1 U7572 ( .A1(n8218), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6385) );
  NAND2_X1 U7573 ( .A1(n8219), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6384) );
  OAI211_X1 U7574 ( .C1(n8223), .C2(n6386), .A(n6385), .B(n6384), .ZN(n6387)
         );
  AOI21_X1 U7575 ( .B1(n8794), .B2(n8191), .A(n6387), .ZN(n8809) );
  NAND2_X1 U7576 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n8708), .ZN(n6388) );
  OAI21_X1 U7577 ( .B1(n8809), .B2(n8708), .A(n6388), .ZN(P2_U3581) );
  INV_X1 U7578 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6390) );
  MUX2_X1 U7579 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n6390), .S(n7411), .Z(n6391)
         );
  INV_X1 U7580 ( .A(n6391), .ZN(n6392) );
  NOR2_X1 U7581 ( .A1(n6393), .A2(n6392), .ZN(n6457) );
  AOI211_X1 U7582 ( .C1(n6393), .C2(n6392), .A(n6457), .B(n10607), .ZN(n6403)
         );
  INV_X1 U7583 ( .A(n7411), .ZN(n6461) );
  NOR2_X1 U7584 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10080), .ZN(n6394) );
  AOI21_X1 U7585 ( .B1(n10606), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n6394), .ZN(
        n6401) );
  OAI21_X1 U7586 ( .B1(n6396), .B2(n6290), .A(n6395), .ZN(n6399) );
  INV_X1 U7587 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6397) );
  MUX2_X1 U7588 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n6397), .S(n7411), .Z(n6398)
         );
  NAND2_X1 U7589 ( .A1(n6398), .A2(n6399), .ZN(n6460) );
  OAI211_X1 U7590 ( .C1(n6399), .C2(n6398), .A(n10615), .B(n6460), .ZN(n6400)
         );
  OAI211_X1 U7591 ( .C1(n10585), .C2(n6461), .A(n6401), .B(n6400), .ZN(n6402)
         );
  OR2_X1 U7592 ( .A1(n6403), .A2(n6402), .ZN(P2_U3255) );
  MUX2_X1 U7593 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n5713), .Z(n6406) );
  NAND2_X1 U7594 ( .A1(n6406), .A2(SI_15_), .ZN(n6441) );
  INV_X1 U7595 ( .A(n6406), .ZN(n6407) );
  NAND2_X1 U7596 ( .A1(n6407), .A2(n10252), .ZN(n6408) );
  OR2_X1 U7597 ( .A1(n6410), .A2(n6409), .ZN(n6411) );
  NAND2_X1 U7598 ( .A1(n6442), .A2(n6411), .ZN(n8085) );
  INV_X1 U7599 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n10401) );
  NAND3_X1 U7600 ( .A1(n10396), .A2(n10397), .A3(n10401), .ZN(n6412) );
  NAND2_X1 U7601 ( .A1(n6454), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6414) );
  XNOR2_X1 U7602 ( .A(n6414), .B(P1_IR_REG_15__SCAN_IN), .ZN(n7756) );
  INV_X1 U7603 ( .A(n7756), .ZN(n7125) );
  INV_X1 U7604 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6415) );
  OAI222_X1 U7605 ( .A1(n10451), .A2(n8085), .B1(n7125), .B2(P1_U3084), .C1(
        n6415), .C2(n10455), .ZN(P1_U3338) );
  NAND2_X1 U7606 ( .A1(n6416), .A2(n6444), .ZN(n6417) );
  NAND2_X1 U7607 ( .A1(n6417), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6418) );
  XNOR2_X1 U7608 ( .A(n6418), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8086) );
  INV_X1 U7609 ( .A(n8086), .ZN(n7837) );
  INV_X1 U7610 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6419) );
  OAI222_X1 U7611 ( .A1(P2_U3152), .A2(n7837), .B1(n9153), .B2(n8085), .C1(
        n6419), .C2(n9151), .ZN(P2_U3343) );
  NOR2_X1 U7612 ( .A1(n7751), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6420) );
  AOI21_X1 U7613 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n7751), .A(n6420), .ZN(
        n6423) );
  AOI21_X1 U7614 ( .B1(n7721), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6421), .ZN(
        n6422) );
  NAND2_X1 U7615 ( .A1(n6423), .A2(n6422), .ZN(n7118) );
  OAI21_X1 U7616 ( .B1(n6423), .B2(n6422), .A(n7118), .ZN(n6424) );
  INV_X1 U7617 ( .A(n6424), .ZN(n6434) );
  INV_X1 U7618 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10856) );
  AOI22_X1 U7619 ( .A1(n7751), .A2(P1_REG1_REG_14__SCAN_IN), .B1(n10856), .B2(
        n6425), .ZN(n6428) );
  OAI21_X1 U7620 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n7721), .A(n6426), .ZN(
        n6427) );
  NAND2_X1 U7621 ( .A1(n6428), .A2(n6427), .ZN(n7122) );
  OAI21_X1 U7622 ( .B1(n6428), .B2(n6427), .A(n7122), .ZN(n6432) );
  INV_X1 U7623 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7620) );
  NOR2_X1 U7624 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6429), .ZN(n9262) );
  AOI21_X1 U7625 ( .B1(n10566), .B2(n7751), .A(n9262), .ZN(n6430) );
  OAI21_X1 U7626 ( .B1(n7620), .B2(n10626), .A(n6430), .ZN(n6431) );
  AOI21_X1 U7627 ( .B1(n6432), .B2(n10573), .A(n6431), .ZN(n6433) );
  OAI21_X1 U7628 ( .B1(n6434), .B2(n7688), .A(n6433), .ZN(P1_U3255) );
  NAND2_X1 U7629 ( .A1(n6031), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6439) );
  NAND2_X1 U7630 ( .A1(n8407), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8421) );
  INV_X1 U7631 ( .A(n8421), .ZN(n6435) );
  NAND2_X1 U7632 ( .A1(n6435), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8429) );
  INV_X1 U7633 ( .A(n8429), .ZN(n8420) );
  NAND2_X1 U7634 ( .A1(n8420), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6602) );
  NAND3_X1 U7635 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .A3(n8445), .ZN(n8448) );
  INV_X1 U7636 ( .A(n8448), .ZN(n9698) );
  NAND2_X1 U7637 ( .A1(n6576), .A2(n9698), .ZN(n6438) );
  NAND2_X1 U7638 ( .A1(n6932), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6437) );
  NAND2_X1 U7639 ( .A1(n9423), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6436) );
  NAND2_X1 U7640 ( .A1(n9674), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6440) );
  OAI21_X1 U7641 ( .B1(n9484), .B2(n9674), .A(n6440), .ZN(P1_U3584) );
  MUX2_X1 U7642 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n7958), .Z(n6589) );
  XNOR2_X1 U7643 ( .A(n6591), .B(n6590), .ZN(n8329) );
  INV_X1 U7644 ( .A(n8329), .ZN(n6456) );
  NOR2_X1 U7645 ( .A1(n6451), .A2(n9146), .ZN(n6448) );
  MUX2_X1 U7646 ( .A(n9146), .B(n6448), .S(P2_IR_REG_16__SCAN_IN), .Z(n6449)
         );
  INV_X1 U7647 ( .A(n6449), .ZN(n6452) );
  NAND2_X1 U7648 ( .A1(n6451), .A2(n6450), .ZN(n6482) );
  AND2_X1 U7649 ( .A1(n6452), .A2(n6482), .ZN(n8092) );
  AOI22_X1 U7650 ( .A1(n8092), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n9149), .ZN(n6453) );
  OAI21_X1 U7651 ( .B1(n6456), .B2(n9153), .A(n6453), .ZN(P2_U3342) );
  OAI21_X1 U7652 ( .B1(n6454), .B2(P1_IR_REG_15__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6596) );
  XNOR2_X1 U7653 ( .A(n6596), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8330) );
  AOI22_X1 U7654 ( .A1(n8330), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n10445), .ZN(n6455) );
  OAI21_X1 U7655 ( .B1(n6456), .B2(n10451), .A(n6455), .ZN(P1_U3337) );
  INV_X1 U7656 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7421) );
  MUX2_X1 U7657 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n7421), .S(n7535), .Z(n6459)
         );
  AOI21_X1 U7658 ( .B1(n7411), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6457), .ZN(
        n6458) );
  NAND2_X1 U7659 ( .A1(n6458), .A2(n6459), .ZN(n7064) );
  OAI21_X1 U7660 ( .B1(n6459), .B2(n6458), .A(n7064), .ZN(n6468) );
  INV_X1 U7661 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7538) );
  NOR2_X1 U7662 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7538), .ZN(n7548) );
  AOI21_X1 U7663 ( .B1(n10606), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7548), .ZN(
        n6466) );
  OAI21_X1 U7664 ( .B1(n6461), .B2(n6397), .A(n6460), .ZN(n6464) );
  INV_X1 U7665 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6462) );
  MUX2_X1 U7666 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n6462), .S(n7535), .Z(n6463)
         );
  NAND2_X1 U7667 ( .A1(n6463), .A2(n6464), .ZN(n7056) );
  OAI211_X1 U7668 ( .C1(n6464), .C2(n6463), .A(n10615), .B(n7056), .ZN(n6465)
         );
  OAI211_X1 U7669 ( .C1(n10585), .C2(n7057), .A(n6466), .B(n6465), .ZN(n6467)
         );
  AOI21_X1 U7670 ( .B1(n10584), .B2(n6468), .A(n6467), .ZN(n6469) );
  INV_X1 U7671 ( .A(n6469), .ZN(P2_U3256) );
  NOR4_X1 U7672 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6473) );
  NOR4_X1 U7673 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6472) );
  NOR4_X1 U7674 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6471) );
  NOR4_X1 U7675 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6470) );
  NAND4_X1 U7676 ( .A1(n6473), .A2(n6472), .A3(n6471), .A4(n6470), .ZN(n6481)
         );
  NOR2_X1 U7677 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6477) );
  NOR4_X1 U7678 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6476) );
  NOR4_X1 U7679 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6475) );
  NOR4_X1 U7680 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6474) );
  NAND4_X1 U7681 ( .A1(n6477), .A2(n6476), .A3(n6475), .A4(n6474), .ZN(n6480)
         );
  INV_X1 U7682 ( .A(P2_B_REG_SCAN_IN), .ZN(n6478) );
  OAI21_X1 U7683 ( .B1(n6481), .B2(n6480), .A(n10461), .ZN(n6608) );
  NAND2_X1 U7684 ( .A1(n7037), .A2(n6483), .ZN(n6484) );
  NAND2_X1 U7685 ( .A1(n6513), .A2(n6499), .ZN(n6615) );
  NAND2_X1 U7686 ( .A1(n6490), .A2(n6489), .ZN(n6491) );
  NAND4_X1 U7687 ( .A1(n6608), .A2(P2_STATE_REG_SCAN_IN), .A3(n6771), .A4(
        n6690), .ZN(n6493) );
  INV_X1 U7688 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10463) );
  NAND2_X1 U7689 ( .A1(n7702), .A2(n7929), .ZN(n10579) );
  NOR2_X1 U7690 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n6494), .ZN(n6495) );
  NAND2_X1 U7691 ( .A1(n6496), .A2(n6495), .ZN(n6497) );
  INV_X1 U7692 ( .A(n6687), .ZN(n6498) );
  INV_X1 U7693 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6529) );
  NAND2_X1 U7694 ( .A1(n6499), .A2(n8324), .ZN(n6753) );
  OAI22_X1 U7695 ( .A1(n6615), .A2(n6522), .B1(n8547), .B2(n6753), .ZN(n6500)
         );
  INV_X1 U7696 ( .A(n6718), .ZN(n6501) );
  NAND2_X1 U7697 ( .A1(n6501), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6504) );
  NAND2_X1 U7698 ( .A1(n6719), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6503) );
  NAND2_X1 U7699 ( .A1(n6516), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6502) );
  NAND4_X1 U7700 ( .A1(n6505), .A2(n6504), .A3(n6503), .A4(n6502), .ZN(n6514)
         );
  NAND2_X1 U7701 ( .A1(n7966), .A2(SI_0_), .ZN(n6506) );
  XNOR2_X1 U7702 ( .A(n6506), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9155) );
  MUX2_X1 U7703 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9155), .S(n6729), .Z(n6756) );
  INV_X1 U7704 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6826) );
  NAND2_X1 U7705 ( .A1(n6516), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6507) );
  NAND4_X2 U7706 ( .A1(n6510), .A2(n6509), .A3(n6508), .A4(n6507), .ZN(n8707)
         );
  NAND2_X1 U7707 ( .A1(n6839), .A2(n6759), .ZN(n8025) );
  NAND2_X1 U7708 ( .A1(n8707), .A2(n6832), .ZN(n8024) );
  NAND2_X1 U7709 ( .A1(n8025), .A2(n8024), .ZN(n6515) );
  XNOR2_X1 U7710 ( .A(n6698), .B(n6515), .ZN(n6829) );
  INV_X1 U7711 ( .A(n6513), .ZN(n8248) );
  OR2_X1 U7712 ( .A1(n6499), .A2(n8252), .ZN(n8246) );
  NAND2_X1 U7713 ( .A1(n6780), .A2(n6756), .ZN(n6731) );
  XNOR2_X1 U7714 ( .A(n6515), .B(n6731), .ZN(n6524) );
  AOI21_X1 U7715 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n6719), .A(n6517), .ZN(
        n6521) );
  INV_X1 U7716 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6518) );
  OR2_X1 U7717 ( .A1(n6707), .A2(n6518), .ZN(n6519) );
  INV_X1 U7718 ( .A(n6756), .ZN(n10639) );
  NAND2_X1 U7719 ( .A1(n6759), .A2(n6756), .ZN(n6525) );
  AND2_X1 U7720 ( .A1(n6873), .A2(n6525), .ZN(n6824) );
  AOI22_X1 U7721 ( .A1(n6824), .A2(n10792), .B1(n9124), .B2(n6759), .ZN(n6527)
         );
  OAI211_X1 U7722 ( .C1(n10841), .C2(n6829), .A(n6835), .B(n6527), .ZN(n6531)
         );
  NAND2_X1 U7723 ( .A1(n6531), .A2(n10873), .ZN(n6528) );
  OAI21_X1 U7724 ( .B1(n10873), .B2(n6529), .A(n6528), .ZN(P2_U3454) );
  INV_X1 U7725 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6533) );
  NAND2_X1 U7726 ( .A1(n6531), .A2(n10870), .ZN(n6532) );
  OAI21_X1 U7727 ( .B1(n10870), .B2(n6533), .A(n6532), .ZN(P2_U3521) );
  OR2_X1 U7728 ( .A1(n6725), .A2(n6231), .ZN(n6535) );
  INV_X4 U7729 ( .A(n6149), .ZN(n8442) );
  NAND2_X1 U7730 ( .A1(n8442), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n6534) );
  OAI211_X1 U7731 ( .C1(n6537), .C2(n6536), .A(n6535), .B(n6534), .ZN(n6860)
         );
  OAI22_X1 U7732 ( .A1(n7046), .A2(n9287), .B1(n7003), .B2(n9289), .ZN(n6538)
         );
  XNOR2_X1 U7733 ( .A(n6538), .B(n9243), .ZN(n6564) );
  OR2_X1 U7734 ( .A1(n7046), .A2(n9286), .ZN(n6540) );
  NAND2_X1 U7735 ( .A1(n6860), .A2(n9198), .ZN(n6539) );
  NAND2_X1 U7736 ( .A1(n6540), .A2(n6539), .ZN(n6563) );
  XNOR2_X1 U7737 ( .A(n6564), .B(n6563), .ZN(n6549) );
  INV_X1 U7738 ( .A(n6541), .ZN(n6542) );
  NAND2_X1 U7739 ( .A1(n6543), .A2(n6542), .ZN(n6544) );
  INV_X1 U7740 ( .A(n6566), .ZN(n6547) );
  AOI211_X1 U7741 ( .C1(n6549), .C2(n6548), .A(n9410), .B(n6547), .ZN(n6562)
         );
  INV_X1 U7742 ( .A(n6550), .ZN(n6679) );
  OAI22_X1 U7743 ( .A1(n6671), .A2(n9402), .B1(n9401), .B2(n6679), .ZN(n6561)
         );
  NAND2_X1 U7744 ( .A1(n6031), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6556) );
  AOI21_X1 U7745 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6551) );
  NOR2_X1 U7746 ( .A1(n6551), .A2(n6578), .ZN(n7074) );
  NAND2_X1 U7747 ( .A1(n6931), .A2(n7074), .ZN(n6555) );
  NAND2_X1 U7748 ( .A1(n6933), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6554) );
  NAND2_X1 U7749 ( .A1(n6552), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6553) );
  NAND4_X1 U7750 ( .A1(n6556), .A2(n6555), .A3(n6554), .A4(n6553), .ZN(n9673)
         );
  INV_X1 U7751 ( .A(n6557), .ZN(n6558) );
  AOI21_X1 U7752 ( .B1(n9406), .B2(n9673), .A(n6558), .ZN(n6559) );
  OAI21_X1 U7753 ( .B1(n9384), .B2(n7003), .A(n6559), .ZN(n6560) );
  OR3_X1 U7754 ( .A1(n6562), .A2(n6561), .A3(n6560), .ZN(P1_U3228) );
  NAND2_X1 U7755 ( .A1(n6564), .A2(n6563), .ZN(n6565) );
  NAND2_X1 U7756 ( .A1(n9673), .A2(n9198), .ZN(n6571) );
  OR2_X1 U7757 ( .A1(n6945), .A2(n6231), .ZN(n6569) );
  AOI22_X1 U7758 ( .A1(n8442), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n8352), .B2(
        n6567), .ZN(n6568) );
  NAND2_X1 U7759 ( .A1(n6571), .A2(n6570), .ZN(n6572) );
  XNOR2_X1 U7760 ( .A(n6572), .B(n9243), .ZN(n6643) );
  NAND2_X1 U7761 ( .A1(n9673), .A2(n9239), .ZN(n6574) );
  NAND2_X1 U7762 ( .A1(n7077), .A2(n9198), .ZN(n6573) );
  NAND2_X1 U7763 ( .A1(n6574), .A2(n6573), .ZN(n6642) );
  INV_X1 U7764 ( .A(n6642), .ZN(n6640) );
  XNOR2_X1 U7765 ( .A(n6643), .B(n6640), .ZN(n6575) );
  XNOR2_X1 U7766 ( .A(n6646), .B(n6575), .ZN(n6588) );
  INV_X1 U7767 ( .A(n9402), .ZN(n9381) );
  AOI22_X1 U7768 ( .A1(n9381), .A2(n6669), .B1(n9347), .B2(n7074), .ZN(n6587)
         );
  OAI21_X1 U7769 ( .B1(n6578), .B2(P1_REG3_REG_6__SCAN_IN), .A(n6577), .ZN(
        n6579) );
  INV_X1 U7770 ( .A(n6579), .ZN(n7031) );
  NAND2_X1 U7771 ( .A1(n6931), .A2(n7031), .ZN(n6583) );
  NAND2_X1 U7772 ( .A1(n6031), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6582) );
  NAND2_X1 U7773 ( .A1(n6933), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6581) );
  NAND2_X1 U7774 ( .A1(n9423), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6580) );
  NOR2_X1 U7775 ( .A1(n9388), .A2(n7047), .ZN(n6584) );
  AOI211_X1 U7776 ( .C1(n7077), .C2(n9407), .A(n6585), .B(n6584), .ZN(n6586)
         );
  OAI211_X1 U7777 ( .C1(n6588), .C2(n9410), .A(n6587), .B(n6586), .ZN(P1_U3225) );
  MUX2_X1 U7778 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n7958), .Z(n6592) );
  NAND2_X1 U7779 ( .A1(n6592), .A2(SI_17_), .ZN(n6984) );
  OAI21_X1 U7780 ( .B1(n6592), .B2(SI_17_), .A(n6984), .ZN(n6593) );
  NAND2_X1 U7781 ( .A1(n6594), .A2(n6593), .ZN(n6595) );
  NAND2_X1 U7782 ( .A1(n6595), .A2(n6985), .ZN(n8334) );
  INV_X1 U7783 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n10405) );
  NAND2_X1 U7784 ( .A1(n6596), .A2(n10405), .ZN(n6597) );
  NAND2_X1 U7785 ( .A1(n6597), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6599) );
  NAND2_X1 U7786 ( .A1(n6599), .A2(n6598), .ZN(n6987) );
  OR2_X1 U7787 ( .A1(n6599), .A2(n6598), .ZN(n6600) );
  AOI22_X1 U7788 ( .A1(n8335), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10445), .ZN(n6601) );
  OAI21_X1 U7789 ( .B1(n8334), .B2(n10451), .A(n6601), .ZN(P1_U3336) );
  INV_X1 U7790 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7944) );
  XNOR2_X1 U7791 ( .A(P1_REG3_REG_27__SCAN_IN), .B(n6602), .ZN(n9715) );
  NAND2_X1 U7792 ( .A1(n6931), .A2(n9715), .ZN(n6606) );
  NAND2_X1 U7793 ( .A1(n6031), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6605) );
  NAND2_X1 U7794 ( .A1(n6932), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6604) );
  NAND2_X1 U7795 ( .A1(n9423), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6603) );
  INV_X1 U7796 ( .A(n9723), .ZN(n8440) );
  NAND2_X1 U7797 ( .A1(n8440), .A2(P1_U4006), .ZN(n6607) );
  OAI21_X1 U7798 ( .B1(n7944), .B2(P1_U4006), .A(n6607), .ZN(P1_U3582) );
  NAND2_X1 U7799 ( .A1(n6771), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6689) );
  INV_X1 U7800 ( .A(n6689), .ZN(n6611) );
  NAND2_X1 U7801 ( .A1(n6609), .A2(n6608), .ZN(n6688) );
  INV_X1 U7802 ( .A(n6688), .ZN(n6610) );
  INV_X1 U7803 ( .A(n6613), .ZN(n6616) );
  NAND2_X1 U7804 ( .A1(n6690), .A2(n6616), .ZN(n6770) );
  NAND2_X1 U7805 ( .A1(n6611), .A2(n6770), .ZN(n6842) );
  INV_X1 U7806 ( .A(n10462), .ZN(n6691) );
  NAND2_X1 U7807 ( .A1(n6691), .A2(n6613), .ZN(n6612) );
  NAND2_X1 U7808 ( .A1(n8676), .A2(n9014), .ZN(n8555) );
  NOR2_X1 U7809 ( .A1(n8547), .A2(n6613), .ZN(n6614) );
  OAI22_X1 U7810 ( .A1(n6839), .A2(n8555), .B1(n8693), .B2(n10639), .ZN(n6621)
         );
  MUX2_X1 U7811 ( .A(n8023), .B(n10639), .S(n6757), .Z(n6619) );
  NOR2_X1 U7812 ( .A1(n6617), .A2(n6616), .ZN(n6618) );
  AOI21_X1 U7813 ( .B1(n6619), .B2(n6731), .A(n8667), .ZN(n6620) );
  AOI211_X1 U7814 ( .C1(P2_REG3_REG_0__SCAN_IN), .C2(n6842), .A(n6621), .B(
        n6620), .ZN(n6622) );
  INV_X1 U7815 ( .A(n6622), .ZN(P2_U3234) );
  NAND3_X1 U7816 ( .A1(n6625), .A2(n6624), .A3(n6623), .ZN(n7015) );
  NOR2_X1 U7817 ( .A1(n6626), .A2(n9812), .ZN(n6627) );
  INV_X1 U7818 ( .A(n6628), .ZN(n6629) );
  AND2_X1 U7819 ( .A1(n6630), .A2(n9659), .ZN(n6631) );
  NAND2_X1 U7820 ( .A1(n10772), .A2(n6632), .ZN(n6635) );
  OAI22_X1 U7821 ( .A1(n10783), .A2(n5831), .B1(n10638), .B2(n9897), .ZN(n6633) );
  INV_X1 U7822 ( .A(n6633), .ZN(n6634) );
  OAI211_X1 U7823 ( .C1(n6160), .C2(n10780), .A(n6635), .B(n6634), .ZN(n6636)
         );
  AOI21_X1 U7824 ( .B1(n10773), .B2(n6637), .A(n6636), .ZN(n6638) );
  OAI21_X1 U7825 ( .B1(n6639), .B2(n10778), .A(n6638), .ZN(P1_U3289) );
  INV_X1 U7826 ( .A(n6643), .ZN(n6641) );
  NAND2_X1 U7827 ( .A1(n6641), .A2(n6640), .ZN(n6645) );
  AND2_X1 U7828 ( .A1(n6643), .A2(n6642), .ZN(n6644) );
  AOI21_X2 U7829 ( .B1(n6646), .B2(n6645), .A(n6644), .ZN(n6921) );
  OR2_X1 U7830 ( .A1(n7089), .A2(n6231), .ZN(n6648) );
  AOI22_X1 U7831 ( .A1(n8442), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n8352), .B2(
        n10513), .ZN(n6647) );
  NAND2_X1 U7832 ( .A1(n6648), .A2(n6647), .ZN(n7164) );
  OR2_X1 U7833 ( .A1(n7047), .A2(n9287), .ZN(n6649) );
  NAND2_X1 U7834 ( .A1(n6650), .A2(n6649), .ZN(n6652) );
  XNOR2_X1 U7835 ( .A(n6652), .B(n9243), .ZN(n6655) );
  NAND2_X1 U7836 ( .A1(n7164), .A2(n9198), .ZN(n6654) );
  OR2_X1 U7837 ( .A1(n7047), .A2(n9286), .ZN(n6653) );
  NAND2_X1 U7838 ( .A1(n6654), .A2(n6653), .ZN(n6656) );
  NAND2_X1 U7839 ( .A1(n6655), .A2(n6656), .ZN(n6920) );
  INV_X1 U7840 ( .A(n6655), .ZN(n6658) );
  INV_X1 U7841 ( .A(n6656), .ZN(n6657) );
  NAND2_X1 U7842 ( .A1(n6658), .A2(n6657), .ZN(n6922) );
  NAND2_X1 U7843 ( .A1(n6920), .A2(n6922), .ZN(n6659) );
  XNOR2_X1 U7844 ( .A(n6921), .B(n6659), .ZN(n6664) );
  AOI22_X1 U7845 ( .A1(n9381), .A2(n9673), .B1(n9347), .B2(n7031), .ZN(n6663)
         );
  NAND2_X1 U7846 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10523) );
  INV_X1 U7847 ( .A(n10523), .ZN(n6661) );
  NOR2_X1 U7848 ( .A1(n9388), .A2(n7198), .ZN(n6660) );
  AOI211_X1 U7849 ( .C1(n7164), .C2(n9407), .A(n6661), .B(n6660), .ZN(n6662)
         );
  OAI211_X1 U7850 ( .C1(n6664), .C2(n9410), .A(n6663), .B(n6662), .ZN(P1_U3237) );
  NAND2_X1 U7851 ( .A1(n6849), .A2(n6160), .ZN(n6665) );
  NAND2_X1 U7852 ( .A1(n6671), .A2(n6813), .ZN(n9451) );
  NAND2_X1 U7853 ( .A1(n9451), .A2(n9453), .ZN(n9625) );
  NAND2_X1 U7854 ( .A1(n6804), .A2(n9625), .ZN(n6803) );
  NAND2_X1 U7855 ( .A1(n6671), .A2(n10662), .ZN(n6668) );
  NAND2_X1 U7856 ( .A1(n6803), .A2(n6668), .ZN(n6670) );
  NAND2_X1 U7857 ( .A1(n7046), .A2(n6860), .ZN(n9456) );
  NAND2_X1 U7858 ( .A1(n6669), .A2(n7003), .ZN(n9454) );
  NAND2_X1 U7859 ( .A1(n9456), .A2(n9454), .ZN(n6674) );
  OAI21_X1 U7860 ( .B1(n6670), .B2(n6674), .A(n7005), .ZN(n6859) );
  INV_X1 U7861 ( .A(n9673), .ZN(n7002) );
  OAI22_X1 U7862 ( .A1(n7002), .A2(n10753), .B1(n6671), .B2(n10755), .ZN(n6677) );
  INV_X1 U7863 ( .A(n9451), .ZN(n6673) );
  INV_X1 U7864 ( .A(n6674), .ZN(n9631) );
  XNOR2_X1 U7865 ( .A(n7001), .B(n9631), .ZN(n6675) );
  NOR2_X1 U7866 ( .A1(n6675), .A2(n9888), .ZN(n6676) );
  AOI211_X1 U7867 ( .C1(n10822), .C2(n6859), .A(n6677), .B(n6676), .ZN(n6863)
         );
  NAND2_X1 U7868 ( .A1(n6678), .A2(n10662), .ZN(n6810) );
  AOI21_X1 U7869 ( .B1(n6860), .B2(n6810), .A(n5351), .ZN(n6861) );
  NOR2_X1 U7870 ( .A1(n10780), .A2(n7003), .ZN(n6682) );
  OAI22_X1 U7871 ( .A1(n10783), .A2(n6680), .B1(n6679), .B2(n9897), .ZN(n6681)
         );
  AOI211_X1 U7872 ( .C1(n6861), .C2(n10772), .A(n6682), .B(n6681), .ZN(n6684)
         );
  NAND2_X1 U7873 ( .A1(n6859), .A2(n10773), .ZN(n6683) );
  OAI211_X1 U7874 ( .C1(n6863), .C2(n10778), .A(n6684), .B(n6683), .ZN(
        P1_U3287) );
  NAND2_X1 U7875 ( .A1(n6482), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6685) );
  XNOR2_X1 U7876 ( .A(n6685), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8720) );
  INV_X1 U7877 ( .A(n8720), .ZN(n8711) );
  INV_X1 U7878 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6686) );
  OAI222_X1 U7879 ( .A1(P2_U3152), .A2(n8711), .B1(n9153), .B2(n8334), .C1(
        n6686), .C2(n9151), .ZN(P2_U3341) );
  AND2_X1 U7880 ( .A1(n6731), .A2(n8023), .ZN(n10641) );
  INV_X1 U7881 ( .A(n6690), .ZN(n6692) );
  OR2_X1 U7882 ( .A1(n8251), .A2(n8314), .ZN(n6872) );
  NAND2_X1 U7883 ( .A1(n8979), .A2(n6872), .ZN(n10809) );
  INV_X1 U7884 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6694) );
  INV_X1 U7885 ( .A(n9014), .ZN(n8808) );
  OAI22_X1 U7886 ( .A1(n10641), .A2(n10797), .B1(n6839), .B2(n8808), .ZN(
        n10643) );
  AOI21_X1 U7887 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n10801), .A(n10643), .ZN(
        n6693) );
  MUX2_X1 U7888 ( .A(n6694), .B(n6693), .S(n10811), .Z(n6697) );
  NOR2_X1 U7889 ( .A1(n8547), .A2(n10640), .ZN(n10803) );
  OAI21_X1 U7890 ( .B1(n9035), .B2(n9020), .A(n6756), .ZN(n6696) );
  OAI211_X1 U7891 ( .C1(n10641), .C2(n9022), .A(n6697), .B(n6696), .ZN(
        P2_U3296) );
  OAI21_X1 U7892 ( .B1(n8707), .B2(n6759), .A(n6698), .ZN(n6700) );
  NAND2_X1 U7893 ( .A1(n8707), .A2(n6759), .ZN(n6699) );
  AND2_X1 U7894 ( .A1(n6700), .A2(n6699), .ZN(n6870) );
  NAND2_X1 U7895 ( .A1(n6791), .A2(n10656), .ZN(n6705) );
  NAND2_X1 U7896 ( .A1(n6871), .A2(n6705), .ZN(n6786) );
  NAND2_X1 U7897 ( .A1(n8192), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6712) );
  NAND2_X1 U7898 ( .A1(n6516), .A2(n10082), .ZN(n6711) );
  INV_X1 U7899 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6706) );
  OR2_X1 U7900 ( .A1(n6707), .A2(n6706), .ZN(n6710) );
  OR2_X1 U7901 ( .A1(n6718), .A2(n6708), .ZN(n6709) );
  NAND4_X2 U7902 ( .A1(n6712), .A2(n6711), .A3(n6710), .A4(n6709), .ZN(n8706)
         );
  OR2_X1 U7903 ( .A1(n6946), .A2(n5199), .ZN(n6717) );
  OR2_X1 U7904 ( .A1(n6702), .A2(n6713), .ZN(n6716) );
  INV_X2 U7905 ( .A(n6729), .ZN(n8134) );
  NAND2_X1 U7906 ( .A1(n8134), .A2(n6714), .ZN(n6715) );
  XNOR2_X1 U7907 ( .A(n8706), .B(n6795), .ZN(n8262) );
  NAND2_X1 U7908 ( .A1(n6786), .A2(n8262), .ZN(n6785) );
  INV_X1 U7909 ( .A(n8706), .ZN(n6910) );
  NAND2_X1 U7910 ( .A1(n6910), .A2(n6795), .ZN(n8030) );
  INV_X1 U7911 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6720) );
  OR2_X1 U7912 ( .A1(n8169), .A2(n6720), .ZN(n6721) );
  OAI21_X1 U7913 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n6737), .ZN(n6911) );
  OR2_X1 U7914 ( .A1(n6946), .A2(n5894), .ZN(n6727) );
  OR2_X1 U7915 ( .A1(n6702), .A2(n6725), .ZN(n6726) );
  OAI211_X1 U7916 ( .C1(n6729), .C2(n6728), .A(n6727), .B(n6726), .ZN(n6914)
         );
  NAND2_X1 U7917 ( .A1(n6961), .A2(n6914), .ZN(n8038) );
  NAND2_X1 U7918 ( .A1(n8705), .A2(n5317), .ZN(n6964) );
  OAI21_X1 U7919 ( .B1(n6730), .B2(n8259), .A(n6944), .ZN(n10673) );
  INV_X1 U7920 ( .A(n10673), .ZN(n6752) );
  NAND2_X1 U7921 ( .A1(n6731), .A2(n8025), .ZN(n8261) );
  NAND2_X1 U7922 ( .A1(n6881), .A2(n8028), .ZN(n6790) );
  INV_X1 U7923 ( .A(n8262), .ZN(n6789) );
  INV_X1 U7924 ( .A(n6788), .ZN(n6733) );
  NOR2_X1 U7925 ( .A1(n8706), .A2(n6795), .ZN(n6734) );
  OAI21_X1 U7926 ( .B1(n6733), .B2(n6734), .A(n8259), .ZN(n6736) );
  NOR2_X1 U7927 ( .A1(n8259), .A2(n6734), .ZN(n6735) );
  NAND3_X1 U7928 ( .A1(n6736), .A2(n7131), .A3(n9017), .ZN(n6746) );
  NAND2_X1 U7929 ( .A1(n8192), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6744) );
  NAND2_X1 U7930 ( .A1(n6737), .A2(n10096), .ZN(n6738) );
  AND2_X1 U7931 ( .A1(n6952), .A2(n6738), .ZN(n6992) );
  NAND2_X1 U7932 ( .A1(n6516), .A2(n6992), .ZN(n6743) );
  INV_X1 U7933 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6739) );
  OR2_X1 U7934 ( .A1(n8169), .A2(n6739), .ZN(n6742) );
  INV_X1 U7935 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6740) );
  OR2_X1 U7936 ( .A1(n8171), .A2(n6740), .ZN(n6741) );
  NAND4_X2 U7937 ( .A1(n6744), .A2(n6743), .A3(n6742), .A4(n6741), .ZN(n8704)
         );
  AOI22_X1 U7938 ( .A1(n9012), .A2(n8706), .B1(n8704), .B2(n9014), .ZN(n6745)
         );
  NAND2_X1 U7939 ( .A1(n6746), .A2(n6745), .ZN(n10671) );
  INV_X1 U7940 ( .A(n10671), .ZN(n6747) );
  MUX2_X1 U7941 ( .A(n6266), .B(n6747), .S(n10811), .Z(n6751) );
  NAND2_X1 U7942 ( .A1(n6797), .A2(n6914), .ZN(n6748) );
  NAND2_X1 U7943 ( .A1(n6962), .A2(n6748), .ZN(n10670) );
  OAI22_X1 U7944 ( .A1(n10670), .A2(n8793), .B1(n6911), .B2(n8981), .ZN(n6749)
         );
  AOI21_X1 U7945 ( .B1(n9035), .B2(n6914), .A(n6749), .ZN(n6750) );
  OAI211_X1 U7946 ( .C1(n6752), .C2(n9022), .A(n6751), .B(n6750), .ZN(P2_U3292) );
  INV_X1 U7947 ( .A(n6698), .ZN(n6758) );
  NAND2_X1 U7948 ( .A1(n6753), .A2(n8314), .ZN(n6754) );
  OAI22_X1 U7949 ( .A1(n6758), .A2(n6757), .B1(n6756), .B2(n6764), .ZN(n6779)
         );
  NAND2_X1 U7950 ( .A1(n8707), .A2(n8531), .ZN(n6761) );
  OAI21_X1 U7951 ( .B1(n6761), .B2(n6760), .A(n6762), .ZN(n6778) );
  INV_X1 U7952 ( .A(n6762), .ZN(n6763) );
  XNOR2_X1 U7953 ( .A(n6765), .B(n6888), .ZN(n6767) );
  NAND2_X1 U7954 ( .A1(n6704), .A2(n8531), .ZN(n6766) );
  OAI21_X1 U7955 ( .B1(n6767), .B2(n6766), .A(n6768), .ZN(n6837) );
  INV_X1 U7956 ( .A(n6768), .ZN(n6769) );
  XNOR2_X1 U7957 ( .A(n6765), .B(n6795), .ZN(n6901) );
  NAND2_X1 U7958 ( .A1(n8706), .A2(n8531), .ZN(n6899) );
  XNOR2_X1 U7959 ( .A(n6901), .B(n6899), .ZN(n6902) );
  XNOR2_X1 U7960 ( .A(n6903), .B(n6902), .ZN(n6776) );
  INV_X1 U7961 ( .A(n8693), .ZN(n8651) );
  INV_X1 U7962 ( .A(n6795), .ZN(n8033) );
  OAI22_X1 U7963 ( .A1(n6791), .A2(n8688), .B1(n6961), .B2(n8555), .ZN(n6774)
         );
  NAND2_X1 U7964 ( .A1(n6771), .A2(n6770), .ZN(n6772) );
  MUX2_X1 U7965 ( .A(P2_U3152), .B(n8690), .S(n10082), .Z(n6773) );
  AOI211_X1 U7966 ( .C1(n8651), .C2(n8033), .A(n6774), .B(n6773), .ZN(n6775)
         );
  OAI21_X1 U7967 ( .B1(n6776), .B2(n8667), .A(n6775), .ZN(P2_U3220) );
  AOI21_X1 U7968 ( .B1(n6779), .B2(n6778), .A(n6777), .ZN(n6784) );
  NOR2_X1 U7969 ( .A1(n8693), .A2(n6832), .ZN(n6782) );
  OAI22_X1 U7970 ( .A1(n6780), .A2(n8688), .B1(n6791), .B2(n8555), .ZN(n6781)
         );
  AOI211_X1 U7971 ( .C1(P2_REG3_REG_1__SCAN_IN), .C2(n6842), .A(n6782), .B(
        n6781), .ZN(n6783) );
  OAI21_X1 U7972 ( .B1(n6784), .B2(n8667), .A(n6783), .ZN(P2_U3224) );
  OAI21_X1 U7973 ( .B1(n6786), .B2(n8262), .A(n6785), .ZN(n6787) );
  INV_X1 U7974 ( .A(n6787), .ZN(n6892) );
  OAI21_X1 U7975 ( .B1(n6790), .B2(n6789), .A(n6788), .ZN(n6794) );
  OAI22_X1 U7976 ( .A1(n6791), .A2(n8806), .B1(n6961), .B2(n8808), .ZN(n6793)
         );
  NOR2_X1 U7977 ( .A1(n6892), .A2(n8979), .ZN(n6792) );
  AOI211_X1 U7978 ( .C1(n9017), .C2(n6794), .A(n6793), .B(n6792), .ZN(n6896)
         );
  OR2_X1 U7979 ( .A1(n6875), .A2(n6795), .ZN(n6796) );
  AND2_X1 U7980 ( .A1(n6797), .A2(n6796), .ZN(n6890) );
  AOI22_X1 U7981 ( .A1(n6890), .A2(n10792), .B1(n9124), .B2(n8033), .ZN(n6798)
         );
  OAI211_X1 U7982 ( .C1(n6892), .C2(n10653), .A(n6896), .B(n6798), .ZN(n6800)
         );
  NAND2_X1 U7983 ( .A1(n6800), .A2(n10873), .ZN(n6799) );
  OAI21_X1 U7984 ( .B1(n10873), .B2(n6706), .A(n6799), .ZN(P2_U3460) );
  NAND2_X1 U7985 ( .A1(n6800), .A2(n10870), .ZN(n6801) );
  OAI21_X1 U7986 ( .B1(n10870), .B2(n6802), .A(n6801), .ZN(P2_U3523) );
  OAI21_X1 U7987 ( .B1(n6804), .B2(n9625), .A(n6803), .ZN(n10666) );
  INV_X1 U7988 ( .A(n10666), .ZN(n6816) );
  INV_X1 U7989 ( .A(n10773), .ZN(n9867) );
  XNOR2_X1 U7990 ( .A(n6805), .B(n9625), .ZN(n6808) );
  OAI22_X1 U7991 ( .A1(n6849), .A2(n10755), .B1(n7046), .B2(n10753), .ZN(n6806) );
  AOI21_X1 U7992 ( .B1(n10666), .B2(n10822), .A(n6806), .ZN(n6807) );
  OAI21_X1 U7993 ( .B1(n9888), .B2(n6808), .A(n6807), .ZN(n10664) );
  NAND2_X1 U7994 ( .A1(n10664), .A2(n10783), .ZN(n6815) );
  INV_X1 U7995 ( .A(n10780), .ZN(n9920) );
  OAI22_X1 U7996 ( .A1(n10783), .A2(n5832), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9897), .ZN(n6812) );
  INV_X1 U7997 ( .A(n10772), .ZN(n7800) );
  OR2_X1 U7998 ( .A1(n6678), .A2(n10662), .ZN(n6809) );
  NAND2_X1 U7999 ( .A1(n6810), .A2(n6809), .ZN(n10663) );
  NOR2_X1 U8000 ( .A1(n7800), .A2(n10663), .ZN(n6811) );
  AOI211_X1 U8001 ( .C1(n9920), .C2(n6813), .A(n6812), .B(n6811), .ZN(n6814)
         );
  OAI211_X1 U8002 ( .C1(n6816), .C2(n9867), .A(n6815), .B(n6814), .ZN(P1_U3288) );
  INV_X1 U8003 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6818) );
  OAI21_X1 U8004 ( .B1(n6818), .B2(n9897), .A(n6817), .ZN(n6819) );
  NAND2_X1 U8005 ( .A1(n6819), .A2(n10783), .ZN(n6822) );
  OAI21_X1 U8006 ( .B1(n9920), .B2(n10772), .A(n6820), .ZN(n6821) );
  OAI211_X1 U8007 ( .C1(n6823), .C2(n10783), .A(n6822), .B(n6821), .ZN(
        P1_U3291) );
  INV_X1 U8008 ( .A(n6824), .ZN(n6825) );
  INV_X1 U8009 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10592) );
  OAI22_X1 U8010 ( .A1(n8793), .A2(n6825), .B1(n10592), .B2(n8981), .ZN(n6828)
         );
  NOR2_X1 U8011 ( .A1(n10811), .A2(n6826), .ZN(n6827) );
  NOR2_X1 U8012 ( .A1(n6828), .A2(n6827), .ZN(n6831) );
  OR2_X1 U8013 ( .A1(n6829), .A2(n9022), .ZN(n6830) );
  OAI211_X1 U8014 ( .C1(n6832), .C2(n9008), .A(n6831), .B(n6830), .ZN(n6833)
         );
  INV_X1 U8015 ( .A(n6833), .ZN(n6834) );
  OAI21_X1 U8016 ( .B1(n6835), .B2(n10813), .A(n6834), .ZN(P2_U3295) );
  AOI21_X1 U8017 ( .B1(n6838), .B2(n6837), .A(n6836), .ZN(n6844) );
  NOR2_X1 U8018 ( .A1(n8693), .A2(n10656), .ZN(n6841) );
  OAI22_X1 U8019 ( .A1(n6910), .A2(n8555), .B1(n6839), .B2(n8688), .ZN(n6840)
         );
  AOI211_X1 U8020 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(n6842), .A(n6841), .B(
        n6840), .ZN(n6843) );
  OAI21_X1 U8021 ( .B1(n6844), .B2(n8667), .A(n6843), .ZN(P2_U3239) );
  INV_X1 U8022 ( .A(n6847), .ZN(n9628) );
  XNOR2_X1 U8023 ( .A(n9628), .B(n6845), .ZN(n10646) );
  OAI21_X1 U8024 ( .B1(n6848), .B2(n6847), .A(n6846), .ZN(n6852) );
  OAI22_X1 U8025 ( .A1(n6850), .A2(n10755), .B1(n6849), .B2(n10753), .ZN(n6851) );
  AOI21_X1 U8026 ( .B1(n6852), .B2(n10758), .A(n6851), .ZN(n6853) );
  OAI21_X1 U8027 ( .B1(n10646), .B2(n10718), .A(n6853), .ZN(n10649) );
  OAI211_X1 U8028 ( .C1(n6855), .C2(n10648), .A(n10878), .B(n6854), .ZN(n10647) );
  INV_X1 U8029 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10567) );
  OAI22_X1 U8030 ( .A1(n10647), .A2(n9760), .B1(n10567), .B2(n9897), .ZN(n6856) );
  OAI21_X1 U8031 ( .B1(n10649), .B2(n6856), .A(n10783), .ZN(n6858) );
  AOI22_X1 U8032 ( .A1(n9920), .A2(n9444), .B1(n10778), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n6857) );
  OAI211_X1 U8033 ( .C1(n10646), .C2(n9867), .A(n6858), .B(n6857), .ZN(
        P1_U3290) );
  INV_X1 U8034 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6866) );
  INV_X1 U8035 ( .A(n6859), .ZN(n6864) );
  AOI22_X1 U8036 ( .A1(n6861), .A2(n10878), .B1(n10877), .B2(n6860), .ZN(n6862) );
  OAI211_X1 U8037 ( .C1(n6864), .C2(n10817), .A(n6863), .B(n6862), .ZN(n6867)
         );
  NAND2_X1 U8038 ( .A1(n6867), .A2(n5045), .ZN(n6865) );
  OAI21_X1 U8039 ( .B1(n5045), .B2(n6866), .A(n6865), .ZN(P1_U3466) );
  INV_X1 U8040 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6869) );
  NAND2_X1 U8041 ( .A1(n6867), .A2(n10722), .ZN(n6868) );
  OAI21_X1 U8042 ( .B1(n10722), .B2(n6869), .A(n6868), .ZN(P1_U3527) );
  OAI21_X1 U8043 ( .B1(n6870), .B2(n6732), .A(n6871), .ZN(n10659) );
  INV_X1 U8044 ( .A(n10659), .ZN(n6877) );
  AND2_X1 U8045 ( .A1(n6873), .A2(n6888), .ZN(n6874) );
  NOR2_X1 U8046 ( .A1(n6875), .A2(n6874), .ZN(n10654) );
  AOI22_X1 U8047 ( .A1(n9020), .A2(n10654), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n10801), .ZN(n6876) );
  OAI21_X1 U8048 ( .B1(n6877), .B2(n8987), .A(n6876), .ZN(n6887) );
  INV_X1 U8049 ( .A(n8979), .ZN(n6878) );
  NAND2_X1 U8050 ( .A1(n10659), .A2(n6878), .ZN(n6885) );
  AOI22_X1 U8051 ( .A1(n9012), .A2(n8707), .B1(n8706), .B2(n9014), .ZN(n6884)
         );
  NAND2_X1 U8052 ( .A1(n6879), .A2(n6732), .ZN(n6880) );
  NAND2_X1 U8053 ( .A1(n6881), .A2(n6880), .ZN(n6882) );
  NAND2_X1 U8054 ( .A1(n6882), .A2(n9017), .ZN(n6883) );
  NAND3_X1 U8055 ( .A1(n6885), .A2(n6884), .A3(n6883), .ZN(n10657) );
  MUX2_X1 U8056 ( .A(n10657), .B(P2_REG2_REG_2__SCAN_IN), .S(n10813), .Z(n6886) );
  AOI211_X1 U8057 ( .C1(n9035), .C2(n6888), .A(n6887), .B(n6886), .ZN(n6889)
         );
  INV_X1 U8058 ( .A(n6889), .ZN(P2_U3294) );
  AOI22_X1 U8059 ( .A1(n6890), .A2(n9020), .B1(n10801), .B2(n10082), .ZN(n6891) );
  OAI21_X1 U8060 ( .B1(n6708), .B2(n10811), .A(n6891), .ZN(n6894) );
  NOR2_X1 U8061 ( .A1(n6892), .A2(n8987), .ZN(n6893) );
  AOI211_X1 U8062 ( .C1(n9035), .C2(n8033), .A(n6894), .B(n6893), .ZN(n6895)
         );
  OAI21_X1 U8063 ( .B1(n6896), .B2(n10813), .A(n6895), .ZN(P2_U3293) );
  XNOR2_X1 U8064 ( .A(n5317), .B(n6765), .ZN(n6898) );
  NOR2_X1 U8065 ( .A1(n6961), .A2(n6757), .ZN(n6897) );
  NOR2_X1 U8066 ( .A1(n6897), .A2(n6898), .ZN(n6973) );
  AOI21_X1 U8067 ( .B1(n6898), .B2(n6897), .A(n6973), .ZN(n6905) );
  INV_X1 U8068 ( .A(n6899), .ZN(n6900) );
  NAND2_X1 U8069 ( .A1(n6904), .A2(n6905), .ZN(n6975) );
  OAI21_X1 U8070 ( .B1(n6905), .B2(n6904), .A(n6975), .ZN(n6906) );
  NAND2_X1 U8071 ( .A1(n6906), .A2(n8683), .ZN(n6916) );
  NAND2_X1 U8072 ( .A1(n8685), .A2(n8704), .ZN(n6909) );
  INV_X1 U8073 ( .A(n6907), .ZN(n6908) );
  OAI211_X1 U8074 ( .C1(n6910), .C2(n8688), .A(n6909), .B(n6908), .ZN(n6913)
         );
  INV_X1 U8075 ( .A(n8690), .ZN(n8674) );
  NOR2_X1 U8076 ( .A1(n8674), .A2(n6911), .ZN(n6912) );
  AOI211_X1 U8077 ( .C1(n8651), .C2(n6914), .A(n6913), .B(n6912), .ZN(n6915)
         );
  NAND2_X1 U8078 ( .A1(n6916), .A2(n6915), .ZN(P2_U3232) );
  NAND2_X1 U8079 ( .A1(n7226), .A2(n9427), .ZN(n6919) );
  AOI22_X1 U8080 ( .A1(n8442), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n8352), .B2(
        n6917), .ZN(n6918) );
  NAND2_X1 U8081 ( .A1(n6919), .A2(n6918), .ZN(n7206) );
  INV_X1 U8082 ( .A(n7206), .ZN(n10685) );
  NAND2_X1 U8083 ( .A1(n6921), .A2(n6920), .ZN(n6923) );
  NAND2_X1 U8084 ( .A1(n6923), .A2(n6922), .ZN(n7175) );
  OR2_X1 U8085 ( .A1(n7198), .A2(n9287), .ZN(n6924) );
  NAND2_X1 U8086 ( .A1(n6925), .A2(n6924), .ZN(n6926) );
  XNOR2_X1 U8087 ( .A(n6926), .B(n9243), .ZN(n7176) );
  NOR2_X1 U8088 ( .A1(n7198), .A2(n9286), .ZN(n6927) );
  AOI21_X1 U8089 ( .B1(n7206), .B2(n9235), .A(n6927), .ZN(n7177) );
  XNOR2_X1 U8090 ( .A(n7176), .B(n7177), .ZN(n7174) );
  XNOR2_X1 U8091 ( .A(n7175), .B(n7174), .ZN(n6928) );
  NAND2_X1 U8092 ( .A1(n6928), .A2(n9376), .ZN(n6942) );
  NAND2_X1 U8093 ( .A1(n6031), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6937) );
  OR2_X1 U8094 ( .A1(n6929), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6930) );
  AND2_X1 U8095 ( .A1(n7190), .A2(n6930), .ZN(n7217) );
  NAND2_X1 U8096 ( .A1(n6931), .A2(n7217), .ZN(n6936) );
  NAND2_X1 U8097 ( .A1(n6933), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6935) );
  NAND2_X1 U8098 ( .A1(n9423), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6934) );
  INV_X1 U8099 ( .A(n10714), .ZN(n9671) );
  INV_X1 U8100 ( .A(n7016), .ZN(n6938) );
  OAI22_X1 U8101 ( .A1(n7047), .A2(n9402), .B1(n9401), .B2(n6938), .ZN(n6939)
         );
  AOI211_X1 U8102 ( .C1(n9406), .C2(n9671), .A(n6940), .B(n6939), .ZN(n6941)
         );
  OAI211_X1 U8103 ( .C1(n10685), .C2(n9384), .A(n6942), .B(n6941), .ZN(
        P1_U3211) );
  NAND2_X1 U8104 ( .A1(n6961), .A2(n5317), .ZN(n6943) );
  OR2_X1 U8105 ( .A1(n6702), .A2(n6945), .ZN(n6951) );
  OR2_X1 U8106 ( .A1(n5137), .A2(n6947), .ZN(n6950) );
  NAND2_X1 U8107 ( .A1(n8134), .A2(n6948), .ZN(n6949) );
  XNOR2_X1 U8108 ( .A(n7141), .B(n8263), .ZN(n6999) );
  NAND2_X1 U8109 ( .A1(n8192), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6959) );
  NAND2_X1 U8110 ( .A1(n6952), .A2(n10331), .ZN(n6953) );
  AND2_X1 U8111 ( .A1(n7103), .A2(n6953), .ZN(n7138) );
  NAND2_X1 U8112 ( .A1(n6516), .A2(n7138), .ZN(n6958) );
  INV_X1 U8113 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n6954) );
  OR2_X1 U8114 ( .A1(n8169), .A2(n6954), .ZN(n6957) );
  INV_X1 U8115 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6955) );
  OR2_X1 U8116 ( .A1(n8171), .A2(n6955), .ZN(n6956) );
  NAND4_X1 U8117 ( .A1(n6959), .A2(n6958), .A3(n6957), .A4(n6956), .ZN(n8703)
         );
  NAND2_X1 U8118 ( .A1(n8703), .A2(n9014), .ZN(n6960) );
  OAI21_X1 U8119 ( .B1(n6961), .B2(n8806), .A(n6960), .ZN(n6991) );
  INV_X1 U8120 ( .A(n7135), .ZN(n7137) );
  AOI211_X1 U8121 ( .C1(n8042), .C2(n6962), .A(n10862), .B(n7137), .ZN(n6990)
         );
  AOI211_X1 U8122 ( .C1(n9124), .C2(n8042), .A(n6991), .B(n6990), .ZN(n6967)
         );
  NAND2_X1 U8123 ( .A1(n8047), .A2(n6964), .ZN(n6963) );
  MUX2_X1 U8124 ( .A(n8047), .B(n6963), .S(n7131), .Z(n6966) );
  INV_X1 U8125 ( .A(n6964), .ZN(n6965) );
  NAND3_X1 U8126 ( .A1(n6966), .A2(n7130), .A3(n9017), .ZN(n6993) );
  OAI211_X1 U8127 ( .C1(n10841), .C2(n6999), .A(n6967), .B(n6993), .ZN(n6969)
         );
  NAND2_X1 U8128 ( .A1(n6969), .A2(n10873), .ZN(n6968) );
  OAI21_X1 U8129 ( .B1(n10873), .B2(n6739), .A(n6968), .ZN(P2_U3466) );
  NAND2_X1 U8130 ( .A1(n6969), .A2(n10870), .ZN(n6970) );
  OAI21_X1 U8131 ( .B1(n10870), .B2(n6286), .A(n6970), .ZN(P2_U3525) );
  INV_X1 U8132 ( .A(n6992), .ZN(n6983) );
  XNOR2_X1 U8133 ( .A(n6765), .B(n7142), .ZN(n6972) );
  AND2_X1 U8134 ( .A1(n8704), .A2(n8531), .ZN(n6971) );
  NOR2_X1 U8135 ( .A1(n6971), .A2(n6972), .ZN(n7097) );
  AOI21_X1 U8136 ( .B1(n6972), .B2(n6971), .A(n7097), .ZN(n6977) );
  INV_X1 U8137 ( .A(n6973), .ZN(n6974) );
  OAI21_X1 U8138 ( .B1(n6977), .B2(n6976), .A(n7099), .ZN(n6978) );
  NAND2_X1 U8139 ( .A1(n6978), .A2(n8683), .ZN(n6982) );
  NOR2_X1 U8140 ( .A1(n8693), .A2(n7142), .ZN(n6980) );
  AOI211_X1 U8141 ( .C1(n6991), .C2(n8676), .A(n6980), .B(n6979), .ZN(n6981)
         );
  OAI211_X1 U8142 ( .C1(n8674), .C2(n6983), .A(n6982), .B(n6981), .ZN(P2_U3229) );
  MUX2_X1 U8143 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7958), .Z(n6986) );
  NAND2_X1 U8144 ( .A1(n6986), .A2(SI_18_), .ZN(n7084) );
  OAI21_X1 U8145 ( .B1(n6986), .B2(SI_18_), .A(n7084), .ZN(n7081) );
  XNOR2_X1 U8146 ( .A(n7083), .B(n7081), .ZN(n8347) );
  INV_X1 U8147 ( .A(n8347), .ZN(n7039) );
  NAND2_X1 U8148 ( .A1(n6987), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6988) );
  XNOR2_X1 U8149 ( .A(n6988), .B(P1_IR_REG_18__SCAN_IN), .ZN(n8348) );
  AOI22_X1 U8150 ( .A1(n8348), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10445), .ZN(n6989) );
  OAI21_X1 U8151 ( .B1(n7039), .B2(n10451), .A(n6989), .ZN(P1_U3335) );
  INV_X1 U8152 ( .A(n6990), .ZN(n6995) );
  AOI21_X1 U8153 ( .B1(n6992), .B2(n10801), .A(n6991), .ZN(n6994) );
  OAI211_X1 U8154 ( .C1(n6995), .C2(n5256), .A(n6994), .B(n6993), .ZN(n6996)
         );
  NAND2_X1 U8155 ( .A1(n6996), .A2(n10811), .ZN(n6998) );
  AOI22_X1 U8156 ( .A1(n9035), .A2(n8042), .B1(P2_REG2_REG_5__SCAN_IN), .B2(
        n10813), .ZN(n6997) );
  OAI211_X1 U8157 ( .C1(n6999), .C2(n9022), .A(n6998), .B(n6997), .ZN(P2_U3291) );
  OR2_X1 U8158 ( .A1(n7206), .A2(n7198), .ZN(n9510) );
  NAND2_X1 U8159 ( .A1(n7206), .A2(n7198), .ZN(n9506) );
  NAND2_X1 U8160 ( .A1(n9510), .A2(n9506), .ZN(n9634) );
  INV_X1 U8161 ( .A(n9454), .ZN(n7000) );
  NAND2_X1 U8162 ( .A1(n7164), .A2(n7047), .ZN(n9507) );
  NAND2_X1 U8163 ( .A1(n7002), .A2(n7077), .ZN(n7022) );
  AND2_X1 U8164 ( .A1(n9507), .A2(n7022), .ZN(n9457) );
  OR2_X1 U8165 ( .A1(n7164), .A2(n7047), .ZN(n9505) );
  XOR2_X1 U8166 ( .A(n9634), .B(n7204), .Z(n7014) );
  NAND2_X1 U8167 ( .A1(n7046), .A2(n7003), .ZN(n7004) );
  NAND2_X1 U8168 ( .A1(n7005), .A2(n7004), .ZN(n7040) );
  INV_X1 U8169 ( .A(n7040), .ZN(n7007) );
  XNOR2_X1 U8170 ( .A(n9673), .B(n7077), .ZN(n9629) );
  INV_X1 U8171 ( .A(n9629), .ZN(n7006) );
  NAND2_X1 U8172 ( .A1(n9673), .A2(n7077), .ZN(n7008) );
  INV_X1 U8173 ( .A(n9632), .ZN(n7009) );
  INV_X1 U8174 ( .A(n7047), .ZN(n9672) );
  OR2_X1 U8175 ( .A1(n7164), .A2(n9672), .ZN(n7010) );
  NAND2_X1 U8176 ( .A1(n7024), .A2(n7010), .ZN(n7011) );
  OAI21_X1 U8177 ( .B1(n7011), .B2(n9634), .A(n7208), .ZN(n10688) );
  OAI22_X1 U8178 ( .A1(n10714), .A2(n10753), .B1(n7047), .B2(n10755), .ZN(
        n7012) );
  AOI21_X1 U8179 ( .B1(n10688), .B2(n10822), .A(n7012), .ZN(n7013) );
  OAI21_X1 U8180 ( .B1(n9888), .B2(n7014), .A(n7013), .ZN(n10686) );
  INV_X1 U8181 ( .A(n10686), .ZN(n7021) );
  OAI211_X1 U8182 ( .C1(n7030), .C2(n10685), .A(n7215), .B(n10878), .ZN(n10684) );
  OR2_X1 U8183 ( .A1(n7015), .A2(n9760), .ZN(n9924) );
  INV_X1 U8184 ( .A(n9897), .ZN(n10776) );
  AOI22_X1 U8185 ( .A1(n10778), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7016), .B2(
        n10776), .ZN(n7018) );
  NAND2_X1 U8186 ( .A1(n9920), .A2(n7206), .ZN(n7017) );
  OAI211_X1 U8187 ( .C1(n10684), .C2(n9924), .A(n7018), .B(n7017), .ZN(n7019)
         );
  AOI21_X1 U8188 ( .B1(n10688), .B2(n10773), .A(n7019), .ZN(n7020) );
  OAI21_X1 U8189 ( .B1(n7021), .B2(n10778), .A(n7020), .ZN(P1_U3284) );
  INV_X1 U8190 ( .A(n7022), .ZN(n7023) );
  OAI21_X1 U8191 ( .B1(n7044), .B2(n7023), .A(n9459), .ZN(n9509) );
  XOR2_X1 U8192 ( .A(n9632), .B(n9509), .Z(n7029) );
  INV_X1 U8193 ( .A(n7024), .ZN(n7025) );
  AOI21_X1 U8194 ( .B1(n9632), .B2(n7026), .A(n7025), .ZN(n7168) );
  AOI22_X1 U8195 ( .A1(n7211), .A2(n9910), .B1(n9912), .B2(n9673), .ZN(n7027)
         );
  OAI21_X1 U8196 ( .B1(n7168), .B2(n10718), .A(n7027), .ZN(n7028) );
  AOI21_X1 U8197 ( .B1(n10758), .B2(n7029), .A(n7028), .ZN(n7167) );
  AOI21_X1 U8198 ( .B1(n7164), .B2(n7048), .A(n7030), .ZN(n7165) );
  INV_X1 U8199 ( .A(n7164), .ZN(n7033) );
  AOI22_X1 U8200 ( .A1(n10778), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7031), .B2(
        n10776), .ZN(n7032) );
  OAI21_X1 U8201 ( .B1(n7033), .B2(n10780), .A(n7032), .ZN(n7035) );
  NOR2_X1 U8202 ( .A1(n7168), .A2(n9867), .ZN(n7034) );
  AOI211_X1 U8203 ( .C1(n7165), .C2(n10772), .A(n7035), .B(n7034), .ZN(n7036)
         );
  OAI21_X1 U8204 ( .B1(n10778), .B2(n7167), .A(n7036), .ZN(P1_U3285) );
  XNOR2_X1 U8205 ( .A(n7037), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8729) );
  INV_X1 U8206 ( .A(n8729), .ZN(n8727) );
  OAI222_X1 U8207 ( .A1(n8727), .A2(P2_U3152), .B1(n9153), .B2(n7039), .C1(
        n9151), .C2(n7038), .ZN(P2_U3340) );
  INV_X1 U8208 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7052) );
  NAND2_X1 U8209 ( .A1(n7040), .A2(n9629), .ZN(n7041) );
  NAND2_X1 U8210 ( .A1(n7042), .A2(n7041), .ZN(n7080) );
  AOI21_X1 U8211 ( .B1(n7043), .B2(n7077), .A(n10833), .ZN(n7049) );
  XOR2_X1 U8212 ( .A(n9629), .B(n7044), .Z(n7045) );
  OAI222_X1 U8213 ( .A1(n10753), .A2(n7047), .B1(n10755), .B2(n7046), .C1(
        n9888), .C2(n7045), .ZN(n7073) );
  AOI21_X1 U8214 ( .B1(n7049), .B2(n7048), .A(n7073), .ZN(n7070) );
  NAND2_X1 U8215 ( .A1(n7077), .A2(n10877), .ZN(n7050) );
  OAI211_X1 U8216 ( .C1(n10831), .C2(n7080), .A(n7070), .B(n7050), .ZN(n7053)
         );
  NAND2_X1 U8217 ( .A1(n7053), .A2(n5045), .ZN(n7051) );
  OAI21_X1 U8218 ( .B1(n5045), .B2(n7052), .A(n7051), .ZN(P1_U3469) );
  INV_X1 U8219 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7055) );
  NAND2_X1 U8220 ( .A1(n7053), .A2(n10722), .ZN(n7054) );
  OAI21_X1 U8221 ( .B1(n10722), .B2(n7055), .A(n7054), .ZN(P1_U3528) );
  OAI21_X1 U8222 ( .B1(n7057), .B2(n6462), .A(n7056), .ZN(n7060) );
  INV_X1 U8223 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7058) );
  MUX2_X1 U8224 ( .A(n7058), .B(P2_REG1_REG_12__SCAN_IN), .S(n7574), .Z(n7059)
         );
  NOR2_X1 U8225 ( .A1(n7059), .A2(n7060), .ZN(n7151) );
  AOI21_X1 U8226 ( .B1(n7060), .B2(n7059), .A(n7151), .ZN(n7063) );
  NAND2_X1 U8227 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7714) );
  INV_X1 U8228 ( .A(n7714), .ZN(n7061) );
  AOI21_X1 U8229 ( .B1(n10606), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7061), .ZN(
        n7062) );
  OAI21_X1 U8230 ( .B1(n10586), .B2(n7063), .A(n7062), .ZN(n7068) );
  INV_X1 U8231 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7542) );
  MUX2_X1 U8232 ( .A(n7542), .B(P2_REG2_REG_12__SCAN_IN), .S(n7574), .Z(n7065)
         );
  NOR2_X1 U8233 ( .A1(n7065), .A2(n7066), .ZN(n7155) );
  AOI211_X1 U8234 ( .C1(n7066), .C2(n7065), .A(n7155), .B(n10607), .ZN(n7067)
         );
  AOI211_X1 U8235 ( .C1(n10613), .C2(n7574), .A(n7068), .B(n7067), .ZN(n7069)
         );
  INV_X1 U8236 ( .A(n7069), .ZN(P2_U3257) );
  OAI21_X1 U8237 ( .B1(n7071), .B2(n7080), .A(n7070), .ZN(n7072) );
  OAI211_X1 U8238 ( .C1(n9812), .C2(n7073), .A(n7072), .B(n10783), .ZN(n7079)
         );
  INV_X1 U8239 ( .A(n7074), .ZN(n7075) );
  OAI22_X1 U8240 ( .A1(n10783), .A2(n5837), .B1(n7075), .B2(n9897), .ZN(n7076)
         );
  AOI21_X1 U8241 ( .B1(n9920), .B2(n7077), .A(n7076), .ZN(n7078) );
  OAI211_X1 U8242 ( .C1(n7080), .C2(n9867), .A(n7079), .B(n7078), .ZN(P1_U3286) );
  INV_X1 U8243 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7086) );
  INV_X1 U8244 ( .A(n7081), .ZN(n7082) );
  NAND2_X1 U8245 ( .A1(n7083), .A2(n7082), .ZN(n7085) );
  MUX2_X1 U8246 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n5713), .Z(n7258) );
  XNOR2_X1 U8247 ( .A(n7258), .B(SI_19_), .ZN(n7261) );
  XNOR2_X1 U8248 ( .A(n7262), .B(n7261), .ZN(n8351) );
  INV_X1 U8249 ( .A(n8351), .ZN(n7088) );
  OAI222_X1 U8250 ( .A1(n10455), .A2(n7086), .B1(n10451), .B2(n7088), .C1(
        P1_U3084), .C2(n9812), .ZN(P1_U3334) );
  INV_X1 U8251 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7087) );
  OAI222_X1 U8252 ( .A1(P2_U3152), .A2(n6499), .B1(n9153), .B2(n7088), .C1(
        n7087), .C2(n9151), .ZN(P2_U3339) );
  INV_X1 U8253 ( .A(n7138), .ZN(n7116) );
  NAND2_X1 U8254 ( .A1(n8134), .A2(n7090), .ZN(n7093) );
  OR2_X1 U8255 ( .A1(n6946), .A2(n7091), .ZN(n7092) );
  XNOR2_X1 U8256 ( .A(n10677), .B(n6765), .ZN(n7096) );
  AND2_X1 U8257 ( .A1(n8703), .A2(n8531), .ZN(n7095) );
  NOR2_X1 U8258 ( .A1(n7095), .A2(n7096), .ZN(n7223) );
  AOI21_X1 U8259 ( .B1(n7096), .B2(n7095), .A(n7223), .ZN(n7101) );
  INV_X1 U8260 ( .A(n7097), .ZN(n7098) );
  OAI21_X1 U8261 ( .B1(n7101), .B2(n7100), .A(n7225), .ZN(n7102) );
  NAND2_X1 U8262 ( .A1(n7102), .A2(n8683), .ZN(n7115) );
  INV_X1 U8263 ( .A(n8704), .ZN(n8043) );
  NAND2_X1 U8264 ( .A1(n7103), .A2(n8554), .ZN(n7104) );
  AND2_X1 U8265 ( .A1(n7236), .A2(n7104), .ZN(n8561) );
  NAND2_X1 U8266 ( .A1(n8191), .A2(n8561), .ZN(n7109) );
  NAND2_X1 U8267 ( .A1(n8192), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7108) );
  INV_X1 U8268 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7105) );
  OR2_X1 U8269 ( .A1(n8169), .A2(n7105), .ZN(n7107) );
  OR2_X1 U8270 ( .A1(n8171), .A2(n6271), .ZN(n7106) );
  NAND4_X1 U8271 ( .A1(n7109), .A2(n7108), .A3(n7107), .A4(n7106), .ZN(n8702)
         );
  NAND2_X1 U8272 ( .A1(n8685), .A2(n8702), .ZN(n7112) );
  INV_X1 U8273 ( .A(n7110), .ZN(n7111) );
  OAI211_X1 U8274 ( .C1(n8043), .C2(n8688), .A(n7112), .B(n7111), .ZN(n7113)
         );
  AOI21_X1 U8275 ( .B1(n8651), .B2(n8049), .A(n7113), .ZN(n7114) );
  OAI211_X1 U8276 ( .C1(n8674), .C2(n7116), .A(n7115), .B(n7114), .ZN(P2_U3241) );
  INV_X1 U8277 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7120) );
  OR2_X1 U8278 ( .A1(n7751), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7117) );
  NAND2_X1 U8279 ( .A1(n7118), .A2(n7117), .ZN(n7349) );
  XOR2_X1 U8280 ( .A(n7756), .B(n7349), .Z(n7119) );
  NOR2_X1 U8281 ( .A1(n7119), .A2(n7120), .ZN(n7350) );
  AOI211_X1 U8282 ( .C1(n7120), .C2(n7119), .A(n7688), .B(n7350), .ZN(n7128)
         );
  INV_X1 U8283 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10883) );
  OR2_X1 U8284 ( .A1(n7751), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7121) );
  NAND2_X1 U8285 ( .A1(n7122), .A2(n7121), .ZN(n7355) );
  XOR2_X1 U8286 ( .A(n7756), .B(n7355), .Z(n7123) );
  NOR2_X1 U8287 ( .A1(n7123), .A2(n10883), .ZN(n7356) );
  AOI211_X1 U8288 ( .C1(n10883), .C2(n7123), .A(n10621), .B(n7356), .ZN(n7127)
         );
  NAND2_X1 U8289 ( .A1(n10550), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n7124) );
  NAND2_X1 U8290 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9399) );
  OAI211_X1 U8291 ( .C1(n10628), .C2(n7125), .A(n7124), .B(n9399), .ZN(n7126)
         );
  OR3_X1 U8292 ( .A1(n7128), .A2(n7127), .A3(n7126), .ZN(P1_U3256) );
  NAND2_X1 U8293 ( .A1(n8704), .A2(n7142), .ZN(n7129) );
  INV_X1 U8294 ( .A(n8703), .ZN(n8557) );
  NAND2_X1 U8295 ( .A1(n8557), .A2(n10677), .ZN(n8050) );
  NAND2_X1 U8296 ( .A1(n8703), .A2(n8049), .ZN(n8052) );
  NAND2_X1 U8297 ( .A1(n8050), .A2(n8052), .ZN(n8264) );
  XNOR2_X1 U8298 ( .A(n7344), .B(n7145), .ZN(n7132) );
  NAND2_X1 U8299 ( .A1(n7132), .A2(n9017), .ZN(n7134) );
  AOI22_X1 U8300 ( .A1(n9012), .A2(n8704), .B1(n8702), .B2(n9014), .ZN(n7133)
         );
  NAND2_X1 U8301 ( .A1(n7134), .A2(n7133), .ZN(n10679) );
  INV_X1 U8302 ( .A(n7340), .ZN(n7136) );
  OAI21_X1 U8303 ( .B1(n10677), .B2(n7137), .A(n7136), .ZN(n10678) );
  AOI22_X1 U8304 ( .A1(n10813), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n7138), .B2(
        n10801), .ZN(n7140) );
  NAND2_X1 U8305 ( .A1(n9035), .A2(n8049), .ZN(n7139) );
  OAI211_X1 U8306 ( .C1(n10678), .C2(n8793), .A(n7140), .B(n7139), .ZN(n7149)
         );
  NAND2_X1 U8307 ( .A1(n8043), .A2(n7142), .ZN(n7143) );
  INV_X1 U8308 ( .A(n10681), .ZN(n7147) );
  AND2_X1 U8309 ( .A1(n8264), .A2(n7146), .ZN(n10676) );
  NOR3_X1 U8310 ( .A1(n7147), .A2(n10676), .A3(n9022), .ZN(n7148) );
  AOI211_X1 U8311 ( .C1(n10811), .C2(n10679), .A(n7149), .B(n7148), .ZN(n7150)
         );
  INV_X1 U8312 ( .A(n7150), .ZN(P2_U3290) );
  AOI21_X1 U8313 ( .B1(n7152), .B2(n7058), .A(n7151), .ZN(n7154) );
  INV_X1 U8314 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10849) );
  AOI22_X1 U8315 ( .A1(n7813), .A2(n10849), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n7287), .ZN(n7153) );
  NOR2_X1 U8316 ( .A1(n7154), .A2(n7153), .ZN(n7286) );
  AOI21_X1 U8317 ( .B1(n7154), .B2(n7153), .A(n7286), .ZN(n7163) );
  INV_X1 U8318 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7156) );
  AOI22_X1 U8319 ( .A1(n7813), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7156), .B2(
        n7287), .ZN(n7157) );
  NAND2_X1 U8320 ( .A1(n7158), .A2(n7157), .ZN(n7291) );
  OAI21_X1 U8321 ( .B1(n7158), .B2(n7157), .A(n7291), .ZN(n7159) );
  NAND2_X1 U8322 ( .A1(n7159), .A2(n10584), .ZN(n7162) );
  INV_X1 U8323 ( .A(n10606), .ZN(n10594) );
  INV_X1 U8324 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7617) );
  NAND2_X1 U8325 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3152), .ZN(n7856) );
  OAI21_X1 U8326 ( .B1(n10594), .B2(n7617), .A(n7856), .ZN(n7160) );
  AOI21_X1 U8327 ( .B1(n7813), .B2(n10613), .A(n7160), .ZN(n7161) );
  OAI211_X1 U8328 ( .C1(n7163), .C2(n10586), .A(n7162), .B(n7161), .ZN(
        P2_U3258) );
  INV_X1 U8329 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7170) );
  AOI22_X1 U8330 ( .A1(n7165), .A2(n10878), .B1(n10877), .B2(n7164), .ZN(n7166) );
  OAI211_X1 U8331 ( .C1(n7168), .C2(n10817), .A(n7167), .B(n7166), .ZN(n7171)
         );
  NAND2_X1 U8332 ( .A1(n7171), .A2(n10722), .ZN(n7169) );
  OAI21_X1 U8333 ( .B1(n10722), .B2(n7170), .A(n7169), .ZN(P1_U3529) );
  INV_X1 U8334 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7173) );
  NAND2_X1 U8335 ( .A1(n7171), .A2(n5045), .ZN(n7172) );
  OAI21_X1 U8336 ( .B1(n5045), .B2(n7173), .A(n7172), .ZN(P1_U3472) );
  INV_X1 U8337 ( .A(n7176), .ZN(n7178) );
  NAND2_X1 U8338 ( .A1(n7178), .A2(n7177), .ZN(n7179) );
  OR2_X1 U8339 ( .A1(n7232), .A2(n6231), .ZN(n7182) );
  AOI22_X1 U8340 ( .A1(n8442), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n8352), .B2(
        n7180), .ZN(n7181) );
  NOR2_X1 U8341 ( .A1(n10714), .A2(n9286), .ZN(n7183) );
  AOI21_X1 U8342 ( .B1(n7393), .B2(n9235), .A(n7183), .ZN(n7184) );
  NAND2_X1 U8343 ( .A1(n7266), .A2(n7267), .ZN(n7188) );
  OR2_X1 U8344 ( .A1(n10714), .A2(n9287), .ZN(n7185) );
  NAND2_X1 U8345 ( .A1(n7186), .A2(n7185), .ZN(n7187) );
  XNOR2_X1 U8346 ( .A(n7187), .B(n9208), .ZN(n7265) );
  XNOR2_X1 U8347 ( .A(n7188), .B(n7265), .ZN(n7202) );
  NAND2_X1 U8348 ( .A1(n6031), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7195) );
  NAND2_X1 U8349 ( .A1(n7190), .A2(n7189), .ZN(n7191) );
  AND2_X1 U8350 ( .A1(n7275), .A2(n7191), .ZN(n10728) );
  NAND2_X1 U8351 ( .A1(n6931), .A2(n10728), .ZN(n7194) );
  NAND2_X1 U8352 ( .A1(n6933), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7193) );
  NAND2_X1 U8353 ( .A1(n9423), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7192) );
  NAND4_X1 U8354 ( .A1(n7195), .A2(n7194), .A3(n7193), .A4(n7192), .ZN(n9670)
         );
  INV_X1 U8355 ( .A(n9670), .ZN(n7397) );
  INV_X1 U8356 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7196) );
  OAI22_X1 U8357 ( .A1(n9388), .A2(n7397), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7196), .ZN(n7200) );
  INV_X1 U8358 ( .A(n7217), .ZN(n7197) );
  OAI22_X1 U8359 ( .A1(n7198), .A2(n9402), .B1(n9401), .B2(n7197), .ZN(n7199)
         );
  AOI211_X1 U8360 ( .C1(n7393), .C2(n9407), .A(n7200), .B(n7199), .ZN(n7201)
         );
  OAI21_X1 U8361 ( .B1(n7202), .B2(n9410), .A(n7201), .ZN(P1_U3219) );
  INV_X1 U8362 ( .A(n9510), .ZN(n7203) );
  INV_X1 U8363 ( .A(n9506), .ZN(n7205) );
  OR2_X1 U8364 ( .A1(n7393), .A2(n10714), .ZN(n9462) );
  NAND2_X1 U8365 ( .A1(n7393), .A2(n10714), .ZN(n9503) );
  XNOR2_X1 U8366 ( .A(n5133), .B(n5538), .ZN(n7214) );
  OR2_X1 U8367 ( .A1(n7206), .A2(n7211), .ZN(n7207) );
  NAND2_X1 U8368 ( .A1(n7209), .A2(n9511), .ZN(n7210) );
  NAND2_X1 U8369 ( .A1(n7395), .A2(n7210), .ZN(n7302) );
  AOI22_X1 U8370 ( .A1(n7211), .A2(n9912), .B1(n9910), .B2(n9670), .ZN(n7212)
         );
  OAI21_X1 U8371 ( .B1(n7302), .B2(n10718), .A(n7212), .ZN(n7213) );
  AOI21_X1 U8372 ( .B1(n7214), .B2(n10758), .A(n7213), .ZN(n7301) );
  NAND2_X1 U8373 ( .A1(n7215), .A2(n7393), .ZN(n7216) );
  AND2_X1 U8374 ( .A1(n10708), .A2(n7216), .ZN(n7299) );
  INV_X1 U8375 ( .A(n7393), .ZN(n7219) );
  AOI22_X1 U8376 ( .A1(n10778), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7217), .B2(
        n10776), .ZN(n7218) );
  OAI21_X1 U8377 ( .B1(n7219), .B2(n10780), .A(n7218), .ZN(n7221) );
  NOR2_X1 U8378 ( .A1(n7302), .A2(n9867), .ZN(n7220) );
  AOI211_X1 U8379 ( .C1(n7299), .C2(n10772), .A(n7221), .B(n7220), .ZN(n7222)
         );
  OAI21_X1 U8380 ( .B1(n10778), .B2(n7301), .A(n7222), .ZN(P1_U3283) );
  INV_X1 U8381 ( .A(n7223), .ZN(n7224) );
  NAND2_X1 U8382 ( .A1(n7225), .A2(n7224), .ZN(n8551) );
  NAND2_X1 U8383 ( .A1(n7226), .A2(n8211), .ZN(n7229) );
  AOI22_X1 U8384 ( .A1(n8135), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8134), .B2(
        n7227), .ZN(n7228) );
  NAND2_X1 U8385 ( .A1(n7229), .A2(n7228), .ZN(n8560) );
  XNOR2_X1 U8386 ( .A(n8560), .B(n6765), .ZN(n7231) );
  NAND2_X1 U8387 ( .A1(n8702), .A2(n8531), .ZN(n7230) );
  XNOR2_X1 U8388 ( .A(n7231), .B(n7230), .ZN(n8552) );
  OR2_X1 U8389 ( .A1(n7232), .A2(n6702), .ZN(n7235) );
  AOI22_X1 U8390 ( .A1(n8135), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8134), .B2(
        n7233), .ZN(n7234) );
  XNOR2_X1 U8391 ( .A(n10702), .B(n6765), .ZN(n7438) );
  NAND2_X1 U8392 ( .A1(n8192), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7243) );
  NAND2_X1 U8393 ( .A1(n7236), .A2(n10293), .ZN(n7237) );
  AND2_X1 U8394 ( .A1(n7244), .A2(n7237), .ZN(n9030) );
  NAND2_X1 U8395 ( .A1(n8191), .A2(n9030), .ZN(n7242) );
  INV_X1 U8396 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7238) );
  OR2_X1 U8397 ( .A1(n8169), .A2(n7238), .ZN(n7241) );
  INV_X1 U8398 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7239) );
  OR2_X1 U8399 ( .A1(n8171), .A2(n7239), .ZN(n7240) );
  NAND4_X1 U8400 ( .A1(n7243), .A2(n7242), .A3(n7241), .A4(n7240), .ZN(n8701)
         );
  NAND2_X1 U8401 ( .A1(n8701), .A2(n8531), .ZN(n7436) );
  XNOR2_X1 U8402 ( .A(n7438), .B(n7436), .ZN(n7439) );
  XNOR2_X1 U8403 ( .A(n7440), .B(n7439), .ZN(n7257) );
  NOR2_X1 U8404 ( .A1(n10702), .A2(n8693), .ZN(n7255) );
  INV_X1 U8405 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10105) );
  NAND2_X1 U8406 ( .A1(n7244), .A2(n10105), .ZN(n7245) );
  AND2_X1 U8407 ( .A1(n7373), .A2(n7245), .ZN(n7450) );
  NAND2_X1 U8408 ( .A1(n6516), .A2(n7450), .ZN(n7251) );
  NAND2_X1 U8409 ( .A1(n8192), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7250) );
  INV_X1 U8410 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7246) );
  OR2_X1 U8411 ( .A1(n8169), .A2(n7246), .ZN(n7249) );
  INV_X1 U8412 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7247) );
  OR2_X1 U8413 ( .A1(n8171), .A2(n7247), .ZN(n7248) );
  NAND4_X1 U8414 ( .A1(n7251), .A2(n7250), .A3(n7249), .A4(n7248), .ZN(n8700)
         );
  NAND2_X1 U8415 ( .A1(n8700), .A2(n9014), .ZN(n7253) );
  NAND2_X1 U8416 ( .A1(n8702), .A2(n9012), .ZN(n7252) );
  AND2_X1 U8417 ( .A1(n7253), .A2(n7252), .ZN(n9024) );
  INV_X1 U8418 ( .A(n8676), .ZN(n8612) );
  OAI22_X1 U8419 ( .A1(n9024), .A2(n8612), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10293), .ZN(n7254) );
  AOI211_X1 U8420 ( .C1(n8690), .C2(n9030), .A(n7255), .B(n7254), .ZN(n7256)
         );
  OAI21_X1 U8421 ( .B1(n7257), .B2(n8667), .A(n7256), .ZN(P2_U3223) );
  INV_X1 U8422 ( .A(n7258), .ZN(n7259) );
  NAND2_X1 U8423 ( .A1(n7259), .A2(n10244), .ZN(n7260) );
  MUX2_X1 U8424 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n7958), .Z(n7310) );
  XNOR2_X1 U8425 ( .A(n7310), .B(n10039), .ZN(n7308) );
  XNOR2_X1 U8426 ( .A(n7309), .B(n7308), .ZN(n8362) );
  INV_X1 U8427 ( .A(n8362), .ZN(n8546) );
  INV_X1 U8428 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7263) );
  OAI222_X1 U8429 ( .A1(n10451), .A2(n8546), .B1(n7264), .B2(P1_U3084), .C1(
        n7263), .C2(n10455), .ZN(P1_U3333) );
  NAND2_X1 U8430 ( .A1(n7370), .A2(n9427), .ZN(n7269) );
  AOI22_X1 U8431 ( .A1(n8442), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8352), .B2(
        n10525), .ZN(n7268) );
  NAND2_X1 U8432 ( .A1(n9670), .A2(n9198), .ZN(n7270) );
  NAND2_X1 U8433 ( .A1(n7271), .A2(n7270), .ZN(n7272) );
  XNOR2_X1 U8434 ( .A(n7272), .B(n9243), .ZN(n7321) );
  AND2_X1 U8435 ( .A1(n9670), .A2(n9239), .ZN(n7273) );
  AOI21_X1 U8436 ( .B1(n7400), .B2(n9235), .A(n7273), .ZN(n7322) );
  XNOR2_X1 U8437 ( .A(n7321), .B(n7322), .ZN(n7319) );
  XOR2_X1 U8438 ( .A(n7320), .B(n7319), .Z(n7285) );
  NAND2_X1 U8439 ( .A1(n6031), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7281) );
  NAND2_X1 U8440 ( .A1(n7275), .A2(n7274), .ZN(n7276) );
  AND2_X1 U8441 ( .A1(n7277), .A2(n7276), .ZN(n7402) );
  NAND2_X1 U8442 ( .A1(n6931), .A2(n7402), .ZN(n7280) );
  NAND2_X1 U8443 ( .A1(n6933), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7279) );
  NAND2_X1 U8444 ( .A1(n9423), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n7278) );
  AOI22_X1 U8445 ( .A1(n9381), .A2(n9671), .B1(n9347), .B2(n10728), .ZN(n7282)
         );
  NAND2_X1 U8446 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3084), .ZN(n10535) );
  OAI211_X1 U8447 ( .C1(n10756), .C2(n9388), .A(n7282), .B(n10535), .ZN(n7283)
         );
  AOI21_X1 U8448 ( .B1(n7400), .B2(n9407), .A(n7283), .ZN(n7284) );
  OAI21_X1 U8449 ( .B1(n7285), .B2(n9410), .A(n7284), .ZN(P1_U3229) );
  AOI21_X1 U8450 ( .B1(n7287), .B2(n10849), .A(n7286), .ZN(n7289) );
  INV_X1 U8451 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10869) );
  AOI22_X1 U8452 ( .A1(n7864), .A2(n10869), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n7559), .ZN(n7288) );
  NOR2_X1 U8453 ( .A1(n7289), .A2(n7288), .ZN(n7558) );
  AOI21_X1 U8454 ( .B1(n7289), .B2(n7288), .A(n7558), .ZN(n7298) );
  INV_X1 U8455 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7290) );
  AOI22_X1 U8456 ( .A1(n7864), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7290), .B2(
        n7559), .ZN(n7293) );
  OAI21_X1 U8457 ( .B1(n7813), .B2(P2_REG2_REG_13__SCAN_IN), .A(n7291), .ZN(
        n7292) );
  NAND2_X1 U8458 ( .A1(n7293), .A2(n7292), .ZN(n7552) );
  OAI21_X1 U8459 ( .B1(n7293), .B2(n7292), .A(n7552), .ZN(n7296) );
  INV_X1 U8460 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7872) );
  NOR2_X1 U8461 ( .A1(n7872), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7901) );
  AOI21_X1 U8462 ( .B1(n10606), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n7901), .ZN(
        n7294) );
  OAI21_X1 U8463 ( .B1(n10585), .B2(n7559), .A(n7294), .ZN(n7295) );
  AOI21_X1 U8464 ( .B1(n7296), .B2(n10584), .A(n7295), .ZN(n7297) );
  OAI21_X1 U8465 ( .B1(n7298), .B2(n10586), .A(n7297), .ZN(P2_U3259) );
  AOI22_X1 U8466 ( .A1(n7299), .A2(n10878), .B1(n10877), .B2(n7393), .ZN(n7300) );
  OAI211_X1 U8467 ( .C1(n10817), .C2(n7302), .A(n7301), .B(n7300), .ZN(n7305)
         );
  NAND2_X1 U8468 ( .A1(n7305), .A2(n10722), .ZN(n7303) );
  OAI21_X1 U8469 ( .B1(n10722), .B2(n7304), .A(n7303), .ZN(P1_U3531) );
  INV_X1 U8470 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7307) );
  NAND2_X1 U8471 ( .A1(n7305), .A2(n5045), .ZN(n7306) );
  OAI21_X1 U8472 ( .B1(n5045), .B2(n7307), .A(n7306), .ZN(P1_U3478) );
  NAND2_X1 U8473 ( .A1(n7309), .A2(n7308), .ZN(n7313) );
  INV_X1 U8474 ( .A(n7310), .ZN(n7311) );
  NAND2_X1 U8475 ( .A1(n7311), .A2(n10039), .ZN(n7312) );
  MUX2_X1 U8476 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n5713), .Z(n7314) );
  NAND2_X1 U8477 ( .A1(n7314), .A2(SI_21_), .ZN(n7471) );
  OAI21_X1 U8478 ( .B1(n7314), .B2(SI_21_), .A(n7471), .ZN(n7315) );
  NAND2_X1 U8479 ( .A1(n7316), .A2(n7315), .ZN(n7317) );
  NAND2_X1 U8480 ( .A1(n7472), .A2(n7317), .ZN(n8372) );
  INV_X1 U8481 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7318) );
  OAI222_X1 U8482 ( .A1(n10451), .A2(n8372), .B1(n9653), .B2(P1_U3084), .C1(
        n7318), .C2(n10455), .ZN(P1_U3332) );
  NAND2_X1 U8483 ( .A1(n7320), .A2(n7319), .ZN(n7325) );
  INV_X1 U8484 ( .A(n7321), .ZN(n7323) );
  NAND2_X1 U8485 ( .A1(n7323), .A2(n7322), .ZN(n7324) );
  NAND2_X1 U8486 ( .A1(n7410), .A2(n9427), .ZN(n7327) );
  AOI22_X1 U8487 ( .A1(n8442), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n8352), .B2(
        n10544), .ZN(n7326) );
  NAND2_X1 U8488 ( .A1(n7327), .A2(n7326), .ZN(n7634) );
  OR2_X1 U8489 ( .A1(n10756), .A2(n9287), .ZN(n7328) );
  NAND2_X1 U8490 ( .A1(n7329), .A2(n7328), .ZN(n7330) );
  XNOR2_X1 U8491 ( .A(n7330), .B(n9208), .ZN(n7489) );
  NOR2_X1 U8492 ( .A1(n10756), .A2(n9286), .ZN(n7331) );
  AOI21_X1 U8493 ( .B1(n7634), .B2(n9235), .A(n7331), .ZN(n7488) );
  XNOR2_X1 U8494 ( .A(n7489), .B(n7488), .ZN(n7332) );
  XNOR2_X1 U8495 ( .A(n7490), .B(n7332), .ZN(n7336) );
  AOI22_X1 U8496 ( .A1(n9381), .A2(n9670), .B1(n9347), .B2(n7402), .ZN(n7333)
         );
  NAND2_X1 U8497 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3084), .ZN(n10547) );
  OAI211_X1 U8498 ( .C1(n7651), .C2(n9388), .A(n7333), .B(n10547), .ZN(n7334)
         );
  AOI21_X1 U8499 ( .B1(n7634), .B2(n9407), .A(n7334), .ZN(n7335) );
  OAI21_X1 U8500 ( .B1(n7336), .B2(n9410), .A(n7335), .ZN(P1_U3215) );
  AND2_X1 U8501 ( .A1(n10681), .A2(n8052), .ZN(n7339) );
  INV_X1 U8502 ( .A(n8702), .ZN(n7366) );
  NAND2_X1 U8503 ( .A1(n7366), .A2(n8560), .ZN(n8055) );
  NAND2_X1 U8504 ( .A1(n10692), .A2(n8702), .ZN(n8056) );
  NAND2_X1 U8505 ( .A1(n8055), .A2(n8056), .ZN(n8268) );
  AND2_X1 U8506 ( .A1(n8268), .A2(n8052), .ZN(n7337) );
  OAI21_X1 U8507 ( .B1(n7339), .B2(n8268), .A(n7368), .ZN(n10696) );
  NAND2_X1 U8508 ( .A1(n7340), .A2(n10692), .ZN(n9026) );
  OR2_X1 U8509 ( .A1(n7340), .A2(n10692), .ZN(n7341) );
  NAND2_X1 U8510 ( .A1(n9026), .A2(n7341), .ZN(n10693) );
  AOI22_X1 U8511 ( .A1(n9035), .A2(n8560), .B1(n8561), .B2(n10801), .ZN(n7342)
         );
  OAI21_X1 U8512 ( .B1(n10693), .B2(n8793), .A(n7342), .ZN(n7347) );
  INV_X1 U8513 ( .A(n8701), .ZN(n8556) );
  AND2_X1 U8514 ( .A1(n8703), .A2(n10677), .ZN(n7343) );
  XNOR2_X1 U8515 ( .A(n7380), .B(n8268), .ZN(n7345) );
  OAI222_X1 U8516 ( .A1(n8808), .A2(n8556), .B1(n7345), .B2(n10797), .C1(n8806), .C2(n8557), .ZN(n10694) );
  MUX2_X1 U8517 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10694), .S(n10811), .Z(n7346) );
  AOI211_X1 U8518 ( .C1(n9033), .C2(n10696), .A(n7347), .B(n7346), .ZN(n7348)
         );
  INV_X1 U8519 ( .A(n7348), .ZN(P2_U3289) );
  INV_X1 U8520 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8164) );
  OAI222_X1 U8521 ( .A1(P2_U3152), .A2(n8314), .B1(n9153), .B2(n8372), .C1(
        n8164), .C2(n9151), .ZN(P2_U3337) );
  INV_X1 U8522 ( .A(n7349), .ZN(n7351) );
  AOI21_X1 U8523 ( .B1(n7351), .B2(n7756), .A(n7350), .ZN(n7354) );
  NAND2_X1 U8524 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n8330), .ZN(n7352) );
  OAI21_X1 U8525 ( .B1(n8330), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7352), .ZN(
        n7353) );
  NOR2_X1 U8526 ( .A1(n7354), .A2(n7353), .ZN(n7480) );
  AOI211_X1 U8527 ( .C1(n7354), .C2(n7353), .A(n7480), .B(n7688), .ZN(n7365)
         );
  INV_X1 U8528 ( .A(n7355), .ZN(n7357) );
  AOI21_X1 U8529 ( .B1(n7357), .B2(n7756), .A(n7356), .ZN(n7360) );
  INV_X1 U8530 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n10895) );
  NOR2_X1 U8531 ( .A1(n8330), .A2(n10895), .ZN(n7358) );
  AOI21_X1 U8532 ( .B1(n8330), .B2(n10895), .A(n7358), .ZN(n7359) );
  NOR2_X1 U8533 ( .A1(n7360), .A2(n7359), .ZN(n7476) );
  AOI211_X1 U8534 ( .C1(n7360), .C2(n7359), .A(n7476), .B(n10621), .ZN(n7364)
         );
  INV_X1 U8535 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7362) );
  NAND2_X1 U8536 ( .A1(n10566), .A2(n8330), .ZN(n7361) );
  NAND2_X1 U8537 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9327) );
  OAI211_X1 U8538 ( .C1(n10626), .C2(n7362), .A(n7361), .B(n9327), .ZN(n7363)
         );
  OR3_X1 U8539 ( .A1(n7365), .A2(n7364), .A3(n7363), .ZN(P1_U3257) );
  NAND2_X1 U8540 ( .A1(n7366), .A2(n10692), .ZN(n7367) );
  NAND2_X1 U8541 ( .A1(n10702), .A2(n8701), .ZN(n8059) );
  NAND2_X1 U8542 ( .A1(n9034), .A2(n8556), .ZN(n8058) );
  NAND2_X1 U8543 ( .A1(n9034), .A2(n8701), .ZN(n7369) );
  AOI22_X1 U8544 ( .A1(n8135), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8134), .B2(
        n7371), .ZN(n7372) );
  INV_X1 U8545 ( .A(n8700), .ZN(n7467) );
  OR2_X1 U8546 ( .A1(n7441), .A2(n7467), .ZN(n8064) );
  NAND2_X1 U8547 ( .A1(n7441), .A2(n7467), .ZN(n8068) );
  NAND2_X1 U8548 ( .A1(n8064), .A2(n8068), .ZN(n8266) );
  OAI21_X1 U8549 ( .B1(n5134), .B2(n8266), .A(n7409), .ZN(n10739) );
  INV_X1 U8550 ( .A(n10739), .ZN(n7391) );
  NAND2_X1 U8551 ( .A1(n7373), .A2(n10080), .ZN(n7374) );
  AND2_X1 U8552 ( .A1(n7539), .A2(n7374), .ZN(n7464) );
  NAND2_X1 U8553 ( .A1(n8191), .A2(n7464), .ZN(n7379) );
  NAND2_X1 U8554 ( .A1(n8192), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7378) );
  INV_X1 U8555 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7375) );
  OR2_X1 U8556 ( .A1(n8169), .A2(n7375), .ZN(n7377) );
  OR2_X1 U8557 ( .A1(n8171), .A2(n6390), .ZN(n7376) );
  NAND4_X1 U8558 ( .A1(n7379), .A2(n7378), .A3(n7377), .A4(n7376), .ZN(n8699)
         );
  AOI22_X1 U8559 ( .A1(n9012), .A2(n8701), .B1(n8699), .B2(n9014), .ZN(n7385)
         );
  NAND2_X1 U8560 ( .A1(n7380), .A2(n5250), .ZN(n7381) );
  OAI211_X1 U8561 ( .C1(n5136), .C2(n7383), .A(n9017), .B(n7418), .ZN(n7384)
         );
  OAI211_X1 U8562 ( .C1(n7391), .C2(n8979), .A(n7385), .B(n7384), .ZN(n10737)
         );
  NAND2_X1 U8563 ( .A1(n10737), .A2(n10811), .ZN(n7390) );
  XNOR2_X1 U8564 ( .A(n9027), .B(n7441), .ZN(n10736) );
  INV_X1 U8565 ( .A(n10736), .ZN(n7388) );
  INV_X1 U8566 ( .A(n7441), .ZN(n10735) );
  AOI22_X1 U8567 ( .A1(n10813), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7450), .B2(
        n10801), .ZN(n7386) );
  OAI21_X1 U8568 ( .B1(n10735), .B2(n9008), .A(n7386), .ZN(n7387) );
  AOI21_X1 U8569 ( .B1(n7388), .B2(n9020), .A(n7387), .ZN(n7389) );
  OAI211_X1 U8570 ( .C1(n7391), .C2(n8987), .A(n7390), .B(n7389), .ZN(P2_U3287) );
  AND2_X1 U8571 ( .A1(n10783), .A2(n10822), .ZN(n7392) );
  OR2_X1 U8572 ( .A1(n10773), .A2(n7392), .ZN(n9926) );
  NAND2_X1 U8573 ( .A1(n7393), .A2(n9671), .ZN(n7394) );
  AND2_X1 U8574 ( .A1(n7400), .A2(n9670), .ZN(n7396) );
  OR2_X1 U8575 ( .A1(n7634), .A2(n10756), .ZN(n9515) );
  NAND2_X1 U8576 ( .A1(n7634), .A2(n10756), .ZN(n9516) );
  XNOR2_X1 U8577 ( .A(n7633), .B(n5067), .ZN(n7456) );
  INV_X1 U8578 ( .A(n7400), .ZN(n10730) );
  AND2_X1 U8579 ( .A1(n10730), .A2(n9670), .ZN(n9513) );
  NAND2_X1 U8580 ( .A1(n7400), .A2(n7397), .ZN(n9504) );
  OAI21_X1 U8581 ( .B1(n5067), .B2(n7398), .A(n7648), .ZN(n7399) );
  AOI222_X1 U8582 ( .A1(n10758), .A2(n7399), .B1(n7637), .B2(n9910), .C1(n9670), .C2(n9912), .ZN(n7455) );
  INV_X1 U8583 ( .A(n7455), .ZN(n7407) );
  INV_X1 U8584 ( .A(n7634), .ZN(n7405) );
  OAI21_X1 U8585 ( .B1(n10709), .B2(n7405), .A(n10878), .ZN(n7401) );
  AND2_X1 U8586 ( .A1(n10709), .A2(n7405), .ZN(n10762) );
  NOR2_X1 U8587 ( .A1(n7401), .A2(n10762), .ZN(n7453) );
  INV_X1 U8588 ( .A(n9924), .ZN(n7647) );
  NAND2_X1 U8589 ( .A1(n7453), .A2(n7647), .ZN(n7404) );
  AOI22_X1 U8590 ( .A1(n10778), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7402), .B2(
        n10776), .ZN(n7403) );
  OAI211_X1 U8591 ( .C1(n7405), .C2(n10780), .A(n7404), .B(n7403), .ZN(n7406)
         );
  AOI21_X1 U8592 ( .B1(n7407), .B2(n10783), .A(n7406), .ZN(n7408) );
  OAI21_X1 U8593 ( .B1(n9885), .B2(n7456), .A(n7408), .ZN(P1_U3281) );
  NAND2_X1 U8594 ( .A1(n7410), .A2(n8211), .ZN(n7413) );
  AOI22_X1 U8595 ( .A1(n8135), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8134), .B2(
        n7411), .ZN(n7412) );
  NAND2_X1 U8596 ( .A1(n7413), .A2(n7412), .ZN(n7579) );
  INV_X1 U8597 ( .A(n8699), .ZN(n7414) );
  OR2_X1 U8598 ( .A1(n7579), .A2(n7414), .ZN(n8070) );
  NAND2_X1 U8599 ( .A1(n7579), .A2(n7414), .ZN(n8067) );
  INV_X1 U8600 ( .A(n7419), .ZN(n7415) );
  NAND2_X1 U8601 ( .A1(n7416), .A2(n7419), .ZN(n7417) );
  XNOR2_X1 U8602 ( .A(n7571), .B(n7415), .ZN(n7427) );
  NAND2_X1 U8603 ( .A1(n8192), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7425) );
  XNOR2_X1 U8604 ( .A(n7539), .B(P2_REG3_REG_11__SCAN_IN), .ZN(n10802) );
  NAND2_X1 U8605 ( .A1(n6516), .A2(n10802), .ZN(n7424) );
  INV_X1 U8606 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7420) );
  OR2_X1 U8607 ( .A1(n8169), .A2(n7420), .ZN(n7423) );
  OR2_X1 U8608 ( .A1(n8171), .A2(n7421), .ZN(n7422) );
  NAND4_X1 U8609 ( .A1(n7425), .A2(n7424), .A3(n7423), .A4(n7422), .ZN(n8698)
         );
  OAI22_X1 U8610 ( .A1(n7716), .A2(n8808), .B1(n7467), .B2(n8806), .ZN(n7426)
         );
  AOI21_X1 U8611 ( .B1(n7427), .B2(n9017), .A(n7426), .ZN(n7428) );
  OAI21_X1 U8612 ( .B1(n10741), .B2(n8979), .A(n7428), .ZN(n10744) );
  NAND2_X1 U8613 ( .A1(n10744), .A2(n10811), .ZN(n7435) );
  INV_X1 U8614 ( .A(n7579), .ZN(n10742) );
  NOR2_X1 U8615 ( .A1(n7429), .A2(n10742), .ZN(n7430) );
  OR2_X1 U8616 ( .A1(n10793), .A2(n7430), .ZN(n10743) );
  INV_X1 U8617 ( .A(n10743), .ZN(n7433) );
  AOI22_X1 U8618 ( .A1(n10813), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n7464), .B2(
        n10801), .ZN(n7431) );
  OAI21_X1 U8619 ( .B1(n10742), .B2(n9008), .A(n7431), .ZN(n7432) );
  AOI21_X1 U8620 ( .B1(n7433), .B2(n9020), .A(n7432), .ZN(n7434) );
  OAI211_X1 U8621 ( .C1(n10741), .C2(n8987), .A(n7435), .B(n7434), .ZN(
        P2_U3286) );
  INV_X1 U8622 ( .A(n7436), .ZN(n7437) );
  XNOR2_X1 U8623 ( .A(n7441), .B(n6764), .ZN(n7443) );
  AND2_X1 U8624 ( .A1(n8700), .A2(n8531), .ZN(n7442) );
  NOR2_X1 U8625 ( .A1(n7443), .A2(n7442), .ZN(n7461) );
  AOI21_X1 U8626 ( .B1(n7443), .B2(n7442), .A(n7461), .ZN(n7444) );
  OAI21_X1 U8627 ( .B1(n7445), .B2(n7444), .A(n7463), .ZN(n7446) );
  NAND2_X1 U8628 ( .A1(n7446), .A2(n8683), .ZN(n7452) );
  NAND2_X1 U8629 ( .A1(n8685), .A2(n8699), .ZN(n7448) );
  OAI211_X1 U8630 ( .C1(n8556), .C2(n8688), .A(n7448), .B(n7447), .ZN(n7449)
         );
  AOI21_X1 U8631 ( .B1(n7450), .B2(n8690), .A(n7449), .ZN(n7451) );
  OAI211_X1 U8632 ( .C1(n10735), .C2(n8693), .A(n7452), .B(n7451), .ZN(
        P2_U3233) );
  INV_X1 U8633 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7458) );
  AOI21_X1 U8634 ( .B1(n10877), .B2(n7634), .A(n7453), .ZN(n7454) );
  OAI211_X1 U8635 ( .C1(n10831), .C2(n7456), .A(n7455), .B(n7454), .ZN(n7459)
         );
  NAND2_X1 U8636 ( .A1(n7459), .A2(n5045), .ZN(n7457) );
  OAI21_X1 U8637 ( .B1(n5045), .B2(n7458), .A(n7457), .ZN(P1_U3484) );
  NAND2_X1 U8638 ( .A1(n7459), .A2(n10722), .ZN(n7460) );
  OAI21_X1 U8639 ( .B1(n10722), .B2(n6103), .A(n7460), .ZN(P1_U3533) );
  INV_X1 U8640 ( .A(n7461), .ZN(n7462) );
  XNOR2_X1 U8641 ( .A(n7579), .B(n6765), .ZN(n7531) );
  NAND2_X1 U8642 ( .A1(n8699), .A2(n8531), .ZN(n7530) );
  XNOR2_X1 U8643 ( .A(n7531), .B(n7530), .ZN(n7532) );
  XNOR2_X1 U8644 ( .A(n7533), .B(n7532), .ZN(n7470) );
  AOI22_X1 U8645 ( .A1(n8685), .A2(n8698), .B1(P2_REG3_REG_10__SCAN_IN), .B2(
        P2_U3152), .ZN(n7466) );
  NAND2_X1 U8646 ( .A1(n8690), .A2(n7464), .ZN(n7465) );
  OAI211_X1 U8647 ( .C1(n7467), .C2(n8688), .A(n7466), .B(n7465), .ZN(n7468)
         );
  AOI21_X1 U8648 ( .B1(n7579), .B2(n8651), .A(n7468), .ZN(n7469) );
  OAI21_X1 U8649 ( .B1(n7470), .B2(n8667), .A(n7469), .ZN(P2_U3219) );
  MUX2_X1 U8650 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n7958), .Z(n7656) );
  XNOR2_X1 U8651 ( .A(n7656), .B(SI_22_), .ZN(n7654) );
  XNOR2_X1 U8652 ( .A(n7655), .B(n7654), .ZN(n8385) );
  INV_X1 U8653 ( .A(n8385), .ZN(n7474) );
  OAI222_X1 U8654 ( .A1(n8252), .A2(P2_U3152), .B1(n9153), .B2(n7474), .C1(
        n9151), .C2(n7473), .ZN(P2_U3336) );
  INV_X1 U8655 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7475) );
  OAI222_X1 U8656 ( .A1(n10455), .A2(n7475), .B1(n10451), .B2(n7474), .C1(
        P1_U3084), .C2(n9596), .ZN(P1_U3331) );
  AOI21_X1 U8657 ( .B1(n8330), .B2(P1_REG1_REG_16__SCAN_IN), .A(n7476), .ZN(
        n7478) );
  XNOR2_X1 U8658 ( .A(n8335), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n7477) );
  NOR2_X1 U8659 ( .A1(n7478), .A2(n7477), .ZN(n7670) );
  AOI211_X1 U8660 ( .C1(n7478), .C2(n7477), .A(n7670), .B(n10621), .ZN(n7479)
         );
  AOI21_X1 U8661 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(n10550), .A(n7479), .ZN(
        n7487) );
  NAND2_X1 U8662 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9334) );
  INV_X1 U8663 ( .A(n9334), .ZN(n7485) );
  AOI21_X1 U8664 ( .B1(n8330), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7480), .ZN(
        n7483) );
  NAND2_X1 U8665 ( .A1(n8335), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7481) );
  OAI21_X1 U8666 ( .B1(n8335), .B2(P1_REG2_REG_17__SCAN_IN), .A(n7481), .ZN(
        n7482) );
  NOR2_X1 U8667 ( .A1(n7483), .A2(n7482), .ZN(n7665) );
  AOI211_X1 U8668 ( .C1(n7483), .C2(n7482), .A(n7665), .B(n7688), .ZN(n7484)
         );
  AOI211_X1 U8669 ( .C1(n8335), .C2(n10566), .A(n7485), .B(n7484), .ZN(n7486)
         );
  NAND2_X1 U8670 ( .A1(n7487), .A2(n7486), .ZN(P1_U3258) );
  NAND2_X1 U8671 ( .A1(n7534), .A2(n9427), .ZN(n7493) );
  AOI22_X1 U8672 ( .A1(n8442), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n8352), .B2(
        n7491), .ZN(n7492) );
  NAND2_X1 U8673 ( .A1(n7493), .A2(n7492), .ZN(n7641) );
  OR2_X1 U8674 ( .A1(n7651), .A2(n9287), .ZN(n7494) );
  NAND2_X1 U8675 ( .A1(n7495), .A2(n7494), .ZN(n7496) );
  XNOR2_X1 U8676 ( .A(n7496), .B(n9243), .ZN(n7512) );
  NOR2_X1 U8677 ( .A1(n7651), .A2(n9286), .ZN(n7497) );
  AOI21_X1 U8678 ( .B1(n7641), .B2(n9235), .A(n7497), .ZN(n7513) );
  XNOR2_X1 U8679 ( .A(n7512), .B(n7513), .ZN(n7510) );
  XOR2_X1 U8680 ( .A(n7511), .B(n7510), .Z(n7509) );
  NAND2_X1 U8681 ( .A1(n6031), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7504) );
  OR2_X1 U8682 ( .A1(n7498), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7500) );
  AND2_X1 U8683 ( .A1(n7500), .A2(n7499), .ZN(n7643) );
  NAND2_X1 U8684 ( .A1(n6931), .A2(n7643), .ZN(n7503) );
  NAND2_X1 U8685 ( .A1(n6933), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7502) );
  NAND2_X1 U8686 ( .A1(n9423), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7501) );
  INV_X1 U8687 ( .A(n10756), .ZN(n9669) );
  AOI22_X1 U8688 ( .A1(n9381), .A2(n9669), .B1(n9347), .B2(n10777), .ZN(n7506)
         );
  OAI211_X1 U8689 ( .C1(n10754), .C2(n9388), .A(n7506), .B(n7505), .ZN(n7507)
         );
  AOI21_X1 U8690 ( .B1(n7641), .B2(n9407), .A(n7507), .ZN(n7508) );
  OAI21_X1 U8691 ( .B1(n7509), .B2(n9410), .A(n7508), .ZN(P1_U3234) );
  INV_X1 U8692 ( .A(n7512), .ZN(n7514) );
  NAND2_X1 U8693 ( .A1(n7514), .A2(n7513), .ZN(n7515) );
  NAND2_X1 U8694 ( .A1(n7516), .A2(n7515), .ZN(n7730) );
  OR2_X1 U8695 ( .A1(n7573), .A2(n6231), .ZN(n7519) );
  AOI22_X1 U8696 ( .A1(n8442), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n8352), .B2(
        n7517), .ZN(n7518) );
  OR2_X1 U8697 ( .A1(n10754), .A2(n9287), .ZN(n7520) );
  NAND2_X1 U8698 ( .A1(n7521), .A2(n7520), .ZN(n7522) );
  XNOR2_X1 U8699 ( .A(n7522), .B(n9208), .ZN(n7724) );
  NOR2_X1 U8700 ( .A1(n10754), .A2(n9286), .ZN(n7523) );
  AOI21_X1 U8701 ( .B1(n10815), .B2(n9235), .A(n7523), .ZN(n7725) );
  XNOR2_X1 U8702 ( .A(n7724), .B(n7725), .ZN(n7524) );
  XNOR2_X1 U8703 ( .A(n7730), .B(n7524), .ZN(n7529) );
  AOI22_X1 U8704 ( .A1(n9381), .A2(n7637), .B1(n9347), .B2(n7643), .ZN(n7526)
         );
  OAI211_X1 U8705 ( .C1(n9260), .C2(n9388), .A(n7526), .B(n7525), .ZN(n7527)
         );
  AOI21_X1 U8706 ( .B1(n10815), .B2(n9407), .A(n7527), .ZN(n7528) );
  OAI21_X1 U8707 ( .B1(n7529), .B2(n9410), .A(n7528), .ZN(P1_U3222) );
  NAND2_X1 U8708 ( .A1(n8698), .A2(n8531), .ZN(n7706) );
  NAND2_X1 U8709 ( .A1(n7534), .A2(n8211), .ZN(n7537) );
  AOI22_X1 U8710 ( .A1(n8135), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8134), .B2(
        n7535), .ZN(n7536) );
  NAND2_X1 U8711 ( .A1(n7537), .A2(n7536), .ZN(n10804) );
  XNOR2_X1 U8712 ( .A(n10804), .B(n6765), .ZN(n7705) );
  XOR2_X1 U8713 ( .A(n7706), .B(n7705), .Z(n7709) );
  XNOR2_X1 U8714 ( .A(n7710), .B(n7709), .ZN(n7551) );
  NAND2_X1 U8715 ( .A1(n8192), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7546) );
  INV_X1 U8716 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10304) );
  OAI21_X1 U8717 ( .B1(n7539), .B2(n7538), .A(n10304), .ZN(n7540) );
  AND2_X1 U8718 ( .A1(n7564), .A2(n7540), .ZN(n7718) );
  NAND2_X1 U8719 ( .A1(n8191), .A2(n7718), .ZN(n7545) );
  INV_X1 U8720 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7541) );
  OR2_X1 U8721 ( .A1(n8169), .A2(n7541), .ZN(n7544) );
  OR2_X1 U8722 ( .A1(n8171), .A2(n7542), .ZN(n7543) );
  NAND4_X1 U8723 ( .A1(n7546), .A2(n7545), .A3(n7544), .A4(n7543), .ZN(n8697)
         );
  AOI22_X1 U8724 ( .A1(n9012), .A2(n8699), .B1(n8697), .B2(n9014), .ZN(n10796)
         );
  NOR2_X1 U8725 ( .A1(n10796), .A2(n8612), .ZN(n7547) );
  AOI211_X1 U8726 ( .C1(n8690), .C2(n10802), .A(n7548), .B(n7547), .ZN(n7550)
         );
  NAND2_X1 U8727 ( .A1(n10804), .A2(n8651), .ZN(n7549) );
  OAI211_X1 U8728 ( .C1(n7551), .C2(n8667), .A(n7550), .B(n7549), .ZN(P2_U3238) );
  XNOR2_X1 U8729 ( .A(n7836), .B(n8086), .ZN(n7554) );
  INV_X1 U8730 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7553) );
  NAND2_X1 U8731 ( .A1(n7554), .A2(n7553), .ZN(n7838) );
  OAI21_X1 U8732 ( .B1(n7554), .B2(n7553), .A(n7838), .ZN(n7555) );
  INV_X1 U8733 ( .A(n7555), .ZN(n7563) );
  INV_X1 U8734 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7556) );
  NAND2_X1 U8735 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8686) );
  OAI21_X1 U8736 ( .B1(n10594), .B2(n7556), .A(n8686), .ZN(n7557) );
  AOI21_X1 U8737 ( .B1(n8086), .B2(n10613), .A(n7557), .ZN(n7562) );
  AOI21_X1 U8738 ( .B1(n7559), .B2(n10869), .A(n7558), .ZN(n7829) );
  XNOR2_X1 U8739 ( .A(n7829), .B(n7837), .ZN(n7560) );
  NAND2_X1 U8740 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n7560), .ZN(n7830) );
  OAI211_X1 U8741 ( .C1(n7560), .C2(P2_REG1_REG_15__SCAN_IN), .A(n10615), .B(
        n7830), .ZN(n7561) );
  OAI211_X1 U8742 ( .C1(n7563), .C2(n10607), .A(n7562), .B(n7561), .ZN(
        P2_U3260) );
  NAND2_X1 U8743 ( .A1(n8192), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7570) );
  NAND2_X1 U8744 ( .A1(n7564), .A2(n10319), .ZN(n7565) );
  AND2_X1 U8745 ( .A1(n7873), .A2(n7565), .ZN(n7860) );
  NAND2_X1 U8746 ( .A1(n8191), .A2(n7860), .ZN(n7569) );
  INV_X1 U8747 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7566) );
  OR2_X1 U8748 ( .A1(n8169), .A2(n7566), .ZN(n7568) );
  OR2_X1 U8749 ( .A1(n8171), .A2(n7156), .ZN(n7567) );
  NAND4_X1 U8750 ( .A1(n7570), .A2(n7569), .A3(n7568), .A4(n7567), .ZN(n8696)
         );
  OR2_X1 U8751 ( .A1(n10804), .A2(n7716), .ZN(n8071) );
  INV_X1 U8752 ( .A(n8071), .ZN(n7572) );
  NAND2_X1 U8753 ( .A1(n10804), .A2(n7716), .ZN(n8066) );
  OAI21_X1 U8754 ( .B1(n7811), .B2(n7572), .A(n8066), .ZN(n7577) );
  OR2_X1 U8755 ( .A1(n7573), .A2(n6702), .ZN(n7576) );
  AOI22_X1 U8756 ( .A1(n8135), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8134), .B2(
        n7574), .ZN(n7575) );
  INV_X1 U8757 ( .A(n8697), .ZN(n7858) );
  OR2_X1 U8758 ( .A1(n7821), .A2(n7858), .ZN(n7809) );
  NAND2_X1 U8759 ( .A1(n7821), .A2(n7858), .ZN(n8076) );
  XNOR2_X1 U8760 ( .A(n7577), .B(n8255), .ZN(n7578) );
  OAI222_X1 U8761 ( .A1(n8808), .A2(n7903), .B1(n7578), .B2(n10797), .C1(n8806), .C2(n7716), .ZN(n10827) );
  INV_X1 U8762 ( .A(n10827), .ZN(n7589) );
  NAND2_X1 U8763 ( .A1(n7579), .A2(n8699), .ZN(n7580) );
  NAND2_X1 U8764 ( .A1(n8071), .A2(n8066), .ZN(n10788) );
  NAND2_X1 U8765 ( .A1(n10804), .A2(n8698), .ZN(n7581) );
  OAI21_X1 U8766 ( .B1(n5135), .B2(n8255), .A(n7582), .ZN(n10829) );
  INV_X1 U8767 ( .A(n10804), .ZN(n10794) );
  NAND2_X1 U8768 ( .A1(n10791), .A2(n7821), .ZN(n7583) );
  NAND2_X1 U8769 ( .A1(n7817), .A2(n7583), .ZN(n10826) );
  INV_X1 U8770 ( .A(n7718), .ZN(n7584) );
  OAI22_X1 U8771 ( .A1(n10811), .A2(n7542), .B1(n7584), .B2(n8981), .ZN(n7585)
         );
  AOI21_X1 U8772 ( .B1(n7821), .B2(n9035), .A(n7585), .ZN(n7586) );
  OAI21_X1 U8773 ( .B1(n10826), .B2(n8793), .A(n7586), .ZN(n7587) );
  AOI21_X1 U8774 ( .B1(n10829), .B2(n9033), .A(n7587), .ZN(n7588) );
  OAI21_X1 U8775 ( .B1(n7589), .B2(n10813), .A(n7588), .ZN(P2_U3284) );
  NOR2_X1 U8776 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7628) );
  NOR2_X1 U8777 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7626) );
  NOR2_X1 U8778 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7624) );
  NOR2_X1 U8779 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7622) );
  NOR2_X1 U8780 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7619) );
  NOR2_X1 U8781 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7616) );
  NAND2_X1 U8782 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7614) );
  XNOR2_X1 U8783 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n7590), .ZN(n10485) );
  NAND2_X1 U8784 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7612) );
  XOR2_X1 U8785 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .Z(n10483) );
  NOR2_X1 U8786 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7596) );
  XNOR2_X1 U8787 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10474) );
  NAND2_X1 U8788 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7594) );
  XOR2_X1 U8789 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(P1_ADDR_REG_3__SCAN_IN), .Z(
        n10472) );
  NAND2_X1 U8790 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7592) );
  XOR2_X1 U8791 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10470) );
  AOI21_X1 U8792 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10465) );
  INV_X1 U8793 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10593) );
  NAND3_X1 U8794 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10467) );
  OAI21_X1 U8795 ( .B1(n10465), .B2(n10593), .A(n10467), .ZN(n10469) );
  NAND2_X1 U8796 ( .A1(n10470), .A2(n10469), .ZN(n7591) );
  NAND2_X1 U8797 ( .A1(n7592), .A2(n7591), .ZN(n10471) );
  NAND2_X1 U8798 ( .A1(n10472), .A2(n10471), .ZN(n7593) );
  NAND2_X1 U8799 ( .A1(n7594), .A2(n7593), .ZN(n10473) );
  NOR2_X1 U8800 ( .A1(n10474), .A2(n10473), .ZN(n7595) );
  NOR2_X1 U8801 ( .A1(n7596), .A2(n7595), .ZN(n7597) );
  NOR2_X1 U8802 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7597), .ZN(n10476) );
  AND2_X1 U8803 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7597), .ZN(n10475) );
  NOR2_X1 U8804 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10475), .ZN(n7598) );
  NAND2_X1 U8805 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n7599), .ZN(n7601) );
  XOR2_X1 U8806 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n7599), .Z(n10478) );
  NAND2_X1 U8807 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10478), .ZN(n7600) );
  NAND2_X1 U8808 ( .A1(n7601), .A2(n7600), .ZN(n7602) );
  NAND2_X1 U8809 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7602), .ZN(n7604) );
  XOR2_X1 U8810 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7602), .Z(n10479) );
  NAND2_X1 U8811 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10479), .ZN(n7603) );
  NAND2_X1 U8812 ( .A1(n7604), .A2(n7603), .ZN(n7605) );
  NAND2_X1 U8813 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7605), .ZN(n7607) );
  XOR2_X1 U8814 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7605), .Z(n10480) );
  NAND2_X1 U8815 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10480), .ZN(n7606) );
  NAND2_X1 U8816 ( .A1(n7607), .A2(n7606), .ZN(n7608) );
  NAND2_X1 U8817 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n7608), .ZN(n7610) );
  XOR2_X1 U8818 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n7608), .Z(n10481) );
  NAND2_X1 U8819 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10481), .ZN(n7609) );
  NAND2_X1 U8820 ( .A1(n7610), .A2(n7609), .ZN(n10482) );
  NAND2_X1 U8821 ( .A1(n10483), .A2(n10482), .ZN(n7611) );
  NAND2_X1 U8822 ( .A1(n7612), .A2(n7611), .ZN(n10484) );
  NAND2_X1 U8823 ( .A1(n10485), .A2(n10484), .ZN(n7613) );
  NAND2_X1 U8824 ( .A1(n7614), .A2(n7613), .ZN(n10487) );
  XNOR2_X1 U8825 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10486) );
  XOR2_X1 U8826 ( .A(n7617), .B(P1_ADDR_REG_13__SCAN_IN), .Z(n10488) );
  XOR2_X1 U8827 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(n7620), .Z(n10490) );
  NOR2_X1 U8828 ( .A1(n10491), .A2(n10490), .ZN(n7621) );
  NOR2_X1 U8829 ( .A1(n7622), .A2(n7621), .ZN(n10493) );
  XNOR2_X1 U8830 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10492) );
  NOR2_X1 U8831 ( .A1(n10493), .A2(n10492), .ZN(n7623) );
  NOR2_X1 U8832 ( .A1(n7624), .A2(n7623), .ZN(n10495) );
  XNOR2_X1 U8833 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10494) );
  NOR2_X1 U8834 ( .A1(n10495), .A2(n10494), .ZN(n7625) );
  NOR2_X1 U8835 ( .A1(n7626), .A2(n7625), .ZN(n10497) );
  XNOR2_X1 U8836 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10496) );
  NOR2_X1 U8837 ( .A1(n10497), .A2(n10496), .ZN(n7627) );
  NOR2_X1 U8838 ( .A1(n7628), .A2(n7627), .ZN(n7629) );
  AND2_X1 U8839 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n7629), .ZN(n10498) );
  NOR2_X1 U8840 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10498), .ZN(n7630) );
  NOR2_X1 U8841 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n7629), .ZN(n10499) );
  NOR2_X1 U8842 ( .A1(n7630), .A2(n10499), .ZN(n7632) );
  XNOR2_X1 U8843 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7631) );
  XNOR2_X1 U8844 ( .A(n7632), .B(n7631), .ZN(ADD_1071_U4) );
  NAND2_X1 U8845 ( .A1(n10815), .A2(n10754), .ZN(n9530) );
  OR2_X1 U8846 ( .A1(n7634), .A2(n9669), .ZN(n7635) );
  NAND2_X1 U8847 ( .A1(n7636), .A2(n7635), .ZN(n10749) );
  OR2_X1 U8848 ( .A1(n7641), .A2(n7651), .ZN(n9526) );
  NAND2_X1 U8849 ( .A1(n7641), .A2(n7651), .ZN(n9519) );
  NAND2_X1 U8850 ( .A1(n9526), .A2(n9519), .ZN(n10750) );
  OR2_X1 U8851 ( .A1(n7641), .A2(n7637), .ZN(n7638) );
  INV_X1 U8852 ( .A(n7779), .ZN(n7639) );
  AOI21_X1 U8853 ( .B1(n9636), .B2(n7640), .A(n7639), .ZN(n10821) );
  INV_X1 U8854 ( .A(n10821), .ZN(n10818) );
  INV_X1 U8855 ( .A(n7641), .ZN(n10781) );
  NAND2_X1 U8856 ( .A1(n10762), .A2(n10781), .ZN(n10764) );
  XNOR2_X1 U8857 ( .A(n10764), .B(n10815), .ZN(n7642) );
  NOR2_X1 U8858 ( .A1(n7642), .A2(n10833), .ZN(n10814) );
  INV_X1 U8859 ( .A(n10815), .ZN(n7645) );
  AOI22_X1 U8860 ( .A1(n10778), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7643), .B2(
        n10776), .ZN(n7644) );
  OAI21_X1 U8861 ( .B1(n7645), .B2(n10780), .A(n7644), .ZN(n7646) );
  AOI21_X1 U8862 ( .B1(n10814), .B2(n7647), .A(n7646), .ZN(n7653) );
  NAND2_X1 U8863 ( .A1(n7648), .A2(n9516), .ZN(n10752) );
  INV_X1 U8864 ( .A(n9519), .ZN(n7649) );
  XNOR2_X1 U8865 ( .A(n7750), .B(n9636), .ZN(n7650) );
  OAI222_X1 U8866 ( .A1(n10753), .A2(n9260), .B1(n10755), .B2(n7651), .C1(
        n9888), .C2(n7650), .ZN(n10819) );
  NAND2_X1 U8867 ( .A1(n10819), .A2(n10783), .ZN(n7652) );
  OAI211_X1 U8868 ( .C1(n10818), .C2(n9885), .A(n7653), .B(n7652), .ZN(
        P1_U3279) );
  INV_X1 U8869 ( .A(n7656), .ZN(n7657) );
  INV_X1 U8870 ( .A(SI_22_), .ZN(n10031) );
  NAND2_X1 U8871 ( .A1(n7657), .A2(n10031), .ZN(n7658) );
  MUX2_X1 U8872 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n5713), .Z(n7692) );
  XNOR2_X1 U8873 ( .A(n7692), .B(n10236), .ZN(n7690) );
  XNOR2_X1 U8874 ( .A(n7691), .B(n7690), .ZN(n8390) );
  INV_X1 U8875 ( .A(n8390), .ZN(n7662) );
  NAND2_X1 U8876 ( .A1(n7660), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9663) );
  NAND2_X1 U8877 ( .A1(n10445), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7661) );
  OAI211_X1 U8878 ( .C1(n7662), .C2(n10451), .A(n9663), .B(n7661), .ZN(
        P1_U3330) );
  INV_X1 U8879 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7999) );
  NAND2_X1 U8880 ( .A1(n8390), .A2(n7663), .ZN(n7664) );
  OAI211_X1 U8881 ( .C1(n7999), .C2(n9151), .A(n7664), .B(n8327), .ZN(P2_U3335) );
  INV_X1 U8882 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n7676) );
  AND2_X1 U8883 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9380) );
  AOI21_X1 U8884 ( .B1(n8335), .B2(P1_REG2_REG_17__SCAN_IN), .A(n7665), .ZN(
        n7668) );
  NAND2_X1 U8885 ( .A1(n8348), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7666) );
  OAI21_X1 U8886 ( .B1(n8348), .B2(P1_REG2_REG_18__SCAN_IN), .A(n7666), .ZN(
        n7667) );
  NOR2_X1 U8887 ( .A1(n7668), .A2(n7667), .ZN(n7677) );
  AOI211_X1 U8888 ( .C1(n7668), .C2(n7667), .A(n7677), .B(n7688), .ZN(n7669)
         );
  AOI211_X1 U8889 ( .C1(n8348), .C2(n10566), .A(n9380), .B(n7669), .ZN(n7675)
         );
  XOR2_X1 U8890 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n8348), .Z(n7672) );
  AOI21_X1 U8891 ( .B1(n8335), .B2(P1_REG1_REG_17__SCAN_IN), .A(n7670), .ZN(
        n7671) );
  NAND2_X1 U8892 ( .A1(n7671), .A2(n7672), .ZN(n7680) );
  OAI21_X1 U8893 ( .B1(n7672), .B2(n7671), .A(n7680), .ZN(n7673) );
  NAND2_X1 U8894 ( .A1(n7673), .A2(n10573), .ZN(n7674) );
  OAI211_X1 U8895 ( .C1(n10626), .C2(n7676), .A(n7675), .B(n7674), .ZN(
        P1_U3259) );
  AOI21_X1 U8896 ( .B1(n8348), .B2(P1_REG2_REG_18__SCAN_IN), .A(n7677), .ZN(
        n7679) );
  XNOR2_X1 U8897 ( .A(n9760), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n7678) );
  XNOR2_X1 U8898 ( .A(n7679), .B(n7678), .ZN(n7689) );
  OAI21_X1 U8899 ( .B1(n8348), .B2(P1_REG1_REG_18__SCAN_IN), .A(n7680), .ZN(
        n7682) );
  XNOR2_X1 U8900 ( .A(n9812), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n7681) );
  XNOR2_X1 U8901 ( .A(n7682), .B(n7681), .ZN(n7686) );
  NAND2_X1 U8902 ( .A1(n10566), .A2(n9760), .ZN(n7683) );
  NAND2_X1 U8903 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9278) );
  OAI211_X1 U8904 ( .C1(n10626), .C2(n7684), .A(n7683), .B(n9278), .ZN(n7685)
         );
  AOI21_X1 U8905 ( .B1(n10573), .B2(n7686), .A(n7685), .ZN(n7687) );
  OAI21_X1 U8906 ( .B1(n7689), .B2(n7688), .A(n7687), .ZN(P1_U3260) );
  INV_X1 U8907 ( .A(n7692), .ZN(n7693) );
  NAND2_X1 U8908 ( .A1(n7693), .A2(n10236), .ZN(n7694) );
  MUX2_X1 U8909 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n5713), .Z(n7696) );
  NAND2_X1 U8910 ( .A1(n7696), .A2(SI_24_), .ZN(n7886) );
  OAI21_X1 U8911 ( .B1(n7696), .B2(SI_24_), .A(n7886), .ZN(n7697) );
  NAND2_X1 U8912 ( .A1(n7698), .A2(n7697), .ZN(n7699) );
  NAND2_X1 U8913 ( .A1(n7887), .A2(n7699), .ZN(n8404) );
  INV_X1 U8914 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7700) );
  OAI222_X1 U8915 ( .A1(n10451), .A2(n8404), .B1(P1_U3084), .B2(n7701), .C1(
        n7700), .C2(n10455), .ZN(P1_U3329) );
  INV_X1 U8916 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7992) );
  OAI222_X1 U8917 ( .A1(P2_U3152), .A2(n7702), .B1(n9153), .B2(n8404), .C1(
        n7992), .C2(n9151), .ZN(P2_U3334) );
  INV_X1 U8918 ( .A(n7821), .ZN(n10825) );
  XNOR2_X1 U8919 ( .A(n7821), .B(n6764), .ZN(n7704) );
  AND2_X1 U8920 ( .A1(n8697), .A2(n8531), .ZN(n7703) );
  NOR2_X1 U8921 ( .A1(n7704), .A2(n7703), .ZN(n7850) );
  AOI21_X1 U8922 ( .B1(n7704), .B2(n7703), .A(n7850), .ZN(n7712) );
  INV_X1 U8923 ( .A(n7705), .ZN(n7708) );
  INV_X1 U8924 ( .A(n7706), .ZN(n7707) );
  OAI21_X1 U8925 ( .B1(n7712), .B2(n7711), .A(n7852), .ZN(n7713) );
  NAND2_X1 U8926 ( .A1(n7713), .A2(n8683), .ZN(n7720) );
  NAND2_X1 U8927 ( .A1(n8685), .A2(n8696), .ZN(n7715) );
  OAI211_X1 U8928 ( .C1(n7716), .C2(n8688), .A(n7715), .B(n7714), .ZN(n7717)
         );
  AOI21_X1 U8929 ( .B1(n7718), .B2(n8690), .A(n7717), .ZN(n7719) );
  OAI211_X1 U8930 ( .C1(n10825), .C2(n8693), .A(n7720), .B(n7719), .ZN(
        P2_U3226) );
  NAND2_X1 U8931 ( .A1(n7812), .A2(n9427), .ZN(n7723) );
  AOI22_X1 U8932 ( .A1(n8442), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n8352), .B2(
        n7721), .ZN(n7722) );
  INV_X1 U8933 ( .A(n7780), .ZN(n10832) );
  AND2_X1 U8934 ( .A1(n7724), .A2(n7725), .ZN(n7729) );
  INV_X1 U8935 ( .A(n7724), .ZN(n7727) );
  INV_X1 U8936 ( .A(n7725), .ZN(n7726) );
  NAND2_X1 U8937 ( .A1(n7727), .A2(n7726), .ZN(n7728) );
  OR2_X1 U8938 ( .A1(n9260), .A2(n9287), .ZN(n7731) );
  NAND2_X1 U8939 ( .A1(n7732), .A2(n7731), .ZN(n7733) );
  XNOR2_X1 U8940 ( .A(n7733), .B(n9243), .ZN(n7736) );
  NAND2_X1 U8941 ( .A1(n7780), .A2(n9235), .ZN(n7735) );
  OR2_X1 U8942 ( .A1(n9260), .A2(n9286), .ZN(n7734) );
  NAND2_X1 U8943 ( .A1(n7735), .A2(n7734), .ZN(n7737) );
  AND2_X1 U8944 ( .A1(n7736), .A2(n7737), .ZN(n7741) );
  INV_X1 U8945 ( .A(n7736), .ZN(n7739) );
  INV_X1 U8946 ( .A(n7737), .ZN(n7738) );
  NAND2_X1 U8947 ( .A1(n7739), .A2(n7738), .ZN(n9158) );
  OAI21_X1 U8948 ( .B1(n7741), .B2(n5599), .A(n7740), .ZN(n7742) );
  OAI21_X1 U8949 ( .B1(n9159), .B2(n5599), .A(n7742), .ZN(n7743) );
  NAND2_X1 U8950 ( .A1(n7743), .A2(n9376), .ZN(n7748) );
  INV_X1 U8951 ( .A(n7744), .ZN(n7746) );
  OAI22_X1 U8952 ( .A1(n10754), .A2(n9402), .B1(n9401), .B2(n7796), .ZN(n7745)
         );
  AOI211_X1 U8953 ( .C1(n9406), .C2(n7782), .A(n7746), .B(n7745), .ZN(n7747)
         );
  OAI211_X1 U8954 ( .C1(n10832), .C2(n9384), .A(n7748), .B(n7747), .ZN(
        P1_U3232) );
  INV_X1 U8955 ( .A(n9524), .ZN(n7749) );
  OR2_X1 U8956 ( .A1(n7780), .A2(n9260), .ZN(n9528) );
  NAND2_X1 U8957 ( .A1(n7780), .A2(n9260), .ZN(n9905) );
  NAND2_X1 U8958 ( .A1(n7863), .A2(n9427), .ZN(n7753) );
  AOI22_X1 U8959 ( .A1(n8442), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n8352), .B2(
        n7751), .ZN(n7752) );
  NAND2_X1 U8960 ( .A1(n9921), .A2(n9403), .ZN(n9536) );
  NAND2_X1 U8961 ( .A1(n9534), .A2(n9536), .ZN(n9915) );
  INV_X1 U8962 ( .A(n9905), .ZN(n9523) );
  NOR2_X1 U8963 ( .A1(n9915), .A2(n9523), .ZN(n7754) );
  NAND2_X1 U8964 ( .A1(n9906), .A2(n7754), .ZN(n7755) );
  AOI22_X1 U8965 ( .A1(n8442), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8352), .B2(
        n7756), .ZN(n7757) );
  NOR2_X1 U8966 ( .A1(n7759), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7760) );
  OR2_X1 U8967 ( .A1(n7767), .A2(n7760), .ZN(n9400) );
  INV_X1 U8968 ( .A(n9400), .ZN(n7775) );
  NAND2_X1 U8969 ( .A1(n6931), .A2(n7775), .ZN(n7764) );
  NAND2_X1 U8970 ( .A1(n6031), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n7763) );
  NAND2_X1 U8971 ( .A1(n6933), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n7762) );
  NAND2_X1 U8972 ( .A1(n9423), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n7761) );
  OR2_X1 U8973 ( .A1(n10876), .A2(n9887), .ZN(n9541) );
  NAND2_X1 U8974 ( .A1(n10876), .A2(n9887), .ZN(n9542) );
  NAND2_X1 U8975 ( .A1(n9541), .A2(n9542), .ZN(n9639) );
  NAND2_X1 U8976 ( .A1(n7765), .A2(n9639), .ZN(n7766) );
  NAND2_X1 U8977 ( .A1(n8455), .A2(n7766), .ZN(n7774) );
  OR2_X1 U8978 ( .A1(n7767), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7768) );
  AND2_X1 U8979 ( .A1(n8339), .A2(n7768), .ZN(n9896) );
  NAND2_X1 U8980 ( .A1(n6931), .A2(n9896), .ZN(n7772) );
  NAND2_X1 U8981 ( .A1(n6031), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n7771) );
  NAND2_X1 U8982 ( .A1(n6933), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7770) );
  NAND2_X1 U8983 ( .A1(n9423), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n7769) );
  OAI22_X1 U8984 ( .A1(n9336), .A2(n10753), .B1(n9403), .B2(n10755), .ZN(n7773) );
  AOI21_X1 U8985 ( .B1(n7774), .B2(n10758), .A(n7773), .ZN(n10881) );
  OR2_X1 U8986 ( .A1(n10764), .A2(n10815), .ZN(n7793) );
  XNOR2_X1 U8987 ( .A(n9916), .B(n10876), .ZN(n10879) );
  INV_X1 U8988 ( .A(n10876), .ZN(n8466) );
  AOI22_X1 U8989 ( .A1(n10778), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n7775), .B2(
        n10776), .ZN(n7776) );
  OAI21_X1 U8990 ( .B1(n8466), .B2(n10780), .A(n7776), .ZN(n7777) );
  AOI21_X1 U8991 ( .B1(n10772), .B2(n10879), .A(n7777), .ZN(n7786) );
  INV_X1 U8992 ( .A(n10754), .ZN(n9668) );
  NAND2_X1 U8993 ( .A1(n10815), .A2(n9668), .ZN(n7778) );
  OR2_X1 U8994 ( .A1(n7780), .A2(n9913), .ZN(n7781) );
  NOR2_X1 U8995 ( .A1(n9921), .A2(n7782), .ZN(n7783) );
  OR2_X1 U8996 ( .A1(n7784), .A2(n9639), .ZN(n10875) );
  NAND2_X1 U8997 ( .A1(n7784), .A2(n9639), .ZN(n10874) );
  NAND3_X1 U8998 ( .A1(n10875), .A2(n10874), .A3(n9926), .ZN(n7785) );
  OAI211_X1 U8999 ( .C1(n10881), .C2(n10778), .A(n7786), .B(n7785), .ZN(
        P1_U3276) );
  XNOR2_X1 U9000 ( .A(n7787), .B(n7789), .ZN(n10837) );
  INV_X1 U9001 ( .A(n10837), .ZN(n7803) );
  INV_X1 U9002 ( .A(n7788), .ZN(n7791) );
  INV_X1 U9003 ( .A(n7789), .ZN(n9638) );
  INV_X1 U9004 ( .A(n9906), .ZN(n7790) );
  AOI21_X1 U9005 ( .B1(n7791), .B2(n9638), .A(n7790), .ZN(n7792) );
  OAI222_X1 U9006 ( .A1(n10753), .A2(n9403), .B1(n10755), .B2(n10754), .C1(
        n9888), .C2(n7792), .ZN(n10835) );
  INV_X1 U9007 ( .A(n7793), .ZN(n7795) );
  INV_X1 U9008 ( .A(n9918), .ZN(n7794) );
  OAI21_X1 U9009 ( .B1(n10832), .B2(n7795), .A(n7794), .ZN(n10834) );
  NOR2_X1 U9010 ( .A1(n9897), .A2(n7796), .ZN(n7798) );
  NOR2_X1 U9011 ( .A1(n10832), .A2(n10780), .ZN(n7797) );
  AOI211_X1 U9012 ( .C1(n10778), .C2(P1_REG2_REG_13__SCAN_IN), .A(n7798), .B(
        n7797), .ZN(n7799) );
  OAI21_X1 U9013 ( .B1(n7800), .B2(n10834), .A(n7799), .ZN(n7801) );
  AOI21_X1 U9014 ( .B1(n10835), .B2(n10783), .A(n7801), .ZN(n7802) );
  OAI21_X1 U9015 ( .B1(n9885), .B2(n7803), .A(n7802), .ZN(P1_U3278) );
  XNOR2_X1 U9016 ( .A(n7873), .B(P2_REG3_REG_14__SCAN_IN), .ZN(n7905) );
  NAND2_X1 U9017 ( .A1(n8191), .A2(n7905), .ZN(n7808) );
  NAND2_X1 U9018 ( .A1(n8192), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7807) );
  INV_X1 U9019 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7804) );
  OR2_X1 U9020 ( .A1(n8169), .A2(n7804), .ZN(n7806) );
  OR2_X1 U9021 ( .A1(n8171), .A2(n7290), .ZN(n7805) );
  NAND4_X1 U9022 ( .A1(n7808), .A2(n7807), .A3(n7806), .A4(n7805), .ZN(n9013)
         );
  NAND2_X1 U9023 ( .A1(n7809), .A2(n8071), .ZN(n8077) );
  NAND2_X1 U9024 ( .A1(n8076), .A2(n8066), .ZN(n7810) );
  NAND2_X1 U9025 ( .A1(n7810), .A2(n7809), .ZN(n8079) );
  NAND2_X1 U9026 ( .A1(n7812), .A2(n8211), .ZN(n7815) );
  AOI22_X1 U9027 ( .A1(n8135), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8134), .B2(
        n7813), .ZN(n7814) );
  NAND2_X1 U9028 ( .A1(n7815), .A2(n7814), .ZN(n7847) );
  OR2_X1 U9029 ( .A1(n7847), .A2(n7903), .ZN(n8081) );
  NAND2_X1 U9030 ( .A1(n7847), .A2(n7903), .ZN(n8082) );
  NAND2_X1 U9031 ( .A1(n8081), .A2(n8082), .ZN(n7869) );
  XNOR2_X1 U9032 ( .A(n7870), .B(n7869), .ZN(n7816) );
  OAI222_X1 U9033 ( .A1(n8808), .A2(n8761), .B1(n7816), .B2(n10797), .C1(n8806), .C2(n7858), .ZN(n10846) );
  INV_X1 U9034 ( .A(n7847), .ZN(n10843) );
  INV_X1 U9035 ( .A(n7817), .ZN(n7818) );
  OAI21_X1 U9036 ( .B1(n10843), .B2(n7818), .A(n5321), .ZN(n10844) );
  AOI22_X1 U9037 ( .A1(n10813), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7860), .B2(
        n10801), .ZN(n7820) );
  NAND2_X1 U9038 ( .A1(n7847), .A2(n9035), .ZN(n7819) );
  OAI211_X1 U9039 ( .C1(n10844), .C2(n8793), .A(n7820), .B(n7819), .ZN(n7827)
         );
  OR2_X1 U9040 ( .A1(n7821), .A2(n8697), .ZN(n7822) );
  NOR2_X1 U9041 ( .A1(n7824), .A2(n7869), .ZN(n10842) );
  INV_X1 U9042 ( .A(n10847), .ZN(n7825) );
  NOR3_X1 U9043 ( .A1(n10842), .A2(n7825), .A3(n9022), .ZN(n7826) );
  AOI211_X1 U9044 ( .C1(n10811), .C2(n10846), .A(n7827), .B(n7826), .ZN(n7828)
         );
  INV_X1 U9045 ( .A(n7828), .ZN(P2_U3283) );
  NAND2_X1 U9046 ( .A1(n8086), .A2(n7829), .ZN(n7831) );
  NAND2_X1 U9047 ( .A1(n7831), .A2(n7830), .ZN(n7833) );
  XNOR2_X1 U9048 ( .A(n8092), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n7832) );
  NOR2_X1 U9049 ( .A1(n7833), .A2(n7832), .ZN(n7913) );
  AOI21_X1 U9050 ( .B1(n7833), .B2(n7832), .A(n7913), .ZN(n7846) );
  INV_X1 U9051 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10308) );
  NOR2_X1 U9052 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10308), .ZN(n7834) );
  AOI21_X1 U9053 ( .B1(n10606), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n7834), .ZN(
        n7835) );
  INV_X1 U9054 ( .A(n7835), .ZN(n7844) );
  NAND2_X1 U9055 ( .A1(n7837), .A2(n7836), .ZN(n7839) );
  NAND2_X1 U9056 ( .A1(n7839), .A2(n7838), .ZN(n7842) );
  NAND2_X1 U9057 ( .A1(n8092), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7840) );
  OAI21_X1 U9058 ( .B1(n8092), .B2(P2_REG2_REG_16__SCAN_IN), .A(n7840), .ZN(
        n7841) );
  NOR2_X1 U9059 ( .A1(n7842), .A2(n7841), .ZN(n7908) );
  AOI211_X1 U9060 ( .C1(n7842), .C2(n7841), .A(n7908), .B(n10607), .ZN(n7843)
         );
  AOI211_X1 U9061 ( .C1(n10613), .C2(n8092), .A(n7844), .B(n7843), .ZN(n7845)
         );
  OAI21_X1 U9062 ( .B1(n7846), .B2(n10586), .A(n7845), .ZN(P2_U3261) );
  XNOR2_X1 U9063 ( .A(n7847), .B(n6764), .ZN(n7849) );
  AND2_X1 U9064 ( .A1(n8696), .A2(n8531), .ZN(n7848) );
  NOR2_X1 U9065 ( .A1(n7849), .A2(n7848), .ZN(n7895) );
  AOI21_X1 U9066 ( .B1(n7849), .B2(n7848), .A(n7895), .ZN(n7854) );
  INV_X1 U9067 ( .A(n7850), .ZN(n7851) );
  NAND2_X1 U9068 ( .A1(n7853), .A2(n7854), .ZN(n7897) );
  OAI21_X1 U9069 ( .B1(n7854), .B2(n7853), .A(n7897), .ZN(n7855) );
  NAND2_X1 U9070 ( .A1(n7855), .A2(n8683), .ZN(n7862) );
  NAND2_X1 U9071 ( .A1(n8685), .A2(n9013), .ZN(n7857) );
  OAI211_X1 U9072 ( .C1(n7858), .C2(n8688), .A(n7857), .B(n7856), .ZN(n7859)
         );
  AOI21_X1 U9073 ( .B1(n7860), .B2(n8690), .A(n7859), .ZN(n7861) );
  OAI211_X1 U9074 ( .C1(n10843), .C2(n8693), .A(n7862), .B(n7861), .ZN(
        P2_U3236) );
  NAND2_X1 U9075 ( .A1(n7863), .A2(n8211), .ZN(n7866) );
  AOI22_X1 U9076 ( .A1(n8135), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8134), .B2(
        n7864), .ZN(n7865) );
  NAND2_X1 U9077 ( .A1(n7866), .A2(n7865), .ZN(n7892) );
  OR2_X1 U9078 ( .A1(n7892), .A2(n8761), .ZN(n8286) );
  NAND2_X1 U9079 ( .A1(n7892), .A2(n8761), .ZN(n8090) );
  AOI21_X1 U9080 ( .B1(n8084), .B2(n7868), .A(n8760), .ZN(n10859) );
  INV_X1 U9081 ( .A(n7869), .ZN(n8270) );
  NAND2_X1 U9082 ( .A1(n7870), .A2(n8270), .ZN(n7871) );
  OAI211_X1 U9083 ( .C1(n5132), .C2(n8084), .A(n9017), .B(n8287), .ZN(n7881)
         );
  NAND2_X1 U9084 ( .A1(n8192), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n7879) );
  INV_X1 U9085 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10121) );
  OAI21_X1 U9086 ( .B1(n7873), .B2(n7872), .A(n10121), .ZN(n7874) );
  AND2_X1 U9087 ( .A1(n7874), .A2(n8095), .ZN(n9006) );
  NAND2_X1 U9088 ( .A1(n6516), .A2(n9006), .ZN(n7878) );
  INV_X1 U9089 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n7875) );
  OR2_X1 U9090 ( .A1(n8169), .A2(n7875), .ZN(n7877) );
  OR2_X1 U9091 ( .A1(n8171), .A2(n7553), .ZN(n7876) );
  NAND4_X1 U9092 ( .A1(n7879), .A2(n7878), .A3(n7877), .A4(n7876), .ZN(n8762)
         );
  AOI22_X1 U9093 ( .A1(n9012), .A2(n8696), .B1(n8762), .B2(n9014), .ZN(n7880)
         );
  NAND2_X1 U9094 ( .A1(n7881), .A2(n7880), .ZN(n10865) );
  XNOR2_X1 U9095 ( .A(n8744), .B(n10861), .ZN(n10863) );
  AOI22_X1 U9096 ( .A1(n10813), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7905), .B2(
        n10801), .ZN(n7883) );
  NAND2_X1 U9097 ( .A1(n7892), .A2(n9035), .ZN(n7882) );
  OAI211_X1 U9098 ( .C1(n10863), .C2(n8793), .A(n7883), .B(n7882), .ZN(n7884)
         );
  AOI21_X1 U9099 ( .B1(n10865), .B2(n10811), .A(n7884), .ZN(n7885) );
  OAI21_X1 U9100 ( .B1(n10859), .B2(n9022), .A(n7885), .ZN(P2_U3282) );
  INV_X1 U9101 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7889) );
  MUX2_X1 U9102 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(P2_DATAO_REG_25__SCAN_IN), 
        .S(n7958), .Z(n7924) );
  XNOR2_X1 U9103 ( .A(n7924), .B(SI_25_), .ZN(n7922) );
  XNOR2_X1 U9104 ( .A(n7923), .B(n7922), .ZN(n8417) );
  INV_X1 U9105 ( .A(n8417), .ZN(n7890) );
  OAI222_X1 U9106 ( .A1(n10455), .A2(n7889), .B1(n10451), .B2(n7890), .C1(
        n7888), .C2(P1_U3084), .ZN(P1_U3328) );
  INV_X1 U9107 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8186) );
  OAI222_X1 U9108 ( .A1(n7891), .A2(P2_U3152), .B1(n9153), .B2(n7890), .C1(
        n8186), .C2(n9151), .ZN(P2_U3333) );
  XNOR2_X1 U9109 ( .A(n7892), .B(n6764), .ZN(n7894) );
  AND2_X1 U9110 ( .A1(n9013), .A2(n8531), .ZN(n7893) );
  NOR2_X1 U9111 ( .A1(n7894), .A2(n7893), .ZN(n8475) );
  AOI21_X1 U9112 ( .B1(n7894), .B2(n7893), .A(n8475), .ZN(n7899) );
  INV_X1 U9113 ( .A(n7895), .ZN(n7896) );
  NAND2_X1 U9114 ( .A1(n7897), .A2(n7896), .ZN(n7898) );
  OAI21_X1 U9115 ( .B1(n7899), .B2(n7898), .A(n8477), .ZN(n7900) );
  NAND2_X1 U9116 ( .A1(n7900), .A2(n8683), .ZN(n7907) );
  AOI21_X1 U9117 ( .B1(n8685), .B2(n8762), .A(n7901), .ZN(n7902) );
  OAI21_X1 U9118 ( .B1(n7903), .B2(n8688), .A(n7902), .ZN(n7904) );
  AOI21_X1 U9119 ( .B1(n7905), .B2(n8690), .A(n7904), .ZN(n7906) );
  OAI211_X1 U9120 ( .C1(n10861), .C2(n8693), .A(n7907), .B(n7906), .ZN(
        P2_U3217) );
  NAND2_X1 U9121 ( .A1(n8720), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7909) );
  OAI21_X1 U9122 ( .B1(n8720), .B2(P2_REG2_REG_17__SCAN_IN), .A(n7909), .ZN(
        n7910) );
  NOR2_X1 U9123 ( .A1(n7911), .A2(n7910), .ZN(n8719) );
  AOI211_X1 U9124 ( .C1(n7911), .C2(n7910), .A(n8719), .B(n10607), .ZN(n7921)
         );
  INV_X1 U9125 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8108) );
  NOR2_X1 U9126 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8108), .ZN(n7912) );
  AOI21_X1 U9127 ( .B1(n10606), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n7912), .ZN(
        n7919) );
  XNOR2_X1 U9128 ( .A(n8711), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n7917) );
  INV_X1 U9129 ( .A(n8092), .ZN(n7915) );
  INV_X1 U9130 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n7914) );
  AOI21_X1 U9131 ( .B1(n7915), .B2(n7914), .A(n7913), .ZN(n7916) );
  NAND2_X1 U9132 ( .A1(n7917), .A2(n7916), .ZN(n8710) );
  OAI211_X1 U9133 ( .C1(n7917), .C2(n7916), .A(n10615), .B(n8710), .ZN(n7918)
         );
  OAI211_X1 U9134 ( .C1(n10585), .C2(n8711), .A(n7919), .B(n7918), .ZN(n7920)
         );
  OR2_X1 U9135 ( .A1(n7921), .A2(n7920), .ZN(P2_U3262) );
  INV_X1 U9136 ( .A(n7924), .ZN(n7926) );
  INV_X1 U9137 ( .A(SI_25_), .ZN(n7925) );
  NAND2_X1 U9138 ( .A1(n7926), .A2(n7925), .ZN(n7927) );
  MUX2_X1 U9139 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .S(n7958), .Z(n7932) );
  XNOR2_X1 U9140 ( .A(n7932), .B(n10027), .ZN(n7930) );
  XNOR2_X1 U9141 ( .A(n7931), .B(n7930), .ZN(n8426) );
  INV_X1 U9142 ( .A(n8426), .ZN(n7942) );
  INV_X1 U9143 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8199) );
  OAI222_X1 U9144 ( .A1(P2_U3152), .A2(n7929), .B1(n9153), .B2(n7942), .C1(
        n8199), .C2(n9151), .ZN(P2_U3332) );
  INV_X1 U9145 ( .A(n7932), .ZN(n7933) );
  NAND2_X1 U9146 ( .A1(n7933), .A2(n10027), .ZN(n7934) );
  MUX2_X1 U9147 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n5713), .Z(n7935) );
  NAND2_X1 U9148 ( .A1(n7935), .A2(SI_27_), .ZN(n7947) );
  INV_X1 U9149 ( .A(n7935), .ZN(n7937) );
  INV_X1 U9150 ( .A(SI_27_), .ZN(n7936) );
  NAND2_X1 U9151 ( .A1(n7937), .A2(n7936), .ZN(n7938) );
  INV_X1 U9152 ( .A(n8437), .ZN(n7943) );
  AOI21_X1 U9153 ( .B1(n10445), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n7939), .ZN(
        n7940) );
  OAI21_X1 U9154 ( .B1(n7943), .B2(n10451), .A(n7940), .ZN(P1_U3326) );
  INV_X1 U9155 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7941) );
  OAI222_X1 U9156 ( .A1(n10451), .A2(n7942), .B1(P1_U3084), .B2(n5750), .C1(
        n7941), .C2(n10455), .ZN(P1_U3327) );
  OAI222_X1 U9157 ( .A1(n6280), .A2(P2_U3152), .B1(n9151), .B2(n7944), .C1(
        n7943), .C2(n9153), .ZN(P2_U3331) );
  NAND2_X1 U9158 ( .A1(n7948), .A2(n7947), .ZN(n7952) );
  INV_X1 U9159 ( .A(n7952), .ZN(n7950) );
  MUX2_X1 U9160 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n7958), .Z(n7954) );
  XNOR2_X1 U9161 ( .A(n7954), .B(SI_28_), .ZN(n7951) );
  INV_X1 U9162 ( .A(n7951), .ZN(n7949) );
  NAND2_X1 U9163 ( .A1(n7952), .A2(n7951), .ZN(n7953) );
  NAND2_X1 U9164 ( .A1(n7957), .A2(n7953), .ZN(n8441) );
  INV_X1 U9165 ( .A(n8441), .ZN(n10453) );
  INV_X1 U9166 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7984) );
  OAI222_X1 U9167 ( .A1(n6278), .A2(P2_U3152), .B1(n9153), .B2(n10453), .C1(
        n7984), .C2(n9151), .ZN(P2_U3330) );
  INV_X1 U9168 ( .A(n7954), .ZN(n7955) );
  INV_X1 U9169 ( .A(SI_28_), .ZN(n10225) );
  NAND2_X1 U9170 ( .A1(n7955), .A2(n10225), .ZN(n7956) );
  INV_X1 U9171 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9152) );
  INV_X1 U9172 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10448) );
  MUX2_X1 U9173 ( .A(n9152), .B(n10448), .S(n7958), .Z(n7959) );
  INV_X1 U9174 ( .A(SI_29_), .ZN(n10229) );
  MUX2_X1 U9175 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n7966), .Z(n7963) );
  XNOR2_X1 U9176 ( .A(n7963), .B(SI_30_), .ZN(n7976) );
  INV_X1 U9177 ( .A(n7976), .ZN(n7962) );
  NAND2_X1 U9178 ( .A1(n7977), .A2(n7962), .ZN(n7965) );
  NAND2_X1 U9179 ( .A1(n7963), .A2(SI_30_), .ZN(n7964) );
  MUX2_X1 U9180 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7966), .Z(n7967) );
  XNOR2_X1 U9181 ( .A(n7967), .B(SI_31_), .ZN(n7968) );
  NAND2_X1 U9182 ( .A1(n9419), .A2(n8211), .ZN(n7972) );
  INV_X1 U9183 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n7970) );
  OR2_X1 U9184 ( .A1(n5137), .A2(n7970), .ZN(n7971) );
  INV_X1 U9185 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8750) );
  NAND2_X1 U9186 ( .A1(n8192), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n7975) );
  INV_X1 U9187 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n7973) );
  OR2_X1 U9188 ( .A1(n8169), .A2(n7973), .ZN(n7974) );
  OAI211_X1 U9189 ( .C1(n8171), .C2(n8750), .A(n7975), .B(n7974), .ZN(n8694)
         );
  INV_X1 U9190 ( .A(n8694), .ZN(n8749) );
  OR2_X1 U9191 ( .A1(n8746), .A2(n8749), .ZN(n8241) );
  NAND2_X1 U9192 ( .A1(n9412), .A2(n8211), .ZN(n7979) );
  INV_X1 U9193 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8548) );
  OR2_X1 U9194 ( .A1(n5137), .A2(n8548), .ZN(n7978) );
  NAND2_X1 U9195 ( .A1(n8757), .A2(n8789), .ZN(n8239) );
  OR2_X1 U9196 ( .A1(n8757), .A2(n8789), .ZN(n8316) );
  INV_X1 U9197 ( .A(n8316), .ZN(n7980) );
  NOR2_X1 U9198 ( .A1(n8318), .A2(n7980), .ZN(n8281) );
  NAND2_X1 U9199 ( .A1(n9428), .A2(n8211), .ZN(n7983) );
  OR2_X1 U9200 ( .A1(n5137), .A2(n9152), .ZN(n7982) );
  OR2_X1 U9201 ( .A1(n8791), .A2(n8809), .ZN(n8313) );
  NAND2_X1 U9202 ( .A1(n8791), .A2(n8809), .ZN(n8312) );
  OR2_X1 U9203 ( .A1(n5137), .A2(n7984), .ZN(n7985) );
  NAND2_X1 U9204 ( .A1(n8216), .A2(n10292), .ZN(n7986) );
  INV_X1 U9205 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n7990) );
  NAND2_X1 U9206 ( .A1(n8218), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n7989) );
  NAND2_X1 U9207 ( .A1(n8219), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7988) );
  OAI211_X1 U9208 ( .C1(n8223), .C2(n7990), .A(n7989), .B(n7988), .ZN(n7991)
         );
  MUX2_X1 U9209 ( .A(n8232), .B(n8311), .S(n5255), .Z(n8237) );
  OR2_X1 U9210 ( .A1(n8404), .A2(n6702), .ZN(n7994) );
  OR2_X1 U9211 ( .A1(n5137), .A2(n7992), .ZN(n7993) );
  INV_X1 U9212 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10314) );
  NAND2_X1 U9213 ( .A1(n8005), .A2(n10314), .ZN(n7995) );
  NAND2_X1 U9214 ( .A1(n8189), .A2(n7995), .ZN(n8632) );
  OR2_X1 U9215 ( .A1(n8632), .A2(n8217), .ZN(n7998) );
  AOI22_X1 U9216 ( .A1(n8192), .A2(P2_REG1_REG_24__SCAN_IN), .B1(n8219), .B2(
        P2_REG0_REG_24__SCAN_IN), .ZN(n7997) );
  NAND2_X1 U9217 ( .A1(n8218), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n7996) );
  NAND2_X1 U9218 ( .A1(n8390), .A2(n8211), .ZN(n8001) );
  OR2_X1 U9219 ( .A1(n5137), .A2(n7999), .ZN(n8000) );
  NAND2_X1 U9220 ( .A1(n8219), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8003) );
  NAND2_X1 U9221 ( .A1(n8218), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8002) );
  AND2_X1 U9222 ( .A1(n8003), .A2(n8002), .ZN(n8008) );
  NAND2_X1 U9223 ( .A1(n8015), .A2(n10291), .ZN(n8004) );
  AND2_X1 U9224 ( .A1(n8005), .A2(n8004), .ZN(n8883) );
  NAND2_X1 U9225 ( .A1(n8883), .A2(n8191), .ZN(n8007) );
  NAND2_X1 U9226 ( .A1(n8192), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8006) );
  OR2_X1 U9227 ( .A1(n9081), .A2(n8773), .ZN(n8277) );
  NAND2_X1 U9228 ( .A1(n8307), .A2(n8277), .ZN(n8010) );
  NAND2_X1 U9229 ( .A1(n9076), .A2(n8601), .ZN(n8254) );
  NAND2_X1 U9230 ( .A1(n9081), .A2(n8773), .ZN(n8868) );
  NAND2_X1 U9231 ( .A1(n8254), .A2(n8868), .ZN(n8009) );
  MUX2_X1 U9232 ( .A(n8010), .B(n8009), .S(n8242), .Z(n8011) );
  INV_X1 U9233 ( .A(n8011), .ZN(n8185) );
  NAND2_X1 U9234 ( .A1(n8385), .A2(n8211), .ZN(n8013) );
  OR2_X1 U9235 ( .A1(n5137), .A2(n7473), .ZN(n8012) );
  NAND2_X1 U9236 ( .A1(n8192), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8022) );
  INV_X1 U9237 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8014) );
  INV_X1 U9238 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10106) );
  OAI21_X1 U9239 ( .B1(n8167), .B2(n8014), .A(n10106), .ZN(n8016) );
  NAND2_X1 U9240 ( .A1(n8016), .A2(n8015), .ZN(n8898) );
  OR2_X1 U9241 ( .A1(n8217), .A2(n8898), .ZN(n8021) );
  INV_X1 U9242 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8017) );
  OR2_X1 U9243 ( .A1(n8169), .A2(n8017), .ZN(n8020) );
  INV_X1 U9244 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8018) );
  OR2_X1 U9245 ( .A1(n8171), .A2(n8018), .ZN(n8019) );
  XNOR2_X1 U9246 ( .A(n9086), .B(n8772), .ZN(n8902) );
  NAND2_X1 U9247 ( .A1(n8024), .A2(n8023), .ZN(n8256) );
  AND2_X1 U9248 ( .A1(n8025), .A2(n8256), .ZN(n8026) );
  MUX2_X1 U9249 ( .A(n8028), .B(n8027), .S(n8242), .Z(n8029) );
  INV_X1 U9250 ( .A(n8030), .ZN(n8032) );
  MUX2_X1 U9251 ( .A(n8033), .B(n8706), .S(n8242), .Z(n8031) );
  NAND2_X1 U9252 ( .A1(n8706), .A2(n8033), .ZN(n8034) );
  NOR2_X1 U9253 ( .A1(n8035), .A2(n8034), .ZN(n8036) );
  OR2_X1 U9254 ( .A1(n8037), .A2(n8036), .ZN(n8041) );
  INV_X1 U9255 ( .A(n8259), .ZN(n8040) );
  NOR2_X1 U9256 ( .A1(n8038), .A2(n5255), .ZN(n8039) );
  AOI21_X1 U9257 ( .B1(n8041), .B2(n8040), .A(n8039), .ZN(n8048) );
  NAND2_X1 U9258 ( .A1(n8043), .A2(n8042), .ZN(n8044) );
  MUX2_X1 U9259 ( .A(n8045), .B(n8044), .S(n8242), .Z(n8046) );
  MUX2_X1 U9260 ( .A(n8703), .B(n8049), .S(n8242), .Z(n8053) );
  INV_X1 U9261 ( .A(n8053), .ZN(n8051) );
  NAND2_X1 U9262 ( .A1(n8051), .A2(n8050), .ZN(n8054) );
  MUX2_X1 U9263 ( .A(n8056), .B(n8055), .S(n8242), .Z(n8057) );
  MUX2_X1 U9264 ( .A(n8059), .B(n8058), .S(n8242), .Z(n8060) );
  NAND2_X1 U9265 ( .A1(n8061), .A2(n8060), .ZN(n8065) );
  AND2_X1 U9266 ( .A1(n8067), .A2(n8068), .ZN(n8062) );
  MUX2_X1 U9267 ( .A(n8064), .B(n8062), .S(n8242), .Z(n8063) );
  NAND2_X1 U9268 ( .A1(n8063), .A2(n8070), .ZN(n8069) );
  AOI21_X1 U9269 ( .B1(n8065), .B2(n8064), .A(n8069), .ZN(n8075) );
  OAI211_X1 U9270 ( .C1(n8069), .C2(n8068), .A(n8067), .B(n8066), .ZN(n8073)
         );
  NAND2_X1 U9271 ( .A1(n8071), .A2(n8070), .ZN(n8072) );
  MUX2_X1 U9272 ( .A(n8073), .B(n8072), .S(n8242), .Z(n8074) );
  NAND2_X1 U9273 ( .A1(n8077), .A2(n8076), .ZN(n8078) );
  MUX2_X1 U9274 ( .A(n8079), .B(n8078), .S(n5255), .Z(n8080) );
  MUX2_X1 U9275 ( .A(n8082), .B(n8081), .S(n8242), .Z(n8083) );
  OR2_X1 U9276 ( .A1(n8085), .A2(n6702), .ZN(n8088) );
  AOI22_X1 U9277 ( .A1(n8135), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8134), .B2(
        n8086), .ZN(n8087) );
  INV_X1 U9278 ( .A(n8762), .ZN(n8089) );
  OR2_X1 U9279 ( .A1(n9123), .A2(n8089), .ZN(n8289) );
  NAND2_X1 U9280 ( .A1(n9123), .A2(n8089), .ZN(n8288) );
  MUX2_X1 U9281 ( .A(n8090), .B(n8286), .S(n5255), .Z(n8091) );
  NAND2_X1 U9282 ( .A1(n8329), .A2(n8211), .ZN(n8094) );
  AOI22_X1 U9283 ( .A1(n8135), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8134), .B2(
        n8092), .ZN(n8093) );
  NAND2_X1 U9284 ( .A1(n8192), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8102) );
  NAND2_X1 U9285 ( .A1(n8095), .A2(n10308), .ZN(n8096) );
  AND2_X1 U9286 ( .A1(n8109), .A2(n8096), .ZN(n8997) );
  NAND2_X1 U9287 ( .A1(n6516), .A2(n8997), .ZN(n8101) );
  INV_X1 U9288 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8097) );
  OR2_X1 U9289 ( .A1(n8169), .A2(n8097), .ZN(n8100) );
  INV_X1 U9290 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8098) );
  OR2_X1 U9291 ( .A1(n8171), .A2(n8098), .ZN(n8099) );
  NAND4_X1 U9292 ( .A1(n8102), .A2(n8101), .A3(n8100), .A4(n8099), .ZN(n9015)
         );
  INV_X1 U9293 ( .A(n9015), .ZN(n8103) );
  OR2_X1 U9294 ( .A1(n9119), .A2(n8103), .ZN(n8292) );
  NAND2_X1 U9295 ( .A1(n9119), .A2(n8103), .ZN(n8291) );
  MUX2_X1 U9296 ( .A(n8288), .B(n8289), .S(n8242), .Z(n8104) );
  NAND3_X1 U9297 ( .A1(n8105), .A2(n8993), .A3(n8104), .ZN(n8117) );
  OR2_X1 U9298 ( .A1(n8334), .A2(n6702), .ZN(n8107) );
  AOI22_X1 U9299 ( .A1(n8135), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8134), .B2(
        n8720), .ZN(n8106) );
  NAND2_X1 U9300 ( .A1(n8192), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8115) );
  NAND2_X1 U9301 ( .A1(n8109), .A2(n8108), .ZN(n8110) );
  AND2_X1 U9302 ( .A1(n8120), .A2(n8110), .ZN(n8622) );
  NAND2_X1 U9303 ( .A1(n8191), .A2(n8622), .ZN(n8114) );
  INV_X1 U9304 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8111) );
  OR2_X1 U9305 ( .A1(n8169), .A2(n8111), .ZN(n8113) );
  INV_X1 U9306 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8983) );
  OR2_X1 U9307 ( .A1(n8171), .A2(n8983), .ZN(n8112) );
  NAND4_X1 U9308 ( .A1(n8115), .A2(n8114), .A3(n8113), .A4(n8112), .ZN(n8965)
         );
  NAND2_X1 U9309 ( .A1(n9114), .A2(n8764), .ZN(n8128) );
  NAND2_X1 U9310 ( .A1(n8295), .A2(n8128), .ZN(n8973) );
  INV_X1 U9311 ( .A(n8973), .ZN(n8294) );
  MUX2_X1 U9312 ( .A(n8291), .B(n8292), .S(n5255), .Z(n8116) );
  NAND3_X1 U9313 ( .A1(n8117), .A2(n8294), .A3(n8116), .ZN(n8130) );
  NAND2_X1 U9314 ( .A1(n8347), .A2(n8211), .ZN(n8119) );
  AOI22_X1 U9315 ( .A1(n8135), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8134), .B2(
        n8729), .ZN(n8118) );
  NAND2_X1 U9316 ( .A1(n8192), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8127) );
  NAND2_X1 U9317 ( .A1(n8120), .A2(n10117), .ZN(n8121) );
  AND2_X1 U9318 ( .A1(n8138), .A2(n8121), .ZN(n8958) );
  NAND2_X1 U9319 ( .A1(n8191), .A2(n8958), .ZN(n8126) );
  INV_X1 U9320 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8122) );
  OR2_X1 U9321 ( .A1(n8169), .A2(n8122), .ZN(n8125) );
  INV_X1 U9322 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8123) );
  OR2_X1 U9323 ( .A1(n8171), .A2(n8123), .ZN(n8124) );
  NAND4_X1 U9324 ( .A1(n8127), .A2(n8126), .A3(n8125), .A4(n8124), .ZN(n8695)
         );
  INV_X1 U9325 ( .A(n8695), .ZN(n8767) );
  NAND2_X1 U9326 ( .A1(n9108), .A2(n8767), .ZN(n8131) );
  NAND2_X1 U9327 ( .A1(n8297), .A2(n8131), .ZN(n8768) );
  MUX2_X1 U9328 ( .A(n8128), .B(n8295), .S(n8242), .Z(n8129) );
  NAND3_X1 U9329 ( .A1(n8130), .A2(n8962), .A3(n8129), .ZN(n8133) );
  MUX2_X1 U9330 ( .A(n8131), .B(n8297), .S(n5255), .Z(n8132) );
  NAND2_X1 U9331 ( .A1(n8133), .A2(n8132), .ZN(n8145) );
  NAND2_X1 U9332 ( .A1(n8351), .A2(n8211), .ZN(n8137) );
  AOI22_X1 U9333 ( .A1(n8135), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5256), .B2(
        n8134), .ZN(n8136) );
  NAND2_X1 U9334 ( .A1(n8192), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n8144) );
  INV_X1 U9335 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10081) );
  NAND2_X1 U9336 ( .A1(n8138), .A2(n10081), .ZN(n8139) );
  AND2_X1 U9337 ( .A1(n8151), .A2(n8139), .ZN(n8583) );
  NAND2_X1 U9338 ( .A1(n6516), .A2(n8583), .ZN(n8143) );
  INV_X1 U9339 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8140) );
  OR2_X1 U9340 ( .A1(n8169), .A2(n8140), .ZN(n8142) );
  INV_X1 U9341 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8730) );
  OR2_X1 U9342 ( .A1(n8171), .A2(n8730), .ZN(n8141) );
  NAND4_X1 U9343 ( .A1(n8144), .A2(n8143), .A3(n8142), .A4(n8141), .ZN(n8964)
         );
  NAND2_X1 U9344 ( .A1(n9103), .A2(n8769), .ZN(n8146) );
  NAND2_X1 U9345 ( .A1(n8299), .A2(n8146), .ZN(n8943) );
  INV_X1 U9346 ( .A(n8943), .ZN(n8298) );
  NAND2_X1 U9347 ( .A1(n8145), .A2(n8298), .ZN(n8148) );
  MUX2_X1 U9348 ( .A(n8146), .B(n8299), .S(n5255), .Z(n8147) );
  NAND2_X1 U9349 ( .A1(n8362), .A2(n8211), .ZN(n8150) );
  INV_X1 U9350 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8545) );
  OR2_X1 U9351 ( .A1(n5137), .A2(n8545), .ZN(n8149) );
  NAND2_X1 U9352 ( .A1(n8151), .A2(n10320), .ZN(n8152) );
  AND2_X1 U9353 ( .A1(n8167), .A2(n8152), .ZN(n8929) );
  NAND2_X1 U9354 ( .A1(n8191), .A2(n8929), .ZN(n8158) );
  NAND2_X1 U9355 ( .A1(n8192), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8157) );
  INV_X1 U9356 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8153) );
  OR2_X1 U9357 ( .A1(n8169), .A2(n8153), .ZN(n8156) );
  INV_X1 U9358 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8154) );
  OR2_X1 U9359 ( .A1(n8171), .A2(n8154), .ZN(n8155) );
  NAND4_X1 U9360 ( .A1(n8158), .A2(n8157), .A3(n8156), .A4(n8155), .ZN(n8920)
         );
  NAND2_X1 U9361 ( .A1(n9096), .A2(n8920), .ZN(n8770) );
  INV_X1 U9362 ( .A(n8770), .ZN(n8159) );
  NAND2_X1 U9363 ( .A1(n8162), .A2(n8159), .ZN(n8161) );
  MUX2_X1 U9364 ( .A(n8920), .B(n9096), .S(n5255), .Z(n8160) );
  NAND2_X1 U9365 ( .A1(n8161), .A2(n8160), .ZN(n8163) );
  OR2_X1 U9366 ( .A1(n8372), .A2(n6702), .ZN(n8166) );
  OR2_X1 U9367 ( .A1(n5137), .A2(n8164), .ZN(n8165) );
  XNOR2_X1 U9368 ( .A(n8167), .B(P2_REG3_REG_21__SCAN_IN), .ZN(n8913) );
  NAND2_X1 U9369 ( .A1(n6516), .A2(n8913), .ZN(n8175) );
  NAND2_X1 U9370 ( .A1(n8192), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8174) );
  INV_X1 U9371 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8168) );
  OR2_X1 U9372 ( .A1(n8169), .A2(n8168), .ZN(n8173) );
  INV_X1 U9373 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8170) );
  OR2_X1 U9374 ( .A1(n8171), .A2(n8170), .ZN(n8172) );
  NAND4_X1 U9375 ( .A1(n8175), .A2(n8174), .A3(n8173), .A4(n8172), .ZN(n8935)
         );
  NAND2_X1 U9376 ( .A1(n9091), .A2(n8935), .ZN(n8176) );
  INV_X1 U9377 ( .A(n8916), .ZN(n8178) );
  NOR2_X1 U9378 ( .A1(n8935), .A2(n8242), .ZN(n8177) );
  AND2_X1 U9379 ( .A1(n9086), .A2(n8772), .ZN(n8180) );
  INV_X1 U9380 ( .A(n8935), .ZN(n8648) );
  OR2_X1 U9381 ( .A1(n9091), .A2(n8648), .ZN(n8302) );
  OR2_X1 U9382 ( .A1(n9086), .A2(n8772), .ZN(n8303) );
  OAI211_X1 U9383 ( .C1(n8902), .C2(n8302), .A(n8277), .B(n8303), .ZN(n8179)
         );
  MUX2_X1 U9384 ( .A(n8180), .B(n8179), .S(n8242), .Z(n8181) );
  INV_X1 U9385 ( .A(n8181), .ZN(n8182) );
  OAI211_X1 U9386 ( .C1(n8902), .C2(n8183), .A(n8182), .B(n8868), .ZN(n8184)
         );
  NAND2_X1 U9387 ( .A1(n8417), .A2(n8211), .ZN(n8188) );
  OR2_X1 U9388 ( .A1(n5137), .A2(n8186), .ZN(n8187) );
  NAND2_X1 U9389 ( .A1(n8189), .A2(n10309), .ZN(n8190) );
  AND2_X1 U9390 ( .A1(n8202), .A2(n8190), .ZN(n8852) );
  NAND2_X1 U9391 ( .A1(n8852), .A2(n8191), .ZN(n8195) );
  AOI22_X1 U9392 ( .A1(n8218), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8219), .B2(
        P2_REG0_REG_25__SCAN_IN), .ZN(n8194) );
  NAND2_X1 U9393 ( .A1(n8192), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8193) );
  NAND2_X1 U9394 ( .A1(n9071), .A2(n8672), .ZN(n8276) );
  INV_X1 U9395 ( .A(n8601), .ZN(n8775) );
  OAI211_X1 U9396 ( .C1(n8775), .C2(n8242), .A(n8196), .B(n8307), .ZN(n8197)
         );
  NAND3_X1 U9397 ( .A1(n8198), .A2(n8276), .A3(n8197), .ZN(n8231) );
  NAND2_X1 U9398 ( .A1(n8426), .A2(n8211), .ZN(n8201) );
  OR2_X1 U9399 ( .A1(n5137), .A2(n8199), .ZN(n8200) );
  INV_X1 U9400 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8673) );
  NAND2_X1 U9401 ( .A1(n8202), .A2(n8673), .ZN(n8203) );
  NAND2_X1 U9402 ( .A1(n8214), .A2(n8203), .ZN(n8840) );
  INV_X1 U9403 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8206) );
  NAND2_X1 U9404 ( .A1(n8219), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8205) );
  NAND2_X1 U9405 ( .A1(n8218), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8204) );
  OAI211_X1 U9406 ( .C1(n8223), .C2(n8206), .A(n8205), .B(n8204), .ZN(n8207)
         );
  INV_X1 U9407 ( .A(n8207), .ZN(n8208) );
  NAND2_X1 U9408 ( .A1(n9065), .A2(n8602), .ZN(n8309) );
  NAND3_X1 U9409 ( .A1(n8231), .A2(n8276), .A3(n8309), .ZN(n8210) );
  NAND3_X1 U9410 ( .A1(n8210), .A2(n5255), .A3(n8253), .ZN(n8229) );
  NAND2_X1 U9411 ( .A1(n8437), .A2(n8211), .ZN(n8213) );
  OR2_X1 U9412 ( .A1(n5137), .A2(n7944), .ZN(n8212) );
  NAND2_X1 U9413 ( .A1(n8214), .A2(n8567), .ZN(n8215) );
  NAND2_X1 U9414 ( .A1(n8216), .A2(n8215), .ZN(n8820) );
  INV_X1 U9415 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8222) );
  NAND2_X1 U9416 ( .A1(n8218), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8221) );
  NAND2_X1 U9417 ( .A1(n8219), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8220) );
  OAI211_X1 U9418 ( .C1(n8223), .C2(n8222), .A(n8221), .B(n8220), .ZN(n8224)
         );
  INV_X1 U9419 ( .A(n8224), .ZN(n8225) );
  NAND2_X1 U9420 ( .A1(n8779), .A2(n5255), .ZN(n8227) );
  NOR2_X1 U9421 ( .A1(n9059), .A2(n8227), .ZN(n8228) );
  AOI21_X1 U9422 ( .B1(n8229), .B2(n8816), .A(n8228), .ZN(n8235) );
  AND2_X1 U9423 ( .A1(n8253), .A2(n8833), .ZN(n8310) );
  NAND2_X1 U9424 ( .A1(n8309), .A2(n8242), .ZN(n8230) );
  AOI21_X1 U9425 ( .B1(n8231), .B2(n8310), .A(n8230), .ZN(n8234) );
  NAND3_X1 U9426 ( .A1(n9059), .A2(n8807), .A3(n8242), .ZN(n8233) );
  OAI211_X1 U9427 ( .C1(n8235), .C2(n8234), .A(n8804), .B(n8233), .ZN(n8236)
         );
  NAND3_X1 U9428 ( .A1(n8785), .A2(n8237), .A3(n8236), .ZN(n8240) );
  MUX2_X1 U9429 ( .A(n8312), .B(n8313), .S(n5255), .Z(n8238) );
  INV_X1 U9430 ( .A(n8241), .ZN(n8243) );
  MUX2_X1 U9431 ( .A(n8318), .B(n8243), .S(n8242), .Z(n8244) );
  AOI21_X1 U9432 ( .B1(n10640), .B2(n8246), .A(n8249), .ZN(n8247) );
  INV_X1 U9433 ( .A(n8247), .ZN(n8323) );
  OAI21_X1 U9434 ( .B1(n8252), .B2(n8251), .A(n8250), .ZN(n8322) );
  INV_X1 U9435 ( .A(n8920), .ZN(n8594) );
  XNOR2_X1 U9436 ( .A(n9096), .B(n8594), .ZN(n8925) );
  INV_X1 U9437 ( .A(n8255), .ZN(n8271) );
  INV_X1 U9438 ( .A(n10788), .ZN(n10795) );
  INV_X1 U9439 ( .A(n8256), .ZN(n8258) );
  INV_X1 U9440 ( .A(n6732), .ZN(n8257) );
  NAND3_X1 U9441 ( .A1(n8258), .A2(n8248), .A3(n8257), .ZN(n8260) );
  NOR4_X1 U9442 ( .A1(n8262), .A2(n8261), .A3(n8260), .A4(n8259), .ZN(n8265)
         );
  NAND4_X1 U9443 ( .A1(n8265), .A2(n9031), .A3(n8264), .A4(n8263), .ZN(n8267)
         );
  NOR4_X1 U9444 ( .A1(n8268), .A2(n7415), .A3(n8267), .A4(n8266), .ZN(n8269)
         );
  NAND4_X1 U9445 ( .A1(n8271), .A2(n8270), .A3(n10795), .A4(n8269), .ZN(n8272)
         );
  NOR4_X1 U9446 ( .A1(n8973), .A2(n8273), .A3(n9010), .A4(n8272), .ZN(n8274)
         );
  NAND4_X1 U9447 ( .A1(n8298), .A2(n8962), .A3(n8993), .A4(n8274), .ZN(n8275)
         );
  NOR4_X1 U9448 ( .A1(n8870), .A2(n8916), .A3(n8925), .A4(n8275), .ZN(n8278)
         );
  NAND2_X1 U9449 ( .A1(n8833), .A2(n8276), .ZN(n8844) );
  INV_X1 U9450 ( .A(n8844), .ZN(n8849) );
  NAND2_X1 U9451 ( .A1(n8277), .A2(n8868), .ZN(n8878) );
  INV_X1 U9452 ( .A(n8902), .ZN(n8893) );
  NAND4_X1 U9453 ( .A1(n8278), .A2(n8849), .A3(n8304), .A4(n8893), .ZN(n8279)
         );
  NOR4_X1 U9454 ( .A1(n8781), .A2(n8824), .A3(n8834), .A4(n8279), .ZN(n8280)
         );
  NAND4_X1 U9455 ( .A1(n8281), .A2(n5077), .A3(n8785), .A4(n8280), .ZN(n8282)
         );
  XNOR2_X1 U9456 ( .A(n8282), .B(n6499), .ZN(n8283) );
  NOR2_X1 U9457 ( .A1(n6755), .A2(n6499), .ZN(n8320) );
  OAI21_X1 U9458 ( .B1(n5256), .B2(n6755), .A(n8531), .ZN(n8319) );
  NAND2_X1 U9459 ( .A1(n8992), .A2(n8291), .ZN(n8293) );
  NAND2_X1 U9460 ( .A1(n8293), .A2(n8292), .ZN(n8974) );
  NAND2_X1 U9461 ( .A1(n8974), .A2(n8294), .ZN(n8296) );
  NAND2_X1 U9462 ( .A1(n8296), .A2(n8295), .ZN(n8963) );
  NAND2_X1 U9463 ( .A1(n8963), .A2(n8962), .ZN(n8961) );
  INV_X1 U9464 ( .A(n8925), .ZN(n8933) );
  OR2_X1 U9465 ( .A1(n9096), .A2(n8594), .ZN(n8300) );
  NAND2_X1 U9466 ( .A1(n9091), .A2(n8648), .ZN(n8301) );
  INV_X1 U9467 ( .A(n8868), .ZN(n8305) );
  NOR2_X1 U9468 ( .A1(n8870), .A2(n8305), .ZN(n8306) );
  NAND2_X1 U9469 ( .A1(n8867), .A2(n8306), .ZN(n8308) );
  NAND2_X1 U9470 ( .A1(n8308), .A2(n8307), .ZN(n8850) );
  NOR4_X1 U9471 ( .A1(n6615), .A2(n10462), .A3(n6280), .A4(n8806), .ZN(n8326)
         );
  OAI21_X1 U9472 ( .B1(n8327), .B2(n8324), .A(P2_B_REG_SCAN_IN), .ZN(n8325) );
  OAI22_X1 U9473 ( .A1(n5086), .A2(n8327), .B1(n8326), .B2(n8325), .ZN(
        P2_U3244) );
  INV_X1 U9474 ( .A(n9887), .ZN(n9911) );
  NAND2_X1 U9475 ( .A1(n10876), .A2(n9911), .ZN(n8328) );
  NAND2_X1 U9476 ( .A1(n10874), .A2(n8328), .ZN(n9893) );
  NAND2_X1 U9477 ( .A1(n8329), .A2(n9427), .ZN(n8332) );
  AOI22_X1 U9478 ( .A1(n8442), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8352), .B2(
        n8330), .ZN(n8331) );
  NAND2_X1 U9479 ( .A1(n10886), .A2(n9336), .ZN(n9545) );
  NAND2_X1 U9480 ( .A1(n9544), .A2(n9545), .ZN(n9892) );
  INV_X1 U9481 ( .A(n9336), .ZN(n9879) );
  NAND2_X1 U9482 ( .A1(n10886), .A2(n9879), .ZN(n8333) );
  OR2_X1 U9483 ( .A1(n8334), .A2(n6231), .ZN(n8337) );
  AOI22_X1 U9484 ( .A1(n8442), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n8352), .B2(
        n8335), .ZN(n8336) );
  NAND2_X1 U9485 ( .A1(n6031), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8345) );
  NAND2_X1 U9486 ( .A1(n8339), .A2(n8338), .ZN(n8340) );
  AND2_X1 U9487 ( .A1(n8341), .A2(n8340), .ZN(n9872) );
  NAND2_X1 U9488 ( .A1(n6576), .A2(n9872), .ZN(n8344) );
  NAND2_X1 U9489 ( .A1(n6933), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8343) );
  NAND2_X1 U9490 ( .A1(n9423), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n8342) );
  NAND2_X1 U9491 ( .A1(n9998), .A2(n9890), .ZN(n9549) );
  INV_X1 U9492 ( .A(n9890), .ZN(n9852) );
  OR2_X1 U9493 ( .A1(n9998), .A2(n9852), .ZN(n8346) );
  NAND2_X1 U9494 ( .A1(n8347), .A2(n9427), .ZN(n8350) );
  AOI22_X1 U9495 ( .A1(n8348), .A2(n8352), .B1(n8442), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n8349) );
  INV_X1 U9496 ( .A(n9878), .ZN(n9837) );
  OR2_X1 U9497 ( .A1(n9993), .A2(n9837), .ZN(n9553) );
  NAND2_X1 U9498 ( .A1(n9993), .A2(n9837), .ZN(n9554) );
  NAND2_X1 U9499 ( .A1(n8351), .A2(n9427), .ZN(n8354) );
  AOI22_X1 U9500 ( .A1(n8442), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9760), .B2(
        n8352), .ZN(n8353) );
  OR2_X1 U9501 ( .A1(n8355), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8356) );
  NAND2_X1 U9502 ( .A1(n8365), .A2(n8356), .ZN(n9842) );
  AOI22_X1 U9503 ( .A1(n6933), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9423), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n8358) );
  NAND2_X1 U9504 ( .A1(n6031), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n8357) );
  OAI211_X1 U9505 ( .C1(n9842), .C2(n8400), .A(n8358), .B(n8357), .ZN(n9853)
         );
  OR2_X1 U9506 ( .A1(n9987), .A2(n9853), .ZN(n8359) );
  NAND2_X1 U9507 ( .A1(n9832), .A2(n8359), .ZN(n8361) );
  NAND2_X1 U9508 ( .A1(n9987), .A2(n9853), .ZN(n8360) );
  NAND2_X1 U9509 ( .A1(n8361), .A2(n8360), .ZN(n9822) );
  NAND2_X1 U9510 ( .A1(n8362), .A2(n9427), .ZN(n8364) );
  NAND2_X1 U9511 ( .A1(n8442), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8363) );
  NAND2_X1 U9512 ( .A1(n8365), .A2(n9356), .ZN(n8366) );
  NAND2_X1 U9513 ( .A1(n8375), .A2(n8366), .ZN(n9826) );
  OR2_X1 U9514 ( .A1(n9826), .A2(n8400), .ZN(n8369) );
  AOI22_X1 U9515 ( .A1(n6031), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n6933), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n8368) );
  NAND2_X1 U9516 ( .A1(n9423), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8367) );
  XNOR2_X1 U9517 ( .A(n9981), .B(n9838), .ZN(n9821) );
  NAND2_X1 U9518 ( .A1(n9822), .A2(n9821), .ZN(n8371) );
  INV_X1 U9519 ( .A(n9838), .ZN(n9667) );
  NAND2_X1 U9520 ( .A1(n9981), .A2(n9667), .ZN(n8370) );
  OR2_X1 U9521 ( .A1(n8372), .A2(n6231), .ZN(n8374) );
  NAND2_X1 U9522 ( .A1(n8442), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8373) );
  NAND2_X1 U9523 ( .A1(n8375), .A2(n9304), .ZN(n8376) );
  AND2_X1 U9524 ( .A1(n8377), .A2(n8376), .ZN(n9305) );
  NAND2_X1 U9525 ( .A1(n9305), .A2(n6576), .ZN(n8383) );
  INV_X1 U9526 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n8380) );
  NAND2_X1 U9527 ( .A1(n9423), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8379) );
  NAND2_X1 U9528 ( .A1(n6933), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8378) );
  OAI211_X1 U9529 ( .C1(n8412), .C2(n8380), .A(n8379), .B(n8378), .ZN(n8381)
         );
  INV_X1 U9530 ( .A(n8381), .ZN(n8382) );
  NAND2_X1 U9531 ( .A1(n9978), .A2(n9820), .ZN(n9565) );
  NAND2_X1 U9532 ( .A1(n8459), .A2(n9565), .ZN(n9806) );
  INV_X1 U9533 ( .A(n9820), .ZN(n9666) );
  NAND2_X1 U9534 ( .A1(n9978), .A2(n9666), .ZN(n8384) );
  NAND2_X1 U9535 ( .A1(n8385), .A2(n9427), .ZN(n8387) );
  NAND2_X1 U9536 ( .A1(n8442), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8386) );
  AND2_X1 U9537 ( .A1(n9971), .A2(n9775), .ZN(n8388) );
  OR2_X1 U9538 ( .A1(n9971), .A2(n9775), .ZN(n8389) );
  INV_X1 U9539 ( .A(n9765), .ZN(n8401) );
  NAND2_X1 U9540 ( .A1(n8390), .A2(n9427), .ZN(n8392) );
  NAND2_X1 U9541 ( .A1(n8442), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8391) );
  NOR2_X1 U9542 ( .A1(n8393), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8394) );
  OR2_X1 U9543 ( .A1(n8407), .A2(n8394), .ZN(n9768) );
  INV_X1 U9544 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n8397) );
  NAND2_X1 U9545 ( .A1(n6933), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8396) );
  NAND2_X1 U9546 ( .A1(n9423), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8395) );
  OAI211_X1 U9547 ( .C1(n8397), .C2(n8412), .A(n8396), .B(n8395), .ZN(n8398)
         );
  INV_X1 U9548 ( .A(n8398), .ZN(n8399) );
  NAND2_X1 U9549 ( .A1(n8401), .A2(n5619), .ZN(n8403) );
  NAND2_X1 U9550 ( .A1(n9966), .A2(n9799), .ZN(n8402) );
  OR2_X1 U9551 ( .A1(n8404), .A2(n6231), .ZN(n8406) );
  NAND2_X1 U9552 ( .A1(n8442), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8405) );
  OR2_X1 U9553 ( .A1(n8407), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8408) );
  AND2_X1 U9554 ( .A1(n8408), .A2(n8421), .ZN(n9758) );
  NAND2_X1 U9555 ( .A1(n9758), .A2(n6576), .ZN(n8415) );
  INV_X1 U9556 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n8411) );
  NAND2_X1 U9557 ( .A1(n6933), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8410) );
  NAND2_X1 U9558 ( .A1(n9423), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8409) );
  OAI211_X1 U9559 ( .C1(n8412), .C2(n8411), .A(n8410), .B(n8409), .ZN(n8413)
         );
  INV_X1 U9560 ( .A(n8413), .ZN(n8414) );
  NAND2_X1 U9561 ( .A1(n8415), .A2(n8414), .ZN(n9776) );
  AND2_X1 U9562 ( .A1(n9963), .A2(n9776), .ZN(n8416) );
  NAND2_X1 U9563 ( .A1(n8417), .A2(n9427), .ZN(n8419) );
  NAND2_X1 U9564 ( .A1(n8442), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8418) );
  INV_X1 U9565 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9314) );
  AOI21_X1 U9566 ( .B1(n9314), .B2(n8421), .A(n8420), .ZN(n9315) );
  NAND2_X1 U9567 ( .A1(n6931), .A2(n9315), .ZN(n8425) );
  NAND2_X1 U9568 ( .A1(n6031), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8424) );
  NAND2_X1 U9569 ( .A1(n6932), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8423) );
  NAND2_X1 U9570 ( .A1(n9423), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8422) );
  NAND2_X1 U9571 ( .A1(n9958), .A2(n9754), .ZN(n9499) );
  NAND2_X1 U9572 ( .A1(n9498), .A2(n9499), .ZN(n9738) );
  INV_X1 U9573 ( .A(n9754), .ZN(n9665) );
  NAND2_X1 U9574 ( .A1(n8426), .A2(n9427), .ZN(n8428) );
  NAND2_X1 U9575 ( .A1(n8442), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8427) );
  INV_X1 U9576 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9387) );
  AOI21_X1 U9577 ( .B1(n9387), .B2(n8429), .A(n8445), .ZN(n9730) );
  NAND2_X1 U9578 ( .A1(n6576), .A2(n9730), .ZN(n8433) );
  NAND2_X1 U9579 ( .A1(n6031), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8432) );
  NAND2_X1 U9580 ( .A1(n6933), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8431) );
  NAND2_X1 U9581 ( .A1(n9423), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8430) );
  NAND4_X1 U9582 ( .A1(n8433), .A2(n8432), .A3(n8431), .A4(n8430), .ZN(n9664)
         );
  NOR2_X1 U9583 ( .A1(n9951), .A2(n9664), .ZN(n8434) );
  OR2_X2 U9584 ( .A1(n9722), .A2(n8434), .ZN(n8436) );
  NAND2_X1 U9585 ( .A1(n9951), .A2(n9664), .ZN(n8435) );
  NAND2_X1 U9586 ( .A1(n8437), .A2(n9427), .ZN(n8439) );
  NAND2_X1 U9587 ( .A1(n8442), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8438) );
  NAND2_X1 U9588 ( .A1(n9948), .A2(n9723), .ZN(n9586) );
  NAND2_X1 U9589 ( .A1(n8441), .A2(n9427), .ZN(n8444) );
  NAND2_X1 U9590 ( .A1(n8442), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8443) );
  NAND2_X1 U9591 ( .A1(n6031), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8452) );
  INV_X1 U9592 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9293) );
  NAND2_X1 U9593 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n8445), .ZN(n8446) );
  NAND2_X1 U9594 ( .A1(n9293), .A2(n8446), .ZN(n8447) );
  NAND2_X1 U9595 ( .A1(n6576), .A2(n9294), .ZN(n8451) );
  NAND2_X1 U9596 ( .A1(n6933), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8450) );
  NAND2_X1 U9597 ( .A1(n9423), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8449) );
  NAND2_X1 U9598 ( .A1(n9941), .A2(n9712), .ZN(n9583) );
  NAND2_X1 U9599 ( .A1(n8453), .A2(n9686), .ZN(n8454) );
  NAND2_X1 U9600 ( .A1(n9702), .A2(n8454), .ZN(n9945) );
  INV_X1 U9601 ( .A(n9545), .ZN(n8456) );
  NAND2_X1 U9602 ( .A1(n9875), .A2(n9548), .ZN(n9856) );
  INV_X1 U9603 ( .A(n9548), .ZN(n8457) );
  NAND2_X1 U9604 ( .A1(n9554), .A2(n8457), .ZN(n8458) );
  AND2_X1 U9605 ( .A1(n8458), .A2(n9553), .ZN(n9434) );
  NAND2_X1 U9606 ( .A1(n9854), .A2(n9434), .ZN(n9834) );
  INV_X1 U9607 ( .A(n9853), .ZN(n9819) );
  OR2_X1 U9608 ( .A1(n9987), .A2(n9819), .ZN(n9559) );
  NAND2_X1 U9609 ( .A1(n9987), .A2(n9819), .ZN(n9560) );
  NAND2_X1 U9610 ( .A1(n9559), .A2(n9560), .ZN(n9835) );
  INV_X1 U9611 ( .A(n9560), .ZN(n9473) );
  OR2_X1 U9612 ( .A1(n9981), .A2(n9838), .ZN(n9804) );
  NAND2_X1 U9613 ( .A1(n8459), .A2(n9804), .ZN(n9566) );
  NAND3_X1 U9614 ( .A1(n8459), .A2(n9838), .A3(n9981), .ZN(n8460) );
  AND2_X1 U9615 ( .A1(n8460), .A2(n9565), .ZN(n9789) );
  INV_X1 U9616 ( .A(n9775), .ZN(n9808) );
  NAND2_X1 U9617 ( .A1(n9971), .A2(n9808), .ZN(n9570) );
  NAND2_X1 U9618 ( .A1(n9789), .A2(n9570), .ZN(n9792) );
  XNOR2_X1 U9619 ( .A(n9966), .B(n9799), .ZN(n9773) );
  NAND2_X1 U9620 ( .A1(n9774), .A2(n9773), .ZN(n9772) );
  OR2_X1 U9621 ( .A1(n9966), .A2(n9752), .ZN(n9432) );
  NAND2_X1 U9622 ( .A1(n9772), .A2(n9432), .ZN(n9751) );
  XNOR2_X1 U9623 ( .A(n9963), .B(n9776), .ZN(n9750) );
  INV_X1 U9624 ( .A(n9776), .ZN(n9741) );
  NOR2_X1 U9625 ( .A1(n9963), .A2(n9741), .ZN(n9574) );
  INV_X1 U9626 ( .A(n9664), .ZN(n9742) );
  OR2_X1 U9627 ( .A1(n9951), .A2(n9742), .ZN(n9496) );
  NAND2_X1 U9628 ( .A1(n9951), .A2(n9742), .ZN(n9497) );
  NAND2_X1 U9629 ( .A1(n9496), .A2(n9497), .ZN(n9726) );
  NAND2_X1 U9630 ( .A1(n9714), .A2(n9497), .ZN(n8461) );
  OAI21_X1 U9631 ( .B1(n9724), .B2(n8461), .A(n9495), .ZN(n9687) );
  INV_X1 U9632 ( .A(n9686), .ZN(n9645) );
  XNOR2_X1 U9633 ( .A(n9687), .B(n9645), .ZN(n8463) );
  OAI22_X1 U9634 ( .A1(n9723), .A2(n10755), .B1(n9484), .B2(n10753), .ZN(n8462) );
  INV_X1 U9635 ( .A(n9945), .ZN(n8472) );
  INV_X1 U9636 ( .A(n9941), .ZN(n9701) );
  INV_X1 U9637 ( .A(n9987), .ZN(n9846) );
  INV_X1 U9638 ( .A(n9993), .ZN(n9862) );
  NOR2_X1 U9639 ( .A1(n9971), .A2(n9810), .ZN(n9783) );
  INV_X1 U9640 ( .A(n9963), .ZN(n9350) );
  NOR2_X2 U9641 ( .A1(n9951), .A2(n9743), .ZN(n9729) );
  NAND2_X1 U9642 ( .A1(n9706), .A2(n9941), .ZN(n8468) );
  NAND2_X1 U9643 ( .A1(n9942), .A2(n10772), .ZN(n8470) );
  AOI22_X1 U9644 ( .A1(n10778), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9294), .B2(
        n10776), .ZN(n8469) );
  OAI211_X1 U9645 ( .C1(n9701), .C2(n10780), .A(n8470), .B(n8469), .ZN(n8471)
         );
  AOI21_X1 U9646 ( .B1(n8472), .B2(n10773), .A(n8471), .ZN(n8473) );
  OAI21_X1 U9647 ( .B1(n9944), .B2(n10778), .A(n8473), .ZN(P1_U3263) );
  INV_X1 U9648 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9413) );
  INV_X1 U9649 ( .A(n9412), .ZN(n8549) );
  OAI222_X1 U9650 ( .A1(n10455), .A2(n9413), .B1(n10451), .B2(n8549), .C1(
        P1_U3084), .C2(n8474), .ZN(P1_U3323) );
  INV_X1 U9651 ( .A(n8475), .ZN(n8476) );
  XNOR2_X1 U9652 ( .A(n9123), .B(n6764), .ZN(n8479) );
  AND2_X1 U9653 ( .A1(n8762), .A2(n8531), .ZN(n8478) );
  NOR2_X1 U9654 ( .A1(n8479), .A2(n8478), .ZN(n8480) );
  AOI21_X1 U9655 ( .B1(n8479), .B2(n8478), .A(n8480), .ZN(n8682) );
  XNOR2_X1 U9656 ( .A(n9119), .B(n6764), .ZN(n8482) );
  AND2_X1 U9657 ( .A1(n9015), .A2(n8531), .ZN(n8481) );
  NOR2_X1 U9658 ( .A1(n8482), .A2(n8481), .ZN(n8483) );
  AOI21_X1 U9659 ( .B1(n8482), .B2(n8481), .A(n8483), .ZN(n8608) );
  INV_X1 U9660 ( .A(n8483), .ZN(n8484) );
  XNOR2_X1 U9661 ( .A(n9114), .B(n6764), .ZN(n8486) );
  AND2_X1 U9662 ( .A1(n8965), .A2(n8531), .ZN(n8485) );
  NOR2_X1 U9663 ( .A1(n8486), .A2(n8485), .ZN(n8617) );
  NAND2_X1 U9664 ( .A1(n8486), .A2(n8485), .ZN(n8618) );
  XNOR2_X1 U9665 ( .A(n9108), .B(n6765), .ZN(n8487) );
  NAND2_X1 U9666 ( .A1(n8695), .A2(n8531), .ZN(n8488) );
  NAND2_X1 U9667 ( .A1(n8487), .A2(n8488), .ZN(n8660) );
  INV_X1 U9668 ( .A(n8487), .ZN(n8490) );
  INV_X1 U9669 ( .A(n8488), .ZN(n8489) );
  NAND2_X1 U9670 ( .A1(n8490), .A2(n8489), .ZN(n8656) );
  XNOR2_X1 U9671 ( .A(n9103), .B(n6765), .ZN(n8492) );
  NAND2_X1 U9672 ( .A1(n8964), .A2(n8531), .ZN(n8491) );
  XNOR2_X1 U9673 ( .A(n8492), .B(n8491), .ZN(n8582) );
  XNOR2_X1 U9674 ( .A(n9096), .B(n6765), .ZN(n8494) );
  NAND2_X1 U9675 ( .A1(n8920), .A2(n8531), .ZN(n8493) );
  NOR2_X1 U9676 ( .A1(n8494), .A2(n8493), .ZN(n8495) );
  AOI21_X1 U9677 ( .B1(n8494), .B2(n8493), .A(n8495), .ZN(n8638) );
  INV_X1 U9678 ( .A(n8495), .ZN(n8496) );
  XNOR2_X1 U9679 ( .A(n9091), .B(n6764), .ZN(n8498) );
  INV_X1 U9680 ( .A(n8498), .ZN(n8500) );
  AND2_X1 U9681 ( .A1(n8935), .A2(n8531), .ZN(n8497) );
  INV_X1 U9682 ( .A(n8497), .ZN(n8499) );
  AOI21_X1 U9683 ( .B1(n8500), .B2(n8499), .A(n8504), .ZN(n8592) );
  XNOR2_X1 U9684 ( .A(n9081), .B(n6765), .ZN(n8510) );
  INV_X1 U9685 ( .A(n8510), .ZN(n8501) );
  XNOR2_X1 U9686 ( .A(n9086), .B(n6764), .ZN(n8508) );
  NOR2_X1 U9687 ( .A1(n8772), .A2(n6757), .ZN(n8515) );
  INV_X1 U9688 ( .A(n8515), .ZN(n8502) );
  NAND2_X1 U9689 ( .A1(n8514), .A2(n8502), .ZN(n8505) );
  NAND2_X1 U9690 ( .A1(n8501), .A2(n8505), .ZN(n8516) );
  INV_X1 U9691 ( .A(n8504), .ZN(n8513) );
  AOI21_X1 U9692 ( .B1(n8513), .B2(n8502), .A(n8514), .ZN(n8503) );
  AOI21_X1 U9693 ( .B1(n8515), .B2(n8504), .A(n8503), .ZN(n8506) );
  MUX2_X1 U9694 ( .A(n8506), .B(n8505), .S(n8510), .Z(n8507) );
  NAND2_X1 U9695 ( .A1(n8508), .A2(n8515), .ZN(n8509) );
  NAND4_X1 U9696 ( .A1(n8590), .A2(n8513), .A3(n8510), .A4(n8509), .ZN(n8511)
         );
  NOR2_X1 U9697 ( .A1(n8773), .A2(n6757), .ZN(n8573) );
  NAND2_X1 U9698 ( .A1(n8590), .A2(n8513), .ZN(n8645) );
  XOR2_X1 U9699 ( .A(n8515), .B(n8514), .Z(n8646) );
  NOR2_X1 U9700 ( .A1(n8645), .A2(n8646), .ZN(n8644) );
  XNOR2_X1 U9701 ( .A(n9076), .B(n6765), .ZN(n8517) );
  NOR2_X1 U9702 ( .A1(n8601), .A2(n6757), .ZN(n8630) );
  INV_X1 U9703 ( .A(n8517), .ZN(n8518) );
  NAND2_X1 U9704 ( .A1(n8519), .A2(n8518), .ZN(n8520) );
  NAND2_X1 U9705 ( .A1(n8629), .A2(n8520), .ZN(n8600) );
  XNOR2_X1 U9706 ( .A(n9071), .B(n6765), .ZN(n8522) );
  OR2_X1 U9707 ( .A1(n8672), .A2(n6757), .ZN(n8521) );
  NOR2_X1 U9708 ( .A1(n8522), .A2(n8521), .ZN(n8523) );
  AOI21_X1 U9709 ( .B1(n8522), .B2(n8521), .A(n8523), .ZN(n8599) );
  NAND2_X1 U9710 ( .A1(n8600), .A2(n8599), .ZN(n8598) );
  INV_X1 U9711 ( .A(n8523), .ZN(n8524) );
  NAND2_X1 U9712 ( .A1(n8598), .A2(n8524), .ZN(n8671) );
  XNOR2_X1 U9713 ( .A(n9065), .B(n6765), .ZN(n8526) );
  NAND2_X1 U9714 ( .A1(n8826), .A2(n8531), .ZN(n8525) );
  NOR2_X1 U9715 ( .A1(n8526), .A2(n8525), .ZN(n8527) );
  AOI21_X1 U9716 ( .B1(n8526), .B2(n8525), .A(n8527), .ZN(n8670) );
  XNOR2_X1 U9717 ( .A(n9059), .B(n6765), .ZN(n8529) );
  NAND2_X1 U9718 ( .A1(n8779), .A2(n8531), .ZN(n8528) );
  NOR2_X1 U9719 ( .A1(n8529), .A2(n8528), .ZN(n8530) );
  AOI21_X1 U9720 ( .B1(n8529), .B2(n8528), .A(n8530), .ZN(n8566) );
  NAND2_X1 U9721 ( .A1(n8531), .A2(n6765), .ZN(n8532) );
  OR2_X1 U9722 ( .A1(n8787), .A2(n8532), .ZN(n8534) );
  NAND2_X1 U9723 ( .A1(n8787), .A2(n6764), .ZN(n8533) );
  NAND2_X1 U9724 ( .A1(n8534), .A2(n8533), .ZN(n8537) );
  NOR3_X1 U9725 ( .A1(n8803), .A2(n9124), .A3(n8537), .ZN(n8535) );
  AOI21_X1 U9726 ( .B1(n8803), .B2(n8537), .A(n8535), .ZN(n8540) );
  NAND3_X1 U9727 ( .A1(n9054), .A2(n8537), .A3(n10860), .ZN(n8536) );
  OAI21_X1 U9728 ( .B1(n9054), .B2(n8537), .A(n8536), .ZN(n8538) );
  OAI21_X1 U9729 ( .B1(n8803), .B2(n8693), .A(n8667), .ZN(n8539) );
  OAI22_X1 U9730 ( .A1(n8807), .A2(n8688), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10292), .ZN(n8542) );
  NOR2_X1 U9731 ( .A1(n8809), .A2(n8555), .ZN(n8541) );
  AOI211_X1 U9732 ( .C1(n8690), .C2(n8801), .A(n8542), .B(n8541), .ZN(n8543)
         );
  NAND2_X1 U9733 ( .A1(n8544), .A2(n8543), .ZN(P2_U3222) );
  OAI222_X1 U9734 ( .A1(n8547), .A2(P2_U3152), .B1(n9153), .B2(n8546), .C1(
        n8545), .C2(n9151), .ZN(P2_U3338) );
  OAI222_X1 U9735 ( .A1(n8550), .A2(P2_U3152), .B1(n9153), .B2(n8549), .C1(
        n8548), .C2(n9151), .ZN(P2_U3328) );
  XOR2_X1 U9736 ( .A(n8552), .B(n8551), .Z(n8553) );
  NAND2_X1 U9737 ( .A1(n8553), .A2(n8683), .ZN(n8565) );
  OAI22_X1 U9738 ( .A1(n8556), .A2(n8555), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8554), .ZN(n8559) );
  NOR2_X1 U9739 ( .A1(n8557), .A2(n8688), .ZN(n8558) );
  NOR2_X1 U9740 ( .A1(n8559), .A2(n8558), .ZN(n8564) );
  NAND2_X1 U9741 ( .A1(n8651), .A2(n8560), .ZN(n8563) );
  NAND2_X1 U9742 ( .A1(n8690), .A2(n8561), .ZN(n8562) );
  NAND4_X1 U9743 ( .A1(n8565), .A2(n8564), .A3(n8563), .A4(n8562), .ZN(
        P2_U3215) );
  INV_X1 U9744 ( .A(n9059), .ZN(n8823) );
  INV_X1 U9745 ( .A(n8787), .ZN(n8827) );
  NOR2_X1 U9746 ( .A1(n8820), .A2(n8674), .ZN(n8569) );
  OAI22_X1 U9747 ( .A1(n8602), .A2(n8688), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8567), .ZN(n8568) );
  AOI211_X1 U9748 ( .C1(n8827), .C2(n8685), .A(n8569), .B(n8568), .ZN(n8570)
         );
  OAI211_X1 U9749 ( .C1(n8823), .C2(n8693), .A(n8571), .B(n8570), .ZN(P2_U3216) );
  INV_X1 U9750 ( .A(n9081), .ZN(n8774) );
  OAI211_X1 U9751 ( .C1(n8574), .C2(n8573), .A(n8572), .B(n8683), .ZN(n8580)
         );
  OR2_X1 U9752 ( .A1(n8601), .A2(n8808), .ZN(n8576) );
  INV_X1 U9753 ( .A(n8772), .ZN(n8919) );
  NAND2_X1 U9754 ( .A1(n8919), .A2(n9012), .ZN(n8575) );
  NAND2_X1 U9755 ( .A1(n8576), .A2(n8575), .ZN(n8881) );
  INV_X1 U9756 ( .A(n8881), .ZN(n8577) );
  OAI22_X1 U9757 ( .A1(n8577), .A2(n8612), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10291), .ZN(n8578) );
  AOI21_X1 U9758 ( .B1(n8883), .B2(n8690), .A(n8578), .ZN(n8579) );
  OAI211_X1 U9759 ( .C1(n8774), .C2(n8693), .A(n8580), .B(n8579), .ZN(P2_U3218) );
  AOI21_X1 U9760 ( .B1(n8582), .B2(n8654), .A(n8581), .ZN(n8589) );
  INV_X1 U9761 ( .A(n8583), .ZN(n8950) );
  NAND2_X1 U9762 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8739) );
  NAND2_X1 U9763 ( .A1(n8695), .A2(n9012), .ZN(n8585) );
  NAND2_X1 U9764 ( .A1(n8920), .A2(n9014), .ZN(n8584) );
  NAND2_X1 U9765 ( .A1(n8585), .A2(n8584), .ZN(n8945) );
  NAND2_X1 U9766 ( .A1(n8945), .A2(n8676), .ZN(n8586) );
  OAI211_X1 U9767 ( .C1(n8674), .C2(n8950), .A(n8739), .B(n8586), .ZN(n8587)
         );
  AOI21_X1 U9768 ( .B1(n9103), .B2(n8651), .A(n8587), .ZN(n8588) );
  OAI21_X1 U9769 ( .B1(n8589), .B2(n8667), .A(n8588), .ZN(P2_U3221) );
  INV_X1 U9770 ( .A(n9091), .ZN(n8915) );
  OAI211_X1 U9771 ( .C1(n8592), .C2(n8591), .A(n8590), .B(n8683), .ZN(n8597)
         );
  AOI22_X1 U9772 ( .A1(n8919), .A2(n8685), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n8593) );
  OAI21_X1 U9773 ( .B1(n8594), .B2(n8688), .A(n8593), .ZN(n8595) );
  AOI21_X1 U9774 ( .B1(n8913), .B2(n8690), .A(n8595), .ZN(n8596) );
  OAI211_X1 U9775 ( .C1(n8915), .C2(n8693), .A(n8597), .B(n8596), .ZN(P2_U3225) );
  OAI211_X1 U9776 ( .C1(n8600), .C2(n8599), .A(n8598), .B(n8683), .ZN(n8605)
         );
  OAI22_X1 U9777 ( .A1(n8602), .A2(n8808), .B1(n8601), .B2(n8806), .ZN(n9070)
         );
  INV_X1 U9778 ( .A(n9070), .ZN(n8851) );
  OAI22_X1 U9779 ( .A1(n8851), .A2(n8612), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10309), .ZN(n8603) );
  AOI21_X1 U9780 ( .B1(n8852), .B2(n8690), .A(n8603), .ZN(n8604) );
  OAI211_X1 U9781 ( .C1(n5327), .C2(n8693), .A(n8605), .B(n8604), .ZN(P2_U3227) );
  INV_X1 U9782 ( .A(n9119), .ZN(n8991) );
  OAI21_X1 U9783 ( .B1(n8608), .B2(n8607), .A(n8606), .ZN(n8609) );
  NAND2_X1 U9784 ( .A1(n8609), .A2(n8683), .ZN(n8616) );
  NAND2_X1 U9785 ( .A1(n8965), .A2(n9014), .ZN(n8611) );
  NAND2_X1 U9786 ( .A1(n8762), .A2(n9012), .ZN(n8610) );
  NAND2_X1 U9787 ( .A1(n8611), .A2(n8610), .ZN(n8994) );
  INV_X1 U9788 ( .A(n8994), .ZN(n8613) );
  OAI22_X1 U9789 ( .A1(n8613), .A2(n8612), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10308), .ZN(n8614) );
  AOI21_X1 U9790 ( .B1(n8997), .B2(n8690), .A(n8614), .ZN(n8615) );
  OAI211_X1 U9791 ( .C1(n8991), .C2(n8693), .A(n8616), .B(n8615), .ZN(P2_U3228) );
  INV_X1 U9792 ( .A(n8617), .ZN(n8619) );
  NAND2_X1 U9793 ( .A1(n8619), .A2(n8618), .ZN(n8620) );
  XNOR2_X1 U9794 ( .A(n8621), .B(n8620), .ZN(n8628) );
  INV_X1 U9795 ( .A(n8622), .ZN(n8982) );
  NAND2_X1 U9796 ( .A1(n9015), .A2(n9012), .ZN(n8624) );
  NAND2_X1 U9797 ( .A1(n8695), .A2(n9014), .ZN(n8623) );
  NAND2_X1 U9798 ( .A1(n8624), .A2(n8623), .ZN(n8975) );
  AOI22_X1 U9799 ( .A1(n8975), .A2(n8676), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3152), .ZN(n8625) );
  OAI21_X1 U9800 ( .B1(n8674), .B2(n8982), .A(n8625), .ZN(n8626) );
  AOI21_X1 U9801 ( .B1(n9114), .B2(n8651), .A(n8626), .ZN(n8627) );
  OAI21_X1 U9802 ( .B1(n8628), .B2(n8667), .A(n8627), .ZN(P2_U3230) );
  OAI211_X1 U9803 ( .C1(n8631), .C2(n8630), .A(n8629), .B(n8683), .ZN(n8636)
         );
  INV_X1 U9804 ( .A(n8632), .ZN(n8864) );
  AOI22_X1 U9805 ( .A1(n8872), .A2(n8685), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3152), .ZN(n8633) );
  OAI21_X1 U9806 ( .B1(n8773), .B2(n8688), .A(n8633), .ZN(n8634) );
  AOI21_X1 U9807 ( .B1(n8864), .B2(n8690), .A(n8634), .ZN(n8635) );
  OAI211_X1 U9808 ( .C1(n8866), .C2(n8693), .A(n8636), .B(n8635), .ZN(P2_U3231) );
  INV_X1 U9809 ( .A(n9096), .ZN(n8931) );
  OAI211_X1 U9810 ( .C1(n8639), .C2(n8638), .A(n8637), .B(n8683), .ZN(n8643)
         );
  AOI22_X1 U9811 ( .A1(n8685), .A2(n8935), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8640) );
  OAI21_X1 U9812 ( .B1(n8769), .B2(n8688), .A(n8640), .ZN(n8641) );
  AOI21_X1 U9813 ( .B1(n8929), .B2(n8690), .A(n8641), .ZN(n8642) );
  OAI211_X1 U9814 ( .C1(n8931), .C2(n8693), .A(n8643), .B(n8642), .ZN(P2_U3235) );
  AOI21_X1 U9815 ( .B1(n8646), .B2(n8645), .A(n8644), .ZN(n8653) );
  NOR2_X1 U9816 ( .A1(n8674), .A2(n8898), .ZN(n8650) );
  INV_X1 U9817 ( .A(n8773), .ZN(n8905) );
  AOI22_X1 U9818 ( .A1(n8905), .A2(n8685), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8647) );
  OAI21_X1 U9819 ( .B1(n8648), .B2(n8688), .A(n8647), .ZN(n8649) );
  AOI211_X1 U9820 ( .C1(n9086), .C2(n8651), .A(n8650), .B(n8649), .ZN(n8652)
         );
  OAI21_X1 U9821 ( .B1(n8653), .B2(n8667), .A(n8652), .ZN(P2_U3237) );
  INV_X1 U9822 ( .A(n8654), .ZN(n8661) );
  INV_X1 U9823 ( .A(n8655), .ZN(n8657) );
  NAND2_X1 U9824 ( .A1(n8657), .A2(n8656), .ZN(n8659) );
  AOI22_X1 U9825 ( .A1(n8661), .A2(n8660), .B1(n8659), .B2(n8658), .ZN(n8668)
         );
  NAND2_X1 U9826 ( .A1(n8685), .A2(n8964), .ZN(n8663) );
  NAND2_X1 U9827 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8709) );
  OAI211_X1 U9828 ( .C1(n8764), .C2(n8688), .A(n8663), .B(n8709), .ZN(n8665)
         );
  NOR2_X1 U9829 ( .A1(n8960), .A2(n8693), .ZN(n8664) );
  AOI211_X1 U9830 ( .C1(n8690), .C2(n8958), .A(n8665), .B(n8664), .ZN(n8666)
         );
  OAI21_X1 U9831 ( .B1(n8668), .B2(n8667), .A(n8666), .ZN(P2_U3240) );
  INV_X1 U9832 ( .A(n9065), .ZN(n8679) );
  OAI211_X1 U9833 ( .C1(n8671), .C2(n8670), .A(n8669), .B(n8683), .ZN(n8678)
         );
  OAI22_X1 U9834 ( .A1(n8807), .A2(n8808), .B1(n8672), .B2(n8806), .ZN(n8836)
         );
  OAI22_X1 U9835 ( .A1(n8674), .A2(n8840), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8673), .ZN(n8675) );
  AOI21_X1 U9836 ( .B1(n8836), .B2(n8676), .A(n8675), .ZN(n8677) );
  OAI211_X1 U9837 ( .C1(n8679), .C2(n8693), .A(n8678), .B(n8677), .ZN(P2_U3242) );
  INV_X1 U9838 ( .A(n9123), .ZN(n9009) );
  OAI21_X1 U9839 ( .B1(n8682), .B2(n8681), .A(n8680), .ZN(n8684) );
  NAND2_X1 U9840 ( .A1(n8684), .A2(n8683), .ZN(n8692) );
  NAND2_X1 U9841 ( .A1(n8685), .A2(n9015), .ZN(n8687) );
  OAI211_X1 U9842 ( .C1(n8761), .C2(n8688), .A(n8687), .B(n8686), .ZN(n8689)
         );
  AOI21_X1 U9843 ( .B1(n9006), .B2(n8690), .A(n8689), .ZN(n8691) );
  OAI211_X1 U9844 ( .C1(n9009), .C2(n8693), .A(n8692), .B(n8691), .ZN(P2_U3243) );
  MUX2_X1 U9845 ( .A(n8694), .B(P2_DATAO_REG_31__SCAN_IN), .S(n8708), .Z(
        P2_U3583) );
  MUX2_X1 U9846 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8827), .S(P2_U3966), .Z(
        P2_U3580) );
  MUX2_X1 U9847 ( .A(n8779), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8708), .Z(
        P2_U3579) );
  MUX2_X1 U9848 ( .A(n8826), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8708), .Z(
        P2_U3578) );
  MUX2_X1 U9849 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8872), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U9850 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8775), .S(P2_U3966), .Z(
        P2_U3576) );
  MUX2_X1 U9851 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8905), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U9852 ( .A(n8919), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8708), .Z(
        P2_U3574) );
  MUX2_X1 U9853 ( .A(n8935), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8708), .Z(
        P2_U3573) );
  MUX2_X1 U9854 ( .A(n8920), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8708), .Z(
        P2_U3572) );
  MUX2_X1 U9855 ( .A(n8964), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8708), .Z(
        P2_U3571) );
  MUX2_X1 U9856 ( .A(n8695), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8708), .Z(
        P2_U3570) );
  MUX2_X1 U9857 ( .A(n8965), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8708), .Z(
        P2_U3569) );
  MUX2_X1 U9858 ( .A(n9015), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8708), .Z(
        P2_U3568) );
  MUX2_X1 U9859 ( .A(n8762), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8708), .Z(
        P2_U3567) );
  MUX2_X1 U9860 ( .A(n9013), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8708), .Z(
        P2_U3566) );
  MUX2_X1 U9861 ( .A(n8696), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8708), .Z(
        P2_U3565) );
  MUX2_X1 U9862 ( .A(n8697), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8708), .Z(
        P2_U3564) );
  MUX2_X1 U9863 ( .A(n8698), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8708), .Z(
        P2_U3563) );
  MUX2_X1 U9864 ( .A(n8699), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8708), .Z(
        P2_U3562) );
  MUX2_X1 U9865 ( .A(n8700), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8708), .Z(
        P2_U3561) );
  MUX2_X1 U9866 ( .A(n8701), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8708), .Z(
        P2_U3560) );
  MUX2_X1 U9867 ( .A(n8702), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8708), .Z(
        P2_U3559) );
  MUX2_X1 U9868 ( .A(n8703), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8708), .Z(
        P2_U3558) );
  MUX2_X1 U9869 ( .A(n8704), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8708), .Z(
        P2_U3557) );
  MUX2_X1 U9870 ( .A(n8705), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8708), .Z(
        P2_U3556) );
  MUX2_X1 U9871 ( .A(n8706), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8708), .Z(
        P2_U3555) );
  MUX2_X1 U9872 ( .A(n6704), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8708), .Z(
        P2_U3554) );
  MUX2_X1 U9873 ( .A(n8707), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8708), .Z(
        P2_U3553) );
  INV_X1 U9874 ( .A(n8709), .ZN(n8718) );
  INV_X1 U9875 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8712) );
  OAI21_X1 U9876 ( .B1(n8712), .B2(n8711), .A(n8710), .ZN(n8715) );
  INV_X1 U9877 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8713) );
  NAND2_X1 U9878 ( .A1(n8727), .A2(n8713), .ZN(n8733) );
  OAI21_X1 U9879 ( .B1(n8727), .B2(n8713), .A(n8733), .ZN(n8714) );
  NOR2_X1 U9880 ( .A1(n8714), .A2(n8715), .ZN(n8735) );
  AOI21_X1 U9881 ( .B1(n8715), .B2(n8714), .A(n8735), .ZN(n8716) );
  NOR2_X1 U9882 ( .A1(n8716), .A2(n10586), .ZN(n8717) );
  AOI211_X1 U9883 ( .C1(n10606), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n8718), .B(
        n8717), .ZN(n8726) );
  MUX2_X1 U9884 ( .A(n8123), .B(P2_REG2_REG_18__SCAN_IN), .S(n8729), .Z(n8721)
         );
  INV_X1 U9885 ( .A(n8721), .ZN(n8722) );
  NAND2_X1 U9886 ( .A1(n8722), .A2(n8723), .ZN(n8728) );
  OAI21_X1 U9887 ( .B1(n8723), .B2(n8722), .A(n8728), .ZN(n8724) );
  NAND2_X1 U9888 ( .A1(n10584), .A2(n8724), .ZN(n8725) );
  OAI211_X1 U9889 ( .C1(n10585), .C2(n8727), .A(n8726), .B(n8725), .ZN(
        P2_U3263) );
  OAI21_X1 U9890 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n8729), .A(n8728), .ZN(
        n8732) );
  XNOR2_X1 U9891 ( .A(n6499), .B(n8730), .ZN(n8731) );
  XNOR2_X1 U9892 ( .A(n8732), .B(n8731), .ZN(n8743) );
  INV_X1 U9893 ( .A(n8733), .ZN(n8734) );
  NOR2_X1 U9894 ( .A1(n8735), .A2(n8734), .ZN(n8737) );
  XNOR2_X1 U9895 ( .A(n6499), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8736) );
  XNOR2_X1 U9896 ( .A(n8737), .B(n8736), .ZN(n8740) );
  NAND2_X1 U9897 ( .A1(n10606), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8738) );
  OAI211_X1 U9898 ( .C1(n8740), .C2(n10586), .A(n8739), .B(n8738), .ZN(n8741)
         );
  AOI21_X1 U9899 ( .B1(n5256), .B2(n10613), .A(n8741), .ZN(n8742) );
  OAI21_X1 U9900 ( .B1(n10607), .B2(n8743), .A(n8742), .ZN(P2_U3264) );
  INV_X1 U9901 ( .A(n9086), .ZN(n8901) );
  NAND2_X1 U9902 ( .A1(n8823), .A2(n8838), .ZN(n8817) );
  NAND2_X1 U9903 ( .A1(n8747), .A2(P2_B_REG_SCAN_IN), .ZN(n8748) );
  NAND2_X1 U9904 ( .A1(n9014), .A2(n8748), .ZN(n8790) );
  NOR2_X1 U9905 ( .A1(n8749), .A2(n8790), .ZN(n9043) );
  NAND2_X1 U9906 ( .A1(n10811), .A2(n9043), .ZN(n8754) );
  OAI21_X1 U9907 ( .B1(n10811), .B2(n8750), .A(n8754), .ZN(n8751) );
  AOI21_X1 U9908 ( .B1(n8746), .B2(n9035), .A(n8751), .ZN(n8752) );
  OAI21_X1 U9909 ( .B1(n9041), .B2(n8793), .A(n8752), .ZN(P2_U3265) );
  AOI21_X1 U9910 ( .B1(n8757), .B2(n8792), .A(n8753), .ZN(n9042) );
  INV_X1 U9911 ( .A(n9042), .ZN(n8759) );
  OAI21_X1 U9912 ( .B1(n10811), .B2(n8755), .A(n8754), .ZN(n8756) );
  AOI21_X1 U9913 ( .B1(n8757), .B2(n9035), .A(n8756), .ZN(n8758) );
  OAI21_X1 U9914 ( .B1(n8759), .B2(n8793), .A(n8758), .ZN(P2_U3266) );
  NAND2_X1 U9915 ( .A1(n8765), .A2(n8764), .ZN(n8766) );
  NAND2_X1 U9916 ( .A1(n8777), .A2(n8776), .ZN(n8832) );
  NAND2_X1 U9917 ( .A1(n8823), .A2(n8807), .ZN(n8780) );
  NAND2_X1 U9918 ( .A1(n8800), .A2(n8781), .ZN(n8782) );
  NAND2_X1 U9919 ( .A1(n8782), .A2(n5625), .ZN(n8784) );
  XNOR2_X1 U9920 ( .A(n8784), .B(n8783), .ZN(n9047) );
  INV_X1 U9921 ( .A(n9047), .ZN(n8799) );
  XOR2_X1 U9922 ( .A(n8786), .B(n8783), .Z(n8788) );
  OAI222_X1 U9923 ( .A1(n8790), .A2(n8789), .B1(n8788), .B2(n10797), .C1(n8806), .C2(n8787), .ZN(n9051) );
  INV_X1 U9924 ( .A(n8791), .ZN(n9048) );
  OAI21_X1 U9925 ( .B1(n9048), .B2(n5315), .A(n8792), .ZN(n9049) );
  NOR2_X1 U9926 ( .A1(n9049), .A2(n8793), .ZN(n8797) );
  AOI22_X1 U9927 ( .A1(n8794), .A2(n10801), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n10813), .ZN(n8795) );
  OAI21_X1 U9928 ( .B1(n9048), .B2(n9008), .A(n8795), .ZN(n8796) );
  AOI211_X1 U9929 ( .C1(n9051), .C2(n10811), .A(n8797), .B(n8796), .ZN(n8798)
         );
  OAI21_X1 U9930 ( .B1(n8799), .B2(n9022), .A(n8798), .ZN(P2_U3267) );
  XNOR2_X1 U9931 ( .A(n8800), .B(n8804), .ZN(n9058) );
  XNOR2_X1 U9932 ( .A(n8803), .B(n8817), .ZN(n9055) );
  AOI22_X1 U9933 ( .A1(n8801), .A2(n10801), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n10813), .ZN(n8802) );
  OAI21_X1 U9934 ( .B1(n8803), .B2(n9008), .A(n8802), .ZN(n8813) );
  XNOR2_X1 U9935 ( .A(n8805), .B(n8804), .ZN(n8811) );
  OAI22_X1 U9936 ( .A1(n8809), .A2(n8808), .B1(n8807), .B2(n8806), .ZN(n8810)
         );
  AOI21_X1 U9937 ( .B1(n8811), .B2(n9017), .A(n8810), .ZN(n9057) );
  NOR2_X1 U9938 ( .A1(n9057), .A2(n10813), .ZN(n8812) );
  AOI211_X1 U9939 ( .C1(n9020), .C2(n9055), .A(n8813), .B(n8812), .ZN(n8814)
         );
  OAI21_X1 U9940 ( .B1(n9058), .B2(n9022), .A(n8814), .ZN(P2_U3268) );
  XNOR2_X1 U9941 ( .A(n8815), .B(n8816), .ZN(n9063) );
  INV_X1 U9942 ( .A(n8838), .ZN(n8819) );
  INV_X1 U9943 ( .A(n8817), .ZN(n8818) );
  AOI21_X1 U9944 ( .B1(n9059), .B2(n8819), .A(n8818), .ZN(n9060) );
  INV_X1 U9945 ( .A(n8820), .ZN(n8821) );
  AOI22_X1 U9946 ( .A1(n8821), .A2(n10801), .B1(n10813), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8822) );
  OAI21_X1 U9947 ( .B1(n8823), .B2(n9008), .A(n8822), .ZN(n8830) );
  XNOR2_X1 U9948 ( .A(n8825), .B(n8824), .ZN(n8828) );
  AOI211_X1 U9949 ( .C1(n9020), .C2(n9060), .A(n8830), .B(n8829), .ZN(n8831)
         );
  OAI21_X1 U9950 ( .B1(n9063), .B2(n9022), .A(n8831), .ZN(P2_U3269) );
  XOR2_X1 U9951 ( .A(n8834), .B(n8832), .Z(n9068) );
  AOI22_X1 U9952 ( .A1(n9065), .A2(n9035), .B1(P2_REG2_REG_26__SCAN_IN), .B2(
        n10813), .ZN(n8843) );
  NAND2_X1 U9953 ( .A1(n8848), .A2(n8833), .ZN(n8835) );
  XNOR2_X1 U9954 ( .A(n8835), .B(n8834), .ZN(n8837) );
  AOI21_X1 U9955 ( .B1(n8837), .B2(n9017), .A(n8836), .ZN(n9067) );
  AOI211_X1 U9956 ( .C1(n9065), .C2(n8846), .A(n10862), .B(n8838), .ZN(n9064)
         );
  NAND2_X1 U9957 ( .A1(n9064), .A2(n6499), .ZN(n8839) );
  OAI211_X1 U9958 ( .C1(n8981), .C2(n8840), .A(n9067), .B(n8839), .ZN(n8841)
         );
  NAND2_X1 U9959 ( .A1(n8841), .A2(n10811), .ZN(n8842) );
  OAI211_X1 U9960 ( .C1(n9068), .C2(n9022), .A(n8843), .B(n8842), .ZN(P2_U3270) );
  XNOR2_X1 U9961 ( .A(n8845), .B(n8844), .ZN(n9069) );
  INV_X1 U9962 ( .A(n9069), .ZN(n8857) );
  AOI21_X1 U9963 ( .B1(n9071), .B2(n8862), .A(n10862), .ZN(n8847) );
  NAND2_X1 U9964 ( .A1(n8847), .A2(n8846), .ZN(n9072) );
  OAI211_X1 U9965 ( .C1(n8850), .C2(n8849), .A(n9017), .B(n8848), .ZN(n9073)
         );
  OAI211_X1 U9966 ( .C1(n5256), .C2(n9072), .A(n9073), .B(n8851), .ZN(n8855)
         );
  AOI22_X1 U9967 ( .A1(n10813), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8852), .B2(
        n10801), .ZN(n8853) );
  OAI21_X1 U9968 ( .B1(n5327), .B2(n9008), .A(n8853), .ZN(n8854) );
  AOI21_X1 U9969 ( .B1(n8855), .B2(n10811), .A(n8854), .ZN(n8856) );
  OAI21_X1 U9970 ( .B1(n8857), .B2(n9022), .A(n8856), .ZN(P2_U3271) );
  INV_X1 U9971 ( .A(n8870), .ZN(n8861) );
  INV_X1 U9972 ( .A(n8858), .ZN(n8859) );
  AOI21_X1 U9973 ( .B1(n8861), .B2(n8860), .A(n8859), .ZN(n9080) );
  INV_X1 U9974 ( .A(n8862), .ZN(n8863) );
  AOI21_X1 U9975 ( .B1(n9076), .B2(n5331), .A(n8863), .ZN(n9077) );
  AOI22_X1 U9976 ( .A1(n10813), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8864), .B2(
        n10801), .ZN(n8865) );
  OAI21_X1 U9977 ( .B1(n8866), .B2(n9008), .A(n8865), .ZN(n8874) );
  NAND2_X1 U9978 ( .A1(n8867), .A2(n8868), .ZN(n8869) );
  XOR2_X1 U9979 ( .A(n8870), .B(n8869), .Z(n8871) );
  AOI222_X1 U9980 ( .A1(n8905), .A2(n9012), .B1(n8872), .B2(n9014), .C1(n9017), 
        .C2(n8871), .ZN(n9079) );
  NOR2_X1 U9981 ( .A1(n9079), .A2(n10813), .ZN(n8873) );
  AOI211_X1 U9982 ( .C1(n9077), .C2(n9020), .A(n8874), .B(n8873), .ZN(n8875)
         );
  OAI21_X1 U9983 ( .B1(n9080), .B2(n9022), .A(n8875), .ZN(P2_U3272) );
  OAI21_X1 U9984 ( .B1(n8877), .B2(n8878), .A(n8876), .ZN(n9085) );
  NAND2_X1 U9985 ( .A1(n8879), .A2(n8878), .ZN(n8880) );
  NAND2_X1 U9986 ( .A1(n8867), .A2(n8880), .ZN(n8882) );
  AOI21_X1 U9987 ( .B1(n8882), .B2(n9017), .A(n8881), .ZN(n9084) );
  INV_X1 U9988 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8885) );
  INV_X1 U9989 ( .A(n8883), .ZN(n8884) );
  OAI22_X1 U9990 ( .A1(n10811), .A2(n8885), .B1(n8884), .B2(n8981), .ZN(n8886)
         );
  AOI21_X1 U9991 ( .B1(n9081), .B2(n9035), .A(n8886), .ZN(n8890) );
  AND2_X1 U9992 ( .A1(n9081), .A2(n8895), .ZN(n8887) );
  NOR2_X1 U9993 ( .A1(n8888), .A2(n8887), .ZN(n9082) );
  NAND2_X1 U9994 ( .A1(n9082), .A2(n9020), .ZN(n8889) );
  OAI211_X1 U9995 ( .C1(n9084), .C2(n10813), .A(n8890), .B(n8889), .ZN(n8891)
         );
  INV_X1 U9996 ( .A(n8891), .ZN(n8892) );
  OAI21_X1 U9997 ( .B1(n9085), .B2(n9022), .A(n8892), .ZN(P2_U3273) );
  XNOR2_X1 U9998 ( .A(n8894), .B(n8893), .ZN(n9090) );
  INV_X1 U9999 ( .A(n8911), .ZN(n8897) );
  INV_X1 U10000 ( .A(n8895), .ZN(n8896) );
  AOI21_X1 U10001 ( .B1(n9086), .B2(n8897), .A(n8896), .ZN(n9087) );
  INV_X1 U10002 ( .A(n8898), .ZN(n8899) );
  AOI22_X1 U10003 ( .A1(n10813), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8899), 
        .B2(n10801), .ZN(n8900) );
  OAI21_X1 U10004 ( .B1(n8901), .B2(n9008), .A(n8900), .ZN(n8907) );
  XNOR2_X1 U10005 ( .A(n8903), .B(n8902), .ZN(n8904) );
  AOI222_X1 U10006 ( .A1(n8935), .A2(n9012), .B1(n8905), .B2(n9014), .C1(n9017), .C2(n8904), .ZN(n9089) );
  NOR2_X1 U10007 ( .A1(n9089), .A2(n10813), .ZN(n8906) );
  AOI211_X1 U10008 ( .C1(n9087), .C2(n9020), .A(n8907), .B(n8906), .ZN(n8908)
         );
  OAI21_X1 U10009 ( .B1(n9090), .B2(n9022), .A(n8908), .ZN(P2_U3274) );
  OAI21_X1 U10010 ( .B1(n5119), .B2(n8916), .A(n8909), .ZN(n8910) );
  INV_X1 U10011 ( .A(n8910), .ZN(n9095) );
  INV_X1 U10012 ( .A(n8928), .ZN(n8912) );
  AOI21_X1 U10013 ( .B1(n9091), .B2(n8912), .A(n8911), .ZN(n9092) );
  AOI22_X1 U10014 ( .A1(n10813), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8913), 
        .B2(n10801), .ZN(n8914) );
  OAI21_X1 U10015 ( .B1(n8915), .B2(n9008), .A(n8914), .ZN(n8922) );
  XNOR2_X1 U10016 ( .A(n8917), .B(n8916), .ZN(n8918) );
  AOI222_X1 U10017 ( .A1(n8920), .A2(n9012), .B1(n8919), .B2(n9014), .C1(n9017), .C2(n8918), .ZN(n9094) );
  NOR2_X1 U10018 ( .A1(n9094), .A2(n10813), .ZN(n8921) );
  AOI211_X1 U10019 ( .C1(n9092), .C2(n9020), .A(n8922), .B(n8921), .ZN(n8923)
         );
  OAI21_X1 U10020 ( .B1(n9095), .B2(n9022), .A(n8923), .ZN(P2_U3275) );
  OAI21_X1 U10021 ( .B1(n8926), .B2(n8925), .A(n8924), .ZN(n9100) );
  INV_X1 U10022 ( .A(n8927), .ZN(n8948) );
  AOI21_X1 U10023 ( .B1(n9096), .B2(n8948), .A(n8928), .ZN(n9097) );
  AOI22_X1 U10024 ( .A1(n10813), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8929), 
        .B2(n10801), .ZN(n8930) );
  OAI21_X1 U10025 ( .B1(n8931), .B2(n9008), .A(n8930), .ZN(n8939) );
  OAI211_X1 U10026 ( .C1(n8934), .C2(n8933), .A(n8932), .B(n9017), .ZN(n8937)
         );
  AOI22_X1 U10027 ( .A1(n9012), .A2(n8964), .B1(n8935), .B2(n9014), .ZN(n8936)
         );
  AND2_X1 U10028 ( .A1(n8937), .A2(n8936), .ZN(n9099) );
  NOR2_X1 U10029 ( .A1(n9099), .A2(n10813), .ZN(n8938) );
  AOI211_X1 U10030 ( .C1(n9097), .C2(n9020), .A(n8939), .B(n8938), .ZN(n8940)
         );
  OAI21_X1 U10031 ( .B1(n9100), .B2(n9022), .A(n8940), .ZN(P2_U3276) );
  OR2_X1 U10032 ( .A1(n8941), .A2(n8943), .ZN(n9102) );
  NAND3_X1 U10033 ( .A1(n9102), .A2(n9101), .A3(n9033), .ZN(n8955) );
  AOI22_X1 U10034 ( .A1(n9103), .A2(n9035), .B1(P2_REG2_REG_19__SCAN_IN), .B2(
        n10813), .ZN(n8954) );
  INV_X1 U10035 ( .A(n8942), .ZN(n8944) );
  AOI21_X1 U10036 ( .B1(n8944), .B2(n8943), .A(n10797), .ZN(n8947) );
  AOI21_X1 U10037 ( .B1(n8947), .B2(n8946), .A(n8945), .ZN(n9106) );
  INV_X1 U10038 ( .A(n9106), .ZN(n8952) );
  OAI211_X1 U10039 ( .C1(n8949), .C2(n8957), .A(n8948), .B(n10792), .ZN(n9104)
         );
  OAI22_X1 U10040 ( .A1(n9104), .A2(n5256), .B1(n8981), .B2(n8950), .ZN(n8951)
         );
  OAI21_X1 U10041 ( .B1(n8952), .B2(n8951), .A(n10811), .ZN(n8953) );
  NAND3_X1 U10042 ( .A1(n8955), .A2(n8954), .A3(n8953), .ZN(P2_U3277) );
  XNOR2_X1 U10043 ( .A(n8956), .B(n8962), .ZN(n9112) );
  AOI21_X1 U10044 ( .B1(n9108), .B2(n5128), .A(n8957), .ZN(n9109) );
  AOI22_X1 U10045 ( .A1(n10813), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8958), 
        .B2(n10801), .ZN(n8959) );
  OAI21_X1 U10046 ( .B1(n8960), .B2(n9008), .A(n8959), .ZN(n8969) );
  OAI211_X1 U10047 ( .C1(n8963), .C2(n8962), .A(n8961), .B(n9017), .ZN(n8967)
         );
  AOI22_X1 U10048 ( .A1(n9012), .A2(n8965), .B1(n8964), .B2(n9014), .ZN(n8966)
         );
  AND2_X1 U10049 ( .A1(n8967), .A2(n8966), .ZN(n9111) );
  NOR2_X1 U10050 ( .A1(n9111), .A2(n10813), .ZN(n8968) );
  AOI211_X1 U10051 ( .C1(n9109), .C2(n9020), .A(n8969), .B(n8968), .ZN(n8970)
         );
  OAI21_X1 U10052 ( .B1(n9112), .B2(n9022), .A(n8970), .ZN(P2_U3278) );
  OAI21_X1 U10053 ( .B1(n5131), .B2(n8973), .A(n8971), .ZN(n8972) );
  INV_X1 U10054 ( .A(n8972), .ZN(n9117) );
  XNOR2_X1 U10055 ( .A(n8974), .B(n8973), .ZN(n8976) );
  AOI21_X1 U10056 ( .B1(n8976), .B2(n9017), .A(n8975), .ZN(n9116) );
  XNOR2_X1 U10057 ( .A(n8996), .B(n9114), .ZN(n8977) );
  NOR2_X1 U10058 ( .A1(n8977), .A2(n10862), .ZN(n9113) );
  NAND2_X1 U10059 ( .A1(n9113), .A2(n6499), .ZN(n8978) );
  OAI211_X1 U10060 ( .C1(n9117), .C2(n8979), .A(n9116), .B(n8978), .ZN(n8980)
         );
  NAND2_X1 U10061 ( .A1(n8980), .A2(n10811), .ZN(n8986) );
  OAI22_X1 U10062 ( .A1(n10811), .A2(n8983), .B1(n8982), .B2(n8981), .ZN(n8984) );
  AOI21_X1 U10063 ( .B1(n9114), .B2(n9035), .A(n8984), .ZN(n8985) );
  OAI211_X1 U10064 ( .C1(n9117), .C2(n8987), .A(n8986), .B(n8985), .ZN(
        P2_U3279) );
  AOI21_X1 U10065 ( .B1(n8993), .B2(n8989), .A(n8988), .ZN(n8990) );
  INV_X1 U10066 ( .A(n8990), .ZN(n9122) );
  NOR2_X1 U10067 ( .A1(n8991), .A2(n9008), .ZN(n9000) );
  XOR2_X1 U10068 ( .A(n8993), .B(n8992), .Z(n8995) );
  AOI21_X1 U10069 ( .B1(n8995), .B2(n9017), .A(n8994), .ZN(n9121) );
  AOI211_X1 U10070 ( .C1(n9119), .C2(n9003), .A(n10862), .B(n5326), .ZN(n9118)
         );
  AOI22_X1 U10071 ( .A1(n9118), .A2(n6499), .B1(n10801), .B2(n8997), .ZN(n8998) );
  AOI21_X1 U10072 ( .B1(n9121), .B2(n8998), .A(n10813), .ZN(n8999) );
  AOI211_X1 U10073 ( .C1(n10813), .C2(P2_REG2_REG_16__SCAN_IN), .A(n9000), .B(
        n8999), .ZN(n9001) );
  OAI21_X1 U10074 ( .B1(n9122), .B2(n9022), .A(n9001), .ZN(P2_U3280) );
  XNOR2_X1 U10075 ( .A(n9002), .B(n9010), .ZN(n9128) );
  INV_X1 U10076 ( .A(n9003), .ZN(n9004) );
  AOI21_X1 U10077 ( .B1(n9123), .B2(n9005), .A(n9004), .ZN(n9125) );
  AOI22_X1 U10078 ( .A1(n10813), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n9006), 
        .B2(n10801), .ZN(n9007) );
  OAI21_X1 U10079 ( .B1(n9009), .B2(n9008), .A(n9007), .ZN(n9019) );
  XNOR2_X1 U10080 ( .A(n9011), .B(n9010), .ZN(n9016) );
  AOI222_X1 U10081 ( .A1(n9017), .A2(n9016), .B1(n9015), .B2(n9014), .C1(n9013), .C2(n9012), .ZN(n9127) );
  NOR2_X1 U10082 ( .A1(n9127), .A2(n10813), .ZN(n9018) );
  AOI211_X1 U10083 ( .C1(n9125), .C2(n9020), .A(n9019), .B(n9018), .ZN(n9021)
         );
  OAI21_X1 U10084 ( .B1(n9128), .B2(n9022), .A(n9021), .ZN(P2_U3281) );
  XOR2_X1 U10085 ( .A(n9023), .B(n9031), .Z(n9025) );
  OAI21_X1 U10086 ( .B1(n9025), .B2(n10797), .A(n9024), .ZN(n10704) );
  INV_X1 U10087 ( .A(n9026), .ZN(n9028) );
  OAI211_X1 U10088 ( .C1(n9028), .C2(n10702), .A(n10792), .B(n9027), .ZN(
        n10700) );
  NOR2_X1 U10089 ( .A1(n10700), .A2(n5256), .ZN(n9029) );
  OAI21_X1 U10090 ( .B1(n10704), .B2(n9029), .A(n10811), .ZN(n9039) );
  AOI22_X1 U10091 ( .A1(n10813), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n9030), .B2(
        n10801), .ZN(n9038) );
  NAND2_X1 U10092 ( .A1(n9032), .A2(n9031), .ZN(n10699) );
  NAND3_X1 U10093 ( .A1(n5624), .A2(n10699), .A3(n9033), .ZN(n9037) );
  NAND2_X1 U10094 ( .A1(n9035), .A2(n9034), .ZN(n9036) );
  NAND4_X1 U10095 ( .A1(n9039), .A2(n9038), .A3(n9037), .A4(n9036), .ZN(
        P2_U3288) );
  AOI21_X1 U10096 ( .B1(n8746), .B2(n9124), .A(n9043), .ZN(n9040) );
  OAI21_X1 U10097 ( .B1(n9041), .B2(n10862), .A(n9040), .ZN(n9129) );
  MUX2_X1 U10098 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9129), .S(n10870), .Z(
        P2_U3551) );
  NAND2_X1 U10099 ( .A1(n9042), .A2(n10792), .ZN(n9045) );
  INV_X1 U10100 ( .A(n9043), .ZN(n9044) );
  OAI211_X1 U10101 ( .C1(n9046), .C2(n10860), .A(n9045), .B(n9044), .ZN(n9130)
         );
  MUX2_X1 U10102 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9130), .S(n10870), .Z(
        P2_U3550) );
  NAND2_X1 U10103 ( .A1(n9047), .A2(n10866), .ZN(n9053) );
  OAI22_X1 U10104 ( .A1(n9049), .A2(n10862), .B1(n9048), .B2(n10860), .ZN(
        n9050) );
  NOR2_X1 U10105 ( .A1(n9051), .A2(n9050), .ZN(n9052) );
  NAND2_X1 U10106 ( .A1(n9053), .A2(n9052), .ZN(n9131) );
  MUX2_X1 U10107 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9131), .S(n10870), .Z(
        P2_U3549) );
  AOI22_X1 U10108 ( .A1(n9055), .A2(n10792), .B1(n9124), .B2(n9054), .ZN(n9056) );
  OAI211_X1 U10109 ( .C1(n9058), .C2(n10841), .A(n9057), .B(n9056), .ZN(n9132)
         );
  MUX2_X1 U10110 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9132), .S(n10870), .Z(
        P2_U3548) );
  AOI22_X1 U10111 ( .A1(n9060), .A2(n10792), .B1(n9124), .B2(n9059), .ZN(n9061) );
  OAI211_X1 U10112 ( .C1(n9063), .C2(n10841), .A(n9062), .B(n9061), .ZN(n9133)
         );
  MUX2_X1 U10113 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9133), .S(n10870), .Z(
        P2_U3547) );
  AOI21_X1 U10114 ( .B1(n9124), .B2(n9065), .A(n9064), .ZN(n9066) );
  OAI211_X1 U10115 ( .C1(n9068), .C2(n10841), .A(n9067), .B(n9066), .ZN(n9134)
         );
  MUX2_X1 U10116 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9134), .S(n10870), .Z(
        P2_U3546) );
  NAND2_X1 U10117 ( .A1(n9069), .A2(n10866), .ZN(n9075) );
  AOI21_X1 U10118 ( .B1(n9071), .B2(n9124), .A(n9070), .ZN(n9074) );
  NAND4_X1 U10119 ( .A1(n9075), .A2(n9074), .A3(n9073), .A4(n9072), .ZN(n9135)
         );
  MUX2_X1 U10120 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9135), .S(n10870), .Z(
        P2_U3545) );
  AOI22_X1 U10121 ( .A1(n9077), .A2(n10792), .B1(n9124), .B2(n9076), .ZN(n9078) );
  OAI211_X1 U10122 ( .C1(n9080), .C2(n10841), .A(n9079), .B(n9078), .ZN(n9136)
         );
  MUX2_X1 U10123 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9136), .S(n10870), .Z(
        P2_U3544) );
  AOI22_X1 U10124 ( .A1(n9082), .A2(n10792), .B1(n9124), .B2(n9081), .ZN(n9083) );
  OAI211_X1 U10125 ( .C1(n9085), .C2(n10841), .A(n9084), .B(n9083), .ZN(n9137)
         );
  MUX2_X1 U10126 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9137), .S(n10870), .Z(
        P2_U3543) );
  AOI22_X1 U10127 ( .A1(n9087), .A2(n10792), .B1(n9124), .B2(n9086), .ZN(n9088) );
  OAI211_X1 U10128 ( .C1(n9090), .C2(n10841), .A(n9089), .B(n9088), .ZN(n9138)
         );
  MUX2_X1 U10129 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9138), .S(n10870), .Z(
        P2_U3542) );
  AOI22_X1 U10130 ( .A1(n9092), .A2(n10792), .B1(n9124), .B2(n9091), .ZN(n9093) );
  OAI211_X1 U10131 ( .C1(n9095), .C2(n10841), .A(n9094), .B(n9093), .ZN(n9139)
         );
  MUX2_X1 U10132 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9139), .S(n10870), .Z(
        P2_U3541) );
  AOI22_X1 U10133 ( .A1(n9097), .A2(n10792), .B1(n9124), .B2(n9096), .ZN(n9098) );
  OAI211_X1 U10134 ( .C1(n9100), .C2(n10841), .A(n9099), .B(n9098), .ZN(n9140)
         );
  MUX2_X1 U10135 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9140), .S(n10870), .Z(
        P2_U3540) );
  NAND3_X1 U10136 ( .A1(n9102), .A2(n9101), .A3(n10866), .ZN(n9107) );
  NAND2_X1 U10137 ( .A1(n9103), .A2(n9124), .ZN(n9105) );
  NAND4_X1 U10138 ( .A1(n9107), .A2(n9106), .A3(n9105), .A4(n9104), .ZN(n9141)
         );
  MUX2_X1 U10139 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9141), .S(n10870), .Z(
        P2_U3539) );
  AOI22_X1 U10140 ( .A1(n9109), .A2(n10792), .B1(n9124), .B2(n9108), .ZN(n9110) );
  OAI211_X1 U10141 ( .C1(n9112), .C2(n10841), .A(n9111), .B(n9110), .ZN(n9142)
         );
  MUX2_X1 U10142 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9142), .S(n10870), .Z(
        P2_U3538) );
  AOI21_X1 U10143 ( .B1(n9124), .B2(n9114), .A(n9113), .ZN(n9115) );
  OAI211_X1 U10144 ( .C1(n9117), .C2(n10841), .A(n9116), .B(n9115), .ZN(n9143)
         );
  MUX2_X1 U10145 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9143), .S(n10870), .Z(
        P2_U3537) );
  AOI21_X1 U10146 ( .B1(n9124), .B2(n9119), .A(n9118), .ZN(n9120) );
  OAI211_X1 U10147 ( .C1(n9122), .C2(n10841), .A(n9121), .B(n9120), .ZN(n9144)
         );
  MUX2_X1 U10148 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9144), .S(n10870), .Z(
        P2_U3536) );
  AOI22_X1 U10149 ( .A1(n9125), .A2(n10792), .B1(n9124), .B2(n9123), .ZN(n9126) );
  OAI211_X1 U10150 ( .C1(n9128), .C2(n10841), .A(n9127), .B(n9126), .ZN(n9145)
         );
  MUX2_X1 U10151 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9145), .S(n10870), .Z(
        P2_U3535) );
  MUX2_X1 U10152 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9129), .S(n10873), .Z(
        P2_U3519) );
  MUX2_X1 U10153 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9130), .S(n10873), .Z(
        P2_U3518) );
  MUX2_X1 U10154 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9131), .S(n10873), .Z(
        P2_U3517) );
  MUX2_X1 U10155 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9132), .S(n10873), .Z(
        P2_U3516) );
  MUX2_X1 U10156 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9133), .S(n10873), .Z(
        P2_U3515) );
  MUX2_X1 U10157 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9134), .S(n10873), .Z(
        P2_U3514) );
  MUX2_X1 U10158 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9135), .S(n10873), .Z(
        P2_U3513) );
  MUX2_X1 U10159 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9136), .S(n10873), .Z(
        P2_U3512) );
  MUX2_X1 U10160 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9137), .S(n10873), .Z(
        P2_U3511) );
  MUX2_X1 U10161 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9138), .S(n10873), .Z(
        P2_U3510) );
  MUX2_X1 U10162 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9139), .S(n10873), .Z(
        P2_U3509) );
  MUX2_X1 U10163 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9140), .S(n10873), .Z(
        P2_U3508) );
  MUX2_X1 U10164 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9141), .S(n10873), .Z(
        P2_U3507) );
  MUX2_X1 U10165 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9142), .S(n10873), .Z(
        P2_U3505) );
  MUX2_X1 U10166 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9143), .S(n10873), .Z(
        P2_U3502) );
  MUX2_X1 U10167 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9144), .S(n10873), .Z(
        P2_U3499) );
  MUX2_X1 U10168 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9145), .S(n10873), .Z(
        P2_U3496) );
  INV_X1 U10169 ( .A(n9419), .ZN(n10447) );
  NOR4_X1 U10170 ( .A1(n9147), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3152), .A4(
        n9146), .ZN(n9148) );
  AOI21_X1 U10171 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n9149), .A(n9148), .ZN(
        n9150) );
  OAI21_X1 U10172 ( .B1(n10447), .B2(n9153), .A(n9150), .ZN(P2_U3327) );
  INV_X1 U10173 ( .A(n9428), .ZN(n10450) );
  OAI222_X1 U10174 ( .A1(P2_U3152), .A2(n9154), .B1(n9153), .B2(n10450), .C1(
        n9152), .C2(n9151), .ZN(P2_U3329) );
  MUX2_X1 U10175 ( .A(n9155), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  AOI22_X1 U10176 ( .A1(n9963), .A2(n9235), .B1(n9239), .B2(n9776), .ZN(n9225)
         );
  INV_X1 U10177 ( .A(n9225), .ZN(n9227) );
  OAI22_X1 U10178 ( .A1(n9350), .A2(n9289), .B1(n9741), .B2(n9287), .ZN(n9156)
         );
  XNOR2_X1 U10179 ( .A(n9156), .B(n9243), .ZN(n9226) );
  OAI22_X1 U10180 ( .A1(n9846), .A2(n9289), .B1(n9819), .B2(n9287), .ZN(n9157)
         );
  XOR2_X1 U10181 ( .A(n9243), .B(n9157), .Z(n9276) );
  INV_X1 U10182 ( .A(n9276), .ZN(n9197) );
  OR2_X1 U10183 ( .A1(n9403), .A2(n9287), .ZN(n9160) );
  NAND2_X1 U10184 ( .A1(n9161), .A2(n9160), .ZN(n9162) );
  XNOR2_X1 U10185 ( .A(n9162), .B(n9208), .ZN(n9165) );
  NAND2_X1 U10186 ( .A1(n9921), .A2(n9235), .ZN(n9164) );
  OR2_X1 U10187 ( .A1(n9403), .A2(n9286), .ZN(n9163) );
  NAND2_X1 U10188 ( .A1(n9164), .A2(n9163), .ZN(n9256) );
  NAND2_X1 U10189 ( .A1(n9254), .A2(n9256), .ZN(n9167) );
  OR2_X1 U10190 ( .A1(n9336), .A2(n9287), .ZN(n9168) );
  NAND2_X1 U10191 ( .A1(n9169), .A2(n9168), .ZN(n9170) );
  XNOR2_X1 U10192 ( .A(n9170), .B(n9208), .ZN(n9324) );
  NOR2_X1 U10193 ( .A1(n9336), .A2(n9286), .ZN(n9171) );
  AOI21_X1 U10194 ( .B1(n10886), .B2(n9235), .A(n9171), .ZN(n9180) );
  NOR2_X1 U10195 ( .A1(n9887), .A2(n9286), .ZN(n9172) );
  AOI21_X1 U10196 ( .B1(n10876), .B2(n9235), .A(n9172), .ZN(n9397) );
  OR2_X1 U10197 ( .A1(n9887), .A2(n9287), .ZN(n9173) );
  NAND2_X1 U10198 ( .A1(n9174), .A2(n9173), .ZN(n9175) );
  XNOR2_X1 U10199 ( .A(n9175), .B(n9208), .ZN(n9321) );
  OAI22_X1 U10200 ( .A1(n9324), .A2(n9180), .B1(n9397), .B2(n9321), .ZN(n9176)
         );
  INV_X1 U10201 ( .A(n9176), .ZN(n9177) );
  NAND2_X1 U10202 ( .A1(n9321), .A2(n9397), .ZN(n9179) );
  INV_X1 U10203 ( .A(n9180), .ZN(n9323) );
  NAND2_X1 U10204 ( .A1(n9179), .A2(n9323), .ZN(n9182) );
  INV_X1 U10205 ( .A(n9179), .ZN(n9181) );
  AOI22_X1 U10206 ( .A1(n9324), .A2(n9182), .B1(n9181), .B2(n9180), .ZN(n9183)
         );
  OR2_X1 U10207 ( .A1(n9890), .A2(n9287), .ZN(n9184) );
  NAND2_X1 U10208 ( .A1(n9185), .A2(n9184), .ZN(n9186) );
  XNOR2_X1 U10209 ( .A(n9186), .B(n9243), .ZN(n9188) );
  NOR2_X1 U10210 ( .A1(n9890), .A2(n9286), .ZN(n9187) );
  AOI21_X1 U10211 ( .B1(n9998), .B2(n9235), .A(n9187), .ZN(n9189) );
  XNOR2_X1 U10212 ( .A(n9188), .B(n9189), .ZN(n9333) );
  INV_X1 U10213 ( .A(n9188), .ZN(n9190) );
  NAND2_X1 U10214 ( .A1(n9878), .A2(n9235), .ZN(n9191) );
  NAND2_X1 U10215 ( .A1(n9192), .A2(n9191), .ZN(n9193) );
  XNOR2_X1 U10216 ( .A(n9193), .B(n9243), .ZN(n9195) );
  AND2_X1 U10217 ( .A1(n9878), .A2(n9239), .ZN(n9194) );
  AOI21_X1 U10218 ( .B1(n9993), .B2(n9235), .A(n9194), .ZN(n9373) );
  NOR2_X1 U10219 ( .A1(n9374), .A2(n9373), .ZN(n9372) );
  AND2_X2 U10220 ( .A1(n9196), .A2(n9195), .ZN(n9377) );
  AOI22_X1 U10221 ( .A1(n9987), .A2(n9235), .B1(n9239), .B2(n9853), .ZN(n9275)
         );
  NAND2_X1 U10222 ( .A1(n9667), .A2(n9198), .ZN(n9199) );
  NAND2_X1 U10223 ( .A1(n9200), .A2(n9199), .ZN(n9201) );
  XNOR2_X1 U10224 ( .A(n9201), .B(n9243), .ZN(n9205) );
  NAND2_X1 U10225 ( .A1(n9981), .A2(n9235), .ZN(n9203) );
  NAND2_X1 U10226 ( .A1(n9667), .A2(n9239), .ZN(n9202) );
  NAND2_X1 U10227 ( .A1(n9203), .A2(n9202), .ZN(n9204) );
  NOR2_X1 U10228 ( .A1(n9205), .A2(n9204), .ZN(n9351) );
  NAND2_X1 U10229 ( .A1(n9205), .A2(n9204), .ZN(n9352) );
  NAND2_X1 U10230 ( .A1(n9666), .A2(n9235), .ZN(n9206) );
  NAND2_X1 U10231 ( .A1(n9207), .A2(n9206), .ZN(n9209) );
  XNOR2_X1 U10232 ( .A(n9209), .B(n9208), .ZN(n9212) );
  NOR2_X1 U10233 ( .A1(n9820), .A2(n9286), .ZN(n9210) );
  AOI21_X1 U10234 ( .B1(n9978), .B2(n9235), .A(n9210), .ZN(n9211) );
  NOR2_X1 U10235 ( .A1(n9212), .A2(n9211), .ZN(n9301) );
  NAND2_X1 U10236 ( .A1(n9212), .A2(n9211), .ZN(n9299) );
  NAND2_X1 U10237 ( .A1(n9775), .A2(n9235), .ZN(n9213) );
  NAND2_X1 U10238 ( .A1(n9214), .A2(n9213), .ZN(n9215) );
  XNOR2_X1 U10239 ( .A(n9215), .B(n9243), .ZN(n9218) );
  NAND2_X1 U10240 ( .A1(n9971), .A2(n9235), .ZN(n9217) );
  NAND2_X1 U10241 ( .A1(n9775), .A2(n9239), .ZN(n9216) );
  NAND2_X1 U10242 ( .A1(n9217), .A2(n9216), .ZN(n9219) );
  NAND2_X1 U10243 ( .A1(n9218), .A2(n9219), .ZN(n9363) );
  INV_X1 U10244 ( .A(n9218), .ZN(n9221) );
  INV_X1 U10245 ( .A(n9219), .ZN(n9220) );
  NAND2_X1 U10246 ( .A1(n9221), .A2(n9220), .ZN(n9365) );
  OAI22_X1 U10247 ( .A1(n9771), .A2(n9289), .B1(n9752), .B2(n9287), .ZN(n9222)
         );
  XOR2_X1 U10248 ( .A(n9243), .B(n9222), .Z(n9223) );
  NAND2_X1 U10249 ( .A1(n9224), .A2(n9223), .ZN(n9265) );
  OAI22_X1 U10250 ( .A1(n9771), .A2(n9287), .B1(n9752), .B2(n9286), .ZN(n9268)
         );
  XNOR2_X1 U10251 ( .A(n9226), .B(n9225), .ZN(n9342) );
  OR2_X1 U10252 ( .A1(n9754), .A2(n9287), .ZN(n9228) );
  NAND2_X1 U10253 ( .A1(n9229), .A2(n9228), .ZN(n9230) );
  XNOR2_X1 U10254 ( .A(n9230), .B(n9243), .ZN(n9311) );
  NAND2_X1 U10255 ( .A1(n9958), .A2(n9235), .ZN(n9232) );
  OR2_X1 U10256 ( .A1(n9754), .A2(n9286), .ZN(n9231) );
  NAND2_X1 U10257 ( .A1(n9232), .A2(n9231), .ZN(n9310) );
  INV_X1 U10258 ( .A(n9311), .ZN(n9234) );
  INV_X1 U10259 ( .A(n9310), .ZN(n9233) );
  NAND2_X1 U10260 ( .A1(n9664), .A2(n9235), .ZN(n9236) );
  NAND2_X1 U10261 ( .A1(n9237), .A2(n9236), .ZN(n9238) );
  XNOR2_X1 U10262 ( .A(n9238), .B(n9243), .ZN(n9241) );
  AOI22_X1 U10263 ( .A1(n9951), .A2(n9235), .B1(n9239), .B2(n9664), .ZN(n9240)
         );
  XNOR2_X1 U10264 ( .A(n9241), .B(n9240), .ZN(n9385) );
  INV_X1 U10265 ( .A(n9240), .ZN(n9242) );
  AOI22_X1 U10266 ( .A1(n9386), .A2(n9385), .B1(n9242), .B2(n9241), .ZN(n9248)
         );
  OAI22_X1 U10267 ( .A1(n9717), .A2(n9289), .B1(n9723), .B2(n9287), .ZN(n9244)
         );
  XNOR2_X1 U10268 ( .A(n9244), .B(n9243), .ZN(n9246) );
  OAI22_X1 U10269 ( .A1(n9717), .A2(n9287), .B1(n9723), .B2(n9286), .ZN(n9245)
         );
  NOR2_X1 U10270 ( .A1(n9246), .A2(n9245), .ZN(n9283) );
  AOI21_X1 U10271 ( .B1(n9246), .B2(n9245), .A(n9283), .ZN(n9247) );
  OAI21_X1 U10272 ( .B1(n9248), .B2(n9247), .A(n9285), .ZN(n9249) );
  NAND2_X1 U10273 ( .A1(n9249), .A2(n9376), .ZN(n9253) );
  AOI22_X1 U10274 ( .A1(n9381), .A2(n9664), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n9252) );
  INV_X1 U10275 ( .A(n9712), .ZN(n9689) );
  AOI22_X1 U10276 ( .A1(n9406), .A2(n9689), .B1(n9347), .B2(n9715), .ZN(n9251)
         );
  NAND2_X1 U10277 ( .A1(n9948), .A2(n9407), .ZN(n9250) );
  NAND4_X1 U10278 ( .A1(n9253), .A2(n9252), .A3(n9251), .A4(n9250), .ZN(
        P1_U3212) );
  NAND2_X1 U10279 ( .A1(n9255), .A2(n9254), .ZN(n9257) );
  XNOR2_X1 U10280 ( .A(n9257), .B(n9256), .ZN(n9258) );
  NAND2_X1 U10281 ( .A1(n9258), .A2(n9376), .ZN(n9264) );
  INV_X1 U10282 ( .A(n9919), .ZN(n9259) );
  OAI22_X1 U10283 ( .A1(n9260), .A2(n9402), .B1(n9401), .B2(n9259), .ZN(n9261)
         );
  AOI211_X1 U10284 ( .C1(n9406), .C2(n9911), .A(n9262), .B(n9261), .ZN(n9263)
         );
  OAI211_X1 U10285 ( .C1(n10853), .C2(n9384), .A(n9264), .B(n9263), .ZN(
        P1_U3213) );
  INV_X1 U10286 ( .A(n9265), .ZN(n9266) );
  NOR2_X1 U10287 ( .A1(n9267), .A2(n9266), .ZN(n9269) );
  XNOR2_X1 U10288 ( .A(n9269), .B(n9268), .ZN(n9274) );
  INV_X1 U10289 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9270) );
  OAI22_X1 U10290 ( .A1(n9808), .A2(n9402), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9270), .ZN(n9272) );
  OAI22_X1 U10291 ( .A1(n9741), .A2(n9388), .B1(n9768), .B2(n9401), .ZN(n9271)
         );
  AOI211_X1 U10292 ( .C1(n9966), .C2(n9407), .A(n9272), .B(n9271), .ZN(n9273)
         );
  OAI21_X1 U10293 ( .B1(n9274), .B2(n9410), .A(n9273), .ZN(P1_U3214) );
  XNOR2_X1 U10294 ( .A(n9276), .B(n9275), .ZN(n9277) );
  XNOR2_X1 U10295 ( .A(n5125), .B(n9277), .ZN(n9282) );
  OAI21_X1 U10296 ( .B1(n9402), .B2(n9837), .A(n9278), .ZN(n9280) );
  OAI22_X1 U10297 ( .A1(n9838), .A2(n9388), .B1(n9401), .B2(n9842), .ZN(n9279)
         );
  AOI211_X1 U10298 ( .C1(n9987), .C2(n9407), .A(n9280), .B(n9279), .ZN(n9281)
         );
  OAI21_X1 U10299 ( .B1(n9282), .B2(n9410), .A(n9281), .ZN(P1_U3217) );
  INV_X1 U10300 ( .A(n9283), .ZN(n9284) );
  OAI22_X1 U10301 ( .A1(n9701), .A2(n9287), .B1(n9712), .B2(n9286), .ZN(n9288)
         );
  XNOR2_X1 U10302 ( .A(n9288), .B(n9243), .ZN(n9291) );
  OAI22_X1 U10303 ( .A1(n9701), .A2(n9289), .B1(n9712), .B2(n9287), .ZN(n9290)
         );
  XNOR2_X1 U10304 ( .A(n9291), .B(n9290), .ZN(n9292) );
  OAI22_X1 U10305 ( .A1(n9402), .A2(n9723), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9293), .ZN(n9297) );
  INV_X1 U10306 ( .A(n9294), .ZN(n9295) );
  OAI22_X1 U10307 ( .A1(n9484), .A2(n9388), .B1(n9401), .B2(n9295), .ZN(n9296)
         );
  AOI211_X1 U10308 ( .C1(n9941), .C2(n9407), .A(n9297), .B(n9296), .ZN(n9298)
         );
  INV_X1 U10309 ( .A(n9299), .ZN(n9300) );
  NOR2_X1 U10310 ( .A1(n9301), .A2(n9300), .ZN(n9302) );
  XNOR2_X1 U10311 ( .A(n9303), .B(n9302), .ZN(n9309) );
  OAI22_X1 U10312 ( .A1(n9838), .A2(n9402), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9304), .ZN(n9307) );
  INV_X1 U10313 ( .A(n9305), .ZN(n9814) );
  OAI22_X1 U10314 ( .A1(n9808), .A2(n9388), .B1(n9401), .B2(n9814), .ZN(n9306)
         );
  AOI211_X1 U10315 ( .C1(n9978), .C2(n9407), .A(n9307), .B(n9306), .ZN(n9308)
         );
  OAI21_X1 U10316 ( .B1(n9309), .B2(n9410), .A(n9308), .ZN(P1_U3221) );
  XNOR2_X1 U10317 ( .A(n9311), .B(n9310), .ZN(n9312) );
  XNOR2_X1 U10318 ( .A(n9313), .B(n9312), .ZN(n9319) );
  OAI22_X1 U10319 ( .A1(n9388), .A2(n9742), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9314), .ZN(n9317) );
  INV_X1 U10320 ( .A(n9315), .ZN(n9744) );
  OAI22_X1 U10321 ( .A1(n9741), .A2(n9402), .B1(n9744), .B2(n9401), .ZN(n9316)
         );
  AOI211_X1 U10322 ( .C1(n9958), .C2(n9407), .A(n9317), .B(n9316), .ZN(n9318)
         );
  OAI21_X1 U10323 ( .B1(n9319), .B2(n9410), .A(n9318), .ZN(P1_U3223) );
  INV_X1 U10324 ( .A(n9321), .ZN(n9322) );
  NOR2_X1 U10325 ( .A1(n9320), .A2(n9322), .ZN(n9394) );
  NAND2_X1 U10326 ( .A1(n9320), .A2(n9322), .ZN(n9395) );
  OAI21_X1 U10327 ( .B1(n9394), .B2(n9397), .A(n9395), .ZN(n9326) );
  XNOR2_X1 U10328 ( .A(n9324), .B(n9323), .ZN(n9325) );
  XNOR2_X1 U10329 ( .A(n9326), .B(n9325), .ZN(n9331) );
  AOI22_X1 U10330 ( .A1(n9381), .A2(n9911), .B1(n9347), .B2(n9896), .ZN(n9328)
         );
  OAI211_X1 U10331 ( .C1(n9890), .C2(n9388), .A(n9328), .B(n9327), .ZN(n9329)
         );
  AOI21_X1 U10332 ( .B1(n10886), .B2(n9407), .A(n9329), .ZN(n9330) );
  OAI21_X1 U10333 ( .B1(n9331), .B2(n9410), .A(n9330), .ZN(P1_U3224) );
  XOR2_X1 U10334 ( .A(n9333), .B(n9332), .Z(n9339) );
  AOI22_X1 U10335 ( .A1(n9406), .A2(n9878), .B1(n9347), .B2(n9872), .ZN(n9335)
         );
  OAI211_X1 U10336 ( .C1(n9336), .C2(n9402), .A(n9335), .B(n9334), .ZN(n9337)
         );
  AOI21_X1 U10337 ( .B1(n9998), .B2(n9407), .A(n9337), .ZN(n9338) );
  OAI21_X1 U10338 ( .B1(n9339), .B2(n9410), .A(n9338), .ZN(P1_U3226) );
  OAI21_X1 U10339 ( .B1(n9342), .B2(n9341), .A(n9340), .ZN(n9343) );
  NAND2_X1 U10340 ( .A1(n9343), .A2(n9376), .ZN(n9349) );
  INV_X1 U10341 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9344) );
  OAI22_X1 U10342 ( .A1(n9388), .A2(n9754), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9344), .ZN(n9346) );
  NOR2_X1 U10343 ( .A1(n9752), .A2(n9402), .ZN(n9345) );
  AOI211_X1 U10344 ( .C1(n9347), .C2(n9758), .A(n9346), .B(n9345), .ZN(n9348)
         );
  OAI211_X1 U10345 ( .C1(n9350), .C2(n9384), .A(n9349), .B(n9348), .ZN(
        P1_U3227) );
  INV_X1 U10346 ( .A(n9351), .ZN(n9353) );
  NAND2_X1 U10347 ( .A1(n9353), .A2(n9352), .ZN(n9354) );
  XNOR2_X1 U10348 ( .A(n9355), .B(n9354), .ZN(n9360) );
  OAI22_X1 U10349 ( .A1(n9402), .A2(n9819), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9356), .ZN(n9358) );
  OAI22_X1 U10350 ( .A1(n9820), .A2(n9388), .B1(n9401), .B2(n9826), .ZN(n9357)
         );
  AOI211_X1 U10351 ( .C1(n9981), .C2(n9407), .A(n9358), .B(n9357), .ZN(n9359)
         );
  OAI21_X1 U10352 ( .B1(n9360), .B2(n9410), .A(n9359), .ZN(P1_U3231) );
  INV_X1 U10353 ( .A(n9361), .ZN(n9366) );
  AOI21_X1 U10354 ( .B1(n9365), .B2(n9363), .A(n9362), .ZN(n9364) );
  AOI21_X1 U10355 ( .B1(n9366), .B2(n9365), .A(n9364), .ZN(n9371) );
  OAI22_X1 U10356 ( .A1(n9752), .A2(n9388), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9367), .ZN(n9369) );
  OAI22_X1 U10357 ( .A1(n9820), .A2(n9402), .B1(n9784), .B2(n9401), .ZN(n9368)
         );
  AOI211_X1 U10358 ( .C1(n9971), .C2(n9407), .A(n9369), .B(n9368), .ZN(n9370)
         );
  OAI21_X1 U10359 ( .B1(n9371), .B2(n9410), .A(n9370), .ZN(P1_U3233) );
  INV_X1 U10360 ( .A(n9372), .ZN(n9378) );
  OAI21_X1 U10361 ( .B1(n9374), .B2(n9377), .A(n9373), .ZN(n9375) );
  OAI211_X1 U10362 ( .C1(n9378), .C2(n9377), .A(n9376), .B(n9375), .ZN(n9383)
         );
  OAI22_X1 U10363 ( .A1(n9819), .A2(n9388), .B1(n9401), .B2(n9859), .ZN(n9379)
         );
  AOI211_X1 U10364 ( .C1(n9381), .C2(n9852), .A(n9380), .B(n9379), .ZN(n9382)
         );
  OAI211_X1 U10365 ( .C1(n9862), .C2(n9384), .A(n9383), .B(n9382), .ZN(
        P1_U3236) );
  XNOR2_X1 U10366 ( .A(n9386), .B(n9385), .ZN(n9393) );
  OAI22_X1 U10367 ( .A1(n9388), .A2(n9723), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9387), .ZN(n9391) );
  INV_X1 U10368 ( .A(n9730), .ZN(n9389) );
  OAI22_X1 U10369 ( .A1(n9754), .A2(n9402), .B1(n9401), .B2(n9389), .ZN(n9390)
         );
  AOI211_X1 U10370 ( .C1(n9951), .C2(n9407), .A(n9391), .B(n9390), .ZN(n9392)
         );
  OAI21_X1 U10371 ( .B1(n9393), .B2(n9410), .A(n9392), .ZN(P1_U3238) );
  INV_X1 U10372 ( .A(n9394), .ZN(n9396) );
  NAND2_X1 U10373 ( .A1(n9396), .A2(n9395), .ZN(n9398) );
  XNOR2_X1 U10374 ( .A(n9398), .B(n9397), .ZN(n9411) );
  INV_X1 U10375 ( .A(n9399), .ZN(n9405) );
  OAI22_X1 U10376 ( .A1(n9403), .A2(n9402), .B1(n9401), .B2(n9400), .ZN(n9404)
         );
  AOI211_X1 U10377 ( .C1(n9406), .C2(n9879), .A(n9405), .B(n9404), .ZN(n9409)
         );
  NAND2_X1 U10378 ( .A1(n10876), .A2(n9407), .ZN(n9408) );
  OAI211_X1 U10379 ( .C1(n9411), .C2(n9410), .A(n9409), .B(n9408), .ZN(
        P1_U3239) );
  NAND2_X1 U10380 ( .A1(n9412), .A2(n9427), .ZN(n9415) );
  OR2_X1 U10381 ( .A1(n6149), .A2(n9413), .ZN(n9414) );
  NAND2_X1 U10382 ( .A1(n6031), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n9418) );
  NAND2_X1 U10383 ( .A1(n6932), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9417) );
  NAND2_X1 U10384 ( .A1(n9423), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9416) );
  NAND3_X1 U10385 ( .A1(n9418), .A2(n9417), .A3(n9416), .ZN(n9691) );
  INV_X1 U10386 ( .A(n9691), .ZN(n9483) );
  OR2_X1 U10387 ( .A1(n9680), .A2(n9483), .ZN(n9591) );
  NAND2_X1 U10388 ( .A1(n9419), .A2(n9427), .ZN(n9422) );
  INV_X1 U10389 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9420) );
  OR2_X1 U10390 ( .A1(n6149), .A2(n9420), .ZN(n9421) );
  NAND2_X1 U10391 ( .A1(n6031), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n9426) );
  NAND2_X1 U10392 ( .A1(n6933), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9425) );
  NAND2_X1 U10393 ( .A1(n9423), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n9424) );
  AND3_X1 U10394 ( .A1(n9426), .A2(n9425), .A3(n9424), .ZN(n9489) );
  NAND2_X1 U10395 ( .A1(n9591), .A2(n9491), .ZN(n9650) );
  INV_X1 U10396 ( .A(n9650), .ZN(n9487) );
  NAND2_X1 U10397 ( .A1(n9428), .A2(n9427), .ZN(n9430) );
  OR2_X1 U10398 ( .A1(n6149), .A2(n10448), .ZN(n9429) );
  NAND2_X1 U10399 ( .A1(n9624), .A2(n9684), .ZN(n9618) );
  AND2_X1 U10400 ( .A1(n9496), .A2(n9498), .ZN(n9431) );
  NAND2_X1 U10401 ( .A1(n9495), .A2(n9431), .ZN(n9479) );
  INV_X1 U10402 ( .A(n9432), .ZN(n9433) );
  OR2_X1 U10403 ( .A1(n9574), .A2(n9433), .ZN(n9502) );
  NOR2_X1 U10404 ( .A1(n9479), .A2(n9502), .ZN(n9616) );
  OAI21_X1 U10405 ( .B1(n9473), .B2(n9434), .A(n9559), .ZN(n9435) );
  NOR2_X1 U10406 ( .A1(n9566), .A2(n9435), .ZN(n9436) );
  OR2_X1 U10407 ( .A1(n9792), .A2(n9436), .ZN(n9437) );
  NAND2_X1 U10408 ( .A1(n9437), .A2(n9791), .ZN(n9608) );
  AND2_X1 U10409 ( .A1(n9549), .A2(n9545), .ZN(n9438) );
  AND2_X1 U10410 ( .A1(n9554), .A2(n9438), .ZN(n9470) );
  INV_X1 U10411 ( .A(n9470), .ZN(n9442) );
  NAND2_X1 U10412 ( .A1(n9536), .A2(n9905), .ZN(n9535) );
  INV_X1 U10413 ( .A(n9515), .ZN(n9439) );
  OAI211_X1 U10414 ( .C1(n9439), .C2(n9504), .A(n9519), .B(n9516), .ZN(n9465)
         );
  INV_X1 U10415 ( .A(n9465), .ZN(n9440) );
  NAND4_X1 U10416 ( .A1(n9440), .A2(n9530), .A3(n9503), .A4(n9506), .ZN(n9441)
         );
  OR4_X1 U10417 ( .A1(n9442), .A2(n5381), .A3(n9535), .A4(n9441), .ZN(n9606)
         );
  OAI211_X1 U10418 ( .C1(n9445), .C2(n9444), .A(n9597), .B(n9443), .ZN(n9447)
         );
  NAND2_X1 U10419 ( .A1(n9447), .A2(n9446), .ZN(n9449) );
  OAI21_X1 U10420 ( .B1(n9450), .B2(n9449), .A(n9448), .ZN(n9452) );
  NAND2_X1 U10421 ( .A1(n9452), .A2(n9451), .ZN(n9455) );
  NAND3_X1 U10422 ( .A1(n9455), .A2(n9454), .A3(n9453), .ZN(n9458) );
  NAND3_X1 U10423 ( .A1(n9458), .A2(n9457), .A3(n9456), .ZN(n9461) );
  NAND2_X1 U10424 ( .A1(n9507), .A2(n5386), .ZN(n9460) );
  AND4_X1 U10425 ( .A1(n9461), .A2(n9510), .A3(n9460), .A4(n9505), .ZN(n9472)
         );
  NAND2_X1 U10426 ( .A1(n9534), .A2(n9528), .ZN(n9537) );
  INV_X1 U10427 ( .A(n9513), .ZN(n9463) );
  AND3_X1 U10428 ( .A1(n9463), .A2(n9515), .A3(n9462), .ZN(n9464) );
  OAI211_X1 U10429 ( .C1(n9465), .C2(n9464), .A(n9526), .B(n9524), .ZN(n9466)
         );
  AND3_X1 U10430 ( .A1(n9905), .A2(n9466), .A3(n9530), .ZN(n9467) );
  OAI211_X1 U10431 ( .C1(n9537), .C2(n9467), .A(n9542), .B(n9536), .ZN(n9468)
         );
  NAND3_X1 U10432 ( .A1(n9544), .A2(n9468), .A3(n9541), .ZN(n9469) );
  AND2_X1 U10433 ( .A1(n9470), .A2(n9469), .ZN(n9609) );
  INV_X1 U10434 ( .A(n9609), .ZN(n9471) );
  OAI21_X1 U10435 ( .B1(n9606), .B2(n9472), .A(n9471), .ZN(n9477) );
  NOR2_X1 U10436 ( .A1(n9792), .A2(n9473), .ZN(n9474) );
  OR2_X1 U10437 ( .A1(n9608), .A2(n9474), .ZN(n9475) );
  NAND2_X1 U10438 ( .A1(n9966), .A2(n9752), .ZN(n9500) );
  NAND2_X1 U10439 ( .A1(n9475), .A2(n9500), .ZN(n9612) );
  INV_X1 U10440 ( .A(n9612), .ZN(n9476) );
  OAI21_X1 U10441 ( .B1(n9608), .B2(n9477), .A(n9476), .ZN(n9482) );
  NAND2_X1 U10442 ( .A1(n9963), .A2(n9741), .ZN(n9573) );
  AND2_X1 U10443 ( .A1(n9499), .A2(n9573), .ZN(n9478) );
  OR2_X1 U10444 ( .A1(n9479), .A2(n9478), .ZN(n9481) );
  INV_X1 U10445 ( .A(n9497), .ZN(n9709) );
  NAND2_X1 U10446 ( .A1(n9495), .A2(n9709), .ZN(n9480) );
  NAND4_X1 U10447 ( .A1(n9481), .A2(n9480), .A3(n9586), .A4(n9583), .ZN(n9614)
         );
  AOI21_X1 U10448 ( .B1(n9616), .B2(n9482), .A(n9614), .ZN(n9485) );
  NAND2_X1 U10449 ( .A1(n9680), .A2(n9483), .ZN(n9646) );
  OAI211_X1 U10450 ( .C1(n9618), .C2(n9485), .A(n9646), .B(n9623), .ZN(n9486)
         );
  INV_X1 U10451 ( .A(n9489), .ZN(n9677) );
  AOI21_X1 U10452 ( .B1(n9487), .B2(n9486), .A(n9651), .ZN(n9488) );
  XNOR2_X1 U10453 ( .A(n9488), .B(n9812), .ZN(n9658) );
  OR2_X1 U10454 ( .A1(n9591), .A2(n9489), .ZN(n9490) );
  NAND2_X1 U10455 ( .A1(n9491), .A2(n9490), .ZN(n9605) );
  NAND2_X1 U10456 ( .A1(n9646), .A2(n9677), .ZN(n9492) );
  NAND2_X1 U10457 ( .A1(n9492), .A2(n9680), .ZN(n9617) );
  NOR2_X1 U10458 ( .A1(n9493), .A2(n9617), .ZN(n9494) );
  INV_X1 U10459 ( .A(n9495), .ZN(n9584) );
  MUX2_X1 U10460 ( .A(n9497), .B(n9496), .S(n9590), .Z(n9581) );
  INV_X1 U10461 ( .A(n9726), .ZN(n9580) );
  INV_X1 U10462 ( .A(n9590), .ZN(n9558) );
  MUX2_X1 U10463 ( .A(n9499), .B(n9498), .S(n9558), .Z(n9579) );
  NAND2_X1 U10464 ( .A1(n9573), .A2(n9500), .ZN(n9501) );
  MUX2_X1 U10465 ( .A(n9502), .B(n9501), .S(n9590), .Z(n9578) );
  INV_X1 U10466 ( .A(n9505), .ZN(n9508) );
  OAI211_X1 U10467 ( .C1(n9509), .C2(n9508), .A(n9507), .B(n9506), .ZN(n9512)
         );
  NAND2_X1 U10468 ( .A1(n9514), .A2(n5067), .ZN(n9522) );
  MUX2_X1 U10469 ( .A(n9516), .B(n9515), .S(n9558), .Z(n9517) );
  INV_X1 U10470 ( .A(n9517), .ZN(n9518) );
  NOR2_X1 U10471 ( .A1(n10750), .A2(n9518), .ZN(n9521) );
  OAI21_X1 U10472 ( .B1(n9519), .B2(n9590), .A(n9636), .ZN(n9520) );
  AOI21_X1 U10473 ( .B1(n9522), .B2(n9521), .A(n9520), .ZN(n9527) );
  INV_X1 U10474 ( .A(n9527), .ZN(n9525) );
  AOI21_X1 U10475 ( .B1(n9525), .B2(n9524), .A(n9523), .ZN(n9533) );
  NAND2_X1 U10476 ( .A1(n9527), .A2(n9526), .ZN(n9531) );
  INV_X1 U10477 ( .A(n9528), .ZN(n9529) );
  AOI21_X1 U10478 ( .B1(n9531), .B2(n9530), .A(n9529), .ZN(n9532) );
  INV_X1 U10479 ( .A(n9915), .ZN(n9907) );
  NAND2_X1 U10480 ( .A1(n9535), .A2(n9534), .ZN(n9539) );
  NAND2_X1 U10481 ( .A1(n9537), .A2(n9536), .ZN(n9538) );
  MUX2_X1 U10482 ( .A(n9539), .B(n9538), .S(n9558), .Z(n9540) );
  INV_X1 U10483 ( .A(n9892), .ZN(n9641) );
  MUX2_X1 U10484 ( .A(n9542), .B(n9541), .S(n9590), .Z(n9543) );
  MUX2_X1 U10485 ( .A(n9545), .B(n9544), .S(n9558), .Z(n9546) );
  NAND3_X1 U10486 ( .A1(n9547), .A2(n9876), .A3(n9546), .ZN(n9551) );
  MUX2_X1 U10487 ( .A(n9549), .B(n9548), .S(n9590), .Z(n9550) );
  NAND2_X1 U10488 ( .A1(n9551), .A2(n9550), .ZN(n9552) );
  NAND2_X1 U10489 ( .A1(n9552), .A2(n9855), .ZN(n9557) );
  INV_X1 U10490 ( .A(n9835), .ZN(n9556) );
  MUX2_X1 U10491 ( .A(n9554), .B(n9553), .S(n9590), .Z(n9555) );
  NAND3_X1 U10492 ( .A1(n9557), .A2(n9556), .A3(n9555), .ZN(n9562) );
  MUX2_X1 U10493 ( .A(n9560), .B(n9559), .S(n9558), .Z(n9561) );
  NAND2_X1 U10494 ( .A1(n9562), .A2(n9561), .ZN(n9564) );
  NOR2_X1 U10495 ( .A1(n9806), .A2(n9821), .ZN(n9563) );
  NAND2_X1 U10496 ( .A1(n9564), .A2(n9563), .ZN(n9569) );
  NAND2_X1 U10497 ( .A1(n9566), .A2(n9565), .ZN(n9567) );
  MUX2_X1 U10498 ( .A(n9567), .B(n9789), .S(n9590), .Z(n9568) );
  NAND3_X1 U10499 ( .A1(n9569), .A2(n9788), .A3(n9568), .ZN(n9572) );
  MUX2_X1 U10500 ( .A(n9570), .B(n9791), .S(n9590), .Z(n9571) );
  INV_X1 U10501 ( .A(n9738), .ZN(n9736) );
  INV_X1 U10502 ( .A(n9573), .ZN(n9575) );
  MUX2_X1 U10503 ( .A(n9575), .B(n9574), .S(n9590), .Z(n9576) );
  INV_X1 U10504 ( .A(n9576), .ZN(n9577) );
  NAND2_X1 U10505 ( .A1(n9686), .A2(n9582), .ZN(n9588) );
  OAI211_X1 U10506 ( .C1(n9584), .C2(n9588), .A(n9623), .B(n9583), .ZN(n9585)
         );
  INV_X1 U10507 ( .A(n9586), .ZN(n9587) );
  NOR2_X1 U10508 ( .A1(n9588), .A2(n9587), .ZN(n9589) );
  NAND3_X1 U10509 ( .A1(n9591), .A2(n9646), .A3(n9677), .ZN(n9592) );
  OAI21_X1 U10510 ( .B1(n9593), .B2(n9680), .A(n9592), .ZN(n9594) );
  AOI21_X1 U10511 ( .B1(n9597), .B2(n9596), .A(n9600), .ZN(n9604) );
  NAND2_X1 U10512 ( .A1(n9598), .A2(n9760), .ZN(n9599) );
  INV_X1 U10513 ( .A(n9605), .ZN(n9621) );
  INV_X1 U10514 ( .A(n9606), .ZN(n9611) );
  AOI211_X1 U10515 ( .C1(n9611), .C2(n9610), .A(n9609), .B(n9608), .ZN(n9613)
         );
  OR2_X1 U10516 ( .A1(n9613), .A2(n9612), .ZN(n9615) );
  AOI21_X1 U10517 ( .B1(n9616), .B2(n9615), .A(n9614), .ZN(n9619) );
  OAI211_X1 U10518 ( .C1(n9619), .C2(n9618), .A(n9617), .B(n9623), .ZN(n9620)
         );
  NAND2_X1 U10519 ( .A1(n9621), .A2(n9620), .ZN(n9622) );
  AOI21_X1 U10520 ( .B1(n9622), .B2(n9601), .A(n9760), .ZN(n9655) );
  NAND2_X1 U10521 ( .A1(n9624), .A2(n9623), .ZN(n9703) );
  INV_X1 U10522 ( .A(n9703), .ZN(n9648) );
  INV_X1 U10523 ( .A(n10750), .ZN(n10751) );
  NOR4_X1 U10524 ( .A1(n9628), .A2(n9627), .A3(n9626), .A4(n9625), .ZN(n9630)
         );
  NAND4_X1 U10525 ( .A1(n9632), .A2(n9631), .A3(n9630), .A4(n9629), .ZN(n9633)
         );
  NOR4_X1 U10526 ( .A1(n5538), .A2(n10712), .A3(n9634), .A4(n9633), .ZN(n9635)
         );
  NAND4_X1 U10527 ( .A1(n9636), .A2(n5067), .A3(n10751), .A4(n9635), .ZN(n9637) );
  NOR4_X1 U10528 ( .A1(n9639), .A2(n9915), .A3(n9638), .A4(n9637), .ZN(n9640)
         );
  NAND4_X1 U10529 ( .A1(n9876), .A2(n9855), .A3(n9641), .A4(n9640), .ZN(n9642)
         );
  NOR4_X1 U10530 ( .A1(n9806), .A2(n9821), .A3(n9835), .A4(n9642), .ZN(n9643)
         );
  NAND4_X1 U10531 ( .A1(n9750), .A2(n9788), .A3(n9643), .A4(n9773), .ZN(n9644)
         );
  NOR4_X1 U10532 ( .A1(n9645), .A2(n9738), .A3(n9726), .A4(n9644), .ZN(n9647)
         );
  NAND4_X1 U10533 ( .A1(n9648), .A2(n9714), .A3(n9647), .A4(n9646), .ZN(n9649)
         );
  NOR3_X1 U10534 ( .A1(n9651), .A2(n9650), .A3(n9649), .ZN(n9652) );
  XNOR2_X1 U10535 ( .A(n9652), .B(n9812), .ZN(n9654) );
  MUX2_X1 U10536 ( .A(n9655), .B(n9654), .S(n9653), .Z(n9656) );
  NAND4_X1 U10537 ( .A1(n10020), .A2(n9912), .A3(n9659), .A4(n9676), .ZN(n9660) );
  OAI211_X1 U10538 ( .C1(n9661), .C2(n9663), .A(n9660), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9662) );
  MUX2_X1 U10539 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9677), .S(P1_U4006), .Z(
        P1_U3586) );
  MUX2_X1 U10540 ( .A(n9691), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9674), .Z(
        P1_U3585) );
  MUX2_X1 U10541 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9689), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10542 ( .A(n9664), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9674), .Z(
        P1_U3581) );
  MUX2_X1 U10543 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9665), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10544 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9776), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10545 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9799), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10546 ( .A(n9666), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9674), .Z(
        P1_U3576) );
  MUX2_X1 U10547 ( .A(n9667), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9674), .Z(
        P1_U3575) );
  MUX2_X1 U10548 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9853), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10549 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9852), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10550 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9879), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10551 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9911), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10552 ( .A(n9668), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9674), .Z(
        P1_U3567) );
  MUX2_X1 U10553 ( .A(n9669), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9674), .Z(
        P1_U3565) );
  MUX2_X1 U10554 ( .A(n9670), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9674), .Z(
        P1_U3564) );
  MUX2_X1 U10555 ( .A(n9671), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9674), .Z(
        P1_U3563) );
  MUX2_X1 U10556 ( .A(n9672), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9674), .Z(
        P1_U3561) );
  MUX2_X1 U10557 ( .A(n9673), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9674), .Z(
        P1_U3560) );
  MUX2_X1 U10558 ( .A(n6208), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9674), .Z(
        P1_U3556) );
  XNOR2_X1 U10559 ( .A(n9930), .B(n9675), .ZN(n9928) );
  NAND2_X1 U10560 ( .A1(n9928), .A2(n10772), .ZN(n9679) );
  AOI21_X1 U10561 ( .B1(n9676), .B2(P1_B_REG_SCAN_IN), .A(n10753), .ZN(n9690)
         );
  NAND2_X1 U10562 ( .A1(n9677), .A2(n9690), .ZN(n9932) );
  NOR2_X1 U10563 ( .A1(n10778), .A2(n9932), .ZN(n9681) );
  AOI21_X1 U10564 ( .B1(n10778), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9681), .ZN(
        n9678) );
  OAI211_X1 U10565 ( .C1(n9930), .C2(n10780), .A(n9679), .B(n9678), .ZN(
        P1_U3261) );
  XNOR2_X1 U10566 ( .A(n9696), .B(n9680), .ZN(n9931) );
  NAND2_X1 U10567 ( .A1(n9931), .A2(n10772), .ZN(n9683) );
  AOI21_X1 U10568 ( .B1(n10778), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9681), .ZN(
        n9682) );
  OAI211_X1 U10569 ( .C1(n9934), .C2(n10780), .A(n9683), .B(n9682), .ZN(
        P1_U3262) );
  INV_X1 U10570 ( .A(n9684), .ZN(n9685) );
  AOI21_X1 U10571 ( .B1(n9687), .B2(n9686), .A(n9685), .ZN(n9688) );
  NAND2_X1 U10572 ( .A1(n9689), .A2(n9912), .ZN(n9693) );
  NAND2_X1 U10573 ( .A1(n9691), .A2(n9690), .ZN(n9692) );
  AOI21_X1 U10574 ( .B1(n9936), .B2(n9697), .A(n9696), .ZN(n9937) );
  INV_X1 U10575 ( .A(n9936), .ZN(n9700) );
  AOI22_X1 U10576 ( .A1(n10778), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9698), 
        .B2(n10776), .ZN(n9699) );
  OAI21_X1 U10577 ( .B1(n9700), .B2(n10780), .A(n9699), .ZN(n9705) );
  INV_X1 U10578 ( .A(n9729), .ZN(n9708) );
  INV_X1 U10579 ( .A(n9706), .ZN(n9707) );
  AOI211_X1 U10580 ( .C1(n9948), .C2(n9708), .A(n10833), .B(n9707), .ZN(n9947)
         );
  AOI21_X1 U10581 ( .B1(n9947), .B2(n9812), .A(n9946), .ZN(n9721) );
  INV_X1 U10582 ( .A(n9949), .ZN(n9719) );
  AOI22_X1 U10583 ( .A1(n10778), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n10776), 
        .B2(n9715), .ZN(n9716) );
  OAI21_X1 U10584 ( .B1(n9717), .B2(n10780), .A(n9716), .ZN(n9718) );
  AOI21_X1 U10585 ( .B1(n9719), .B2(n9926), .A(n9718), .ZN(n9720) );
  OAI21_X1 U10586 ( .B1(n9721), .B2(n10778), .A(n9720), .ZN(P1_U3264) );
  XNOR2_X1 U10587 ( .A(n9722), .B(n9726), .ZN(n9950) );
  OAI22_X1 U10588 ( .A1(n9723), .A2(n10753), .B1(n9754), .B2(n10755), .ZN(
        n9728) );
  AOI21_X1 U10589 ( .B1(n9726), .B2(n9725), .A(n9724), .ZN(n9727) );
  INV_X1 U10590 ( .A(n9951), .ZN(n9733) );
  AOI21_X1 U10591 ( .B1(n9951), .B2(n9743), .A(n9729), .ZN(n9952) );
  NAND2_X1 U10592 ( .A1(n9952), .A2(n10772), .ZN(n9732) );
  AOI22_X1 U10593 ( .A1(n10778), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9730), 
        .B2(n10776), .ZN(n9731) );
  OAI211_X1 U10594 ( .C1(n9733), .C2(n10780), .A(n9732), .B(n9731), .ZN(n9734)
         );
  AOI21_X1 U10595 ( .B1(n9950), .B2(n10773), .A(n9734), .ZN(n9735) );
  OAI21_X1 U10596 ( .B1(n9954), .B2(n10778), .A(n9735), .ZN(P1_U3265) );
  XNOR2_X1 U10597 ( .A(n9737), .B(n9736), .ZN(n9960) );
  XNOR2_X1 U10598 ( .A(n9739), .B(n9738), .ZN(n9740) );
  OAI222_X1 U10599 ( .A1(n10753), .A2(n9742), .B1(n10755), .B2(n9741), .C1(
        n9888), .C2(n9740), .ZN(n9956) );
  AOI211_X1 U10600 ( .C1(n9958), .C2(n9755), .A(n10833), .B(n8467), .ZN(n9957)
         );
  INV_X1 U10601 ( .A(n9957), .ZN(n9745) );
  OAI22_X1 U10602 ( .A1(n9745), .A2(n9760), .B1(n9897), .B2(n9744), .ZN(n9746)
         );
  OAI21_X1 U10603 ( .B1(n9956), .B2(n9746), .A(n10783), .ZN(n9748) );
  AOI22_X1 U10604 ( .A1(n9958), .A2(n9920), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n10778), .ZN(n9747) );
  OAI211_X1 U10605 ( .C1(n9885), .C2(n9960), .A(n9748), .B(n9747), .ZN(
        P1_U3266) );
  XOR2_X1 U10606 ( .A(n9750), .B(n9749), .Z(n9965) );
  XNOR2_X1 U10607 ( .A(n9751), .B(n9750), .ZN(n9753) );
  OAI222_X1 U10608 ( .A1(n10753), .A2(n9754), .B1(n9753), .B2(n9888), .C1(
        n10755), .C2(n9752), .ZN(n9961) );
  INV_X1 U10609 ( .A(n9766), .ZN(n9757) );
  INV_X1 U10610 ( .A(n9755), .ZN(n9756) );
  AOI211_X1 U10611 ( .C1(n9963), .C2(n9757), .A(n10833), .B(n9756), .ZN(n9962)
         );
  INV_X1 U10612 ( .A(n9962), .ZN(n9761) );
  INV_X1 U10613 ( .A(n9758), .ZN(n9759) );
  OAI22_X1 U10614 ( .A1(n9761), .A2(n9760), .B1(n9897), .B2(n9759), .ZN(n9762)
         );
  OAI21_X1 U10615 ( .B1(n9961), .B2(n9762), .A(n10783), .ZN(n9764) );
  AOI22_X1 U10616 ( .A1(n9963), .A2(n9920), .B1(n10778), .B2(
        P1_REG2_REG_24__SCAN_IN), .ZN(n9763) );
  OAI211_X1 U10617 ( .C1(n9885), .C2(n9965), .A(n9764), .B(n9763), .ZN(
        P1_U3267) );
  XNOR2_X1 U10618 ( .A(n9765), .B(n9773), .ZN(n9970) );
  INV_X1 U10619 ( .A(n9783), .ZN(n9767) );
  AOI21_X1 U10620 ( .B1(n9966), .B2(n9767), .A(n9766), .ZN(n9967) );
  INV_X1 U10621 ( .A(n9768), .ZN(n9769) );
  AOI22_X1 U10622 ( .A1(n9769), .A2(n10776), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n10778), .ZN(n9770) );
  OAI21_X1 U10623 ( .B1(n9771), .B2(n10780), .A(n9770), .ZN(n9780) );
  OAI211_X1 U10624 ( .C1(n9774), .C2(n9773), .A(n9772), .B(n10758), .ZN(n9778)
         );
  AOI22_X1 U10625 ( .A1(n9776), .A2(n9910), .B1(n9912), .B2(n9775), .ZN(n9777)
         );
  AND2_X1 U10626 ( .A1(n9778), .A2(n9777), .ZN(n9969) );
  NOR2_X1 U10627 ( .A1(n9969), .A2(n10778), .ZN(n9779) );
  AOI211_X1 U10628 ( .C1(n9967), .C2(n10772), .A(n9780), .B(n9779), .ZN(n9781)
         );
  OAI21_X1 U10629 ( .B1(n9885), .B2(n9970), .A(n9781), .ZN(P1_U3268) );
  XOR2_X1 U10630 ( .A(n9782), .B(n9788), .Z(n9975) );
  AOI21_X1 U10631 ( .B1(n9971), .B2(n9810), .A(n9783), .ZN(n9972) );
  INV_X1 U10632 ( .A(n9971), .ZN(n9787) );
  INV_X1 U10633 ( .A(n9784), .ZN(n9785) );
  AOI22_X1 U10634 ( .A1(n9785), .A2(n10776), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n10778), .ZN(n9786) );
  OAI21_X1 U10635 ( .B1(n9787), .B2(n10780), .A(n9786), .ZN(n9801) );
  NOR2_X1 U10636 ( .A1(n9820), .A2(n10755), .ZN(n9798) );
  INV_X1 U10637 ( .A(n9794), .ZN(n9790) );
  AOI21_X1 U10638 ( .B1(n9790), .B2(n9789), .A(n9788), .ZN(n9796) );
  INV_X1 U10639 ( .A(n9791), .ZN(n9793) );
  NOR3_X1 U10640 ( .A1(n9794), .A2(n9793), .A3(n9792), .ZN(n9795) );
  NOR3_X1 U10641 ( .A1(n9796), .A2(n9795), .A3(n9888), .ZN(n9797) );
  AOI211_X1 U10642 ( .C1(n9910), .C2(n9799), .A(n9798), .B(n9797), .ZN(n9974)
         );
  NOR2_X1 U10643 ( .A1(n9974), .A2(n10778), .ZN(n9800) );
  AOI211_X1 U10644 ( .C1(n9972), .C2(n10772), .A(n9801), .B(n9800), .ZN(n9802)
         );
  OAI21_X1 U10645 ( .B1(n9885), .B2(n9975), .A(n9802), .ZN(P1_U3269) );
  XNOR2_X1 U10646 ( .A(n9803), .B(n9806), .ZN(n9980) );
  OAI21_X1 U10647 ( .B1(n5365), .B2(n9821), .A(n9804), .ZN(n9805) );
  XOR2_X1 U10648 ( .A(n9806), .B(n9805), .Z(n9807) );
  OAI222_X1 U10649 ( .A1(n10753), .A2(n9808), .B1(n10755), .B2(n9838), .C1(
        n9888), .C2(n9807), .ZN(n9976) );
  AOI21_X1 U10650 ( .B1(n9978), .B2(n5349), .A(n10833), .ZN(n9811) );
  AND2_X1 U10651 ( .A1(n9811), .A2(n9810), .ZN(n9977) );
  NAND2_X1 U10652 ( .A1(n9977), .A2(n9812), .ZN(n9813) );
  OAI21_X1 U10653 ( .B1(n9897), .B2(n9814), .A(n9813), .ZN(n9815) );
  OAI21_X1 U10654 ( .B1(n9976), .B2(n9815), .A(n10783), .ZN(n9817) );
  AOI22_X1 U10655 ( .A1(n9978), .A2(n9920), .B1(n10778), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9816) );
  OAI211_X1 U10656 ( .C1(n9885), .C2(n9980), .A(n9817), .B(n9816), .ZN(
        P1_U3270) );
  XNOR2_X1 U10657 ( .A(n9818), .B(n9821), .ZN(n9825) );
  OAI22_X1 U10658 ( .A1(n9820), .A2(n10753), .B1(n9819), .B2(n10755), .ZN(
        n9824) );
  XNOR2_X1 U10659 ( .A(n9822), .B(n9821), .ZN(n9985) );
  NOR2_X1 U10660 ( .A1(n9985), .A2(n10718), .ZN(n9823) );
  AOI211_X1 U10661 ( .C1(n10758), .C2(n9825), .A(n9824), .B(n9823), .ZN(n9984)
         );
  AOI21_X1 U10662 ( .B1(n9981), .B2(n9839), .A(n9809), .ZN(n9982) );
  INV_X1 U10663 ( .A(n9826), .ZN(n9827) );
  AOI22_X1 U10664 ( .A1(n10778), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9827), 
        .B2(n10776), .ZN(n9828) );
  OAI21_X1 U10665 ( .B1(n5347), .B2(n10780), .A(n9828), .ZN(n9830) );
  NOR2_X1 U10666 ( .A1(n9985), .A2(n9867), .ZN(n9829) );
  AOI211_X1 U10667 ( .C1(n9982), .C2(n10772), .A(n9830), .B(n9829), .ZN(n9831)
         );
  OAI21_X1 U10668 ( .B1(n9984), .B2(n10778), .A(n9831), .ZN(P1_U3271) );
  XNOR2_X1 U10669 ( .A(n9832), .B(n9835), .ZN(n9991) );
  AOI21_X1 U10670 ( .B1(n9835), .B2(n9834), .A(n9833), .ZN(n9836) );
  OAI222_X1 U10671 ( .A1(n10753), .A2(n9838), .B1(n10755), .B2(n9837), .C1(
        n9888), .C2(n9836), .ZN(n9986) );
  INV_X1 U10672 ( .A(n9863), .ZN(n9841) );
  INV_X1 U10673 ( .A(n9839), .ZN(n9840) );
  AOI21_X1 U10674 ( .B1(n9987), .B2(n9841), .A(n9840), .ZN(n9988) );
  NAND2_X1 U10675 ( .A1(n9988), .A2(n10772), .ZN(n9845) );
  INV_X1 U10676 ( .A(n9842), .ZN(n9843) );
  AOI22_X1 U10677 ( .A1(n10778), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9843), 
        .B2(n10776), .ZN(n9844) );
  OAI211_X1 U10678 ( .C1(n9846), .C2(n10780), .A(n9845), .B(n9844), .ZN(n9847)
         );
  AOI21_X1 U10679 ( .B1(n9986), .B2(n10783), .A(n9847), .ZN(n9848) );
  OAI21_X1 U10680 ( .B1(n9885), .B2(n9991), .A(n9848), .ZN(P1_U3272) );
  NAND2_X1 U10681 ( .A1(n9849), .A2(n9855), .ZN(n9850) );
  NAND2_X1 U10682 ( .A1(n9851), .A2(n9850), .ZN(n9997) );
  AOI22_X1 U10683 ( .A1(n9853), .A2(n9910), .B1(n9852), .B2(n9912), .ZN(n9858)
         );
  OAI211_X1 U10684 ( .C1(n9856), .C2(n9855), .A(n9854), .B(n10758), .ZN(n9857)
         );
  OAI211_X1 U10685 ( .C1(n9997), .C2(n10718), .A(n9858), .B(n9857), .ZN(n9992)
         );
  INV_X1 U10686 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9860) );
  OAI22_X1 U10687 ( .A1(n10783), .A2(n9860), .B1(n9859), .B2(n9897), .ZN(n9861) );
  AOI21_X1 U10688 ( .B1(n9993), .B2(n9920), .A(n9861), .ZN(n9866) );
  NOR2_X1 U10689 ( .A1(n9862), .A2(n9871), .ZN(n9864) );
  NOR2_X1 U10690 ( .A1(n9864), .A2(n9863), .ZN(n9994) );
  NAND2_X1 U10691 ( .A1(n9994), .A2(n10772), .ZN(n9865) );
  OAI211_X1 U10692 ( .C1(n9997), .C2(n9867), .A(n9866), .B(n9865), .ZN(n9868)
         );
  AOI21_X1 U10693 ( .B1(n9992), .B2(n10783), .A(n9868), .ZN(n9869) );
  INV_X1 U10694 ( .A(n9869), .ZN(P1_U3273) );
  XOR2_X1 U10695 ( .A(n9870), .B(n9876), .Z(n10002) );
  AOI21_X1 U10696 ( .B1(n9998), .B2(n5075), .A(n9871), .ZN(n9999) );
  INV_X1 U10697 ( .A(n9998), .ZN(n9874) );
  AOI22_X1 U10698 ( .A1(n10778), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9872), 
        .B2(n10776), .ZN(n9873) );
  OAI21_X1 U10699 ( .B1(n9874), .B2(n10780), .A(n9873), .ZN(n9883) );
  OAI211_X1 U10700 ( .C1(n9877), .C2(n9876), .A(n9875), .B(n10758), .ZN(n9881)
         );
  AOI22_X1 U10701 ( .A1(n9912), .A2(n9879), .B1(n9878), .B2(n9910), .ZN(n9880)
         );
  AND2_X1 U10702 ( .A1(n9881), .A2(n9880), .ZN(n10001) );
  NOR2_X1 U10703 ( .A1(n10001), .A2(n10778), .ZN(n9882) );
  AOI211_X1 U10704 ( .C1(n9999), .C2(n10772), .A(n9883), .B(n9882), .ZN(n9884)
         );
  OAI21_X1 U10705 ( .B1(n9885), .B2(n10002), .A(n9884), .ZN(P1_U3274) );
  XNOR2_X1 U10706 ( .A(n9886), .B(n9892), .ZN(n9889) );
  OAI222_X1 U10707 ( .A1(n10753), .A2(n9890), .B1(n9889), .B2(n9888), .C1(
        n10755), .C2(n9887), .ZN(n10890) );
  INV_X1 U10708 ( .A(n10890), .ZN(n9904) );
  OAI21_X1 U10709 ( .B1(n9893), .B2(n9892), .A(n9891), .ZN(n9894) );
  INV_X1 U10710 ( .A(n9894), .ZN(n10893) );
  AOI21_X1 U10711 ( .B1(n10886), .B2(n5130), .A(n10833), .ZN(n9895) );
  NAND2_X1 U10712 ( .A1(n9895), .A2(n5075), .ZN(n10887) );
  INV_X1 U10713 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9899) );
  INV_X1 U10714 ( .A(n9896), .ZN(n9898) );
  OAI22_X1 U10715 ( .A1(n10783), .A2(n9899), .B1(n9898), .B2(n9897), .ZN(n9900) );
  AOI21_X1 U10716 ( .B1(n10886), .B2(n9920), .A(n9900), .ZN(n9901) );
  OAI21_X1 U10717 ( .B1(n10887), .B2(n9924), .A(n9901), .ZN(n9902) );
  AOI21_X1 U10718 ( .B1(n10893), .B2(n9926), .A(n9902), .ZN(n9903) );
  OAI21_X1 U10719 ( .B1(n9904), .B2(n10778), .A(n9903), .ZN(P1_U3275) );
  NAND2_X1 U10720 ( .A1(n9906), .A2(n9905), .ZN(n9908) );
  XNOR2_X1 U10721 ( .A(n9908), .B(n9907), .ZN(n9909) );
  AOI222_X1 U10722 ( .A1(n9913), .A2(n9912), .B1(n9911), .B2(n9910), .C1(
        n10758), .C2(n9909), .ZN(n10852) );
  XNOR2_X1 U10723 ( .A(n9914), .B(n9915), .ZN(n10855) );
  INV_X1 U10724 ( .A(n9916), .ZN(n9917) );
  OAI211_X1 U10725 ( .C1(n10853), .C2(n9918), .A(n9917), .B(n10878), .ZN(
        n10851) );
  AOI22_X1 U10726 ( .A1(n10778), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9919), 
        .B2(n10776), .ZN(n9923) );
  NAND2_X1 U10727 ( .A1(n9921), .A2(n9920), .ZN(n9922) );
  OAI211_X1 U10728 ( .C1(n10851), .C2(n9924), .A(n9923), .B(n9922), .ZN(n9925)
         );
  AOI21_X1 U10729 ( .B1(n10855), .B2(n9926), .A(n9925), .ZN(n9927) );
  OAI21_X1 U10730 ( .B1(n10852), .B2(n10778), .A(n9927), .ZN(P1_U3277) );
  NAND2_X1 U10731 ( .A1(n9928), .A2(n10878), .ZN(n9929) );
  OAI211_X1 U10732 ( .C1(n9930), .C2(n10888), .A(n9929), .B(n9932), .ZN(n10003) );
  MUX2_X1 U10733 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n10003), .S(n10722), .Z(
        P1_U3554) );
  NAND2_X1 U10734 ( .A1(n9931), .A2(n10878), .ZN(n9933) );
  OAI211_X1 U10735 ( .C1(n9934), .C2(n10888), .A(n9933), .B(n9932), .ZN(n10004) );
  MUX2_X1 U10736 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n10004), .S(n10722), .Z(
        P1_U3553) );
  AOI22_X1 U10737 ( .A1(n9937), .A2(n10878), .B1(n10877), .B2(n9936), .ZN(
        n9938) );
  NAND3_X1 U10738 ( .A1(n9940), .A2(n9939), .A3(n9938), .ZN(n10005) );
  MUX2_X1 U10739 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n10005), .S(n10722), .Z(
        P1_U3552) );
  AOI22_X1 U10740 ( .A1(n9942), .A2(n10878), .B1(n10877), .B2(n9941), .ZN(
        n9943) );
  OAI211_X1 U10741 ( .C1(n10817), .C2(n9945), .A(n9944), .B(n9943), .ZN(n10006) );
  MUX2_X1 U10742 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n10006), .S(n10722), .Z(
        P1_U3551) );
  INV_X1 U10743 ( .A(n9950), .ZN(n9955) );
  AOI22_X1 U10744 ( .A1(n9952), .A2(n10878), .B1(n10877), .B2(n9951), .ZN(
        n9953) );
  OAI211_X1 U10745 ( .C1(n9955), .C2(n10817), .A(n9954), .B(n9953), .ZN(n10008) );
  MUX2_X1 U10746 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10008), .S(n10722), .Z(
        P1_U3549) );
  OAI21_X1 U10747 ( .B1(n10831), .B2(n9960), .A(n9959), .ZN(n10009) );
  MUX2_X1 U10748 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10009), .S(n10722), .Z(
        P1_U3548) );
  AOI211_X1 U10749 ( .C1(n10877), .C2(n9963), .A(n9962), .B(n9961), .ZN(n9964)
         );
  OAI21_X1 U10750 ( .B1(n10831), .B2(n9965), .A(n9964), .ZN(n10010) );
  MUX2_X1 U10751 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10010), .S(n10722), .Z(
        P1_U3547) );
  AOI22_X1 U10752 ( .A1(n9967), .A2(n10878), .B1(n10877), .B2(n9966), .ZN(
        n9968) );
  OAI211_X1 U10753 ( .C1(n9970), .C2(n10831), .A(n9969), .B(n9968), .ZN(n10011) );
  MUX2_X1 U10754 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10011), .S(n10722), .Z(
        P1_U3546) );
  AOI22_X1 U10755 ( .A1(n9972), .A2(n10878), .B1(n10877), .B2(n9971), .ZN(
        n9973) );
  OAI211_X1 U10756 ( .C1(n10831), .C2(n9975), .A(n9974), .B(n9973), .ZN(n10012) );
  MUX2_X1 U10757 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10012), .S(n10722), .Z(
        P1_U3545) );
  AOI211_X1 U10758 ( .C1(n10877), .C2(n9978), .A(n9977), .B(n9976), .ZN(n9979)
         );
  OAI21_X1 U10759 ( .B1(n10831), .B2(n9980), .A(n9979), .ZN(n10013) );
  MUX2_X1 U10760 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10013), .S(n10722), .Z(
        P1_U3544) );
  AOI22_X1 U10761 ( .A1(n9982), .A2(n10878), .B1(n10877), .B2(n9981), .ZN(
        n9983) );
  OAI211_X1 U10762 ( .C1(n9985), .C2(n10817), .A(n9984), .B(n9983), .ZN(n10014) );
  MUX2_X1 U10763 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10014), .S(n10722), .Z(
        P1_U3543) );
  INV_X1 U10764 ( .A(n9986), .ZN(n9990) );
  AOI22_X1 U10765 ( .A1(n9988), .A2(n10878), .B1(n10877), .B2(n9987), .ZN(
        n9989) );
  OAI211_X1 U10766 ( .C1(n10831), .C2(n9991), .A(n9990), .B(n9989), .ZN(n10015) );
  MUX2_X1 U10767 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10015), .S(n10722), .Z(
        P1_U3542) );
  INV_X1 U10768 ( .A(n9992), .ZN(n9996) );
  AOI22_X1 U10769 ( .A1(n9994), .A2(n10878), .B1(n10877), .B2(n9993), .ZN(
        n9995) );
  OAI211_X1 U10770 ( .C1(n10817), .C2(n9997), .A(n9996), .B(n9995), .ZN(n10016) );
  MUX2_X1 U10771 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10016), .S(n10722), .Z(
        P1_U3541) );
  AOI22_X1 U10772 ( .A1(n9999), .A2(n10878), .B1(n10877), .B2(n9998), .ZN(
        n10000) );
  OAI211_X1 U10773 ( .C1(n10002), .C2(n10831), .A(n10001), .B(n10000), .ZN(
        n10017) );
  MUX2_X1 U10774 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10017), .S(n10722), .Z(
        P1_U3540) );
  MUX2_X1 U10775 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n10003), .S(n5045), .Z(
        P1_U3522) );
  MUX2_X1 U10776 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10004), .S(n5045), .Z(
        P1_U3521) );
  MUX2_X1 U10777 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10005), .S(n5045), .Z(
        P1_U3520) );
  MUX2_X1 U10778 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n10006), .S(n5045), .Z(
        P1_U3519) );
  MUX2_X1 U10779 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10007), .S(n5045), .Z(
        P1_U3518) );
  MUX2_X1 U10780 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10008), .S(n5045), .Z(
        P1_U3517) );
  MUX2_X1 U10781 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10009), .S(n5045), .Z(
        P1_U3516) );
  MUX2_X1 U10782 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10010), .S(n5045), .Z(
        P1_U3515) );
  MUX2_X1 U10783 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10011), .S(n5045), .Z(
        P1_U3514) );
  MUX2_X1 U10784 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10012), .S(n5045), .Z(
        P1_U3513) );
  MUX2_X1 U10785 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10013), .S(n5045), .Z(
        P1_U3512) );
  MUX2_X1 U10786 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10014), .S(n5045), .Z(
        P1_U3511) );
  MUX2_X1 U10787 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10015), .S(n5045), .Z(
        P1_U3510) );
  MUX2_X1 U10788 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10016), .S(n5045), .Z(
        P1_U3508) );
  MUX2_X1 U10789 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10017), .S(n5045), .Z(
        P1_U3505) );
  INV_X1 U10790 ( .A(n10018), .ZN(n10019) );
  NAND2_X1 U10791 ( .A1(n10460), .A2(P1_D_REG_9__SCAN_IN), .ZN(n10440) );
  XOR2_X1 U10792 ( .A(SI_31_), .B(keyinput_1), .Z(n10023) );
  XNOR2_X1 U10793 ( .A(SI_28_), .B(keyinput_4), .ZN(n10022) );
  XNOR2_X1 U10794 ( .A(SI_30_), .B(keyinput_2), .ZN(n10021) );
  NAND3_X1 U10795 ( .A1(n10023), .A2(n10022), .A3(n10021), .ZN(n10026) );
  XNOR2_X1 U10796 ( .A(SI_29_), .B(keyinput_3), .ZN(n10025) );
  XNOR2_X1 U10797 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_0), .ZN(n10024) );
  NOR3_X1 U10798 ( .A1(n10026), .A2(n10025), .A3(n10024), .ZN(n10030) );
  XNOR2_X1 U10799 ( .A(SI_27_), .B(keyinput_5), .ZN(n10029) );
  XNOR2_X1 U10800 ( .A(n10027), .B(keyinput_6), .ZN(n10028) );
  OAI21_X1 U10801 ( .B1(n10030), .B2(n10029), .A(n10028), .ZN(n10038) );
  XNOR2_X1 U10802 ( .A(SI_25_), .B(keyinput_7), .ZN(n10037) );
  XOR2_X1 U10803 ( .A(SI_21_), .B(keyinput_11), .Z(n10035) );
  XOR2_X1 U10804 ( .A(SI_24_), .B(keyinput_8), .Z(n10034) );
  XNOR2_X1 U10805 ( .A(n10031), .B(keyinput_10), .ZN(n10033) );
  XNOR2_X1 U10806 ( .A(SI_23_), .B(keyinput_9), .ZN(n10032) );
  NAND4_X1 U10807 ( .A1(n10035), .A2(n10034), .A3(n10033), .A4(n10032), .ZN(
        n10036) );
  AOI21_X1 U10808 ( .B1(n10038), .B2(n10037), .A(n10036), .ZN(n10043) );
  XNOR2_X1 U10809 ( .A(n10039), .B(keyinput_12), .ZN(n10042) );
  XOR2_X1 U10810 ( .A(SI_18_), .B(keyinput_14), .Z(n10041) );
  XNOR2_X1 U10811 ( .A(SI_19_), .B(keyinput_13), .ZN(n10040) );
  OAI211_X1 U10812 ( .C1(n10043), .C2(n10042), .A(n10041), .B(n10040), .ZN(
        n10046) );
  XOR2_X1 U10813 ( .A(SI_17_), .B(keyinput_15), .Z(n10045) );
  XNOR2_X1 U10814 ( .A(SI_16_), .B(keyinput_16), .ZN(n10044) );
  AOI21_X1 U10815 ( .B1(n10046), .B2(n10045), .A(n10044), .ZN(n10056) );
  XNOR2_X1 U10816 ( .A(SI_15_), .B(keyinput_17), .ZN(n10055) );
  XNOR2_X1 U10817 ( .A(n10047), .B(keyinput_22), .ZN(n10050) );
  XNOR2_X1 U10818 ( .A(SI_14_), .B(keyinput_18), .ZN(n10049) );
  XNOR2_X1 U10819 ( .A(SI_11_), .B(keyinput_21), .ZN(n10048) );
  NAND3_X1 U10820 ( .A1(n10050), .A2(n10049), .A3(n10048), .ZN(n10053) );
  XNOR2_X1 U10821 ( .A(SI_13_), .B(keyinput_19), .ZN(n10052) );
  XNOR2_X1 U10822 ( .A(SI_12_), .B(keyinput_20), .ZN(n10051) );
  NOR3_X1 U10823 ( .A1(n10053), .A2(n10052), .A3(n10051), .ZN(n10054) );
  OAI21_X1 U10824 ( .B1(n10056), .B2(n10055), .A(n10054), .ZN(n10059) );
  XNOR2_X1 U10825 ( .A(n10263), .B(keyinput_23), .ZN(n10058) );
  XNOR2_X1 U10826 ( .A(n10264), .B(keyinput_24), .ZN(n10057) );
  AOI21_X1 U10827 ( .B1(n10059), .B2(n10058), .A(n10057), .ZN(n10062) );
  XNOR2_X1 U10828 ( .A(SI_7_), .B(keyinput_25), .ZN(n10061) );
  XNOR2_X1 U10829 ( .A(SI_6_), .B(keyinput_26), .ZN(n10060) );
  OAI21_X1 U10830 ( .B1(n10062), .B2(n10061), .A(n10060), .ZN(n10067) );
  XNOR2_X1 U10831 ( .A(SI_5_), .B(keyinput_27), .ZN(n10066) );
  XNOR2_X1 U10832 ( .A(n10063), .B(keyinput_29), .ZN(n10065) );
  XNOR2_X1 U10833 ( .A(SI_4_), .B(keyinput_28), .ZN(n10064) );
  AOI211_X1 U10834 ( .C1(n10067), .C2(n10066), .A(n10065), .B(n10064), .ZN(
        n10070) );
  INV_X1 U10835 ( .A(SI_1_), .ZN(n10277) );
  XNOR2_X1 U10836 ( .A(n10277), .B(keyinput_31), .ZN(n10069) );
  XNOR2_X1 U10837 ( .A(SI_2_), .B(keyinput_30), .ZN(n10068) );
  NOR3_X1 U10838 ( .A1(n10070), .A2(n10069), .A3(n10068), .ZN(n10074) );
  XNOR2_X1 U10839 ( .A(SI_0_), .B(keyinput_32), .ZN(n10073) );
  INV_X1 U10840 ( .A(P2_RD_REG_SCAN_IN), .ZN(n10281) );
  XNOR2_X1 U10841 ( .A(n10281), .B(keyinput_33), .ZN(n10072) );
  XNOR2_X1 U10842 ( .A(P2_U3152), .B(keyinput_34), .ZN(n10071) );
  OAI211_X1 U10843 ( .C1(n10074), .C2(n10073), .A(n10072), .B(n10071), .ZN(
        n10079) );
  INV_X1 U10844 ( .A(keyinput_35), .ZN(n10075) );
  XNOR2_X1 U10845 ( .A(n10075), .B(P2_REG3_REG_7__SCAN_IN), .ZN(n10078) );
  XNOR2_X1 U10846 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_36), .ZN(n10077)
         );
  XNOR2_X1 U10847 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_37), .ZN(n10076)
         );
  NAND4_X1 U10848 ( .A1(n10079), .A2(n10078), .A3(n10077), .A4(n10076), .ZN(
        n10092) );
  XNOR2_X1 U10849 ( .A(n10291), .B(keyinput_38), .ZN(n10091) );
  XNOR2_X1 U10850 ( .A(n10080), .B(keyinput_39), .ZN(n10086) );
  XOR2_X1 U10851 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_44), .Z(n10085) );
  XNOR2_X1 U10852 ( .A(n10081), .B(keyinput_41), .ZN(n10084) );
  XNOR2_X1 U10853 ( .A(n10082), .B(keyinput_40), .ZN(n10083) );
  NOR4_X1 U10854 ( .A1(n10086), .A2(n10085), .A3(n10084), .A4(n10083), .ZN(
        n10089) );
  XNOR2_X1 U10855 ( .A(n10293), .B(keyinput_43), .ZN(n10088) );
  XNOR2_X1 U10856 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_42), .ZN(n10087)
         );
  NAND3_X1 U10857 ( .A1(n10089), .A2(n10088), .A3(n10087), .ZN(n10090) );
  AOI21_X1 U10858 ( .B1(n10092), .B2(n10091), .A(n10090), .ZN(n10095) );
  XNOR2_X1 U10859 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput_46), .ZN(n10094)
         );
  XNOR2_X1 U10860 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput_45), .ZN(n10093)
         );
  NOR3_X1 U10861 ( .A1(n10095), .A2(n10094), .A3(n10093), .ZN(n10100) );
  XNOR2_X1 U10862 ( .A(n10096), .B(keyinput_49), .ZN(n10099) );
  XNOR2_X1 U10863 ( .A(n10309), .B(keyinput_47), .ZN(n10098) );
  XNOR2_X1 U10864 ( .A(n10308), .B(keyinput_48), .ZN(n10097) );
  NOR4_X1 U10865 ( .A1(n10100), .A2(n10099), .A3(n10098), .A4(n10097), .ZN(
        n10104) );
  XNOR2_X1 U10866 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput_50), .ZN(n10103)
         );
  XNOR2_X1 U10867 ( .A(n10314), .B(keyinput_51), .ZN(n10102) );
  XNOR2_X1 U10868 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_52), .ZN(n10101)
         );
  OAI211_X1 U10869 ( .C1(n10104), .C2(n10103), .A(n10102), .B(n10101), .ZN(
        n10113) );
  XNOR2_X1 U10870 ( .A(n10105), .B(keyinput_53), .ZN(n10112) );
  XNOR2_X1 U10871 ( .A(n10106), .B(keyinput_57), .ZN(n10110) );
  XNOR2_X1 U10872 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput_55), .ZN(n10109)
         );
  XNOR2_X1 U10873 ( .A(P2_REG3_REG_13__SCAN_IN), .B(keyinput_56), .ZN(n10108)
         );
  XNOR2_X1 U10874 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_54), .ZN(n10107)
         );
  NAND4_X1 U10875 ( .A1(n10110), .A2(n10109), .A3(n10108), .A4(n10107), .ZN(
        n10111) );
  AOI21_X1 U10876 ( .B1(n10113), .B2(n10112), .A(n10111), .ZN(n10116) );
  XOR2_X1 U10877 ( .A(P2_REG3_REG_11__SCAN_IN), .B(keyinput_58), .Z(n10115) );
  XNOR2_X1 U10878 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_59), .ZN(n10114)
         );
  NOR3_X1 U10879 ( .A1(n10116), .A2(n10115), .A3(n10114), .ZN(n10120) );
  XNOR2_X1 U10880 ( .A(n10117), .B(keyinput_60), .ZN(n10119) );
  XNOR2_X1 U10881 ( .A(n10331), .B(keyinput_61), .ZN(n10118) );
  OAI21_X1 U10882 ( .B1(n10120), .B2(n10119), .A(n10118), .ZN(n10124) );
  XNOR2_X1 U10883 ( .A(n10121), .B(keyinput_63), .ZN(n10123) );
  XNOR2_X1 U10884 ( .A(P2_REG3_REG_26__SCAN_IN), .B(keyinput_62), .ZN(n10122)
         );
  NAND3_X1 U10885 ( .A1(n10124), .A2(n10123), .A3(n10122), .ZN(n10127) );
  XNOR2_X1 U10886 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_64), .ZN(n10126) );
  XNOR2_X1 U10887 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_65), .ZN(n10125)
         );
  NAND3_X1 U10888 ( .A1(n10127), .A2(n10126), .A3(n10125), .ZN(n10130) );
  XOR2_X1 U10889 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(keyinput_66), .Z(n10129)
         );
  XNOR2_X1 U10890 ( .A(n10448), .B(keyinput_67), .ZN(n10128) );
  AOI21_X1 U10891 ( .B1(n10130), .B2(n10129), .A(n10128), .ZN(n10134) );
  XOR2_X1 U10892 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_68), .Z(n10133)
         );
  XOR2_X1 U10893 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput_69), .Z(n10132)
         );
  XNOR2_X1 U10894 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(keyinput_70), .ZN(n10131)
         );
  NOR4_X1 U10895 ( .A1(n10134), .A2(n10133), .A3(n10132), .A4(n10131), .ZN(
        n10137) );
  XOR2_X1 U10896 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_71), .Z(n10136)
         );
  XOR2_X1 U10897 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_72), .Z(n10135)
         );
  NOR3_X1 U10898 ( .A1(n10137), .A2(n10136), .A3(n10135), .ZN(n10140) );
  XNOR2_X1 U10899 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput_73), .ZN(n10139)
         );
  XOR2_X1 U10900 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_74), .Z(n10138)
         );
  OAI21_X1 U10901 ( .B1(n10140), .B2(n10139), .A(n10138), .ZN(n10143) );
  XNOR2_X1 U10902 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_75), .ZN(n10142)
         );
  XNOR2_X1 U10903 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(keyinput_76), .ZN(n10141)
         );
  NAND3_X1 U10904 ( .A1(n10143), .A2(n10142), .A3(n10141), .ZN(n10146) );
  XOR2_X1 U10905 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_78), .Z(n10145)
         );
  XNOR2_X1 U10906 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_77), .ZN(n10144)
         );
  NAND3_X1 U10907 ( .A1(n10146), .A2(n10145), .A3(n10144), .ZN(n10153) );
  XOR2_X1 U10908 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_79), .Z(n10150)
         );
  XOR2_X1 U10909 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(keyinput_80), .Z(n10149)
         );
  XOR2_X1 U10910 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_81), .Z(n10148)
         );
  XOR2_X1 U10911 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput_82), .Z(n10147)
         );
  NOR4_X1 U10912 ( .A1(n10150), .A2(n10149), .A3(n10148), .A4(n10147), .ZN(
        n10152) );
  XNOR2_X1 U10913 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_83), .ZN(n10151)
         );
  AOI21_X1 U10914 ( .B1(n10153), .B2(n10152), .A(n10151), .ZN(n10156) );
  XOR2_X1 U10915 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_84), .Z(n10155)
         );
  XNOR2_X1 U10916 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_85), .ZN(n10154)
         );
  OAI21_X1 U10917 ( .B1(n10156), .B2(n10155), .A(n10154), .ZN(n10159) );
  XOR2_X1 U10918 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_86), .Z(n10158)
         );
  XOR2_X1 U10919 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput_87), .Z(n10157) );
  AOI21_X1 U10920 ( .B1(n10159), .B2(n10158), .A(n10157), .ZN(n10163) );
  XOR2_X1 U10921 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_89), .Z(n10162) );
  XOR2_X1 U10922 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_88), .Z(n10161) );
  XNOR2_X1 U10923 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput_90), .ZN(n10160)
         );
  NOR4_X1 U10924 ( .A1(n10163), .A2(n10162), .A3(n10161), .A4(n10160), .ZN(
        n10173) );
  XNOR2_X1 U10925 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_91), .ZN(n10172) );
  XOR2_X1 U10926 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_92), .Z(n10170) );
  XNOR2_X1 U10927 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_96), .ZN(n10166) );
  XNOR2_X1 U10928 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_95), .ZN(n10165) );
  XNOR2_X1 U10929 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_94), .ZN(n10164) );
  NAND3_X1 U10930 ( .A1(n10166), .A2(n10165), .A3(n10164), .ZN(n10169) );
  XNOR2_X1 U10931 ( .A(n10167), .B(keyinput_93), .ZN(n10168) );
  NOR3_X1 U10932 ( .A1(n10170), .A2(n10169), .A3(n10168), .ZN(n10171) );
  OAI21_X1 U10933 ( .B1(n10173), .B2(n10172), .A(n10171), .ZN(n10178) );
  XNOR2_X1 U10934 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_97), .ZN(n10177) );
  XNOR2_X1 U10935 ( .A(n10174), .B(keyinput_99), .ZN(n10176) );
  XNOR2_X1 U10936 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_98), .ZN(n10175) );
  AOI211_X1 U10937 ( .C1(n10178), .C2(n10177), .A(n10176), .B(n10175), .ZN(
        n10182) );
  XOR2_X1 U10938 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_100), .Z(n10181) );
  XNOR2_X1 U10939 ( .A(n10390), .B(keyinput_101), .ZN(n10180) );
  XNOR2_X1 U10940 ( .A(n10391), .B(keyinput_102), .ZN(n10179) );
  NOR4_X1 U10941 ( .A1(n10182), .A2(n10181), .A3(n10180), .A4(n10179), .ZN(
        n10185) );
  XNOR2_X1 U10942 ( .A(n10396), .B(keyinput_103), .ZN(n10184) );
  XNOR2_X1 U10943 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_104), .ZN(n10183)
         );
  NOR3_X1 U10944 ( .A1(n10185), .A2(n10184), .A3(n10183), .ZN(n10188) );
  XNOR2_X1 U10945 ( .A(n10401), .B(keyinput_105), .ZN(n10187) );
  XOR2_X1 U10946 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_106), .Z(n10186) );
  NOR3_X1 U10947 ( .A1(n10188), .A2(n10187), .A3(n10186), .ZN(n10191) );
  XNOR2_X1 U10948 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_107), .ZN(n10190)
         );
  XNOR2_X1 U10949 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_108), .ZN(n10189)
         );
  OAI21_X1 U10950 ( .B1(n10191), .B2(n10190), .A(n10189), .ZN(n10195) );
  XNOR2_X1 U10951 ( .A(n10192), .B(keyinput_109), .ZN(n10194) );
  XNOR2_X1 U10952 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_110), .ZN(n10193)
         );
  NAND3_X1 U10953 ( .A1(n10195), .A2(n10194), .A3(n10193), .ZN(n10199) );
  XNOR2_X1 U10954 ( .A(n10196), .B(keyinput_112), .ZN(n10198) );
  XNOR2_X1 U10955 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_111), .ZN(n10197)
         );
  NAND3_X1 U10956 ( .A1(n10199), .A2(n10198), .A3(n10197), .ZN(n10203) );
  XNOR2_X1 U10957 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_113), .ZN(n10202)
         );
  XNOR2_X1 U10958 ( .A(n10200), .B(keyinput_114), .ZN(n10201) );
  AOI21_X1 U10959 ( .B1(n10203), .B2(n10202), .A(n10201), .ZN(n10207) );
  XNOR2_X1 U10960 ( .A(n10204), .B(keyinput_115), .ZN(n10206) );
  XNOR2_X1 U10961 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_116), .ZN(n10205)
         );
  OAI21_X1 U10962 ( .B1(n10207), .B2(n10206), .A(n10205), .ZN(n10212) );
  XNOR2_X1 U10963 ( .A(n10208), .B(keyinput_118), .ZN(n10211) );
  XOR2_X1 U10964 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_119), .Z(n10210) );
  XNOR2_X1 U10965 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_117), .ZN(n10209)
         );
  NAND4_X1 U10966 ( .A1(n10212), .A2(n10211), .A3(n10210), .A4(n10209), .ZN(
        n10224) );
  XNOR2_X1 U10967 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_120), .ZN(n10223)
         );
  XNOR2_X1 U10968 ( .A(n10213), .B(keyinput_123), .ZN(n10218) );
  INV_X1 U10969 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10457) );
  XNOR2_X1 U10970 ( .A(n10457), .B(keyinput_125), .ZN(n10217) );
  INV_X1 U10971 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10458) );
  XNOR2_X1 U10972 ( .A(n10458), .B(keyinput_126), .ZN(n10216) );
  XNOR2_X1 U10973 ( .A(n10214), .B(keyinput_124), .ZN(n10215) );
  NOR4_X1 U10974 ( .A1(n10218), .A2(n10217), .A3(n10216), .A4(n10215), .ZN(
        n10221) );
  XOR2_X1 U10975 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_121), .Z(n10220) );
  XOR2_X1 U10976 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_122), .Z(n10219) );
  NAND3_X1 U10977 ( .A1(n10221), .A2(n10220), .A3(n10219), .ZN(n10222) );
  AOI21_X1 U10978 ( .B1(n10224), .B2(n10223), .A(n10222), .ZN(n10438) );
  XNOR2_X1 U10979 ( .A(keyinput_255), .B(keyinput_127), .ZN(n10437) );
  XOR2_X1 U10980 ( .A(keyinput_255), .B(P1_D_REG_4__SCAN_IN), .Z(n10436) );
  XOR2_X1 U10981 ( .A(SI_30_), .B(keyinput_130), .Z(n10228) );
  XNOR2_X1 U10982 ( .A(n10225), .B(keyinput_132), .ZN(n10227) );
  XNOR2_X1 U10983 ( .A(SI_31_), .B(keyinput_129), .ZN(n10226) );
  NOR3_X1 U10984 ( .A1(n10228), .A2(n10227), .A3(n10226), .ZN(n10232) );
  XNOR2_X1 U10985 ( .A(n10229), .B(keyinput_131), .ZN(n10231) );
  XOR2_X1 U10986 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_128), .Z(n10230) );
  NAND3_X1 U10987 ( .A1(n10232), .A2(n10231), .A3(n10230), .ZN(n10235) );
  XNOR2_X1 U10988 ( .A(SI_27_), .B(keyinput_133), .ZN(n10234) );
  XNOR2_X1 U10989 ( .A(SI_26_), .B(keyinput_134), .ZN(n10233) );
  AOI21_X1 U10990 ( .B1(n10235), .B2(n10234), .A(n10233), .ZN(n10243) );
  XNOR2_X1 U10991 ( .A(SI_25_), .B(keyinput_135), .ZN(n10242) );
  XOR2_X1 U10992 ( .A(SI_24_), .B(keyinput_136), .Z(n10240) );
  XOR2_X1 U10993 ( .A(SI_21_), .B(keyinput_139), .Z(n10239) );
  XNOR2_X1 U10994 ( .A(n10236), .B(keyinput_137), .ZN(n10238) );
  XNOR2_X1 U10995 ( .A(SI_22_), .B(keyinput_138), .ZN(n10237) );
  NOR4_X1 U10996 ( .A1(n10240), .A2(n10239), .A3(n10238), .A4(n10237), .ZN(
        n10241) );
  OAI21_X1 U10997 ( .B1(n10243), .B2(n10242), .A(n10241), .ZN(n10248) );
  XNOR2_X1 U10998 ( .A(SI_20_), .B(keyinput_140), .ZN(n10247) );
  XNOR2_X1 U10999 ( .A(n10244), .B(keyinput_141), .ZN(n10246) );
  XNOR2_X1 U11000 ( .A(SI_18_), .B(keyinput_142), .ZN(n10245) );
  AOI211_X1 U11001 ( .C1(n10248), .C2(n10247), .A(n10246), .B(n10245), .ZN(
        n10251) );
  XOR2_X1 U11002 ( .A(SI_17_), .B(keyinput_143), .Z(n10250) );
  XOR2_X1 U11003 ( .A(SI_16_), .B(keyinput_144), .Z(n10249) );
  OAI21_X1 U11004 ( .B1(n10251), .B2(n10250), .A(n10249), .ZN(n10262) );
  XNOR2_X1 U11005 ( .A(n10252), .B(keyinput_145), .ZN(n10261) );
  OAI22_X1 U11006 ( .A1(n10254), .A2(keyinput_148), .B1(SI_14_), .B2(
        keyinput_146), .ZN(n10253) );
  AOI221_X1 U11007 ( .B1(n10254), .B2(keyinput_148), .C1(keyinput_146), .C2(
        SI_14_), .A(n10253), .ZN(n10259) );
  XNOR2_X1 U11008 ( .A(n10255), .B(keyinput_147), .ZN(n10258) );
  XNOR2_X1 U11009 ( .A(SI_10_), .B(keyinput_150), .ZN(n10257) );
  XNOR2_X1 U11010 ( .A(SI_11_), .B(keyinput_149), .ZN(n10256) );
  NAND4_X1 U11011 ( .A1(n10259), .A2(n10258), .A3(n10257), .A4(n10256), .ZN(
        n10260) );
  AOI21_X1 U11012 ( .B1(n10262), .B2(n10261), .A(n10260), .ZN(n10267) );
  XNOR2_X1 U11013 ( .A(n10263), .B(keyinput_151), .ZN(n10266) );
  XNOR2_X1 U11014 ( .A(n10264), .B(keyinput_152), .ZN(n10265) );
  OAI21_X1 U11015 ( .B1(n10267), .B2(n10266), .A(n10265), .ZN(n10270) );
  XOR2_X1 U11016 ( .A(SI_7_), .B(keyinput_153), .Z(n10269) );
  XNOR2_X1 U11017 ( .A(SI_6_), .B(keyinput_154), .ZN(n10268) );
  AOI21_X1 U11018 ( .B1(n10270), .B2(n10269), .A(n10268), .ZN(n10275) );
  XNOR2_X1 U11019 ( .A(SI_5_), .B(keyinput_155), .ZN(n10274) );
  XNOR2_X1 U11020 ( .A(n10271), .B(keyinput_156), .ZN(n10273) );
  XNOR2_X1 U11021 ( .A(SI_3_), .B(keyinput_157), .ZN(n10272) );
  OAI211_X1 U11022 ( .C1(n10275), .C2(n10274), .A(n10273), .B(n10272), .ZN(
        n10280) );
  XNOR2_X1 U11023 ( .A(n10276), .B(keyinput_158), .ZN(n10279) );
  XNOR2_X1 U11024 ( .A(n10277), .B(keyinput_159), .ZN(n10278) );
  NAND3_X1 U11025 ( .A1(n10280), .A2(n10279), .A3(n10278), .ZN(n10285) );
  XOR2_X1 U11026 ( .A(SI_0_), .B(keyinput_160), .Z(n10284) );
  XNOR2_X1 U11027 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_161), .ZN(n10283) );
  XNOR2_X1 U11028 ( .A(P2_STATE_REG_SCAN_IN), .B(keyinput_162), .ZN(n10282) );
  AOI211_X1 U11029 ( .C1(n10285), .C2(n10284), .A(n10283), .B(n10282), .ZN(
        n10290) );
  XNOR2_X1 U11030 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput_163), .ZN(n10289)
         );
  XNOR2_X1 U11031 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_164), .ZN(n10287)
         );
  XNOR2_X1 U11032 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_165), .ZN(n10286)
         );
  NAND2_X1 U11033 ( .A1(n10287), .A2(n10286), .ZN(n10288) );
  NOR3_X1 U11034 ( .A1(n10290), .A2(n10289), .A3(n10288), .ZN(n10303) );
  XNOR2_X1 U11035 ( .A(n10291), .B(keyinput_166), .ZN(n10302) );
  XOR2_X1 U11036 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_172), .Z(n10297) );
  XNOR2_X1 U11037 ( .A(n10292), .B(keyinput_170), .ZN(n10296) );
  XNOR2_X1 U11038 ( .A(n10293), .B(keyinput_171), .ZN(n10295) );
  XNOR2_X1 U11039 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_168), .ZN(n10294)
         );
  NAND4_X1 U11040 ( .A1(n10297), .A2(n10296), .A3(n10295), .A4(n10294), .ZN(
        n10300) );
  XNOR2_X1 U11041 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_167), .ZN(n10299)
         );
  XNOR2_X1 U11042 ( .A(P2_REG3_REG_19__SCAN_IN), .B(keyinput_169), .ZN(n10298)
         );
  NOR3_X1 U11043 ( .A1(n10300), .A2(n10299), .A3(n10298), .ZN(n10301) );
  OAI21_X1 U11044 ( .B1(n10303), .B2(n10302), .A(n10301), .ZN(n10307) );
  XNOR2_X1 U11045 ( .A(n10304), .B(keyinput_174), .ZN(n10306) );
  XOR2_X1 U11046 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput_173), .Z(n10305)
         );
  NAND3_X1 U11047 ( .A1(n10307), .A2(n10306), .A3(n10305), .ZN(n10313) );
  XNOR2_X1 U11048 ( .A(n10308), .B(keyinput_176), .ZN(n10312) );
  XNOR2_X1 U11049 ( .A(n10309), .B(keyinput_175), .ZN(n10311) );
  XNOR2_X1 U11050 ( .A(P2_REG3_REG_5__SCAN_IN), .B(keyinput_177), .ZN(n10310)
         );
  NAND4_X1 U11051 ( .A1(n10313), .A2(n10312), .A3(n10311), .A4(n10310), .ZN(
        n10318) );
  XNOR2_X1 U11052 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput_178), .ZN(n10317)
         );
  XOR2_X1 U11053 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_180), .Z(n10316) );
  XNOR2_X1 U11054 ( .A(n10314), .B(keyinput_179), .ZN(n10315) );
  AOI211_X1 U11055 ( .C1(n10318), .C2(n10317), .A(n10316), .B(n10315), .ZN(
        n10327) );
  XNOR2_X1 U11056 ( .A(P2_REG3_REG_9__SCAN_IN), .B(keyinput_181), .ZN(n10326)
         );
  XOR2_X1 U11057 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_182), .Z(n10324) );
  XNOR2_X1 U11058 ( .A(n10319), .B(keyinput_184), .ZN(n10323) );
  XNOR2_X1 U11059 ( .A(n10320), .B(keyinput_183), .ZN(n10322) );
  XNOR2_X1 U11060 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput_185), .ZN(n10321)
         );
  NOR4_X1 U11061 ( .A1(n10324), .A2(n10323), .A3(n10322), .A4(n10321), .ZN(
        n10325) );
  OAI21_X1 U11062 ( .B1(n10327), .B2(n10326), .A(n10325), .ZN(n10330) );
  XOR2_X1 U11063 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_187), .Z(n10329) );
  XNOR2_X1 U11064 ( .A(P2_REG3_REG_11__SCAN_IN), .B(keyinput_186), .ZN(n10328)
         );
  NAND3_X1 U11065 ( .A1(n10330), .A2(n10329), .A3(n10328), .ZN(n10334) );
  XNOR2_X1 U11066 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_188), .ZN(n10333)
         );
  XNOR2_X1 U11067 ( .A(n10331), .B(keyinput_189), .ZN(n10332) );
  AOI21_X1 U11068 ( .B1(n10334), .B2(n10333), .A(n10332), .ZN(n10337) );
  XNOR2_X1 U11069 ( .A(P2_REG3_REG_15__SCAN_IN), .B(keyinput_191), .ZN(n10336)
         );
  XNOR2_X1 U11070 ( .A(P2_REG3_REG_26__SCAN_IN), .B(keyinput_190), .ZN(n10335)
         );
  NOR3_X1 U11071 ( .A1(n10337), .A2(n10336), .A3(n10335), .ZN(n10340) );
  XOR2_X1 U11072 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_192), .Z(n10339) );
  XNOR2_X1 U11073 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_193), .ZN(n10338) );
  NOR3_X1 U11074 ( .A1(n10340), .A2(n10339), .A3(n10338), .ZN(n10343) );
  XNOR2_X1 U11075 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(keyinput_194), .ZN(n10342) );
  XNOR2_X1 U11076 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput_195), .ZN(n10341) );
  OAI21_X1 U11077 ( .B1(n10343), .B2(n10342), .A(n10341), .ZN(n10347) );
  XOR2_X1 U11078 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput_197), .Z(n10346)
         );
  XNOR2_X1 U11079 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(keyinput_198), .ZN(n10345) );
  XNOR2_X1 U11080 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_196), .ZN(n10344) );
  NAND4_X1 U11081 ( .A1(n10347), .A2(n10346), .A3(n10345), .A4(n10344), .ZN(
        n10350) );
  XOR2_X1 U11082 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_200), .Z(n10349)
         );
  XOR2_X1 U11083 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_199), .Z(n10348)
         );
  NAND3_X1 U11084 ( .A1(n10350), .A2(n10349), .A3(n10348), .ZN(n10353) );
  XOR2_X1 U11085 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput_201), .Z(n10352)
         );
  XNOR2_X1 U11086 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_202), .ZN(n10351) );
  AOI21_X1 U11087 ( .B1(n10353), .B2(n10352), .A(n10351), .ZN(n10356) );
  XOR2_X1 U11088 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_203), .Z(n10355)
         );
  XNOR2_X1 U11089 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(keyinput_204), .ZN(n10354) );
  NOR3_X1 U11090 ( .A1(n10356), .A2(n10355), .A3(n10354), .ZN(n10359) );
  XOR2_X1 U11091 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_205), .Z(n10358)
         );
  XOR2_X1 U11092 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_206), .Z(n10357)
         );
  NOR3_X1 U11093 ( .A1(n10359), .A2(n10358), .A3(n10357), .ZN(n10366) );
  XOR2_X1 U11094 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_209), .Z(n10363)
         );
  XOR2_X1 U11095 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput_210), .Z(n10362)
         );
  XNOR2_X1 U11096 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(keyinput_208), .ZN(n10361) );
  XNOR2_X1 U11097 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_207), .ZN(n10360) );
  NAND4_X1 U11098 ( .A1(n10363), .A2(n10362), .A3(n10361), .A4(n10360), .ZN(
        n10365) );
  XNOR2_X1 U11099 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_211), .ZN(n10364) );
  OAI21_X1 U11100 ( .B1(n10366), .B2(n10365), .A(n10364), .ZN(n10369) );
  XOR2_X1 U11101 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_212), .Z(n10368)
         );
  XNOR2_X1 U11102 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_213), .ZN(n10367) );
  AOI21_X1 U11103 ( .B1(n10369), .B2(n10368), .A(n10367), .ZN(n10372) );
  XOR2_X1 U11104 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_214), .Z(n10371)
         );
  XOR2_X1 U11105 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput_215), .Z(n10370)
         );
  OAI21_X1 U11106 ( .B1(n10372), .B2(n10371), .A(n10370), .ZN(n10376) );
  XOR2_X1 U11107 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_216), .Z(n10375)
         );
  XNOR2_X1 U11108 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_217), .ZN(n10374)
         );
  XNOR2_X1 U11109 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput_218), .ZN(n10373)
         );
  NAND4_X1 U11110 ( .A1(n10376), .A2(n10375), .A3(n10374), .A4(n10373), .ZN(
        n10385) );
  XNOR2_X1 U11111 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_219), .ZN(n10384) );
  INV_X1 U11112 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n10378) );
  AOI22_X1 U11113 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(keyinput_221), .B1(n10378), 
        .B2(keyinput_222), .ZN(n10377) );
  OAI221_X1 U11114 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(keyinput_221), .C1(n10378), 
        .C2(keyinput_222), .A(n10377), .ZN(n10383) );
  XOR2_X1 U11115 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_224), .Z(n10381) );
  XNOR2_X1 U11116 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_220), .ZN(n10380) );
  XNOR2_X1 U11117 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_223), .ZN(n10379) );
  NAND3_X1 U11118 ( .A1(n10381), .A2(n10380), .A3(n10379), .ZN(n10382) );
  AOI211_X1 U11119 ( .C1(n10385), .C2(n10384), .A(n10383), .B(n10382), .ZN(
        n10389) );
  XNOR2_X1 U11120 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_225), .ZN(n10388) );
  XNOR2_X1 U11121 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_226), .ZN(n10387) );
  XNOR2_X1 U11122 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_227), .ZN(n10386) );
  OAI211_X1 U11123 ( .C1(n10389), .C2(n10388), .A(n10387), .B(n10386), .ZN(
        n10395) );
  XNOR2_X1 U11124 ( .A(n10390), .B(keyinput_229), .ZN(n10394) );
  XOR2_X1 U11125 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_228), .Z(n10393) );
  XNOR2_X1 U11126 ( .A(n10391), .B(keyinput_230), .ZN(n10392) );
  NAND4_X1 U11127 ( .A1(n10395), .A2(n10394), .A3(n10393), .A4(n10392), .ZN(
        n10400) );
  XNOR2_X1 U11128 ( .A(n10396), .B(keyinput_231), .ZN(n10399) );
  XNOR2_X1 U11129 ( .A(n10397), .B(keyinput_232), .ZN(n10398) );
  NAND3_X1 U11130 ( .A1(n10400), .A2(n10399), .A3(n10398), .ZN(n10404) );
  XNOR2_X1 U11131 ( .A(n10401), .B(keyinput_233), .ZN(n10403) );
  XNOR2_X1 U11132 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_234), .ZN(n10402)
         );
  NAND3_X1 U11133 ( .A1(n10404), .A2(n10403), .A3(n10402), .ZN(n10408) );
  XNOR2_X1 U11134 ( .A(n10405), .B(keyinput_235), .ZN(n10407) );
  XNOR2_X1 U11135 ( .A(n6598), .B(keyinput_236), .ZN(n10406) );
  AOI21_X1 U11136 ( .B1(n10408), .B2(n10407), .A(n10406), .ZN(n10411) );
  XNOR2_X1 U11137 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_237), .ZN(n10410)
         );
  XNOR2_X1 U11138 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_238), .ZN(n10409)
         );
  NOR3_X1 U11139 ( .A1(n10411), .A2(n10410), .A3(n10409), .ZN(n10414) );
  XNOR2_X1 U11140 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_239), .ZN(n10413)
         );
  XNOR2_X1 U11141 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_240), .ZN(n10412)
         );
  NOR3_X1 U11142 ( .A1(n10414), .A2(n10413), .A3(n10412), .ZN(n10417) );
  XNOR2_X1 U11143 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_241), .ZN(n10416)
         );
  XNOR2_X1 U11144 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_242), .ZN(n10415)
         );
  OAI21_X1 U11145 ( .B1(n10417), .B2(n10416), .A(n10415), .ZN(n10420) );
  XNOR2_X1 U11146 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_243), .ZN(n10419)
         );
  XNOR2_X1 U11147 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_244), .ZN(n10418)
         );
  AOI21_X1 U11148 ( .B1(n10420), .B2(n10419), .A(n10418), .ZN(n10424) );
  XNOR2_X1 U11149 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_247), .ZN(n10423)
         );
  XNOR2_X1 U11150 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_246), .ZN(n10422)
         );
  XNOR2_X1 U11151 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_245), .ZN(n10421)
         );
  NOR4_X1 U11152 ( .A1(n10424), .A2(n10423), .A3(n10422), .A4(n10421), .ZN(
        n10434) );
  XOR2_X1 U11153 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_248), .Z(n10433) );
  XOR2_X1 U11154 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_250), .Z(n10428) );
  XOR2_X1 U11155 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_249), .Z(n10427) );
  XNOR2_X1 U11156 ( .A(P1_D_REG_3__SCAN_IN), .B(keyinput_254), .ZN(n10426) );
  XNOR2_X1 U11157 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput_251), .ZN(n10425) );
  NAND4_X1 U11158 ( .A1(n10428), .A2(n10427), .A3(n10426), .A4(n10425), .ZN(
        n10431) );
  XNOR2_X1 U11159 ( .A(P1_D_REG_2__SCAN_IN), .B(keyinput_253), .ZN(n10430) );
  XNOR2_X1 U11160 ( .A(P1_D_REG_1__SCAN_IN), .B(keyinput_252), .ZN(n10429) );
  NOR3_X1 U11161 ( .A1(n10431), .A2(n10430), .A3(n10429), .ZN(n10432) );
  OAI21_X1 U11162 ( .B1(n10434), .B2(n10433), .A(n10432), .ZN(n10435) );
  OAI211_X1 U11163 ( .C1(n10438), .C2(n10437), .A(n10436), .B(n10435), .ZN(
        n10439) );
  XOR2_X1 U11164 ( .A(n10440), .B(n10439), .Z(P1_U3314) );
  MUX2_X1 U11165 ( .A(n10442), .B(P1_D_REG_0__SCAN_IN), .S(n10441), .Z(
        P1_U3440) );
  NOR4_X1 U11166 ( .A1(n10443), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), 
        .A4(n5884), .ZN(n10444) );
  AOI21_X1 U11167 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n10445), .A(n10444), 
        .ZN(n10446) );
  OAI21_X1 U11168 ( .B1(n10447), .B2(n10451), .A(n10446), .ZN(P1_U3322) );
  OAI222_X1 U11169 ( .A1(n10451), .A2(n10450), .B1(n10449), .B2(P1_U3084), 
        .C1(n10448), .C2(n10455), .ZN(P1_U3324) );
  INV_X1 U11170 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10454) );
  OAI222_X1 U11171 ( .A1(n10455), .A2(n10454), .B1(n10451), .B2(n10453), .C1(
        P1_U3084), .C2(n10452), .ZN(P1_U3325) );
  MUX2_X1 U11172 ( .A(n10456), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U11173 ( .A(n10460), .ZN(n10459) );
  NOR2_X1 U11174 ( .A1(n10459), .A2(n10457), .ZN(P1_U3321) );
  NOR2_X1 U11175 ( .A1(n10459), .A2(n10458), .ZN(P1_U3320) );
  AND2_X1 U11176 ( .A1(n10460), .A2(P1_D_REG_4__SCAN_IN), .ZN(P1_U3319) );
  AND2_X1 U11177 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10460), .ZN(P1_U3318) );
  AND2_X1 U11178 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10460), .ZN(P1_U3317) );
  AND2_X1 U11179 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10460), .ZN(P1_U3316) );
  AND2_X1 U11180 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10460), .ZN(P1_U3315) );
  AND2_X1 U11181 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10460), .ZN(P1_U3313) );
  AND2_X1 U11182 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10460), .ZN(P1_U3312) );
  AND2_X1 U11183 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10460), .ZN(P1_U3311) );
  AND2_X1 U11184 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10460), .ZN(P1_U3310) );
  AND2_X1 U11185 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10460), .ZN(P1_U3309) );
  AND2_X1 U11186 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10460), .ZN(P1_U3308) );
  AND2_X1 U11187 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10460), .ZN(P1_U3307) );
  AND2_X1 U11188 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10460), .ZN(P1_U3306) );
  AND2_X1 U11189 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10460), .ZN(P1_U3305) );
  AND2_X1 U11190 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10460), .ZN(P1_U3304) );
  AND2_X1 U11191 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10460), .ZN(P1_U3303) );
  AND2_X1 U11192 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10460), .ZN(P1_U3302) );
  AND2_X1 U11193 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10460), .ZN(P1_U3301) );
  AND2_X1 U11194 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10460), .ZN(P1_U3300) );
  AND2_X1 U11195 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10460), .ZN(P1_U3299) );
  AND2_X1 U11196 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10460), .ZN(P1_U3298) );
  AND2_X1 U11197 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10460), .ZN(P1_U3297) );
  AND2_X1 U11198 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10460), .ZN(P1_U3296) );
  AND2_X1 U11199 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10460), .ZN(P1_U3295) );
  AND2_X1 U11200 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10460), .ZN(P1_U3294) );
  AND2_X1 U11201 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10460), .ZN(P1_U3293) );
  AND2_X1 U11202 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10460), .ZN(P1_U3292) );
  AOI22_X1 U11203 ( .A1(n10583), .A2(n10464), .B1(n10463), .B2(n10580), .ZN(
        P2_U3438) );
  AND2_X1 U11204 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10580), .ZN(P2_U3326) );
  AND2_X1 U11205 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10580), .ZN(P2_U3325) );
  AND2_X1 U11206 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10580), .ZN(P2_U3324) );
  AND2_X1 U11207 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10580), .ZN(P2_U3323) );
  AND2_X1 U11208 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10580), .ZN(P2_U3322) );
  AND2_X1 U11209 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10580), .ZN(P2_U3321) );
  AND2_X1 U11210 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10580), .ZN(P2_U3320) );
  AND2_X1 U11211 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10580), .ZN(P2_U3319) );
  AND2_X1 U11212 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10580), .ZN(P2_U3318) );
  AND2_X1 U11213 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10580), .ZN(P2_U3317) );
  AND2_X1 U11214 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10580), .ZN(P2_U3316) );
  AND2_X1 U11215 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10580), .ZN(P2_U3315) );
  AND2_X1 U11216 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10580), .ZN(P2_U3314) );
  AND2_X1 U11217 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10580), .ZN(P2_U3313) );
  AND2_X1 U11218 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10580), .ZN(P2_U3312) );
  AND2_X1 U11219 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10580), .ZN(P2_U3311) );
  AND2_X1 U11220 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10580), .ZN(P2_U3310) );
  AND2_X1 U11221 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10580), .ZN(P2_U3309) );
  AND2_X1 U11222 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10580), .ZN(P2_U3308) );
  AND2_X1 U11223 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10580), .ZN(P2_U3307) );
  AND2_X1 U11224 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10580), .ZN(P2_U3306) );
  AND2_X1 U11225 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10580), .ZN(P2_U3305) );
  AND2_X1 U11226 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10580), .ZN(P2_U3304) );
  AND2_X1 U11227 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10580), .ZN(P2_U3303) );
  AND2_X1 U11228 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10580), .ZN(P2_U3302) );
  AND2_X1 U11229 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10580), .ZN(P2_U3301) );
  AND2_X1 U11230 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10580), .ZN(P2_U3300) );
  AND2_X1 U11231 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10580), .ZN(P2_U3299) );
  AND2_X1 U11232 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10580), .ZN(P2_U3298) );
  AND2_X1 U11233 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10580), .ZN(P2_U3297) );
  XOR2_X1 U11234 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  INV_X1 U11235 ( .A(n10465), .ZN(n10466) );
  NAND2_X1 U11236 ( .A1(n10467), .A2(n10466), .ZN(n10468) );
  XOR2_X1 U11237 ( .A(n10593), .B(n10468), .Z(ADD_1071_U5) );
  XOR2_X1 U11238 ( .A(n10470), .B(n10469), .Z(ADD_1071_U54) );
  XOR2_X1 U11239 ( .A(n10472), .B(n10471), .Z(ADD_1071_U53) );
  XNOR2_X1 U11240 ( .A(n10474), .B(n10473), .ZN(ADD_1071_U52) );
  NOR2_X1 U11241 ( .A1(n10476), .A2(n10475), .ZN(n10477) );
  XOR2_X1 U11242 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n10477), .Z(ADD_1071_U51) );
  XOR2_X1 U11243 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10478), .Z(ADD_1071_U50) );
  XOR2_X1 U11244 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10479), .Z(ADD_1071_U49) );
  XOR2_X1 U11245 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10480), .Z(ADD_1071_U48) );
  XOR2_X1 U11246 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n10481), .Z(ADD_1071_U47) );
  XOR2_X1 U11247 ( .A(n10483), .B(n10482), .Z(ADD_1071_U63) );
  XOR2_X1 U11248 ( .A(n10485), .B(n10484), .Z(ADD_1071_U62) );
  XNOR2_X1 U11249 ( .A(n10487), .B(n10486), .ZN(ADD_1071_U61) );
  XNOR2_X1 U11250 ( .A(n10489), .B(n10488), .ZN(ADD_1071_U60) );
  XNOR2_X1 U11251 ( .A(n10491), .B(n10490), .ZN(ADD_1071_U59) );
  XNOR2_X1 U11252 ( .A(n10493), .B(n10492), .ZN(ADD_1071_U58) );
  XNOR2_X1 U11253 ( .A(n10495), .B(n10494), .ZN(ADD_1071_U57) );
  XNOR2_X1 U11254 ( .A(n10497), .B(n10496), .ZN(ADD_1071_U56) );
  NOR2_X1 U11255 ( .A1(n10499), .A2(n10498), .ZN(n10500) );
  XOR2_X1 U11256 ( .A(P1_ADDR_REG_18__SCAN_IN), .B(n10500), .Z(ADD_1071_U55)
         );
  INV_X1 U11257 ( .A(n10501), .ZN(n10508) );
  NAND2_X1 U11258 ( .A1(n10503), .A2(n10502), .ZN(n10506) );
  NAND2_X1 U11259 ( .A1(n10504), .A2(n10506), .ZN(n10505) );
  MUX2_X1 U11260 ( .A(n10506), .B(n10505), .S(P1_IR_REG_0__SCAN_IN), .Z(n10507) );
  NAND2_X1 U11261 ( .A1(n10508), .A2(n10507), .ZN(n10511) );
  AOI22_X1 U11262 ( .A1(n10550), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .ZN(n10510) );
  OAI21_X1 U11263 ( .B1(n10512), .B2(n10511), .A(n10510), .ZN(P1_U3241) );
  AOI22_X1 U11264 ( .A1(n10550), .A2(P1_ADDR_REG_6__SCAN_IN), .B1(n10513), 
        .B2(n10566), .ZN(n10524) );
  AOI211_X1 U11265 ( .C1(n10516), .C2(n10515), .A(n10514), .B(n10621), .ZN(
        n10517) );
  INV_X1 U11266 ( .A(n10517), .ZN(n10522) );
  OAI211_X1 U11267 ( .C1(n10520), .C2(n10519), .A(n10633), .B(n10518), .ZN(
        n10521) );
  NAND4_X1 U11268 ( .A1(n10524), .A2(n10523), .A3(n10522), .A4(n10521), .ZN(
        P1_U3247) );
  AOI22_X1 U11269 ( .A1(n10550), .A2(P1_ADDR_REG_9__SCAN_IN), .B1(n10525), 
        .B2(n10566), .ZN(n10536) );
  OAI21_X1 U11270 ( .B1(n10528), .B2(n10527), .A(n10526), .ZN(n10529) );
  NAND2_X1 U11271 ( .A1(n10529), .A2(n10573), .ZN(n10534) );
  OAI211_X1 U11272 ( .C1(n10532), .C2(n10531), .A(n10633), .B(n10530), .ZN(
        n10533) );
  NAND4_X1 U11273 ( .A1(n10536), .A2(n10535), .A3(n10534), .A4(n10533), .ZN(
        P1_U3250) );
  OAI21_X1 U11274 ( .B1(n10539), .B2(n10538), .A(n10537), .ZN(n10540) );
  AOI22_X1 U11275 ( .A1(n10540), .A2(n10573), .B1(n10550), .B2(
        P1_ADDR_REG_10__SCAN_IN), .ZN(n10548) );
  OAI211_X1 U11276 ( .C1(n10543), .C2(n10542), .A(n10541), .B(n10633), .ZN(
        n10546) );
  NAND2_X1 U11277 ( .A1(n10566), .A2(n10544), .ZN(n10545) );
  NAND4_X1 U11278 ( .A1(n10548), .A2(n10547), .A3(n10546), .A4(n10545), .ZN(
        P1_U3251) );
  AOI22_X1 U11279 ( .A1(n10550), .A2(P1_ADDR_REG_3__SCAN_IN), .B1(n10549), 
        .B2(n10566), .ZN(n10561) );
  INV_X1 U11280 ( .A(n10551), .ZN(n10552) );
  OAI211_X1 U11281 ( .C1(n10554), .C2(n10553), .A(n10573), .B(n10552), .ZN(
        n10559) );
  OAI211_X1 U11282 ( .C1(n10557), .C2(n10556), .A(n10633), .B(n10555), .ZN(
        n10558) );
  NAND4_X1 U11283 ( .A1(n10561), .A2(n10560), .A3(n10559), .A4(n10558), .ZN(
        P1_U3244) );
  NAND2_X1 U11284 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n10563) );
  AOI21_X1 U11285 ( .B1(n10564), .B2(n10563), .A(n10562), .ZN(n10572) );
  INV_X1 U11286 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10570) );
  NAND2_X1 U11287 ( .A1(n10566), .A2(n10565), .ZN(n10569) );
  NAND2_X1 U11288 ( .A1(P1_U3084), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n10568) );
  OAI211_X1 U11289 ( .C1(n10626), .C2(n10570), .A(n10569), .B(n10568), .ZN(
        n10571) );
  AOI21_X1 U11290 ( .B1(n10573), .B2(n10572), .A(n10571), .ZN(n10578) );
  OAI211_X1 U11291 ( .C1(n10576), .C2(n10575), .A(n10633), .B(n10574), .ZN(
        n10577) );
  NAND2_X1 U11292 ( .A1(n10578), .A2(n10577), .ZN(P1_U3242) );
  INV_X1 U11293 ( .A(n10579), .ZN(n10582) );
  INV_X1 U11294 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10581) );
  AOI22_X1 U11295 ( .A1(n10583), .A2(n10582), .B1(n10581), .B2(n10580), .ZN(
        P2_U3437) );
  AOI22_X1 U11296 ( .A1(n10584), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10615), .ZN(n10591) );
  AOI22_X1 U11297 ( .A1(n10606), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10590) );
  OAI21_X1 U11298 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(n10586), .A(n10585), .ZN(
        n10588) );
  NOR2_X1 U11299 ( .A1(n10607), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10587) );
  OAI21_X1 U11300 ( .B1(n10588), .B2(n10587), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n10589) );
  OAI211_X1 U11301 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n10591), .A(n10590), .B(
        n10589), .ZN(P2_U3245) );
  OAI22_X1 U11302 ( .A1(n10594), .A2(n10593), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10592), .ZN(n10599) );
  AOI211_X1 U11303 ( .C1(n10597), .C2(n10596), .A(n10595), .B(n10607), .ZN(
        n10598) );
  AOI211_X1 U11304 ( .C1(n10613), .C2(n10600), .A(n10599), .B(n10598), .ZN(
        n10605) );
  INV_X1 U11305 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10644) );
  NOR2_X1 U11306 ( .A1(n5421), .A2(n10644), .ZN(n10603) );
  OAI211_X1 U11307 ( .C1(n10603), .C2(n10602), .A(n10615), .B(n10601), .ZN(
        n10604) );
  NAND2_X1 U11308 ( .A1(n10605), .A2(n10604), .ZN(P2_U3246) );
  AOI22_X1 U11309 ( .A1(n10606), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n10620) );
  AOI211_X1 U11310 ( .C1(n10610), .C2(n10609), .A(n10608), .B(n10607), .ZN(
        n10611) );
  AOI21_X1 U11311 ( .B1(n10613), .B2(n10612), .A(n10611), .ZN(n10619) );
  OAI211_X1 U11312 ( .C1(n10617), .C2(n10616), .A(n10615), .B(n10614), .ZN(
        n10618) );
  NAND3_X1 U11313 ( .A1(n10620), .A2(n10619), .A3(n10618), .ZN(P2_U3247) );
  XNOR2_X1 U11314 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AOI211_X1 U11315 ( .C1(n10624), .C2(n10623), .A(n10622), .B(n10621), .ZN(
        n10630) );
  INV_X1 U11316 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10625) );
  OAI22_X1 U11317 ( .A1(n10628), .A2(n10627), .B1(n10626), .B2(n10625), .ZN(
        n10629) );
  NOR3_X1 U11318 ( .A1(n10631), .A2(n10630), .A3(n10629), .ZN(n10637) );
  OAI211_X1 U11319 ( .C1(n10635), .C2(n10634), .A(n10633), .B(n10632), .ZN(
        n10636) );
  OAI211_X1 U11320 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n10638), .A(n10637), .B(
        n10636), .ZN(P1_U3243) );
  OAI22_X1 U11321 ( .A1(n10641), .A2(n10841), .B1(n10640), .B2(n10639), .ZN(
        n10642) );
  NOR2_X1 U11322 ( .A1(n10643), .A2(n10642), .ZN(n10645) );
  AOI22_X1 U11323 ( .A1(n10870), .A2(n10645), .B1(n10644), .B2(n10868), .ZN(
        P2_U3520) );
  AOI22_X1 U11324 ( .A1(n10873), .A2(n10645), .B1(n5200), .B2(n10871), .ZN(
        P2_U3451) );
  INV_X1 U11325 ( .A(n10817), .ZN(n10766) );
  INV_X1 U11326 ( .A(n10646), .ZN(n10651) );
  OAI21_X1 U11327 ( .B1(n10648), .B2(n10888), .A(n10647), .ZN(n10650) );
  AOI211_X1 U11328 ( .C1(n10766), .C2(n10651), .A(n10650), .B(n10649), .ZN(
        n10652) );
  AOI22_X1 U11329 ( .A1(n10722), .A2(n10652), .B1(n5849), .B2(n10894), .ZN(
        P1_U3524) );
  AOI22_X1 U11330 ( .A1(n5045), .A2(n10652), .B1(n5368), .B2(n10896), .ZN(
        P1_U3457) );
  INV_X1 U11331 ( .A(n10653), .ZN(n10747) );
  NAND2_X1 U11332 ( .A1(n10654), .A2(n10792), .ZN(n10655) );
  OAI21_X1 U11333 ( .B1(n10656), .B2(n10860), .A(n10655), .ZN(n10658) );
  AOI211_X1 U11334 ( .C1(n10747), .C2(n10659), .A(n10658), .B(n10657), .ZN(
        n10661) );
  AOI22_X1 U11335 ( .A1(n10870), .A2(n10661), .B1(n10660), .B2(n10868), .ZN(
        P2_U3522) );
  AOI22_X1 U11336 ( .A1(n10873), .A2(n10661), .B1(n6518), .B2(n10871), .ZN(
        P2_U3457) );
  OAI22_X1 U11337 ( .A1(n10663), .A2(n10833), .B1(n10662), .B2(n10888), .ZN(
        n10665) );
  AOI211_X1 U11338 ( .C1(n10766), .C2(n10666), .A(n10665), .B(n10664), .ZN(
        n10669) );
  INV_X1 U11339 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10667) );
  AOI22_X1 U11340 ( .A1(n10722), .A2(n10669), .B1(n10667), .B2(n10894), .ZN(
        P1_U3526) );
  INV_X1 U11341 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10668) );
  AOI22_X1 U11342 ( .A1(n5045), .A2(n10669), .B1(n10668), .B2(n10896), .ZN(
        P1_U3463) );
  OAI22_X1 U11343 ( .A1(n10670), .A2(n10862), .B1(n5317), .B2(n10860), .ZN(
        n10672) );
  AOI211_X1 U11344 ( .C1(n10866), .C2(n10673), .A(n10672), .B(n10671), .ZN(
        n10675) );
  AOI22_X1 U11345 ( .A1(n10870), .A2(n10675), .B1(n10674), .B2(n10868), .ZN(
        P2_U3524) );
  AOI22_X1 U11346 ( .A1(n10873), .A2(n10675), .B1(n6720), .B2(n10871), .ZN(
        P2_U3463) );
  NOR2_X1 U11347 ( .A1(n10676), .A2(n10841), .ZN(n10682) );
  OAI22_X1 U11348 ( .A1(n10678), .A2(n10862), .B1(n10677), .B2(n10860), .ZN(
        n10680) );
  AOI211_X1 U11349 ( .C1(n10682), .C2(n10681), .A(n10680), .B(n10679), .ZN(
        n10683) );
  AOI22_X1 U11350 ( .A1(n10870), .A2(n10683), .B1(n6285), .B2(n10868), .ZN(
        P2_U3526) );
  AOI22_X1 U11351 ( .A1(n10873), .A2(n10683), .B1(n6954), .B2(n10871), .ZN(
        P2_U3469) );
  OAI21_X1 U11352 ( .B1(n10685), .B2(n10888), .A(n10684), .ZN(n10687) );
  AOI211_X1 U11353 ( .C1(n10766), .C2(n10688), .A(n10687), .B(n10686), .ZN(
        n10691) );
  INV_X1 U11354 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10689) );
  AOI22_X1 U11355 ( .A1(n10722), .A2(n10691), .B1(n10689), .B2(n10894), .ZN(
        P1_U3530) );
  INV_X1 U11356 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10690) );
  AOI22_X1 U11357 ( .A1(n5045), .A2(n10691), .B1(n10690), .B2(n10896), .ZN(
        P1_U3475) );
  OAI22_X1 U11358 ( .A1(n10693), .A2(n10862), .B1(n10692), .B2(n10860), .ZN(
        n10695) );
  AOI211_X1 U11359 ( .C1(n10866), .C2(n10696), .A(n10695), .B(n10694), .ZN(
        n10698) );
  AOI22_X1 U11360 ( .A1(n10870), .A2(n10698), .B1(n10697), .B2(n10868), .ZN(
        P2_U3527) );
  AOI22_X1 U11361 ( .A1(n10873), .A2(n10698), .B1(n7105), .B2(n10871), .ZN(
        P2_U3472) );
  NAND3_X1 U11362 ( .A1(n5624), .A2(n10699), .A3(n10866), .ZN(n10701) );
  OAI211_X1 U11363 ( .C1(n10702), .C2(n10860), .A(n10701), .B(n10700), .ZN(
        n10703) );
  NOR2_X1 U11364 ( .A1(n10704), .A2(n10703), .ZN(n10706) );
  AOI22_X1 U11365 ( .A1(n10870), .A2(n10706), .B1(n10705), .B2(n10868), .ZN(
        P2_U3528) );
  AOI22_X1 U11366 ( .A1(n10873), .A2(n10706), .B1(n7238), .B2(n10871), .ZN(
        P2_U3475) );
  XNOR2_X1 U11367 ( .A(n10707), .B(n10712), .ZN(n10719) );
  INV_X1 U11368 ( .A(n10719), .ZN(n10727) );
  INV_X1 U11369 ( .A(n10708), .ZN(n10711) );
  INV_X1 U11370 ( .A(n10709), .ZN(n10710) );
  OAI21_X1 U11371 ( .B1(n10730), .B2(n10711), .A(n10710), .ZN(n10725) );
  OAI22_X1 U11372 ( .A1(n10725), .A2(n10833), .B1(n10730), .B2(n10888), .ZN(
        n10720) );
  XNOR2_X1 U11373 ( .A(n10713), .B(n10712), .ZN(n10716) );
  OAI22_X1 U11374 ( .A1(n10756), .A2(n10753), .B1(n10714), .B2(n10755), .ZN(
        n10715) );
  AOI21_X1 U11375 ( .B1(n10716), .B2(n10758), .A(n10715), .ZN(n10717) );
  OAI21_X1 U11376 ( .B1(n10719), .B2(n10718), .A(n10717), .ZN(n10732) );
  AOI211_X1 U11377 ( .C1(n10766), .C2(n10727), .A(n10720), .B(n10732), .ZN(
        n10724) );
  AOI22_X1 U11378 ( .A1(n10722), .A2(n10724), .B1(n10721), .B2(n10894), .ZN(
        P1_U3532) );
  INV_X1 U11379 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10723) );
  AOI22_X1 U11380 ( .A1(n5045), .A2(n10724), .B1(n10723), .B2(n10896), .ZN(
        P1_U3481) );
  INV_X1 U11381 ( .A(n10725), .ZN(n10726) );
  AOI22_X1 U11382 ( .A1(n10727), .A2(n10773), .B1(n10772), .B2(n10726), .ZN(
        n10734) );
  AOI22_X1 U11383 ( .A1(n10778), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n10728), 
        .B2(n10776), .ZN(n10729) );
  OAI21_X1 U11384 ( .B1(n10730), .B2(n10780), .A(n10729), .ZN(n10731) );
  AOI21_X1 U11385 ( .B1(n10732), .B2(n10783), .A(n10731), .ZN(n10733) );
  NAND2_X1 U11386 ( .A1(n10734), .A2(n10733), .ZN(P1_U3282) );
  OAI22_X1 U11387 ( .A1(n10736), .A2(n10862), .B1(n10735), .B2(n10860), .ZN(
        n10738) );
  AOI211_X1 U11388 ( .C1(n10747), .C2(n10739), .A(n10738), .B(n10737), .ZN(
        n10740) );
  AOI22_X1 U11389 ( .A1(n10870), .A2(n10740), .B1(n6290), .B2(n10868), .ZN(
        P2_U3529) );
  AOI22_X1 U11390 ( .A1(n10873), .A2(n10740), .B1(n7246), .B2(n10871), .ZN(
        P2_U3478) );
  INV_X1 U11391 ( .A(n10741), .ZN(n10746) );
  OAI22_X1 U11392 ( .A1(n10743), .A2(n10862), .B1(n10742), .B2(n10860), .ZN(
        n10745) );
  AOI211_X1 U11393 ( .C1(n10747), .C2(n10746), .A(n10745), .B(n10744), .ZN(
        n10748) );
  AOI22_X1 U11394 ( .A1(n10870), .A2(n10748), .B1(n6397), .B2(n10868), .ZN(
        P2_U3530) );
  AOI22_X1 U11395 ( .A1(n10873), .A2(n10748), .B1(n7375), .B2(n10871), .ZN(
        P2_U3481) );
  XNOR2_X1 U11396 ( .A(n10749), .B(n10750), .ZN(n10774) );
  NAND2_X1 U11397 ( .A1(n10774), .A2(n10822), .ZN(n10761) );
  XNOR2_X1 U11398 ( .A(n10752), .B(n10751), .ZN(n10759) );
  OAI22_X1 U11399 ( .A1(n10756), .A2(n10755), .B1(n10754), .B2(n10753), .ZN(
        n10757) );
  AOI21_X1 U11400 ( .B1(n10759), .B2(n10758), .A(n10757), .ZN(n10760) );
  AND2_X1 U11401 ( .A1(n10761), .A2(n10760), .ZN(n10775) );
  OR2_X1 U11402 ( .A1(n10762), .A2(n10781), .ZN(n10763) );
  NAND2_X1 U11403 ( .A1(n10764), .A2(n10763), .ZN(n10770) );
  OAI22_X1 U11404 ( .A1(n10770), .A2(n10833), .B1(n10781), .B2(n10888), .ZN(
        n10765) );
  AOI21_X1 U11405 ( .B1(n10774), .B2(n10766), .A(n10765), .ZN(n10767) );
  AOI22_X1 U11406 ( .A1(n10722), .A2(n10769), .B1(n6100), .B2(n10894), .ZN(
        P1_U3534) );
  INV_X1 U11407 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10768) );
  AOI22_X1 U11408 ( .A1(n5045), .A2(n10769), .B1(n10768), .B2(n10896), .ZN(
        P1_U3487) );
  INV_X1 U11409 ( .A(n10770), .ZN(n10771) );
  AOI22_X1 U11410 ( .A1(n10774), .A2(n10773), .B1(n10772), .B2(n10771), .ZN(
        n10786) );
  INV_X1 U11411 ( .A(n10775), .ZN(n10784) );
  AOI22_X1 U11412 ( .A1(n10778), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n10777), 
        .B2(n10776), .ZN(n10779) );
  OAI21_X1 U11413 ( .B1(n10781), .B2(n10780), .A(n10779), .ZN(n10782) );
  AOI21_X1 U11414 ( .B1(n10784), .B2(n10783), .A(n10782), .ZN(n10785) );
  NAND2_X1 U11415 ( .A1(n10786), .A2(n10785), .ZN(P1_U3280) );
  OAI21_X1 U11416 ( .B1(n10789), .B2(n10788), .A(n10787), .ZN(n10790) );
  INV_X1 U11417 ( .A(n10790), .ZN(n10810) );
  OAI211_X1 U11418 ( .C1(n10793), .C2(n10794), .A(n10792), .B(n10791), .ZN(
        n10806) );
  OAI21_X1 U11419 ( .B1(n10794), .B2(n10860), .A(n10806), .ZN(n10799) );
  XNOR2_X1 U11420 ( .A(n7811), .B(n10795), .ZN(n10798) );
  OAI21_X1 U11421 ( .B1(n10798), .B2(n10797), .A(n10796), .ZN(n10807) );
  AOI211_X1 U11422 ( .C1(n10810), .C2(n10866), .A(n10799), .B(n10807), .ZN(
        n10800) );
  AOI22_X1 U11423 ( .A1(n10870), .A2(n10800), .B1(n6462), .B2(n10868), .ZN(
        P2_U3531) );
  AOI22_X1 U11424 ( .A1(n10873), .A2(n10800), .B1(n7420), .B2(n10871), .ZN(
        P2_U3484) );
  AOI22_X1 U11425 ( .A1(n10804), .A2(n10803), .B1(n10802), .B2(n10801), .ZN(
        n10805) );
  OAI21_X1 U11426 ( .B1(n10806), .B2(n5256), .A(n10805), .ZN(n10808) );
  AOI211_X1 U11427 ( .C1(n10810), .C2(n10809), .A(n10808), .B(n10807), .ZN(
        n10812) );
  AOI22_X1 U11428 ( .A1(n10813), .A2(n7421), .B1(n10812), .B2(n10811), .ZN(
        P2_U3285) );
  AOI21_X1 U11429 ( .B1(n10877), .B2(n10815), .A(n10814), .ZN(n10816) );
  OAI21_X1 U11430 ( .B1(n10818), .B2(n10817), .A(n10816), .ZN(n10820) );
  AOI211_X1 U11431 ( .C1(n10822), .C2(n10821), .A(n10820), .B(n10819), .ZN(
        n10824) );
  AOI22_X1 U11432 ( .A1(n10722), .A2(n10824), .B1(n6183), .B2(n10894), .ZN(
        P1_U3535) );
  INV_X1 U11433 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10823) );
  AOI22_X1 U11434 ( .A1(n5045), .A2(n10824), .B1(n10823), .B2(n10896), .ZN(
        P1_U3490) );
  OAI22_X1 U11435 ( .A1(n10826), .A2(n10862), .B1(n10825), .B2(n10860), .ZN(
        n10828) );
  AOI211_X1 U11436 ( .C1(n10866), .C2(n10829), .A(n10828), .B(n10827), .ZN(
        n10830) );
  AOI22_X1 U11437 ( .A1(n10870), .A2(n10830), .B1(n7058), .B2(n10868), .ZN(
        P2_U3532) );
  AOI22_X1 U11438 ( .A1(n10873), .A2(n10830), .B1(n7541), .B2(n10871), .ZN(
        P2_U3487) );
  INV_X1 U11439 ( .A(n10831), .ZN(n10892) );
  OAI22_X1 U11440 ( .A1(n10834), .A2(n10833), .B1(n10832), .B2(n10888), .ZN(
        n10836) );
  AOI211_X1 U11441 ( .C1(n10837), .C2(n10892), .A(n10836), .B(n10835), .ZN(
        n10840) );
  INV_X1 U11442 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10838) );
  AOI22_X1 U11443 ( .A1(n10722), .A2(n10840), .B1(n10838), .B2(n10894), .ZN(
        P1_U3536) );
  INV_X1 U11444 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10839) );
  AOI22_X1 U11445 ( .A1(n5045), .A2(n10840), .B1(n10839), .B2(n10896), .ZN(
        P1_U3493) );
  NOR2_X1 U11446 ( .A1(n10842), .A2(n10841), .ZN(n10848) );
  OAI22_X1 U11447 ( .A1(n10844), .A2(n10862), .B1(n10843), .B2(n10860), .ZN(
        n10845) );
  AOI211_X1 U11448 ( .C1(n10848), .C2(n10847), .A(n10846), .B(n10845), .ZN(
        n10850) );
  AOI22_X1 U11449 ( .A1(n10870), .A2(n10850), .B1(n10849), .B2(n10868), .ZN(
        P2_U3533) );
  AOI22_X1 U11450 ( .A1(n10873), .A2(n10850), .B1(n7566), .B2(n10871), .ZN(
        P2_U3490) );
  OAI211_X1 U11451 ( .C1(n10853), .C2(n10888), .A(n10852), .B(n10851), .ZN(
        n10854) );
  AOI21_X1 U11452 ( .B1(n10892), .B2(n10855), .A(n10854), .ZN(n10858) );
  AOI22_X1 U11453 ( .A1(n10722), .A2(n10858), .B1(n10856), .B2(n10894), .ZN(
        P1_U3537) );
  INV_X1 U11454 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10857) );
  AOI22_X1 U11455 ( .A1(n5045), .A2(n10858), .B1(n10857), .B2(n10896), .ZN(
        P1_U3496) );
  INV_X1 U11456 ( .A(n10859), .ZN(n10867) );
  OAI22_X1 U11457 ( .A1(n10863), .A2(n10862), .B1(n10861), .B2(n10860), .ZN(
        n10864) );
  AOI211_X1 U11458 ( .C1(n10867), .C2(n10866), .A(n10865), .B(n10864), .ZN(
        n10872) );
  AOI22_X1 U11459 ( .A1(n10870), .A2(n10872), .B1(n10869), .B2(n10868), .ZN(
        P2_U3534) );
  AOI22_X1 U11460 ( .A1(n10873), .A2(n10872), .B1(n7804), .B2(n10871), .ZN(
        P2_U3493) );
  NAND3_X1 U11461 ( .A1(n10875), .A2(n10874), .A3(n10892), .ZN(n10882) );
  AOI22_X1 U11462 ( .A1(n10879), .A2(n10878), .B1(n10877), .B2(n10876), .ZN(
        n10880) );
  AOI22_X1 U11463 ( .A1(n10722), .A2(n10885), .B1(n10883), .B2(n10894), .ZN(
        P1_U3538) );
  INV_X1 U11464 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10884) );
  AOI22_X1 U11465 ( .A1(n5045), .A2(n10885), .B1(n10884), .B2(n10896), .ZN(
        P1_U3499) );
  INV_X1 U11466 ( .A(n10886), .ZN(n10889) );
  OAI21_X1 U11467 ( .B1(n10889), .B2(n10888), .A(n10887), .ZN(n10891) );
  AOI211_X1 U11468 ( .C1(n10893), .C2(n10892), .A(n10891), .B(n10890), .ZN(
        n10898) );
  AOI22_X1 U11469 ( .A1(n10722), .A2(n10898), .B1(n10895), .B2(n10894), .ZN(
        P1_U3539) );
  INV_X1 U11470 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10897) );
  AOI22_X1 U11471 ( .A1(n5045), .A2(n10898), .B1(n10897), .B2(n10896), .ZN(
        P1_U3502) );
  XNOR2_X1 U11472 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  CLKBUF_X2 U5146 ( .A(n6718), .Z(n8171) );
  CLKBUF_X1 U5279 ( .A(n6516), .Z(n8191) );
endmodule

