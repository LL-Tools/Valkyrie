

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, keyinput58, 
        keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, keyinput52, 
        keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, keyinput46, 
        keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, keyinput40, 
        keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, keyinput34, 
        keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, keyinput28, 
        keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, keyinput22, 
        keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, keyinput16, 
        keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, 
        keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, 
        keyinput3, keyinput2, keyinput1, keyinput0 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput63,
         keyinput62, keyinput61, keyinput60, keyinput59, keyinput58,
         keyinput57, keyinput56, keyinput55, keyinput54, keyinput53,
         keyinput52, keyinput51, keyinput50, keyinput49, keyinput48,
         keyinput47, keyinput46, keyinput45, keyinput44, keyinput43,
         keyinput42, keyinput41, keyinput40, keyinput39, keyinput38,
         keyinput37, keyinput36, keyinput35, keyinput34, keyinput33,
         keyinput32, keyinput31, keyinput30, keyinput29, keyinput28,
         keyinput27, keyinput26, keyinput25, keyinput24, keyinput23,
         keyinput22, keyinput21, keyinput20, keyinput19, keyinput18,
         keyinput17, keyinput16, keyinput15, keyinput14, keyinput13,
         keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, keyinput7,
         keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, keyinput1,
         keyinput0;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180;

  OAI21_X1 U7170 ( .B1(n12038), .B2(n9253), .A(n9576), .ZN(n14058) );
  NOR2_X1 U7171 ( .A1(n7898), .A2(n7897), .ZN(n7915) );
  INV_X1 U7172 ( .A(n8738), .ZN(n8828) );
  CLKBUF_X1 U7173 ( .A(n10629), .Z(n6434) );
  INV_X1 U7174 ( .A(n9695), .ZN(n9672) );
  INV_X1 U7175 ( .A(n9253), .ZN(n9715) );
  NAND2_X1 U7176 ( .A1(n7395), .A2(n13422), .ZN(n13427) );
  INV_X2 U7177 ( .A(n8096), .ZN(n8061) );
  CLKBUF_X3 U7178 ( .A(n12152), .Z(n6435) );
  AND2_X1 U7179 ( .A1(n8408), .A2(n8407), .ZN(n8454) );
  AND2_X1 U7180 ( .A1(n6592), .A2(n6591), .ZN(n9155) );
  AOI21_X1 U7181 ( .B1(n12627), .B2(n9839), .A(n9838), .ZN(n12608) );
  NAND2_X1 U7182 ( .A1(n15062), .A2(n15085), .ZN(n10559) );
  INV_X1 U7183 ( .A(n12152), .ZN(n10900) );
  INV_X2 U7184 ( .A(n10629), .ZN(n10625) );
  AND2_X1 U7185 ( .A1(n12152), .A2(n13958), .ZN(n10634) );
  NAND2_X1 U7186 ( .A1(n11085), .A2(n9720), .ZN(n10591) );
  INV_X1 U7187 ( .A(n12284), .ZN(n11386) );
  XNOR2_X1 U7188 ( .A(n9147), .B(n9148), .ZN(n15010) );
  OR2_X1 U7189 ( .A1(n12525), .A2(n12524), .ZN(n6995) );
  BUF_X1 U7190 ( .A(n8448), .Z(n8738) );
  BUF_X1 U7191 ( .A(n8449), .Z(n8829) );
  INV_X1 U7192 ( .A(n9799), .ZN(n8438) );
  INV_X1 U7193 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8479) );
  INV_X1 U7194 ( .A(n11598), .ZN(n8293) );
  INV_X1 U7195 ( .A(n10712), .ZN(n11018) );
  NAND2_X1 U7196 ( .A1(n13187), .A2(n9942), .ZN(n13175) );
  INV_X2 U7197 ( .A(n10634), .ZN(n12159) );
  NAND2_X1 U7199 ( .A1(n9465), .A2(n9464), .ZN(n13946) );
  INV_X1 U7200 ( .A(n13398), .ZN(n13162) );
  NAND2_X1 U7201 ( .A1(n10293), .A2(n11532), .ZN(n7799) );
  NAND2_X1 U7202 ( .A1(n7537), .A2(n7536), .ZN(n11168) );
  INV_X1 U7203 ( .A(n14898), .ZN(n14896) );
  AND4_X1 U7204 ( .A1(n8371), .A2(n8370), .A3(n8369), .A4(n14207), .ZN(n6422)
         );
  AND2_X1 U7205 ( .A1(n10596), .A2(n10591), .ZN(n12152) );
  NAND2_X1 U7206 ( .A1(n7325), .A2(n10638), .ZN(n10718) );
  OR2_X1 U7207 ( .A1(n7388), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n7661) );
  NAND2_X2 U7208 ( .A1(n11477), .A2(n11476), .ZN(n11585) );
  AOI21_X2 U7209 ( .B1(n12582), .B2(n8844), .A(n8971), .ZN(n12563) );
  INV_X4 U7210 ( .A(n10694), .ZN(n10967) );
  AND3_X4 U7211 ( .A1(n6833), .A2(n7380), .A3(n7379), .ZN(n10694) );
  NAND2_X2 U7212 ( .A1(n9038), .A2(n7332), .ZN(n9040) );
  NAND2_X2 U7213 ( .A1(n6951), .A2(n10899), .ZN(n10946) );
  NAND2_X2 U7214 ( .A1(n10734), .A2(n10733), .ZN(n6951) );
  NOR2_X2 U7215 ( .A1(n14936), .A2(n9135), .ZN(n9137) );
  OR2_X1 U7216 ( .A1(n7467), .A2(n7466), .ZN(n10712) );
  AND2_X4 U7217 ( .A1(n6589), .A2(n6956), .ZN(n12130) );
  XNOR2_X2 U7218 ( .A(n9043), .B(n9136), .ZN(n10789) );
  CLKBUF_X1 U7219 ( .A(n9693), .Z(n6423) );
  NAND2_X2 U7221 ( .A1(n14270), .A2(n9182), .ZN(n9693) );
  XNOR2_X2 U7222 ( .A(n9151), .B(n9150), .ZN(n14439) );
  BUF_X4 U7223 ( .A(n8454), .Z(n6426) );
  XNOR2_X2 U7224 ( .A(n9140), .B(n14959), .ZN(n14955) );
  NOR2_X2 U7225 ( .A1(n10508), .A2(n15093), .ZN(n10511) );
  NOR2_X2 U7226 ( .A1(n10988), .A2(n10987), .ZN(n10986) );
  XNOR2_X2 U7227 ( .A(n7384), .B(n7383), .ZN(n11598) );
  XNOR2_X2 U7228 ( .A(n8271), .B(n10967), .ZN(n9915) );
  AOI21_X2 U7229 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n10993), .A(n10986), .ZN(
        n9046) );
  XNOR2_X2 U7230 ( .A(n9056), .B(n12516), .ZN(n12508) );
  AND3_X4 U7231 ( .A1(n7008), .A2(n7009), .A3(n6573), .ZN(n9056) );
  INV_X2 U7232 ( .A(n7479), .ZN(n7438) );
  XNOR2_X2 U7233 ( .A(n9050), .B(n9148), .ZN(n15003) );
  AOI21_X4 U7234 ( .B1(n6599), .B2(n6598), .A(n6597), .ZN(n9050) );
  AOI21_X2 U7235 ( .B1(P3_REG1_REG_8__SCAN_IN), .B2(n10993), .A(n10994), .ZN(
        n9140) );
  NAND2_X1 U7236 ( .A1(n13471), .A2(n12140), .ZN(n13535) );
  AND2_X1 U7237 ( .A1(n13124), .A2(n13389), .ZN(n13114) );
  NOR2_X2 U7238 ( .A1(n6768), .A2(n13162), .ZN(n13158) );
  AND2_X1 U7239 ( .A1(n7876), .A2(n7875), .ZN(n13174) );
  OAI21_X1 U7240 ( .B1(n14991), .B2(n7069), .A(n7068), .ZN(n12462) );
  CLKBUF_X2 U7241 ( .A(n6434), .Z(n12162) );
  CLKBUF_X2 U7242 ( .A(n6434), .Z(n12071) );
  NOR2_X2 U7243 ( .A1(n15077), .A2(n10582), .ZN(n10566) );
  INV_X1 U7244 ( .A(n8453), .ZN(n8832) );
  CLKBUF_X2 U7245 ( .A(P2_U3947), .Z(n6427) );
  BUF_X1 U7246 ( .A(n10594), .Z(n11060) );
  INV_X4 U7247 ( .A(n13083), .ZN(n7779) );
  CLKBUF_X2 U7248 ( .A(n9247), .Z(n9716) );
  NAND2_X1 U7250 ( .A1(n7392), .A2(n12239), .ZN(n9954) );
  NAND2_X1 U7251 ( .A1(n14861), .A2(n11815), .ZN(n11535) );
  INV_X8 U7252 ( .A(n7438), .ZN(n10049) );
  INV_X8 U7253 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n7677) );
  OR2_X1 U7254 ( .A1(n7082), .A2(n6744), .ZN(n6742) );
  AOI211_X1 U7255 ( .C1(n14623), .C2(n14027), .A(n13789), .B(n13788), .ZN(
        n13790) );
  AND2_X1 U7256 ( .A1(n14025), .A2(n7331), .ZN(n6632) );
  OAI21_X1 U7257 ( .B1(n13314), .B2(n13362), .A(n13312), .ZN(n6610) );
  AND2_X1 U7258 ( .A1(n13330), .A2(n13329), .ZN(n13396) );
  OR2_X1 U7259 ( .A1(n13796), .A2(n6630), .ZN(n6624) );
  AND2_X1 U7260 ( .A1(n13154), .A2(n13153), .ZN(n13329) );
  NAND2_X1 U7261 ( .A1(n13797), .A2(n6699), .ZN(n13796) );
  OR2_X1 U7262 ( .A1(n8159), .A2(n8160), .ZN(n8161) );
  AND2_X1 U7263 ( .A1(n6625), .A2(n14729), .ZN(n6622) );
  NAND2_X1 U7264 ( .A1(n13499), .A2(n12131), .ZN(n13470) );
  AND2_X1 U7265 ( .A1(n13810), .A2(n13729), .ZN(n13797) );
  OR2_X1 U7266 ( .A1(n13151), .A2(n13279), .ZN(n13154) );
  NAND2_X1 U7267 ( .A1(n12623), .A2(n12626), .ZN(n12625) );
  NAND2_X1 U7268 ( .A1(n8748), .A2(n8852), .ZN(n12623) );
  AND2_X1 U7269 ( .A1(n13142), .A2(n13129), .ZN(n13124) );
  OAI21_X2 U7270 ( .B1(n13175), .B2(n7059), .A(n9944), .ZN(n13156) );
  NAND2_X1 U7271 ( .A1(n12916), .A2(n7845), .ZN(n7865) );
  AND2_X1 U7272 ( .A1(n13158), .A2(n13394), .ZN(n13142) );
  NAND2_X1 U7273 ( .A1(n12942), .A2(n7232), .ZN(n12916) );
  INV_X1 U7274 ( .A(n13174), .ZN(n6769) );
  NAND2_X1 U7275 ( .A1(n12690), .A2(n9834), .ZN(n12674) );
  OAI21_X1 U7276 ( .B1(n7900), .B2(n7899), .A(n7915), .ZN(n12019) );
  NAND2_X1 U7277 ( .A1(n6882), .A2(n6879), .ZN(n12690) );
  AND2_X1 U7278 ( .A1(n7721), .A2(n7739), .ZN(n7231) );
  NAND2_X1 U7279 ( .A1(n7895), .A2(n7873), .ZN(n7894) );
  OAI21_X1 U7280 ( .B1(n14439), .B2(n7072), .A(n7071), .ZN(n12498) );
  AND2_X1 U7281 ( .A1(n12917), .A2(n7825), .ZN(n7232) );
  NAND2_X1 U7282 ( .A1(n11886), .A2(n11885), .ZN(n11924) );
  NAND2_X1 U7283 ( .A1(n11787), .A2(n6458), .ZN(n11878) );
  AND2_X1 U7284 ( .A1(n9103), .A2(n9150), .ZN(n9104) );
  NAND2_X1 U7285 ( .A1(n7849), .A2(n7848), .ZN(n7851) );
  NAND2_X1 U7286 ( .A1(n7850), .A2(SI_22_), .ZN(n7869) );
  NAND2_X1 U7287 ( .A1(n11585), .A2(n11584), .ZN(n11586) );
  NAND2_X1 U7288 ( .A1(n9448), .A2(n9447), .ZN(n14522) );
  NAND2_X1 U7289 ( .A1(n7847), .A2(n7846), .ZN(n7850) );
  NAND2_X1 U7290 ( .A1(n7831), .A2(n7830), .ZN(n7847) );
  NAND2_X1 U7291 ( .A1(n9824), .A2(n9823), .ZN(n14451) );
  NAND2_X1 U7292 ( .A1(n9423), .A2(n9422), .ZN(n11934) );
  NAND2_X1 U7293 ( .A1(n7665), .A2(n7664), .ZN(n11666) );
  NAND2_X1 U7294 ( .A1(n9476), .A2(n9475), .ZN(n14232) );
  OR2_X1 U7295 ( .A1(n7807), .A2(n11210), .ZN(n7826) );
  NAND2_X1 U7296 ( .A1(n7643), .A2(n7642), .ZN(n11643) );
  XNOR2_X1 U7297 ( .A(n9144), .B(n9143), .ZN(n14991) );
  NAND2_X1 U7298 ( .A1(n11158), .A2(n11157), .ZN(n11156) );
  OAI21_X1 U7299 ( .B1(n14955), .B2(n7066), .A(n7065), .ZN(n14974) );
  OR2_X1 U7300 ( .A1(n11239), .A2(n14881), .ZN(n11331) );
  NOR2_X1 U7301 ( .A1(n13540), .A2(n13991), .ZN(n13551) );
  NAND2_X1 U7302 ( .A1(n6690), .A2(n7511), .ZN(n11096) );
  NAND2_X1 U7303 ( .A1(n6715), .A2(n6717), .ZN(n7553) );
  CLKBUF_X1 U7304 ( .A(n10634), .Z(n6594) );
  INV_X1 U7305 ( .A(n11389), .ZN(n12448) );
  INV_X1 U7306 ( .A(n11176), .ZN(n12450) );
  INV_X2 U7307 ( .A(n15094), .ZN(n15071) );
  NAND2_X1 U7308 ( .A1(n9255), .A2(n9254), .ZN(n14668) );
  NAND4_X1 U7309 ( .A1(n8425), .A2(n8424), .A3(n8423), .A4(n8422), .ZN(n15077)
         );
  BUF_X1 U7310 ( .A(n8271), .Z(n6429) );
  NAND2_X1 U7311 ( .A1(n9704), .A2(n9213), .ZN(n9310) );
  AND3_X1 U7312 ( .A1(n8468), .A2(n8467), .A3(n8466), .ZN(n10845) );
  CLKBUF_X1 U7313 ( .A(n7535), .Z(n8236) );
  INV_X4 U7314 ( .A(n7987), .ZN(n7918) );
  NAND4_X1 U7315 ( .A1(n9246), .A2(n9245), .A3(n9244), .A4(n9243), .ZN(n13571)
         );
  AND4_X1 U7316 ( .A1(n9189), .A2(n9188), .A3(n9187), .A4(n9186), .ZN(n10594)
         );
  AOI22_X1 U7317 ( .A1(n9506), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n10162), .B2(
        n13607), .ZN(n9255) );
  INV_X2 U7318 ( .A(n9558), .ZN(n10162) );
  NAND2_X1 U7319 ( .A1(n9719), .A2(n11268), .ZN(n10315) );
  NAND2_X2 U7320 ( .A1(n9558), .A2(n7438), .ZN(n9253) );
  NAND2_X2 U7321 ( .A1(n12029), .A2(n6431), .ZN(n9799) );
  INV_X1 U7322 ( .A(n13427), .ZN(n7399) );
  NAND2_X1 U7323 ( .A1(n6812), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6811) );
  NAND2_X2 U7324 ( .A1(n6604), .A2(n6602), .ZN(n12882) );
  NAND2_X2 U7325 ( .A1(n9784), .A2(n9783), .ZN(n9558) );
  NAND2_X1 U7326 ( .A1(n9210), .A2(n9209), .ZN(n11268) );
  XNOR2_X1 U7327 ( .A(n9205), .B(P1_IR_REG_20__SCAN_IN), .ZN(n11257) );
  XNOR2_X1 U7328 ( .A(n9203), .B(n9206), .ZN(n11650) );
  AND2_X1 U7329 ( .A1(n8022), .A2(n11532), .ZN(n14861) );
  MUX2_X1 U7330 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7393), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n7395) );
  MUX2_X1 U7331 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7359), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n6855) );
  NAND2_X1 U7332 ( .A1(n9194), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9196) );
  INV_X1 U7333 ( .A(n8382), .ZN(n6428) );
  MUX2_X1 U7334 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7360), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n6854) );
  OR2_X1 U7335 ( .A1(n10511), .A2(n9032), .ZN(n10447) );
  OAI21_X1 U7336 ( .B1(n7385), .B2(n7229), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n7360) );
  NAND2_X2 U7337 ( .A1(n10049), .A2(P3_U3151), .ZN(n12040) );
  AND2_X1 U7338 ( .A1(n7287), .A2(n6994), .ZN(n6993) );
  AND2_X1 U7339 ( .A1(n9199), .A2(n9200), .ZN(n7287) );
  AND2_X1 U7340 ( .A1(n7389), .A2(n7352), .ZN(n7353) );
  NAND2_X1 U7341 ( .A1(n8436), .A2(n8435), .ZN(n10066) );
  NOR2_X1 U7342 ( .A1(n6866), .A2(n6867), .ZN(n6863) );
  AND3_X1 U7343 ( .A1(n8375), .A2(n7201), .A3(n8445), .ZN(n6864) );
  AND4_X1 U7344 ( .A1(n7348), .A2(n7347), .A3(n7531), .A4(n7346), .ZN(n7349)
         );
  AND2_X1 U7345 ( .A1(n9172), .A2(n9171), .ZN(n9200) );
  AND2_X1 U7346 ( .A1(n7386), .A2(n7228), .ZN(n7226) );
  AND3_X1 U7347 ( .A1(n7351), .A2(n7350), .A3(n7679), .ZN(n7389) );
  AND2_X1 U7348 ( .A1(n9170), .A2(n9169), .ZN(n9199) );
  INV_X1 U7349 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n7509) );
  INV_X1 U7350 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n7991) );
  INV_X1 U7351 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9195) );
  INV_X1 U7352 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7459) );
  NOR2_X1 U7353 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n9172) );
  NOR2_X1 U7354 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n9171) );
  INV_X4 U7355 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7356 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n7614) );
  NOR3_X1 U7357 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .A3(
        P1_IR_REG_24__SCAN_IN), .ZN(n9176) );
  NOR3_X1 U7358 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .A3(
        P2_IR_REG_13__SCAN_IN), .ZN(n7352) );
  NOR2_X1 U7359 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n9166) );
  INV_X1 U7360 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9284) );
  NOR2_X1 U7361 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n9165) );
  NOR2_X1 U7362 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n9169) );
  NOR2_X1 U7363 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n9170) );
  INV_X4 U7364 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7365 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n8405) );
  INV_X4 U7366 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7367 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n12243) );
  INV_X1 U7368 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7365) );
  NOR2_X1 U7369 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n8372) );
  NOR2_X1 U7370 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n8370) );
  NOR2_X1 U7371 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n8369) );
  NOR2_X1 U7372 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n7201) );
  NOR2_X2 U7373 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n8445) );
  NOR2_X1 U7374 ( .A1(P3_IR_REG_11__SCAN_IN), .A2(P3_IR_REG_12__SCAN_IN), .ZN(
        n8375) );
  NOR2_X1 U7375 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_13__SCAN_IN), .ZN(
        n8373) );
  NOR2_X1 U7376 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n8374) );
  INV_X2 U7377 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7294) );
  OAI21_X1 U7378 ( .B1(n13301), .B2(n14478), .A(n10029), .ZN(n10030) );
  NAND4_X1 U7379 ( .A1(n7402), .A2(n7400), .A3(n7401), .A4(n7403), .ZN(n8271)
         );
  NAND2_X1 U7380 ( .A1(n6604), .A2(n6602), .ZN(n6430) );
  NAND2_X1 U7381 ( .A1(n6604), .A2(n6602), .ZN(n6431) );
  NAND2_X2 U7382 ( .A1(n10640), .A2(n10641), .ZN(n10734) );
  INV_X2 U7383 ( .A(n11141), .ZN(n10631) );
  XNOR2_X2 U7384 ( .A(n10630), .B(n11141), .ZN(n11131) );
  NAND2_X2 U7385 ( .A1(n11769), .A2(n11768), .ZN(n11787) );
  NAND2_X2 U7386 ( .A1(n10906), .A2(n10905), .ZN(n10945) );
  AND2_X4 U7387 ( .A1(n8408), .A2(n12042), .ZN(n8455) );
  AOI21_X2 U7388 ( .B1(P3_REG1_REG_14__SCAN_IN), .B2(n12474), .A(n12469), .ZN(
        n9151) );
  NAND2_X1 U7389 ( .A1(n8032), .A2(n12024), .ZN(n6432) );
  NAND2_X1 U7390 ( .A1(n8032), .A2(n12024), .ZN(n6433) );
  AND2_X2 U7391 ( .A1(n12033), .A2(n7399), .ZN(n8204) );
  INV_X4 U7392 ( .A(n8204), .ZN(n7452) );
  NAND2_X2 U7393 ( .A1(n11586), .A2(n11587), .ZN(n11769) );
  NAND2_X2 U7394 ( .A1(n6855), .A2(n7394), .ZN(n8032) );
  OAI22_X2 U7395 ( .A1(n13136), .A2(n9945), .B1(n10001), .B2(n13006), .ZN(
        n13130) );
  OAI21_X1 U7396 ( .B1(n13130), .B2(n7037), .A(n7034), .ZN(n13091) );
  NAND2_X2 U7397 ( .A1(n13535), .A2(n13536), .ZN(n13534) );
  OAI21_X2 U7398 ( .B1(n13234), .B2(n6860), .A(n6858), .ZN(n13180) );
  INV_X2 U7399 ( .A(n10630), .ZN(n9224) );
  NAND4_X2 U7400 ( .A1(n9217), .A2(n9216), .A3(n9215), .A4(n9214), .ZN(n10630)
         );
  AOI21_X2 U7401 ( .B1(P3_REG1_REG_12__SCAN_IN), .B2(n10100), .A(n12462), .ZN(
        n9147) );
  NAND2_X2 U7402 ( .A1(n13482), .A2(n13483), .ZN(n13481) );
  XNOR2_X2 U7403 ( .A(n9779), .B(P1_IR_REG_24__SCAN_IN), .ZN(n10102) );
  XNOR2_X2 U7404 ( .A(n9777), .B(P1_IR_REG_25__SCAN_IN), .ZN(n10103) );
  INV_X1 U7405 ( .A(n8457), .ZN(n8504) );
  NOR2_X1 U7406 ( .A1(n12838), .A2(n12595), .ZN(n9840) );
  NAND2_X1 U7407 ( .A1(n12735), .A2(n9832), .ZN(n6882) );
  NAND2_X1 U7408 ( .A1(n6869), .A2(n6868), .ZN(n12627) );
  AOI21_X1 U7409 ( .B1(n6871), .B2(n6873), .A(n6496), .ZN(n6868) );
  NAND2_X1 U7410 ( .A1(n13964), .A2(n6641), .ZN(n6640) );
  NOR2_X1 U7411 ( .A1(n7309), .A2(n6642), .ZN(n6641) );
  INV_X1 U7412 ( .A(n13714), .ZN(n6642) );
  NAND2_X1 U7413 ( .A1(n13928), .A2(n13940), .ZN(n7309) );
  NAND2_X1 U7414 ( .A1(n6750), .A2(n6751), .ZN(n8188) );
  NAND2_X1 U7415 ( .A1(n7935), .A2(n6752), .ZN(n6750) );
  NAND2_X1 U7416 ( .A1(n9799), .A2(n10049), .ZN(n8449) );
  INV_X1 U7417 ( .A(n6426), .ZN(n8835) );
  XNOR2_X1 U7418 ( .A(n12602), .B(n12583), .ZN(n12599) );
  AOI21_X1 U7419 ( .B1(n6784), .B2(n6787), .A(n6783), .ZN(n6782) );
  INV_X1 U7420 ( .A(n7182), .ZN(n7180) );
  NOR2_X1 U7421 ( .A1(n7108), .A2(n8093), .ZN(n7109) );
  NAND2_X1 U7422 ( .A1(n8113), .A2(n7091), .ZN(n7090) );
  AOI21_X1 U7423 ( .B1(n7103), .B2(n7101), .A(n7100), .ZN(n7099) );
  INV_X1 U7424 ( .A(n6736), .ZN(n6733) );
  AOI21_X1 U7425 ( .B1(n6752), .B2(n7934), .A(n6564), .ZN(n6751) );
  INV_X1 U7426 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9768) );
  NOR2_X1 U7427 ( .A1(n8985), .A2(n8840), .ZN(n6807) );
  NAND2_X1 U7428 ( .A1(n10446), .A2(n9034), .ZN(n9035) );
  NAND2_X1 U7429 ( .A1(n12591), .A2(n12596), .ZN(n9842) );
  AND2_X1 U7430 ( .A1(n12591), .A2(n12570), .ZN(n8971) );
  NOR2_X1 U7431 ( .A1(n12599), .A2(n6898), .ZN(n6897) );
  INV_X1 U7432 ( .A(n6900), .ZN(n6898) );
  OR2_X1 U7433 ( .A1(n12771), .A2(n12643), .ZN(n8963) );
  INV_X1 U7434 ( .A(n9836), .ZN(n6877) );
  NOR2_X1 U7435 ( .A1(n7329), .A2(n6549), .ZN(n6881) );
  OR2_X1 U7436 ( .A1(n12862), .A2(n12724), .ZN(n8932) );
  INV_X1 U7437 ( .A(n8899), .ZN(n6791) );
  AND2_X1 U7438 ( .A1(n8561), .A2(n8560), .ZN(n8905) );
  INV_X1 U7439 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8379) );
  OR2_X1 U7440 ( .A1(n8345), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8347) );
  AND2_X1 U7441 ( .A1(n8695), .A2(n8338), .ZN(n7164) );
  NAND2_X1 U7442 ( .A1(n8590), .A2(n8324), .ZN(n8325) );
  OR2_X1 U7443 ( .A1(n8541), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8543) );
  INV_X1 U7444 ( .A(n8314), .ZN(n7134) );
  OR2_X1 U7445 ( .A1(n8267), .A2(n12889), .ZN(n10005) );
  NAND2_X1 U7446 ( .A1(n6515), .A2(n9997), .ZN(n6860) );
  NAND2_X1 U7447 ( .A1(n6470), .A2(n9940), .ZN(n7030) );
  NAND2_X1 U7448 ( .A1(n13236), .A2(n13235), .ZN(n13234) );
  NAND2_X1 U7449 ( .A1(n7049), .A2(n13258), .ZN(n7048) );
  INV_X1 U7450 ( .A(n7050), .ZN(n7049) );
  INV_X1 U7451 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7228) );
  NAND2_X1 U7452 ( .A1(n6702), .A2(n7254), .ZN(n6701) );
  NOR2_X1 U7453 ( .A1(n6943), .A2(n13727), .ZN(n6942) );
  INV_X1 U7454 ( .A(n6945), .ZN(n6943) );
  AOI21_X1 U7455 ( .B1(n13928), .B2(n7311), .A(n6494), .ZN(n7310) );
  INV_X1 U7456 ( .A(n13716), .ZN(n7311) );
  INV_X1 U7457 ( .A(n11650), .ZN(n11085) );
  OAI21_X1 U7458 ( .B1(n7746), .B2(n6724), .A(n6721), .ZN(n7807) );
  AOI21_X1 U7459 ( .B1(n7236), .B2(n6723), .A(n6722), .ZN(n6721) );
  NAND2_X1 U7460 ( .A1(n7236), .A2(n6725), .ZN(n6724) );
  NOR2_X1 U7461 ( .A1(n7804), .A2(SI_19_), .ZN(n6722) );
  NAND2_X1 U7462 ( .A1(n7762), .A2(n7238), .ZN(n7237) );
  XNOR2_X1 U7463 ( .A(n7804), .B(SI_19_), .ZN(n7805) );
  NAND2_X1 U7464 ( .A1(n7743), .A2(n7742), .ZN(n7746) );
  OAI21_X1 U7465 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(n14291), .A(n14290), .ZN(
        n14292) );
  OAI22_X1 U7466 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(n14988), .B1(n14312), 
        .B2(n14363), .ZN(n14366) );
  NOR2_X1 U7467 ( .A1(n6445), .A2(n6655), .ZN(n6654) );
  INV_X1 U7468 ( .A(n6663), .ZN(n6655) );
  INV_X1 U7469 ( .A(n7178), .ZN(n7177) );
  NAND2_X1 U7470 ( .A1(n15077), .A2(n10818), .ZN(n15073) );
  NAND2_X1 U7471 ( .A1(n12380), .A2(n6552), .ZN(n12334) );
  AND2_X1 U7472 ( .A1(n14973), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7021) );
  OR2_X1 U7473 ( .A1(n12442), .A2(n12558), .ZN(n7340) );
  XNOR2_X1 U7474 ( .A(n12289), .B(n12422), .ZN(n12568) );
  OR2_X1 U7475 ( .A1(n8790), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8804) );
  AND2_X1 U7476 ( .A1(n8770), .A2(n8769), .ZN(n12595) );
  NAND2_X1 U7477 ( .A1(n12793), .A2(n12407), .ZN(n9834) );
  AOI21_X1 U7478 ( .B1(n6779), .B2(n6780), .A(n6776), .ZN(n6775) );
  INV_X1 U7479 ( .A(n8895), .ZN(n6776) );
  INV_X1 U7480 ( .A(n11339), .ZN(n9884) );
  INV_X1 U7481 ( .A(n8829), .ZN(n8699) );
  INV_X1 U7482 ( .A(n7335), .ZN(n6815) );
  OAI21_X1 U7483 ( .B1(n8761), .B2(n12016), .A(n8347), .ZN(n8772) );
  INV_X1 U7484 ( .A(n8736), .ZN(n7147) );
  AOI21_X1 U7485 ( .B1(n8736), .B2(n7146), .A(n7145), .ZN(n7144) );
  INV_X1 U7486 ( .A(n8343), .ZN(n7145) );
  INV_X1 U7487 ( .A(n8340), .ZN(n7146) );
  AND2_X1 U7488 ( .A1(n7197), .A2(n8376), .ZN(n7196) );
  AND2_X1 U7489 ( .A1(n7201), .A2(n7198), .ZN(n7197) );
  NAND2_X1 U7490 ( .A1(n8720), .A2(n8721), .ZN(n8725) );
  NAND2_X1 U7491 ( .A1(n8633), .A2(n8329), .ZN(n8649) );
  NAND2_X1 U7492 ( .A1(n8649), .A2(n8648), .ZN(n8647) );
  NAND2_X1 U7493 ( .A1(n7126), .A2(n7124), .ZN(n8633) );
  AND2_X1 U7494 ( .A1(n7123), .A2(n7122), .ZN(n7124) );
  AND2_X1 U7495 ( .A1(n7125), .A2(n6546), .ZN(n7122) );
  INV_X1 U7496 ( .A(n8630), .ZN(n7125) );
  OAI21_X1 U7497 ( .B1(n8558), .B2(n8557), .A(n8319), .ZN(n8565) );
  INV_X1 U7498 ( .A(n8312), .ZN(n7138) );
  NAND2_X1 U7499 ( .A1(n7152), .A2(n7150), .ZN(n7156) );
  NOR2_X1 U7500 ( .A1(n8307), .A2(n7151), .ZN(n7150) );
  INV_X1 U7501 ( .A(n7522), .ZN(n11042) );
  AND2_X1 U7502 ( .A1(n7611), .A2(n7590), .ZN(n7230) );
  AOI21_X1 U7503 ( .B1(n13115), .B2(n7966), .A(n7965), .ZN(n12985) );
  OAI21_X1 U7504 ( .B1(n11749), .B2(n9932), .A(n9933), .ZN(n14482) );
  INV_X1 U7505 ( .A(n6835), .ZN(n6834) );
  NAND2_X1 U7506 ( .A1(n10011), .A2(n10010), .ZN(n14475) );
  NAND3_X1 U7507 ( .A1(n7851), .A2(n7869), .A3(n7852), .ZN(n7872) );
  INV_X1 U7508 ( .A(n7854), .ZN(n7852) );
  OAI211_X1 U7509 ( .C1(n10602), .C2(n10596), .A(n10601), .B(n10600), .ZN(
        n10637) );
  OAI211_X1 U7510 ( .C1(n13577), .C2(n10324), .A(n10325), .B(n6621), .ZN(
        n13592) );
  NAND2_X1 U7511 ( .A1(n13577), .A2(n10324), .ZN(n6621) );
  OR2_X1 U7512 ( .A1(n9407), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n9420) );
  NOR3_X1 U7513 ( .A1(n13798), .A2(n6442), .A3(n14028), .ZN(n6820) );
  OR2_X1 U7514 ( .A1(n13800), .A2(n14034), .ZN(n13798) );
  NAND2_X1 U7515 ( .A1(n6636), .A2(n6637), .ZN(n6635) );
  NAND2_X1 U7516 ( .A1(n9632), .A2(n9631), .ZN(n13817) );
  AND2_X1 U7517 ( .A1(n14045), .A2(n13748), .ZN(n7254) );
  OR2_X1 U7518 ( .A1(n13856), .A2(n6946), .ZN(n6944) );
  INV_X1 U7519 ( .A(n6947), .ZN(n6946) );
  NOR2_X1 U7520 ( .A1(n13876), .A2(n14058), .ZN(n6831) );
  AND2_X1 U7521 ( .A1(n13897), .A2(n13718), .ZN(n7316) );
  OR2_X1 U7522 ( .A1(n13946), .A2(n13955), .ZN(n13741) );
  NAND2_X1 U7523 ( .A1(n6643), .A2(n13710), .ZN(n6644) );
  AND2_X1 U7524 ( .A1(n7299), .A2(n13710), .ZN(n6646) );
  INV_X1 U7525 ( .A(n13565), .ZN(n11582) );
  NAND2_X1 U7526 ( .A1(n6931), .A2(n11438), .ZN(n6933) );
  INV_X1 U7527 ( .A(n6939), .ZN(n6931) );
  NAND2_X1 U7528 ( .A1(n9558), .A2(n10049), .ZN(n9247) );
  NAND2_X1 U7529 ( .A1(n10594), .A2(n11125), .ZN(n11071) );
  AOI21_X1 U7530 ( .B1(n10310), .B2(n10308), .A(n10307), .ZN(n10748) );
  NAND2_X1 U7531 ( .A1(n8230), .A2(n8197), .ZN(n8234) );
  NOR2_X1 U7532 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n7318) );
  NAND2_X1 U7533 ( .A1(n14353), .A2(n14352), .ZN(n14354) );
  OAI21_X1 U7534 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n14307), .A(n14306), .ZN(
        n14356) );
  AOI21_X1 U7535 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n14309), .A(n14308), .ZN(
        n14358) );
  NOR2_X1 U7536 ( .A1(n14357), .A2(n14356), .ZN(n14308) );
  NAND2_X1 U7537 ( .A1(n6666), .A2(n6665), .ZN(n7041) );
  NAND2_X1 U7538 ( .A1(n14364), .A2(n14365), .ZN(n6665) );
  INV_X1 U7539 ( .A(n14552), .ZN(n6666) );
  INV_X1 U7540 ( .A(n12629), .ZN(n12654) );
  NAND2_X1 U7541 ( .A1(n8778), .A2(n8777), .ZN(n12602) );
  INV_X1 U7542 ( .A(n12838), .ZN(n12377) );
  NAND2_X1 U7543 ( .A1(n8785), .A2(n8784), .ZN(n12583) );
  NOR2_X1 U7544 ( .A1(n12535), .A2(n7075), .ZN(n7074) );
  AND2_X1 U7545 ( .A1(n14960), .A2(n12536), .ZN(n7075) );
  AOI21_X1 U7546 ( .B1(n9116), .B2(n14963), .A(n9115), .ZN(n9120) );
  XNOR2_X1 U7547 ( .A(n6608), .B(n6607), .ZN(n9116) );
  INV_X1 U7548 ( .A(n9111), .ZN(n6607) );
  NAND2_X1 U7549 ( .A1(n8264), .A2(n7342), .ZN(n8265) );
  OR2_X1 U7550 ( .A1(n14402), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n6670) );
  XNOR2_X1 U7551 ( .A(n7041), .B(n14369), .ZN(n7040) );
  AND2_X1 U7552 ( .A1(n9240), .A2(n11064), .ZN(n9242) );
  NAND2_X1 U7553 ( .A1(n9225), .A2(n10631), .ZN(n9226) );
  NAND2_X1 U7554 ( .A1(n9224), .A2(n9223), .ZN(n9227) );
  INV_X1 U7555 ( .A(n8055), .ZN(n8058) );
  MUX2_X1 U7556 ( .A(n13028), .B(n10712), .S(n8074), .Z(n8072) );
  NAND2_X1 U7557 ( .A1(n7280), .A2(n9411), .ZN(n7279) );
  INV_X1 U7558 ( .A(n9461), .ZN(n7266) );
  NAND2_X1 U7559 ( .A1(n8093), .A2(n7108), .ZN(n7107) );
  OAI21_X1 U7560 ( .B1(n9523), .B2(n7261), .A(n9522), .ZN(n9534) );
  NAND2_X1 U7561 ( .A1(n9520), .A2(n9519), .ZN(n9523) );
  OR2_X1 U7562 ( .A1(n9546), .A2(n9548), .ZN(n7289) );
  NAND2_X1 U7563 ( .A1(n8102), .A2(n8104), .ZN(n7084) );
  NOR2_X1 U7564 ( .A1(n7102), .A2(n8121), .ZN(n7103) );
  NAND2_X1 U7565 ( .A1(n8121), .A2(n7102), .ZN(n7101) );
  OAI21_X1 U7566 ( .B1(n8114), .B2(n6501), .A(n6576), .ZN(n8119) );
  NOR2_X1 U7567 ( .A1(n8118), .A2(n6577), .ZN(n6576) );
  NOR2_X1 U7568 ( .A1(n7118), .A2(n8154), .ZN(n7119) );
  NAND2_X1 U7569 ( .A1(n7118), .A2(n8154), .ZN(n7117) );
  OR2_X1 U7570 ( .A1(n9719), .A2(n11268), .ZN(n9211) );
  NAND2_X1 U7571 ( .A1(n7639), .A2(n7638), .ZN(n6728) );
  NAND2_X1 U7572 ( .A1(n8978), .A2(n8977), .ZN(n7176) );
  OAI21_X1 U7573 ( .B1(n8771), .B2(n6802), .A(n12599), .ZN(n6801) );
  NAND2_X1 U7574 ( .A1(n12451), .A2(n10772), .ZN(n8874) );
  AOI21_X1 U7575 ( .B1(n7028), .B2(n7027), .A(n7026), .ZN(n7025) );
  INV_X1 U7576 ( .A(n7031), .ZN(n7027) );
  INV_X1 U7577 ( .A(n13203), .ZN(n7026) );
  INV_X1 U7578 ( .A(n9682), .ZN(n7275) );
  INV_X1 U7579 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7364) );
  INV_X1 U7580 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7362) );
  OAI21_X1 U7581 ( .B1(n11738), .B2(n7212), .A(n7210), .ZN(n11940) );
  OR2_X1 U7582 ( .A1(n6472), .A2(n7211), .ZN(n7210) );
  NAND2_X1 U7583 ( .A1(n7213), .A2(n11938), .ZN(n7212) );
  INV_X1 U7584 ( .A(n11938), .ZN(n7211) );
  NAND2_X1 U7585 ( .A1(n9906), .A2(n8980), .ZN(n6808) );
  INV_X1 U7586 ( .A(n7002), .ZN(n6999) );
  AOI21_X1 U7587 ( .B1(n8479), .B2(P3_IR_REG_2__SCAN_IN), .A(n7005), .ZN(n7001) );
  NAND2_X1 U7588 ( .A1(n6596), .A2(n14923), .ZN(n7017) );
  NAND3_X1 U7589 ( .A1(n6441), .A2(n9131), .A3(P3_REG1_REG_3__SCAN_IN), .ZN(
        n7064) );
  NAND2_X1 U7590 ( .A1(n7017), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7015) );
  AND2_X1 U7591 ( .A1(n10468), .A2(n7080), .ZN(n9133) );
  NAND2_X1 U7592 ( .A1(n10478), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7080) );
  AND2_X1 U7593 ( .A1(n10035), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n9135) );
  AND2_X1 U7594 ( .A1(n12478), .A2(n12477), .ZN(n12475) );
  NAND2_X1 U7595 ( .A1(n12497), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n6591) );
  INV_X1 U7596 ( .A(n12498), .ZN(n6592) );
  NOR2_X1 U7597 ( .A1(n12511), .A2(n9108), .ZN(n9109) );
  OR2_X1 U7598 ( .A1(n9910), .A2(n12327), .ZN(n8980) );
  NOR2_X1 U7599 ( .A1(n6797), .A2(n6796), .ZN(n6795) );
  INV_X1 U7600 ( .A(n8954), .ZN(n6796) );
  NOR2_X1 U7601 ( .A1(n8718), .A2(n6798), .ZN(n6797) );
  INV_X1 U7602 ( .A(n8951), .ZN(n6798) );
  OR2_X1 U7603 ( .A1(n8728), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8741) );
  INV_X1 U7604 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n12354) );
  NAND2_X1 U7605 ( .A1(n14457), .A2(n6892), .ZN(n6891) );
  INV_X1 U7606 ( .A(n9887), .ZN(n9883) );
  NAND2_X1 U7607 ( .A1(n10564), .A2(n10559), .ZN(n15052) );
  INV_X1 U7608 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9017) );
  AND2_X1 U7609 ( .A1(n8846), .A2(n7183), .ZN(n7182) );
  INV_X1 U7610 ( .A(n8664), .ZN(n7159) );
  INV_X1 U7611 ( .A(n8331), .ZN(n7158) );
  NOR2_X1 U7612 ( .A1(n7137), .A2(n8314), .ZN(n7132) );
  NAND2_X1 U7613 ( .A1(n8435), .A2(n7006), .ZN(n7003) );
  AND2_X1 U7614 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n7007), .ZN(n7006) );
  NAND2_X1 U7615 ( .A1(n8172), .A2(n6491), .ZN(n6578) );
  NAND2_X1 U7616 ( .A1(n6438), .A2(n6451), .ZN(n7120) );
  NAND2_X1 U7617 ( .A1(n8173), .A2(n8174), .ZN(n7121) );
  OR2_X1 U7618 ( .A1(n8251), .A2(n8250), .ZN(n8252) );
  AOI211_X1 U7619 ( .C1(n8225), .C2(n8223), .A(n8250), .B(n8224), .ZN(n8254)
         );
  INV_X1 U7620 ( .A(n10004), .ZN(n6848) );
  NOR2_X1 U7621 ( .A1(n6449), .A2(n7330), .ZN(n6851) );
  NAND2_X1 U7622 ( .A1(n13155), .A2(n6464), .ZN(n6852) );
  OR2_X1 U7623 ( .A1(n6769), .A2(n13008), .ZN(n9944) );
  NAND2_X1 U7624 ( .A1(n13192), .A2(n6767), .ZN(n6766) );
  AND2_X1 U7625 ( .A1(n10019), .A2(n6773), .ZN(n6772) );
  NOR2_X1 U7626 ( .A1(n11643), .A2(n12208), .ZN(n6773) );
  INV_X1 U7627 ( .A(n9971), .ZN(n6837) );
  AND2_X1 U7628 ( .A1(n11231), .A2(n9923), .ZN(n7060) );
  AND2_X1 U7629 ( .A1(n8293), .A2(n11532), .ZN(n9955) );
  NAND2_X1 U7630 ( .A1(n6584), .A2(n13181), .ZN(n13187) );
  INV_X1 U7631 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n7993) );
  INV_X1 U7632 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n7348) );
  NOR2_X1 U7633 ( .A1(n11832), .A2(n11709), .ZN(n7299) );
  NAND2_X1 U7634 ( .A1(n6932), .A2(n6473), .ZN(n6939) );
  NAND2_X1 U7635 ( .A1(n11302), .A2(n11301), .ZN(n6941) );
  NAND2_X1 U7636 ( .A1(n6473), .A2(n11301), .ZN(n6938) );
  INV_X1 U7637 ( .A(n11075), .ZN(n6930) );
  NAND2_X1 U7638 ( .A1(n10631), .A2(n10630), .ZN(n6916) );
  INV_X1 U7639 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n14287) );
  NAND2_X1 U7640 ( .A1(n11184), .A2(n11066), .ZN(n7305) );
  OAI21_X1 U7641 ( .B1(n7915), .B2(n6749), .A(n6565), .ZN(n8210) );
  INV_X1 U7642 ( .A(n6752), .ZN(n6749) );
  NAND2_X1 U7643 ( .A1(n6752), .A2(n6748), .ZN(n6747) );
  NAND2_X1 U7644 ( .A1(n7915), .A2(n7914), .ZN(n7935) );
  AOI21_X1 U7645 ( .B1(n6440), .B2(n7239), .A(n6511), .ZN(n7236) );
  INV_X1 U7646 ( .A(n7762), .ZN(n7239) );
  OR2_X1 U7647 ( .A1(n9491), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n9493) );
  NAND2_X1 U7648 ( .A1(n7240), .A2(n7241), .ZN(n7743) );
  AOI21_X1 U7649 ( .B1(n7243), .B2(n7245), .A(n6510), .ZN(n7241) );
  NOR2_X1 U7650 ( .A1(n7702), .A2(n7247), .ZN(n7246) );
  INV_X1 U7651 ( .A(n7674), .ZN(n7247) );
  AND2_X1 U7652 ( .A1(n7658), .A2(n6474), .ZN(n6736) );
  NAND2_X1 U7653 ( .A1(n6737), .A2(n7638), .ZN(n7656) );
  NAND2_X1 U7654 ( .A1(n7613), .A2(n7612), .ZN(n7640) );
  INV_X1 U7655 ( .A(n7549), .ZN(n6718) );
  OAI21_X1 U7656 ( .B1(n7479), .B2(n7367), .A(n7366), .ZN(n7368) );
  XNOR2_X1 U7657 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n14329) );
  NAND2_X1 U7658 ( .A1(n14294), .A2(n14295), .ZN(n14325) );
  NOR2_X1 U7659 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n6660), .ZN(n6657) );
  NOR2_X1 U7660 ( .A1(n7192), .A2(n7190), .ZN(n7189) );
  AOI21_X1 U7661 ( .B1(n7194), .B2(n7193), .A(n12407), .ZN(n7192) );
  INV_X1 U7662 ( .A(n12408), .ZN(n7194) );
  AND2_X1 U7663 ( .A1(n12362), .A2(n12264), .ZN(n7193) );
  AND2_X1 U7664 ( .A1(n7191), .A2(n12408), .ZN(n7190) );
  NAND2_X1 U7665 ( .A1(n12362), .A2(n12264), .ZN(n7191) );
  OR2_X1 U7666 ( .A1(n8804), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8817) );
  OR2_X1 U7667 ( .A1(n8597), .A2(n8387), .ZN(n8610) );
  AOI21_X1 U7668 ( .B1(n12399), .B2(n12654), .A(n12304), .ZN(n12369) );
  AND2_X1 U7669 ( .A1(n11010), .A2(n11008), .ZN(n7186) );
  NAND2_X1 U7670 ( .A1(n7214), .A2(n7213), .ZN(n11803) );
  NAND2_X1 U7671 ( .A1(n10565), .A2(n10562), .ZN(n7178) );
  INV_X1 U7672 ( .A(n11980), .ZN(n7203) );
  AND2_X1 U7673 ( .A1(n12292), .A2(n7206), .ZN(n7205) );
  NAND2_X1 U7674 ( .A1(n7208), .A2(n7207), .ZN(n7206) );
  INV_X1 U7675 ( .A(n12430), .ZN(n12256) );
  AND2_X1 U7676 ( .A1(n8838), .A2(n8420), .ZN(n9901) );
  AND4_X1 U7677 ( .A1(n8473), .A2(n8472), .A3(n8471), .A4(n8470), .ZN(n11176)
         );
  AND2_X1 U7678 ( .A1(n8407), .A2(n8406), .ZN(n8457) );
  OAI21_X1 U7679 ( .B1(n10066), .B2(n9031), .A(n9030), .ZN(n10508) );
  NOR2_X1 U7680 ( .A1(n10820), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9031) );
  AND2_X1 U7681 ( .A1(n9035), .A2(n10054), .ZN(n9036) );
  OR2_X1 U7682 ( .A1(n14929), .A2(n14928), .ZN(n6997) );
  AND2_X1 U7683 ( .A1(n6997), .A2(n6996), .ZN(n9043) );
  NAND2_X1 U7684 ( .A1(n10035), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n6996) );
  INV_X1 U7685 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11945) );
  AND2_X1 U7686 ( .A1(n7020), .A2(n6519), .ZN(n12454) );
  AOI21_X1 U7687 ( .B1(P3_REG2_REG_14__SCAN_IN), .B2(n12474), .A(n9052), .ZN(
        n9053) );
  NAND2_X1 U7688 ( .A1(n9100), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7019) );
  NAND2_X1 U7689 ( .A1(n9051), .A2(n9100), .ZN(n7018) );
  XNOR2_X1 U7690 ( .A(n9155), .B(n12516), .ZN(n12518) );
  NOR2_X1 U7691 ( .A1(n12513), .A2(n12512), .ZN(n12511) );
  NAND2_X1 U7692 ( .A1(n8980), .A2(n8979), .ZN(n9907) );
  OAI21_X1 U7693 ( .B1(n6896), .B2(n6895), .A(n6505), .ZN(n6894) );
  INV_X1 U7694 ( .A(n9842), .ZN(n6895) );
  AOI21_X1 U7695 ( .B1(n12568), .B2(n12565), .A(n12564), .ZN(n12574) );
  OR2_X1 U7696 ( .A1(n8764), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8779) );
  OR2_X1 U7697 ( .A1(n12377), .A2(n12630), .ZN(n6900) );
  AND2_X1 U7698 ( .A1(n6899), .A2(n6897), .ZN(n12597) );
  INV_X1 U7699 ( .A(n12583), .ZN(n12614) );
  INV_X1 U7700 ( .A(n12663), .ZN(n12642) );
  NAND2_X1 U7701 ( .A1(n6516), .A2(n6877), .ZN(n6874) );
  AND2_X1 U7702 ( .A1(n8852), .A2(n8851), .ZN(n12645) );
  OR2_X1 U7703 ( .A1(n8702), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8713) );
  NAND2_X1 U7704 ( .A1(n8719), .A2(n8718), .ZN(n12665) );
  NOR2_X1 U7705 ( .A1(n6880), .A2(n12687), .ZN(n6879) );
  INV_X1 U7706 ( .A(n6881), .ZN(n6880) );
  OR2_X1 U7707 ( .A1(n8670), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8687) );
  OR2_X1 U7708 ( .A1(n8640), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8657) );
  OAI21_X1 U7709 ( .B1(n11865), .B2(n8616), .A(n8921), .ZN(n11915) );
  AND2_X1 U7710 ( .A1(n8918), .A2(n8917), .ZN(n11818) );
  AOI21_X1 U7711 ( .B1(n6790), .B2(n6786), .A(n6785), .ZN(n6784) );
  INV_X1 U7712 ( .A(n8904), .ZN(n6785) );
  AND2_X1 U7713 ( .A1(n8911), .A2(n8910), .ZN(n14455) );
  NAND2_X1 U7714 ( .A1(n9818), .A2(n9817), .ZN(n11313) );
  NAND2_X1 U7715 ( .A1(n8550), .A2(n8899), .ZN(n15038) );
  AND3_X1 U7716 ( .A1(n8532), .A2(n8531), .A3(n8530), .ZN(n9814) );
  AND4_X1 U7717 ( .A1(n8540), .A2(n8539), .A3(n8538), .A4(n8537), .ZN(n11566)
         );
  AND4_X1 U7718 ( .A1(n8510), .A2(n8509), .A3(n8508), .A4(n8507), .ZN(n11389)
         );
  NAND2_X1 U7719 ( .A1(n11026), .A2(n9812), .ZN(n11197) );
  AND2_X1 U7720 ( .A1(n8888), .A2(n8884), .ZN(n11030) );
  AND3_X1 U7721 ( .A1(n8485), .A2(n8484), .A3(n8483), .ZN(n11005) );
  INV_X1 U7722 ( .A(n15061), .ZN(n15076) );
  INV_X1 U7723 ( .A(n12736), .ZN(n15074) );
  INV_X1 U7724 ( .A(n11211), .ZN(n9886) );
  NAND2_X1 U7725 ( .A1(n8712), .A2(n8711), .ZN(n12784) );
  NAND2_X1 U7726 ( .A1(n8701), .A2(n8700), .ZN(n12788) );
  OR2_X1 U7727 ( .A1(n15083), .A2(n15143), .ZN(n15099) );
  OR2_X1 U7728 ( .A1(n9880), .A2(n9869), .ZN(n10570) );
  AND2_X1 U7729 ( .A1(n10537), .A2(n10542), .ZN(n10573) );
  INV_X1 U7730 ( .A(n15079), .ZN(n15059) );
  INV_X1 U7731 ( .A(n11955), .ZN(n9851) );
  AND2_X1 U7732 ( .A1(n9061), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10542) );
  AND2_X1 U7733 ( .A1(n8381), .A2(n6810), .ZN(n6809) );
  INV_X1 U7734 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n6810) );
  NAND2_X1 U7735 ( .A1(n8775), .A2(n8350), .ZN(n8787) );
  NAND2_X1 U7736 ( .A1(n8347), .A2(n8346), .ZN(n8761) );
  AND2_X1 U7737 ( .A1(n8343), .A2(n8342), .ZN(n8736) );
  NAND2_X1 U7738 ( .A1(n7163), .A2(n7162), .ZN(n8720) );
  NAND2_X1 U7739 ( .A1(n6562), .A2(n8338), .ZN(n7162) );
  NAND2_X1 U7740 ( .A1(n8696), .A2(n8695), .ZN(n8694) );
  NAND2_X1 U7741 ( .A1(n8682), .A2(n8335), .ZN(n8696) );
  NAND2_X1 U7742 ( .A1(n8326), .A2(n7128), .ZN(n7123) );
  NOR2_X1 U7743 ( .A1(n8327), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7128) );
  NAND2_X1 U7744 ( .A1(n7129), .A2(n8604), .ZN(n7126) );
  AND2_X1 U7745 ( .A1(n8326), .A2(n8617), .ZN(n7129) );
  NAND2_X1 U7746 ( .A1(n8325), .A2(n10443), .ZN(n8326) );
  OAI21_X1 U7747 ( .B1(n8325), .B2(n10443), .A(n8326), .ZN(n8604) );
  NAND2_X1 U7748 ( .A1(n7130), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8606) );
  INV_X1 U7749 ( .A(n8604), .ZN(n7130) );
  AND2_X1 U7750 ( .A1(n8324), .A2(n8323), .ZN(n8587) );
  NAND2_X1 U7751 ( .A1(n8322), .A2(n6460), .ZN(n7161) );
  OR2_X1 U7752 ( .A1(n8543), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n8566) );
  OAI21_X1 U7753 ( .B1(n8546), .B2(n8317), .A(n8316), .ZN(n8558) );
  INV_X1 U7754 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8513) );
  AOI21_X1 U7755 ( .B1(n7137), .B2(n8494), .A(n6455), .ZN(n7135) );
  XNOR2_X1 U7756 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n8516) );
  NAND2_X1 U7757 ( .A1(n8493), .A2(n8311), .ZN(n8496) );
  NAND2_X1 U7758 ( .A1(n8477), .A2(n8309), .ZN(n8493) );
  NAND2_X1 U7759 ( .A1(n7156), .A2(n7148), .ZN(n8477) );
  AND2_X1 U7760 ( .A1(n7155), .A2(n8306), .ZN(n7148) );
  INV_X1 U7761 ( .A(n8474), .ZN(n7155) );
  NOR2_X1 U7762 ( .A1(n10081), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7151) );
  NAND2_X1 U7763 ( .A1(n8304), .A2(n7153), .ZN(n7152) );
  NOR2_X1 U7764 ( .A1(n8305), .A2(n7154), .ZN(n7153) );
  INV_X1 U7765 ( .A(n8303), .ZN(n7154) );
  AOI21_X1 U7766 ( .B1(n6675), .B2(n6680), .A(n6674), .ZN(n6673) );
  INV_X1 U7767 ( .A(n7951), .ZN(n6674) );
  INV_X1 U7768 ( .A(n7761), .ZN(n6689) );
  NAND2_X1 U7769 ( .A1(n10764), .A2(n7524), .ZN(n7225) );
  AOI21_X1 U7770 ( .B1(n12955), .B2(n12954), .A(n7866), .ZN(n7887) );
  NAND2_X1 U7771 ( .A1(n12902), .A2(n6486), .ZN(n12942) );
  XNOR2_X1 U7772 ( .A(n11096), .B(n7918), .ZN(n7522) );
  NAND2_X1 U7773 ( .A1(n6677), .A2(n6675), .ZN(n12983) );
  NAND2_X1 U7774 ( .A1(n6682), .A2(n7913), .ZN(n6678) );
  AND2_X1 U7775 ( .A1(n7985), .A2(n7984), .ZN(n12889) );
  AND4_X1 U7776 ( .A1(n7756), .A2(n7755), .A3(n7754), .A4(n7753), .ZN(n12968)
         );
  OR2_X1 U7777 ( .A1(n8205), .A2(n7405), .ZN(n7407) );
  NAND2_X1 U7778 ( .A1(n9948), .A2(n9947), .ZN(n7037) );
  INV_X1 U7779 ( .A(n7035), .ZN(n7034) );
  OAI22_X1 U7780 ( .A1(n13109), .A2(n7036), .B1(n12985), .B2(n13389), .ZN(
        n7035) );
  AOI22_X2 U7781 ( .A1(n13166), .A2(n10000), .B1(n6769), .B2(n12959), .ZN(
        n13149) );
  NOR2_X1 U7782 ( .A1(n9941), .A2(n7032), .ZN(n7031) );
  INV_X1 U7783 ( .A(n9940), .ZN(n7032) );
  NAND2_X1 U7784 ( .A1(n6593), .A2(n6469), .ZN(n13211) );
  NAND2_X1 U7786 ( .A1(n13250), .A2(n9939), .ZN(n13226) );
  AOI21_X1 U7787 ( .B1(n7051), .B2(n11902), .A(n6488), .ZN(n7050) );
  AND2_X1 U7788 ( .A1(n13277), .A2(n9936), .ZN(n7051) );
  NAND2_X1 U7789 ( .A1(n9985), .A2(n14480), .ZN(n6841) );
  NAND2_X1 U7790 ( .A1(n9987), .A2(n9986), .ZN(n6840) );
  NAND3_X1 U7791 ( .A1(n6841), .A2(n6840), .A3(n11902), .ZN(n11896) );
  NAND2_X1 U7792 ( .A1(n7061), .A2(n9931), .ZN(n11749) );
  AND2_X1 U7793 ( .A1(n11620), .A2(n9979), .ZN(n6856) );
  NAND2_X1 U7794 ( .A1(n9968), .A2(n9967), .ZN(n10975) );
  NOR2_X1 U7795 ( .A1(n13030), .A2(n10018), .ZN(n10484) );
  OR2_X1 U7796 ( .A1(n11535), .A2(n8293), .ZN(n10287) );
  NAND2_X1 U7797 ( .A1(n7938), .A2(n7937), .ZN(n13318) );
  OR2_X1 U7798 ( .A1(n11649), .A2(n8235), .ZN(n7834) );
  AND2_X1 U7799 ( .A1(n8000), .A2(n13434), .ZN(n14870) );
  OR2_X1 U7800 ( .A1(n8006), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n7998) );
  AND2_X1 U7801 ( .A1(n7382), .A2(n7383), .ZN(n7992) );
  NOR2_X1 U7802 ( .A1(n7385), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n7382) );
  INV_X1 U7803 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7383) );
  NAND2_X1 U7804 ( .A1(n7354), .A2(n7353), .ZN(n7385) );
  NAND2_X1 U7805 ( .A1(n6964), .A2(n6962), .ZN(n6961) );
  INV_X1 U7806 ( .A(n6965), .ZN(n6962) );
  INV_X1 U7807 ( .A(n12110), .ZN(n6958) );
  INV_X1 U7808 ( .A(n12111), .ZN(n6959) );
  NAND2_X1 U7809 ( .A1(n6964), .A2(n12111), .ZN(n6960) );
  AOI21_X1 U7810 ( .B1(n13444), .B2(n12149), .A(n6976), .ZN(n6975) );
  INV_X1 U7811 ( .A(n12158), .ZN(n6976) );
  NOR2_X1 U7812 ( .A1(n13462), .A2(n6966), .ZN(n6965) );
  INV_X1 U7813 ( .A(n6968), .ZN(n6966) );
  NAND2_X1 U7814 ( .A1(n6980), .A2(n6444), .ZN(n6977) );
  NAND2_X1 U7815 ( .A1(n10627), .A2(n10626), .ZN(n10628) );
  INV_X1 U7816 ( .A(n9621), .ZN(n9697) );
  AND4_X1 U7817 ( .A1(n9456), .A2(n9455), .A3(n9454), .A4(n9453), .ZN(n12051)
         );
  AND4_X1 U7818 ( .A1(n9272), .A2(n9271), .A3(n9270), .A4(n9269), .ZN(n11077)
         );
  AND2_X1 U7819 ( .A1(n10163), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10033) );
  NAND2_X1 U7820 ( .A1(n13591), .A2(n13592), .ZN(n10326) );
  OR2_X1 U7821 ( .A1(n11608), .A2(n11609), .ZN(n6616) );
  AND2_X1 U7822 ( .A1(n13779), .A2(n14020), .ZN(n13756) );
  NAND2_X1 U7823 ( .A1(n6944), .A2(n6477), .ZN(n6695) );
  INV_X1 U7824 ( .A(n6697), .ZN(n6696) );
  XOR2_X1 U7825 ( .A(n13773), .B(n13758), .Z(n13754) );
  NOR2_X1 U7826 ( .A1(n13784), .A2(n7314), .ZN(n7313) );
  INV_X1 U7827 ( .A(n13730), .ZN(n7314) );
  INV_X1 U7828 ( .A(n13811), .ZN(n6704) );
  INV_X1 U7829 ( .A(n6944), .ZN(n6700) );
  AOI21_X1 U7830 ( .B1(n6947), .B2(n13863), .A(n6504), .ZN(n6945) );
  NAND2_X1 U7831 ( .A1(n13724), .A2(n13723), .ZN(n13848) );
  NAND2_X1 U7832 ( .A1(n6831), .A2(n6830), .ZN(n13843) );
  AND2_X1 U7833 ( .A1(n13851), .A2(n6479), .ZN(n6947) );
  NAND2_X1 U7834 ( .A1(n13856), .A2(n13855), .ZN(n6948) );
  OAI22_X1 U7835 ( .A1(n13871), .A2(n13873), .B1(n13745), .B2(n14066), .ZN(
        n13856) );
  NAND2_X1 U7836 ( .A1(n6950), .A2(n6949), .ZN(n13901) );
  AND2_X1 U7837 ( .A1(n13909), .A2(n13742), .ZN(n6949) );
  AOI22_X1 U7838 ( .A1(n13951), .A2(n13740), .B1(n13739), .B2(n14232), .ZN(
        n13936) );
  NAND2_X1 U7839 ( .A1(n13997), .A2(n13977), .ZN(n13974) );
  NAND2_X1 U7840 ( .A1(n11842), .A2(n11841), .ZN(n13998) );
  OR2_X1 U7841 ( .A1(n6648), .A2(n11850), .ZN(n6643) );
  NAND2_X1 U7842 ( .A1(n11715), .A2(n7299), .ZN(n6649) );
  AND2_X1 U7843 ( .A1(n6714), .A2(n11850), .ZN(n6903) );
  NAND2_X1 U7844 ( .A1(n11846), .A2(n11834), .ZN(n6714) );
  INV_X1 U7845 ( .A(n11834), .ZN(n6904) );
  OAI21_X1 U7846 ( .B1(n6902), .B2(n11846), .A(n11834), .ZN(n11836) );
  INV_X1 U7847 ( .A(n11833), .ZN(n6902) );
  OR2_X1 U7848 ( .A1(n11688), .A2(n11884), .ZN(n11717) );
  NAND3_X1 U7849 ( .A1(n6936), .A2(n6933), .A3(n6448), .ZN(n11547) );
  NAND2_X1 U7850 ( .A1(n6921), .A2(n6925), .ZN(n6920) );
  INV_X1 U7851 ( .A(n11076), .ZN(n6921) );
  NAND2_X1 U7852 ( .A1(n11076), .A2(n6929), .ZN(n6926) );
  INV_X1 U7853 ( .A(n14636), .ZN(n14618) );
  NAND2_X1 U7854 ( .A1(n6913), .A2(n11074), .ZN(n11185) );
  NAND2_X1 U7855 ( .A1(n14628), .A2(n14630), .ZN(n6913) );
  OR2_X1 U7856 ( .A1(n9695), .A2(n9185), .ZN(n9187) );
  NAND2_X1 U7857 ( .A1(n9651), .A2(n9650), .ZN(n14034) );
  NOR2_X1 U7858 ( .A1(n13909), .A2(n6639), .ZN(n6638) );
  INV_X1 U7859 ( .A(n7310), .ZN(n6639) );
  OR2_X1 U7860 ( .A1(n11086), .A2(n11085), .ZN(n14636) );
  INV_X1 U7861 ( .A(n13977), .ZN(n14240) );
  OR2_X1 U7862 ( .A1(n14704), .A2(n11085), .ZN(n11054) );
  NAND2_X1 U7863 ( .A1(n10318), .A2(n10317), .ZN(n14708) );
  AND2_X1 U7864 ( .A1(n10106), .A2(n10105), .ZN(n10310) );
  AND2_X1 U7865 ( .A1(n10596), .A2(n10033), .ZN(n11056) );
  NAND2_X1 U7866 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n6912) );
  AND2_X1 U7867 ( .A1(n14263), .A2(n9180), .ZN(n6911) );
  NAND2_X1 U7868 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(n9445), .ZN(n6909) );
  OAI21_X1 U7869 ( .B1(n14263), .B2(n9180), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6910) );
  OR2_X1 U7870 ( .A1(n8188), .A2(n8187), .ZN(n8230) );
  INV_X1 U7871 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9180) );
  NAND2_X1 U7872 ( .A1(n7867), .A2(n7868), .ZN(n7895) );
  OR2_X1 U7873 ( .A1(n7894), .A2(n11578), .ZN(n7891) );
  AND2_X1 U7874 ( .A1(n9201), .A2(n9206), .ZN(n7276) );
  NAND2_X1 U7875 ( .A1(n7808), .A2(n7809), .ZN(n7256) );
  INV_X1 U7876 ( .A(n7810), .ZN(n7809) );
  INV_X1 U7877 ( .A(n7826), .ZN(n7255) );
  XNOR2_X1 U7878 ( .A(n6710), .B(n7702), .ZN(n10645) );
  NAND2_X1 U7879 ( .A1(n7675), .A2(n7674), .ZN(n6710) );
  NAND2_X1 U7880 ( .A1(n6711), .A2(n6736), .ZN(n7675) );
  NAND2_X1 U7881 ( .A1(n7656), .A2(n7655), .ZN(n6711) );
  NAND2_X1 U7882 ( .A1(n7250), .A2(n7248), .ZN(n7598) );
  AOI21_X1 U7883 ( .B1(n7251), .B2(n7253), .A(n7249), .ZN(n7248) );
  INV_X1 U7884 ( .A(n7594), .ZN(n7249) );
  NAND2_X1 U7885 ( .A1(n7598), .A2(n7597), .ZN(n7613) );
  NAND2_X1 U7886 ( .A1(n7573), .A2(n7572), .ZN(n7593) );
  NAND2_X1 U7887 ( .A1(n7553), .A2(n7552), .ZN(n7573) );
  OR2_X1 U7888 ( .A1(n9339), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9354) );
  NAND2_X1 U7889 ( .A1(n6650), .A2(SI_6_), .ZN(n7525) );
  INV_X1 U7890 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9163) );
  AND2_X1 U7891 ( .A1(n6672), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14330) );
  NOR2_X1 U7892 ( .A1(n14344), .A2(n14345), .ZN(n14346) );
  AOI21_X1 U7893 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(n14311), .A(n14310), .ZN(
        n14363) );
  NOR2_X1 U7894 ( .A1(n14561), .A2(n6660), .ZN(n6659) );
  NAND2_X1 U7895 ( .A1(n6664), .A2(n14371), .ZN(n6663) );
  INV_X1 U7896 ( .A(n14557), .ZN(n6664) );
  OAI21_X1 U7897 ( .B1(n14387), .B2(n11423), .A(n14419), .ZN(n14425) );
  AOI21_X1 U7898 ( .B1(n12556), .B2(n8806), .A(n8821), .ZN(n12442) );
  AND3_X1 U7899 ( .A1(n8717), .A2(n8716), .A3(n8715), .ZN(n12653) );
  NAND2_X1 U7900 ( .A1(n8816), .A2(n8815), .ZN(n12330) );
  NAND2_X1 U7901 ( .A1(n6861), .A2(n8439), .ZN(n15085) );
  INV_X1 U7902 ( .A(n6862), .ZN(n6861) );
  NAND2_X1 U7903 ( .A1(n8438), .A2(n8437), .ZN(n8439) );
  OAI22_X1 U7904 ( .A1(n7369), .A2(n8449), .B1(n8448), .B2(n10065), .ZN(n6862)
         );
  AND2_X1 U7905 ( .A1(n8797), .A2(n8796), .ZN(n12596) );
  NAND2_X1 U7906 ( .A1(n12281), .A2(n12280), .ZN(n12344) );
  NAND2_X1 U7907 ( .A1(n8656), .A2(n8655), .ZN(n12803) );
  AND2_X1 U7908 ( .A1(n8759), .A2(n8758), .ZN(n12643) );
  NAND2_X1 U7909 ( .A1(n8740), .A2(n8739), .ZN(n12403) );
  INV_X1 U7910 ( .A(n12591), .ZN(n12758) );
  INV_X1 U7911 ( .A(n9845), .ZN(n7168) );
  INV_X1 U7912 ( .A(n12595), .ZN(n12630) );
  INV_X1 U7913 ( .A(n12653), .ZN(n12675) );
  INV_X1 U7914 ( .A(n11566), .ZN(n15040) );
  XNOR2_X1 U7915 ( .A(n9070), .B(n8437), .ZN(n10505) );
  OR2_X1 U7916 ( .A1(n14987), .A2(n9068), .ZN(n7020) );
  OAI21_X1 U7917 ( .B1(n12532), .B2(n6450), .A(n9160), .ZN(n7076) );
  NOR2_X1 U7918 ( .A1(n12506), .A2(n9057), .ZN(n12525) );
  NAND2_X1 U7919 ( .A1(n6995), .A2(n9058), .ZN(n9059) );
  NAND2_X1 U7920 ( .A1(n12612), .A2(n8966), .ZN(n12594) );
  NAND2_X1 U7921 ( .A1(n8752), .A2(n8751), .ZN(n12771) );
  CLKBUF_X1 U7922 ( .A(n12714), .Z(n12715) );
  AOI21_X1 U7923 ( .B1(n15143), .B2(n12755), .A(n12754), .ZN(n12826) );
  NAND2_X1 U7924 ( .A1(n8669), .A2(n8668), .ZN(n12857) );
  NAND2_X1 U7925 ( .A1(n8639), .A2(n8638), .ZN(n12862) );
  NAND2_X1 U7926 ( .A1(n8622), .A2(n8621), .ZN(n12866) );
  NAND2_X1 U7927 ( .A1(n8402), .A2(n8384), .ZN(n12029) );
  MUX2_X1 U7928 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8383), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n8384) );
  OR2_X1 U7929 ( .A1(n8385), .A2(n6901), .ZN(n6604) );
  NOR2_X1 U7930 ( .A1(n6428), .A2(n6603), .ZN(n6602) );
  AND2_X1 U7931 ( .A1(n8847), .A2(n6480), .ZN(n11339) );
  INV_X1 U7932 ( .A(n11669), .ZN(n7220) );
  AND2_X1 U7933 ( .A1(n7695), .A2(n7218), .ZN(n7217) );
  NAND2_X1 U7934 ( .A1(n11669), .A2(n7219), .ZN(n7218) );
  INV_X1 U7935 ( .A(n11653), .ZN(n7219) );
  NAND2_X1 U7936 ( .A1(n12210), .A2(n6683), .ZN(n11651) );
  NOR2_X1 U7937 ( .A1(n6499), .A2(n6684), .ZN(n6683) );
  INV_X1 U7938 ( .A(n7635), .ZN(n6684) );
  NAND2_X1 U7939 ( .A1(n7792), .A2(n7791), .ZN(n13229) );
  NAND2_X1 U7940 ( .A1(n11668), .A2(n11669), .ZN(n11667) );
  XNOR2_X1 U7941 ( .A(n7865), .B(n7863), .ZN(n12955) );
  NAND2_X1 U7942 ( .A1(n11451), .A2(n7631), .ZN(n12210) );
  AND2_X1 U7943 ( .A1(n12204), .A2(n7630), .ZN(n7631) );
  OR3_X1 U7944 ( .A1(n8035), .A2(n10113), .A3(n14490), .ZN(n12971) );
  NAND2_X1 U7945 ( .A1(n7708), .A2(n7707), .ZN(n11860) );
  AND2_X1 U7946 ( .A1(n7081), .A2(n8294), .ZN(n6746) );
  INV_X1 U7947 ( .A(n8300), .ZN(n6741) );
  NAND2_X1 U7948 ( .A1(n6739), .A2(n8300), .ZN(n6738) );
  NAND2_X1 U7949 ( .A1(n6745), .A2(n12034), .ZN(n6739) );
  OR2_X1 U7950 ( .A1(n7081), .A2(n8295), .ZN(n6745) );
  AND2_X1 U7951 ( .A1(n8238), .A2(n8237), .ZN(n13086) );
  AOI21_X2 U7952 ( .B1(n10017), .B2(n14475), .A(n10016), .ZN(n13301) );
  NAND2_X1 U7953 ( .A1(n10015), .A2(n10014), .ZN(n10016) );
  AOI21_X1 U7954 ( .B1(n13299), .B2(n14847), .A(n10028), .ZN(n10029) );
  AND2_X2 U7955 ( .A1(n10493), .A2(n10492), .ZN(n14903) );
  NAND2_X1 U7956 ( .A1(n8203), .A2(n8202), .ZN(n13378) );
  NAND2_X1 U7957 ( .A1(n7814), .A2(n7813), .ZN(n13406) );
  OR2_X1 U7958 ( .A1(n11534), .A2(n8235), .ZN(n7814) );
  NAND2_X1 U7959 ( .A1(n9662), .A2(n9661), .ZN(n14028) );
  AND3_X1 U7960 ( .A1(n9471), .A2(n9470), .A3(n9469), .ZN(n13955) );
  INV_X1 U7961 ( .A(n13557), .ZN(n13537) );
  AND2_X1 U7962 ( .A1(n10164), .A2(n13587), .ZN(n13981) );
  AND2_X1 U7963 ( .A1(n11056), .A2(n10735), .ZN(n10747) );
  INV_X1 U7964 ( .A(n9681), .ZN(n13773) );
  AND2_X1 U7965 ( .A1(n9408), .A2(n9420), .ZN(n10532) );
  NAND2_X1 U7966 ( .A1(n6620), .A2(n6619), .ZN(n6618) );
  OR2_X1 U7967 ( .A1(n13689), .A2(n13688), .ZN(n6620) );
  AOI21_X1 U7968 ( .B1(n13690), .B2(n14602), .A(n14595), .ZN(n6619) );
  OAI21_X1 U7969 ( .B1(n13724), .B2(n6637), .A(n6636), .ZN(n13812) );
  NOR2_X1 U7970 ( .A1(n13822), .A2(n7254), .ZN(n13807) );
  NOR2_X1 U7971 ( .A1(n13966), .A2(n7307), .ZN(n7306) );
  INV_X1 U7972 ( .A(n13712), .ZN(n7307) );
  NAND2_X1 U7973 ( .A1(n13962), .A2(n11089), .ZN(n14002) );
  NAND2_X1 U7974 ( .A1(n6668), .A2(n6667), .ZN(n14409) );
  NAND2_X1 U7975 ( .A1(n14404), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n6667) );
  NAND2_X1 U7976 ( .A1(n6670), .A2(n6492), .ZN(n6668) );
  AOI21_X1 U7977 ( .B1(n7040), .B2(n7039), .A(n14370), .ZN(n14558) );
  INV_X1 U7978 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7039) );
  INV_X1 U7979 ( .A(n7041), .ZN(n14368) );
  INV_X1 U7980 ( .A(n6661), .ZN(n6658) );
  INV_X1 U7981 ( .A(n6659), .ZN(n6656) );
  INV_X1 U7982 ( .A(n7042), .ZN(n14569) );
  INV_X1 U7983 ( .A(n14565), .ZN(n7043) );
  XNOR2_X1 U7984 ( .A(n14425), .B(n14424), .ZN(n14423) );
  NOR2_X1 U7985 ( .A1(n9310), .A2(n10631), .ZN(n9223) );
  NAND2_X1 U7986 ( .A1(n9311), .A2(n7286), .ZN(n7285) );
  NAND2_X1 U7987 ( .A1(n9343), .A2(n9345), .ZN(n6586) );
  OR2_X1 U7988 ( .A1(n7283), .A2(n9379), .ZN(n7282) );
  INV_X1 U7989 ( .A(n9378), .ZN(n7283) );
  OR2_X1 U7990 ( .A1(n8072), .A2(n7096), .ZN(n7095) );
  INV_X1 U7991 ( .A(n8070), .ZN(n7096) );
  NOR2_X1 U7992 ( .A1(n8073), .A2(n8070), .ZN(n7097) );
  NAND2_X1 U7993 ( .A1(n8082), .A2(n8084), .ZN(n7086) );
  AND2_X1 U7994 ( .A1(n9498), .A2(n7266), .ZN(n7260) );
  NAND2_X1 U7995 ( .A1(n9498), .A2(n7263), .ZN(n7262) );
  INV_X1 U7996 ( .A(n7264), .ZN(n7263) );
  AOI21_X1 U7997 ( .B1(n7266), .B2(n11835), .A(n7265), .ZN(n7264) );
  INV_X1 U7998 ( .A(n9460), .ZN(n7265) );
  OAI21_X1 U7999 ( .B1(n8094), .B2(n7109), .A(n6503), .ZN(n8100) );
  OR2_X1 U8000 ( .A1(n7291), .A2(n9547), .ZN(n7290) );
  INV_X1 U8001 ( .A(n9546), .ZN(n7291) );
  MUX2_X1 U8002 ( .A(n13745), .B(n13875), .S(n9289), .Z(n9562) );
  INV_X1 U8003 ( .A(n7090), .ZN(n6577) );
  AOI21_X1 U8004 ( .B1(n6501), .B2(n7090), .A(n7089), .ZN(n7088) );
  INV_X1 U8005 ( .A(n8118), .ZN(n7089) );
  OAI21_X1 U8006 ( .B1(n8122), .B2(n7103), .A(n6502), .ZN(n8127) );
  INV_X1 U8007 ( .A(n8749), .ZN(n7143) );
  NAND2_X1 U8008 ( .A1(n7119), .A2(n7117), .ZN(n7116) );
  NAND2_X1 U8009 ( .A1(n9652), .A2(n9654), .ZN(n7269) );
  INV_X1 U8010 ( .A(n15085), .ZN(n9802) );
  INV_X1 U8011 ( .A(n6874), .ZN(n6873) );
  INV_X1 U8012 ( .A(n6872), .ZN(n6871) );
  OAI21_X1 U8013 ( .B1(n6467), .B2(n6873), .A(n9837), .ZN(n6872) );
  OR2_X1 U8014 ( .A1(n12403), .A2(n12629), .ZN(n9837) );
  NOR2_X1 U8015 ( .A1(n7112), .A2(n6554), .ZN(n7111) );
  INV_X1 U8016 ( .A(n8171), .ZN(n7112) );
  NOR2_X1 U8017 ( .A1(n8166), .A2(n8163), .ZN(n7114) );
  NAND2_X1 U8018 ( .A1(n8163), .A2(n8166), .ZN(n7113) );
  MUX2_X1 U8019 ( .A(n8219), .B(n10027), .S(n8262), .Z(n8249) );
  NOR2_X1 U8020 ( .A1(n8249), .A2(n8248), .ZN(n8224) );
  MUX2_X1 U8021 ( .A(n13306), .B(n12889), .S(n8096), .Z(n8225) );
  NOR2_X1 U8022 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n6595) );
  INV_X1 U8023 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n7347) );
  INV_X1 U8024 ( .A(n7914), .ZN(n6748) );
  NOR2_X1 U8025 ( .A1(n7954), .A2(n6753), .ZN(n6752) );
  INV_X1 U8026 ( .A(n7933), .ZN(n6753) );
  INV_X1 U8027 ( .A(n7805), .ZN(n6725) );
  NOR2_X1 U8028 ( .A1(n6440), .A2(n7805), .ZN(n6723) );
  INV_X1 U8029 ( .A(n7745), .ZN(n7238) );
  INV_X1 U8030 ( .A(n7784), .ZN(n7789) );
  AND2_X1 U8031 ( .A1(n6730), .A2(n6535), .ZN(n6727) );
  AND2_X1 U8032 ( .A1(n7243), .A2(n6731), .ZN(n6730) );
  NAND2_X1 U8033 ( .A1(n6736), .A2(n6732), .ZN(n6731) );
  INV_X1 U8034 ( .A(n7244), .ZN(n7243) );
  OAI21_X1 U8035 ( .B1(n7246), .B2(n7245), .A(n7722), .ZN(n7244) );
  INV_X1 U8036 ( .A(n7701), .ZN(n7245) );
  INV_X1 U8037 ( .A(n11739), .ZN(n7213) );
  AND3_X1 U8038 ( .A1(n8502), .A2(n8501), .A3(n8500), .ZN(n11175) );
  AND3_X1 U8039 ( .A1(n7078), .A2(n7077), .A3(P3_REG1_REG_0__SCAN_IN), .ZN(
        n9126) );
  INV_X1 U8040 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n7078) );
  INV_X1 U8041 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7077) );
  NOR2_X1 U8042 ( .A1(n10682), .A2(n9134), .ZN(n14938) );
  INV_X1 U8043 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11981) );
  INV_X1 U8044 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n12294) );
  AND2_X1 U8045 ( .A1(n8824), .A2(n8823), .ZN(n8982) );
  NAND2_X1 U8046 ( .A1(n6803), .A2(n8966), .ZN(n6799) );
  INV_X1 U8047 ( .A(n6801), .ZN(n6800) );
  INV_X1 U8048 ( .A(n12580), .ZN(n12581) );
  OR2_X1 U8049 ( .A1(n12857), .A2(n12725), .ZN(n8858) );
  INV_X1 U8050 ( .A(n14455), .ZN(n6783) );
  AOI21_X1 U8051 ( .B1(n11198), .B2(n8890), .A(n11387), .ZN(n6779) );
  INV_X1 U8052 ( .A(n8890), .ZN(n6780) );
  AOI21_X1 U8053 ( .B1(n6566), .B2(n7144), .A(n7142), .ZN(n7141) );
  NOR2_X1 U8054 ( .A1(n9575), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7142) );
  INV_X1 U8055 ( .A(n8337), .ZN(n7165) );
  NOR2_X1 U8056 ( .A1(n6865), .A2(n6867), .ZN(n8376) );
  NAND2_X1 U8057 ( .A1(n8375), .A2(n8373), .ZN(n6865) );
  OR2_X1 U8058 ( .A1(n8650), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n8651) );
  INV_X1 U8059 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n8318) );
  AND2_X1 U8060 ( .A1(n7771), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n7793) );
  NOR2_X1 U8061 ( .A1(n7751), .A2(n7750), .ZN(n7771) );
  INV_X1 U8062 ( .A(n12926), .ZN(n6682) );
  INV_X1 U8063 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n7679) );
  INV_X1 U8064 ( .A(n9946), .ZN(n7036) );
  NAND2_X1 U8065 ( .A1(n6765), .A2(n6764), .ZN(n6768) );
  NOR2_X1 U8066 ( .A1(n6769), .A2(n6766), .ZN(n6764) );
  INV_X1 U8067 ( .A(n13215), .ZN(n6765) );
  NOR2_X1 U8068 ( .A1(n7688), .A2(n7685), .ZN(n7709) );
  NOR2_X1 U8069 ( .A1(n7580), .A2(n7579), .ZN(n7624) );
  AOI21_X1 U8070 ( .B1(n7025), .B2(n7029), .A(n6495), .ZN(n7022) );
  NAND2_X1 U8071 ( .A1(n13226), .A2(n7025), .ZN(n7023) );
  NAND2_X1 U8072 ( .A1(n9960), .A2(n9959), .ZN(n10705) );
  OR2_X1 U8073 ( .A1(n7575), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n7600) );
  OR3_X1 U8074 ( .A1(n7556), .A2(P2_IR_REG_7__SCAN_IN), .A3(
        P2_IR_REG_6__SCAN_IN), .ZN(n7575) );
  INV_X1 U8075 ( .A(n9586), .ZN(n9587) );
  NOR2_X1 U8076 ( .A1(n12070), .A2(n12062), .ZN(n6984) );
  NAND2_X1 U8077 ( .A1(n7272), .A2(n7271), .ZN(n9711) );
  OR2_X1 U8078 ( .A1(n7275), .A2(n9684), .ZN(n7271) );
  OAI21_X1 U8079 ( .B1(n6701), .B2(n6699), .A(n6698), .ZN(n6697) );
  AOI21_X1 U8080 ( .B1(n13791), .B2(n6707), .A(n6705), .ZN(n6698) );
  AND2_X1 U8081 ( .A1(n14034), .A2(n13751), .ZN(n6705) );
  AND2_X1 U8082 ( .A1(n13942), .A2(n6821), .ZN(n13874) );
  AND2_X1 U8083 ( .A1(n6823), .A2(n6822), .ZN(n6821) );
  NOR2_X1 U8084 ( .A1(n13915), .A2(n6825), .ZN(n6823) );
  NOR2_X1 U8085 ( .A1(n13974), .A2(n14232), .ZN(n13942) );
  OR2_X1 U8086 ( .A1(n14522), .A2(n12051), .ZN(n13735) );
  NOR2_X1 U8087 ( .A1(n11717), .A2(n11934), .ZN(n11842) );
  OAI21_X1 U8088 ( .B1(n11506), .B2(n7298), .A(n11291), .ZN(n7297) );
  NAND2_X1 U8089 ( .A1(n11294), .A2(n6918), .ZN(n6917) );
  INV_X1 U8090 ( .A(n6925), .ZN(n6918) );
  NAND2_X1 U8091 ( .A1(n14638), .A2(n13572), .ZN(n11063) );
  NAND2_X1 U8092 ( .A1(n13826), .A2(n13750), .ZN(n13800) );
  NAND2_X1 U8093 ( .A1(n11511), .A2(n6436), .ZN(n11434) );
  AND2_X1 U8094 ( .A1(n9720), .A2(n11268), .ZN(n10592) );
  XNOR2_X1 U8095 ( .A(n9771), .B(n9770), .ZN(n10163) );
  NAND2_X1 U8096 ( .A1(n7828), .A2(SI_21_), .ZN(n7846) );
  OR2_X1 U8097 ( .A1(n9493), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n9473) );
  AND2_X1 U8098 ( .A1(n7317), .A2(n9199), .ZN(n9444) );
  INV_X1 U8099 ( .A(n7252), .ZN(n7251) );
  OAI21_X1 U8100 ( .B1(n7552), .B2(n7253), .A(n7592), .ZN(n7252) );
  INV_X1 U8101 ( .A(n7572), .ZN(n7253) );
  AND2_X2 U8102 ( .A1(n7258), .A2(n7257), .ZN(n7479) );
  INV_X1 U8103 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7363) );
  NAND2_X1 U8104 ( .A1(n7056), .A2(n14296), .ZN(n14297) );
  NAND2_X1 U8105 ( .A1(n14325), .A2(n14324), .ZN(n7056) );
  XNOR2_X1 U8106 ( .A(n14297), .B(n7055), .ZN(n14340) );
  INV_X1 U8107 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n7055) );
  OR2_X1 U8108 ( .A1(n12249), .A2(n6544), .ZN(n7208) );
  NAND2_X1 U8109 ( .A1(n8389), .A2(n8388), .ZN(n8623) );
  INV_X1 U8110 ( .A(n8610), .ZN(n8389) );
  INV_X1 U8111 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n8533) );
  NAND2_X1 U8112 ( .A1(n9799), .A2(n7438), .ZN(n8448) );
  INV_X1 U8113 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n10679) );
  NAND2_X1 U8114 ( .A1(n12334), .A2(n12273), .ZN(n12303) );
  XNOR2_X1 U8115 ( .A(n6804), .B(n9885), .ZN(n7169) );
  NAND2_X1 U8116 ( .A1(n6806), .A2(n6805), .ZN(n6804) );
  NAND2_X1 U8117 ( .A1(n8983), .A2(n12818), .ZN(n6805) );
  NAND2_X1 U8118 ( .A1(n6808), .A2(n6807), .ZN(n6806) );
  AND4_X1 U8119 ( .A1(n8602), .A2(n8601), .A3(n8600), .A4(n8599), .ZN(n12247)
         );
  AOI21_X1 U8120 ( .B1(n8440), .B2(P3_REG2_REG_3__SCAN_IN), .A(n8461), .ZN(
        n10780) );
  NOR2_X1 U8121 ( .A1(n10507), .A2(n15147), .ZN(n10506) );
  NOR2_X1 U8122 ( .A1(n10506), .A2(n9126), .ZN(n10449) );
  INV_X1 U8123 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n14291) );
  NAND2_X1 U8124 ( .A1(n6999), .A2(n7005), .ZN(n6998) );
  INV_X1 U8125 ( .A(n7017), .ZN(n7016) );
  NOR2_X1 U8126 ( .A1(n7015), .A2(n9036), .ZN(n14911) );
  NAND2_X1 U8127 ( .A1(n7064), .A2(n6441), .ZN(n10469) );
  NAND2_X1 U8128 ( .A1(n10469), .A2(n10470), .ZN(n10468) );
  AND2_X1 U8129 ( .A1(n7015), .A2(n7014), .ZN(n10467) );
  NOR2_X1 U8130 ( .A1(n10466), .A2(n10467), .ZN(n10465) );
  NAND2_X1 U8131 ( .A1(n10462), .A2(n6600), .ZN(n10678) );
  NAND2_X1 U8132 ( .A1(n6601), .A2(n9132), .ZN(n6600) );
  INV_X1 U8133 ( .A(n9074), .ZN(n6601) );
  XNOR2_X1 U8134 ( .A(n9133), .B(n7079), .ZN(n10683) );
  NOR2_X1 U8135 ( .A1(n10683), .A2(n15155), .ZN(n10682) );
  AOI21_X1 U8136 ( .B1(n14933), .B2(n14932), .A(n14931), .ZN(n14930) );
  NOR2_X1 U8137 ( .A1(n10790), .A2(n9138), .ZN(n10996) );
  NOR2_X1 U8138 ( .A1(n10996), .A2(n10995), .ZN(n10994) );
  NOR2_X1 U8139 ( .A1(n14977), .A2(n14978), .ZN(n14976) );
  NAND2_X1 U8140 ( .A1(n7067), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n7066) );
  NAND2_X1 U8141 ( .A1(n9141), .A2(n7067), .ZN(n7065) );
  NOR2_X1 U8142 ( .A1(n14976), .A2(n9092), .ZN(n14993) );
  NAND2_X1 U8143 ( .A1(n7070), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n7069) );
  NAND2_X1 U8144 ( .A1(n9145), .A2(n7070), .ZN(n7068) );
  INV_X1 U8145 ( .A(n12463), .ZN(n7070) );
  NOR2_X1 U8146 ( .A1(n14991), .A2(n9067), .ZN(n14990) );
  AND2_X1 U8147 ( .A1(n10100), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n6597) );
  INV_X1 U8148 ( .A(n12453), .ZN(n6598) );
  NAND2_X1 U8149 ( .A1(n9096), .A2(n9097), .ZN(n15013) );
  OR2_X1 U8150 ( .A1(n12456), .A2(n12455), .ZN(n9096) );
  NOR2_X1 U8151 ( .A1(n15010), .A2(n15011), .ZN(n15009) );
  NAND2_X1 U8152 ( .A1(n9102), .A2(n6605), .ZN(n14442) );
  NAND2_X1 U8153 ( .A1(n6606), .A2(n14437), .ZN(n6605) );
  NOR2_X1 U8154 ( .A1(n14442), .A2(n14443), .ZN(n14441) );
  NAND2_X1 U8155 ( .A1(n7073), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n7072) );
  NAND2_X1 U8156 ( .A1(n9152), .A2(n7073), .ZN(n7071) );
  INV_X1 U8157 ( .A(n12499), .ZN(n7073) );
  NOR2_X1 U8158 ( .A1(n14439), .A2(n14440), .ZN(n14438) );
  OR2_X1 U8159 ( .A1(n12489), .A2(n14435), .ZN(n7011) );
  NAND2_X1 U8160 ( .A1(n9054), .A2(n7010), .ZN(n7009) );
  INV_X1 U8161 ( .A(n12489), .ZN(n7010) );
  NOR2_X1 U8162 ( .A1(n12517), .A2(n9156), .ZN(n12534) );
  NAND2_X1 U8163 ( .A1(n12526), .A2(n9110), .ZN(n6608) );
  XNOR2_X1 U8164 ( .A(n12330), .B(n12442), .ZN(n9797) );
  OR2_X1 U8165 ( .A1(n8971), .A2(n8970), .ZN(n12580) );
  NAND2_X1 U8166 ( .A1(n9841), .A2(n6897), .ZN(n6893) );
  AOI21_X1 U8167 ( .B1(n6897), .B2(n9840), .A(n7343), .ZN(n6896) );
  INV_X1 U8168 ( .A(n8779), .ZN(n8399) );
  AND2_X1 U8169 ( .A1(n12771), .A2(n12444), .ZN(n9838) );
  NAND2_X1 U8170 ( .A1(n12625), .A2(n8771), .ZN(n12612) );
  NAND2_X1 U8171 ( .A1(n8397), .A2(n8396), .ZN(n8753) );
  INV_X1 U8172 ( .A(n8741), .ZN(n8397) );
  AOI21_X1 U8173 ( .B1(n6795), .B2(n6798), .A(n6794), .ZN(n6793) );
  INV_X1 U8174 ( .A(n8955), .ZN(n6794) );
  NAND2_X1 U8175 ( .A1(n8395), .A2(n8394), .ZN(n8728) );
  NAND2_X1 U8176 ( .A1(n8393), .A2(n8392), .ZN(n8702) );
  INV_X1 U8177 ( .A(n8687), .ZN(n8393) );
  NAND2_X1 U8178 ( .A1(n6882), .A2(n6881), .ZN(n12688) );
  NAND2_X1 U8179 ( .A1(n8391), .A2(n12354), .ZN(n8670) );
  NAND2_X1 U8180 ( .A1(n11910), .A2(n9827), .ZN(n12735) );
  INV_X1 U8181 ( .A(n12710), .ZN(n12738) );
  NAND2_X1 U8182 ( .A1(n11911), .A2(n11914), .ZN(n11910) );
  NAND2_X1 U8183 ( .A1(n6890), .A2(n6888), .ZN(n11820) );
  NAND2_X1 U8184 ( .A1(n6889), .A2(n12447), .ZN(n6888) );
  INV_X1 U8185 ( .A(n14457), .ZN(n6889) );
  OR2_X1 U8186 ( .A1(n8571), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8597) );
  AOI21_X1 U8187 ( .B1(n6886), .B2(n11317), .A(n6885), .ZN(n6884) );
  INV_X1 U8188 ( .A(n9821), .ZN(n6885) );
  NAND2_X1 U8189 ( .A1(n6788), .A2(n8562), .ZN(n15025) );
  NAND2_X1 U8190 ( .A1(n8550), .A2(n6789), .ZN(n6788) );
  AND2_X1 U8191 ( .A1(n8534), .A2(n8533), .ZN(n8551) );
  NAND2_X1 U8192 ( .A1(n8551), .A2(n11740), .ZN(n8571) );
  INV_X1 U8193 ( .A(n8905), .ZN(n15046) );
  NAND2_X1 U8194 ( .A1(n11194), .A2(n8989), .ZN(n6778) );
  OR2_X1 U8195 ( .A1(n8505), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8520) );
  NAND2_X1 U8196 ( .A1(n9810), .A2(n9809), .ZN(n11028) );
  AND4_X1 U8197 ( .A1(n8492), .A2(n8491), .A3(n8490), .A4(n8489), .ZN(n11377)
         );
  NAND2_X1 U8198 ( .A1(n10817), .A2(n10816), .ZN(n10819) );
  INV_X1 U8199 ( .A(n10984), .ZN(n9885) );
  NAND2_X1 U8200 ( .A1(n8831), .A2(n8830), .ZN(n9910) );
  OR2_X1 U8201 ( .A1(n9855), .A2(P3_D_REG_0__SCAN_IN), .ZN(n7179) );
  NAND2_X1 U8202 ( .A1(n8362), .A2(n8361), .ZN(n8827) );
  NAND2_X1 U8203 ( .A1(n6814), .A2(n6813), .ZN(n8382) );
  AND2_X1 U8204 ( .A1(n7335), .A2(n6529), .ZN(n6813) );
  NOR2_X1 U8205 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_27__SCAN_IN), .ZN(
        n6603) );
  NAND2_X1 U8206 ( .A1(n8772), .A2(n8349), .ZN(n8775) );
  NAND2_X1 U8207 ( .A1(n7182), .A2(n9017), .ZN(n7181) );
  XNOR2_X1 U8208 ( .A(n9015), .B(n9017), .ZN(n9061) );
  XNOR2_X1 U8209 ( .A(n8842), .B(P3_IR_REG_21__SCAN_IN), .ZN(n10832) );
  AND2_X1 U8210 ( .A1(n8340), .A2(n8339), .ZN(n8721) );
  AND2_X1 U8211 ( .A1(n8337), .A2(n8336), .ZN(n8695) );
  AND2_X1 U8212 ( .A1(n8376), .A2(n7200), .ZN(n7199) );
  INV_X1 U8213 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7200) );
  AND2_X1 U8214 ( .A1(n8333), .A2(n8332), .ZN(n8677) );
  NOR2_X1 U8215 ( .A1(n7159), .A2(n7158), .ZN(n7157) );
  AND2_X1 U8216 ( .A1(n8335), .A2(n8334), .ZN(n8678) );
  AND2_X1 U8217 ( .A1(n8331), .A2(n8330), .ZN(n8648) );
  INV_X1 U8218 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8636) );
  INV_X1 U8219 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8634) );
  AND2_X1 U8220 ( .A1(n8587), .A2(n6545), .ZN(n7160) );
  OR2_X1 U8221 ( .A1(n8593), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n8619) );
  AND2_X1 U8222 ( .A1(n8544), .A2(n8566), .ZN(n9139) );
  AND2_X1 U8223 ( .A1(n8316), .A2(n8315), .ZN(n8545) );
  NAND2_X1 U8224 ( .A1(n7133), .A2(n7131), .ZN(n8546) );
  AOI21_X1 U8225 ( .B1(n7132), .B2(n7135), .A(n6556), .ZN(n7131) );
  AND2_X1 U8226 ( .A1(n8515), .A2(n8541), .ZN(n14942) );
  NAND2_X1 U8227 ( .A1(n7002), .A2(n7003), .ZN(n9122) );
  NAND2_X1 U8228 ( .A1(n8426), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8433) );
  AND2_X1 U8229 ( .A1(n7992), .A2(n7991), .ZN(n8003) );
  OR2_X1 U8230 ( .A1(n7539), .A2(n7538), .ZN(n7561) );
  XNOR2_X1 U8231 ( .A(n7410), .B(n7412), .ZN(n10695) );
  OR2_X1 U8232 ( .A1(n7733), .A2(n11971), .ZN(n7751) );
  NAND2_X1 U8233 ( .A1(n10857), .A2(n7435), .ZN(n10407) );
  NAND2_X1 U8234 ( .A1(n7793), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n7816) );
  INV_X1 U8235 ( .A(n12967), .ZN(n12986) );
  INV_X1 U8236 ( .A(n12984), .ZN(n12946) );
  NAND3_X1 U8237 ( .A1(n10695), .A2(n10689), .A3(n10665), .ZN(n10690) );
  NAND2_X1 U8238 ( .A1(n7216), .A2(n7215), .ZN(n7720) );
  AOI21_X1 U8239 ( .B1(n7217), .B2(n7220), .A(n6507), .ZN(n7215) );
  AND2_X1 U8240 ( .A1(n8252), .A2(n8253), .ZN(n6755) );
  NAND2_X1 U8241 ( .A1(n6478), .A2(n7120), .ZN(n6757) );
  NOR2_X1 U8242 ( .A1(n6485), .A2(n6578), .ZN(n6756) );
  AND2_X1 U8243 ( .A1(n7926), .A2(n7925), .ZN(n12979) );
  AND2_X1 U8244 ( .A1(n7911), .A2(n7910), .ZN(n12924) );
  AND2_X1 U8245 ( .A1(n7886), .A2(n7885), .ZN(n12959) );
  AND2_X1 U8246 ( .A1(n7862), .A2(n7861), .ZN(n12896) );
  NAND2_X1 U8247 ( .A1(n8204), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7401) );
  INV_X1 U8248 ( .A(n10006), .ZN(n10007) );
  NAND2_X1 U8249 ( .A1(n10005), .A2(n8268), .ZN(n13090) );
  AND2_X1 U8250 ( .A1(n13114), .A2(n13306), .ZN(n13102) );
  AND2_X1 U8251 ( .A1(n13318), .A2(n13005), .ZN(n9946) );
  NAND2_X1 U8252 ( .A1(n6850), .A2(n6848), .ZN(n6844) );
  AND2_X1 U8253 ( .A1(n10002), .A2(n13109), .ZN(n6842) );
  NOR2_X1 U8254 ( .A1(n6851), .A2(n6847), .ZN(n6846) );
  NOR2_X1 U8255 ( .A1(n10002), .A2(n10004), .ZN(n13131) );
  INV_X1 U8257 ( .A(n6851), .ZN(n6850) );
  INV_X1 U8258 ( .A(n9943), .ZN(n7059) );
  XNOR2_X1 U8259 ( .A(n13162), .B(n13007), .ZN(n13150) );
  INV_X1 U8260 ( .A(n6768), .ZN(n13169) );
  INV_X1 U8261 ( .A(n6859), .ZN(n6858) );
  OAI21_X1 U8262 ( .B1(n6469), .B2(n6860), .A(n9998), .ZN(n6859) );
  NOR2_X1 U8263 ( .A1(n13215), .A2(n6766), .ZN(n13189) );
  NOR2_X1 U8264 ( .A1(n13215), .A2(n13344), .ZN(n13198) );
  OR2_X1 U8265 ( .A1(n13406), .A2(n13228), .ZN(n13215) );
  NAND2_X1 U8266 ( .A1(n10020), .A2(n6763), .ZN(n6762) );
  NAND2_X1 U8267 ( .A1(n7048), .A2(n7047), .ZN(n7046) );
  INV_X1 U8268 ( .A(n9937), .ZN(n7047) );
  NAND2_X1 U8269 ( .A1(n11896), .A2(n9988), .ZN(n13276) );
  AND2_X1 U8270 ( .A1(n6456), .A2(n11625), .ZN(n14484) );
  NAND2_X1 U8271 ( .A1(n11625), .A2(n6772), .ZN(n14483) );
  AND2_X1 U8272 ( .A1(n9934), .A2(n9935), .ZN(n14481) );
  OR2_X1 U8273 ( .A1(n10444), .A2(n8235), .ZN(n7665) );
  AND2_X1 U8274 ( .A1(n9982), .A2(n8270), .ZN(n11636) );
  NAND2_X1 U8275 ( .A1(n6857), .A2(n9979), .ZN(n11618) );
  AND2_X1 U8276 ( .A1(n14890), .A2(n11497), .ZN(n11625) );
  NAND2_X1 U8277 ( .A1(n11156), .A2(n9923), .ZN(n11227) );
  NAND2_X1 U8278 ( .A1(n11159), .A2(n6839), .ZN(n11239) );
  INV_X1 U8279 ( .A(n10756), .ZN(n6760) );
  NAND2_X1 U8280 ( .A1(n6759), .A2(n6758), .ZN(n10973) );
  NOR2_X1 U8281 ( .A1(n10613), .A2(n10622), .ZN(n10704) );
  NAND2_X1 U8282 ( .A1(n10694), .A2(n10018), .ZN(n10613) );
  NOR2_X1 U8283 ( .A1(n8021), .A2(n14879), .ZN(n9952) );
  NAND2_X1 U8284 ( .A1(n7917), .A2(n7916), .ZN(n10001) );
  AND2_X1 U8285 ( .A1(n9954), .A2(n11535), .ZN(n13362) );
  NAND2_X1 U8286 ( .A1(n7052), .A2(n9936), .ZN(n13283) );
  OR2_X1 U8287 ( .A1(n11903), .A2(n11902), .ZN(n7052) );
  INV_X1 U8288 ( .A(n13362), .ZN(n14511) );
  AND2_X1 U8289 ( .A1(n10118), .A2(n10112), .ZN(n8041) );
  INV_X1 U8290 ( .A(n7358), .ZN(n7361) );
  OR2_X1 U8291 ( .A1(n7485), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n7508) );
  INV_X1 U8292 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7345) );
  INV_X1 U8293 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8426) );
  AND2_X1 U8294 ( .A1(n12004), .A2(n12003), .ZN(n6991) );
  INV_X1 U8295 ( .A(n9568), .ZN(n9569) );
  NAND2_X1 U8296 ( .A1(n10729), .A2(n10728), .ZN(n10730) );
  NAND2_X1 U8297 ( .A1(n12084), .A2(n12083), .ZN(n6968) );
  OR2_X1 U8298 ( .A1(n13510), .A2(n13509), .ZN(n6967) );
  INV_X1 U8299 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9483) );
  NOR2_X1 U8300 ( .A1(n9484), .A2(n9483), .ZN(n9486) );
  NAND2_X1 U8301 ( .A1(n6463), .A2(n10637), .ZN(n10638) );
  NOR2_X1 U8302 ( .A1(n9510), .A2(n9509), .ZN(n9524) );
  NAND2_X1 U8303 ( .A1(n6955), .A2(n6468), .ZN(n13517) );
  OR2_X1 U8304 ( .A1(n13510), .A2(n6963), .ZN(n6955) );
  INV_X1 U8305 ( .A(n13527), .ZN(n6981) );
  NAND2_X1 U8306 ( .A1(n13490), .A2(n12069), .ZN(n6983) );
  NAND2_X1 U8307 ( .A1(n13481), .A2(n6984), .ZN(n6982) );
  NAND2_X1 U8308 ( .A1(n9749), .A2(n9748), .ZN(n9764) );
  AND4_X2 U8309 ( .A1(n9233), .A2(n9232), .A3(n9231), .A4(n9230), .ZN(n11073)
         );
  OR2_X1 U8310 ( .A1(n9675), .A2(n9229), .ZN(n9232) );
  INV_X1 U8311 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14341) );
  NOR2_X1 U8312 ( .A1(n14571), .A2(n6471), .ZN(n13627) );
  NAND2_X1 U8313 ( .A1(n13627), .A2(n13628), .ZN(n13626) );
  OR2_X1 U8314 ( .A1(n9321), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n9339) );
  INV_X1 U8315 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14309) );
  OR2_X1 U8316 ( .A1(n9420), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n9430) );
  OAI22_X1 U8317 ( .A1(n6616), .A2(n11695), .B1(n11697), .B2(n11696), .ZN(
        n11698) );
  NAND2_X1 U8318 ( .A1(n11698), .A2(n11699), .ZN(n13667) );
  NAND2_X1 U8319 ( .A1(n6631), .A2(n13732), .ZN(n6630) );
  INV_X1 U8320 ( .A(n13754), .ZN(n6631) );
  INV_X1 U8321 ( .A(n7315), .ZN(n6637) );
  AOI21_X1 U8322 ( .B1(n7315), .B2(n13851), .A(n6482), .ZN(n6636) );
  AND2_X1 U8323 ( .A1(n13727), .A2(n13726), .ZN(n7315) );
  NOR2_X1 U8324 ( .A1(n14045), .A2(n13843), .ZN(n13826) );
  AND2_X1 U8325 ( .A1(n14283), .A2(n9558), .ZN(n13875) );
  NAND2_X1 U8326 ( .A1(n13885), .A2(n6708), .ZN(n13871) );
  NAND2_X1 U8327 ( .A1(n6822), .A2(n13904), .ZN(n6708) );
  NAND2_X1 U8328 ( .A1(n13901), .A2(n6709), .ZN(n13887) );
  NAND2_X1 U8329 ( .A1(n14082), .A2(n13559), .ZN(n6709) );
  NAND2_X1 U8330 ( .A1(n13887), .A2(n13886), .ZN(n13885) );
  NAND2_X1 U8331 ( .A1(n13942), .A2(n6823), .ZN(n13907) );
  NAND2_X1 U8332 ( .A1(n13942), .A2(n13695), .ZN(n13943) );
  OR2_X1 U8333 ( .A1(n9478), .A2(n9466), .ZN(n9510) );
  INV_X1 U8334 ( .A(n13737), .ZN(n13980) );
  NOR2_X1 U8335 ( .A1(n13998), .A2(n14522), .ZN(n13997) );
  AND4_X1 U8336 ( .A1(n9490), .A2(n9489), .A3(n9488), .A4(n9487), .ZN(n13994)
         );
  NAND2_X1 U8337 ( .A1(n6903), .A2(n6904), .ZN(n6713) );
  NAND2_X1 U8338 ( .A1(n6903), .A2(n11833), .ZN(n6712) );
  OR2_X1 U8339 ( .A1(n9435), .A2(n9434), .ZN(n9450) );
  AND2_X1 U8340 ( .A1(n7301), .A2(n11848), .ZN(n7300) );
  NAND2_X1 U8341 ( .A1(n11846), .A2(n7302), .ZN(n7301) );
  INV_X1 U8342 ( .A(n11716), .ZN(n7302) );
  AND4_X1 U8343 ( .A1(n9441), .A2(n9440), .A3(n9439), .A4(n9438), .ZN(n13992)
         );
  NOR2_X1 U8344 ( .A1(n9368), .A2(n10335), .ZN(n9399) );
  INV_X1 U8345 ( .A(n13563), .ZN(n11781) );
  NAND3_X1 U8346 ( .A1(n6437), .A2(n14541), .A3(n11511), .ZN(n11688) );
  OR2_X1 U8347 ( .A1(n9347), .A2(n9346), .ZN(n9368) );
  NAND2_X1 U8348 ( .A1(n6939), .A2(n6934), .ZN(n11439) );
  INV_X1 U8349 ( .A(n6938), .ZN(n6935) );
  INV_X1 U8350 ( .A(n13564), .ZN(n11763) );
  OR2_X1 U8351 ( .A1(n10604), .A2(n13587), .ZN(n13993) );
  NAND2_X1 U8352 ( .A1(n11511), .A2(n11481), .ZN(n11362) );
  NAND2_X1 U8353 ( .A1(n11507), .A2(n11506), .ZN(n11505) );
  AND2_X1 U8354 ( .A1(n14701), .A2(n14620), .ZN(n11511) );
  AND2_X1 U8355 ( .A1(n6454), .A2(n14680), .ZN(n6817) );
  NAND2_X1 U8356 ( .A1(n11076), .A2(n11075), .ZN(n11280) );
  AND2_X1 U8357 ( .A1(n12160), .A2(n10316), .ZN(n11058) );
  NAND2_X1 U8358 ( .A1(n11063), .A2(n11064), .ZN(n14630) );
  NAND2_X1 U8359 ( .A1(n6914), .A2(n11072), .ZN(n14628) );
  NAND2_X1 U8360 ( .A1(n6916), .A2(n6915), .ZN(n6914) );
  INV_X1 U8361 ( .A(n11071), .ZN(n6915) );
  NAND2_X1 U8362 ( .A1(n11084), .A2(n14661), .ZN(n14639) );
  NOR2_X1 U8363 ( .A1(n11060), .A2(n11059), .ZN(n11132) );
  INV_X1 U8364 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n14207) );
  INV_X1 U8365 ( .A(n14017), .ZN(n14023) );
  NAND2_X1 U8366 ( .A1(n6640), .A2(n7310), .ZN(n13910) );
  NAND2_X1 U8367 ( .A1(n6940), .A2(n11301), .ZN(n11366) );
  OR2_X1 U8368 ( .A1(n11510), .A2(n11302), .ZN(n6940) );
  AND2_X1 U8369 ( .A1(n11069), .A2(n11068), .ZN(n7304) );
  INV_X1 U8370 ( .A(n14726), .ZN(n14669) );
  XNOR2_X1 U8371 ( .A(n8215), .B(n8214), .ZN(n9669) );
  XNOR2_X1 U8372 ( .A(n7975), .B(n7974), .ZN(n12021) );
  XNOR2_X1 U8373 ( .A(n6816), .B(n9197), .ZN(n9783) );
  NAND2_X1 U8374 ( .A1(n9781), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6816) );
  OAI21_X1 U8375 ( .B1(n7935), .B2(n7934), .A(n7933), .ZN(n7955) );
  XNOR2_X1 U8376 ( .A(n7935), .B(n7934), .ZN(n13436) );
  NAND2_X1 U8377 ( .A1(n9778), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9779) );
  INV_X1 U8378 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6994) );
  INV_X1 U8379 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9206) );
  INV_X1 U8380 ( .A(n9204), .ZN(n9209) );
  NAND2_X1 U8381 ( .A1(n6720), .A2(n7236), .ZN(n7806) );
  NAND2_X1 U8382 ( .A1(n7746), .A2(n6440), .ZN(n6720) );
  XNOR2_X1 U8383 ( .A(n7766), .B(n7765), .ZN(n11206) );
  NAND2_X1 U8384 ( .A1(n7763), .A2(n7762), .ZN(n7788) );
  NAND2_X1 U8385 ( .A1(n7242), .A2(n7701), .ZN(n7723) );
  NAND2_X1 U8386 ( .A1(n7675), .A2(n7246), .ZN(n7242) );
  NAND2_X1 U8387 ( .A1(n7655), .A2(n6729), .ZN(n6734) );
  NAND2_X1 U8388 ( .A1(n6693), .A2(n6692), .ZN(n6737) );
  AOI21_X1 U8389 ( .B1(n7529), .B2(n6719), .A(n6718), .ZN(n6717) );
  INV_X1 U8390 ( .A(n7525), .ZN(n6719) );
  NAND2_X1 U8391 ( .A1(n7478), .A2(n7477), .ZN(n7483) );
  INV_X1 U8392 ( .A(n7481), .ZN(n7482) );
  NAND2_X1 U8393 ( .A1(n7483), .A2(n7482), .ZN(n7504) );
  OAI21_X1 U8394 ( .B1(n7421), .B2(SI_2_), .A(n7436), .ZN(n7423) );
  XNOR2_X1 U8395 ( .A(n14329), .B(n14330), .ZN(n14331) );
  NAND2_X1 U8396 ( .A1(n14289), .A2(n7053), .ZN(n14328) );
  NAND2_X1 U8397 ( .A1(n7054), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7053) );
  INV_X1 U8398 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7054) );
  XOR2_X1 U8399 ( .A(n14292), .B(P3_ADDR_REG_3__SCAN_IN), .Z(n14336) );
  NAND2_X1 U8400 ( .A1(n6651), .A2(n14349), .ZN(n14351) );
  NAND2_X1 U8401 ( .A1(n14401), .A2(n14400), .ZN(n6651) );
  OR2_X1 U8402 ( .A1(n14404), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n6669) );
  OAI21_X1 U8403 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n14314), .A(n14313), .ZN(
        n14320) );
  NAND2_X1 U8404 ( .A1(n6653), .A2(n6497), .ZN(n14376) );
  NAND2_X1 U8405 ( .A1(n7204), .A2(n7207), .ZN(n12293) );
  OR2_X1 U8406 ( .A1(n7209), .A2(n7208), .ZN(n7204) );
  AOI22_X1 U8407 ( .A1(n7192), .A2(n6543), .B1(n7190), .B2(n7195), .ZN(n7188)
         );
  OR2_X1 U8408 ( .A1(n12361), .A2(n7189), .ZN(n7187) );
  NAND2_X1 U8409 ( .A1(n7177), .A2(n10774), .ZN(n10775) );
  NAND2_X1 U8410 ( .A1(n12380), .A2(n12270), .ZN(n12336) );
  NAND2_X1 U8411 ( .A1(n8727), .A2(n8726), .ZN(n12341) );
  OAI21_X1 U8412 ( .B1(n10784), .B2(n7185), .A(n7184), .ZN(n11376) );
  AOI21_X1 U8413 ( .B1(n7186), .B2(n10782), .A(n6483), .ZN(n7184) );
  INV_X1 U8414 ( .A(n7186), .ZN(n7185) );
  OR2_X1 U8415 ( .A1(n12361), .A2(n12362), .ZN(n12363) );
  OAI21_X1 U8416 ( .B1(n12370), .B2(n12444), .A(n7326), .ZN(n12373) );
  OR2_X1 U8417 ( .A1(n12369), .A2(n6538), .ZN(n7326) );
  NAND2_X1 U8418 ( .A1(n11009), .A2(n7186), .ZN(n11174) );
  NAND2_X1 U8419 ( .A1(n11736), .A2(n11735), .ZN(n11738) );
  AND4_X2 U8420 ( .A1(n8431), .A2(n8430), .A3(n8429), .A4(n8428), .ZN(n15062)
         );
  NAND2_X1 U8421 ( .A1(n8457), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8431) );
  CLKBUF_X1 U8422 ( .A(n10780), .Z(n15060) );
  OR2_X1 U8423 ( .A1(n10570), .A2(n10550), .ZN(n12433) );
  AND4_X1 U8424 ( .A1(n8525), .A2(n8524), .A3(n8523), .A4(n8522), .ZN(n11569)
         );
  AND2_X1 U8425 ( .A1(n8811), .A2(n8810), .ZN(n12422) );
  NAND2_X1 U8426 ( .A1(n10545), .A2(n15056), .ZN(n12424) );
  AOI22_X1 U8427 ( .A1(n12344), .A2(n12345), .B1(n12614), .B2(n12283), .ZN(
        n12416) );
  OAI21_X1 U8428 ( .B1(n11979), .B2(n7202), .A(n7205), .ZN(n12252) );
  NAND2_X1 U8429 ( .A1(n7207), .A2(n7203), .ZN(n7202) );
  AND2_X1 U8430 ( .A1(n8838), .A2(n8837), .ZN(n12327) );
  INV_X1 U8431 ( .A(n12643), .ZN(n12444) );
  OR2_X1 U8432 ( .A1(n10537), .A2(n10208), .ZN(n12443) );
  INV_X1 U8433 ( .A(n12357), .ZN(n12724) );
  INV_X1 U8434 ( .A(n11569), .ZN(n11562) );
  INV_X1 U8435 ( .A(n11377), .ZN(n12449) );
  NAND2_X1 U8436 ( .A1(n8457), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8424) );
  INV_X1 U8437 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14910) );
  AOI22_X1 U8438 ( .A1(n10505), .A2(n14907), .B1(n9071), .B2(n8437), .ZN(
        n10456) );
  OR2_X1 U8439 ( .A1(n7016), .A2(n9036), .ZN(n14913) );
  OR3_X1 U8440 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n8464) );
  NAND2_X1 U8441 ( .A1(n10463), .A2(n10464), .ZN(n10462) );
  INV_X1 U8442 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n14948) );
  INV_X1 U8443 ( .A(n9040), .ZN(n9039) );
  INV_X1 U8444 ( .A(n6997), .ZN(n14927) );
  OAI21_X1 U8445 ( .B1(n14930), .B2(n10794), .A(n10793), .ZN(n10796) );
  NOR2_X1 U8446 ( .A1(n15003), .A2(n15004), .ZN(n15002) );
  NAND2_X1 U8447 ( .A1(n9099), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7063) );
  NAND2_X1 U8448 ( .A1(n9149), .A2(n9099), .ZN(n7062) );
  OR2_X1 U8449 ( .A1(n14434), .A2(n14435), .ZN(n7013) );
  AND2_X1 U8450 ( .A1(P3_U3897), .A2(n12029), .ZN(n14963) );
  NAND2_X1 U8451 ( .A1(n7009), .A2(n7008), .ZN(n12488) );
  NOR2_X1 U8452 ( .A1(n9903), .A2(n9902), .ZN(n9904) );
  NOR2_X1 U8453 ( .A1(n12442), .A2(n15061), .ZN(n9903) );
  AND2_X1 U8454 ( .A1(n8789), .A2(n8788), .ZN(n12591) );
  NAND2_X1 U8455 ( .A1(n6899), .A2(n6900), .ZN(n12598) );
  NAND2_X1 U8456 ( .A1(n6870), .A2(n6874), .ZN(n12640) );
  NAND2_X1 U8457 ( .A1(n12662), .A2(n6467), .ZN(n6870) );
  AND2_X1 U8458 ( .A1(n6875), .A2(n6878), .ZN(n12651) );
  NAND2_X1 U8459 ( .A1(n12662), .A2(n12668), .ZN(n6875) );
  NAND2_X1 U8460 ( .A1(n12665), .A2(n8951), .ZN(n12656) );
  NAND2_X1 U8461 ( .A1(n12699), .A2(n8855), .ZN(n12679) );
  AND2_X1 U8462 ( .A1(n8686), .A2(n8685), .ZN(n12793) );
  CLKBUF_X1 U8463 ( .A(n12727), .Z(n12729) );
  OAI21_X1 U8464 ( .B1(n8550), .B2(n6787), .A(n6784), .ZN(n14456) );
  NAND2_X1 U8465 ( .A1(n11313), .A2(n6886), .ZN(n15042) );
  NAND2_X1 U8466 ( .A1(n15048), .A2(n15084), .ZN(n12744) );
  NAND2_X1 U8467 ( .A1(n10819), .A2(n15056), .ZN(n15094) );
  AND2_X1 U8468 ( .A1(n15094), .A2(n15069), .ZN(n15091) );
  AND2_X2 U8469 ( .A1(n10573), .A2(n10544), .ZN(n15090) );
  AOI21_X1 U8470 ( .B1(n12244), .B2(n8828), .A(n8415), .ZN(n12753) );
  NOR2_X1 U8471 ( .A1(n12558), .A2(n12817), .ZN(n9895) );
  INV_X1 U8472 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10503) );
  INV_X1 U8473 ( .A(n9910), .ZN(n12548) );
  AND2_X1 U8474 ( .A1(n8763), .A2(n8762), .ZN(n12838) );
  INV_X1 U8475 ( .A(n12403), .ZN(n12846) );
  INV_X1 U8476 ( .A(n12341), .ZN(n12850) );
  AND2_X1 U8477 ( .A1(n12800), .A2(n12799), .ZN(n12854) );
  NAND2_X1 U8478 ( .A1(n8609), .A2(n8608), .ZN(n12870) );
  INV_X1 U8479 ( .A(n10818), .ZN(n10582) );
  INV_X1 U8480 ( .A(n10542), .ZN(n10208) );
  NAND2_X1 U8481 ( .A1(n9022), .A2(n9025), .ZN(n11955) );
  XNOR2_X1 U8482 ( .A(n9019), .B(n9018), .ZN(n11908) );
  INV_X1 U8483 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n9018) );
  OAI21_X1 U8484 ( .B1(n6462), .B2(P3_IR_REG_24__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9019) );
  XNOR2_X1 U8485 ( .A(n9021), .B(n9020), .ZN(n9849) );
  INV_X1 U8486 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n9020) );
  NAND2_X1 U8487 ( .A1(n6462), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9021) );
  OAI21_X1 U8488 ( .B1(n8725), .B2(n7147), .A(n7144), .ZN(n8750) );
  NAND2_X1 U8489 ( .A1(n8737), .A2(n8736), .ZN(n8735) );
  NAND2_X1 U8490 ( .A1(n8725), .A2(n8340), .ZN(n8737) );
  INV_X1 U8491 ( .A(n10832), .ZN(n11360) );
  INV_X1 U8492 ( .A(SI_20_), .ZN(n11210) );
  NAND2_X1 U8493 ( .A1(n8694), .A2(n8337), .ZN(n8710) );
  XNOR2_X1 U8494 ( .A(n8843), .B(n7198), .ZN(n11211) );
  NAND2_X1 U8495 ( .A1(n8647), .A2(n8331), .ZN(n8665) );
  INV_X1 U8496 ( .A(SI_16_), .ZN(n10587) );
  INV_X1 U8497 ( .A(n9154), .ZN(n12497) );
  INV_X1 U8498 ( .A(SI_15_), .ZN(n10441) );
  NAND2_X1 U8499 ( .A1(n7126), .A2(n7127), .ZN(n8631) );
  AND2_X1 U8500 ( .A1(n7123), .A2(n6546), .ZN(n7127) );
  INV_X1 U8501 ( .A(SI_14_), .ZN(n10321) );
  NAND2_X1 U8502 ( .A1(n8606), .A2(n8326), .ZN(n8618) );
  NAND2_X1 U8503 ( .A1(n8322), .A2(n8321), .ZN(n8578) );
  XNOR2_X1 U8504 ( .A(n8568), .B(n8567), .ZN(n14973) );
  INV_X1 U8505 ( .A(n9139), .ZN(n10993) );
  OAI21_X1 U8506 ( .B1(n8493), .B2(n7136), .A(n7135), .ZN(n8527) );
  INV_X1 U8507 ( .A(n14942), .ZN(n10035) );
  NAND2_X1 U8508 ( .A1(n8496), .A2(n8312), .ZN(n8517) );
  NAND2_X1 U8509 ( .A1(n7156), .A2(n8306), .ZN(n8475) );
  NAND2_X1 U8510 ( .A1(n7152), .A2(n7149), .ZN(n8463) );
  INV_X1 U8511 ( .A(n7151), .ZN(n7149) );
  NAND2_X1 U8512 ( .A1(n8304), .A2(n8303), .ZN(n8447) );
  MUX2_X1 U8513 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8434), .S(
        P3_IR_REG_1__SCAN_IN), .Z(n8436) );
  INV_X1 U8514 ( .A(SI_1_), .ZN(n7369) );
  NAND2_X1 U8515 ( .A1(n12983), .A2(n7224), .ZN(n12885) );
  OAI21_X1 U8516 ( .B1(n12937), .B2(n6676), .A(n6673), .ZN(n6681) );
  NAND2_X1 U8517 ( .A1(n11155), .A2(n7590), .ZN(n11452) );
  NAND2_X1 U8518 ( .A1(n7602), .A2(n7601), .ZN(n11500) );
  AOI21_X1 U8519 ( .B1(n6687), .B2(n6686), .A(n6453), .ZN(n6685) );
  AND2_X1 U8520 ( .A1(n8037), .A2(n8036), .ZN(n12992) );
  AOI21_X1 U8521 ( .B1(n7224), .B2(n7223), .A(n7969), .ZN(n7222) );
  INV_X1 U8522 ( .A(n6489), .ZN(n7223) );
  AND2_X1 U8523 ( .A1(n12219), .A2(n7567), .ZN(n7568) );
  NAND2_X1 U8524 ( .A1(n7559), .A2(n7558), .ZN(n14881) );
  AND2_X1 U8525 ( .A1(n12942), .A2(n7825), .ZN(n12918) );
  NAND2_X1 U8526 ( .A1(n12210), .A2(n7635), .ZN(n11652) );
  NAND2_X1 U8527 ( .A1(n11854), .A2(n7721), .ZN(n11968) );
  NAND2_X1 U8528 ( .A1(n7757), .A2(n11960), .ZN(n11966) );
  NAND2_X1 U8529 ( .A1(n12937), .A2(n12936), .ZN(n12935) );
  INV_X1 U8530 ( .A(n10018), .ZN(n10668) );
  NAND2_X1 U8531 ( .A1(n12902), .A2(n12903), .ZN(n12944) );
  NAND2_X1 U8532 ( .A1(n11651), .A2(n11653), .ZN(n11668) );
  NAND2_X1 U8533 ( .A1(n11966), .A2(n7761), .ZN(n12972) );
  AND2_X1 U8534 ( .A1(n7523), .A2(n7524), .ZN(n10765) );
  NAND2_X1 U8535 ( .A1(n10667), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12990) );
  INV_X1 U8536 ( .A(n12971), .ZN(n12996) );
  INV_X1 U8537 ( .A(n12978), .ZN(n12953) );
  NAND2_X1 U8538 ( .A1(n8291), .A2(n12034), .ZN(n6744) );
  INV_X1 U8539 ( .A(n12889), .ZN(n13003) );
  INV_X1 U8540 ( .A(n12979), .ZN(n13006) );
  INV_X1 U8541 ( .A(n12924), .ZN(n13007) );
  INV_X1 U8542 ( .A(n12959), .ZN(n13008) );
  NAND2_X1 U8543 ( .A1(n8204), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7406) );
  OR2_X1 U8544 ( .A1(n13077), .A2(n7799), .ZN(n13292) );
  OR3_X1 U8545 ( .A1(n13114), .A2(n13113), .A3(n7799), .ZN(n13312) );
  AND2_X1 U8546 ( .A1(n7979), .A2(n7962), .ZN(n13115) );
  INV_X1 U8547 ( .A(n13318), .ZN(n13129) );
  OR2_X1 U8548 ( .A1(n11816), .A2(n8235), .ZN(n7857) );
  NAND2_X1 U8549 ( .A1(n13211), .A2(n9997), .ZN(n13204) );
  NAND2_X1 U8550 ( .A1(n7024), .A2(n7028), .ZN(n13197) );
  NAND2_X1 U8551 ( .A1(n13226), .A2(n7031), .ZN(n7024) );
  OAI21_X1 U8552 ( .B1(n13226), .B2(n6470), .A(n9940), .ZN(n13210) );
  CLKBUF_X1 U8553 ( .A(n13242), .Z(n13243) );
  NAND2_X1 U8554 ( .A1(n7045), .A2(n7050), .ZN(n13267) );
  NAND2_X1 U8555 ( .A1(n11903), .A2(n7051), .ZN(n7045) );
  NAND2_X1 U8556 ( .A1(n7732), .A2(n7731), .ZN(n13285) );
  NAND2_X1 U8557 ( .A1(n6841), .A2(n6840), .ZN(n11894) );
  INV_X1 U8558 ( .A(n11666), .ZN(n10019) );
  NAND2_X1 U8559 ( .A1(n6838), .A2(n9971), .ZN(n11163) );
  NAND2_X1 U8560 ( .A1(n10975), .A2(n9969), .ZN(n6838) );
  NAND2_X1 U8561 ( .A1(n14868), .A2(n10023), .ZN(n14853) );
  INV_X1 U8562 ( .A(n14847), .ZN(n13221) );
  AND2_X1 U8563 ( .A1(n14868), .A2(n12239), .ZN(n14847) );
  INV_X1 U8564 ( .A(n14853), .ZN(n14479) );
  NAND2_X1 U8565 ( .A1(n14880), .A2(n8023), .ZN(n14863) );
  INV_X1 U8566 ( .A(n13086), .ZN(n13382) );
  INV_X1 U8567 ( .A(n10001), .ZN(n13394) );
  INV_X1 U8568 ( .A(n13229), .ZN(n10020) );
  NAND2_X1 U8569 ( .A1(n7578), .A2(n7577), .ZN(n11543) );
  OR2_X1 U8570 ( .A1(n10075), .A2(n8235), .ZN(n6690) );
  AND2_X1 U8571 ( .A1(n8041), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14880) );
  XNOR2_X1 U8572 ( .A(n7999), .B(P2_IR_REG_26__SCAN_IN), .ZN(n13434) );
  OAI21_X1 U8573 ( .B1(n7998), .B2(P2_IR_REG_25__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7999) );
  AND2_X1 U8574 ( .A1(n7995), .A2(n7998), .ZN(n12015) );
  OR2_X1 U8575 ( .A1(n7992), .A2(n7677), .ZN(n7381) );
  OR2_X1 U8576 ( .A1(n7382), .A2(n7677), .ZN(n7384) );
  XNOR2_X1 U8577 ( .A(n7387), .B(n7386), .ZN(n11532) );
  INV_X1 U8578 ( .A(n8022), .ZN(n12239) );
  INV_X1 U8579 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n14112) );
  INV_X1 U8580 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n14123) );
  INV_X1 U8581 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10982) );
  INV_X1 U8582 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10283) );
  INV_X1 U8583 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10094) );
  INV_X1 U8584 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10090) );
  INV_X1 U8585 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10078) );
  INV_X1 U8586 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10083) );
  INV_X1 U8587 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10076) );
  NOR2_X1 U8588 ( .A1(n10049), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13433) );
  NAND2_X1 U8589 ( .A1(n6989), .A2(n11212), .ZN(n6988) );
  NAND2_X1 U8590 ( .A1(n6992), .A2(n12003), .ZN(n12006) );
  INV_X1 U8591 ( .A(n6957), .ZN(n6956) );
  OAI21_X1 U8592 ( .B1(n6468), .B2(n6959), .A(n6958), .ZN(n6957) );
  INV_X1 U8593 ( .A(n6975), .ZN(n6971) );
  NAND2_X1 U8594 ( .A1(n10718), .A2(n7344), .ZN(n10717) );
  NAND2_X1 U8595 ( .A1(n6967), .A2(n6968), .ZN(n13463) );
  AOI21_X1 U8596 ( .B1(n13481), .B2(n13491), .A(n13490), .ZN(n13493) );
  NAND2_X1 U8597 ( .A1(n11787), .A2(n11786), .ZN(n11790) );
  OR2_X1 U8598 ( .A1(n10606), .A2(n10590), .ZN(n13540) );
  NAND2_X1 U8599 ( .A1(n6982), .A2(n6983), .ZN(n13528) );
  OR2_X1 U8600 ( .A1(n10606), .A2(n10605), .ZN(n13557) );
  XNOR2_X1 U8601 ( .A(n12052), .B(n12054), .ZN(n13548) );
  AND2_X1 U8602 ( .A1(n13529), .A2(n14669), .ZN(n13555) );
  OR3_X1 U8603 ( .A1(n9700), .A2(n9699), .A3(n9698), .ZN(n13699) );
  NOR2_X1 U8604 ( .A1(n10413), .A2(n10412), .ZN(n13635) );
  NAND2_X1 U8605 ( .A1(n13626), .A2(n6611), .ZN(n10413) );
  NAND2_X1 U8606 ( .A1(n6613), .A2(n6612), .ZN(n6611) );
  NOR2_X1 U8607 ( .A1(n10423), .A2(n6615), .ZN(n10424) );
  AND2_X1 U8608 ( .A1(n10426), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6615) );
  NAND2_X1 U8609 ( .A1(n10424), .A2(n10425), .ZN(n10528) );
  AOI21_X1 U8610 ( .B1(n10528), .B2(n10526), .A(n10527), .ZN(n10923) );
  NOR2_X1 U8611 ( .A1(n10923), .A2(n6614), .ZN(n14600) );
  AND2_X1 U8612 ( .A1(n10931), .A2(n10525), .ZN(n6614) );
  INV_X1 U8613 ( .A(n6616), .ZN(n11694) );
  INV_X1 U8614 ( .A(n6820), .ZN(n13702) );
  INV_X1 U8615 ( .A(n6626), .ZN(n6625) );
  OAI21_X1 U8616 ( .B1(n7313), .B2(n6630), .A(n6627), .ZN(n6626) );
  NAND2_X1 U8617 ( .A1(n13754), .A2(n6628), .ZN(n6627) );
  INV_X1 U8618 ( .A(n13732), .ZN(n6628) );
  AND2_X1 U8619 ( .A1(n7313), .A2(n13754), .ZN(n6629) );
  AOI21_X1 U8620 ( .B1(n13778), .B2(n14708), .A(n13777), .ZN(n14030) );
  NAND2_X1 U8621 ( .A1(n13776), .A2(n13775), .ZN(n13777) );
  OAI21_X1 U8622 ( .B1(n6700), .B2(n6703), .A(n6508), .ZN(n13792) );
  NAND2_X1 U8623 ( .A1(n13848), .A2(n13726), .ZN(n13836) );
  NAND2_X1 U8624 ( .A1(n13848), .A2(n7315), .ZN(n13834) );
  NAND2_X1 U8625 ( .A1(n6944), .A2(n6945), .ZN(n13823) );
  INV_X1 U8626 ( .A(n6831), .ZN(n13845) );
  NAND2_X1 U8627 ( .A1(n6948), .A2(n6947), .ZN(n13839) );
  AND2_X1 U8628 ( .A1(n6948), .A2(n6479), .ZN(n13840) );
  AND2_X1 U8629 ( .A1(n13908), .A2(n13718), .ZN(n13898) );
  AND2_X1 U8630 ( .A1(n6950), .A2(n13742), .ZN(n13902) );
  NAND2_X1 U8631 ( .A1(n13934), .A2(n13741), .ZN(n13927) );
  AND2_X1 U8632 ( .A1(n9496), .A2(n9495), .ZN(n13977) );
  NAND2_X1 U8633 ( .A1(n9433), .A2(n9432), .ZN(n14528) );
  INV_X1 U8634 ( .A(n6643), .ZN(n6647) );
  OAI21_X1 U8635 ( .B1(n11833), .B2(n6904), .A(n6903), .ZN(n13734) );
  NAND2_X1 U8636 ( .A1(n11715), .A2(n11714), .ZN(n7303) );
  NAND2_X1 U8637 ( .A1(n9410), .A2(n9409), .ZN(n11884) );
  AND3_X1 U8638 ( .A1(n6936), .A2(n6933), .A3(n6443), .ZN(n11441) );
  NAND2_X1 U8639 ( .A1(n6922), .A2(n6920), .ZN(n14612) );
  AOI21_X1 U8640 ( .B1(n6924), .B2(n6925), .A(n6923), .ZN(n6922) );
  NAND2_X1 U8641 ( .A1(n6926), .A2(n6927), .ZN(n11296) );
  NAND2_X1 U8642 ( .A1(n11056), .A2(n11055), .ZN(n13913) );
  INV_X1 U8643 ( .A(n14002), .ZN(n14634) );
  INV_X1 U8644 ( .A(n14643), .ZN(n14623) );
  NAND2_X1 U8645 ( .A1(n7334), .A2(n11071), .ZN(n11258) );
  INV_X1 U8646 ( .A(n14008), .ZN(n13967) );
  AND4_X2 U8647 ( .A1(n10314), .A2(n10748), .A3(n10747), .A4(n13761), .ZN(
        n14745) );
  OR2_X1 U8648 ( .A1(n14042), .A2(n14041), .ZN(n14249) );
  XNOR2_X1 U8649 ( .A(n8201), .B(n8200), .ZN(n14268) );
  NAND2_X1 U8650 ( .A1(n8234), .A2(n8198), .ZN(n8201) );
  NAND2_X1 U8651 ( .A1(n6910), .A2(n6909), .ZN(n6908) );
  NAND2_X1 U8652 ( .A1(n9179), .A2(n6911), .ZN(n6905) );
  OR2_X1 U8653 ( .A1(n9179), .A2(n6912), .ZN(n6906) );
  NAND2_X1 U8654 ( .A1(n8234), .A2(n8233), .ZN(n14272) );
  CLKBUF_X1 U8655 ( .A(n9783), .Z(n6588) );
  NAND2_X1 U8656 ( .A1(n7891), .A2(n7874), .ZN(n12038) );
  NAND2_X1 U8657 ( .A1(n9767), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7277) );
  OR2_X1 U8658 ( .A1(n7255), .A2(n7256), .ZN(n7827) );
  INV_X1 U8659 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11171) );
  INV_X1 U8660 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n14181) );
  INV_X1 U8661 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10894) );
  INV_X1 U8662 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10646) );
  INV_X1 U8663 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10443) );
  INV_X1 U8664 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10461) );
  INV_X1 U8665 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10284) );
  AND2_X1 U8666 ( .A1(n9357), .A2(n9374), .ZN(n13656) );
  INV_X1 U8667 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10095) );
  INV_X1 U8668 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10092) );
  NAND2_X1 U8669 ( .A1(n7526), .A2(n7525), .ZN(n7530) );
  INV_X1 U8670 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10061) );
  INV_X1 U8671 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10063) );
  CLKBUF_X1 U8672 ( .A(n9248), .Z(n9249) );
  NOR2_X1 U8673 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n9234) );
  XNOR2_X1 U8674 ( .A(n9218), .B(n9219), .ZN(n13577) );
  CLKBUF_X1 U8675 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n14284) );
  XNOR2_X1 U8676 ( .A(n14331), .B(n6671), .ZN(n15179) );
  INV_X1 U8677 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6671) );
  XNOR2_X1 U8678 ( .A(n14346), .B(n7058), .ZN(n14401) );
  INV_X1 U8679 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7058) );
  XNOR2_X1 U8680 ( .A(n14351), .B(n7057), .ZN(n15172) );
  AOI21_X1 U8681 ( .B1(n14361), .B2(n14360), .A(n14407), .ZN(n14554) );
  AOI21_X1 U8682 ( .B1(n14383), .B2(n14382), .A(n14567), .ZN(n14420) );
  OAI21_X1 U8683 ( .B1(n9013), .B2(n7166), .A(n9016), .ZN(n9029) );
  INV_X1 U8684 ( .A(n7020), .ZN(n14986) );
  AND2_X1 U8685 ( .A1(n7076), .A2(n7074), .ZN(n12537) );
  INV_X1 U8686 ( .A(n6995), .ZN(n12523) );
  AND2_X1 U8687 ( .A1(n9120), .A2(n9119), .ZN(n7339) );
  NAND2_X1 U8688 ( .A1(n12289), .A2(n12748), .ZN(n6580) );
  OAI21_X1 U8689 ( .B1(n12558), .B2(n12871), .A(n9874), .ZN(n9875) );
  NAND2_X1 U8690 ( .A1(n12289), .A2(n12821), .ZN(n6581) );
  OAI21_X1 U8691 ( .B1(n11651), .B2(n7220), .A(n7217), .ZN(n12196) );
  OR2_X1 U8692 ( .A1(n6746), .A2(n6741), .ZN(n6740) );
  INV_X1 U8693 ( .A(n10030), .ZN(n10031) );
  NAND2_X1 U8694 ( .A1(n13116), .A2(n13351), .ZN(n6583) );
  NAND2_X1 U8695 ( .A1(n13116), .A2(n13407), .ZN(n6582) );
  OAI211_X1 U8696 ( .C1(n13692), .C2(n13691), .A(n13694), .B(n6617), .ZN(
        P1_U3262) );
  NAND2_X1 U8697 ( .A1(n6618), .A2(n13691), .ZN(n6617) );
  NOR2_X1 U8698 ( .A1(n14405), .A2(n14404), .ZN(n14403) );
  AND2_X1 U8699 ( .A1(n6670), .A2(n6475), .ZN(n14405) );
  INV_X1 U8700 ( .A(n7040), .ZN(n14556) );
  NAND2_X1 U8701 ( .A1(n6661), .A2(n6662), .ZN(n14562) );
  NOR2_X1 U8702 ( .A1(n6658), .A2(n6656), .ZN(n14560) );
  XNOR2_X1 U8703 ( .A(n6652), .B(n6542), .ZN(SUB_1596_U4) );
  OAI21_X1 U8704 ( .B1(n14423), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n6481), .ZN(
        n6652) );
  OR2_X2 U8705 ( .A1(n11535), .A2(n11598), .ZN(n8096) );
  INV_X2 U8706 ( .A(n8061), .ZN(n8262) );
  AND2_X1 U8707 ( .A1(n11481), .A2(n6828), .ZN(n6436) );
  INV_X2 U8708 ( .A(n8096), .ZN(n8074) );
  AND2_X1 U8709 ( .A1(n6436), .A2(n6827), .ZN(n6437) );
  AND2_X1 U8710 ( .A1(n8185), .A2(n8184), .ZN(n6438) );
  INV_X1 U8711 ( .A(n11290), .ZN(n7298) );
  AND2_X1 U8712 ( .A1(n6422), .A2(n8478), .ZN(n6439) );
  AND2_X1 U8713 ( .A1(n7787), .A2(n7237), .ZN(n6440) );
  NAND2_X1 U8714 ( .A1(n9130), .A2(n10054), .ZN(n6441) );
  INV_X1 U8715 ( .A(n12171), .ZN(n6758) );
  INV_X1 U8716 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7007) );
  XNOR2_X1 U8717 ( .A(n7653), .B(SI_12_), .ZN(n7655) );
  INV_X1 U8718 ( .A(n7655), .ZN(n6732) );
  INV_X1 U8719 ( .A(n14020), .ZN(n13758) );
  OR2_X1 U8720 ( .A1(n13758), .A2(n13707), .ZN(n6442) );
  NAND2_X1 U8721 ( .A1(n14557), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n6662) );
  INV_X1 U8722 ( .A(n6662), .ZN(n6660) );
  NAND2_X1 U8723 ( .A1(n11594), .A2(n11582), .ZN(n6443) );
  INV_X1 U8724 ( .A(n11294), .ZN(n6923) );
  NOR2_X1 U8725 ( .A1(n13452), .A2(n13453), .ZN(n6444) );
  NOR2_X1 U8726 ( .A1(n14561), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n6445) );
  XNOR2_X1 U8727 ( .A(n14058), .B(n13746), .ZN(n13863) );
  INV_X1 U8728 ( .A(n7029), .ZN(n7028) );
  OAI22_X1 U8729 ( .A1(n9941), .A2(n7030), .B1(n13011), .B2(n13406), .ZN(n7029) );
  OR2_X1 U8730 ( .A1(n13939), .A2(n13935), .ZN(n6446) );
  INV_X1 U8731 ( .A(n9948), .ZN(n13109) );
  AND2_X1 U8732 ( .A1(n6882), .A2(n6883), .ZN(n12707) );
  AND4_X1 U8733 ( .A1(n6595), .A2(n7614), .A3(n7459), .A4(n7509), .ZN(n6447)
         );
  AND2_X1 U8734 ( .A1(n11440), .A2(n6443), .ZN(n6448) );
  AND2_X1 U8735 ( .A1(n13135), .A2(n6852), .ZN(n6449) );
  AND2_X1 U8736 ( .A1(n12534), .A2(n12533), .ZN(n6450) );
  NAND2_X1 U8737 ( .A1(n8175), .A2(n7121), .ZN(n6451) );
  INV_X1 U8738 ( .A(n6703), .ZN(n6702) );
  OAI21_X1 U8739 ( .B1(n6942), .B2(n7254), .A(n6704), .ZN(n6703) );
  OAI21_X1 U8740 ( .B1(n6737), .B2(n6732), .A(n6509), .ZN(n6735) );
  NAND2_X1 U8741 ( .A1(n7161), .A2(n6545), .ZN(n6452) );
  AND2_X1 U8742 ( .A1(n7783), .A2(n7782), .ZN(n6453) );
  AND2_X1 U8743 ( .A1(n14661), .A2(n11190), .ZN(n6454) );
  AND2_X1 U8744 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n7139), .ZN(n6455) );
  XNOR2_X1 U8745 ( .A(n12369), .B(n6538), .ZN(n12370) );
  AND2_X1 U8746 ( .A1(n6772), .A2(n6771), .ZN(n6456) );
  AND2_X1 U8747 ( .A1(n9811), .A2(n9809), .ZN(n6457) );
  AND2_X1 U8748 ( .A1(n11788), .A2(n11786), .ZN(n6458) );
  OR2_X1 U8749 ( .A1(n11469), .A2(n13566), .ZN(n6459) );
  OR2_X1 U8750 ( .A1(n7209), .A2(n6544), .ZN(n12388) );
  INV_X1 U8751 ( .A(n12264), .ZN(n7195) );
  AND2_X1 U8752 ( .A1(n7958), .A2(n7957), .ZN(n13389) );
  INV_X1 U8753 ( .A(n13389), .ZN(n13116) );
  NAND2_X1 U8754 ( .A1(n11803), .A2(n6472), .ZN(n11939) );
  NOR3_X1 U8755 ( .A1(n13286), .A2(n13265), .A3(n13359), .ZN(n13227) );
  AND2_X1 U8756 ( .A1(n6557), .A2(n8321), .ZN(n6460) );
  INV_X1 U8757 ( .A(n12289), .ZN(n12829) );
  NAND2_X1 U8758 ( .A1(n8803), .A2(n8802), .ZN(n12289) );
  NAND2_X1 U8759 ( .A1(n9377), .A2(n9376), .ZN(n11776) );
  INV_X1 U8760 ( .A(n11776), .ZN(n6827) );
  NAND2_X1 U8761 ( .A1(n11625), .A2(n6773), .ZN(n6774) );
  NAND2_X1 U8762 ( .A1(n7196), .A2(n6439), .ZN(n6461) );
  INV_X1 U8763 ( .A(n13791), .ZN(n6699) );
  OR2_X1 U8764 ( .A1(n6461), .A2(n7181), .ZN(n6462) );
  INV_X1 U8765 ( .A(n7447), .ZN(n7555) );
  INV_X1 U8766 ( .A(n10039), .ZN(n7079) );
  INV_X1 U8767 ( .A(n8455), .ZN(n8707) );
  AND2_X1 U8768 ( .A1(n10599), .A2(n10598), .ZN(n6463) );
  OR2_X1 U8769 ( .A1(n13398), .A2(n13007), .ZN(n6464) );
  INV_X1 U8770 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n14263) );
  AND2_X1 U8771 ( .A1(n7857), .A2(n7856), .ZN(n13192) );
  INV_X1 U8772 ( .A(n13192), .ZN(n6770) );
  AND2_X1 U8773 ( .A1(n7977), .A2(n7976), .ZN(n13306) );
  AND2_X1 U8774 ( .A1(n6982), .A2(n6979), .ZN(n6465) );
  NOR2_X1 U8775 ( .A1(n13142), .A2(n13141), .ZN(n6466) );
  INV_X1 U8776 ( .A(n11293), .ZN(n6819) );
  AND2_X1 U8777 ( .A1(n6877), .A2(n12668), .ZN(n6467) );
  INV_X1 U8778 ( .A(n6787), .ZN(n6786) );
  NAND2_X1 U8779 ( .A1(n8562), .A2(n8903), .ZN(n6787) );
  AND2_X1 U8780 ( .A1(n13518), .A2(n6961), .ZN(n6468) );
  AND2_X1 U8781 ( .A1(n13212), .A2(n9995), .ZN(n6469) );
  NOR2_X1 U8782 ( .A1(n13229), .A2(n13012), .ZN(n6470) );
  AND2_X1 U8783 ( .A1(n7427), .A2(n7345), .ZN(n7448) );
  AND2_X1 U8784 ( .A1(n14579), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6471) );
  AND2_X1 U8785 ( .A1(n11802), .A2(n11804), .ZN(n6472) );
  INV_X1 U8786 ( .A(n9122), .ZN(n9121) );
  OR2_X1 U8787 ( .A1(n11469), .A2(n11467), .ZN(n6473) );
  OR2_X1 U8788 ( .A1(n7654), .A2(SI_12_), .ZN(n6474) );
  AND2_X1 U8789 ( .A1(n7902), .A2(n7901), .ZN(n13398) );
  AND2_X1 U8790 ( .A1(n7749), .A2(n7748), .ZN(n13416) );
  INV_X1 U8791 ( .A(n13416), .ZN(n13265) );
  AND2_X1 U8792 ( .A1(n7317), .A2(n6993), .ZN(n9204) );
  NAND2_X1 U8793 ( .A1(n7746), .A2(n7745), .ZN(n7763) );
  NAND2_X1 U8794 ( .A1(n13896), .A2(n13719), .ZN(n13872) );
  OR2_X1 U8795 ( .A1(n14355), .A2(n14354), .ZN(n6475) );
  INV_X1 U8796 ( .A(n7638), .ZN(n6729) );
  NAND2_X1 U8797 ( .A1(n6446), .A2(n13716), .ZN(n13920) );
  AND2_X1 U8798 ( .A1(n6893), .A2(n6896), .ZN(n6476) );
  INV_X1 U8799 ( .A(n13928), .ZN(n7312) );
  AND2_X1 U8800 ( .A1(n6702), .A2(n13791), .ZN(n6477) );
  INV_X1 U8801 ( .A(n11168), .ZN(n6839) );
  INV_X1 U8802 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9445) );
  OAI21_X1 U8803 ( .B1(n9905), .B2(n12736), .A(n9904), .ZN(n12547) );
  AND2_X1 U8804 ( .A1(n8254), .A2(n8222), .ZN(n6478) );
  NAND2_X1 U8805 ( .A1(n14058), .A2(n13746), .ZN(n6479) );
  NAND2_X1 U8806 ( .A1(n7317), .A2(n7287), .ZN(n9207) );
  INV_X1 U8807 ( .A(n8123), .ZN(n7102) );
  INV_X1 U8808 ( .A(n8115), .ZN(n7091) );
  INV_X1 U8809 ( .A(n8095), .ZN(n7108) );
  INV_X1 U8810 ( .A(n9312), .ZN(n7286) );
  INV_X1 U8811 ( .A(n8126), .ZN(n7100) );
  INV_X1 U8812 ( .A(n8099), .ZN(n7106) );
  OR2_X1 U8813 ( .A1(n6461), .A2(n7180), .ZN(n6480) );
  INV_X1 U8814 ( .A(n7639), .ZN(n6692) );
  NAND2_X1 U8815 ( .A1(n7619), .A2(n7618), .ZN(n12208) );
  OR2_X1 U8816 ( .A1(n14425), .A2(n14424), .ZN(n6481) );
  INV_X1 U8817 ( .A(n8966), .ZN(n6802) );
  AND2_X1 U8818 ( .A1(n8899), .A2(n8900), .ZN(n11317) );
  AND2_X1 U8819 ( .A1(n14045), .A2(n13728), .ZN(n6482) );
  AND2_X1 U8820 ( .A1(n11173), .A2(n11176), .ZN(n6483) );
  NOR2_X1 U8821 ( .A1(n14438), .A2(n9152), .ZN(n6484) );
  INV_X1 U8822 ( .A(n6707), .ZN(n6706) );
  NOR2_X1 U8823 ( .A1(n13750), .A2(n13749), .ZN(n6707) );
  INV_X1 U8824 ( .A(n6694), .ZN(n13772) );
  NOR2_X1 U8825 ( .A1(n8170), .A2(n8171), .ZN(n6485) );
  INV_X1 U8826 ( .A(n8078), .ZN(n7094) );
  INV_X1 U8827 ( .A(n7137), .ZN(n7136) );
  NOR2_X1 U8828 ( .A1(n8313), .A2(n7138), .ZN(n7137) );
  AND2_X1 U8829 ( .A1(n7822), .A2(n12903), .ZN(n6486) );
  INV_X1 U8830 ( .A(n9412), .ZN(n7280) );
  INV_X1 U8831 ( .A(n6680), .ZN(n6679) );
  NAND2_X1 U8832 ( .A1(n6682), .A2(n12936), .ZN(n6680) );
  OR2_X1 U8833 ( .A1(n8173), .A2(n8174), .ZN(n6487) );
  AND2_X1 U8834 ( .A1(n13285), .A2(n13015), .ZN(n6488) );
  NOR2_X1 U8835 ( .A1(n12982), .A2(n7948), .ZN(n6489) );
  OR2_X1 U8836 ( .A1(n9683), .A2(n9682), .ZN(n6490) );
  AND2_X1 U8837 ( .A1(n9686), .A2(n9685), .ZN(n14016) );
  AND2_X1 U8838 ( .A1(n13714), .A2(n9482), .ZN(n13713) );
  AND2_X1 U8839 ( .A1(n6438), .A2(n6487), .ZN(n6491) );
  AND2_X1 U8840 ( .A1(n6475), .A2(n6669), .ZN(n6492) );
  OR2_X1 U8841 ( .A1(n6659), .A2(n6657), .ZN(n6493) );
  INV_X1 U8842 ( .A(n11429), .ZN(n11438) );
  INV_X1 U8843 ( .A(n9947), .ZN(n7038) );
  NOR2_X1 U8844 ( .A1(n14221), .A2(n13903), .ZN(n6494) );
  NOR2_X1 U8845 ( .A1(n13344), .A2(n13010), .ZN(n6495) );
  NOR2_X1 U8846 ( .A1(n12846), .A2(n12654), .ZN(n6496) );
  OR2_X1 U8847 ( .A1(n6445), .A2(n6493), .ZN(n6497) );
  OR2_X1 U8848 ( .A1(n8082), .A2(n8084), .ZN(n6498) );
  INV_X1 U8849 ( .A(n6928), .ZN(n6927) );
  NOR2_X1 U8850 ( .A1(n11274), .A2(n11077), .ZN(n6928) );
  AND2_X1 U8851 ( .A1(n7650), .A2(n7651), .ZN(n6499) );
  OR2_X1 U8852 ( .A1(n6461), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n6500) );
  INV_X1 U8853 ( .A(n12687), .ZN(n12696) );
  AND2_X1 U8854 ( .A1(n8855), .A2(n8941), .ZN(n12687) );
  NOR2_X1 U8855 ( .A1(n7091), .A2(n8113), .ZN(n6501) );
  AND2_X1 U8856 ( .A1(n7101), .A2(n7100), .ZN(n6502) );
  AND2_X1 U8857 ( .A1(n7107), .A2(n7106), .ZN(n6503) );
  NOR2_X1 U8858 ( .A1(n14051), .A2(n13747), .ZN(n6504) );
  NAND2_X1 U8859 ( .A1(n12758), .A2(n12570), .ZN(n6505) );
  INV_X1 U8860 ( .A(n7330), .ZN(n6853) );
  NAND2_X1 U8861 ( .A1(n7317), .A2(n9177), .ZN(n6506) );
  AND2_X1 U8862 ( .A1(n7698), .A2(n7697), .ZN(n6507) );
  AND2_X1 U8863 ( .A1(n6701), .A2(n6706), .ZN(n6508) );
  INV_X1 U8864 ( .A(n6825), .ZN(n6824) );
  NAND2_X1 U8865 ( .A1(n13695), .A2(n6826), .ZN(n6825) );
  INV_X1 U8866 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9197) );
  INV_X1 U8867 ( .A(n6964), .ZN(n6963) );
  AOI21_X1 U8868 ( .B1(n6965), .B2(n13509), .A(n13519), .ZN(n6964) );
  AND2_X1 U8869 ( .A1(n6734), .A2(n6474), .ZN(n6509) );
  NAND2_X1 U8870 ( .A1(n9389), .A2(n9388), .ZN(n11797) );
  INV_X1 U8871 ( .A(n6887), .ZN(n6886) );
  NAND2_X1 U8872 ( .A1(n9820), .A2(n9819), .ZN(n6887) );
  INV_X1 U8873 ( .A(n6676), .ZN(n6675) );
  NAND2_X1 U8874 ( .A1(n6489), .A2(n6678), .ZN(n6676) );
  AND2_X1 U8875 ( .A1(n7725), .A2(n10441), .ZN(n6510) );
  INV_X1 U8876 ( .A(n6688), .ZN(n6687) );
  OR2_X1 U8877 ( .A1(n12973), .A2(n6689), .ZN(n6688) );
  AND2_X1 U8878 ( .A1(n7789), .A2(SI_18_), .ZN(n6511) );
  AND2_X1 U8879 ( .A1(n6967), .A2(n6965), .ZN(n13461) );
  AND2_X1 U8880 ( .A1(n6635), .A2(n13811), .ZN(n6512) );
  NAND2_X1 U8881 ( .A1(n6839), .A2(n13024), .ZN(n6513) );
  AND2_X1 U8882 ( .A1(n8445), .A2(n8372), .ZN(n8478) );
  AND2_X1 U8883 ( .A1(n12341), .A2(n12663), .ZN(n6514) );
  NAND2_X1 U8884 ( .A1(n13344), .A2(n12958), .ZN(n6515) );
  INV_X1 U8885 ( .A(n6790), .ZN(n6789) );
  OR2_X1 U8886 ( .A1(n8563), .A2(n6791), .ZN(n6790) );
  INV_X1 U8887 ( .A(n6980), .ZN(n6979) );
  NAND2_X1 U8888 ( .A1(n6983), .A2(n6981), .ZN(n6980) );
  OR2_X1 U8889 ( .A1(n6876), .A2(n6514), .ZN(n6516) );
  INV_X1 U8890 ( .A(n9652), .ZN(n7268) );
  INV_X1 U8891 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10074) );
  INV_X1 U8892 ( .A(n9755), .ZN(n14013) );
  NAND2_X1 U8893 ( .A1(n9718), .A2(n9717), .ZN(n9755) );
  AND2_X1 U8894 ( .A1(n7135), .A2(n7134), .ZN(n6517) );
  AND2_X1 U8895 ( .A1(n6897), .A2(n9842), .ZN(n6518) );
  OR2_X1 U8896 ( .A1(n9143), .A2(n9048), .ZN(n6519) );
  AND2_X1 U8897 ( .A1(n6975), .A2(n12157), .ZN(n6520) );
  NOR3_X1 U8898 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .A3(
        n10820), .ZN(n9032) );
  AND2_X1 U8899 ( .A1(n13258), .A2(n7051), .ZN(n6521) );
  NAND2_X1 U8900 ( .A1(n8403), .A2(n6812), .ZN(n12042) );
  AND2_X1 U8901 ( .A1(n9265), .A2(n9264), .ZN(n14680) );
  INV_X1 U8902 ( .A(n14680), .ZN(n11274) );
  AND2_X1 U8903 ( .A1(n9856), .A2(n10555), .ZN(n6522) );
  INV_X1 U8904 ( .A(n6929), .ZN(n6924) );
  NOR2_X1 U8905 ( .A1(n11078), .A2(n6930), .ZN(n6929) );
  AND2_X1 U8906 ( .A1(n8708), .A2(n8855), .ZN(n6523) );
  AND2_X1 U8907 ( .A1(n9671), .A2(n9670), .ZN(n14020) );
  AND2_X1 U8908 ( .A1(n6444), .A2(n6984), .ZN(n6524) );
  AND2_X1 U8909 ( .A1(n6593), .A2(n9995), .ZN(n6525) );
  OR2_X1 U8910 ( .A1(n7280), .A2(n9411), .ZN(n6526) );
  OR2_X1 U8911 ( .A1(n9345), .A2(n9343), .ZN(n6527) );
  OR2_X1 U8912 ( .A1(n9380), .A2(n9378), .ZN(n6528) );
  AND2_X1 U8913 ( .A1(n8379), .A2(n6901), .ZN(n6529) );
  OR2_X1 U8914 ( .A1(n7286), .A2(n9311), .ZN(n6530) );
  AND2_X1 U8915 ( .A1(n7013), .A2(n7012), .ZN(n6531) );
  AND2_X1 U8916 ( .A1(n7312), .A2(n13741), .ZN(n6532) );
  INV_X1 U8917 ( .A(n13717), .ZN(n13909) );
  OR2_X1 U8918 ( .A1(n8102), .A2(n8104), .ZN(n6533) );
  AND2_X1 U8919 ( .A1(n6853), .A2(n6464), .ZN(n6534) );
  OR2_X1 U8920 ( .A1(n6733), .A2(n6728), .ZN(n6535) );
  NOR2_X1 U8921 ( .A1(n6733), .A2(n6729), .ZN(n6536) );
  AND2_X1 U8922 ( .A1(n12886), .A2(n7951), .ZN(n7224) );
  INV_X1 U8923 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n6901) );
  OR2_X1 U8924 ( .A1(n14528), .A2(n13992), .ZN(n13733) );
  NAND2_X1 U8925 ( .A1(n6439), .A2(n7199), .ZN(n6537) );
  INV_X1 U8926 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n7183) );
  XOR2_X1 U8927 ( .A(n12771), .B(n12284), .Z(n6538) );
  NAND2_X1 U8928 ( .A1(n14558), .A2(n6663), .ZN(n6661) );
  INV_X1 U8929 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6612) );
  INV_X1 U8930 ( .A(n14051), .ZN(n6830) );
  NAND2_X1 U8931 ( .A1(n11854), .A2(n7231), .ZN(n11959) );
  NAND2_X1 U8932 ( .A1(n7308), .A2(n7306), .ZN(n13964) );
  NAND2_X1 U8933 ( .A1(n6647), .A2(n6649), .ZN(n6539) );
  AND2_X1 U8934 ( .A1(n13942), .A2(n6824), .ZN(n6540) );
  INV_X1 U8935 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10438) );
  NAND2_X1 U8936 ( .A1(n7303), .A2(n11716), .ZN(n11847) );
  NOR2_X1 U8937 ( .A1(n15002), .A2(n9051), .ZN(n6541) );
  XOR2_X1 U8938 ( .A(n14432), .B(n14431), .Z(n6542) );
  OR2_X1 U8939 ( .A1(n12408), .A2(n7195), .ZN(n6543) );
  INV_X1 U8940 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7198) );
  NAND2_X1 U8941 ( .A1(n9545), .A2(n9544), .ZN(n14073) );
  INV_X1 U8942 ( .A(n14073), .ZN(n6822) );
  AND2_X1 U8943 ( .A1(n12248), .A2(n12247), .ZN(n6544) );
  NAND2_X1 U8944 ( .A1(n10283), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n6545) );
  NAND2_X1 U8945 ( .A1(n11820), .A2(n11822), .ZN(n11821) );
  OR2_X1 U8946 ( .A1(n10646), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n6546) );
  NAND2_X1 U8947 ( .A1(n12383), .A2(n12382), .ZN(n12380) );
  NOR3_X1 U8948 ( .A1(n13286), .A2(n13265), .A3(n6762), .ZN(n6761) );
  NAND2_X1 U8949 ( .A1(n7308), .A2(n13712), .ZN(n13965) );
  NAND2_X1 U8950 ( .A1(n6649), .A2(n7300), .ZN(n11849) );
  NOR2_X1 U8951 ( .A1(n14990), .A2(n9145), .ZN(n6547) );
  NOR2_X1 U8952 ( .A1(n15009), .A2(n9149), .ZN(n6548) );
  NOR2_X1 U8953 ( .A1(n12857), .A2(n12693), .ZN(n6549) );
  NAND2_X1 U8954 ( .A1(n13964), .A2(n13714), .ZN(n13939) );
  AND2_X1 U8955 ( .A1(n11966), .A2(n6687), .ZN(n6550) );
  NOR2_X1 U8956 ( .A1(n14558), .A2(n14557), .ZN(n6551) );
  INV_X1 U8957 ( .A(n8156), .ZN(n7118) );
  AND2_X1 U8958 ( .A1(n12271), .A2(n12270), .ZN(n6552) );
  NOR2_X1 U8959 ( .A1(n13416), .A2(n13014), .ZN(n6553) );
  NOR2_X1 U8960 ( .A1(n11979), .A2(n11980), .ZN(n7209) );
  AND2_X1 U8961 ( .A1(n7114), .A2(n7113), .ZN(n6554) );
  AND2_X1 U8962 ( .A1(n7052), .A2(n7051), .ZN(n6555) );
  AND2_X1 U8963 ( .A1(n12059), .A2(n12058), .ZN(n12062) );
  INV_X1 U8964 ( .A(n13940), .ZN(n13935) );
  INV_X1 U8965 ( .A(n14082), .ZN(n13915) );
  AND2_X1 U8966 ( .A1(n9531), .A2(n9530), .ZN(n14082) );
  AND2_X1 U8967 ( .A1(n10092), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n6556) );
  NAND2_X1 U8968 ( .A1(n10284), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n6557) );
  OR2_X1 U8969 ( .A1(n13286), .A2(n13265), .ZN(n6558) );
  OR2_X1 U8970 ( .A1(n12390), .A2(n12389), .ZN(n7207) );
  NAND2_X1 U8971 ( .A1(n12363), .A2(n12264), .ZN(n12406) );
  AND2_X1 U8972 ( .A1(n8160), .A2(n7116), .ZN(n6559) );
  INV_X1 U8973 ( .A(n6878), .ZN(n6876) );
  NAND2_X1 U8974 ( .A1(n12784), .A2(n12675), .ZN(n6878) );
  NOR2_X1 U8975 ( .A1(n11295), .A2(n6928), .ZN(n6925) );
  NAND2_X1 U8976 ( .A1(n7684), .A2(n7683), .ZN(n14480) );
  INV_X1 U8977 ( .A(n14480), .ZN(n6771) );
  NAND2_X1 U8978 ( .A1(n7179), .A2(n9856), .ZN(n10553) );
  NAND2_X1 U8979 ( .A1(n15166), .A2(n15084), .ZN(n12817) );
  NAND2_X1 U8980 ( .A1(n15146), .A2(n15084), .ZN(n12871) );
  NAND2_X1 U8981 ( .A1(n7834), .A2(n7833), .ZN(n13344) );
  INV_X1 U8982 ( .A(n13344), .ZN(n6767) );
  NAND2_X1 U8983 ( .A1(n9359), .A2(n9358), .ZN(n11594) );
  INV_X1 U8984 ( .A(n11594), .ZN(n6828) );
  INV_X1 U8985 ( .A(n11960), .ZN(n6686) );
  NAND2_X1 U8986 ( .A1(n9508), .A2(n9507), .ZN(n14221) );
  INV_X1 U8987 ( .A(n14221), .ZN(n6826) );
  AND2_X1 U8988 ( .A1(n11625), .A2(n11729), .ZN(n6560) );
  AND2_X1 U8989 ( .A1(n14898), .A2(n14490), .ZN(n13407) );
  NAND2_X1 U8990 ( .A1(n7770), .A2(n7769), .ZN(n13359) );
  INV_X1 U8991 ( .A(n13359), .ZN(n6763) );
  NAND2_X1 U8992 ( .A1(n11130), .A2(n11062), .ZN(n14629) );
  NAND2_X1 U8993 ( .A1(n6778), .A2(n8890), .ZN(n11246) );
  NAND2_X1 U8994 ( .A1(n6987), .A2(n11105), .ZN(n11213) );
  NAND2_X1 U8995 ( .A1(n11505), .A2(n11290), .ZN(n11361) );
  XNOR2_X1 U8996 ( .A(n11776), .B(n11763), .ZN(n11549) );
  AND2_X1 U8997 ( .A1(n14903), .A2(n14490), .ZN(n13351) );
  INV_X1 U8998 ( .A(n11105), .ZN(n6989) );
  NOR2_X1 U8999 ( .A1(n14954), .A2(n9141), .ZN(n6561) );
  NAND2_X1 U9000 ( .A1(n6439), .A2(n8376), .ZN(n8683) );
  OR2_X1 U9001 ( .A1(n8709), .A2(n7165), .ZN(n6562) );
  AND2_X1 U9002 ( .A1(n6751), .A2(n6754), .ZN(n6563) );
  NAND2_X1 U9003 ( .A1(n6437), .A2(n11511), .ZN(n6829) );
  AND2_X1 U9004 ( .A1(n7953), .A2(SI_26_), .ZN(n6564) );
  AND2_X1 U9005 ( .A1(n6563), .A2(n6747), .ZN(n6565) );
  AND2_X1 U9006 ( .A1(n7147), .A2(n7143), .ZN(n6566) );
  AND2_X1 U9007 ( .A1(n7144), .A2(n7143), .ZN(n6567) );
  NAND2_X1 U9008 ( .A1(n7305), .A2(n7304), .ZN(n11275) );
  AND2_X1 U9009 ( .A1(n12184), .A2(n7502), .ZN(n6568) );
  AND2_X1 U9010 ( .A1(n11803), .A2(n11802), .ZN(n6569) );
  AND2_X1 U9011 ( .A1(n11313), .A2(n9819), .ZN(n6570) );
  NAND4_X1 U9012 ( .A1(n8585), .A2(n8584), .A3(n8583), .A4(n8582), .ZN(n12447)
         );
  INV_X1 U9013 ( .A(n12447), .ZN(n6892) );
  AND2_X1 U9014 ( .A1(n11339), .A2(n10832), .ZN(n9887) );
  AND2_X1 U9015 ( .A1(n11084), .A2(n6454), .ZN(n6571) );
  INV_X1 U9016 ( .A(n14525), .ZN(n14729) );
  NAND2_X1 U9017 ( .A1(n7178), .A2(n10774), .ZN(n10805) );
  NAND2_X1 U9018 ( .A1(n10784), .A2(n10783), .ZN(n11009) );
  NAND2_X1 U9019 ( .A1(n7305), .A2(n11068), .ZN(n11276) );
  NAND2_X1 U9020 ( .A1(n6760), .A2(n10887), .ZN(n10861) );
  INV_X1 U9021 ( .A(n10861), .ZN(n6759) );
  AND2_X1 U9022 ( .A1(n10774), .A2(n10562), .ZN(n6572) );
  NAND2_X1 U9023 ( .A1(n12497), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n6573) );
  AND2_X1 U9024 ( .A1(n11009), .A2(n11008), .ZN(n6574) );
  INV_X1 U9025 ( .A(n13621), .ZN(n6613) );
  XOR2_X1 U9026 ( .A(n9885), .B(P3_REG1_REG_19__SCAN_IN), .Z(n6575) );
  NAND2_X1 U9027 ( .A1(n6907), .A2(n9180), .ZN(n14262) );
  OAI211_X1 U9028 ( .C1(n7003), .C2(P3_REG2_REG_2__SCAN_IN), .A(n7000), .B(
        n6998), .ZN(n10445) );
  INV_X1 U9029 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7139) );
  INV_X1 U9030 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6672) );
  INV_X1 U9031 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7057) );
  NAND2_X1 U9032 ( .A1(n8136), .A2(n8135), .ZN(n8139) );
  OAI21_X1 U9033 ( .B1(n8145), .B2(n8144), .A(n8143), .ZN(n8148) );
  NAND2_X1 U9034 ( .A1(n10755), .A2(n10757), .ZN(n10754) );
  NAND2_X1 U9035 ( .A1(n10612), .A2(n10611), .ZN(n10610) );
  NAND2_X1 U9036 ( .A1(n10972), .A2(n10974), .ZN(n10971) );
  NAND2_X1 U9037 ( .A1(n6579), .A2(n9935), .ZN(n11903) );
  INV_X1 U9038 ( .A(n7388), .ZN(n7354) );
  INV_X1 U9039 ( .A(n13185), .ZN(n6584) );
  NAND2_X1 U9040 ( .A1(n13252), .A2(n13251), .ZN(n13250) );
  OAI21_X2 U9041 ( .B1(n11621), .B2(n9930), .A(n9929), .ZN(n11634) );
  NAND2_X1 U9042 ( .A1(n14482), .A2(n9934), .ZN(n6579) );
  NAND2_X1 U9043 ( .A1(n12757), .A2(n6580), .ZN(P3_U3486) );
  NAND2_X1 U9044 ( .A1(n12828), .A2(n6581), .ZN(P3_U3454) );
  NAND2_X1 U9045 ( .A1(n13388), .A2(n6582), .ZN(P2_U3494) );
  NAND2_X1 U9046 ( .A1(n13316), .A2(n6583), .ZN(P2_U3526) );
  NAND2_X1 U9047 ( .A1(n8374), .A2(n8636), .ZN(n6867) );
  INV_X4 U9048 ( .A(n8504), .ZN(n8806) );
  NAND2_X1 U9049 ( .A1(n8693), .A2(n12687), .ZN(n12699) );
  NAND2_X1 U9050 ( .A1(n6428), .A2(n8381), .ZN(n8402) );
  NAND2_X1 U9051 ( .A1(n6777), .A2(n6775), .ZN(n11316) );
  NAND2_X1 U9052 ( .A1(n8603), .A2(n8917), .ZN(n11865) );
  NAND2_X1 U9053 ( .A1(n8676), .A2(n8858), .ZN(n12697) );
  OAI21_X1 U9054 ( .B1(n6757), .B2(n6756), .A(n6755), .ZN(n8261) );
  OAI21_X1 U9055 ( .B1(n11915), .B2(n8629), .A(n8926), .ZN(n12741) );
  NAND2_X1 U9056 ( .A1(n11634), .A2(n11633), .ZN(n7061) );
  NAND3_X1 U9057 ( .A1(n9443), .A2(n9442), .A3(n7260), .ZN(n6585) );
  NAND2_X2 U9058 ( .A1(n9184), .A2(n12031), .ZN(n9695) );
  XNOR2_X2 U9059 ( .A(n9181), .B(n9180), .ZN(n12031) );
  AOI21_X1 U9060 ( .B1(n9257), .B2(n9256), .A(n11066), .ZN(n9258) );
  NAND2_X1 U9061 ( .A1(n6587), .A2(n6586), .ZN(n9362) );
  NAND2_X1 U9062 ( .A1(n9584), .A2(n9583), .ZN(n9597) );
  NAND2_X1 U9063 ( .A1(n9620), .A2(n9619), .ZN(n9635) );
  NAND2_X1 U9064 ( .A1(n9262), .A2(n9261), .ZN(n9275) );
  NAND2_X1 U9065 ( .A1(n6585), .A2(n7262), .ZN(n7261) );
  NAND3_X1 U9066 ( .A1(n9177), .A2(n9178), .A3(n7317), .ZN(n9781) );
  NOR2_X2 U9067 ( .A1(n9251), .A2(n9168), .ZN(n9198) );
  NAND3_X1 U9068 ( .A1(n9331), .A2(n9330), .A3(n6527), .ZN(n6587) );
  NOR2_X2 U9069 ( .A1(n9193), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n9179) );
  NAND3_X1 U9070 ( .A1(n9177), .A2(n9198), .A3(n7318), .ZN(n9193) );
  OAI21_X2 U9071 ( .B1(n11463), .B2(n11462), .A(n11461), .ZN(n11475) );
  NAND2_X1 U9072 ( .A1(n12049), .A2(n12048), .ZN(n12052) );
  XNOR2_X1 U9073 ( .A(n13443), .B(n13444), .ZN(n13445) );
  NAND2_X1 U9074 ( .A1(n11999), .A2(n11998), .ZN(n6992) );
  NAND2_X1 U9075 ( .A1(n6978), .A2(n6977), .ZN(n13451) );
  OR2_X2 U9076 ( .A1(n13510), .A2(n6960), .ZN(n6589) );
  INV_X1 U9077 ( .A(n7376), .ZN(n7373) );
  NAND2_X1 U9078 ( .A1(n7371), .A2(n7419), .ZN(n7376) );
  NAND3_X1 U9079 ( .A1(n6691), .A2(n7529), .A3(n7233), .ZN(n6715) );
  NAND2_X1 U9080 ( .A1(n6716), .A2(n7503), .ZN(n6691) );
  NAND2_X1 U9081 ( .A1(n7807), .A2(n11210), .ZN(n7808) );
  NOR2_X1 U9082 ( .A1(n12534), .A2(n12533), .ZN(n12532) );
  NAND2_X1 U9083 ( .A1(n6590), .A2(n9160), .ZN(n9161) );
  XNOR2_X1 U9084 ( .A(n9157), .B(n6575), .ZN(n6590) );
  NOR2_X1 U9085 ( .A1(n14950), .A2(n15050), .ZN(n14949) );
  XNOR2_X1 U9086 ( .A(n9046), .B(n14959), .ZN(n14950) );
  INV_X1 U9087 ( .A(n9035), .ZN(n6596) );
  INV_X1 U9088 ( .A(n12454), .ZN(n6599) );
  NAND2_X1 U9089 ( .A1(n6992), .A2(n6991), .ZN(n12049) );
  NAND2_X1 U9090 ( .A1(n11924), .A2(n11923), .ZN(n11999) );
  OAI21_X2 U9091 ( .B1(n12130), .B2(n13501), .A(n13500), .ZN(n13499) );
  CLKBUF_X3 U9092 ( .A(n9198), .Z(n7317) );
  MUX2_X1 U9093 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n7479), .Z(n7439) );
  INV_X1 U9094 ( .A(n7640), .ZN(n6693) );
  OAI21_X2 U9095 ( .B1(n9714), .B2(n9713), .A(n9712), .ZN(n9766) );
  NAND2_X2 U9096 ( .A1(n8032), .A2(n12024), .ZN(n10114) );
  NAND2_X1 U9097 ( .A1(n11229), .A2(n9924), .ZN(n11325) );
  NAND2_X1 U9098 ( .A1(n7023), .A2(n7022), .ZN(n13185) );
  OAI22_X2 U9099 ( .A1(n13156), .A2(n13150), .B1(n13398), .B2(n12924), .ZN(
        n13136) );
  NOR2_X1 U9100 ( .A1(n6610), .A2(n6609), .ZN(n13386) );
  NOR2_X1 U9101 ( .A1(n7033), .A2(n9946), .ZN(n13107) );
  OAI21_X2 U9102 ( .B1(n13259), .B2(n6553), .A(n9992), .ZN(n13242) );
  NAND2_X1 U9103 ( .A1(n11492), .A2(n11489), .ZN(n6857) );
  NAND2_X1 U9104 ( .A1(n9962), .A2(n9961), .ZN(n6832) );
  NAND2_X1 U9105 ( .A1(n9958), .A2(n10483), .ZN(n10617) );
  OR2_X1 U9106 ( .A1(n8235), .A2(n10050), .ZN(n6833) );
  AOI21_X1 U9107 ( .B1(n13180), .B2(n13184), .A(n9999), .ZN(n13166) );
  AOI21_X2 U9108 ( .B1(n12081), .B2(n12080), .A(n13451), .ZN(n13510) );
  NAND2_X1 U9109 ( .A1(n11635), .A2(n9982), .ZN(n11745) );
  INV_X1 U9110 ( .A(n13313), .ZN(n6609) );
  NAND2_X4 U9111 ( .A1(n6433), .A2(n10049), .ZN(n8235) );
  XNOR2_X1 U9112 ( .A(n9048), .B(n9143), .ZN(n14987) );
  NOR2_X1 U9113 ( .A1(n14949), .A2(n9047), .ZN(n14971) );
  NOR2_X1 U9114 ( .A1(n10673), .A2(n9041), .ZN(n14929) );
  NAND2_X1 U9115 ( .A1(n9094), .A2(n9095), .ZN(n12455) );
  NOR2_X1 U9116 ( .A1(n15013), .A2(n15014), .ZN(n15012) );
  INV_X1 U9117 ( .A(n9103), .ZN(n6606) );
  AND3_X2 U9118 ( .A1(n7354), .A2(n7353), .A3(n7227), .ZN(n7358) );
  NAND2_X1 U9119 ( .A1(n13274), .A2(n9991), .ZN(n13259) );
  OAI21_X1 U9120 ( .B1(n6845), .B2(n6844), .A(n10003), .ZN(n13110) );
  INV_X4 U9121 ( .A(n10114), .ZN(n7790) );
  NAND2_X1 U9122 ( .A1(n13796), .A2(n6629), .ZN(n6623) );
  NAND2_X1 U9123 ( .A1(n13796), .A2(n7313), .ZN(n13787) );
  NAND3_X1 U9124 ( .A1(n6624), .A2(n6623), .A3(n6625), .ZN(n14026) );
  NAND3_X1 U9125 ( .A1(n6624), .A2(n6623), .A3(n6622), .ZN(n6633) );
  NAND2_X1 U9126 ( .A1(n6633), .A2(n6632), .ZN(n14246) );
  NAND2_X1 U9127 ( .A1(n13724), .A2(n6636), .ZN(n6634) );
  NAND2_X1 U9128 ( .A1(n6634), .A2(n6512), .ZN(n13810) );
  NAND2_X1 U9129 ( .A1(n6640), .A2(n6638), .ZN(n13908) );
  NAND2_X1 U9130 ( .A1(n6646), .A2(n11715), .ZN(n6645) );
  NAND2_X1 U9131 ( .A1(n6645), .A2(n6644), .ZN(n7292) );
  INV_X1 U9132 ( .A(n7300), .ZN(n6648) );
  INV_X1 U9133 ( .A(n7297), .ZN(n7296) );
  NAND2_X1 U9134 ( .A1(n11430), .A2(n11429), .ZN(n11432) );
  OAI211_X1 U9135 ( .C1(n7297), .C2(n11290), .A(n7295), .B(n6459), .ZN(n11430)
         );
  OAI21_X2 U9136 ( .B1(n10093), .B2(n9253), .A(n9323), .ZN(n11517) );
  XNOR2_X2 U9137 ( .A(n7530), .B(n7529), .ZN(n10093) );
  OAI21_X1 U9138 ( .B1(SI_6_), .B2(n6650), .A(n7525), .ZN(n7505) );
  MUX2_X1 U9139 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7438), .Z(n6650) );
  NAND2_X1 U9140 ( .A1(n14558), .A2(n6654), .ZN(n6653) );
  NAND3_X1 U9141 ( .A1(n7504), .A2(n7503), .A3(n7505), .ZN(n7507) );
  NAND2_X1 U9142 ( .A1(n12937), .A2(n6679), .ZN(n6677) );
  NAND2_X1 U9143 ( .A1(n6677), .A2(n6678), .ZN(n12927) );
  INV_X1 U9144 ( .A(n6681), .ZN(n12887) );
  OAI21_X2 U9145 ( .B1(n7757), .B2(n6688), .A(n6685), .ZN(n12905) );
  NAND3_X1 U9146 ( .A1(n10765), .A2(n12184), .A3(n7502), .ZN(n10764) );
  NAND2_X1 U9147 ( .A1(n6691), .A2(n7233), .ZN(n7526) );
  NAND2_X1 U9148 ( .A1(n6695), .A2(n6696), .ZN(n6694) );
  AND2_X1 U9149 ( .A1(n6944), .A2(n6942), .ZN(n13822) );
  NAND3_X1 U9150 ( .A1(n6713), .A2(n6712), .A3(n13733), .ZN(n13990) );
  INV_X1 U9151 ( .A(n7483), .ZN(n6716) );
  NAND2_X1 U9152 ( .A1(n6726), .A2(n6727), .ZN(n7240) );
  NAND2_X1 U9153 ( .A1(n7640), .A2(n6536), .ZN(n6726) );
  OAI21_X1 U9154 ( .B1(n6740), .B2(n7082), .A(n6738), .ZN(n6743) );
  NAND2_X1 U9155 ( .A1(n6743), .A2(n6742), .ZN(P2_U3328) );
  INV_X1 U9156 ( .A(n8186), .ZN(n6754) );
  AND2_X2 U9157 ( .A1(n13102), .A2(n10027), .ZN(n13082) );
  NOR2_X2 U9158 ( .A1(n10973), .A2(n11096), .ZN(n11159) );
  INV_X1 U9159 ( .A(n6761), .ZN(n13228) );
  INV_X1 U9160 ( .A(n13286), .ZN(n13268) );
  INV_X1 U9161 ( .A(n6774), .ZN(n11642) );
  NAND2_X1 U9162 ( .A1(n11194), .A2(n6779), .ZN(n6777) );
  NAND2_X1 U9163 ( .A1(n8550), .A2(n6784), .ZN(n6781) );
  NAND2_X1 U9164 ( .A1(n6781), .A2(n6782), .ZN(n8586) );
  NAND2_X1 U9165 ( .A1(n8719), .A2(n6795), .ZN(n6792) );
  NAND2_X1 U9166 ( .A1(n6792), .A2(n6793), .ZN(n12644) );
  OAI22_X1 U9167 ( .A1(n12625), .A2(n6799), .B1(n6800), .B2(n8849), .ZN(n12582) );
  INV_X1 U9168 ( .A(n8849), .ZN(n6803) );
  NAND2_X1 U9169 ( .A1(n6428), .A2(n6809), .ZN(n6812) );
  INV_X1 U9170 ( .A(n6812), .ZN(n8404) );
  XNOR2_X2 U9171 ( .A(n6811), .B(n8405), .ZN(n8408) );
  NAND2_X1 U9172 ( .A1(n12699), .A2(n6523), .ZN(n12677) );
  INV_X1 U9173 ( .A(n8841), .ZN(n6814) );
  NOR2_X1 U9174 ( .A1(n8841), .A2(n6815), .ZN(n8380) );
  INV_X1 U9175 ( .A(n8380), .ZN(n9023) );
  INV_X1 U9176 ( .A(n11271), .ZN(n6818) );
  NAND2_X1 U9177 ( .A1(n6817), .A2(n11084), .ZN(n11271) );
  NAND2_X1 U9178 ( .A1(n6818), .A2(n6819), .ZN(n14617) );
  XNOR2_X1 U9179 ( .A(n6820), .B(n9755), .ZN(n13696) );
  NOR2_X1 U9180 ( .A1(n13798), .A2(n14028), .ZN(n13779) );
  INV_X1 U9181 ( .A(n6829), .ZN(n11553) );
  NAND2_X1 U9182 ( .A1(n6832), .A2(n9963), .ZN(n9965) );
  XNOR2_X1 U9183 ( .A(n6832), .B(n10757), .ZN(n10759) );
  NAND2_X1 U9184 ( .A1(n10484), .A2(n9915), .ZN(n10483) );
  NAND4_X2 U9185 ( .A1(n7409), .A2(n7407), .A3(n7406), .A4(n7408), .ZN(n13030)
         );
  OAI21_X2 U9186 ( .B1(n10975), .B2(n6836), .A(n6834), .ZN(n11230) );
  OAI21_X1 U9187 ( .B1(n6836), .B2(n9969), .A(n6513), .ZN(n6835) );
  OR2_X1 U9188 ( .A1(n6837), .A2(n9972), .ZN(n6836) );
  NAND2_X1 U9189 ( .A1(n11230), .A2(n11226), .ZN(n9974) );
  NAND2_X1 U9190 ( .A1(n13149), .A2(n6534), .ZN(n6849) );
  AOI21_X2 U9191 ( .B1(n6849), .B2(n6846), .A(n6842), .ZN(n13108) );
  NAND2_X1 U9192 ( .A1(n6843), .A2(n6850), .ZN(n13121) );
  INV_X1 U9193 ( .A(n6843), .ZN(n6845) );
  NAND2_X1 U9194 ( .A1(n13109), .A2(n6848), .ZN(n6847) );
  OAI21_X1 U9195 ( .B1(n13149), .B2(n13155), .A(n6464), .ZN(n13137) );
  NAND2_X2 U9196 ( .A1(n6854), .A2(n7361), .ZN(n12024) );
  NAND2_X1 U9197 ( .A1(n6857), .A2(n6856), .ZN(n11616) );
  NAND2_X1 U9198 ( .A1(n8373), .A2(n8372), .ZN(n6866) );
  NAND3_X1 U9199 ( .A1(n6864), .A2(n6422), .A3(n6863), .ZN(n8841) );
  NAND2_X1 U9200 ( .A1(n12662), .A2(n6871), .ZN(n6869) );
  NAND2_X1 U9201 ( .A1(n9810), .A2(n6457), .ZN(n11026) );
  INV_X1 U9202 ( .A(n7329), .ZN(n6883) );
  OAI21_X2 U9203 ( .B1(n9818), .B2(n6887), .A(n6884), .ZN(n15027) );
  NAND2_X1 U9204 ( .A1(n14451), .A2(n6891), .ZN(n6890) );
  OR2_X1 U9205 ( .A1(n9840), .A2(n9841), .ZN(n6899) );
  AOI21_X1 U9206 ( .B1(n9841), .B2(n6518), .A(n6894), .ZN(n12567) );
  NAND2_X1 U9207 ( .A1(n8380), .A2(n8379), .ZN(n9022) );
  NAND2_X1 U9208 ( .A1(n8382), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8383) );
  NAND3_X2 U9209 ( .A1(n6906), .A2(n6905), .A3(n6908), .ZN(n14270) );
  CLKBUF_X1 U9210 ( .A(n9179), .Z(n6907) );
  INV_X2 U9211 ( .A(n14270), .ZN(n9184) );
  NAND3_X1 U9212 ( .A1(n6919), .A2(n6917), .A3(n14611), .ZN(n11299) );
  NAND3_X1 U9213 ( .A1(n11294), .A2(n11076), .A3(n6929), .ZN(n6919) );
  NAND2_X1 U9214 ( .A1(n11303), .A2(n6941), .ZN(n6932) );
  NAND2_X1 U9215 ( .A1(n11510), .A2(n6935), .ZN(n6934) );
  NAND2_X1 U9216 ( .A1(n11510), .A2(n6937), .ZN(n6936) );
  NOR2_X1 U9217 ( .A1(n11429), .A2(n6938), .ZN(n6937) );
  NAND2_X1 U9218 ( .A1(n13934), .A2(n6532), .ZN(n6950) );
  INV_X1 U9219 ( .A(n6950), .ZN(n13926) );
  AOI21_X1 U9220 ( .B1(n13990), .B2(n14007), .A(n13736), .ZN(n13979) );
  NAND2_X1 U9221 ( .A1(n11299), .A2(n11298), .ZN(n11510) );
  AND3_X2 U9222 ( .A1(n9239), .A2(n9238), .A3(n9237), .ZN(n14661) );
  OR2_X1 U9223 ( .A1(n6423), .A2(n10324), .ZN(n9217) );
  OR2_X2 U9224 ( .A1(n9179), .A2(n9445), .ZN(n9181) );
  NAND2_X4 U9225 ( .A1(n9184), .A2(n9182), .ZN(n9675) );
  OR2_X1 U9226 ( .A1(n9253), .A2(n10050), .ZN(n9220) );
  NAND2_X1 U9227 ( .A1(n7169), .A2(n7168), .ZN(n7167) );
  INV_X1 U9228 ( .A(n9808), .ZN(n10828) );
  NAND2_X1 U9229 ( .A1(n9014), .A2(n7167), .ZN(n7166) );
  NAND2_X1 U9230 ( .A1(n6951), .A2(n10903), .ZN(n10906) );
  NAND2_X1 U9231 ( .A1(n6951), .A2(n13537), .ZN(n10744) );
  AND2_X2 U9232 ( .A1(n6952), .A2(n10639), .ZN(n7344) );
  NAND2_X1 U9233 ( .A1(n6954), .A2(n10635), .ZN(n10639) );
  NAND2_X1 U9234 ( .A1(n6953), .A2(n10636), .ZN(n6952) );
  INV_X1 U9235 ( .A(n6954), .ZN(n6953) );
  XNOR2_X1 U9236 ( .A(n10632), .B(n12122), .ZN(n6954) );
  NAND2_X1 U9237 ( .A1(n13534), .A2(n12150), .ZN(n13443) );
  OAI211_X1 U9238 ( .C1(n13534), .C2(n6974), .A(n6972), .B(n6969), .ZN(n12170)
         );
  NAND2_X1 U9239 ( .A1(n13534), .A2(n6970), .ZN(n6969) );
  NOR2_X1 U9240 ( .A1(n12165), .A2(n6971), .ZN(n6970) );
  OAI21_X1 U9241 ( .B1(n12165), .B2(n6520), .A(n6973), .ZN(n6972) );
  NAND2_X1 U9242 ( .A1(n12165), .A2(n6975), .ZN(n6973) );
  NAND2_X1 U9243 ( .A1(n12165), .A2(n13444), .ZN(n6974) );
  NAND2_X1 U9244 ( .A1(n13481), .A2(n6524), .ZN(n6978) );
  NAND4_X1 U9245 ( .A1(n10907), .A2(n10945), .A3(n11212), .A4(n6990), .ZN(
        n6985) );
  NAND2_X1 U9246 ( .A1(n6985), .A2(n6986), .ZN(n11463) );
  AND2_X1 U9247 ( .A1(n6988), .A2(n11214), .ZN(n6986) );
  NAND3_X1 U9248 ( .A1(n10907), .A2(n10945), .A3(n6990), .ZN(n6987) );
  NAND2_X1 U9249 ( .A1(n10907), .A2(n10945), .ZN(n11107) );
  INV_X1 U9250 ( .A(n11106), .ZN(n6990) );
  NAND3_X1 U9251 ( .A1(n7317), .A2(n6993), .A3(n9201), .ZN(n9202) );
  NAND3_X1 U9252 ( .A1(n7003), .A2(n7004), .A3(n7001), .ZN(n7000) );
  OAI21_X1 U9253 ( .B1(n8445), .B2(n8479), .A(P3_IR_REG_2__SCAN_IN), .ZN(n7002) );
  NAND2_X1 U9254 ( .A1(n8445), .A2(P3_IR_REG_2__SCAN_IN), .ZN(n7004) );
  INV_X1 U9255 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n7005) );
  OR2_X2 U9256 ( .A1(n14434), .A2(n7011), .ZN(n7008) );
  INV_X1 U9257 ( .A(n7013), .ZN(n14433) );
  INV_X1 U9258 ( .A(n9054), .ZN(n7012) );
  INV_X1 U9259 ( .A(n9036), .ZN(n7014) );
  OAI21_X1 U9260 ( .B1(n15003), .B2(n7019), .A(n7018), .ZN(n9052) );
  NOR2_X2 U9261 ( .A1(n14969), .A2(n7021), .ZN(n9048) );
  NOR2_X1 U9262 ( .A1(n13130), .A2(n7038), .ZN(n7033) );
  XNOR2_X1 U9263 ( .A(n13091), .B(n13090), .ZN(n13303) );
  INV_X1 U9264 ( .A(n14376), .ZN(n14380) );
  OAI21_X1 U9265 ( .B1(n14564), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7043), .ZN(
        n7042) );
  AND2_X1 U9266 ( .A1(n14376), .A2(n7044), .ZN(n14564) );
  INV_X1 U9267 ( .A(n14381), .ZN(n7044) );
  AOI21_X1 U9268 ( .B1(n11903), .B2(n6521), .A(n7046), .ZN(n13252) );
  NAND2_X1 U9269 ( .A1(n11156), .A2(n7060), .ZN(n11229) );
  OAI21_X2 U9270 ( .B1(n15010), .B2(n7063), .A(n7062), .ZN(n12469) );
  INV_X1 U9271 ( .A(n7064), .ZN(n14914) );
  NAND2_X1 U9272 ( .A1(n6441), .A2(n9131), .ZN(n14915) );
  NOR2_X1 U9273 ( .A1(n14955), .A2(n15161), .ZN(n14954) );
  INV_X1 U9274 ( .A(n14975), .ZN(n7067) );
  MUX2_X1 U9275 ( .A(n10967), .B(n6429), .S(n8096), .Z(n8055) );
  NOR2_X1 U9276 ( .A1(n8288), .A2(n8293), .ZN(n7081) );
  NAND2_X1 U9277 ( .A1(n8266), .A2(n8265), .ZN(n7082) );
  NAND2_X1 U9278 ( .A1(n7083), .A2(n7084), .ZN(n8107) );
  NAND3_X1 U9279 ( .A1(n8101), .A2(n6533), .A3(n8100), .ZN(n7083) );
  NAND2_X1 U9280 ( .A1(n7085), .A2(n7086), .ZN(n8087) );
  NAND3_X1 U9281 ( .A1(n8081), .A2(n6498), .A3(n8080), .ZN(n7085) );
  NAND2_X1 U9282 ( .A1(n8114), .A2(n7090), .ZN(n7087) );
  NAND2_X1 U9283 ( .A1(n7087), .A2(n7088), .ZN(n8117) );
  NAND2_X1 U9284 ( .A1(n8071), .A2(n7095), .ZN(n7093) );
  NAND2_X1 U9285 ( .A1(n7093), .A2(n7092), .ZN(n8076) );
  AOI21_X1 U9286 ( .B1(n7097), .B2(n7095), .A(n7094), .ZN(n7092) );
  OAI21_X1 U9287 ( .B1(n8071), .B2(n7097), .A(n7095), .ZN(n8077) );
  NAND2_X1 U9288 ( .A1(n8122), .A2(n7101), .ZN(n7098) );
  NAND2_X1 U9289 ( .A1(n7098), .A2(n7099), .ZN(n8125) );
  NAND2_X1 U9290 ( .A1(n8094), .A2(n7107), .ZN(n7104) );
  NAND2_X1 U9291 ( .A1(n7104), .A2(n7105), .ZN(n8098) );
  AOI21_X1 U9292 ( .B1(n7109), .B2(n7107), .A(n7106), .ZN(n7105) );
  NAND2_X1 U9293 ( .A1(n8164), .A2(n7113), .ZN(n7110) );
  OAI21_X1 U9294 ( .B1(n8164), .B2(n7114), .A(n7113), .ZN(n8170) );
  NAND2_X1 U9295 ( .A1(n7110), .A2(n7111), .ZN(n8169) );
  NAND2_X1 U9296 ( .A1(n8155), .A2(n7117), .ZN(n7115) );
  OAI21_X1 U9297 ( .B1(n8155), .B2(n7119), .A(n7117), .ZN(n8159) );
  NAND2_X1 U9298 ( .A1(n7115), .A2(n6559), .ZN(n8158) );
  NAND2_X1 U9299 ( .A1(n8493), .A2(n6517), .ZN(n7133) );
  NAND2_X1 U9300 ( .A1(n8725), .A2(n6567), .ZN(n7140) );
  NAND2_X1 U9301 ( .A1(n7140), .A2(n7141), .ZN(n8345) );
  NAND2_X1 U9302 ( .A1(n8647), .A2(n7157), .ZN(n8333) );
  NAND2_X1 U9303 ( .A1(n7161), .A2(n7160), .ZN(n8590) );
  NAND2_X1 U9304 ( .A1(n8696), .A2(n7164), .ZN(n7163) );
  NAND2_X1 U9305 ( .A1(n7170), .A2(n8984), .ZN(n8986) );
  NAND3_X1 U9306 ( .A1(n7174), .A2(n7171), .A3(n9007), .ZN(n7170) );
  OAI21_X1 U9307 ( .B1(n7176), .B2(n7173), .A(n7172), .ZN(n7171) );
  NOR2_X1 U9308 ( .A1(n8981), .A2(n9883), .ZN(n7172) );
  INV_X1 U9309 ( .A(n8982), .ZN(n7173) );
  NAND2_X1 U9310 ( .A1(n7175), .A2(n9883), .ZN(n7174) );
  NAND2_X1 U9311 ( .A1(n7176), .A2(n8979), .ZN(n7175) );
  NAND2_X1 U9312 ( .A1(n10805), .A2(n10806), .ZN(n10779) );
  NAND2_X1 U9313 ( .A1(n7179), .A2(n6522), .ZN(n10557) );
  NAND2_X1 U9314 ( .A1(n7187), .A2(n7188), .ZN(n12312) );
  INV_X1 U9315 ( .A(n11738), .ZN(n7214) );
  NAND2_X1 U9316 ( .A1(n11651), .A2(n7217), .ZN(n7216) );
  NAND2_X1 U9317 ( .A1(n7221), .A2(n7222), .ZN(n7990) );
  NAND2_X1 U9318 ( .A1(n12927), .A2(n7224), .ZN(n7221) );
  NAND2_X1 U9319 ( .A1(n7225), .A2(n11044), .ZN(n11046) );
  AND2_X1 U9320 ( .A1(n7336), .A2(n7226), .ZN(n7227) );
  NAND2_X1 U9321 ( .A1(n7336), .A2(n7386), .ZN(n7229) );
  NAND2_X1 U9322 ( .A1(n11155), .A2(n7230), .ZN(n11451) );
  NAND2_X1 U9323 ( .A1(n11853), .A2(n7717), .ZN(n11854) );
  NAND3_X1 U9324 ( .A1(n10857), .A2(n7435), .A3(n7324), .ZN(n7498) );
  NAND2_X1 U9325 ( .A1(n7431), .A2(n10850), .ZN(n10857) );
  INV_X1 U9326 ( .A(n7503), .ZN(n7235) );
  INV_X1 U9327 ( .A(n7234), .ZN(n7233) );
  OAI21_X1 U9328 ( .B1(n7482), .B2(n7235), .A(n7506), .ZN(n7234) );
  NAND2_X1 U9329 ( .A1(n7553), .A2(n7251), .ZN(n7250) );
  NAND2_X1 U9330 ( .A1(n7826), .A2(n7256), .ZN(n7831) );
  NAND2_X1 U9331 ( .A1(n7826), .A2(n7808), .ZN(n7811) );
  NAND2_X1 U9332 ( .A1(n7851), .A2(n7869), .ZN(n7853) );
  NAND2_X1 U9333 ( .A1(n7872), .A2(n7869), .ZN(n7867) );
  NAND2_X1 U9334 ( .A1(n7479), .A2(n8426), .ZN(n7259) );
  NAND4_X1 U9335 ( .A1(n7365), .A2(n7364), .A3(P2_ADDR_REG_19__SCAN_IN), .A4(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n7257) );
  NAND4_X1 U9336 ( .A1(n12243), .A2(n7363), .A3(n7362), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7258) );
  OAI21_X1 U9337 ( .B1(n7479), .B2(P2_DATAO_REG_0__SCAN_IN), .A(n7259), .ZN(
        n7372) );
  NAND3_X1 U9338 ( .A1(n9640), .A2(n9639), .A3(n7267), .ZN(n7270) );
  NAND2_X1 U9339 ( .A1(n9653), .A2(n7268), .ZN(n7267) );
  NAND2_X1 U9340 ( .A1(n7270), .A2(n7269), .ZN(n9665) );
  NAND2_X1 U9341 ( .A1(n9668), .A2(n9667), .ZN(n7273) );
  NAND2_X1 U9342 ( .A1(n9664), .A2(n9663), .ZN(n7274) );
  NAND3_X1 U9343 ( .A1(n7274), .A2(n7273), .A3(n6490), .ZN(n7272) );
  NAND2_X1 U9344 ( .A1(n9204), .A2(n7276), .ZN(n9767) );
  XNOR2_X2 U9345 ( .A(n7277), .B(P1_IR_REG_22__SCAN_IN), .ZN(n9719) );
  NAND2_X1 U9346 ( .A1(n9362), .A2(n9363), .ZN(n9361) );
  NAND3_X1 U9347 ( .A1(n9397), .A2(n9396), .A3(n6526), .ZN(n7278) );
  NAND2_X1 U9348 ( .A1(n7278), .A2(n7279), .ZN(n9426) );
  NAND3_X1 U9349 ( .A1(n9367), .A2(n9366), .A3(n6528), .ZN(n7281) );
  NAND2_X1 U9350 ( .A1(n7281), .A2(n7282), .ZN(n9392) );
  NAND3_X1 U9351 ( .A1(n9297), .A2(n9296), .A3(n6530), .ZN(n7284) );
  NAND2_X1 U9352 ( .A1(n7284), .A2(n7285), .ZN(n9326) );
  NAND2_X1 U9353 ( .A1(n7288), .A2(n7290), .ZN(n9561) );
  NAND3_X1 U9354 ( .A1(n9536), .A2(n9535), .A3(n7289), .ZN(n7288) );
  NAND2_X1 U9355 ( .A1(n11128), .A2(n11061), .ZN(n11130) );
  INV_X1 U9356 ( .A(n7292), .ZN(n14006) );
  NAND2_X1 U9357 ( .A1(n7292), .A2(n13989), .ZN(n14004) );
  INV_X1 U9358 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7293) );
  NAND3_X1 U9359 ( .A1(n9235), .A2(n7294), .A3(n7293), .ZN(n9248) );
  INV_X2 U9360 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9235) );
  NAND2_X1 U9361 ( .A1(n11507), .A2(n7296), .ZN(n7295) );
  NAND2_X1 U9362 ( .A1(n13972), .A2(n13737), .ZN(n7308) );
  NAND2_X1 U9363 ( .A1(n13796), .A2(n13730), .ZN(n13785) );
  NAND2_X1 U9364 ( .A1(n13908), .A2(n7316), .ZN(n13896) );
  AOI21_X1 U9365 ( .B1(n13872), .B2(n13873), .A(n13720), .ZN(n13864) );
  XNOR2_X2 U9366 ( .A(n10887), .B(n13027), .ZN(n10757) );
  NAND4_X2 U9367 ( .A1(n7458), .A2(n7457), .A3(n7456), .A4(n7455), .ZN(n13027)
         );
  NAND2_X1 U9368 ( .A1(n7966), .A2(n10129), .ZN(n7470) );
  BUF_X4 U9369 ( .A(n7453), .Z(n7966) );
  INV_X1 U9370 ( .A(n15062), .ZN(n12452) );
  NAND2_X1 U9371 ( .A1(n9128), .A2(n9127), .ZN(n10451) );
  NAND2_X1 U9372 ( .A1(n15062), .A2(n9802), .ZN(n10558) );
  NAND2_X1 U9373 ( .A1(n12452), .A2(n9802), .ZN(n8865) );
  NAND2_X1 U9374 ( .A1(n8865), .A2(n10559), .ZN(n9801) );
  NAND2_X1 U9375 ( .A1(n12284), .A2(n10559), .ZN(n10560) );
  NAND2_X1 U9376 ( .A1(n8677), .A2(n8678), .ZN(n8682) );
  NAND2_X1 U9377 ( .A1(n7453), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n7402) );
  INV_X1 U9378 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n7531) );
  INV_X1 U9379 ( .A(n8493), .ZN(n8495) );
  INV_X1 U9380 ( .A(n7368), .ZN(n7370) );
  INV_X1 U9381 ( .A(n14473), .ZN(n9987) );
  NAND2_X1 U9382 ( .A1(n8210), .A2(n8190), .ZN(n7975) );
  INV_X1 U9383 ( .A(n12983), .ZN(n12997) );
  NAND2_X1 U9384 ( .A1(n12905), .A2(n7800), .ZN(n12902) );
  NOR2_X1 U9385 ( .A1(n13306), .A2(n13305), .ZN(n13308) );
  NAND2_X1 U9386 ( .A1(n9916), .A2(n10696), .ZN(n10479) );
  NAND2_X1 U9387 ( .A1(n12303), .A2(n7327), .ZN(n12281) );
  NAND4_X2 U9388 ( .A1(n8444), .A2(n8443), .A3(n8442), .A4(n8441), .ZN(n15078)
         );
  CLKBUF_X1 U9389 ( .A(n10764), .Z(n11043) );
  INV_X1 U9390 ( .A(n11815), .ZN(n10009) );
  AND2_X1 U9391 ( .A1(n11815), .A2(n11598), .ZN(n10293) );
  INV_X1 U9392 ( .A(n7512), .ZN(n7821) );
  NOR2_X2 U9393 ( .A1(n8408), .A2(n8407), .ZN(n8440) );
  NAND4_X2 U9394 ( .A1(n7471), .A2(n7470), .A3(n7469), .A4(n7468), .ZN(n13028)
         );
  OR2_X1 U9395 ( .A1(n13303), .A2(n13362), .ZN(n13311) );
  OR2_X1 U9396 ( .A1(n9675), .A2(n11139), .ZN(n9216) );
  INV_X1 U9397 ( .A(n12330), .ZN(n12558) );
  INV_X1 U9398 ( .A(n10449), .ZN(n9127) );
  NAND2_X1 U9399 ( .A1(n9012), .A2(n9791), .ZN(n9014) );
  OAI22_X1 U9400 ( .A1(n9012), .A2(n15086), .B1(n9011), .B2(n10554), .ZN(n9013) );
  NAND2_X1 U9401 ( .A1(n8801), .A2(n8357), .ZN(n8814) );
  OR2_X1 U9402 ( .A1(n12038), .A2(n8235), .ZN(n7876) );
  CLKBUF_X1 U9403 ( .A(n11475), .Z(n11480) );
  NAND2_X1 U9404 ( .A1(n7479), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7366) );
  NAND2_X1 U9405 ( .A1(n8218), .A2(n8217), .ZN(n8282) );
  INV_X1 U9406 ( .A(n9248), .ZN(n9164) );
  OR3_X1 U9408 ( .A1(n11908), .A2(n9849), .A3(n11955), .ZN(n10537) );
  XNOR2_X1 U9409 ( .A(n11071), .B(n9310), .ZN(n9222) );
  XNOR2_X1 U9410 ( .A(n8188), .B(n7956), .ZN(n12023) );
  OAI21_X1 U9411 ( .B1(n9711), .B2(n9710), .A(n9709), .ZN(n9712) );
  OR2_X1 U9412 ( .A1(n14272), .A2(n9253), .ZN(n9686) );
  OR2_X1 U9413 ( .A1(n6425), .A2(n10328), .ZN(n9245) );
  OR2_X1 U9414 ( .A1(n6423), .A2(n10602), .ZN(n9189) );
  AND2_X1 U9415 ( .A1(n13359), .A2(n9993), .ZN(n7319) );
  OR2_X1 U9416 ( .A1(n13359), .A2(n9993), .ZN(n7320) );
  NAND2_X1 U9417 ( .A1(n12803), .A2(n12710), .ZN(n7321) );
  INV_X1 U9418 ( .A(n11835), .ZN(n11850) );
  OR2_X1 U9419 ( .A1(n12548), .A2(n12817), .ZN(n7322) );
  OR2_X1 U9420 ( .A1(n12548), .A2(n12871), .ZN(n7323) );
  AND2_X2 U9421 ( .A1(n9872), .A2(n10573), .ZN(n15146) );
  AND2_X1 U9422 ( .A1(n7476), .A2(n10402), .ZN(n7324) );
  OR2_X1 U9423 ( .A1(n10637), .A2(n12122), .ZN(n7325) );
  AND2_X1 U9424 ( .A1(n12274), .A2(n7328), .ZN(n7327) );
  OR2_X1 U9425 ( .A1(n12302), .A2(n12654), .ZN(n7328) );
  NOR2_X1 U9426 ( .A1(n9831), .A2(n12705), .ZN(n7329) );
  AND2_X1 U9427 ( .A1(n10001), .A2(n12979), .ZN(n7330) );
  AND2_X1 U9428 ( .A1(n14023), .A2(n14022), .ZN(n7331) );
  OR2_X1 U9429 ( .A1(n9132), .A2(n9037), .ZN(n7332) );
  AND2_X1 U9430 ( .A1(n13008), .A2(n7799), .ZN(n7333) );
  OR2_X1 U9431 ( .A1(n10594), .A2(n11125), .ZN(n7334) );
  AND4_X1 U9432 ( .A1(n8378), .A2(n8377), .A3(n8846), .A4(n7183), .ZN(n7335)
         );
  INV_X1 U9433 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7367) );
  AND4_X1 U9434 ( .A1(n7356), .A2(n7355), .A3(n7993), .A4(n7991), .ZN(n7336)
         );
  AND2_X2 U9435 ( .A1(n11057), .A2(n13913), .ZN(n14647) );
  INV_X1 U9436 ( .A(n14647), .ZN(n13962) );
  OR2_X1 U9437 ( .A1(n13302), .A2(n13254), .ZN(n7337) );
  NAND2_X2 U9438 ( .A1(n9953), .A2(n14863), .ZN(n14868) );
  INV_X1 U9439 ( .A(n12668), .ZN(n8718) );
  INV_X1 U9440 ( .A(n10161), .ZN(n9772) );
  INV_X1 U9441 ( .A(n9132), .ZN(n10478) );
  AND2_X1 U9442 ( .A1(n10293), .A2(n8296), .ZN(n14490) );
  AND2_X1 U9443 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7338) );
  XNOR2_X1 U9444 ( .A(n10967), .B(n7987), .ZN(n7410) );
  AND2_X1 U9445 ( .A1(n9764), .A2(n9763), .ZN(n7341) );
  OR2_X1 U9446 ( .A1(n13378), .A2(n13079), .ZN(n7342) );
  AND2_X1 U9447 ( .A1(n12602), .A2(n12583), .ZN(n7343) );
  INV_X1 U9448 ( .A(n15041), .ZN(n9820) );
  AND2_X1 U9449 ( .A1(n9242), .A2(n14638), .ZN(n9256) );
  NAND2_X1 U9450 ( .A1(n8069), .A2(n8068), .ZN(n8071) );
  MUX2_X1 U9451 ( .A(n13567), .B(n11517), .S(n9707), .Z(n9327) );
  NAND2_X1 U9452 ( .A1(n8092), .A2(n8091), .ZN(n8094) );
  MUX2_X1 U9453 ( .A(n13565), .B(n11594), .S(n9289), .Z(n9363) );
  MUX2_X1 U9454 ( .A(n13563), .B(n11797), .S(n9289), .Z(n9393) );
  NAND2_X1 U9455 ( .A1(n8112), .A2(n8111), .ZN(n8114) );
  AND2_X1 U9456 ( .A1(n9499), .A2(n9497), .ZN(n9498) );
  NAND2_X1 U9457 ( .A1(n8128), .A2(n8127), .ZN(n8131) );
  MUX2_X1 U9458 ( .A(n13721), .B(n14058), .S(n9725), .Z(n9580) );
  MUX2_X1 U9459 ( .A(n13725), .B(n14051), .S(n9289), .Z(n9598) );
  MUX2_X1 U9460 ( .A(n13749), .B(n13817), .S(n9707), .Z(n9636) );
  NAND2_X1 U9461 ( .A1(n8162), .A2(n8161), .ZN(n8164) );
  INV_X1 U9462 ( .A(n8221), .ZN(n8182) );
  INV_X1 U9463 ( .A(n8167), .ZN(n8168) );
  NAND2_X1 U9464 ( .A1(n8183), .A2(n8182), .ZN(n8184) );
  INV_X1 U9465 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n7346) );
  INV_X1 U9466 ( .A(n9032), .ZN(n9030) );
  INV_X1 U9467 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n9037) );
  INV_X1 U9468 ( .A(n11030), .ZN(n9811) );
  INV_X1 U9469 ( .A(n13277), .ZN(n9989) );
  AOI22_X1 U9470 ( .A1(n10625), .A2(n11125), .B1(n10597), .B2(n14284), .ZN(
        n10598) );
  OAI22_X1 U9471 ( .A1(n10900), .A2(n10631), .B1(n9224), .B2(n6434), .ZN(
        n10632) );
  OR4_X1 U9472 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n10302) );
  INV_X1 U9473 ( .A(n10066), .ZN(n8437) );
  INV_X1 U9474 ( .A(n10782), .ZN(n10783) );
  INV_X1 U9475 ( .A(n8657), .ZN(n8391) );
  INV_X1 U9476 ( .A(n10799), .ZN(n9136) );
  INV_X1 U9477 ( .A(n14437), .ZN(n9150) );
  AND2_X1 U9478 ( .A1(n9797), .A2(n9843), .ZN(n9844) );
  INV_X1 U9479 ( .A(n9839), .ZN(n12626) );
  INV_X1 U9480 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8846) );
  NOR2_X1 U9481 ( .A1(n7939), .A2(n12989), .ZN(n7959) );
  NOR2_X1 U9482 ( .A1(n7879), .A2(n7877), .ZN(n7903) );
  INV_X1 U9483 ( .A(n9955), .ZN(n8290) );
  AND2_X1 U9484 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n7623) );
  INV_X1 U9485 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7357) );
  NAND2_X1 U9486 ( .A1(n10625), .A2(n13572), .ZN(n10626) );
  INV_X1 U9487 ( .A(n13835), .ZN(n13727) );
  INV_X1 U9488 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9434) );
  INV_X1 U9489 ( .A(n13851), .ZN(n13723) );
  INV_X1 U9490 ( .A(n7952), .ZN(n7953) );
  INV_X1 U9491 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9201) );
  NAND2_X1 U9492 ( .A1(n9164), .A2(n9163), .ZN(n9251) );
  INV_X1 U9493 ( .A(n11526), .ZN(n11382) );
  INV_X1 U9494 ( .A(n8623), .ZN(n8390) );
  INV_X1 U9495 ( .A(n12337), .ZN(n12271) );
  INV_X1 U9496 ( .A(n8713), .ZN(n8395) );
  NAND2_X1 U9497 ( .A1(n8399), .A2(n8398), .ZN(n8790) );
  INV_X1 U9498 ( .A(n8408), .ZN(n8406) );
  NAND2_X1 U9499 ( .A1(n8874), .A2(n8875), .ZN(n9805) );
  INV_X1 U9500 ( .A(n9822), .ZN(n15026) );
  OR2_X1 U9501 ( .A1(n9855), .A2(n9866), .ZN(n9878) );
  INV_X1 U9502 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n8320) );
  AND2_X1 U9503 ( .A1(n7959), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n7978) );
  OR2_X1 U9504 ( .A1(n7561), .A2(n7560), .ZN(n7580) );
  INV_X1 U9505 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7489) );
  OR2_X1 U9506 ( .A1(n7816), .A2(n7815), .ZN(n7835) );
  INV_X1 U9507 ( .A(n8282), .ZN(n10027) );
  INV_X1 U9508 ( .A(n13306), .ZN(n8267) );
  NAND2_X1 U9509 ( .A1(n13001), .A2(n13078), .ZN(n10014) );
  AND2_X1 U9510 ( .A1(n7680), .A2(n7679), .ZN(n7705) );
  INV_X1 U9511 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n9575) );
  INV_X1 U9512 ( .A(n11791), .ZN(n11788) );
  OR2_X1 U9513 ( .A1(n9450), .A2(n14183), .ZN(n9484) );
  INV_X1 U9514 ( .A(n9604), .ZN(n9605) );
  AND2_X1 U9515 ( .A1(n9524), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n9537) );
  INV_X1 U9516 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10335) );
  NOR2_X1 U9517 ( .A1(n13783), .A2(n13765), .ZN(n13753) );
  NAND2_X1 U9518 ( .A1(n13874), .A2(n14066), .ZN(n13876) );
  INV_X1 U9519 ( .A(n14528), .ZN(n11841) );
  AND2_X1 U9520 ( .A1(n9399), .A2(n9398), .ZN(n9413) );
  AND2_X1 U9521 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9279) );
  OR2_X1 U9522 ( .A1(n11141), .A2(n11125), .ZN(n14637) );
  INV_X1 U9523 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9770) );
  INV_X1 U9524 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9178) );
  INV_X1 U9525 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n14307) );
  NAND2_X1 U9526 ( .A1(n8390), .A2(n12294), .ZN(n8640) );
  AND2_X1 U9527 ( .A1(n12279), .A2(n12278), .ZN(n12280) );
  INV_X1 U9528 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n11740) );
  OR2_X1 U9529 ( .A1(n10570), .A2(n10546), .ZN(n12421) );
  AND2_X1 U9530 ( .A1(n10573), .A2(n9026), .ZN(n10549) );
  INV_X1 U9531 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14988) );
  OR2_X1 U9532 ( .A1(n8753), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8764) );
  OR2_X1 U9533 ( .A1(n9836), .A2(n6514), .ZN(n12655) );
  AND2_X1 U9534 ( .A1(n8932), .A2(n8929), .ZN(n12740) );
  OR2_X1 U9535 ( .A1(n10547), .A2(n9883), .ZN(n15061) );
  NOR2_X1 U9536 ( .A1(n8520), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8534) );
  OR2_X1 U9537 ( .A1(n10813), .A2(n10553), .ZN(n9881) );
  INV_X1 U9538 ( .A(n11269), .ZN(n12540) );
  AND2_X1 U9539 ( .A1(n9868), .A2(n9845), .ZN(n12736) );
  INV_X1 U9540 ( .A(n15083), .ZN(n15067) );
  NAND2_X1 U9541 ( .A1(n9884), .A2(n11360), .ZN(n15130) );
  AND2_X1 U9542 ( .A1(n10090), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8314) );
  NAND2_X1 U9543 ( .A1(n8003), .A2(n7993), .ZN(n8006) );
  OR2_X1 U9544 ( .A1(n7919), .A2(n12931), .ZN(n7939) );
  NAND2_X1 U9545 ( .A1(n7887), .A2(n7889), .ZN(n7890) );
  OR2_X1 U9546 ( .A1(n7644), .A2(n11657), .ZN(n7688) );
  INV_X1 U9547 ( .A(n11453), .ZN(n7611) );
  OR2_X1 U9548 ( .A1(n7835), .A2(n12919), .ZN(n7879) );
  INV_X1 U9549 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n11657) );
  INV_X1 U9550 ( .A(n14820), .ZN(n14838) );
  INV_X1 U9551 ( .A(n13227), .ZN(n13246) );
  INV_X1 U9552 ( .A(n9938), .ZN(n13251) );
  INV_X1 U9553 ( .A(n10611), .ZN(n10616) );
  AND2_X1 U9554 ( .A1(n10113), .A2(n8296), .ZN(n10490) );
  AOI22_X1 U9555 ( .A1(n13091), .A2(n13090), .B1(n8267), .B2(n13003), .ZN(
        n9949) );
  INV_X1 U9556 ( .A(n11860), .ZN(n14493) );
  INV_X1 U9557 ( .A(n11636), .ZN(n11633) );
  INV_X1 U9558 ( .A(n14475), .ZN(n13279) );
  OR2_X1 U9559 ( .A1(n11056), .A2(n9772), .ZN(n10275) );
  OAI22_X1 U9560 ( .A1(n12159), .A2(n11067), .B1(n11190), .B2(n12162), .ZN(
        n10896) );
  AND2_X1 U9561 ( .A1(n9537), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9549) );
  INV_X1 U9562 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14293) );
  INV_X1 U9563 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n14183) );
  INV_X1 U9564 ( .A(n9784), .ZN(n13587) );
  INV_X1 U9565 ( .A(n13713), .ZN(n13966) );
  OR2_X1 U9566 ( .A1(n10103), .A2(n10311), .ZN(n10312) );
  AND2_X1 U9567 ( .A1(n8229), .A2(n8196), .ZN(n8197) );
  XNOR2_X1 U9568 ( .A(n7764), .B(SI_17_), .ZN(n7762) );
  AOI22_X1 U9569 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14301), .B1(n14348), .B2(
        n14300), .ZN(n14303) );
  NAND2_X1 U9570 ( .A1(n11978), .A2(n11977), .ZN(n11979) );
  XNOR2_X1 U9571 ( .A(n11378), .B(n12449), .ZN(n11375) );
  INV_X1 U9572 ( .A(n12433), .ZN(n12418) );
  NAND2_X1 U9573 ( .A1(n10771), .A2(n11576), .ZN(n12437) );
  OR2_X1 U9574 ( .A1(n12541), .A2(n8504), .ZN(n8838) );
  AND4_X1 U9575 ( .A1(n8645), .A2(n8644), .A3(n8643), .A4(n8642), .ZN(n12357)
         );
  NOR2_X1 U9576 ( .A1(n9044), .A2(n10788), .ZN(n10988) );
  INV_X1 U9577 ( .A(n15017), .ZN(n9160) );
  NAND2_X1 U9578 ( .A1(n9794), .A2(n9882), .ZN(n15083) );
  AND2_X1 U9579 ( .A1(n12699), .A2(n12698), .ZN(n12795) );
  INV_X1 U9580 ( .A(n12553), .ZN(n14458) );
  AND2_X1 U9581 ( .A1(n10547), .A2(n9887), .ZN(n15079) );
  NOR2_X1 U9582 ( .A1(n10819), .A2(n15054), .ZN(n15048) );
  INV_X1 U9583 ( .A(n15090), .ZN(n15056) );
  AND3_X1 U9584 ( .A1(n9881), .A2(n9880), .A3(n9879), .ZN(n10817) );
  AND2_X1 U9585 ( .A1(n9884), .A2(n15054), .ZN(n15143) );
  INV_X1 U9586 ( .A(n15130), .ZN(n15084) );
  NOR2_X1 U9587 ( .A1(n10209), .A2(n10208), .ZN(n10213) );
  INV_X1 U9588 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8591) );
  AND2_X1 U9589 ( .A1(n8018), .A2(n12015), .ZN(n8002) );
  AND2_X1 U9590 ( .A1(n12187), .A2(n7694), .ZN(n7695) );
  AND2_X1 U9591 ( .A1(n7496), .A2(n12177), .ZN(n7497) );
  NAND2_X1 U9592 ( .A1(n13030), .A2(n10668), .ZN(n10696) );
  NAND2_X1 U9593 ( .A1(n8024), .A2(n14863), .ZN(n12976) );
  AND2_X1 U9594 ( .A1(n7946), .A2(n7945), .ZN(n12888) );
  NAND2_X2 U9595 ( .A1(n7399), .A2(n7398), .ZN(n8025) );
  INV_X1 U9596 ( .A(n14836), .ZN(n14825) );
  AND2_X1 U9597 ( .A1(n10133), .A2(n10132), .ZN(n14820) );
  AND2_X1 U9598 ( .A1(n14746), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14841) );
  INV_X1 U9599 ( .A(n13254), .ZN(n14856) );
  INV_X1 U9600 ( .A(n10696), .ZN(n10481) );
  AND2_X1 U9601 ( .A1(n9951), .A2(n14880), .ZN(n10290) );
  INV_X1 U9602 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7386) );
  AND2_X1 U9603 ( .A1(n10737), .A2(n11056), .ZN(n13529) );
  AND4_X1 U9604 ( .A1(n9680), .A2(n9679), .A3(n9678), .A4(n9677), .ZN(n9681)
         );
  INV_X1 U9605 ( .A(n13688), .ZN(n14597) );
  INV_X1 U9606 ( .A(n13993), .ZN(n13983) );
  NAND2_X1 U9607 ( .A1(n10313), .A2(n10312), .ZN(n13761) );
  NAND2_X1 U9608 ( .A1(n10593), .A2(n10589), .ZN(n14726) );
  INV_X1 U9609 ( .A(n14708), .ZN(n14077) );
  AND2_X1 U9610 ( .A1(n14703), .A2(n14704), .ZN(n14525) );
  OR2_X1 U9611 ( .A1(n10749), .A2(n10748), .ZN(n13762) );
  INV_X1 U9612 ( .A(n14277), .ZN(n10311) );
  INV_X1 U9613 ( .A(n11257), .ZN(n9720) );
  AND2_X1 U9614 ( .A1(n9421), .A2(n9430), .ZN(n14596) );
  AND2_X1 U9615 ( .A1(n14380), .A2(n14381), .ZN(n14565) );
  AND2_X1 U9616 ( .A1(n9114), .A2(n9113), .ZN(n14983) );
  INV_X1 U9617 ( .A(n12437), .ZN(n11810) );
  INV_X1 U9618 ( .A(n12424), .ZN(n12434) );
  NAND2_X1 U9619 ( .A1(n10574), .A2(n10573), .ZN(n12439) );
  INV_X1 U9620 ( .A(n12596), .ZN(n12570) );
  NAND2_X1 U9621 ( .A1(n8734), .A2(n8733), .ZN(n12663) );
  INV_X1 U9622 ( .A(n12247), .ZN(n14452) );
  INV_X1 U9623 ( .A(n14963), .ZN(n15015) );
  INV_X1 U9624 ( .A(n14983), .ZN(n15005) );
  OR2_X1 U9625 ( .A1(n9159), .A2(n9158), .ZN(n15017) );
  NOR2_X1 U9626 ( .A1(n9895), .A2(n9894), .ZN(n9896) );
  INV_X1 U9627 ( .A(n15166), .ZN(n15163) );
  AND2_X2 U9628 ( .A1(n10817), .A2(n9891), .ZN(n15166) );
  INV_X1 U9629 ( .A(n15146), .ZN(n15144) );
  NAND2_X1 U9630 ( .A1(n9854), .A2(n9853), .ZN(n10813) );
  INV_X1 U9631 ( .A(SI_23_), .ZN(n11578) );
  INV_X1 U9632 ( .A(SI_17_), .ZN(n10723) );
  INV_X1 U9633 ( .A(SI_11_), .ZN(n10088) );
  INV_X1 U9634 ( .A(n14923), .ZN(n10054) );
  NAND2_X1 U9635 ( .A1(n8002), .A2(n13434), .ZN(n10118) );
  AND2_X1 U9636 ( .A1(n8047), .A2(n8046), .ZN(n8048) );
  INV_X1 U9637 ( .A(n12992), .ZN(n12961) );
  INV_X1 U9638 ( .A(n12976), .ZN(n12994) );
  OR2_X1 U9639 ( .A1(n8299), .A2(n8298), .ZN(n8300) );
  INV_X1 U9640 ( .A(n12888), .ZN(n13005) );
  INV_X1 U9641 ( .A(n12968), .ZN(n13014) );
  INV_X1 U9642 ( .A(n14841), .ZN(n10396) );
  OR2_X1 U9643 ( .A1(n10133), .A2(P2_U3088), .ZN(n14845) );
  AND2_X1 U9644 ( .A1(n11496), .A2(n11495), .ZN(n14895) );
  AND2_X1 U9645 ( .A1(n11236), .A2(n11235), .ZN(n14887) );
  NAND2_X1 U9646 ( .A1(n14868), .A2(n9956), .ZN(n13254) );
  INV_X1 U9647 ( .A(n13351), .ZN(n13374) );
  INV_X2 U9648 ( .A(n14903), .ZN(n14900) );
  AND2_X1 U9649 ( .A1(n14895), .A2(n14894), .ZN(n14902) );
  AND2_X2 U9650 ( .A1(n10290), .A2(n10289), .ZN(n14898) );
  NOR2_X1 U9651 ( .A1(n14877), .A2(n14870), .ZN(n14873) );
  INV_X1 U9652 ( .A(n14873), .ZN(n14874) );
  INV_X1 U9653 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11531) );
  INV_X1 U9654 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10440) );
  INV_X1 U9655 ( .A(n13875), .ZN(n14066) );
  INV_X1 U9656 ( .A(n13555), .ZN(n13526) );
  OR2_X1 U9657 ( .A1(n9481), .A2(n9480), .ZN(n13984) );
  INV_X1 U9658 ( .A(n12051), .ZN(n13982) );
  OR2_X1 U9659 ( .A1(n10596), .A2(n10034), .ZN(n13573) );
  INV_X1 U9660 ( .A(n14595), .ZN(n13677) );
  AND2_X1 U9661 ( .A1(n13842), .A2(n13841), .ZN(n14052) );
  AND2_X1 U9662 ( .A1(n11838), .A2(n11837), .ZN(n14534) );
  NAND2_X1 U9663 ( .A1(n13962), .A2(n11058), .ZN(n14008) );
  INV_X1 U9664 ( .A(n14745), .ZN(n14742) );
  AND3_X1 U9665 ( .A1(n14534), .A2(n14533), .A3(n14532), .ZN(n14548) );
  OR2_X1 U9666 ( .A1(n13762), .A2(n10750), .ZN(n14731) );
  NAND2_X1 U9667 ( .A1(n10107), .A2(n11056), .ZN(n14651) );
  INV_X1 U9668 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11207) );
  INV_X2 U9669 ( .A(n12443), .ZN(P3_U3897) );
  NOR2_X1 U9670 ( .A1(n10118), .A2(n10032), .ZN(P2_U3947) );
  NAND2_X1 U9671 ( .A1(n7337), .A2(n10031), .ZN(P2_U3236) );
  INV_X1 U9672 ( .A(n13573), .ZN(P1_U4016) );
  NOR2_X2 U9673 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7427) );
  NAND3_X1 U9674 ( .A1(n6447), .A2(n7448), .A3(n7349), .ZN(n7388) );
  NOR2_X1 U9675 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n7351) );
  NOR2_X1 U9676 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n7350) );
  NOR2_X1 U9677 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n7356) );
  NOR2_X1 U9678 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n7355) );
  NAND2_X1 U9679 ( .A1(n7358), .A2(n7357), .ZN(n7394) );
  NAND2_X1 U9680 ( .A1(n7361), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7359) );
  NAND2_X1 U9681 ( .A1(n7368), .A2(SI_1_), .ZN(n7419) );
  NAND2_X1 U9682 ( .A1(n7370), .A2(n7369), .ZN(n7371) );
  INV_X1 U9683 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9191) );
  INV_X1 U9684 ( .A(SI_0_), .ZN(n9190) );
  NOR2_X1 U9685 ( .A1(n7372), .A2(n9190), .ZN(n7374) );
  NAND2_X1 U9686 ( .A1(n7373), .A2(n7374), .ZN(n7420) );
  INV_X1 U9687 ( .A(n7374), .ZN(n7375) );
  NAND2_X1 U9688 ( .A1(n7376), .A2(n7375), .ZN(n7377) );
  NAND2_X1 U9689 ( .A1(n7420), .A2(n7377), .ZN(n10050) );
  AND2_X2 U9690 ( .A1(n6432), .A2(n7438), .ZN(n7447) );
  NAND2_X1 U9691 ( .A1(n7447), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7380) );
  NAND2_X1 U9692 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7378) );
  XNOR2_X1 U9693 ( .A(n7378), .B(P2_IR_REG_1__SCAN_IN), .ZN(n14749) );
  NAND2_X1 U9694 ( .A1(n7790), .A2(n14749), .ZN(n7379) );
  XNOR2_X2 U9695 ( .A(n7381), .B(n7991), .ZN(n11815) );
  NAND2_X1 U9696 ( .A1(n7385), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7387) );
  XNOR2_X1 U9697 ( .A(n11815), .B(n9955), .ZN(n7392) );
  NOR2_X2 U9698 ( .A1(n7661), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n7680) );
  AOI21_X1 U9699 ( .B1(n7680), .B2(n7389), .A(n7677), .ZN(n7390) );
  INV_X1 U9700 ( .A(n7390), .ZN(n7391) );
  XNOR2_X1 U9701 ( .A(n7391), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8022) );
  NAND2_X4 U9702 ( .A1(n9954), .A2(n8290), .ZN(n7987) );
  NAND2_X1 U9703 ( .A1(n7394), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7393) );
  NOR2_X2 U9704 ( .A1(n7394), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n7396) );
  INV_X1 U9705 ( .A(n7396), .ZN(n13422) );
  OR2_X2 U9706 ( .A1(n7396), .A2(n7677), .ZN(n7397) );
  XNOR2_X2 U9707 ( .A(n7397), .B(P2_IR_REG_30__SCAN_IN), .ZN(n7398) );
  NAND2_X2 U9708 ( .A1(n7398), .A2(n13427), .ZN(n8205) );
  INV_X1 U9709 ( .A(n8205), .ZN(n7921) );
  NAND2_X1 U9710 ( .A1(n7921), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7403) );
  INV_X2 U9711 ( .A(n8025), .ZN(n7453) );
  INV_X2 U9712 ( .A(n7398), .ZN(n12033) );
  AND2_X2 U9713 ( .A1(n12033), .A2(n13427), .ZN(n7512) );
  NAND2_X1 U9714 ( .A1(n7512), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7400) );
  NAND2_X1 U9715 ( .A1(n6429), .A2(n7799), .ZN(n7412) );
  INV_X1 U9716 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n14750) );
  NAND2_X1 U9717 ( .A1(n10049), .A2(SI_0_), .ZN(n7404) );
  XNOR2_X1 U9718 ( .A(n8426), .B(n7404), .ZN(n13441) );
  MUX2_X1 U9719 ( .A(n14750), .B(n13441), .S(n10114), .Z(n10018) );
  NAND2_X1 U9720 ( .A1(n10018), .A2(n7918), .ZN(n10689) );
  NAND2_X1 U9721 ( .A1(n7453), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7409) );
  NAND2_X1 U9722 ( .A1(n7512), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7408) );
  INV_X1 U9723 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7405) );
  NAND2_X1 U9724 ( .A1(n10481), .A2(n7779), .ZN(n10665) );
  INV_X1 U9725 ( .A(n7410), .ZN(n7411) );
  NAND2_X1 U9726 ( .A1(n7412), .A2(n7411), .ZN(n7413) );
  NAND2_X1 U9727 ( .A1(n10690), .A2(n7413), .ZN(n7431) );
  NAND2_X1 U9728 ( .A1(n8204), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7418) );
  NAND2_X1 U9729 ( .A1(n7453), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7417) );
  INV_X1 U9730 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7414) );
  OR2_X1 U9731 ( .A1(n8205), .A2(n7414), .ZN(n7416) );
  NAND2_X1 U9732 ( .A1(n7512), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n7415) );
  NAND4_X2 U9733 ( .A1(n7418), .A2(n7417), .A3(n7416), .A4(n7415), .ZN(n13029)
         );
  NAND2_X1 U9734 ( .A1(n13029), .A2(n7799), .ZN(n7434) );
  NAND2_X1 U9735 ( .A1(n7420), .A2(n7419), .ZN(n7425) );
  INV_X1 U9736 ( .A(n7425), .ZN(n7422) );
  MUX2_X1 U9737 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n7479), .Z(n7421) );
  NAND2_X1 U9738 ( .A1(n7421), .A2(SI_2_), .ZN(n7436) );
  NAND2_X1 U9739 ( .A1(n7422), .A2(n7423), .ZN(n7426) );
  INV_X1 U9740 ( .A(n7423), .ZN(n7424) );
  NAND2_X1 U9741 ( .A1(n7425), .A2(n7424), .ZN(n7437) );
  NAND2_X1 U9742 ( .A1(n7426), .A2(n7437), .ZN(n10082) );
  NAND2_X1 U9743 ( .A1(n7447), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7430) );
  OR2_X1 U9744 ( .A1(n7427), .A2(n7677), .ZN(n7428) );
  XNOR2_X1 U9745 ( .A(n7428), .B(P2_IR_REG_2__SCAN_IN), .ZN(n10143) );
  NAND2_X1 U9746 ( .A1(n7790), .A2(n10143), .ZN(n7429) );
  OAI211_X2 U9747 ( .C1(n8235), .C2(n10082), .A(n7430), .B(n7429), .ZN(n10622)
         );
  XNOR2_X1 U9748 ( .A(n10622), .B(n7987), .ZN(n7432) );
  XNOR2_X1 U9749 ( .A(n7434), .B(n7432), .ZN(n10850) );
  INV_X1 U9750 ( .A(n7432), .ZN(n7433) );
  NAND2_X1 U9751 ( .A1(n7434), .A2(n7433), .ZN(n7435) );
  NAND2_X1 U9752 ( .A1(n7437), .A2(n7436), .ZN(n7461) );
  NAND2_X1 U9753 ( .A1(n7439), .A2(SI_3_), .ZN(n7441) );
  OAI21_X1 U9754 ( .B1(n7439), .B2(SI_3_), .A(n7441), .ZN(n7462) );
  INV_X1 U9755 ( .A(n7462), .ZN(n7440) );
  NAND2_X1 U9756 ( .A1(n7461), .A2(n7440), .ZN(n7464) );
  NAND2_X1 U9757 ( .A1(n7464), .A2(n7441), .ZN(n7445) );
  MUX2_X1 U9758 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n7479), .Z(n7442) );
  NAND2_X1 U9759 ( .A1(n7442), .A2(SI_4_), .ZN(n7477) );
  OAI21_X1 U9760 ( .B1(n7442), .B2(SI_4_), .A(n7477), .ZN(n7443) );
  INV_X1 U9761 ( .A(n7443), .ZN(n7444) );
  NAND2_X1 U9762 ( .A1(n7445), .A2(n7444), .ZN(n7478) );
  OR2_X1 U9763 ( .A1(n7445), .A2(n7444), .ZN(n7446) );
  AND2_X1 U9764 ( .A1(n7478), .A2(n7446), .ZN(n10062) );
  INV_X2 U9765 ( .A(n8235), .ZN(n8216) );
  NAND2_X1 U9766 ( .A1(n10062), .A2(n8216), .ZN(n7451) );
  INV_X1 U9767 ( .A(n7555), .ZN(n7535) );
  NAND2_X1 U9768 ( .A1(n7448), .A2(n7459), .ZN(n7485) );
  NAND2_X1 U9769 ( .A1(n7485), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7449) );
  XNOR2_X1 U9770 ( .A(n7449), .B(P2_IR_REG_4__SCAN_IN), .ZN(n14763) );
  AOI22_X1 U9771 ( .A1(n7535), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n7790), .B2(
        n14763), .ZN(n7450) );
  NAND2_X1 U9772 ( .A1(n7451), .A2(n7450), .ZN(n10761) );
  XNOR2_X1 U9773 ( .A(n10761), .B(n7918), .ZN(n10649) );
  NAND2_X1 U9774 ( .A1(n7512), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n7458) );
  INV_X2 U9775 ( .A(n7452), .ZN(n8239) );
  NAND2_X1 U9776 ( .A1(n8239), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7457) );
  INV_X1 U9777 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10129) );
  INV_X1 U9778 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n14761) );
  NAND2_X1 U9779 ( .A1(n10129), .A2(n14761), .ZN(n7454) );
  NAND2_X1 U9780 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7490) );
  AND2_X1 U9781 ( .A1(n7454), .A2(n7490), .ZN(n10885) );
  NAND2_X1 U9782 ( .A1(n7966), .A2(n10885), .ZN(n7456) );
  INV_X4 U9783 ( .A(n8205), .ZN(n8240) );
  NAND2_X1 U9784 ( .A1(n8240), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7455) );
  NAND2_X1 U9785 ( .A1(n13027), .A2(n7779), .ZN(n10648) );
  NAND2_X1 U9786 ( .A1(n10649), .A2(n10648), .ZN(n7476) );
  OR2_X1 U9787 ( .A1(n7448), .A2(n7677), .ZN(n7460) );
  XNOR2_X1 U9788 ( .A(n7460), .B(n7459), .ZN(n10172) );
  OAI22_X1 U9789 ( .A1(n7555), .A2(n10076), .B1(n10114), .B2(n10172), .ZN(
        n7467) );
  INV_X1 U9790 ( .A(n7461), .ZN(n7463) );
  NAND2_X1 U9791 ( .A1(n7463), .A2(n7462), .ZN(n7465) );
  NAND2_X1 U9792 ( .A1(n7465), .A2(n7464), .ZN(n10077) );
  NOR2_X1 U9793 ( .A1(n10077), .A2(n8235), .ZN(n7466) );
  XNOR2_X1 U9794 ( .A(n10712), .B(n7918), .ZN(n10659) );
  NAND2_X1 U9795 ( .A1(n8204), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7471) );
  NAND2_X1 U9796 ( .A1(n8240), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7469) );
  INV_X2 U9797 ( .A(n7821), .ZN(n8241) );
  NAND2_X1 U9798 ( .A1(n7512), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n7468) );
  NAND2_X1 U9799 ( .A1(n13028), .A2(n7779), .ZN(n7472) );
  NAND2_X1 U9800 ( .A1(n10659), .A2(n7472), .ZN(n10402) );
  INV_X1 U9801 ( .A(n7472), .ZN(n7474) );
  INV_X1 U9802 ( .A(n10659), .ZN(n7473) );
  AND2_X1 U9803 ( .A1(n7474), .A2(n7473), .ZN(n10650) );
  INV_X1 U9804 ( .A(n10648), .ZN(n7475) );
  INV_X1 U9805 ( .A(n10649), .ZN(n12176) );
  AOI22_X1 U9806 ( .A1(n7476), .A2(n10650), .B1(n7475), .B2(n12176), .ZN(n7496) );
  MUX2_X1 U9807 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n10049), .Z(n7480) );
  NAND2_X1 U9808 ( .A1(n7480), .A2(SI_5_), .ZN(n7503) );
  OAI21_X1 U9809 ( .B1(n7480), .B2(SI_5_), .A(n7503), .ZN(n7481) );
  OR2_X1 U9810 ( .A1(n7483), .A2(n7482), .ZN(n7484) );
  NAND2_X1 U9811 ( .A1(n7504), .A2(n7484), .ZN(n10080) );
  OR2_X1 U9812 ( .A1(n10080), .A2(n8235), .ZN(n7488) );
  NAND2_X1 U9813 ( .A1(n7508), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7486) );
  XNOR2_X1 U9814 ( .A(n7486), .B(P2_IR_REG_5__SCAN_IN), .ZN(n13036) );
  AOI22_X1 U9815 ( .A1(n7535), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n7790), .B2(
        n13036), .ZN(n7487) );
  NAND2_X1 U9816 ( .A1(n7488), .A2(n7487), .ZN(n12171) );
  XNOR2_X1 U9817 ( .A(n12171), .B(n7987), .ZN(n7499) );
  NAND2_X1 U9818 ( .A1(n7512), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n7495) );
  NAND2_X1 U9819 ( .A1(n8239), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7494) );
  NOR2_X1 U9820 ( .A1(n7490), .A2(n7489), .ZN(n7513) );
  INV_X1 U9821 ( .A(n7513), .ZN(n7514) );
  NAND2_X1 U9822 ( .A1(n7490), .A2(n7489), .ZN(n7491) );
  AND2_X1 U9823 ( .A1(n7514), .A2(n7491), .ZN(n12182) );
  NAND2_X1 U9824 ( .A1(n7966), .A2(n12182), .ZN(n7493) );
  NAND2_X1 U9825 ( .A1(n8240), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7492) );
  NAND4_X1 U9826 ( .A1(n7495), .A2(n7494), .A3(n7493), .A4(n7492), .ZN(n13026)
         );
  NAND2_X1 U9827 ( .A1(n13026), .A2(n7779), .ZN(n7500) );
  XNOR2_X1 U9828 ( .A(n7499), .B(n7500), .ZN(n12177) );
  NAND2_X1 U9829 ( .A1(n7498), .A2(n7497), .ZN(n12184) );
  INV_X1 U9830 ( .A(n7499), .ZN(n7501) );
  NAND2_X1 U9831 ( .A1(n7501), .A2(n7500), .ZN(n7502) );
  INV_X1 U9832 ( .A(n7505), .ZN(n7506) );
  NAND2_X1 U9833 ( .A1(n7526), .A2(n7507), .ZN(n10075) );
  INV_X1 U9834 ( .A(n7508), .ZN(n7510) );
  NAND2_X1 U9835 ( .A1(n7510), .A2(n7509), .ZN(n7556) );
  NAND2_X1 U9836 ( .A1(n7556), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7532) );
  XNOR2_X1 U9837 ( .A(n7532), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10182) );
  AOI22_X1 U9838 ( .A1(n7535), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7790), .B2(
        n10182), .ZN(n7511) );
  NAND2_X1 U9839 ( .A1(n8241), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n7519) );
  NAND2_X1 U9840 ( .A1(n8239), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7518) );
  NAND2_X1 U9841 ( .A1(n7513), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7539) );
  INV_X1 U9842 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10766) );
  NAND2_X1 U9843 ( .A1(n7514), .A2(n10766), .ZN(n7515) );
  AND2_X1 U9844 ( .A1(n7539), .A2(n7515), .ZN(n11095) );
  NAND2_X1 U9845 ( .A1(n7966), .A2(n11095), .ZN(n7517) );
  NAND2_X1 U9846 ( .A1(n8240), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7516) );
  NAND4_X1 U9847 ( .A1(n7519), .A2(n7518), .A3(n7517), .A4(n7516), .ZN(n13025)
         );
  AND2_X1 U9848 ( .A1(n13025), .A2(n7779), .ZN(n7520) );
  NAND2_X1 U9849 ( .A1(n11042), .A2(n7520), .ZN(n7524) );
  INV_X1 U9850 ( .A(n7520), .ZN(n7521) );
  NAND2_X1 U9851 ( .A1(n7522), .A2(n7521), .ZN(n7523) );
  MUX2_X1 U9852 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n10049), .Z(n7527) );
  NAND2_X1 U9853 ( .A1(n7527), .A2(SI_7_), .ZN(n7549) );
  OAI21_X1 U9854 ( .B1(n7527), .B2(SI_7_), .A(n7549), .ZN(n7528) );
  INV_X1 U9855 ( .A(n7528), .ZN(n7529) );
  OR2_X1 U9856 ( .A1(n10093), .A2(n8235), .ZN(n7537) );
  NAND2_X1 U9857 ( .A1(n7532), .A2(n7531), .ZN(n7533) );
  NAND2_X1 U9858 ( .A1(n7533), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7534) );
  XNOR2_X1 U9859 ( .A(n7534), .B(P2_IR_REG_7__SCAN_IN), .ZN(n13052) );
  AOI22_X1 U9860 ( .A1(n7535), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7790), .B2(
        n13052), .ZN(n7536) );
  XNOR2_X1 U9861 ( .A(n11168), .B(n7987), .ZN(n7545) );
  NAND2_X1 U9862 ( .A1(n8241), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7544) );
  NAND2_X1 U9863 ( .A1(n8239), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7543) );
  INV_X1 U9864 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7538) );
  NAND2_X1 U9865 ( .A1(n7539), .A2(n7538), .ZN(n7540) );
  AND2_X1 U9866 ( .A1(n7561), .A2(n7540), .ZN(n14850) );
  NAND2_X1 U9867 ( .A1(n7966), .A2(n14850), .ZN(n7542) );
  NAND2_X1 U9868 ( .A1(n8240), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7541) );
  NAND4_X1 U9869 ( .A1(n7544), .A2(n7543), .A3(n7542), .A4(n7541), .ZN(n13024)
         );
  AND2_X1 U9870 ( .A1(n13024), .A2(n7779), .ZN(n7546) );
  NAND2_X1 U9871 ( .A1(n7545), .A2(n7546), .ZN(n7567) );
  INV_X1 U9872 ( .A(n7545), .ZN(n12216) );
  INV_X1 U9873 ( .A(n7546), .ZN(n7547) );
  NAND2_X1 U9874 ( .A1(n12216), .A2(n7547), .ZN(n7548) );
  AND2_X1 U9875 ( .A1(n7567), .A2(n7548), .ZN(n11044) );
  MUX2_X1 U9876 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n10049), .Z(n7550) );
  NAND2_X1 U9877 ( .A1(n7550), .A2(SI_8_), .ZN(n7572) );
  OAI21_X1 U9878 ( .B1(n7550), .B2(SI_8_), .A(n7572), .ZN(n7551) );
  INV_X1 U9879 ( .A(n7551), .ZN(n7552) );
  OR2_X1 U9880 ( .A1(n7553), .A2(n7552), .ZN(n7554) );
  NAND2_X1 U9881 ( .A1(n7573), .A2(n7554), .ZN(n10096) );
  OR2_X1 U9882 ( .A1(n10096), .A2(n8235), .ZN(n7559) );
  NAND2_X1 U9883 ( .A1(n7575), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7557) );
  XNOR2_X1 U9884 ( .A(n7557), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10188) );
  AOI22_X1 U9885 ( .A1(n7535), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7790), .B2(
        n10188), .ZN(n7558) );
  XNOR2_X1 U9886 ( .A(n14881), .B(n7987), .ZN(n11148) );
  NAND2_X1 U9887 ( .A1(n8241), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n7566) );
  NAND2_X1 U9888 ( .A1(n8239), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7565) );
  INV_X1 U9889 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7560) );
  NAND2_X1 U9890 ( .A1(n7561), .A2(n7560), .ZN(n7562) );
  NAND2_X1 U9891 ( .A1(n7580), .A2(n7562), .ZN(n12214) );
  INV_X1 U9892 ( .A(n12214), .ZN(n11241) );
  NAND2_X1 U9893 ( .A1(n7966), .A2(n11241), .ZN(n7564) );
  NAND2_X1 U9894 ( .A1(n8240), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7563) );
  NAND4_X1 U9895 ( .A1(n7566), .A2(n7565), .A3(n7564), .A4(n7563), .ZN(n13023)
         );
  NAND2_X1 U9896 ( .A1(n13023), .A2(n7779), .ZN(n7569) );
  XNOR2_X1 U9897 ( .A(n11148), .B(n7569), .ZN(n12219) );
  NAND2_X1 U9898 ( .A1(n11046), .A2(n7568), .ZN(n12224) );
  INV_X1 U9899 ( .A(n11148), .ZN(n7570) );
  NAND2_X1 U9900 ( .A1(n7570), .A2(n7569), .ZN(n7571) );
  NAND2_X1 U9901 ( .A1(n12224), .A2(n7571), .ZN(n7586) );
  MUX2_X1 U9902 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n10049), .Z(n7574) );
  NAND2_X1 U9903 ( .A1(n7574), .A2(SI_9_), .ZN(n7594) );
  OAI21_X1 U9904 ( .B1(n7574), .B2(SI_9_), .A(n7594), .ZN(n7591) );
  XNOR2_X1 U9905 ( .A(n7593), .B(n7591), .ZN(n10110) );
  NAND2_X1 U9906 ( .A1(n10110), .A2(n8216), .ZN(n7578) );
  NAND2_X1 U9907 ( .A1(n7600), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7576) );
  XNOR2_X1 U9908 ( .A(n7576), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10266) );
  AOI22_X1 U9909 ( .A1(n7535), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7790), .B2(
        n10266), .ZN(n7577) );
  XNOR2_X1 U9910 ( .A(n11543), .B(n7987), .ZN(n7587) );
  NAND2_X1 U9911 ( .A1(n8241), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7585) );
  NAND2_X1 U9912 ( .A1(n8239), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7584) );
  INV_X1 U9913 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7579) );
  INV_X1 U9914 ( .A(n7624), .ZN(n7622) );
  NAND2_X1 U9915 ( .A1(n7580), .A2(n7579), .ZN(n7581) );
  AND2_X1 U9916 ( .A1(n7622), .A2(n7581), .ZN(n11332) );
  NAND2_X1 U9917 ( .A1(n7966), .A2(n11332), .ZN(n7583) );
  NAND2_X1 U9918 ( .A1(n8240), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7582) );
  NAND4_X1 U9919 ( .A1(n7585), .A2(n7584), .A3(n7583), .A4(n7582), .ZN(n13022)
         );
  NAND2_X1 U9920 ( .A1(n13022), .A2(n7779), .ZN(n7588) );
  XNOR2_X1 U9921 ( .A(n7587), .B(n7588), .ZN(n11149) );
  NAND2_X1 U9922 ( .A1(n7586), .A2(n11149), .ZN(n11155) );
  INV_X1 U9923 ( .A(n7587), .ZN(n7589) );
  NAND2_X1 U9924 ( .A1(n7589), .A2(n7588), .ZN(n7590) );
  INV_X1 U9925 ( .A(n7591), .ZN(n7592) );
  MUX2_X1 U9926 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n10049), .Z(n7595) );
  NAND2_X1 U9927 ( .A1(n7595), .A2(SI_10_), .ZN(n7612) );
  OAI21_X1 U9928 ( .B1(n7595), .B2(SI_10_), .A(n7612), .ZN(n7596) );
  INV_X1 U9929 ( .A(n7596), .ZN(n7597) );
  OR2_X1 U9930 ( .A1(n7598), .A2(n7597), .ZN(n7599) );
  NAND2_X1 U9931 ( .A1(n7613), .A2(n7599), .ZN(n10207) );
  OR2_X1 U9932 ( .A1(n10207), .A2(n8235), .ZN(n7602) );
  OAI21_X1 U9933 ( .B1(n7600), .B2(P2_IR_REG_9__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7615) );
  XNOR2_X1 U9934 ( .A(n7615), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10386) );
  AOI22_X1 U9935 ( .A1(n8236), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7790), .B2(
        n10386), .ZN(n7601) );
  XNOR2_X1 U9936 ( .A(n11500), .B(n7987), .ZN(n7607) );
  NAND2_X1 U9937 ( .A1(n8241), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7606) );
  NAND2_X1 U9938 ( .A1(n8239), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7605) );
  XNOR2_X1 U9939 ( .A(n7622), .B(P2_REG3_REG_10__SCAN_IN), .ZN(n11499) );
  NAND2_X1 U9940 ( .A1(n7966), .A2(n11499), .ZN(n7604) );
  NAND2_X1 U9941 ( .A1(n8240), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7603) );
  NAND4_X1 U9942 ( .A1(n7606), .A2(n7605), .A3(n7604), .A4(n7603), .ZN(n13021)
         );
  AND2_X1 U9943 ( .A1(n13021), .A2(n7799), .ZN(n7608) );
  NAND2_X1 U9944 ( .A1(n7607), .A2(n7608), .ZN(n7630) );
  INV_X1 U9945 ( .A(n7607), .ZN(n12201) );
  INV_X1 U9946 ( .A(n7608), .ZN(n7609) );
  NAND2_X1 U9947 ( .A1(n12201), .A2(n7609), .ZN(n7610) );
  NAND2_X1 U9948 ( .A1(n7630), .A2(n7610), .ZN(n11453) );
  MUX2_X1 U9949 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n10049), .Z(n7636) );
  XNOR2_X1 U9950 ( .A(n7636), .B(SI_11_), .ZN(n7639) );
  XNOR2_X1 U9951 ( .A(n7640), .B(n7639), .ZN(n10282) );
  NAND2_X1 U9952 ( .A1(n10282), .A2(n8216), .ZN(n7619) );
  NAND2_X1 U9953 ( .A1(n7615), .A2(n7614), .ZN(n7616) );
  NAND2_X1 U9954 ( .A1(n7616), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7617) );
  XNOR2_X1 U9955 ( .A(n7617), .B(P2_IR_REG_11__SCAN_IN), .ZN(n13066) );
  AOI22_X1 U9956 ( .A1(n7447), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n13066), 
        .B2(n7790), .ZN(n7618) );
  XNOR2_X1 U9957 ( .A(n12208), .B(n7987), .ZN(n7632) );
  NAND2_X1 U9958 ( .A1(n8241), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n7629) );
  NAND2_X1 U9959 ( .A1(n8239), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7628) );
  INV_X1 U9960 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7621) );
  INV_X1 U9961 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7620) );
  OAI21_X1 U9962 ( .B1(n7622), .B2(n7621), .A(n7620), .ZN(n7625) );
  NAND2_X1 U9963 ( .A1(n7624), .A2(n7623), .ZN(n7644) );
  AND2_X1 U9964 ( .A1(n7625), .A2(n7644), .ZN(n12197) );
  NAND2_X1 U9965 ( .A1(n7966), .A2(n12197), .ZN(n7627) );
  NAND2_X1 U9966 ( .A1(n8240), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7626) );
  NAND4_X1 U9967 ( .A1(n7629), .A2(n7628), .A3(n7627), .A4(n7626), .ZN(n13020)
         );
  NAND2_X1 U9968 ( .A1(n13020), .A2(n7779), .ZN(n7633) );
  XNOR2_X1 U9969 ( .A(n7632), .B(n7633), .ZN(n12204) );
  INV_X1 U9970 ( .A(n7632), .ZN(n7634) );
  NAND2_X1 U9971 ( .A1(n7634), .A2(n7633), .ZN(n7635) );
  INV_X1 U9972 ( .A(n7636), .ZN(n7637) );
  NAND2_X1 U9973 ( .A1(n7637), .A2(n10088), .ZN(n7638) );
  MUX2_X1 U9974 ( .A(n10461), .B(n10440), .S(n10049), .Z(n7653) );
  XNOR2_X1 U9975 ( .A(n7656), .B(n7655), .ZN(n10439) );
  NAND2_X1 U9976 ( .A1(n10439), .A2(n8216), .ZN(n7643) );
  NAND2_X1 U9977 ( .A1(n7388), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7641) );
  XNOR2_X1 U9978 ( .A(n7641), .B(P2_IR_REG_12__SCAN_IN), .ZN(n10390) );
  AOI22_X1 U9979 ( .A1(n7447), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7790), .B2(
        n10390), .ZN(n7642) );
  XNOR2_X1 U9980 ( .A(n11643), .B(n7918), .ZN(n7650) );
  NAND2_X1 U9981 ( .A1(n8241), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7649) );
  NAND2_X1 U9982 ( .A1(n8239), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7648) );
  NAND2_X1 U9983 ( .A1(n7644), .A2(n11657), .ZN(n7645) );
  AND2_X1 U9984 ( .A1(n7688), .A2(n7645), .ZN(n11661) );
  NAND2_X1 U9985 ( .A1(n7966), .A2(n11661), .ZN(n7647) );
  NAND2_X1 U9986 ( .A1(n8240), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7646) );
  NAND4_X1 U9987 ( .A1(n7649), .A2(n7648), .A3(n7647), .A4(n7646), .ZN(n13019)
         );
  NAND2_X1 U9988 ( .A1(n13019), .A2(n7779), .ZN(n7651) );
  INV_X1 U9989 ( .A(n7650), .ZN(n11656) );
  INV_X1 U9990 ( .A(n7651), .ZN(n7652) );
  NAND2_X1 U9991 ( .A1(n11656), .A2(n7652), .ZN(n11653) );
  INV_X1 U9992 ( .A(n7653), .ZN(n7654) );
  MUX2_X1 U9993 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n10049), .Z(n7657) );
  NAND2_X1 U9994 ( .A1(n7657), .A2(SI_13_), .ZN(n7674) );
  OAI21_X1 U9995 ( .B1(n7657), .B2(SI_13_), .A(n7674), .ZN(n7659) );
  INV_X1 U9996 ( .A(n7659), .ZN(n7658) );
  NAND2_X1 U9997 ( .A1(n6735), .A2(n7659), .ZN(n7660) );
  NAND2_X1 U9998 ( .A1(n7675), .A2(n7660), .ZN(n10444) );
  NAND2_X1 U9999 ( .A1(n7661), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7663) );
  INV_X1 U10000 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n7662) );
  XNOR2_X1 U10001 ( .A(n7663), .B(n7662), .ZN(n11412) );
  INV_X1 U10002 ( .A(n11412), .ZN(n14794) );
  AOI22_X1 U10003 ( .A1(n7447), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7790), 
        .B2(n14794), .ZN(n7664) );
  XNOR2_X1 U10004 ( .A(n11666), .B(n7987), .ZN(n12185) );
  NAND2_X1 U10005 ( .A1(n8239), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7669) );
  XNOR2_X1 U10006 ( .A(n7688), .B(P2_REG3_REG_13__SCAN_IN), .ZN(n11750) );
  NAND2_X1 U10007 ( .A1(n7966), .A2(n11750), .ZN(n7668) );
  NAND2_X1 U10008 ( .A1(n8240), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7667) );
  NAND2_X1 U10009 ( .A1(n8241), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n7666) );
  NAND4_X1 U10010 ( .A1(n7669), .A2(n7668), .A3(n7667), .A4(n7666), .ZN(n13018) );
  AND2_X1 U10011 ( .A1(n13018), .A2(n7799), .ZN(n7670) );
  NAND2_X1 U10012 ( .A1(n12185), .A2(n7670), .ZN(n7694) );
  INV_X1 U10013 ( .A(n12185), .ZN(n7672) );
  INV_X1 U10014 ( .A(n7670), .ZN(n7671) );
  NAND2_X1 U10015 ( .A1(n7672), .A2(n7671), .ZN(n7673) );
  AND2_X1 U10016 ( .A1(n7694), .A2(n7673), .ZN(n11669) );
  MUX2_X1 U10017 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n10049), .Z(n7699) );
  XNOR2_X1 U10018 ( .A(n7699), .B(SI_14_), .ZN(n7702) );
  NAND2_X1 U10019 ( .A1(n10645), .A2(n8216), .ZN(n7684) );
  NOR2_X1 U10020 ( .A1(n7680), .A2(n7677), .ZN(n7676) );
  MUX2_X1 U10021 ( .A(n7677), .B(n7676), .S(P2_IR_REG_14__SCAN_IN), .Z(n7678)
         );
  INV_X1 U10022 ( .A(n7678), .ZN(n7682) );
  INV_X1 U10023 ( .A(n7705), .ZN(n7681) );
  AND2_X1 U10024 ( .A1(n7682), .A2(n7681), .ZN(n14801) );
  AOI22_X1 U10025 ( .A1(n7447), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7790), 
        .B2(n14801), .ZN(n7683) );
  XNOR2_X1 U10026 ( .A(n14480), .B(n7987), .ZN(n7696) );
  NAND2_X1 U10027 ( .A1(n8241), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n7693) );
  NAND2_X1 U10028 ( .A1(n8239), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7692) );
  NAND2_X1 U10029 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), 
        .ZN(n7685) );
  INV_X1 U10030 ( .A(n7709), .ZN(n7711) );
  INV_X1 U10031 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7687) );
  INV_X1 U10032 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7686) );
  OAI21_X1 U10033 ( .B1(n7688), .B2(n7687), .A(n7686), .ZN(n7689) );
  AND2_X1 U10034 ( .A1(n7711), .A2(n7689), .ZN(n14477) );
  NAND2_X1 U10035 ( .A1(n7966), .A2(n14477), .ZN(n7691) );
  NAND2_X1 U10036 ( .A1(n8240), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7690) );
  NAND4_X1 U10037 ( .A1(n7693), .A2(n7692), .A3(n7691), .A4(n7690), .ZN(n13017) );
  NAND2_X1 U10038 ( .A1(n13017), .A2(n7779), .ZN(n7697) );
  XNOR2_X1 U10039 ( .A(n7696), .B(n7697), .ZN(n12187) );
  INV_X1 U10040 ( .A(n7696), .ZN(n7698) );
  INV_X1 U10041 ( .A(n7699), .ZN(n7700) );
  NAND2_X1 U10042 ( .A1(n7700), .A2(n10321), .ZN(n7701) );
  MUX2_X1 U10043 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n10049), .Z(n7724) );
  XNOR2_X1 U10044 ( .A(n7724), .B(n10441), .ZN(n7722) );
  XNOR2_X1 U10045 ( .A(n7723), .B(n7722), .ZN(n10893) );
  NAND2_X1 U10046 ( .A1(n10893), .A2(n8216), .ZN(n7708) );
  NOR2_X1 U10047 ( .A1(n7705), .A2(n7677), .ZN(n7703) );
  MUX2_X1 U10048 ( .A(n7677), .B(n7703), .S(P2_IR_REG_15__SCAN_IN), .Z(n7706)
         );
  INV_X1 U10049 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n7704) );
  AND2_X1 U10050 ( .A1(n7705), .A2(n7704), .ZN(n7729) );
  NOR2_X1 U10051 ( .A1(n7706), .A2(n7729), .ZN(n14809) );
  AOI22_X1 U10052 ( .A1(n7447), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n7790), 
        .B2(n14809), .ZN(n7707) );
  XNOR2_X1 U10053 ( .A(n11860), .B(n7987), .ZN(n7718) );
  XNOR2_X1 U10054 ( .A(n7720), .B(n7718), .ZN(n11853) );
  NAND2_X1 U10055 ( .A1(n8241), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n7716) );
  NAND2_X1 U10056 ( .A1(n8239), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n7715) );
  NAND2_X1 U10057 ( .A1(n7709), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7733) );
  INV_X1 U10058 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7710) );
  NAND2_X1 U10059 ( .A1(n7711), .A2(n7710), .ZN(n7712) );
  AND2_X1 U10060 ( .A1(n7733), .A2(n7712), .ZN(n11898) );
  NAND2_X1 U10061 ( .A1(n7966), .A2(n11898), .ZN(n7714) );
  NAND2_X1 U10062 ( .A1(n8240), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n7713) );
  NAND4_X1 U10063 ( .A1(n7716), .A2(n7715), .A3(n7714), .A4(n7713), .ZN(n13016) );
  AND2_X1 U10064 ( .A1(n13016), .A2(n7799), .ZN(n7717) );
  INV_X1 U10065 ( .A(n7718), .ZN(n7719) );
  OR2_X1 U10066 ( .A1(n7720), .A2(n7719), .ZN(n7721) );
  INV_X1 U10067 ( .A(n7724), .ZN(n7725) );
  MUX2_X1 U10068 ( .A(n14181), .B(n10982), .S(n10049), .Z(n7744) );
  XNOR2_X1 U10069 ( .A(n7744), .B(SI_16_), .ZN(n7742) );
  XNOR2_X1 U10070 ( .A(n7743), .B(n7742), .ZN(n10981) );
  NAND2_X1 U10071 ( .A1(n10981), .A2(n8216), .ZN(n7732) );
  NOR2_X1 U10072 ( .A1(n7729), .A2(n7677), .ZN(n7726) );
  MUX2_X1 U10073 ( .A(n7677), .B(n7726), .S(P2_IR_REG_16__SCAN_IN), .Z(n7727)
         );
  INV_X1 U10074 ( .A(n7727), .ZN(n7730) );
  INV_X1 U10075 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n7728) );
  NAND2_X1 U10076 ( .A1(n7729), .A2(n7728), .ZN(n7767) );
  AND2_X1 U10077 ( .A1(n7730), .A2(n7767), .ZN(n14823) );
  AOI22_X1 U10078 ( .A1(n7790), .A2(n14823), .B1(n8236), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n7731) );
  XNOR2_X1 U10079 ( .A(n13285), .B(n7918), .ZN(n11962) );
  NAND2_X1 U10080 ( .A1(n8239), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7738) );
  NAND2_X1 U10081 ( .A1(n8240), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7737) );
  INV_X1 U10082 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n11971) );
  NAND2_X1 U10083 ( .A1(n7733), .A2(n11971), .ZN(n7734) );
  AND2_X1 U10084 ( .A1(n7751), .A2(n7734), .ZN(n11970) );
  NAND2_X1 U10085 ( .A1(n7966), .A2(n11970), .ZN(n7736) );
  NAND2_X1 U10086 ( .A1(n8241), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n7735) );
  NAND4_X1 U10087 ( .A1(n7738), .A2(n7737), .A3(n7736), .A4(n7735), .ZN(n13015) );
  NAND2_X1 U10088 ( .A1(n13015), .A2(n7779), .ZN(n7740) );
  XNOR2_X1 U10089 ( .A(n11962), .B(n7740), .ZN(n11969) );
  INV_X1 U10090 ( .A(n11969), .ZN(n7739) );
  NAND2_X1 U10091 ( .A1(n11962), .A2(n7740), .ZN(n7741) );
  NAND2_X1 U10092 ( .A1(n11959), .A2(n7741), .ZN(n7757) );
  NAND2_X1 U10093 ( .A1(n7744), .A2(n10587), .ZN(n7745) );
  MUX2_X1 U10094 ( .A(n11171), .B(n14123), .S(n10049), .Z(n7764) );
  XNOR2_X1 U10095 ( .A(n7763), .B(n7762), .ZN(n11104) );
  NAND2_X1 U10096 ( .A1(n11104), .A2(n8216), .ZN(n7749) );
  NAND2_X1 U10097 ( .A1(n7767), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7747) );
  XNOR2_X1 U10098 ( .A(n7747), .B(P2_IR_REG_17__SCAN_IN), .ZN(n11425) );
  AOI22_X1 U10099 ( .A1(n7447), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7790), 
        .B2(n11425), .ZN(n7748) );
  XNOR2_X1 U10100 ( .A(n13416), .B(n7918), .ZN(n7758) );
  INV_X1 U10101 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7750) );
  INV_X1 U10102 ( .A(n7771), .ZN(n7773) );
  NAND2_X1 U10103 ( .A1(n7751), .A2(n7750), .ZN(n7752) );
  NAND2_X1 U10104 ( .A1(n7773), .A2(n7752), .ZN(n13262) );
  OR2_X1 U10105 ( .A1(n8025), .A2(n13262), .ZN(n7756) );
  NAND2_X1 U10106 ( .A1(n8239), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7755) );
  NAND2_X1 U10107 ( .A1(n8241), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n7754) );
  INV_X1 U10108 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13263) );
  OR2_X1 U10109 ( .A1(n8205), .A2(n13263), .ZN(n7753) );
  NAND2_X1 U10110 ( .A1(n13014), .A2(n7779), .ZN(n7759) );
  XNOR2_X1 U10111 ( .A(n7758), .B(n7759), .ZN(n11960) );
  INV_X1 U10112 ( .A(n7758), .ZN(n7760) );
  NAND2_X1 U10113 ( .A1(n7760), .A2(n7759), .ZN(n7761) );
  NAND2_X1 U10114 ( .A1(n7764), .A2(n10723), .ZN(n7785) );
  NAND2_X1 U10115 ( .A1(n7788), .A2(n7785), .ZN(n7766) );
  MUX2_X1 U10116 ( .A(n11207), .B(n14112), .S(n10049), .Z(n7784) );
  XNOR2_X1 U10117 ( .A(n7784), .B(SI_18_), .ZN(n7765) );
  NAND2_X1 U10118 ( .A1(n11206), .A2(n8216), .ZN(n7770) );
  OAI21_X1 U10119 ( .B1(n7767), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7768) );
  XNOR2_X1 U10120 ( .A(n7768), .B(P2_IR_REG_18__SCAN_IN), .ZN(n14842) );
  AOI22_X1 U10121 ( .A1(n7790), .A2(n14842), .B1(n8236), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n7769) );
  XNOR2_X1 U10122 ( .A(n13359), .B(n7918), .ZN(n7780) );
  INV_X1 U10123 ( .A(n7793), .ZN(n7795) );
  INV_X1 U10124 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n7772) );
  NAND2_X1 U10125 ( .A1(n7773), .A2(n7772), .ZN(n7774) );
  NAND2_X1 U10126 ( .A1(n7795), .A2(n7774), .ZN(n13247) );
  NAND2_X1 U10127 ( .A1(n8241), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n7776) );
  NAND2_X1 U10128 ( .A1(n8239), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n7775) );
  AND2_X1 U10129 ( .A1(n7776), .A2(n7775), .ZN(n7778) );
  NAND2_X1 U10130 ( .A1(n8240), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n7777) );
  OAI211_X1 U10131 ( .C1(n13247), .C2(n8025), .A(n7778), .B(n7777), .ZN(n13013) );
  NAND2_X1 U10132 ( .A1(n13013), .A2(n7779), .ZN(n7781) );
  XNOR2_X1 U10133 ( .A(n7780), .B(n7781), .ZN(n12973) );
  INV_X1 U10134 ( .A(n7780), .ZN(n7783) );
  INV_X1 U10135 ( .A(n7781), .ZN(n7782) );
  OAI21_X1 U10136 ( .B1(n7789), .B2(SI_18_), .A(n7785), .ZN(n7786) );
  INV_X1 U10137 ( .A(n7786), .ZN(n7787) );
  MUX2_X1 U10138 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n10049), .Z(n7804) );
  XNOR2_X1 U10139 ( .A(n7806), .B(n7805), .ZN(n11264) );
  NAND2_X1 U10140 ( .A1(n11264), .A2(n8216), .ZN(n7792) );
  AOI22_X1 U10141 ( .A1(n7447), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7790), 
        .B2(n8022), .ZN(n7791) );
  XNOR2_X1 U10142 ( .A(n13229), .B(n7918), .ZN(n7801) );
  INV_X1 U10143 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n13231) );
  INV_X1 U10144 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n7794) );
  NAND2_X1 U10145 ( .A1(n7795), .A2(n7794), .ZN(n7796) );
  NAND2_X1 U10146 ( .A1(n7816), .A2(n7796), .ZN(n13230) );
  OR2_X1 U10147 ( .A1(n13230), .A2(n8025), .ZN(n7798) );
  AOI22_X1 U10148 ( .A1(n8204), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n8241), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n7797) );
  OAI211_X1 U10149 ( .C1(n8205), .C2(n13231), .A(n7798), .B(n7797), .ZN(n13012) );
  NAND2_X1 U10150 ( .A1(n13012), .A2(n7799), .ZN(n7802) );
  NAND2_X1 U10151 ( .A1(n7801), .A2(n7802), .ZN(n7800) );
  INV_X1 U10152 ( .A(n7801), .ZN(n12907) );
  INV_X1 U10153 ( .A(n7802), .ZN(n7803) );
  NAND2_X1 U10154 ( .A1(n12907), .A2(n7803), .ZN(n12903) );
  INV_X1 U10155 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11533) );
  MUX2_X1 U10156 ( .A(n11533), .B(n11531), .S(n10049), .Z(n7810) );
  NAND2_X1 U10157 ( .A1(n7811), .A2(n7810), .ZN(n7812) );
  NAND2_X1 U10158 ( .A1(n7827), .A2(n7812), .ZN(n11534) );
  NAND2_X1 U10159 ( .A1(n8236), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7813) );
  XNOR2_X1 U10160 ( .A(n13406), .B(n7918), .ZN(n7824) );
  INV_X1 U10161 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n7820) );
  INV_X1 U10162 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7815) );
  NAND2_X1 U10163 ( .A1(n7816), .A2(n7815), .ZN(n7817) );
  NAND2_X1 U10164 ( .A1(n7835), .A2(n7817), .ZN(n13217) );
  OR2_X1 U10165 ( .A1(n13217), .A2(n8025), .ZN(n7819) );
  AOI22_X1 U10166 ( .A1(n8239), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n8240), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n7818) );
  OAI211_X1 U10167 ( .C1(n7821), .C2(n7820), .A(n7819), .B(n7818), .ZN(n13011)
         );
  NAND2_X1 U10168 ( .A1(n13011), .A2(n7799), .ZN(n7823) );
  XNOR2_X1 U10169 ( .A(n7824), .B(n7823), .ZN(n12945) );
  INV_X1 U10170 ( .A(n12945), .ZN(n7822) );
  NAND2_X1 U10171 ( .A1(n7824), .A2(n7823), .ZN(n7825) );
  MUX2_X1 U10172 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n10049), .Z(n7828) );
  OAI21_X1 U10173 ( .B1(n7828), .B2(SI_21_), .A(n7846), .ZN(n7829) );
  INV_X1 U10174 ( .A(n7829), .ZN(n7830) );
  OR2_X1 U10175 ( .A1(n7831), .A2(n7830), .ZN(n7832) );
  NAND2_X1 U10176 ( .A1(n7847), .A2(n7832), .ZN(n11649) );
  NAND2_X1 U10177 ( .A1(n8236), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7833) );
  XNOR2_X1 U10178 ( .A(n13344), .B(n7987), .ZN(n7844) );
  INV_X1 U10179 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n12919) );
  NAND2_X1 U10180 ( .A1(n7835), .A2(n12919), .ZN(n7836) );
  NAND2_X1 U10181 ( .A1(n7879), .A2(n7836), .ZN(n13199) );
  INV_X1 U10182 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n7839) );
  NAND2_X1 U10183 ( .A1(n8241), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n7838) );
  NAND2_X1 U10184 ( .A1(n8240), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n7837) );
  OAI211_X1 U10185 ( .C1(n7452), .C2(n7839), .A(n7838), .B(n7837), .ZN(n7840)
         );
  INV_X1 U10186 ( .A(n7840), .ZN(n7841) );
  OAI21_X1 U10187 ( .B1(n13199), .B2(n8025), .A(n7841), .ZN(n13010) );
  NAND2_X1 U10188 ( .A1(n13010), .A2(n7799), .ZN(n7842) );
  XNOR2_X1 U10189 ( .A(n7844), .B(n7842), .ZN(n12917) );
  INV_X1 U10190 ( .A(n7842), .ZN(n7843) );
  NAND2_X1 U10191 ( .A1(n7844), .A2(n7843), .ZN(n7845) );
  INV_X1 U10192 ( .A(n7850), .ZN(n7849) );
  INV_X1 U10193 ( .A(SI_22_), .ZN(n7848) );
  INV_X1 U10194 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8341) );
  INV_X1 U10195 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11814) );
  MUX2_X1 U10196 ( .A(n8341), .B(n11814), .S(n10049), .Z(n7854) );
  NAND2_X1 U10197 ( .A1(n7853), .A2(n7854), .ZN(n7855) );
  NAND2_X1 U10198 ( .A1(n7872), .A2(n7855), .ZN(n11816) );
  NAND2_X1 U10199 ( .A1(n8236), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n7856) );
  XNOR2_X1 U10200 ( .A(n13192), .B(n7987), .ZN(n7863) );
  XNOR2_X1 U10201 ( .A(n7879), .B(P2_REG3_REG_22__SCAN_IN), .ZN(n13190) );
  NAND2_X1 U10202 ( .A1(n13190), .A2(n7966), .ZN(n7862) );
  INV_X1 U10203 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n14196) );
  NAND2_X1 U10204 ( .A1(n8241), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n7859) );
  NAND2_X1 U10205 ( .A1(n8240), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n7858) );
  OAI211_X1 U10206 ( .C1(n7452), .C2(n14196), .A(n7859), .B(n7858), .ZN(n7860)
         );
  INV_X1 U10207 ( .A(n7860), .ZN(n7861) );
  INV_X1 U10208 ( .A(n12896), .ZN(n13009) );
  NAND2_X1 U10209 ( .A1(n13009), .A2(n7799), .ZN(n12954) );
  INV_X1 U10210 ( .A(n7863), .ZN(n7864) );
  NOR2_X1 U10211 ( .A1(n7865), .A2(n7864), .ZN(n7866) );
  MUX2_X1 U10212 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n10049), .Z(n7868) );
  INV_X1 U10213 ( .A(n7868), .ZN(n7870) );
  AND2_X1 U10214 ( .A1(n7870), .A2(n7869), .ZN(n7871) );
  NAND2_X1 U10215 ( .A1(n7872), .A2(n7871), .ZN(n7873) );
  NAND2_X1 U10216 ( .A1(n7894), .A2(n11578), .ZN(n7874) );
  NAND2_X1 U10217 ( .A1(n8236), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7875) );
  XNOR2_X1 U10218 ( .A(n13174), .B(n7987), .ZN(n7888) );
  XNOR2_X1 U10219 ( .A(n7887), .B(n7888), .ZN(n12895) );
  NAND2_X1 U10220 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(P2_REG3_REG_23__SCAN_IN), 
        .ZN(n7877) );
  INV_X1 U10221 ( .A(n7903), .ZN(n7905) );
  INV_X1 U10222 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n12960) );
  INV_X1 U10223 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n7878) );
  OAI21_X1 U10224 ( .B1(n7879), .B2(n12960), .A(n7878), .ZN(n7880) );
  NAND2_X1 U10225 ( .A1(n7905), .A2(n7880), .ZN(n13171) );
  OR2_X1 U10226 ( .A1(n13171), .A2(n8025), .ZN(n7886) );
  INV_X1 U10227 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n7883) );
  NAND2_X1 U10228 ( .A1(n8241), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n7882) );
  NAND2_X1 U10229 ( .A1(n8240), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n7881) );
  OAI211_X1 U10230 ( .C1(n7452), .C2(n7883), .A(n7882), .B(n7881), .ZN(n7884)
         );
  INV_X1 U10231 ( .A(n7884), .ZN(n7885) );
  NAND2_X1 U10232 ( .A1(n12895), .A2(n7333), .ZN(n12894) );
  INV_X1 U10233 ( .A(n7888), .ZN(n7889) );
  NAND2_X2 U10234 ( .A1(n12894), .A2(n7890), .ZN(n12937) );
  NAND2_X1 U10235 ( .A1(n7891), .A2(n7895), .ZN(n7900) );
  MUX2_X1 U10236 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n10049), .Z(n7892) );
  NAND2_X1 U10237 ( .A1(n7892), .A2(SI_24_), .ZN(n7914) );
  OAI21_X1 U10238 ( .B1(SI_24_), .B2(n7892), .A(n7914), .ZN(n7896) );
  INV_X1 U10239 ( .A(n7896), .ZN(n7899) );
  OR2_X1 U10240 ( .A1(n11578), .A2(n7896), .ZN(n7893) );
  NOR2_X1 U10241 ( .A1(n7894), .A2(n7893), .ZN(n7898) );
  NOR2_X1 U10242 ( .A1(n7896), .A2(n7895), .ZN(n7897) );
  OR2_X1 U10243 ( .A1(n12019), .A2(n8235), .ZN(n7902) );
  NAND2_X1 U10244 ( .A1(n8236), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n7901) );
  XNOR2_X1 U10245 ( .A(n13398), .B(n7987), .ZN(n12925) );
  NAND2_X1 U10246 ( .A1(n7903), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n7919) );
  INV_X1 U10247 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n7904) );
  NAND2_X1 U10248 ( .A1(n7905), .A2(n7904), .ZN(n7906) );
  NAND2_X1 U10249 ( .A1(n7919), .A2(n7906), .ZN(n13159) );
  OR2_X1 U10250 ( .A1(n13159), .A2(n8025), .ZN(n7911) );
  INV_X1 U10251 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n13331) );
  NAND2_X1 U10252 ( .A1(n8241), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n7908) );
  NAND2_X1 U10253 ( .A1(n8240), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n7907) );
  OAI211_X1 U10254 ( .C1(n7452), .C2(n13331), .A(n7908), .B(n7907), .ZN(n7909)
         );
  INV_X1 U10255 ( .A(n7909), .ZN(n7910) );
  NAND2_X1 U10256 ( .A1(n13007), .A2(n7799), .ZN(n7912) );
  NOR2_X1 U10257 ( .A1(n12925), .A2(n7912), .ZN(n7913) );
  AOI21_X1 U10258 ( .B1(n12925), .B2(n7912), .A(n7913), .ZN(n12936) );
  MUX2_X1 U10259 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n10049), .Z(n7931) );
  XNOR2_X1 U10260 ( .A(n7931), .B(SI_25_), .ZN(n7934) );
  NAND2_X1 U10261 ( .A1(n13436), .A2(n8216), .ZN(n7917) );
  NAND2_X1 U10262 ( .A1(n8236), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7916) );
  XNOR2_X1 U10263 ( .A(n13394), .B(n7918), .ZN(n7927) );
  INV_X1 U10264 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n12931) );
  NAND2_X1 U10265 ( .A1(n7919), .A2(n12931), .ZN(n7920) );
  AND2_X1 U10266 ( .A1(n7939), .A2(n7920), .ZN(n13143) );
  NAND2_X1 U10267 ( .A1(n13143), .A2(n7966), .ZN(n7926) );
  INV_X1 U10268 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n13324) );
  NAND2_X1 U10269 ( .A1(n7921), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n7923) );
  NAND2_X1 U10270 ( .A1(n8241), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n7922) );
  OAI211_X1 U10271 ( .C1(n7452), .C2(n13324), .A(n7923), .B(n7922), .ZN(n7924)
         );
  INV_X1 U10272 ( .A(n7924), .ZN(n7925) );
  NOR2_X1 U10273 ( .A1(n12979), .A2(n13083), .ZN(n7928) );
  NAND2_X1 U10274 ( .A1(n7927), .A2(n7928), .ZN(n7947) );
  INV_X1 U10275 ( .A(n7927), .ZN(n12980) );
  INV_X1 U10276 ( .A(n7928), .ZN(n7929) );
  NAND2_X1 U10277 ( .A1(n12980), .A2(n7929), .ZN(n7930) );
  NAND2_X1 U10278 ( .A1(n7947), .A2(n7930), .ZN(n12926) );
  INV_X1 U10279 ( .A(n7931), .ZN(n7932) );
  INV_X1 U10280 ( .A(SI_25_), .ZN(n11907) );
  NAND2_X1 U10281 ( .A1(n7932), .A2(n11907), .ZN(n7933) );
  INV_X1 U10282 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14275) );
  INV_X1 U10283 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8351) );
  MUX2_X1 U10284 ( .A(n14275), .B(n8351), .S(n10049), .Z(n7952) );
  XNOR2_X1 U10285 ( .A(n7952), .B(SI_26_), .ZN(n7936) );
  XNOR2_X1 U10286 ( .A(n7955), .B(n7936), .ZN(n13432) );
  NAND2_X1 U10287 ( .A1(n13432), .A2(n8216), .ZN(n7938) );
  NAND2_X1 U10288 ( .A1(n8236), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n7937) );
  XNOR2_X1 U10289 ( .A(n13129), .B(n7987), .ZN(n7950) );
  INV_X1 U10290 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n12989) );
  INV_X1 U10291 ( .A(n7959), .ZN(n7961) );
  NAND2_X1 U10292 ( .A1(n7939), .A2(n12989), .ZN(n7940) );
  NAND2_X1 U10293 ( .A1(n7961), .A2(n7940), .ZN(n13126) );
  OR2_X1 U10294 ( .A1(n13126), .A2(n8025), .ZN(n7946) );
  INV_X1 U10295 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n7943) );
  NAND2_X1 U10296 ( .A1(n8241), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n7942) );
  NAND2_X1 U10297 ( .A1(n8240), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n7941) );
  OAI211_X1 U10298 ( .C1(n7452), .C2(n7943), .A(n7942), .B(n7941), .ZN(n7944)
         );
  INV_X1 U10299 ( .A(n7944), .ZN(n7945) );
  NAND2_X1 U10300 ( .A1(n13005), .A2(n7779), .ZN(n7949) );
  XNOR2_X1 U10301 ( .A(n7950), .B(n7949), .ZN(n12982) );
  INV_X1 U10302 ( .A(n7947), .ZN(n7948) );
  NAND2_X1 U10303 ( .A1(n7950), .A2(n7949), .ZN(n7951) );
  NOR2_X1 U10304 ( .A1(n7953), .A2(SI_26_), .ZN(n7954) );
  MUX2_X1 U10305 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n10049), .Z(n7970) );
  XNOR2_X1 U10306 ( .A(n7970), .B(SI_27_), .ZN(n7956) );
  NAND2_X1 U10307 ( .A1(n12023), .A2(n8216), .ZN(n7958) );
  NAND2_X1 U10308 ( .A1(n8236), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7957) );
  XNOR2_X1 U10309 ( .A(n13389), .B(n7987), .ZN(n7968) );
  INV_X1 U10310 ( .A(n7978), .ZN(n7979) );
  INV_X1 U10311 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n7960) );
  NAND2_X1 U10312 ( .A1(n7961), .A2(n7960), .ZN(n7962) );
  INV_X1 U10313 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n13315) );
  NAND2_X1 U10314 ( .A1(n8240), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n7964) );
  NAND2_X1 U10315 ( .A1(n8241), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n7963) );
  OAI211_X1 U10316 ( .C1(n7452), .C2(n13315), .A(n7964), .B(n7963), .ZN(n7965)
         );
  OR2_X1 U10317 ( .A1(n12985), .A2(n13083), .ZN(n7967) );
  NOR2_X1 U10318 ( .A1(n7968), .A2(n7967), .ZN(n7969) );
  AOI21_X1 U10319 ( .B1(n7968), .B2(n7967), .A(n7969), .ZN(n12886) );
  INV_X1 U10320 ( .A(n7970), .ZN(n7971) );
  INV_X1 U10321 ( .A(SI_27_), .ZN(n12881) );
  NOR2_X1 U10322 ( .A1(n7971), .A2(n12881), .ZN(n8186) );
  NAND2_X1 U10323 ( .A1(n7971), .A2(n12881), .ZN(n8190) );
  INV_X1 U10324 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12022) );
  INV_X1 U10325 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8358) );
  MUX2_X1 U10326 ( .A(n12022), .B(n8358), .S(n10049), .Z(n7972) );
  INV_X1 U10327 ( .A(SI_28_), .ZN(n12027) );
  NAND2_X1 U10328 ( .A1(n7972), .A2(n12027), .ZN(n8189) );
  INV_X1 U10329 ( .A(n7972), .ZN(n7973) );
  NAND2_X1 U10330 ( .A1(n7973), .A2(SI_28_), .ZN(n8211) );
  AND2_X1 U10331 ( .A1(n8189), .A2(n8211), .ZN(n7974) );
  NAND2_X1 U10332 ( .A1(n12021), .A2(n8216), .ZN(n7977) );
  NAND2_X1 U10333 ( .A1(n8236), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7976) );
  NAND2_X1 U10334 ( .A1(n7978), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n10024) );
  INV_X1 U10335 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8044) );
  NAND2_X1 U10336 ( .A1(n7979), .A2(n8044), .ZN(n7980) );
  NAND2_X1 U10337 ( .A1(n10024), .A2(n7980), .ZN(n13099) );
  OR2_X1 U10338 ( .A1(n13099), .A2(n8025), .ZN(n7985) );
  INV_X1 U10339 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13103) );
  NAND2_X1 U10340 ( .A1(n8241), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7982) );
  NAND2_X1 U10341 ( .A1(n8239), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n7981) );
  OAI211_X1 U10342 ( .C1(n13103), .C2(n8205), .A(n7982), .B(n7981), .ZN(n7983)
         );
  INV_X1 U10343 ( .A(n7983), .ZN(n7984) );
  NAND2_X1 U10344 ( .A1(n13003), .A2(n7799), .ZN(n7986) );
  XOR2_X1 U10345 ( .A(n7987), .B(n7986), .Z(n7988) );
  XNOR2_X1 U10346 ( .A(n13306), .B(n7988), .ZN(n7989) );
  XNOR2_X1 U10347 ( .A(n7990), .B(n7989), .ZN(n8049) );
  NAND2_X1 U10348 ( .A1(n8006), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7994) );
  MUX2_X1 U10349 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7994), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n7995) );
  INV_X1 U10350 ( .A(P2_B_REG_SCAN_IN), .ZN(n10012) );
  XNOR2_X1 U10351 ( .A(n12015), .B(n10012), .ZN(n7997) );
  NAND2_X1 U10352 ( .A1(n7998), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7996) );
  XNOR2_X1 U10353 ( .A(n7996), .B(P2_IR_REG_25__SCAN_IN), .ZN(n8018) );
  INV_X1 U10354 ( .A(n8018), .ZN(n13437) );
  NAND2_X1 U10355 ( .A1(n7997), .A2(n13437), .ZN(n8000) );
  INV_X1 U10356 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14876) );
  NOR2_X1 U10357 ( .A1(n13434), .A2(n12015), .ZN(n8001) );
  AOI21_X1 U10358 ( .B1(n14870), .B2(n14876), .A(n8001), .ZN(n9950) );
  INV_X1 U10359 ( .A(n8003), .ZN(n8004) );
  NAND2_X1 U10360 ( .A1(n8004), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8005) );
  MUX2_X1 U10361 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8005), .S(
        P2_IR_REG_23__SCAN_IN), .Z(n8007) );
  NAND2_X1 U10362 ( .A1(n8007), .A2(n8006), .ZN(n10112) );
  NAND2_X1 U10363 ( .A1(n9950), .A2(n14880), .ZN(n14875) );
  INV_X1 U10364 ( .A(n14875), .ZN(n10492) );
  NOR4_X1 U10365 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n8011) );
  NOR4_X1 U10366 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n8010) );
  NOR4_X1 U10367 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8009) );
  NOR4_X1 U10368 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n8008) );
  NAND4_X1 U10369 ( .A1(n8011), .A2(n8010), .A3(n8009), .A4(n8008), .ZN(n8017)
         );
  NOR2_X1 U10370 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .ZN(
        n8015) );
  NOR4_X1 U10371 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n8014) );
  NOR4_X1 U10372 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n8013) );
  NOR4_X1 U10373 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n8012) );
  NAND4_X1 U10374 ( .A1(n8015), .A2(n8014), .A3(n8013), .A4(n8012), .ZN(n8016)
         );
  OAI21_X1 U10375 ( .B1(n8017), .B2(n8016), .A(n14870), .ZN(n10288) );
  INV_X1 U10376 ( .A(n10288), .ZN(n8021) );
  INV_X1 U10377 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14878) );
  NAND2_X1 U10378 ( .A1(n14870), .A2(n14878), .ZN(n8020) );
  OR2_X1 U10379 ( .A1(n13434), .A2(n8018), .ZN(n8019) );
  NAND2_X1 U10380 ( .A1(n8020), .A2(n8019), .ZN(n14879) );
  NAND2_X1 U10381 ( .A1(n10492), .A2(n9952), .ZN(n8035) );
  AND2_X1 U10382 ( .A1(n10009), .A2(n8293), .ZN(n10113) );
  NAND2_X1 U10383 ( .A1(n12239), .A2(n11532), .ZN(n8296) );
  INV_X1 U10384 ( .A(n11532), .ZN(n8292) );
  AND2_X1 U10385 ( .A1(n11598), .A2(n8292), .ZN(n8289) );
  NAND2_X1 U10386 ( .A1(n11815), .A2(n8289), .ZN(n10022) );
  OR2_X1 U10387 ( .A1(n8035), .A2(n10022), .ZN(n8024) );
  INV_X1 U10388 ( .A(n10287), .ZN(n8023) );
  NAND2_X1 U10389 ( .A1(n8267), .A2(n12976), .ZN(n8047) );
  OR2_X1 U10390 ( .A1(n10024), .A2(n8025), .ZN(n8031) );
  INV_X1 U10391 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8028) );
  NAND2_X1 U10392 ( .A1(n8241), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8027) );
  NAND2_X1 U10393 ( .A1(n8240), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8026) );
  OAI211_X1 U10394 ( .C1(n7452), .C2(n8028), .A(n8027), .B(n8026), .ZN(n8029)
         );
  INV_X1 U10395 ( .A(n8029), .ZN(n8030) );
  AND2_X1 U10396 ( .A1(n8031), .A2(n8030), .ZN(n8219) );
  NAND2_X1 U10397 ( .A1(n10113), .A2(n8032), .ZN(n12984) );
  INV_X1 U10398 ( .A(n8032), .ZN(n8033) );
  NAND2_X1 U10399 ( .A1(n8033), .A2(n10113), .ZN(n12967) );
  OR2_X1 U10400 ( .A1(n12985), .A2(n12967), .ZN(n8034) );
  OAI21_X1 U10401 ( .B1(n8219), .B2(n12984), .A(n8034), .ZN(n13095) );
  INV_X1 U10402 ( .A(n8035), .ZN(n8037) );
  INV_X1 U10403 ( .A(n8296), .ZN(n8036) );
  INV_X1 U10404 ( .A(n9952), .ZN(n8039) );
  INV_X1 U10405 ( .A(n9950), .ZN(n8038) );
  OAI21_X1 U10406 ( .B1(n8039), .B2(n8038), .A(n10287), .ZN(n8043) );
  INV_X1 U10407 ( .A(n10490), .ZN(n8040) );
  AND2_X1 U10408 ( .A1(n8041), .A2(n8040), .ZN(n8042) );
  NAND2_X1 U10409 ( .A1(n8043), .A2(n8042), .ZN(n10667) );
  OAI22_X1 U10410 ( .A1(n13099), .A2(n12990), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8044), .ZN(n8045) );
  AOI21_X1 U10411 ( .B1(n13095), .B2(n12992), .A(n8045), .ZN(n8046) );
  OAI21_X1 U10412 ( .B1(n8049), .B2(n12971), .A(n8048), .ZN(P2_U3192) );
  NAND2_X1 U10413 ( .A1(n11815), .A2(n8022), .ZN(n8050) );
  AND2_X1 U10414 ( .A1(n8050), .A2(n9955), .ZN(n8051) );
  AOI21_X1 U10415 ( .B1(n10668), .B2(n8096), .A(n8051), .ZN(n8054) );
  NAND3_X1 U10416 ( .A1(n13030), .A2(n8061), .A3(n10018), .ZN(n8053) );
  NAND2_X1 U10417 ( .A1(n10668), .A2(n8051), .ZN(n8052) );
  OAI211_X1 U10418 ( .C1(n13030), .C2(n8054), .A(n8053), .B(n8052), .ZN(n8057)
         );
  MUX2_X1 U10419 ( .A(n6429), .B(n10967), .S(n8096), .Z(n8056) );
  OAI21_X1 U10420 ( .B1(n8057), .B2(n8058), .A(n8056), .ZN(n8060) );
  NAND2_X1 U10421 ( .A1(n8058), .A2(n8057), .ZN(n8059) );
  NAND2_X1 U10422 ( .A1(n8060), .A2(n8059), .ZN(n8064) );
  MUX2_X1 U10423 ( .A(n13029), .B(n10622), .S(n8262), .Z(n8065) );
  NAND2_X1 U10424 ( .A1(n8064), .A2(n8065), .ZN(n8063) );
  MUX2_X1 U10425 ( .A(n13029), .B(n10622), .S(n8074), .Z(n8062) );
  NAND2_X1 U10426 ( .A1(n8063), .A2(n8062), .ZN(n8069) );
  INV_X1 U10427 ( .A(n8064), .ZN(n8067) );
  INV_X1 U10428 ( .A(n8065), .ZN(n8066) );
  NAND2_X1 U10429 ( .A1(n8067), .A2(n8066), .ZN(n8068) );
  MUX2_X1 U10430 ( .A(n10712), .B(n13028), .S(n8074), .Z(n8070) );
  INV_X1 U10431 ( .A(n8072), .ZN(n8073) );
  MUX2_X1 U10432 ( .A(n13027), .B(n10761), .S(n8262), .Z(n8078) );
  MUX2_X1 U10433 ( .A(n13027), .B(n10761), .S(n8074), .Z(n8075) );
  NAND2_X1 U10434 ( .A1(n8076), .A2(n8075), .ZN(n8081) );
  INV_X1 U10435 ( .A(n8077), .ZN(n8079) );
  NAND2_X1 U10436 ( .A1(n8079), .A2(n7094), .ZN(n8080) );
  MUX2_X1 U10437 ( .A(n12171), .B(n13026), .S(n8262), .Z(n8083) );
  MUX2_X1 U10438 ( .A(n12171), .B(n13026), .S(n8074), .Z(n8082) );
  INV_X1 U10439 ( .A(n8083), .ZN(n8084) );
  MUX2_X1 U10440 ( .A(n11096), .B(n13025), .S(n8074), .Z(n8088) );
  NAND2_X1 U10441 ( .A1(n8087), .A2(n8088), .ZN(n8086) );
  MUX2_X1 U10442 ( .A(n11096), .B(n13025), .S(n8262), .Z(n8085) );
  NAND2_X1 U10443 ( .A1(n8086), .A2(n8085), .ZN(n8092) );
  INV_X1 U10444 ( .A(n8087), .ZN(n8090) );
  INV_X1 U10445 ( .A(n8088), .ZN(n8089) );
  NAND2_X1 U10446 ( .A1(n8090), .A2(n8089), .ZN(n8091) );
  MUX2_X1 U10447 ( .A(n13024), .B(n11168), .S(n8074), .Z(n8095) );
  MUX2_X1 U10448 ( .A(n11168), .B(n13024), .S(n8074), .Z(n8093) );
  MUX2_X1 U10449 ( .A(n13023), .B(n14881), .S(n8262), .Z(n8099) );
  MUX2_X1 U10450 ( .A(n13023), .B(n14881), .S(n8074), .Z(n8097) );
  NAND2_X1 U10451 ( .A1(n8098), .A2(n8097), .ZN(n8101) );
  MUX2_X1 U10452 ( .A(n13022), .B(n11543), .S(n8074), .Z(n8103) );
  MUX2_X1 U10453 ( .A(n13022), .B(n11543), .S(n8262), .Z(n8102) );
  INV_X1 U10454 ( .A(n8103), .ZN(n8104) );
  MUX2_X1 U10455 ( .A(n13021), .B(n11500), .S(n8262), .Z(n8108) );
  NAND2_X1 U10456 ( .A1(n8107), .A2(n8108), .ZN(n8106) );
  MUX2_X1 U10457 ( .A(n13021), .B(n11500), .S(n8074), .Z(n8105) );
  NAND2_X1 U10458 ( .A1(n8106), .A2(n8105), .ZN(n8112) );
  INV_X1 U10459 ( .A(n8107), .ZN(n8110) );
  INV_X1 U10460 ( .A(n8108), .ZN(n8109) );
  NAND2_X1 U10461 ( .A1(n8110), .A2(n8109), .ZN(n8111) );
  MUX2_X1 U10462 ( .A(n13020), .B(n12208), .S(n8061), .Z(n8115) );
  MUX2_X1 U10463 ( .A(n13020), .B(n12208), .S(n8262), .Z(n8113) );
  MUX2_X1 U10464 ( .A(n13019), .B(n11643), .S(n8262), .Z(n8118) );
  MUX2_X1 U10465 ( .A(n13019), .B(n11643), .S(n8061), .Z(n8116) );
  NAND2_X1 U10466 ( .A1(n8117), .A2(n8116), .ZN(n8120) );
  NAND2_X1 U10467 ( .A1(n8120), .A2(n8119), .ZN(n8122) );
  MUX2_X1 U10468 ( .A(n13018), .B(n11666), .S(n8074), .Z(n8123) );
  MUX2_X1 U10469 ( .A(n13018), .B(n11666), .S(n8262), .Z(n8121) );
  MUX2_X1 U10470 ( .A(n13017), .B(n14480), .S(n8262), .Z(n8126) );
  MUX2_X1 U10471 ( .A(n13017), .B(n14480), .S(n8074), .Z(n8124) );
  NAND2_X1 U10472 ( .A1(n8125), .A2(n8124), .ZN(n8128) );
  MUX2_X1 U10473 ( .A(n13016), .B(n11860), .S(n8061), .Z(n8132) );
  NAND2_X1 U10474 ( .A1(n8131), .A2(n8132), .ZN(n8130) );
  MUX2_X1 U10475 ( .A(n13016), .B(n11860), .S(n8262), .Z(n8129) );
  NAND2_X1 U10476 ( .A1(n8130), .A2(n8129), .ZN(n8136) );
  INV_X1 U10477 ( .A(n8131), .ZN(n8134) );
  INV_X1 U10478 ( .A(n8132), .ZN(n8133) );
  NAND2_X1 U10479 ( .A1(n8134), .A2(n8133), .ZN(n8135) );
  MUX2_X1 U10480 ( .A(n13015), .B(n13285), .S(n8262), .Z(n8138) );
  MUX2_X1 U10481 ( .A(n12968), .B(n13416), .S(n8074), .Z(n8140) );
  AND2_X1 U10482 ( .A1(n13265), .A2(n13014), .ZN(n9937) );
  OAI22_X1 U10483 ( .A1(n8139), .A2(n8138), .B1(n8140), .B2(n9937), .ZN(n8145)
         );
  INV_X1 U10484 ( .A(n13015), .ZN(n11961) );
  INV_X1 U10485 ( .A(n13285), .ZN(n13421) );
  MUX2_X1 U10486 ( .A(n11961), .B(n13421), .S(n8074), .Z(n8137) );
  AOI21_X1 U10487 ( .B1(n8139), .B2(n8138), .A(n8137), .ZN(n8144) );
  INV_X1 U10488 ( .A(n8140), .ZN(n8142) );
  NOR2_X1 U10489 ( .A1(n13265), .A2(n13014), .ZN(n8141) );
  OR2_X1 U10490 ( .A1(n8142), .A2(n8141), .ZN(n8143) );
  MUX2_X1 U10491 ( .A(n13013), .B(n13359), .S(n8262), .Z(n8149) );
  NAND2_X1 U10492 ( .A1(n8148), .A2(n8149), .ZN(n8147) );
  MUX2_X1 U10493 ( .A(n13013), .B(n13359), .S(n8074), .Z(n8146) );
  NAND2_X1 U10494 ( .A1(n8147), .A2(n8146), .ZN(n8153) );
  INV_X1 U10495 ( .A(n8148), .ZN(n8151) );
  INV_X1 U10496 ( .A(n8149), .ZN(n8150) );
  NAND2_X1 U10497 ( .A1(n8151), .A2(n8150), .ZN(n8152) );
  NAND2_X1 U10498 ( .A1(n8153), .A2(n8152), .ZN(n8155) );
  MUX2_X1 U10499 ( .A(n13012), .B(n13229), .S(n8061), .Z(n8156) );
  MUX2_X1 U10500 ( .A(n13012), .B(n13229), .S(n8262), .Z(n8154) );
  MUX2_X1 U10501 ( .A(n13011), .B(n13406), .S(n8262), .Z(n8160) );
  MUX2_X1 U10502 ( .A(n13011), .B(n13406), .S(n8074), .Z(n8157) );
  NAND2_X1 U10503 ( .A1(n8158), .A2(n8157), .ZN(n8162) );
  MUX2_X1 U10504 ( .A(n13010), .B(n13344), .S(n8061), .Z(n8165) );
  MUX2_X1 U10505 ( .A(n13010), .B(n13344), .S(n8262), .Z(n8163) );
  INV_X1 U10506 ( .A(n8165), .ZN(n8166) );
  MUX2_X1 U10507 ( .A(n13009), .B(n6770), .S(n8262), .Z(n8171) );
  MUX2_X1 U10508 ( .A(n13192), .B(n12896), .S(n8262), .Z(n8167) );
  NAND2_X1 U10509 ( .A1(n8169), .A2(n8168), .ZN(n8172) );
  MUX2_X1 U10510 ( .A(n13174), .B(n12959), .S(n8262), .Z(n8174) );
  MUX2_X1 U10511 ( .A(n13008), .B(n6769), .S(n8262), .Z(n8173) );
  MUX2_X1 U10512 ( .A(n13398), .B(n12924), .S(n8262), .Z(n8177) );
  MUX2_X1 U10513 ( .A(n13007), .B(n13162), .S(n8262), .Z(n8176) );
  MUX2_X1 U10514 ( .A(n12979), .B(n13394), .S(n8262), .Z(n8181) );
  MUX2_X1 U10515 ( .A(n13006), .B(n10001), .S(n8061), .Z(n8180) );
  NOR2_X1 U10516 ( .A1(n8181), .A2(n8180), .ZN(n8178) );
  AOI21_X1 U10517 ( .B1(n8177), .B2(n8176), .A(n8178), .ZN(n8175) );
  NOR3_X1 U10518 ( .A1(n8178), .A2(n8177), .A3(n8176), .ZN(n8179) );
  AOI21_X1 U10519 ( .B1(n8181), .B2(n8180), .A(n8179), .ZN(n8185) );
  MUX2_X1 U10520 ( .A(n13005), .B(n13318), .S(n8262), .Z(n8220) );
  INV_X1 U10521 ( .A(n8220), .ZN(n8183) );
  MUX2_X1 U10522 ( .A(n12888), .B(n13129), .S(n8061), .Z(n8221) );
  MUX2_X1 U10523 ( .A(n13003), .B(n8267), .S(n8262), .Z(n8223) );
  INV_X1 U10524 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n12030) );
  INV_X1 U10525 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13426) );
  MUX2_X1 U10526 ( .A(n12030), .B(n13426), .S(n10049), .Z(n8192) );
  XNOR2_X1 U10527 ( .A(n8192), .B(SI_29_), .ZN(n8213) );
  NAND2_X1 U10528 ( .A1(n8211), .A2(n8213), .ZN(n8191) );
  OR2_X1 U10529 ( .A1(n8186), .A2(n8191), .ZN(n8187) );
  AND2_X1 U10530 ( .A1(n8190), .A2(n8189), .ZN(n8209) );
  OR2_X1 U10531 ( .A1(n8191), .A2(n8209), .ZN(n8194) );
  INV_X1 U10532 ( .A(SI_29_), .ZN(n12041) );
  NAND2_X1 U10533 ( .A1(n8192), .A2(n12041), .ZN(n8193) );
  AND2_X1 U10534 ( .A1(n8194), .A2(n8193), .ZN(n8229) );
  MUX2_X1 U10535 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n10049), .Z(n8195) );
  NAND2_X1 U10536 ( .A1(n8195), .A2(SI_30_), .ZN(n8198) );
  OAI21_X1 U10537 ( .B1(n8195), .B2(SI_30_), .A(n8198), .ZN(n8231) );
  INV_X1 U10538 ( .A(n8231), .ZN(n8196) );
  MUX2_X1 U10539 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n10049), .Z(n8199) );
  XNOR2_X1 U10540 ( .A(n8199), .B(SI_31_), .ZN(n8200) );
  NAND2_X1 U10541 ( .A1(n14268), .A2(n8216), .ZN(n8203) );
  NAND2_X1 U10542 ( .A1(n7447), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8202) );
  NAND2_X1 U10543 ( .A1(n8204), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8208) );
  NAND2_X1 U10544 ( .A1(n8241), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8207) );
  OR2_X1 U10545 ( .A1(n8205), .A2(n14205), .ZN(n8206) );
  AND3_X1 U10546 ( .A1(n8208), .A2(n8207), .A3(n8206), .ZN(n8245) );
  XNOR2_X1 U10547 ( .A(n13378), .B(n8245), .ZN(n8250) );
  NAND2_X1 U10548 ( .A1(n8210), .A2(n8209), .ZN(n8212) );
  NAND2_X1 U10549 ( .A1(n8212), .A2(n8211), .ZN(n8215) );
  INV_X1 U10550 ( .A(n8213), .ZN(n8214) );
  NAND2_X1 U10551 ( .A1(n9669), .A2(n8216), .ZN(n8218) );
  NAND2_X1 U10552 ( .A1(n7447), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8217) );
  INV_X1 U10553 ( .A(n8219), .ZN(n13002) );
  MUX2_X1 U10554 ( .A(n8282), .B(n13002), .S(n8262), .Z(n8248) );
  MUX2_X1 U10555 ( .A(n12985), .B(n13389), .S(n8074), .Z(n8256) );
  INV_X1 U10556 ( .A(n12985), .ZN(n13004) );
  MUX2_X1 U10557 ( .A(n13004), .B(n13116), .S(n8096), .Z(n8255) );
  AOI22_X1 U10558 ( .A1(n8256), .A2(n8255), .B1(n8221), .B2(n8220), .ZN(n8222)
         );
  INV_X1 U10559 ( .A(n8250), .ZN(n8286) );
  INV_X1 U10560 ( .A(n8223), .ZN(n8228) );
  INV_X1 U10561 ( .A(n8224), .ZN(n8227) );
  INV_X1 U10562 ( .A(n8225), .ZN(n8226) );
  NAND4_X1 U10563 ( .A1(n8286), .A2(n8228), .A3(n8227), .A4(n8226), .ZN(n8253)
         );
  NAND2_X1 U10564 ( .A1(n8230), .A2(n8229), .ZN(n8232) );
  NAND2_X1 U10565 ( .A1(n8232), .A2(n8231), .ZN(n8233) );
  OR2_X1 U10566 ( .A1(n14272), .A2(n8235), .ZN(n8238) );
  NAND2_X1 U10567 ( .A1(n8236), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8237) );
  NAND2_X1 U10568 ( .A1(n8239), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8244) );
  NAND2_X1 U10569 ( .A1(n8240), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8243) );
  NAND2_X1 U10570 ( .A1(n8241), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8242) );
  AND3_X1 U10571 ( .A1(n8244), .A2(n8243), .A3(n8242), .ZN(n8283) );
  INV_X1 U10572 ( .A(n8245), .ZN(n13079) );
  OAI211_X1 U10573 ( .C1(n11815), .C2(n8292), .A(n8293), .B(n8296), .ZN(n8246)
         );
  AOI21_X1 U10574 ( .B1(n13079), .B2(n8262), .A(n8246), .ZN(n8247) );
  OAI22_X1 U10575 ( .A1(n13086), .A2(n8262), .B1(n8283), .B2(n8247), .ZN(n8258) );
  MUX2_X1 U10576 ( .A(n8283), .B(n13086), .S(n8262), .Z(n8259) );
  AOI22_X1 U10577 ( .A1(n8258), .A2(n8259), .B1(n8249), .B2(n8248), .ZN(n8251)
         );
  INV_X1 U10578 ( .A(n8254), .ZN(n8257) );
  NOR3_X1 U10579 ( .A1(n8257), .A2(n8256), .A3(n8255), .ZN(n8260) );
  OAI22_X1 U10580 ( .A1(n8261), .A2(n8260), .B1(n8259), .B2(n8258), .ZN(n8266)
         );
  MUX2_X1 U10581 ( .A(n13378), .B(n13079), .S(n8262), .Z(n8263) );
  INV_X1 U10582 ( .A(n8263), .ZN(n8264) );
  NAND2_X1 U10583 ( .A1(n8267), .A2(n12889), .ZN(n8268) );
  NOR2_X1 U10584 ( .A1(n13129), .A2(n13005), .ZN(n10002) );
  NOR2_X1 U10585 ( .A1(n13318), .A2(n12888), .ZN(n10004) );
  XNOR2_X1 U10586 ( .A(n6770), .B(n12896), .ZN(n13181) );
  INV_X1 U10587 ( .A(n13010), .ZN(n12958) );
  XNOR2_X1 U10588 ( .A(n13344), .B(n12958), .ZN(n13203) );
  INV_X1 U10589 ( .A(n13011), .ZN(n9996) );
  XNOR2_X1 U10590 ( .A(n13406), .B(n9996), .ZN(n13209) );
  INV_X1 U10591 ( .A(n13016), .ZN(n12188) );
  XNOR2_X1 U10592 ( .A(n11860), .B(n12188), .ZN(n11893) );
  XNOR2_X1 U10593 ( .A(n13285), .B(n11961), .ZN(n13277) );
  OR2_X1 U10594 ( .A1(n14480), .A2(n13017), .ZN(n9934) );
  NAND2_X1 U10595 ( .A1(n14480), .A2(n13017), .ZN(n9935) );
  INV_X1 U10596 ( .A(n13019), .ZN(n8269) );
  OR2_X1 U10597 ( .A1(n11643), .A2(n8269), .ZN(n9982) );
  NAND2_X1 U10598 ( .A1(n11643), .A2(n8269), .ZN(n8270) );
  INV_X1 U10599 ( .A(n13021), .ZN(n12200) );
  XNOR2_X1 U10600 ( .A(n11500), .B(n12200), .ZN(n11491) );
  INV_X1 U10601 ( .A(n13022), .ZN(n9976) );
  XNOR2_X1 U10602 ( .A(n11543), .B(n9976), .ZN(n11327) );
  INV_X1 U10603 ( .A(n13023), .ZN(n11144) );
  XNOR2_X1 U10604 ( .A(n14881), .B(n11144), .ZN(n11231) );
  XNOR2_X1 U10605 ( .A(n11168), .B(n13024), .ZN(n11162) );
  INV_X1 U10606 ( .A(n10761), .ZN(n10887) );
  XNOR2_X2 U10607 ( .A(n13028), .B(n11018), .ZN(n10702) );
  OAI21_X1 U10608 ( .B1(n13030), .B2(n10668), .A(n10696), .ZN(n14859) );
  NAND3_X1 U10609 ( .A1(n9915), .A2(n8292), .A3(n14859), .ZN(n8273) );
  INV_X1 U10610 ( .A(n10622), .ZN(n10956) );
  INV_X2 U10611 ( .A(n13029), .ZN(n8272) );
  XNOR2_X2 U10612 ( .A(n10622), .B(n8272), .ZN(n10611) );
  NOR4_X1 U10613 ( .A1(n10757), .A2(n10702), .A3(n8273), .A4(n10611), .ZN(
        n8274) );
  XNOR2_X1 U10614 ( .A(n11096), .B(n13025), .ZN(n9969) );
  XNOR2_X1 U10615 ( .A(n12171), .B(n13026), .ZN(n10863) );
  NAND4_X1 U10616 ( .A1(n11162), .A2(n8274), .A3(n9969), .A4(n10863), .ZN(
        n8275) );
  NOR4_X1 U10617 ( .A1(n11491), .A2(n11327), .A3(n11231), .A4(n8275), .ZN(
        n8276) );
  XNOR2_X1 U10618 ( .A(n11666), .B(n13018), .ZN(n11748) );
  XNOR2_X1 U10619 ( .A(n12208), .B(n13020), .ZN(n11620) );
  NAND4_X1 U10620 ( .A1(n11636), .A2(n8276), .A3(n11748), .A4(n11620), .ZN(
        n8277) );
  NOR4_X1 U10621 ( .A1(n11893), .A2(n13277), .A3(n14481), .A4(n8277), .ZN(
        n8278) );
  XNOR2_X1 U10622 ( .A(n13229), .B(n13012), .ZN(n13235) );
  XNOR2_X1 U10623 ( .A(n13359), .B(n13013), .ZN(n9938) );
  XNOR2_X1 U10624 ( .A(n13265), .B(n13014), .ZN(n13266) );
  NAND4_X1 U10625 ( .A1(n8278), .A2(n13235), .A3(n9938), .A4(n13266), .ZN(
        n8279) );
  NOR4_X1 U10626 ( .A1(n13181), .A2(n13203), .A3(n13209), .A4(n8279), .ZN(
        n8280) );
  NAND2_X1 U10627 ( .A1(n6769), .A2(n13008), .ZN(n9943) );
  NAND2_X1 U10628 ( .A1(n9944), .A2(n9943), .ZN(n13176) );
  NAND4_X1 U10629 ( .A1(n13131), .A2(n8280), .A3(n13176), .A4(n13150), .ZN(
        n8281) );
  XNOR2_X1 U10630 ( .A(n13116), .B(n12985), .ZN(n9948) );
  XOR2_X1 U10631 ( .A(n13006), .B(n10001), .Z(n13138) );
  NOR4_X1 U10632 ( .A1(n13090), .A2(n8281), .A3(n9948), .A4(n13138), .ZN(n8285) );
  XNOR2_X1 U10633 ( .A(n8282), .B(n13002), .ZN(n10006) );
  INV_X1 U10634 ( .A(n8283), .ZN(n13001) );
  XNOR2_X1 U10635 ( .A(n13382), .B(n13001), .ZN(n8284) );
  NAND4_X1 U10636 ( .A1(n8286), .A2(n8285), .A3(n10006), .A4(n8284), .ZN(n8287) );
  XOR2_X1 U10637 ( .A(n8287), .B(n8022), .Z(n8288) );
  OAI22_X1 U10638 ( .A1(n10009), .A2(n8290), .B1(n8289), .B2(n8022), .ZN(n8291) );
  INV_X1 U10639 ( .A(n14861), .ZN(n8294) );
  NAND2_X1 U10640 ( .A1(n8293), .A2(n8292), .ZN(n10010) );
  OAI22_X1 U10641 ( .A1(n8294), .A2(n11815), .B1(n10010), .B2(n12239), .ZN(
        n8295) );
  NOR2_X1 U10642 ( .A1(n10112), .A2(P2_U3088), .ZN(n12034) );
  INV_X1 U10643 ( .A(n14880), .ZN(n14877) );
  NOR4_X1 U10644 ( .A1(n14877), .A2(n12967), .A3(n12024), .A4(n8296), .ZN(
        n8299) );
  INV_X1 U10645 ( .A(n12034), .ZN(n8297) );
  OAI21_X1 U10646 ( .B1(n8297), .B2(n10009), .A(P2_B_REG_SCAN_IN), .ZN(n8298)
         );
  INV_X1 U10647 ( .A(n8433), .ZN(n8301) );
  XNOR2_X1 U10648 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8432) );
  NAND2_X1 U10649 ( .A1(n8301), .A2(n8432), .ZN(n8304) );
  INV_X1 U10650 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n8302) );
  NAND2_X1 U10651 ( .A1(n8302), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8303) );
  INV_X1 U10652 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10060) );
  NOR2_X1 U10653 ( .A1(n10060), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8305) );
  INV_X1 U10654 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10081) );
  NOR2_X1 U10655 ( .A1(n10076), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8307) );
  NAND2_X1 U10656 ( .A1(n10076), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8306) );
  NAND2_X1 U10657 ( .A1(n10063), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8309) );
  NAND2_X1 U10658 ( .A1(n10083), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8308) );
  NAND2_X1 U10659 ( .A1(n8309), .A2(n8308), .ZN(n8474) );
  NAND2_X1 U10660 ( .A1(n10061), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8312) );
  NAND2_X1 U10661 ( .A1(n10078), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8310) );
  NAND2_X1 U10662 ( .A1(n8312), .A2(n8310), .ZN(n8494) );
  INV_X1 U10663 ( .A(n8494), .ZN(n8311) );
  INV_X1 U10664 ( .A(n8516), .ZN(n8313) );
  NAND2_X1 U10665 ( .A1(n10094), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8316) );
  NAND2_X1 U10666 ( .A1(n10095), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8315) );
  INV_X1 U10667 ( .A(n8545), .ZN(n8317) );
  XNOR2_X1 U10668 ( .A(n8318), .B(P1_DATAO_REG_9__SCAN_IN), .ZN(n8557) );
  NAND2_X1 U10669 ( .A1(n8318), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8319) );
  XNOR2_X1 U10670 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n8564) );
  NAND2_X1 U10671 ( .A1(n8565), .A2(n8564), .ZN(n8322) );
  NAND2_X1 U10672 ( .A1(n8320), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8321) );
  NAND2_X1 U10673 ( .A1(n10461), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8324) );
  NAND2_X1 U10674 ( .A1(n10440), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n8323) );
  XNOR2_X1 U10675 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n8617) );
  INV_X1 U10676 ( .A(n8617), .ZN(n8327) );
  NAND2_X1 U10677 ( .A1(n10894), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8329) );
  INV_X1 U10678 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10940) );
  NAND2_X1 U10679 ( .A1(n10940), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8328) );
  NAND2_X1 U10680 ( .A1(n8329), .A2(n8328), .ZN(n8630) );
  NAND2_X1 U10681 ( .A1(n14181), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8331) );
  NAND2_X1 U10682 ( .A1(n10982), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8330) );
  XNOR2_X1 U10683 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .ZN(n8664) );
  NAND2_X1 U10684 ( .A1(n14123), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8332) );
  NAND2_X1 U10685 ( .A1(n11207), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8335) );
  NAND2_X1 U10686 ( .A1(n14112), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8334) );
  INV_X1 U10687 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11266) );
  NAND2_X1 U10688 ( .A1(n11266), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8337) );
  INV_X1 U10689 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11265) );
  NAND2_X1 U10690 ( .A1(n11265), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8336) );
  XNOR2_X1 U10691 ( .A(n11531), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n8709) );
  NAND2_X1 U10692 ( .A1(n11531), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8338) );
  INV_X1 U10693 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n14126) );
  NAND2_X1 U10694 ( .A1(n14126), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8340) );
  INV_X1 U10695 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11597) );
  NAND2_X1 U10696 ( .A1(n11597), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8339) );
  NAND2_X1 U10697 ( .A1(n8341), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8343) );
  NAND2_X1 U10698 ( .A1(n11814), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8342) );
  INV_X1 U10699 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8344) );
  XNOR2_X1 U10700 ( .A(n8344), .B(P2_DATAO_REG_23__SCAN_IN), .ZN(n8749) );
  NAND2_X1 U10701 ( .A1(n8345), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8346) );
  INV_X1 U10702 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n12016) );
  INV_X1 U10703 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14279) );
  NAND2_X1 U10704 ( .A1(n14279), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8350) );
  INV_X1 U10705 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13439) );
  NAND2_X1 U10706 ( .A1(n13439), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8348) );
  NAND2_X1 U10707 ( .A1(n8350), .A2(n8348), .ZN(n8773) );
  INV_X1 U10708 ( .A(n8773), .ZN(n8349) );
  NAND2_X1 U10709 ( .A1(n14275), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8354) );
  NAND2_X1 U10710 ( .A1(n8351), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8352) );
  NAND2_X1 U10711 ( .A1(n8354), .A2(n8352), .ZN(n8786) );
  INV_X1 U10712 ( .A(n8786), .ZN(n8353) );
  NAND2_X1 U10713 ( .A1(n8787), .A2(n8353), .ZN(n8355) );
  NAND2_X1 U10714 ( .A1(n8355), .A2(n8354), .ZN(n8799) );
  INV_X1 U10715 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14273) );
  NAND2_X1 U10716 ( .A1(n14273), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8357) );
  INV_X1 U10717 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n12025) );
  NAND2_X1 U10718 ( .A1(n12025), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8356) );
  AND2_X1 U10719 ( .A1(n8357), .A2(n8356), .ZN(n8798) );
  NAND2_X1 U10720 ( .A1(n8799), .A2(n8798), .ZN(n8801) );
  NAND2_X1 U10721 ( .A1(n12022), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8361) );
  NAND2_X1 U10722 ( .A1(n8358), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8359) );
  NAND2_X1 U10723 ( .A1(n8361), .A2(n8359), .ZN(n8813) );
  INV_X1 U10724 ( .A(n8813), .ZN(n8360) );
  NAND2_X1 U10725 ( .A1(n8814), .A2(n8360), .ZN(n8362) );
  NAND2_X1 U10726 ( .A1(n13426), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8363) );
  NAND2_X1 U10727 ( .A1(n8827), .A2(n8363), .ZN(n8365) );
  NAND2_X1 U10728 ( .A1(n12030), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8364) );
  NAND2_X1 U10729 ( .A1(n8365), .A2(n8364), .ZN(n8414) );
  INV_X1 U10730 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14271) );
  AND2_X1 U10731 ( .A1(n14271), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8366) );
  OAI22_X1 U10732 ( .A1(n8414), .A2(n8366), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n14271), .ZN(n8368) );
  XNOR2_X1 U10733 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n8367) );
  XNOR2_X1 U10734 ( .A(n8368), .B(n8367), .ZN(n12873) );
  NOR2_X1 U10735 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .ZN(
        n8371) );
  NOR2_X1 U10736 ( .A1(P3_IR_REG_25__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), 
        .ZN(n8378) );
  NOR2_X1 U10737 ( .A1(P3_IR_REG_24__SCAN_IN), .A2(P3_IR_REG_20__SCAN_IN), 
        .ZN(n8377) );
  INV_X1 U10738 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8381) );
  NAND2_X1 U10739 ( .A1(n9022), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8385) );
  INV_X1 U10740 ( .A(SI_31_), .ZN(n12877) );
  NOR2_X1 U10741 ( .A1(n8829), .A2(n12877), .ZN(n8386) );
  AOI21_X1 U10742 ( .B1(n12873), .B2(n8828), .A(n8386), .ZN(n12543) );
  INV_X1 U10743 ( .A(n12543), .ZN(n12818) );
  NOR2_X1 U10744 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8487) );
  NAND2_X1 U10745 ( .A1(n8487), .A2(n10679), .ZN(n8505) );
  NAND2_X1 U10746 ( .A1(n11945), .A2(n11981), .ZN(n8387) );
  INV_X1 U10747 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8388) );
  INV_X1 U10748 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n8392) );
  INV_X1 U10749 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n8394) );
  INV_X1 U10750 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n8396) );
  INV_X1 U10751 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8398) );
  INV_X1 U10752 ( .A(n8817), .ZN(n8400) );
  INV_X1 U10753 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n12326) );
  NAND2_X1 U10754 ( .A1(n8400), .A2(n12326), .ZN(n12541) );
  NAND2_X1 U10755 ( .A1(n8402), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8401) );
  MUX2_X1 U10756 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8401), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n8403) );
  NAND2_X1 U10757 ( .A1(n6426), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n8411) );
  NAND2_X1 U10758 ( .A1(n8455), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n8410) );
  INV_X1 U10759 ( .A(n12042), .ZN(n8407) );
  INV_X1 U10760 ( .A(n8440), .ZN(n8453) );
  NAND2_X1 U10761 ( .A1(n8440), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n8409) );
  AND3_X1 U10762 ( .A1(n8411), .A2(n8410), .A3(n8409), .ZN(n8412) );
  NAND2_X1 U10763 ( .A1(n8838), .A2(n8412), .ZN(n11269) );
  NAND2_X1 U10764 ( .A1(n12818), .A2(n12540), .ZN(n8987) );
  INV_X1 U10765 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12032) );
  XNOR2_X1 U10766 ( .A(n12032), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n8413) );
  XNOR2_X1 U10767 ( .A(n8414), .B(n8413), .ZN(n12244) );
  INV_X1 U10768 ( .A(SI_30_), .ZN(n12246) );
  NOR2_X1 U10769 ( .A1(n8829), .A2(n12246), .ZN(n8415) );
  INV_X1 U10770 ( .A(n12753), .ZN(n12822) );
  INV_X1 U10771 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n8418) );
  NAND2_X1 U10772 ( .A1(n8455), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8417) );
  NAND2_X1 U10773 ( .A1(n8440), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8416) );
  OAI211_X1 U10774 ( .C1(n8835), .C2(n8418), .A(n8417), .B(n8416), .ZN(n8419)
         );
  INV_X1 U10775 ( .A(n8419), .ZN(n8420) );
  OR2_X1 U10776 ( .A1(n12822), .A2(n9901), .ZN(n8421) );
  NAND2_X1 U10777 ( .A1(n8987), .A2(n8421), .ZN(n8983) );
  NAND2_X1 U10778 ( .A1(n6426), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8425) );
  NAND2_X1 U10779 ( .A1(n8440), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8423) );
  NAND2_X1 U10780 ( .A1(n8455), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8422) );
  OAI21_X1 U10781 ( .B1(P2_DATAO_REG_0__SCAN_IN), .B2(n8426), .A(n8433), .ZN(
        n8427) );
  MUX2_X1 U10782 ( .A(n8427), .B(SI_0_), .S(n10049), .Z(n12884) );
  MUX2_X1 U10783 ( .A(P3_IR_REG_0__SCAN_IN), .B(n12884), .S(n9799), .Z(n10818)
         );
  NAND2_X1 U10784 ( .A1(n6426), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8430) );
  NAND2_X1 U10785 ( .A1(n8440), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8429) );
  NAND2_X1 U10786 ( .A1(n8455), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8428) );
  XNOR2_X1 U10787 ( .A(n8433), .B(n8432), .ZN(n10065) );
  NAND2_X1 U10788 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n8434) );
  INV_X1 U10789 ( .A(n8445), .ZN(n8435) );
  NAND2_X1 U10790 ( .A1(n10566), .A2(n8865), .ZN(n10564) );
  NAND2_X1 U10791 ( .A1(n8457), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8444) );
  NAND2_X1 U10792 ( .A1(n6426), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8443) );
  NAND2_X1 U10793 ( .A1(n8440), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8442) );
  NAND2_X1 U10794 ( .A1(n8455), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8441) );
  XNOR2_X1 U10795 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8446) );
  XNOR2_X1 U10796 ( .A(n8447), .B(n8446), .ZN(n10042) );
  OR2_X1 U10797 ( .A1(n8448), .A2(n10042), .ZN(n8451) );
  OR2_X1 U10798 ( .A1(n8449), .A2(SI_2_), .ZN(n8450) );
  OAI211_X1 U10799 ( .C1(n9122), .C2(n9799), .A(n8451), .B(n8450), .ZN(n9804)
         );
  XNOR2_X1 U10800 ( .A(n15078), .B(n9804), .ZN(n9803) );
  INV_X1 U10801 ( .A(n9803), .ZN(n8993) );
  NAND2_X1 U10802 ( .A1(n15052), .A2(n8993), .ZN(n8452) );
  INV_X1 U10803 ( .A(n15078), .ZN(n10776) );
  INV_X1 U10804 ( .A(n9804), .ZN(n15053) );
  NAND2_X1 U10805 ( .A1(n10776), .A2(n15053), .ZN(n8868) );
  NAND2_X1 U10806 ( .A1(n8452), .A2(n8868), .ZN(n10836) );
  NAND2_X1 U10807 ( .A1(n6426), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8460) );
  NAND2_X1 U10808 ( .A1(n8455), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8459) );
  INV_X1 U10809 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n8456) );
  NAND2_X1 U10810 ( .A1(n8457), .A2(n8456), .ZN(n8458) );
  NAND3_X1 U10811 ( .A1(n8460), .A2(n8459), .A3(n8458), .ZN(n8461) );
  INV_X1 U10812 ( .A(n10780), .ZN(n12451) );
  OR2_X1 U10813 ( .A1(n8449), .A2(SI_3_), .ZN(n8468) );
  XNOR2_X1 U10814 ( .A(n10076), .B(P2_DATAO_REG_3__SCAN_IN), .ZN(n8462) );
  XNOR2_X1 U10815 ( .A(n8463), .B(n8462), .ZN(n10051) );
  OR2_X1 U10816 ( .A1(n8738), .A2(n10051), .ZN(n8467) );
  NAND2_X1 U10817 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n8464), .ZN(n8465) );
  XNOR2_X1 U10818 ( .A(n8465), .B(P3_IR_REG_3__SCAN_IN), .ZN(n14923) );
  OR2_X1 U10819 ( .A1(n9799), .A2(n14923), .ZN(n8466) );
  INV_X1 U10820 ( .A(n10845), .ZN(n10772) );
  NAND2_X1 U10821 ( .A1(n10780), .A2(n10845), .ZN(n8875) );
  INV_X1 U10822 ( .A(n9805), .ZN(n10838) );
  NAND2_X1 U10823 ( .A1(n10836), .A2(n10838), .ZN(n8469) );
  NAND2_X1 U10824 ( .A1(n8469), .A2(n8875), .ZN(n10827) );
  NAND2_X1 U10825 ( .A1(n6426), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8473) );
  OR2_X1 U10826 ( .A1(n7338), .A2(n8487), .ZN(n11004) );
  NAND2_X1 U10827 ( .A1(n8806), .A2(n11004), .ZN(n8472) );
  NAND2_X1 U10828 ( .A1(n8440), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8471) );
  NAND2_X1 U10829 ( .A1(n8455), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8470) );
  OR2_X1 U10830 ( .A1(n8829), .A2(SI_4_), .ZN(n8485) );
  NAND2_X1 U10831 ( .A1(n8475), .A2(n8474), .ZN(n8476) );
  AND2_X1 U10832 ( .A1(n8477), .A2(n8476), .ZN(n10055) );
  OR2_X1 U10833 ( .A1(n8738), .A2(n10055), .ZN(n8484) );
  NOR2_X1 U10834 ( .A1(n8478), .A2(n8479), .ZN(n8480) );
  MUX2_X1 U10835 ( .A(n8479), .B(n8480), .S(P3_IR_REG_4__SCAN_IN), .Z(n8482)
         );
  NAND2_X1 U10836 ( .A1(n8478), .A2(n14207), .ZN(n8511) );
  INV_X1 U10837 ( .A(n8511), .ZN(n8481) );
  NOR2_X2 U10838 ( .A1(n8482), .A2(n8481), .ZN(n9132) );
  OR2_X1 U10839 ( .A1(n9799), .A2(n9132), .ZN(n8483) );
  NAND2_X1 U10840 ( .A1(n11176), .A2(n11005), .ZN(n8880) );
  INV_X1 U10841 ( .A(n11005), .ZN(n11012) );
  NAND2_X1 U10842 ( .A1(n12450), .A2(n11012), .ZN(n8881) );
  NAND2_X1 U10843 ( .A1(n8880), .A2(n8881), .ZN(n9808) );
  NAND2_X1 U10844 ( .A1(n10827), .A2(n10828), .ZN(n8486) );
  NAND2_X1 U10845 ( .A1(n8486), .A2(n8880), .ZN(n11029) );
  OR2_X1 U10846 ( .A1(n8487), .A2(n10679), .ZN(n8488) );
  NAND2_X1 U10847 ( .A1(n8505), .A2(n8488), .ZN(n11180) );
  NAND2_X1 U10848 ( .A1(n8806), .A2(n11180), .ZN(n8492) );
  NAND2_X1 U10849 ( .A1(n6426), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8491) );
  NAND2_X1 U10850 ( .A1(n8440), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8490) );
  NAND2_X1 U10851 ( .A1(n8455), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8489) );
  OR2_X1 U10852 ( .A1(n8829), .A2(SI_5_), .ZN(n8502) );
  NAND2_X1 U10853 ( .A1(n8495), .A2(n8494), .ZN(n8497) );
  AND2_X1 U10854 ( .A1(n8497), .A2(n8496), .ZN(n10038) );
  OR2_X1 U10855 ( .A1(n8738), .A2(n10038), .ZN(n8501) );
  NAND2_X1 U10856 ( .A1(n8511), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8499) );
  INV_X1 U10857 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8498) );
  XNOR2_X1 U10858 ( .A(n8499), .B(n8498), .ZN(n10039) );
  OR2_X1 U10859 ( .A1(n9799), .A2(n7079), .ZN(n8500) );
  NAND2_X1 U10860 ( .A1(n11377), .A2(n11175), .ZN(n8888) );
  INV_X1 U10861 ( .A(n11175), .ZN(n11177) );
  NAND2_X1 U10862 ( .A1(n12449), .A2(n11177), .ZN(n8884) );
  NAND2_X1 U10863 ( .A1(n11029), .A2(n11030), .ZN(n8503) );
  NAND2_X1 U10864 ( .A1(n8503), .A2(n8888), .ZN(n11194) );
  NAND2_X1 U10865 ( .A1(n8505), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8506) );
  NAND2_X1 U10866 ( .A1(n8520), .A2(n8506), .ZN(n11529) );
  NAND2_X1 U10867 ( .A1(n8806), .A2(n11529), .ZN(n8510) );
  NAND2_X1 U10868 ( .A1(n6426), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8509) );
  INV_X1 U10869 ( .A(n8453), .ZN(n8536) );
  NAND2_X1 U10870 ( .A1(n8536), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8508) );
  NAND2_X1 U10871 ( .A1(n8455), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8507) );
  NOR2_X1 U10872 ( .A1(n8511), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n8514) );
  OR2_X1 U10873 ( .A1(n8514), .A2(n8479), .ZN(n8512) );
  MUX2_X1 U10874 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8512), .S(
        P3_IR_REG_6__SCAN_IN), .Z(n8515) );
  NAND2_X1 U10875 ( .A1(n8514), .A2(n8513), .ZN(n8541) );
  XNOR2_X1 U10876 ( .A(n8517), .B(n8516), .ZN(n10037) );
  OR2_X1 U10877 ( .A1(n8738), .A2(n10037), .ZN(n8519) );
  INV_X1 U10878 ( .A(SI_6_), .ZN(n10036) );
  OR2_X1 U10879 ( .A1(n8829), .A2(n10036), .ZN(n8518) );
  OAI211_X1 U10880 ( .C1(n9799), .C2(n10035), .A(n8519), .B(n8518), .ZN(n11521) );
  NAND2_X1 U10881 ( .A1(n11389), .A2(n11521), .ZN(n8890) );
  INV_X1 U10882 ( .A(n11521), .ZN(n11381) );
  NAND2_X1 U10883 ( .A1(n12448), .A2(n11381), .ZN(n8892) );
  NAND2_X1 U10884 ( .A1(n8890), .A2(n8892), .ZN(n11198) );
  INV_X1 U10885 ( .A(n11198), .ZN(n8989) );
  NAND2_X1 U10886 ( .A1(n6426), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8525) );
  AND2_X1 U10887 ( .A1(n8520), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8521) );
  OR2_X1 U10888 ( .A1(n8521), .A2(n8534), .ZN(n11374) );
  NAND2_X1 U10889 ( .A1(n8806), .A2(n11374), .ZN(n8524) );
  NAND2_X1 U10890 ( .A1(n8832), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8523) );
  NAND2_X1 U10891 ( .A1(n8455), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8522) );
  XNOR2_X1 U10892 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n8526) );
  XNOR2_X1 U10893 ( .A(n8527), .B(n8526), .ZN(n10045) );
  OR2_X1 U10894 ( .A1(n8738), .A2(n10045), .ZN(n8532) );
  OR2_X1 U10895 ( .A1(n8829), .A2(SI_7_), .ZN(n8531) );
  NAND2_X1 U10896 ( .A1(n8541), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8529) );
  INV_X1 U10897 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8528) );
  XNOR2_X1 U10898 ( .A(n8529), .B(n8528), .ZN(n10799) );
  OR2_X1 U10899 ( .A1(n9799), .A2(n9136), .ZN(n8530) );
  NAND2_X1 U10900 ( .A1(n11569), .A2(n9814), .ZN(n8895) );
  INV_X1 U10901 ( .A(n9814), .ZN(n15125) );
  NAND2_X1 U10902 ( .A1(n11562), .A2(n15125), .ZN(n8896) );
  NAND2_X1 U10903 ( .A1(n8895), .A2(n8896), .ZN(n11387) );
  INV_X1 U10904 ( .A(n11387), .ZN(n11247) );
  NAND2_X1 U10905 ( .A1(n6426), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8540) );
  NOR2_X1 U10906 ( .A1(n8534), .A2(n8533), .ZN(n8535) );
  OR2_X1 U10907 ( .A1(n8551), .A2(n8535), .ZN(n11560) );
  NAND2_X1 U10908 ( .A1(n8806), .A2(n11560), .ZN(n8539) );
  NAND2_X1 U10909 ( .A1(n8536), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8538) );
  NAND2_X1 U10910 ( .A1(n8455), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8537) );
  NAND2_X1 U10911 ( .A1(n8543), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8542) );
  MUX2_X1 U10912 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8542), .S(
        P3_IR_REG_8__SCAN_IN), .Z(n8544) );
  XNOR2_X1 U10913 ( .A(n8546), .B(n8545), .ZN(n10068) );
  OR2_X1 U10914 ( .A1(n10068), .A2(n8738), .ZN(n8548) );
  INV_X1 U10915 ( .A(SI_8_), .ZN(n10067) );
  OR2_X1 U10916 ( .A1(n8829), .A2(n10067), .ZN(n8547) );
  OAI211_X1 U10917 ( .C1(n9799), .C2(n10993), .A(n8548), .B(n8547), .ZN(n8549)
         );
  NAND2_X1 U10918 ( .A1(n11566), .A2(n8549), .ZN(n8899) );
  INV_X1 U10919 ( .A(n8549), .ZN(n15131) );
  NAND2_X1 U10920 ( .A1(n15040), .A2(n15131), .ZN(n8900) );
  NAND2_X1 U10921 ( .A1(n11316), .A2(n11317), .ZN(n8550) );
  NAND2_X1 U10922 ( .A1(n6426), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8556) );
  OR2_X1 U10923 ( .A1(n8551), .A2(n11740), .ZN(n8552) );
  NAND2_X1 U10924 ( .A1(n8571), .A2(n8552), .ZN(n15047) );
  NAND2_X1 U10925 ( .A1(n8806), .A2(n15047), .ZN(n8555) );
  NAND2_X1 U10926 ( .A1(n8832), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8554) );
  NAND2_X1 U10927 ( .A1(n8455), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8553) );
  NAND4_X1 U10928 ( .A1(n8556), .A2(n8555), .A3(n8554), .A4(n8553), .ZN(n11807) );
  XNOR2_X1 U10929 ( .A(n8558), .B(n8557), .ZN(n10070) );
  NAND2_X1 U10930 ( .A1(n10070), .A2(n8828), .ZN(n8561) );
  INV_X1 U10931 ( .A(SI_9_), .ZN(n10069) );
  NAND2_X1 U10932 ( .A1(n8566), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8559) );
  XNOR2_X1 U10933 ( .A(n8559), .B(P3_IR_REG_9__SCAN_IN), .ZN(n14959) );
  INV_X1 U10934 ( .A(n14959), .ZN(n10071) );
  AOI22_X1 U10935 ( .A1(n8699), .A2(n10069), .B1(n8438), .B2(n10071), .ZN(
        n8560) );
  NOR2_X1 U10936 ( .A1(n11807), .A2(n15046), .ZN(n8563) );
  NAND2_X1 U10937 ( .A1(n11807), .A2(n15046), .ZN(n8562) );
  XNOR2_X1 U10938 ( .A(n8565), .B(n8564), .ZN(n10073) );
  NAND2_X1 U10939 ( .A1(n10073), .A2(n8828), .ZN(n8570) );
  INV_X1 U10940 ( .A(SI_10_), .ZN(n10072) );
  OAI21_X1 U10941 ( .B1(n8566), .B2(P3_IR_REG_9__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8568) );
  INV_X1 U10942 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8567) );
  AOI22_X1 U10943 ( .A1(n8699), .A2(n10072), .B1(n8438), .B2(n14973), .ZN(
        n8569) );
  NAND2_X1 U10944 ( .A1(n8570), .A2(n8569), .ZN(n15033) );
  NAND2_X1 U10945 ( .A1(n8571), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8572) );
  NAND2_X1 U10946 ( .A1(n8597), .A2(n8572), .ZN(n15034) );
  NAND2_X1 U10947 ( .A1(n8806), .A2(n15034), .ZN(n8576) );
  NAND2_X1 U10948 ( .A1(n6426), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8575) );
  NAND2_X1 U10949 ( .A1(n8536), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8574) );
  NAND2_X1 U10950 ( .A1(n8455), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8573) );
  NAND4_X1 U10951 ( .A1(n8576), .A2(n8575), .A3(n8574), .A4(n8573), .ZN(n15039) );
  NAND2_X1 U10952 ( .A1(n15033), .A2(n15039), .ZN(n8903) );
  OR2_X1 U10953 ( .A1(n15039), .A2(n15033), .ZN(n8904) );
  XNOR2_X1 U10954 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8577) );
  XNOR2_X1 U10955 ( .A(n8578), .B(n8577), .ZN(n10089) );
  NAND2_X1 U10956 ( .A1(n10089), .A2(n8828), .ZN(n8581) );
  OR2_X1 U10957 ( .A1(n6439), .A2(n8479), .ZN(n8579) );
  XNOR2_X1 U10958 ( .A(n8579), .B(n8591), .ZN(n14989) );
  AOI22_X1 U10959 ( .A1(n8699), .A2(n10088), .B1(n8438), .B2(n14989), .ZN(
        n8580) );
  NAND2_X1 U10960 ( .A1(n8581), .A2(n8580), .ZN(n14457) );
  XNOR2_X1 U10961 ( .A(n8597), .B(P3_REG3_REG_11__SCAN_IN), .ZN(n14454) );
  NAND2_X1 U10962 ( .A1(n8806), .A2(n14454), .ZN(n8585) );
  NAND2_X1 U10963 ( .A1(n6426), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8584) );
  NAND2_X1 U10964 ( .A1(n8536), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8583) );
  NAND2_X1 U10965 ( .A1(n8455), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8582) );
  OR2_X1 U10966 ( .A1(n14457), .A2(n12447), .ZN(n8911) );
  NAND2_X1 U10967 ( .A1(n14457), .A2(n12447), .ZN(n8910) );
  NAND2_X1 U10968 ( .A1(n8586), .A2(n8911), .ZN(n11817) );
  INV_X1 U10969 ( .A(n8587), .ZN(n8588) );
  NAND2_X1 U10970 ( .A1(n6452), .A2(n8588), .ZN(n8589) );
  AND2_X1 U10971 ( .A1(n8590), .A2(n8589), .ZN(n10098) );
  NAND2_X1 U10972 ( .A1(n10098), .A2(n8828), .ZN(n8596) );
  NAND2_X1 U10973 ( .A1(n6439), .A2(n8591), .ZN(n8593) );
  NAND2_X1 U10974 ( .A1(n8593), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8592) );
  MUX2_X1 U10975 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8592), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n8594) );
  NAND2_X1 U10976 ( .A1(n8594), .A2(n8619), .ZN(n10100) );
  INV_X1 U10977 ( .A(n10100), .ZN(n12457) );
  AOI22_X1 U10978 ( .A1(n8699), .A2(SI_12_), .B1(n8438), .B2(n12457), .ZN(
        n8595) );
  NAND2_X1 U10979 ( .A1(n8596), .A2(n8595), .ZN(n11982) );
  NAND2_X1 U10980 ( .A1(n6426), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8602) );
  OAI21_X1 U10981 ( .B1(n8597), .B2(P3_REG3_REG_11__SCAN_IN), .A(
        P3_REG3_REG_12__SCAN_IN), .ZN(n8598) );
  NAND2_X1 U10982 ( .A1(n8598), .A2(n8610), .ZN(n11986) );
  NAND2_X1 U10983 ( .A1(n8806), .A2(n11986), .ZN(n8601) );
  NAND2_X1 U10984 ( .A1(n8832), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8600) );
  NAND2_X1 U10985 ( .A1(n8455), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8599) );
  OR2_X1 U10986 ( .A1(n11982), .A2(n12247), .ZN(n8918) );
  NAND2_X1 U10987 ( .A1(n11982), .A2(n12247), .ZN(n8917) );
  NAND2_X1 U10988 ( .A1(n11817), .A2(n11818), .ZN(n8603) );
  NAND2_X1 U10989 ( .A1(n8604), .A2(n10438), .ZN(n8605) );
  NAND2_X1 U10990 ( .A1(n8606), .A2(n8605), .ZN(n10258) );
  NAND2_X1 U10991 ( .A1(n10258), .A2(n8828), .ZN(n8609) );
  INV_X1 U10992 ( .A(SI_13_), .ZN(n10257) );
  NAND2_X1 U10993 ( .A1(n8619), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8607) );
  XNOR2_X1 U10994 ( .A(n8607), .B(P3_IR_REG_13__SCAN_IN), .ZN(n9148) );
  INV_X1 U10995 ( .A(n9148), .ZN(n15007) );
  AOI22_X1 U10996 ( .A1(n8699), .A2(n10257), .B1(n8438), .B2(n15007), .ZN(
        n8608) );
  NAND2_X1 U10997 ( .A1(n6426), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8615) );
  NAND2_X1 U10998 ( .A1(n8610), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8611) );
  NAND2_X1 U10999 ( .A1(n8623), .A2(n8611), .ZN(n12392) );
  NAND2_X1 U11000 ( .A1(n8806), .A2(n12392), .ZN(n8614) );
  NAND2_X1 U11001 ( .A1(n8536), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8613) );
  NAND2_X1 U11002 ( .A1(n8455), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8612) );
  NAND4_X1 U11003 ( .A1(n8615), .A2(n8614), .A3(n8613), .A4(n8612), .ZN(n12446) );
  OR2_X1 U11004 ( .A1(n12870), .A2(n12446), .ZN(n8922) );
  INV_X1 U11005 ( .A(n8922), .ZN(n8616) );
  NAND2_X1 U11006 ( .A1(n12870), .A2(n12446), .ZN(n8921) );
  XNOR2_X1 U11007 ( .A(n8618), .B(n8617), .ZN(n10322) );
  NAND2_X1 U11008 ( .A1(n10322), .A2(n8828), .ZN(n8622) );
  NOR2_X1 U11009 ( .A1(n8619), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n8635) );
  OR2_X1 U11010 ( .A1(n8635), .A2(n8479), .ZN(n8620) );
  XNOR2_X1 U11011 ( .A(n8620), .B(n8634), .ZN(n12474) );
  AOI22_X1 U11012 ( .A1(n8699), .A2(n10321), .B1(n8438), .B2(n12474), .ZN(
        n8621) );
  NAND2_X1 U11013 ( .A1(n6426), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8628) );
  NAND2_X1 U11014 ( .A1(n8623), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8624) );
  NAND2_X1 U11015 ( .A1(n8640), .A2(n8624), .ZN(n12298) );
  NAND2_X1 U11016 ( .A1(n8806), .A2(n12298), .ZN(n8627) );
  NAND2_X1 U11017 ( .A1(n8536), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8626) );
  NAND2_X1 U11018 ( .A1(n8455), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8625) );
  NAND4_X1 U11019 ( .A1(n8628), .A2(n8627), .A3(n8626), .A4(n8625), .ZN(n12445) );
  NAND2_X1 U11020 ( .A1(n12866), .A2(n12445), .ZN(n8925) );
  INV_X1 U11021 ( .A(n8925), .ZN(n8629) );
  OR2_X1 U11022 ( .A1(n12866), .A2(n12445), .ZN(n8926) );
  NAND2_X1 U11023 ( .A1(n8631), .A2(n8630), .ZN(n8632) );
  NAND2_X1 U11024 ( .A1(n8633), .A2(n8632), .ZN(n10442) );
  NAND2_X1 U11025 ( .A1(n10442), .A2(n8828), .ZN(n8639) );
  NAND2_X1 U11026 ( .A1(n8635), .A2(n8634), .ZN(n8650) );
  NAND2_X1 U11027 ( .A1(n8650), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8637) );
  XNOR2_X1 U11028 ( .A(n8637), .B(n8636), .ZN(n14437) );
  AOI22_X1 U11029 ( .A1(n8699), .A2(n10441), .B1(n8438), .B2(n14437), .ZN(
        n8638) );
  NAND2_X1 U11030 ( .A1(n6426), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8645) );
  NAND2_X1 U11031 ( .A1(n8640), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8641) );
  NAND2_X1 U11032 ( .A1(n8657), .A2(n8641), .ZN(n12742) );
  NAND2_X1 U11033 ( .A1(n8806), .A2(n12742), .ZN(n8644) );
  NAND2_X1 U11034 ( .A1(n8832), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8643) );
  NAND2_X1 U11035 ( .A1(n8455), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8642) );
  NAND2_X1 U11036 ( .A1(n12862), .A2(n12724), .ZN(n8929) );
  NAND2_X1 U11037 ( .A1(n12741), .A2(n12740), .ZN(n8646) );
  NAND2_X1 U11038 ( .A1(n8646), .A2(n8932), .ZN(n12727) );
  OAI21_X1 U11039 ( .B1(n8649), .B2(n8648), .A(n8647), .ZN(n10588) );
  OR2_X1 U11040 ( .A1(n10588), .A2(n8738), .ZN(n8656) );
  NAND2_X1 U11041 ( .A1(n8651), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8653) );
  INV_X1 U11042 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8652) );
  OR2_X1 U11043 ( .A1(n8653), .A2(n8652), .ZN(n8654) );
  NAND2_X1 U11044 ( .A1(n8653), .A2(n8652), .ZN(n8666) );
  AND2_X1 U11045 ( .A1(n8654), .A2(n8666), .ZN(n9154) );
  AOI22_X1 U11046 ( .A1(n8699), .A2(SI_16_), .B1(n8438), .B2(n9154), .ZN(n8655) );
  NAND2_X1 U11047 ( .A1(n6426), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8662) );
  NAND2_X1 U11048 ( .A1(n8657), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8658) );
  NAND2_X1 U11049 ( .A1(n8670), .A2(n8658), .ZN(n12730) );
  NAND2_X1 U11050 ( .A1(n8806), .A2(n12730), .ZN(n8661) );
  NAND2_X1 U11051 ( .A1(n8536), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8660) );
  NAND2_X1 U11052 ( .A1(n8455), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8659) );
  NAND4_X1 U11053 ( .A1(n8662), .A2(n8661), .A3(n8660), .A4(n8659), .ZN(n12710) );
  XNOR2_X1 U11054 ( .A(n12803), .B(n12710), .ZN(n12728) );
  NAND2_X1 U11055 ( .A1(n12727), .A2(n12728), .ZN(n8663) );
  NAND2_X1 U11056 ( .A1(n12803), .A2(n12738), .ZN(n8933) );
  NAND2_X1 U11057 ( .A1(n8663), .A2(n8933), .ZN(n12714) );
  XNOR2_X1 U11058 ( .A(n8665), .B(n8664), .ZN(n10724) );
  NAND2_X1 U11059 ( .A1(n10724), .A2(n8828), .ZN(n8669) );
  NAND2_X1 U11060 ( .A1(n8666), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8667) );
  XNOR2_X1 U11061 ( .A(n8667), .B(P3_IR_REG_17__SCAN_IN), .ZN(n12516) );
  INV_X1 U11062 ( .A(n12516), .ZN(n10722) );
  AOI22_X1 U11063 ( .A1(n8699), .A2(n10723), .B1(n8438), .B2(n10722), .ZN(
        n8668) );
  NAND2_X1 U11064 ( .A1(n6426), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8675) );
  NAND2_X1 U11065 ( .A1(n8670), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8671) );
  NAND2_X1 U11066 ( .A1(n8687), .A2(n8671), .ZN(n12716) );
  NAND2_X1 U11067 ( .A1(n8806), .A2(n12716), .ZN(n8674) );
  NAND2_X1 U11068 ( .A1(n8832), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8673) );
  NAND2_X1 U11069 ( .A1(n8455), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8672) );
  NAND4_X1 U11070 ( .A1(n8675), .A2(n8674), .A3(n8673), .A4(n8672), .ZN(n12725) );
  NAND2_X1 U11071 ( .A1(n12857), .A2(n12725), .ZN(n8853) );
  NAND2_X1 U11072 ( .A1(n8858), .A2(n8853), .ZN(n12708) );
  NAND2_X1 U11073 ( .A1(n12714), .A2(n9831), .ZN(n8676) );
  INV_X1 U11074 ( .A(n12697), .ZN(n8693) );
  INV_X1 U11075 ( .A(n8677), .ZN(n8680) );
  INV_X1 U11076 ( .A(n8678), .ZN(n8679) );
  NAND2_X1 U11077 ( .A1(n8680), .A2(n8679), .ZN(n8681) );
  AND2_X1 U11078 ( .A1(n8682), .A2(n8681), .ZN(n10941) );
  NAND2_X1 U11079 ( .A1(n10941), .A2(n8828), .ZN(n8686) );
  NAND2_X1 U11080 ( .A1(n8683), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8684) );
  XNOR2_X1 U11081 ( .A(n8684), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12536) );
  AOI22_X1 U11082 ( .A1(n8699), .A2(SI_18_), .B1(n8438), .B2(n12536), .ZN(
        n8685) );
  NAND2_X1 U11083 ( .A1(n8687), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8688) );
  NAND2_X1 U11084 ( .A1(n8702), .A2(n8688), .ZN(n12700) );
  NAND2_X1 U11085 ( .A1(n12700), .A2(n8806), .ZN(n8692) );
  NAND2_X1 U11086 ( .A1(n6426), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8691) );
  NAND2_X1 U11087 ( .A1(n8832), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8690) );
  NAND2_X1 U11088 ( .A1(n8455), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8689) );
  NAND4_X1 U11089 ( .A1(n8692), .A2(n8691), .A3(n8690), .A4(n8689), .ZN(n12711) );
  NAND2_X1 U11090 ( .A1(n12793), .A2(n12711), .ZN(n8855) );
  INV_X1 U11091 ( .A(n12793), .ZN(n9833) );
  INV_X1 U11092 ( .A(n12711), .ZN(n12407) );
  NAND2_X1 U11093 ( .A1(n9833), .A2(n12407), .ZN(n8941) );
  OAI21_X1 U11094 ( .B1(n8696), .B2(n8695), .A(n8694), .ZN(n10985) );
  OR2_X1 U11095 ( .A1(n10985), .A2(n8738), .ZN(n8701) );
  NAND2_X1 U11096 ( .A1(n6537), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8697) );
  MUX2_X1 U11097 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8697), .S(
        P3_IR_REG_19__SCAN_IN), .Z(n8698) );
  NAND2_X1 U11098 ( .A1(n8698), .A2(n8841), .ZN(n10984) );
  AOI22_X1 U11099 ( .A1(n8699), .A2(SI_19_), .B1(n9885), .B2(n8438), .ZN(n8700) );
  INV_X1 U11100 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n8706) );
  NAND2_X1 U11101 ( .A1(n8702), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8703) );
  NAND2_X1 U11102 ( .A1(n8713), .A2(n8703), .ZN(n12681) );
  NAND2_X1 U11103 ( .A1(n12681), .A2(n8806), .ZN(n8705) );
  AOI22_X1 U11104 ( .A1(n6426), .A2(P3_REG1_REG_19__SCAN_IN), .B1(n8832), .B2(
        P3_REG2_REG_19__SCAN_IN), .ZN(n8704) );
  OAI211_X1 U11105 ( .C1(n8707), .C2(n8706), .A(n8705), .B(n8704), .ZN(n12691)
         );
  INV_X1 U11106 ( .A(n12691), .ZN(n12411) );
  XNOR2_X1 U11107 ( .A(n12788), .B(n12411), .ZN(n12680) );
  INV_X1 U11108 ( .A(n12680), .ZN(n8708) );
  NAND2_X1 U11109 ( .A1(n12788), .A2(n12411), .ZN(n8946) );
  NAND2_X1 U11110 ( .A1(n12677), .A2(n8946), .ZN(n12667) );
  INV_X1 U11111 ( .A(n12667), .ZN(n8719) );
  XNOR2_X1 U11112 ( .A(n8710), .B(n8709), .ZN(n11208) );
  NAND2_X1 U11113 ( .A1(n11208), .A2(n8828), .ZN(n8712) );
  OR2_X1 U11114 ( .A1(n8829), .A2(n11210), .ZN(n8711) );
  NAND2_X1 U11115 ( .A1(n8713), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8714) );
  NAND2_X1 U11116 ( .A1(n8728), .A2(n8714), .ZN(n12669) );
  NAND2_X1 U11117 ( .A1(n12669), .A2(n8806), .ZN(n8717) );
  AOI22_X1 U11118 ( .A1(n8455), .A2(P3_REG0_REG_20__SCAN_IN), .B1(n8536), .B2(
        P3_REG2_REG_20__SCAN_IN), .ZN(n8716) );
  NAND2_X1 U11119 ( .A1(n6426), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n8715) );
  XNOR2_X1 U11120 ( .A(n12784), .B(n12653), .ZN(n12668) );
  OR2_X1 U11121 ( .A1(n12784), .A2(n12653), .ZN(n8951) );
  INV_X1 U11122 ( .A(n8720), .ZN(n8723) );
  INV_X1 U11123 ( .A(n8721), .ZN(n8722) );
  NAND2_X1 U11124 ( .A1(n8723), .A2(n8722), .ZN(n8724) );
  AND2_X1 U11125 ( .A1(n8725), .A2(n8724), .ZN(n11357) );
  NAND2_X1 U11126 ( .A1(n11357), .A2(n8828), .ZN(n8727) );
  INV_X1 U11127 ( .A(SI_21_), .ZN(n11359) );
  OR2_X1 U11128 ( .A1(n8829), .A2(n11359), .ZN(n8726) );
  NAND2_X1 U11129 ( .A1(n8728), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8729) );
  NAND2_X1 U11130 ( .A1(n8741), .A2(n8729), .ZN(n12657) );
  NAND2_X1 U11131 ( .A1(n12657), .A2(n8806), .ZN(n8734) );
  INV_X1 U11132 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12782) );
  NAND2_X1 U11133 ( .A1(n8536), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8731) );
  NAND2_X1 U11134 ( .A1(n8455), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8730) );
  OAI211_X1 U11135 ( .C1(n12782), .C2(n8835), .A(n8731), .B(n8730), .ZN(n8732)
         );
  INV_X1 U11136 ( .A(n8732), .ZN(n8733) );
  NAND2_X1 U11137 ( .A1(n12341), .A2(n12642), .ZN(n8954) );
  NAND2_X1 U11138 ( .A1(n12850), .A2(n12663), .ZN(n8955) );
  OAI21_X1 U11139 ( .B1(n8737), .B2(n8736), .A(n8735), .ZN(n11341) );
  OR2_X1 U11140 ( .A1(n11341), .A2(n8738), .ZN(n8740) );
  OR2_X1 U11141 ( .A1(n8829), .A2(n7848), .ZN(n8739) );
  NAND2_X1 U11142 ( .A1(n8741), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8742) );
  NAND2_X1 U11143 ( .A1(n8753), .A2(n8742), .ZN(n12646) );
  NAND2_X1 U11144 ( .A1(n12646), .A2(n8806), .ZN(n8747) );
  INV_X1 U11145 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12778) );
  NAND2_X1 U11146 ( .A1(n8832), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8744) );
  NAND2_X1 U11147 ( .A1(n8455), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8743) );
  OAI211_X1 U11148 ( .C1(n12778), .C2(n8835), .A(n8744), .B(n8743), .ZN(n8745)
         );
  INV_X1 U11149 ( .A(n8745), .ZN(n8746) );
  NAND2_X1 U11150 ( .A1(n8747), .A2(n8746), .ZN(n12629) );
  NAND2_X1 U11151 ( .A1(n12403), .A2(n12654), .ZN(n8851) );
  NAND2_X1 U11152 ( .A1(n12644), .A2(n8851), .ZN(n8748) );
  NAND2_X1 U11153 ( .A1(n12846), .A2(n12629), .ZN(n8852) );
  XNOR2_X1 U11154 ( .A(n8750), .B(n8749), .ZN(n11575) );
  NAND2_X1 U11155 ( .A1(n11575), .A2(n8828), .ZN(n8752) );
  OR2_X1 U11156 ( .A1(n8829), .A2(n11578), .ZN(n8751) );
  NAND2_X1 U11157 ( .A1(n8753), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8754) );
  NAND2_X1 U11158 ( .A1(n8764), .A2(n8754), .ZN(n12633) );
  NAND2_X1 U11159 ( .A1(n12633), .A2(n8806), .ZN(n8759) );
  INV_X1 U11160 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12774) );
  NAND2_X1 U11161 ( .A1(n8455), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8756) );
  NAND2_X1 U11162 ( .A1(n8440), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8755) );
  OAI211_X1 U11163 ( .C1(n8835), .C2(n12774), .A(n8756), .B(n8755), .ZN(n8757)
         );
  INV_X1 U11164 ( .A(n8757), .ZN(n8758) );
  NAND2_X1 U11165 ( .A1(n12771), .A2(n12643), .ZN(n8760) );
  NAND2_X1 U11166 ( .A1(n8963), .A2(n8760), .ZN(n9839) );
  XNOR2_X1 U11167 ( .A(n8761), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n11812) );
  NAND2_X1 U11168 ( .A1(n11812), .A2(n8828), .ZN(n8763) );
  INV_X1 U11169 ( .A(SI_24_), .ZN(n14087) );
  OR2_X1 U11170 ( .A1(n8829), .A2(n14087), .ZN(n8762) );
  NAND2_X1 U11171 ( .A1(n8764), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8765) );
  NAND2_X1 U11172 ( .A1(n8779), .A2(n8765), .ZN(n12618) );
  NAND2_X1 U11173 ( .A1(n12618), .A2(n8806), .ZN(n8770) );
  INV_X1 U11174 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12769) );
  NAND2_X1 U11175 ( .A1(n8455), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8767) );
  NAND2_X1 U11176 ( .A1(n8832), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8766) );
  OAI211_X1 U11177 ( .C1(n8835), .C2(n12769), .A(n8767), .B(n8766), .ZN(n8768)
         );
  INV_X1 U11178 ( .A(n8768), .ZN(n8769) );
  OR2_X1 U11179 ( .A1(n12377), .A2(n12595), .ZN(n8964) );
  NAND2_X1 U11180 ( .A1(n12377), .A2(n12595), .ZN(n8966) );
  NAND2_X1 U11181 ( .A1(n8964), .A2(n8966), .ZN(n12609) );
  INV_X1 U11182 ( .A(n8963), .ZN(n12610) );
  NOR2_X1 U11183 ( .A1(n12609), .A2(n12610), .ZN(n8771) );
  INV_X1 U11184 ( .A(n8772), .ZN(n8774) );
  NAND2_X1 U11185 ( .A1(n8774), .A2(n8773), .ZN(n8776) );
  AND2_X1 U11186 ( .A1(n8776), .A2(n8775), .ZN(n11906) );
  NAND2_X1 U11187 ( .A1(n11906), .A2(n8828), .ZN(n8778) );
  OR2_X1 U11188 ( .A1(n8829), .A2(n11907), .ZN(n8777) );
  NAND2_X1 U11189 ( .A1(n8779), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8780) );
  NAND2_X1 U11190 ( .A1(n8790), .A2(n8780), .ZN(n12603) );
  NAND2_X1 U11191 ( .A1(n12603), .A2(n8806), .ZN(n8785) );
  INV_X1 U11192 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12765) );
  NAND2_X1 U11193 ( .A1(n8455), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8782) );
  NAND2_X1 U11194 ( .A1(n8832), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8781) );
  OAI211_X1 U11195 ( .C1(n8835), .C2(n12765), .A(n8782), .B(n8781), .ZN(n8783)
         );
  INV_X1 U11196 ( .A(n8783), .ZN(n8784) );
  AND2_X1 U11197 ( .A1(n12602), .A2(n12614), .ZN(n8849) );
  XNOR2_X1 U11198 ( .A(n8787), .B(n8786), .ZN(n11952) );
  NAND2_X1 U11199 ( .A1(n11952), .A2(n8828), .ZN(n8789) );
  INV_X1 U11200 ( .A(SI_26_), .ZN(n11953) );
  OR2_X1 U11201 ( .A1(n8829), .A2(n11953), .ZN(n8788) );
  NAND2_X1 U11202 ( .A1(n8790), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8791) );
  NAND2_X1 U11203 ( .A1(n8804), .A2(n8791), .ZN(n12589) );
  NAND2_X1 U11204 ( .A1(n12589), .A2(n8806), .ZN(n8797) );
  INV_X1 U11205 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n8794) );
  NAND2_X1 U11206 ( .A1(n8832), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8793) );
  NAND2_X1 U11207 ( .A1(n8455), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8792) );
  OAI211_X1 U11208 ( .C1(n8835), .C2(n8794), .A(n8793), .B(n8792), .ZN(n8795)
         );
  INV_X1 U11209 ( .A(n8795), .ZN(n8796) );
  NAND2_X1 U11210 ( .A1(n12758), .A2(n12596), .ZN(n8844) );
  OR2_X1 U11211 ( .A1(n8799), .A2(n8798), .ZN(n8800) );
  AND2_X1 U11212 ( .A1(n8801), .A2(n8800), .ZN(n12878) );
  NAND2_X1 U11213 ( .A1(n12878), .A2(n8828), .ZN(n8803) );
  OR2_X1 U11214 ( .A1(n8829), .A2(n12881), .ZN(n8802) );
  NAND2_X1 U11215 ( .A1(n8804), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8805) );
  NAND2_X1 U11216 ( .A1(n8817), .A2(n8805), .ZN(n12575) );
  NAND2_X1 U11217 ( .A1(n12575), .A2(n8806), .ZN(n8811) );
  INV_X1 U11218 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12756) );
  NAND2_X1 U11219 ( .A1(n8455), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8808) );
  NAND2_X1 U11220 ( .A1(n8440), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8807) );
  OAI211_X1 U11221 ( .C1(n8835), .C2(n12756), .A(n8808), .B(n8807), .ZN(n8809)
         );
  INV_X1 U11222 ( .A(n8809), .ZN(n8810) );
  INV_X1 U11223 ( .A(n12568), .ZN(n8812) );
  NAND2_X1 U11224 ( .A1(n12563), .A2(n8812), .ZN(n9795) );
  XNOR2_X1 U11225 ( .A(n8814), .B(n8813), .ZN(n12026) );
  NAND2_X1 U11226 ( .A1(n12026), .A2(n8828), .ZN(n8816) );
  OR2_X1 U11227 ( .A1(n8829), .A2(n12027), .ZN(n8815) );
  NAND2_X1 U11228 ( .A1(n8817), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8818) );
  NAND2_X1 U11229 ( .A1(n12541), .A2(n8818), .ZN(n12556) );
  INV_X1 U11230 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n9893) );
  NAND2_X1 U11231 ( .A1(n8536), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8820) );
  NAND2_X1 U11232 ( .A1(n8455), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8819) );
  OAI211_X1 U11233 ( .C1(n8835), .C2(n9893), .A(n8820), .B(n8819), .ZN(n8821)
         );
  OR2_X1 U11234 ( .A1(n12330), .A2(n12442), .ZN(n8822) );
  INV_X1 U11235 ( .A(n8822), .ZN(n8825) );
  AND2_X1 U11236 ( .A1(n12289), .A2(n12422), .ZN(n9796) );
  NAND2_X1 U11237 ( .A1(n8822), .A2(n9796), .ZN(n8824) );
  NAND2_X1 U11238 ( .A1(n12330), .A2(n12442), .ZN(n8823) );
  OAI21_X2 U11239 ( .B1(n9795), .B2(n8825), .A(n8982), .ZN(n9906) );
  XNOR2_X1 U11240 ( .A(n13426), .B(P2_DATAO_REG_29__SCAN_IN), .ZN(n8826) );
  XNOR2_X1 U11241 ( .A(n8827), .B(n8826), .ZN(n12039) );
  NAND2_X1 U11242 ( .A1(n12039), .A2(n8828), .ZN(n8831) );
  OR2_X1 U11243 ( .A1(n8829), .A2(n12041), .ZN(n8830) );
  INV_X1 U11244 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9909) );
  NAND2_X1 U11245 ( .A1(n8832), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8834) );
  NAND2_X1 U11246 ( .A1(n8455), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8833) );
  OAI211_X1 U11247 ( .C1(n9909), .C2(n8835), .A(n8834), .B(n8833), .ZN(n8836)
         );
  INV_X1 U11248 ( .A(n8836), .ZN(n8837) );
  AND2_X1 U11249 ( .A1(n12543), .A2(n11269), .ZN(n8985) );
  NOR2_X1 U11250 ( .A1(n12540), .A2(n9901), .ZN(n8839) );
  NAND2_X1 U11251 ( .A1(n9910), .A2(n12327), .ZN(n8979) );
  OAI21_X1 U11252 ( .B1(n12753), .B2(n8839), .A(n8979), .ZN(n8840) );
  NAND2_X1 U11253 ( .A1(n6461), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8842) );
  NAND2_X1 U11254 ( .A1(n8841), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8843) );
  NAND2_X1 U11255 ( .A1(n10832), .A2(n9886), .ZN(n9845) );
  INV_X1 U11256 ( .A(n8844), .ZN(n8970) );
  NOR2_X1 U11257 ( .A1(n12602), .A2(n12614), .ZN(n8848) );
  NAND2_X1 U11258 ( .A1(n6500), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8845) );
  MUX2_X1 U11259 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8845), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n8847) );
  MUX2_X1 U11260 ( .A(n8849), .B(n8848), .S(n9887), .Z(n8850) );
  NOR2_X1 U11261 ( .A1(n12580), .A2(n8850), .ZN(n8974) );
  MUX2_X1 U11262 ( .A(n8851), .B(n8852), .S(n9887), .Z(n8959) );
  NOR2_X1 U11263 ( .A1(n12341), .A2(n12663), .ZN(n9836) );
  INV_X1 U11264 ( .A(n12788), .ZN(n12683) );
  NAND2_X1 U11265 ( .A1(n12683), .A2(n12691), .ZN(n8947) );
  INV_X1 U11266 ( .A(n8853), .ZN(n8854) );
  NAND2_X1 U11267 ( .A1(n8941), .A2(n8854), .ZN(n8856) );
  AND3_X1 U11268 ( .A1(n8856), .A2(n8855), .A3(n9887), .ZN(n8857) );
  NAND2_X1 U11269 ( .A1(n8947), .A2(n8857), .ZN(n8943) );
  INV_X1 U11270 ( .A(n8858), .ZN(n8940) );
  AND2_X1 U11271 ( .A1(n15077), .A2(n10582), .ZN(n8988) );
  INV_X1 U11272 ( .A(n8988), .ZN(n8859) );
  NAND2_X1 U11273 ( .A1(n8859), .A2(n11339), .ZN(n8862) );
  NAND2_X1 U11274 ( .A1(n8859), .A2(n10832), .ZN(n8860) );
  NAND3_X1 U11275 ( .A1(n10559), .A2(n9883), .A3(n8860), .ZN(n8861) );
  OAI21_X1 U11276 ( .B1(n9801), .B2(n8862), .A(n8861), .ZN(n8864) );
  NAND2_X1 U11277 ( .A1(n10566), .A2(n11360), .ZN(n8863) );
  NAND2_X1 U11278 ( .A1(n8864), .A2(n8863), .ZN(n8867) );
  MUX2_X1 U11279 ( .A(n8865), .B(n10559), .S(n9887), .Z(n8866) );
  NAND3_X1 U11280 ( .A1(n8867), .A2(n8993), .A3(n8866), .ZN(n8872) );
  NAND2_X1 U11281 ( .A1(n8875), .A2(n8868), .ZN(n8869) );
  NAND2_X1 U11282 ( .A1(n8869), .A2(n9883), .ZN(n8871) );
  INV_X1 U11283 ( .A(n8874), .ZN(n8870) );
  AOI21_X1 U11284 ( .B1(n8872), .B2(n8871), .A(n8870), .ZN(n8879) );
  NAND2_X1 U11285 ( .A1(n15078), .A2(n9804), .ZN(n8873) );
  AOI21_X1 U11286 ( .B1(n8874), .B2(n8873), .A(n9883), .ZN(n8878) );
  NOR2_X1 U11287 ( .A1(n8875), .A2(n9883), .ZN(n8876) );
  NOR2_X1 U11288 ( .A1(n8876), .A2(n9808), .ZN(n8877) );
  OAI21_X1 U11289 ( .B1(n8879), .B2(n8878), .A(n8877), .ZN(n8883) );
  MUX2_X1 U11290 ( .A(n8881), .B(n8880), .S(n9883), .Z(n8882) );
  NAND3_X1 U11291 ( .A1(n8883), .A2(n11030), .A3(n8882), .ZN(n8887) );
  NAND2_X1 U11292 ( .A1(n8892), .A2(n8884), .ZN(n8885) );
  NAND2_X1 U11293 ( .A1(n8885), .A2(n9883), .ZN(n8886) );
  NAND2_X1 U11294 ( .A1(n8887), .A2(n8886), .ZN(n8891) );
  AOI21_X1 U11295 ( .B1(n8890), .B2(n8888), .A(n9883), .ZN(n8889) );
  AOI21_X1 U11296 ( .B1(n8891), .B2(n8890), .A(n8889), .ZN(n8894) );
  NOR2_X1 U11297 ( .A1(n8892), .A2(n9883), .ZN(n8893) );
  OR3_X1 U11298 ( .A1(n8894), .A2(n8893), .A3(n11387), .ZN(n8898) );
  MUX2_X1 U11299 ( .A(n8896), .B(n8895), .S(n9887), .Z(n8897) );
  NAND3_X1 U11300 ( .A1(n8898), .A2(n11317), .A3(n8897), .ZN(n8902) );
  XNOR2_X1 U11301 ( .A(n8905), .B(n11807), .ZN(n15041) );
  NAND2_X1 U11302 ( .A1(n8904), .A2(n8903), .ZN(n9822) );
  MUX2_X1 U11303 ( .A(n8900), .B(n8899), .S(n9883), .Z(n8901) );
  NAND4_X1 U11304 ( .A1(n8902), .A2(n15041), .A3(n15026), .A4(n8901), .ZN(
        n8909) );
  MUX2_X1 U11305 ( .A(n8904), .B(n8903), .S(n9883), .Z(n8908) );
  NAND2_X1 U11306 ( .A1(n8905), .A2(n11807), .ZN(n9821) );
  MUX2_X1 U11307 ( .A(n11807), .B(n8905), .S(n9887), .Z(n8906) );
  NAND3_X1 U11308 ( .A1(n15026), .A2(n9821), .A3(n8906), .ZN(n8907) );
  NAND4_X1 U11309 ( .A1(n8909), .A2(n14455), .A3(n8908), .A4(n8907), .ZN(n8916) );
  NAND2_X1 U11310 ( .A1(n8918), .A2(n8910), .ZN(n8913) );
  NAND2_X1 U11311 ( .A1(n8917), .A2(n8911), .ZN(n8912) );
  MUX2_X1 U11312 ( .A(n8913), .B(n8912), .S(n9883), .Z(n8914) );
  INV_X1 U11313 ( .A(n8914), .ZN(n8915) );
  NAND2_X1 U11314 ( .A1(n8916), .A2(n8915), .ZN(n8920) );
  NAND2_X1 U11315 ( .A1(n8922), .A2(n8921), .ZN(n11868) );
  INV_X1 U11316 ( .A(n11868), .ZN(n11864) );
  MUX2_X1 U11317 ( .A(n8918), .B(n8917), .S(n9887), .Z(n8919) );
  NAND3_X1 U11318 ( .A1(n8920), .A2(n11864), .A3(n8919), .ZN(n8924) );
  NAND2_X1 U11319 ( .A1(n8926), .A2(n8925), .ZN(n11914) );
  INV_X1 U11320 ( .A(n11914), .ZN(n8998) );
  MUX2_X1 U11321 ( .A(n8922), .B(n8921), .S(n9887), .Z(n8923) );
  NAND3_X1 U11322 ( .A1(n8924), .A2(n8998), .A3(n8923), .ZN(n8928) );
  MUX2_X1 U11323 ( .A(n8926), .B(n8925), .S(n9883), .Z(n8927) );
  NAND2_X1 U11324 ( .A1(n8928), .A2(n8927), .ZN(n8931) );
  OAI21_X1 U11325 ( .B1(n12803), .B2(n12738), .A(n8929), .ZN(n8930) );
  AOI22_X1 U11326 ( .A1(n8931), .A2(n12740), .B1(n9883), .B2(n8930), .ZN(n8936) );
  INV_X1 U11327 ( .A(n8933), .ZN(n8935) );
  AND2_X1 U11328 ( .A1(n8933), .A2(n8932), .ZN(n8934) );
  OAI22_X1 U11329 ( .A1(n8936), .A2(n8935), .B1(n8934), .B2(n9883), .ZN(n8938)
         );
  INV_X1 U11330 ( .A(n12803), .ZN(n12732) );
  NAND3_X1 U11331 ( .A1(n12732), .A2(n9887), .A3(n12710), .ZN(n8937) );
  AOI21_X1 U11332 ( .B1(n8938), .B2(n8937), .A(n12708), .ZN(n8939) );
  AOI21_X1 U11333 ( .B1(n8943), .B2(n8940), .A(n8939), .ZN(n8945) );
  NAND3_X1 U11334 ( .A1(n8946), .A2(n9883), .A3(n8941), .ZN(n8942) );
  NAND2_X1 U11335 ( .A1(n8943), .A2(n8942), .ZN(n8944) );
  OAI21_X1 U11336 ( .B1(n8945), .B2(n12696), .A(n8944), .ZN(n8949) );
  MUX2_X1 U11337 ( .A(n8947), .B(n8946), .S(n9887), .Z(n8948) );
  NAND3_X1 U11338 ( .A1(n8949), .A2(n8718), .A3(n8948), .ZN(n8953) );
  NAND2_X1 U11339 ( .A1(n12784), .A2(n12653), .ZN(n8950) );
  MUX2_X1 U11340 ( .A(n8951), .B(n8950), .S(n9883), .Z(n8952) );
  NAND3_X1 U11341 ( .A1(n12655), .A2(n8953), .A3(n8952), .ZN(n8957) );
  MUX2_X1 U11342 ( .A(n8955), .B(n8954), .S(n9887), .Z(n8956) );
  NAND3_X1 U11343 ( .A1(n12645), .A2(n8957), .A3(n8956), .ZN(n8958) );
  NAND2_X1 U11344 ( .A1(n8959), .A2(n8958), .ZN(n8961) );
  NAND3_X1 U11345 ( .A1(n12771), .A2(n12643), .A3(n9887), .ZN(n8960) );
  OAI21_X1 U11346 ( .B1(n8961), .B2(n9839), .A(n8960), .ZN(n8962) );
  INV_X1 U11347 ( .A(n8962), .ZN(n8969) );
  NAND2_X1 U11348 ( .A1(n8964), .A2(n8963), .ZN(n8965) );
  NAND2_X1 U11349 ( .A1(n8965), .A2(n8966), .ZN(n8967) );
  MUX2_X1 U11350 ( .A(n8967), .B(n8966), .S(n9887), .Z(n8968) );
  OAI211_X1 U11351 ( .C1(n8969), .C2(n12609), .A(n12599), .B(n8968), .ZN(n8973) );
  MUX2_X1 U11352 ( .A(n8971), .B(n8970), .S(n9887), .Z(n8972) );
  AOI21_X1 U11353 ( .B1(n8974), .B2(n8973), .A(n8972), .ZN(n8976) );
  NAND2_X1 U11354 ( .A1(n8982), .A2(n9883), .ZN(n8975) );
  OR2_X1 U11355 ( .A1(n9797), .A2(n12568), .ZN(n9005) );
  MUX2_X1 U11356 ( .A(n8976), .B(n8975), .S(n9005), .Z(n8978) );
  INV_X1 U11357 ( .A(n9907), .ZN(n8977) );
  INV_X1 U11358 ( .A(n8980), .ZN(n8981) );
  INV_X1 U11359 ( .A(n9901), .ZN(n12441) );
  XNOR2_X1 U11360 ( .A(n12822), .B(n12441), .ZN(n9007) );
  INV_X1 U11361 ( .A(n8983), .ZN(n8984) );
  INV_X1 U11362 ( .A(n8985), .ZN(n9008) );
  NAND2_X1 U11363 ( .A1(n8986), .A2(n9008), .ZN(n9012) );
  NAND2_X1 U11364 ( .A1(n11211), .A2(n10984), .ZN(n9888) );
  INV_X1 U11365 ( .A(n9888), .ZN(n9791) );
  AND2_X1 U11366 ( .A1(n9885), .A2(n11211), .ZN(n15054) );
  INV_X1 U11367 ( .A(n15054), .ZN(n15086) );
  INV_X1 U11368 ( .A(n8987), .ZN(n9006) );
  INV_X1 U11369 ( .A(n12609), .ZN(n12607) );
  INV_X1 U11370 ( .A(n9801), .ZN(n8990) );
  NOR2_X1 U11371 ( .A1(n10566), .A2(n8988), .ZN(n10581) );
  NAND4_X1 U11372 ( .A1(n8990), .A2(n10581), .A3(n10838), .A4(n8989), .ZN(
        n8992) );
  NAND3_X1 U11373 ( .A1(n11247), .A2(n10828), .A3(n11030), .ZN(n8991) );
  NOR2_X1 U11374 ( .A1(n8992), .A2(n8991), .ZN(n8994) );
  AND4_X1 U11375 ( .A1(n8994), .A2(n8993), .A3(n11317), .A4(n15026), .ZN(n8995) );
  NAND4_X1 U11376 ( .A1(n11818), .A2(n15041), .A3(n14455), .A4(n8995), .ZN(
        n8996) );
  NOR2_X1 U11377 ( .A1(n11868), .A2(n8996), .ZN(n8997) );
  AND4_X1 U11378 ( .A1(n12728), .A2(n8998), .A3(n12740), .A4(n8997), .ZN(n8999) );
  NAND3_X1 U11379 ( .A1(n12687), .A2(n9831), .A3(n8999), .ZN(n9000) );
  NOR2_X1 U11380 ( .A1(n12680), .A2(n9000), .ZN(n9001) );
  NAND4_X1 U11381 ( .A1(n12645), .A2(n9001), .A3(n8718), .A4(n12655), .ZN(
        n9002) );
  NOR2_X1 U11382 ( .A1(n9839), .A2(n9002), .ZN(n9003) );
  NAND4_X1 U11383 ( .A1(n12581), .A2(n12607), .A3(n9003), .A4(n12599), .ZN(
        n9004) );
  NOR4_X1 U11384 ( .A1(n9006), .A2(n9005), .A3(n9907), .A4(n9004), .ZN(n9009)
         );
  NAND3_X1 U11385 ( .A1(n9009), .A2(n9008), .A3(n9007), .ZN(n9010) );
  XNOR2_X1 U11386 ( .A(n9010), .B(n10984), .ZN(n9011) );
  OR2_X1 U11387 ( .A1(n10832), .A2(n11211), .ZN(n10554) );
  NAND2_X1 U11388 ( .A1(n6480), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9015) );
  OR2_X1 U11389 ( .A1(n9061), .A2(P3_U3151), .ZN(n11576) );
  INV_X1 U11390 ( .A(n11576), .ZN(n9016) );
  NAND2_X1 U11391 ( .A1(n9023), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9024) );
  MUX2_X1 U11392 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9024), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n9025) );
  NAND2_X1 U11393 ( .A1(n9887), .A2(n9791), .ZN(n10499) );
  INV_X1 U11394 ( .A(n10499), .ZN(n9026) );
  INV_X1 U11395 ( .A(n12029), .ZN(n9117) );
  NAND3_X1 U11396 ( .A1(n10549), .A2(n9117), .A3(n12882), .ZN(n9027) );
  OAI211_X1 U11397 ( .C1(n11339), .C2(n11576), .A(n9027), .B(P3_B_REG_SCAN_IN), 
        .ZN(n9028) );
  NAND2_X1 U11398 ( .A1(n9029), .A2(n9028), .ZN(P3_U3296) );
  INV_X1 U11399 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14435) );
  INV_X1 U11400 ( .A(n14989), .ZN(n9143) );
  MUX2_X1 U11401 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n9037), .S(n9132), .Z(n10466) );
  INV_X1 U11402 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10820) );
  INV_X1 U11403 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15093) );
  INV_X1 U11404 ( .A(n10445), .ZN(n9033) );
  NAND2_X1 U11405 ( .A1(n10447), .A2(n9033), .ZN(n10446) );
  NAND2_X1 U11406 ( .A1(n9121), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9034) );
  INV_X1 U11407 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n14912) );
  INV_X1 U11408 ( .A(n10465), .ZN(n9038) );
  NOR2_X1 U11409 ( .A1(n7079), .A2(n9039), .ZN(n9041) );
  INV_X1 U11410 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10675) );
  XNOR2_X1 U11411 ( .A(n9040), .B(n10039), .ZN(n10674) );
  NOR2_X1 U11412 ( .A1(n10675), .A2(n10674), .ZN(n10673) );
  INV_X1 U11413 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n9042) );
  AOI22_X1 U11414 ( .A1(n14942), .A2(P3_REG2_REG_6__SCAN_IN), .B1(n9042), .B2(
        n10035), .ZN(n14928) );
  NOR2_X1 U11415 ( .A1(n9136), .A2(n9043), .ZN(n9044) );
  INV_X1 U11416 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11253) );
  NOR2_X1 U11417 ( .A1(n11253), .A2(n10789), .ZN(n10788) );
  INV_X1 U11418 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n9045) );
  AOI22_X1 U11419 ( .A1(n9139), .A2(P3_REG2_REG_8__SCAN_IN), .B1(n9045), .B2(
        n10993), .ZN(n10987) );
  NOR2_X1 U11420 ( .A1(n14959), .A2(n9046), .ZN(n9047) );
  INV_X1 U11421 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n15050) );
  INV_X1 U11422 ( .A(n14973), .ZN(n9142) );
  INV_X1 U11423 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n15036) );
  AOI22_X1 U11424 ( .A1(n9142), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n15036), 
        .B2(n14973), .ZN(n14970) );
  NOR2_X1 U11425 ( .A1(n14971), .A2(n14970), .ZN(n14969) );
  NAND2_X1 U11426 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n10100), .ZN(n9049) );
  OAI21_X1 U11427 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n10100), .A(n9049), .ZN(
        n12453) );
  NOR2_X1 U11428 ( .A1(n9148), .A2(n9050), .ZN(n9051) );
  INV_X1 U11429 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n15004) );
  XNOR2_X1 U11430 ( .A(n12474), .B(P3_REG2_REG_14__SCAN_IN), .ZN(n12471) );
  XNOR2_X1 U11431 ( .A(n9150), .B(n9053), .ZN(n14434) );
  NOR2_X1 U11432 ( .A1(n9150), .A2(n9053), .ZN(n9054) );
  INV_X1 U11433 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n9055) );
  AOI22_X1 U11434 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n9154), .B1(n12497), 
        .B2(n9055), .ZN(n12489) );
  INV_X1 U11435 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12507) );
  NOR2_X2 U11436 ( .A1(n12508), .A2(n12507), .ZN(n12506) );
  NOR2_X1 U11437 ( .A1(n12516), .A2(n9056), .ZN(n9057) );
  INV_X1 U11438 ( .A(n12536), .ZN(n10942) );
  NAND2_X1 U11439 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n10942), .ZN(n9058) );
  OAI21_X1 U11440 ( .B1(P3_REG2_REG_18__SCAN_IN), .B2(n10942), .A(n9058), .ZN(
        n12524) );
  XNOR2_X1 U11441 ( .A(n10984), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n9063) );
  XNOR2_X1 U11442 ( .A(n9059), .B(n9063), .ZN(n9162) );
  INV_X1 U11443 ( .A(n10573), .ZN(n9060) );
  NAND2_X1 U11444 ( .A1(n9060), .A2(n11576), .ZN(n9114) );
  NAND2_X1 U11445 ( .A1(n9887), .A2(n9061), .ZN(n9062) );
  AND2_X1 U11446 ( .A1(n9062), .A2(n9799), .ZN(n9112) );
  NAND2_X1 U11447 ( .A1(n9114), .A2(n9112), .ZN(n9159) );
  INV_X1 U11448 ( .A(n12882), .ZN(n9158) );
  NAND2_X1 U11449 ( .A1(n9117), .A2(n9158), .ZN(n9800) );
  OR2_X1 U11450 ( .A1(n9159), .A2(n9800), .ZN(n15023) );
  MUX2_X1 U11451 ( .A(n9063), .B(n6575), .S(n12882), .Z(n9111) );
  INV_X1 U11452 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n9064) );
  INV_X1 U11453 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n14200) );
  MUX2_X1 U11454 ( .A(n9064), .B(n14200), .S(n12882), .Z(n12527) );
  INV_X1 U11455 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12801) );
  MUX2_X1 U11456 ( .A(n12507), .B(n12801), .S(n12882), .Z(n9106) );
  NOR2_X1 U11457 ( .A1(n9106), .A2(n12516), .ZN(n9108) );
  MUX2_X1 U11458 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n12882), .Z(n9065) );
  AND2_X1 U11459 ( .A1(n9065), .A2(n12497), .ZN(n12490) );
  MUX2_X1 U11460 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n12882), .Z(n9101) );
  INV_X1 U11461 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n15011) );
  MUX2_X1 U11462 ( .A(n15004), .B(n15011), .S(n12882), .Z(n9098) );
  XNOR2_X1 U11463 ( .A(n9098), .B(n9148), .ZN(n15014) );
  MUX2_X1 U11464 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12882), .Z(n9066) );
  NAND2_X1 U11465 ( .A1(n9066), .A2(n10100), .ZN(n9097) );
  XNOR2_X1 U11466 ( .A(n9066), .B(n10100), .ZN(n12456) );
  INV_X1 U11467 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n9068) );
  INV_X1 U11468 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n9067) );
  MUX2_X1 U11469 ( .A(n9068), .B(n9067), .S(n12882), .Z(n9093) );
  NAND2_X1 U11470 ( .A1(n9093), .A2(n9143), .ZN(n9095) );
  MUX2_X1 U11471 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n12882), .Z(n9090) );
  NOR2_X1 U11472 ( .A1(n9090), .A2(n14973), .ZN(n9092) );
  MUX2_X1 U11473 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n12882), .Z(n9088) );
  NOR2_X1 U11474 ( .A1(n9088), .A2(n10071), .ZN(n9089) );
  MUX2_X1 U11475 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12882), .Z(n9087) );
  MUX2_X1 U11476 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12882), .Z(n9074) );
  XNOR2_X1 U11477 ( .A(n9074), .B(n9132), .ZN(n10464) );
  MUX2_X1 U11478 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n12882), .Z(n9069) );
  OR2_X1 U11479 ( .A1(n9069), .A2(n10054), .ZN(n9073) );
  XNOR2_X1 U11480 ( .A(n9069), .B(n14923), .ZN(n14921) );
  MUX2_X1 U11481 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n6430), .Z(n9070) );
  MUX2_X1 U11482 ( .A(n10820), .B(n10503), .S(n6430), .Z(n14904) );
  AND2_X1 U11483 ( .A1(n14904), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n14907) );
  INV_X1 U11484 ( .A(n9070), .ZN(n9071) );
  MUX2_X1 U11485 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n6431), .Z(n9072) );
  XOR2_X1 U11486 ( .A(n9122), .B(n9072), .Z(n10455) );
  OAI22_X1 U11487 ( .A1(n10456), .A2(n10455), .B1(n9072), .B2(n9121), .ZN(
        n14922) );
  NAND2_X1 U11488 ( .A1(n14921), .A2(n14922), .ZN(n14920) );
  NAND2_X1 U11489 ( .A1(n9073), .A2(n14920), .ZN(n10463) );
  MUX2_X1 U11490 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12882), .Z(n9075) );
  NAND2_X1 U11491 ( .A1(n9075), .A2(n10039), .ZN(n10676) );
  NAND2_X1 U11492 ( .A1(n10678), .A2(n10676), .ZN(n14933) );
  INV_X1 U11493 ( .A(n9075), .ZN(n9076) );
  NAND2_X1 U11494 ( .A1(n9076), .A2(n7079), .ZN(n14932) );
  INV_X1 U11495 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n9077) );
  MUX2_X1 U11496 ( .A(n9042), .B(n9077), .S(n12882), .Z(n9078) );
  NAND2_X1 U11497 ( .A1(n9078), .A2(n14942), .ZN(n9081) );
  INV_X1 U11498 ( .A(n9078), .ZN(n9079) );
  NAND2_X1 U11499 ( .A1(n9079), .A2(n10035), .ZN(n9080) );
  NAND2_X1 U11500 ( .A1(n9081), .A2(n9080), .ZN(n14931) );
  INV_X1 U11501 ( .A(n9081), .ZN(n10794) );
  INV_X1 U11502 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n9082) );
  MUX2_X1 U11503 ( .A(n11253), .B(n9082), .S(n12882), .Z(n9083) );
  NAND2_X1 U11504 ( .A1(n9083), .A2(n9136), .ZN(n9086) );
  INV_X1 U11505 ( .A(n9083), .ZN(n9084) );
  NAND2_X1 U11506 ( .A1(n9084), .A2(n10799), .ZN(n9085) );
  AND2_X1 U11507 ( .A1(n9086), .A2(n9085), .ZN(n10793) );
  NAND2_X1 U11508 ( .A1(n10796), .A2(n9086), .ZN(n10991) );
  XNOR2_X1 U11509 ( .A(n9087), .B(n9139), .ZN(n10990) );
  NAND2_X1 U11510 ( .A1(n10991), .A2(n10990), .ZN(n10989) );
  OAI21_X1 U11511 ( .B1(n9087), .B2(n10993), .A(n10989), .ZN(n14962) );
  AOI21_X1 U11512 ( .B1(n9088), .B2(n10071), .A(n9089), .ZN(n14961) );
  AND2_X1 U11513 ( .A1(n14962), .A2(n14961), .ZN(n14965) );
  NOR2_X1 U11514 ( .A1(n9089), .A2(n14965), .ZN(n14977) );
  AOI21_X1 U11515 ( .B1(n9090), .B2(n14973), .A(n9092), .ZN(n9091) );
  INV_X1 U11516 ( .A(n9091), .ZN(n14978) );
  OAI21_X1 U11517 ( .B1(n9093), .B2(n9143), .A(n9095), .ZN(n14994) );
  NOR2_X1 U11518 ( .A1(n14993), .A2(n14994), .ZN(n14992) );
  INV_X1 U11519 ( .A(n14992), .ZN(n9094) );
  AOI21_X1 U11520 ( .B1(n9098), .B2(n9148), .A(n15012), .ZN(n12478) );
  INV_X1 U11521 ( .A(n12471), .ZN(n9100) );
  XNOR2_X1 U11522 ( .A(n12474), .B(P3_REG1_REG_14__SCAN_IN), .ZN(n12470) );
  INV_X1 U11523 ( .A(n12470), .ZN(n9099) );
  MUX2_X1 U11524 ( .A(n9100), .B(n9099), .S(n12882), .Z(n12477) );
  AOI21_X1 U11525 ( .B1(n12474), .B2(n9101), .A(n12475), .ZN(n9103) );
  INV_X1 U11526 ( .A(n9104), .ZN(n9102) );
  MUX2_X1 U11527 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12882), .Z(n14443) );
  NOR2_X1 U11528 ( .A1(n9104), .A2(n14441), .ZN(n12494) );
  INV_X1 U11529 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n9153) );
  MUX2_X1 U11530 ( .A(n9055), .B(n9153), .S(n12882), .Z(n9105) );
  NAND2_X1 U11531 ( .A1(n9105), .A2(n9154), .ZN(n12492) );
  OAI21_X1 U11532 ( .B1(n12490), .B2(n12494), .A(n12492), .ZN(n12513) );
  AOI21_X1 U11533 ( .B1(n12516), .B2(n9106), .A(n9108), .ZN(n9107) );
  INV_X1 U11534 ( .A(n9107), .ZN(n12512) );
  XNOR2_X1 U11535 ( .A(n10942), .B(n9109), .ZN(n12528) );
  NAND2_X1 U11536 ( .A1(n12527), .A2(n12528), .ZN(n12526) );
  NAND2_X1 U11537 ( .A1(n12536), .A2(n9109), .ZN(n9110) );
  INV_X1 U11538 ( .A(n9112), .ZN(n9113) );
  NAND2_X1 U11539 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12314)
         );
  OAI21_X1 U11540 ( .B1(n15005), .B2(n7365), .A(n12314), .ZN(n9115) );
  INV_X1 U11541 ( .A(n9159), .ZN(n9118) );
  MUX2_X1 U11542 ( .A(n9118), .B(P3_U3897), .S(n9117), .Z(n14960) );
  NAND2_X1 U11543 ( .A1(n14960), .A2(n9885), .ZN(n9119) );
  NAND2_X1 U11544 ( .A1(n9121), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n9129) );
  INV_X1 U11545 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n15149) );
  NAND2_X1 U11546 ( .A1(n9122), .A2(n15149), .ZN(n9123) );
  NAND2_X1 U11547 ( .A1(n9129), .A2(n9123), .ZN(n10448) );
  INV_X1 U11548 ( .A(n10448), .ZN(n9128) );
  INV_X1 U11549 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n15147) );
  NOR2_X1 U11550 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n10503), .ZN(n9125) );
  INV_X1 U11551 ( .A(n9126), .ZN(n9124) );
  OAI21_X1 U11552 ( .B1(n10066), .B2(n9125), .A(n9124), .ZN(n10507) );
  NAND2_X1 U11553 ( .A1(n10451), .A2(n9129), .ZN(n9130) );
  OR2_X1 U11554 ( .A1(n9130), .A2(n10054), .ZN(n9131) );
  INV_X1 U11555 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15151) );
  INV_X1 U11556 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15153) );
  MUX2_X1 U11557 ( .A(n15153), .B(P3_REG1_REG_4__SCAN_IN), .S(n9132), .Z(
        n10470) );
  NOR2_X1 U11558 ( .A1(n7079), .A2(n9133), .ZN(n9134) );
  INV_X1 U11559 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15155) );
  AOI22_X1 U11560 ( .A1(n14942), .A2(P3_REG1_REG_6__SCAN_IN), .B1(n9077), .B2(
        n10035), .ZN(n14937) );
  NOR2_X1 U11561 ( .A1(n14938), .A2(n14937), .ZN(n14936) );
  NOR2_X1 U11562 ( .A1(n9136), .A2(n9137), .ZN(n9138) );
  XNOR2_X1 U11563 ( .A(n9137), .B(n9136), .ZN(n10791) );
  NOR2_X1 U11564 ( .A1(n9082), .A2(n10791), .ZN(n10790) );
  INV_X1 U11565 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15159) );
  AOI22_X1 U11566 ( .A1(n9139), .A2(P3_REG1_REG_8__SCAN_IN), .B1(n15159), .B2(
        n10993), .ZN(n10995) );
  NOR2_X1 U11567 ( .A1(n14959), .A2(n9140), .ZN(n9141) );
  INV_X1 U11568 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15161) );
  INV_X1 U11569 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n15164) );
  AOI22_X1 U11570 ( .A1(n9142), .A2(P3_REG1_REG_10__SCAN_IN), .B1(n15164), 
        .B2(n14973), .ZN(n14975) );
  AOI21_X2 U11571 ( .B1(P3_REG1_REG_10__SCAN_IN), .B2(n14973), .A(n14974), 
        .ZN(n9144) );
  NOR2_X1 U11572 ( .A1(n9143), .A2(n9144), .ZN(n9145) );
  NAND2_X1 U11573 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n10100), .ZN(n9146) );
  OAI21_X1 U11574 ( .B1(P3_REG1_REG_12__SCAN_IN), .B2(n10100), .A(n9146), .ZN(
        n12463) );
  NOR2_X1 U11575 ( .A1(n9148), .A2(n9147), .ZN(n9149) );
  NOR2_X1 U11576 ( .A1(n9150), .A2(n9151), .ZN(n9152) );
  INV_X1 U11577 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n14440) );
  AOI22_X1 U11578 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n9154), .B1(n12497), 
        .B2(n9153), .ZN(n12499) );
  NOR2_X1 U11579 ( .A1(n12518), .A2(n12801), .ZN(n12517) );
  NOR2_X1 U11580 ( .A1(n12516), .A2(n9155), .ZN(n9156) );
  AOI22_X1 U11581 ( .A1(P3_REG1_REG_18__SCAN_IN), .A2(n12536), .B1(n10942), 
        .B2(n14200), .ZN(n12533) );
  AOI21_X1 U11582 ( .B1(P3_REG1_REG_18__SCAN_IN), .B2(n10942), .A(n12532), 
        .ZN(n9157) );
  OAI211_X1 U11583 ( .C1(n9162), .C2(n15023), .A(n7339), .B(n9161), .ZN(
        P3_U3201) );
  NOR2_X1 U11584 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n9167) );
  NAND4_X1 U11585 ( .A1(n9167), .A2(n9166), .A3(n9165), .A4(n9284), .ZN(n9168)
         );
  NOR2_X1 U11586 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), 
        .ZN(n9174) );
  NOR2_X1 U11587 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n9173) );
  AND2_X1 U11588 ( .A1(n9174), .A2(n9173), .ZN(n9175) );
  AND4_X2 U11589 ( .A1(n9199), .A2(n9200), .A3(n9176), .A4(n9175), .ZN(n9177)
         );
  INV_X2 U11590 ( .A(n12031), .ZN(n9182) );
  INV_X1 U11591 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10602) );
  INV_X1 U11592 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9183) );
  OR2_X1 U11593 ( .A1(n9675), .A2(n9183), .ZN(n9188) );
  INV_X1 U11594 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9185) );
  AND2_X4 U11595 ( .A1(n14270), .A2(n12031), .ZN(n9621) );
  NAND2_X1 U11596 ( .A1(n9621), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9186) );
  NOR2_X1 U11597 ( .A1(n10049), .A2(n9190), .ZN(n9192) );
  XNOR2_X1 U11598 ( .A(n9192), .B(n9191), .ZN(n14285) );
  XNOR2_X2 U11599 ( .A(n9196), .B(n9195), .ZN(n9784) );
  MUX2_X1 U11600 ( .A(n14284), .B(n14285), .S(n9558), .Z(n11125) );
  NAND2_X1 U11601 ( .A1(n9202), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9203) );
  NAND2_X1 U11602 ( .A1(n9209), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9205) );
  NAND2_X1 U11603 ( .A1(n9207), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9208) );
  MUX2_X1 U11604 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9208), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n9210) );
  NAND2_X1 U11605 ( .A1(n9211), .A2(n10315), .ZN(n9212) );
  NAND2_X1 U11606 ( .A1(n9212), .A2(n11650), .ZN(n9701) );
  NAND2_X1 U11607 ( .A1(n11085), .A2(n11257), .ZN(n10317) );
  NAND2_X1 U11608 ( .A1(n9701), .A2(n10317), .ZN(n9704) );
  NAND2_X1 U11609 ( .A1(n9212), .A2(n11257), .ZN(n9213) );
  INV_X1 U11610 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10324) );
  INV_X1 U11611 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n11139) );
  OR2_X1 U11612 ( .A1(n9695), .A2(n14202), .ZN(n9215) );
  NAND2_X1 U11613 ( .A1(n9621), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n9214) );
  INV_X1 U11614 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n9219) );
  NAND2_X1 U11615 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n14284), .ZN(n9218) );
  OR2_X1 U11616 ( .A1(n9247), .A2(n7367), .ZN(n9221) );
  OAI211_X2 U11617 ( .C1(n9558), .C2(n13577), .A(n9221), .B(n9220), .ZN(n11141) );
  OAI211_X1 U11618 ( .C1(n11258), .C2(n10591), .A(n9222), .B(n11131), .ZN(
        n9228) );
  AND2_X1 U11619 ( .A1(n9310), .A2(n10630), .ZN(n9225) );
  NAND3_X1 U11620 ( .A1(n9228), .A2(n9227), .A3(n9226), .ZN(n9257) );
  NAND2_X1 U11621 ( .A1(n9621), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9233) );
  INV_X1 U11622 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9229) );
  INV_X1 U11623 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10323) );
  OR2_X1 U11624 ( .A1(n6424), .A2(n10323), .ZN(n9231) );
  INV_X1 U11625 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10339) );
  OR2_X1 U11626 ( .A1(n9695), .A2(n10339), .ZN(n9230) );
  NAND2_X1 U11627 ( .A1(n9310), .A2(n11073), .ZN(n9240) );
  OR2_X1 U11628 ( .A1(n10082), .A2(n9253), .ZN(n9239) );
  OR2_X1 U11629 ( .A1(n9716), .A2(n10060), .ZN(n9238) );
  OR2_X1 U11630 ( .A1(n9234), .A2(n9445), .ZN(n9236) );
  XNOR2_X1 U11631 ( .A(n9236), .B(n9235), .ZN(n13598) );
  OR2_X1 U11632 ( .A1(n9558), .A2(n13598), .ZN(n9237) );
  NAND2_X1 U11633 ( .A1(n11073), .A2(n14661), .ZN(n11064) );
  INV_X2 U11634 ( .A(n9310), .ZN(n9724) );
  MUX2_X1 U11635 ( .A(n11073), .B(n14661), .S(n9310), .Z(n9241) );
  OAI21_X1 U11636 ( .B1(n9257), .B2(n9242), .A(n9241), .ZN(n9259) );
  INV_X1 U11637 ( .A(n14661), .ZN(n14638) );
  NAND2_X1 U11638 ( .A1(n9621), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9246) );
  INV_X1 U11639 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10328) );
  OR2_X1 U11640 ( .A1(n9675), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9244) );
  INV_X1 U11641 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10338) );
  OR2_X1 U11642 ( .A1(n9695), .A2(n10338), .ZN(n9243) );
  INV_X2 U11643 ( .A(n9247), .ZN(n9506) );
  NAND2_X1 U11644 ( .A1(n9249), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9250) );
  MUX2_X1 U11645 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9250), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n9252) );
  AND2_X1 U11646 ( .A1(n9252), .A2(n9251), .ZN(n13607) );
  OR2_X1 U11647 ( .A1(n10077), .A2(n9253), .ZN(n9254) );
  XNOR2_X2 U11648 ( .A(n13571), .B(n14668), .ZN(n11186) );
  INV_X1 U11649 ( .A(n11186), .ZN(n11066) );
  NAND2_X1 U11650 ( .A1(n9259), .A2(n9258), .ZN(n9262) );
  INV_X1 U11651 ( .A(n14668), .ZN(n11190) );
  NAND2_X1 U11652 ( .A1(n13571), .A2(n11190), .ZN(n9260) );
  INV_X1 U11653 ( .A(n13571), .ZN(n11067) );
  NAND2_X1 U11654 ( .A1(n11067), .A2(n14668), .ZN(n11075) );
  INV_X4 U11655 ( .A(n9724), .ZN(n9707) );
  MUX2_X1 U11656 ( .A(n9260), .B(n11075), .S(n9707), .Z(n9261) );
  NAND2_X1 U11657 ( .A1(n10062), .A2(n9715), .ZN(n9265) );
  NAND2_X1 U11658 ( .A1(n9251), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9263) );
  XNOR2_X1 U11659 ( .A(n9263), .B(P1_IR_REG_4__SCAN_IN), .ZN(n14579) );
  AOI22_X1 U11660 ( .A1(n9506), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n10162), 
        .B2(n14579), .ZN(n9264) );
  NAND2_X1 U11661 ( .A1(n9621), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9272) );
  INV_X1 U11662 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10344) );
  OR2_X1 U11663 ( .A1(n9695), .A2(n10344), .ZN(n9271) );
  INV_X1 U11664 ( .A(n9279), .ZN(n9268) );
  INV_X1 U11665 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9266) );
  INV_X1 U11666 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n10949) );
  NAND2_X1 U11667 ( .A1(n9266), .A2(n10949), .ZN(n9267) );
  NAND2_X1 U11668 ( .A1(n9268), .A2(n9267), .ZN(n11272) );
  OR2_X1 U11669 ( .A1(n9675), .A2(n11272), .ZN(n9270) );
  OR2_X1 U11670 ( .A1(n6424), .A2(n14735), .ZN(n9269) );
  INV_X4 U11671 ( .A(n9724), .ZN(n9289) );
  MUX2_X1 U11672 ( .A(n14680), .B(n11077), .S(n9289), .Z(n9274) );
  INV_X1 U11673 ( .A(n11077), .ZN(n13570) );
  MUX2_X1 U11674 ( .A(n13570), .B(n11274), .S(n9707), .Z(n9273) );
  OAI21_X1 U11675 ( .B1(n9275), .B2(n9274), .A(n9273), .ZN(n9277) );
  NAND2_X1 U11676 ( .A1(n9275), .A2(n9274), .ZN(n9276) );
  NAND2_X1 U11677 ( .A1(n9277), .A2(n9276), .ZN(n9292) );
  NAND2_X1 U11678 ( .A1(n9672), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9283) );
  INV_X1 U11679 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9278) );
  OR2_X1 U11680 ( .A1(n9697), .A2(n9278), .ZN(n9282) );
  NAND2_X1 U11681 ( .A1(n9279), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9315) );
  OAI21_X1 U11682 ( .B1(n9279), .B2(P1_REG3_REG_5__SCAN_IN), .A(n9315), .ZN(
        n11090) );
  OR2_X1 U11683 ( .A1(n9675), .A2(n11090), .ZN(n9281) );
  OR2_X1 U11684 ( .A1(n6425), .A2(n6612), .ZN(n9280) );
  NAND4_X1 U11685 ( .A1(n9283), .A2(n9282), .A3(n9281), .A4(n9280), .ZN(n13569) );
  OR2_X1 U11686 ( .A1(n10080), .A2(n9253), .ZN(n9288) );
  INV_X1 U11687 ( .A(n9251), .ZN(n9285) );
  NAND2_X1 U11688 ( .A1(n9285), .A2(n9284), .ZN(n9298) );
  NAND2_X1 U11689 ( .A1(n9298), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9286) );
  XNOR2_X1 U11690 ( .A(n9286), .B(P1_IR_REG_5__SCAN_IN), .ZN(n13621) );
  AOI22_X1 U11691 ( .A1(n9506), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n10162), 
        .B2(n13621), .ZN(n9287) );
  NAND2_X1 U11692 ( .A1(n9288), .A2(n9287), .ZN(n11293) );
  MUX2_X1 U11693 ( .A(n13569), .B(n11293), .S(n9289), .Z(n9293) );
  NAND2_X1 U11694 ( .A1(n9292), .A2(n9293), .ZN(n9291) );
  MUX2_X1 U11695 ( .A(n11293), .B(n13569), .S(n9707), .Z(n9290) );
  NAND2_X1 U11696 ( .A1(n9291), .A2(n9290), .ZN(n9297) );
  INV_X1 U11697 ( .A(n9292), .ZN(n9295) );
  INV_X1 U11698 ( .A(n9293), .ZN(n9294) );
  NAND2_X1 U11699 ( .A1(n9295), .A2(n9294), .ZN(n9296) );
  OR2_X1 U11700 ( .A1(n10075), .A2(n9253), .ZN(n9303) );
  INV_X1 U11701 ( .A(n9298), .ZN(n9300) );
  INV_X1 U11702 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9299) );
  NAND2_X1 U11703 ( .A1(n9300), .A2(n9299), .ZN(n9321) );
  NAND2_X1 U11704 ( .A1(n9321), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9301) );
  XNOR2_X1 U11705 ( .A(n9301), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10414) );
  AOI22_X1 U11706 ( .A1(n9506), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n10162), 
        .B2(n10414), .ZN(n9302) );
  NAND2_X1 U11707 ( .A1(n9303), .A2(n9302), .ZN(n14616) );
  NAND2_X1 U11708 ( .A1(n9621), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n9309) );
  INV_X1 U11709 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10349) );
  OR2_X1 U11710 ( .A1(n9695), .A2(n10349), .ZN(n9308) );
  INV_X1 U11711 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9304) );
  XNOR2_X1 U11712 ( .A(n9315), .B(n9304), .ZN(n14614) );
  OR2_X1 U11713 ( .A1(n9675), .A2(n14614), .ZN(n9307) );
  INV_X1 U11714 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9305) );
  OR2_X1 U11715 ( .A1(n6424), .A2(n9305), .ZN(n9306) );
  NAND4_X1 U11716 ( .A1(n9309), .A2(n9308), .A3(n9307), .A4(n9306), .ZN(n13568) );
  MUX2_X1 U11717 ( .A(n14616), .B(n13568), .S(n9289), .Z(n9312) );
  INV_X2 U11718 ( .A(n9310), .ZN(n9725) );
  MUX2_X1 U11719 ( .A(n14616), .B(n13568), .S(n9725), .Z(n9311) );
  NAND2_X1 U11720 ( .A1(n9621), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n9320) );
  INV_X1 U11721 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n11513) );
  OR2_X1 U11722 ( .A1(n9695), .A2(n11513), .ZN(n9319) );
  INV_X1 U11723 ( .A(n9315), .ZN(n9313) );
  AOI21_X1 U11724 ( .B1(n9313), .B2(P1_REG3_REG_6__SCAN_IN), .A(
        P1_REG3_REG_7__SCAN_IN), .ZN(n9316) );
  NAND2_X1 U11725 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n9314) );
  NOR2_X1 U11726 ( .A1(n9315), .A2(n9314), .ZN(n9333) );
  OR2_X1 U11727 ( .A1(n9316), .A2(n9333), .ZN(n11515) );
  OR2_X1 U11728 ( .A1(n9675), .A2(n11515), .ZN(n9318) );
  INV_X1 U11729 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10329) );
  OR2_X1 U11730 ( .A1(n6424), .A2(n10329), .ZN(n9317) );
  NAND4_X1 U11731 ( .A1(n9320), .A2(n9319), .A3(n9318), .A4(n9317), .ZN(n13567) );
  NAND2_X1 U11732 ( .A1(n9339), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9322) );
  XNOR2_X1 U11733 ( .A(n9322), .B(P1_IR_REG_7__SCAN_IN), .ZN(n13638) );
  AOI22_X1 U11734 ( .A1(n9506), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n10162), 
        .B2(n13638), .ZN(n9323) );
  NAND2_X1 U11735 ( .A1(n9326), .A2(n9327), .ZN(n9325) );
  MUX2_X1 U11736 ( .A(n11517), .B(n13567), .S(n9289), .Z(n9324) );
  NAND2_X1 U11737 ( .A1(n9325), .A2(n9324), .ZN(n9331) );
  INV_X1 U11738 ( .A(n9326), .ZN(n9329) );
  INV_X1 U11739 ( .A(n9327), .ZN(n9328) );
  NAND2_X1 U11740 ( .A1(n9329), .A2(n9328), .ZN(n9330) );
  NAND2_X1 U11741 ( .A1(n9672), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9338) );
  INV_X1 U11742 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9332) );
  OR2_X1 U11743 ( .A1(n9697), .A2(n9332), .ZN(n9337) );
  NAND2_X1 U11744 ( .A1(n9333), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9347) );
  OR2_X1 U11745 ( .A1(n9333), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9334) );
  NAND2_X1 U11746 ( .A1(n9347), .A2(n9334), .ZN(n11485) );
  OR2_X1 U11747 ( .A1(n9675), .A2(n11485), .ZN(n9336) );
  INV_X1 U11748 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10331) );
  OR2_X1 U11749 ( .A1(n6424), .A2(n10331), .ZN(n9335) );
  NAND4_X1 U11750 ( .A1(n9338), .A2(n9337), .A3(n9336), .A4(n9335), .ZN(n13566) );
  OR2_X1 U11751 ( .A1(n10096), .A2(n9253), .ZN(n9342) );
  NAND2_X1 U11752 ( .A1(n9354), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9340) );
  XNOR2_X1 U11753 ( .A(n9340), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10372) );
  AOI22_X1 U11754 ( .A1(n9506), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n10162), 
        .B2(n10372), .ZN(n9341) );
  NAND2_X1 U11755 ( .A1(n9342), .A2(n9341), .ZN(n11469) );
  MUX2_X1 U11756 ( .A(n13566), .B(n11469), .S(n9725), .Z(n9344) );
  MUX2_X1 U11757 ( .A(n13566), .B(n11469), .S(n9707), .Z(n9343) );
  INV_X1 U11758 ( .A(n9344), .ZN(n9345) );
  NAND2_X1 U11759 ( .A1(n9621), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n9353) );
  INV_X1 U11760 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n11307) );
  OR2_X1 U11761 ( .A1(n9695), .A2(n11307), .ZN(n9352) );
  INV_X1 U11762 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9346) );
  NAND2_X1 U11763 ( .A1(n9347), .A2(n9346), .ZN(n9348) );
  NAND2_X1 U11764 ( .A1(n9368), .A2(n9348), .ZN(n11592) );
  OR2_X1 U11765 ( .A1(n9675), .A2(n11592), .ZN(n9351) );
  INV_X1 U11766 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9349) );
  OR2_X1 U11767 ( .A1(n6424), .A2(n9349), .ZN(n9350) );
  NAND4_X1 U11768 ( .A1(n9353), .A2(n9352), .A3(n9351), .A4(n9350), .ZN(n13565) );
  NAND2_X1 U11769 ( .A1(n10110), .A2(n9715), .ZN(n9359) );
  OAI21_X1 U11770 ( .B1(n9354), .B2(P1_IR_REG_8__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9356) );
  INV_X1 U11771 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9355) );
  OR2_X1 U11772 ( .A1(n9356), .A2(n9355), .ZN(n9357) );
  NAND2_X1 U11773 ( .A1(n9356), .A2(n9355), .ZN(n9374) );
  AOI22_X1 U11774 ( .A1(n9506), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n10162), 
        .B2(n13656), .ZN(n9358) );
  MUX2_X1 U11775 ( .A(n13565), .B(n11594), .S(n9725), .Z(n9360) );
  NAND2_X1 U11776 ( .A1(n9361), .A2(n9360), .ZN(n9367) );
  INV_X1 U11777 ( .A(n9362), .ZN(n9365) );
  INV_X1 U11778 ( .A(n9363), .ZN(n9364) );
  NAND2_X1 U11779 ( .A1(n9365), .A2(n9364), .ZN(n9366) );
  INV_X1 U11780 ( .A(n6425), .ZN(n9512) );
  NAND2_X1 U11781 ( .A1(n9512), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9373) );
  INV_X1 U11782 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14206) );
  OR2_X1 U11783 ( .A1(n9697), .A2(n14206), .ZN(n9372) );
  INV_X1 U11784 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n11433) );
  OR2_X1 U11785 ( .A1(n9695), .A2(n11433), .ZN(n9371) );
  AND2_X1 U11786 ( .A1(n9368), .A2(n10335), .ZN(n9369) );
  OR2_X1 U11787 ( .A1(n9369), .A2(n9399), .ZN(n11759) );
  OR2_X1 U11788 ( .A1(n9675), .A2(n11759), .ZN(n9370) );
  NAND4_X1 U11789 ( .A1(n9373), .A2(n9372), .A3(n9371), .A4(n9370), .ZN(n13564) );
  OR2_X1 U11790 ( .A1(n10207), .A2(n9253), .ZN(n9377) );
  NAND2_X1 U11791 ( .A1(n9374), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9375) );
  XNOR2_X1 U11792 ( .A(n9375), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10426) );
  AOI22_X1 U11793 ( .A1(n10162), .A2(n10426), .B1(n9506), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n9376) );
  MUX2_X1 U11794 ( .A(n13564), .B(n11776), .S(n9725), .Z(n9379) );
  MUX2_X1 U11795 ( .A(n13564), .B(n11776), .S(n9707), .Z(n9378) );
  INV_X1 U11796 ( .A(n9379), .ZN(n9380) );
  NAND2_X1 U11797 ( .A1(n9672), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9386) );
  INV_X1 U11798 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9381) );
  OR2_X1 U11799 ( .A1(n9697), .A2(n9381), .ZN(n9385) );
  XNOR2_X1 U11800 ( .A(n9399), .B(P1_REG3_REG_11__SCAN_IN), .ZN(n11795) );
  OR2_X1 U11801 ( .A1(n9675), .A2(n11795), .ZN(n9384) );
  INV_X1 U11802 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9382) );
  OR2_X1 U11803 ( .A1(n6425), .A2(n9382), .ZN(n9383) );
  NAND4_X1 U11804 ( .A1(n9386), .A2(n9385), .A3(n9384), .A4(n9383), .ZN(n13563) );
  NAND2_X1 U11805 ( .A1(n10282), .A2(n9715), .ZN(n9389) );
  OR2_X1 U11806 ( .A1(n7317), .A2(n9445), .ZN(n9387) );
  XNOR2_X1 U11807 ( .A(n9387), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10519) );
  AOI22_X1 U11808 ( .A1(n9506), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n10162), 
        .B2(n10519), .ZN(n9388) );
  NAND2_X1 U11809 ( .A1(n9392), .A2(n9393), .ZN(n9391) );
  MUX2_X1 U11810 ( .A(n13563), .B(n11797), .S(n9725), .Z(n9390) );
  NAND2_X1 U11811 ( .A1(n9391), .A2(n9390), .ZN(n9397) );
  INV_X1 U11812 ( .A(n9392), .ZN(n9395) );
  INV_X1 U11813 ( .A(n9393), .ZN(n9394) );
  NAND2_X1 U11814 ( .A1(n9395), .A2(n9394), .ZN(n9396) );
  NAND2_X1 U11815 ( .A1(n9621), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n9404) );
  AND2_X1 U11816 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .ZN(n9398) );
  AOI21_X1 U11817 ( .B1(n9399), .B2(P1_REG3_REG_11__SCAN_IN), .A(
        P1_REG3_REG_12__SCAN_IN), .ZN(n9400) );
  OR2_X1 U11818 ( .A1(n9413), .A2(n9400), .ZN(n11887) );
  OR2_X1 U11819 ( .A1(n9675), .A2(n11887), .ZN(n9403) );
  INV_X1 U11820 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10525) );
  OR2_X1 U11821 ( .A1(n6425), .A2(n10525), .ZN(n9402) );
  INV_X1 U11822 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11687) );
  OR2_X1 U11823 ( .A1(n9695), .A2(n11687), .ZN(n9401) );
  NAND4_X1 U11824 ( .A1(n9404), .A2(n9403), .A3(n9402), .A4(n9401), .ZN(n13562) );
  NAND2_X1 U11825 ( .A1(n10439), .A2(n9715), .ZN(n9410) );
  INV_X1 U11826 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9405) );
  NAND2_X1 U11827 ( .A1(n7317), .A2(n9405), .ZN(n9407) );
  NAND2_X1 U11828 ( .A1(n9407), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9406) );
  MUX2_X1 U11829 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9406), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n9408) );
  AOI22_X1 U11830 ( .A1(n9506), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n10162), 
        .B2(n10532), .ZN(n9409) );
  MUX2_X1 U11831 ( .A(n13562), .B(n11884), .S(n9725), .Z(n9412) );
  MUX2_X1 U11832 ( .A(n13562), .B(n11884), .S(n9707), .Z(n9411) );
  NAND2_X1 U11833 ( .A1(n9621), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n9418) );
  INV_X1 U11834 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10924) );
  OR2_X1 U11835 ( .A1(n6425), .A2(n10924), .ZN(n9417) );
  NAND2_X1 U11836 ( .A1(n9413), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9435) );
  OR2_X1 U11837 ( .A1(n9413), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9414) );
  NAND2_X1 U11838 ( .A1(n9435), .A2(n9414), .ZN(n11932) );
  OR2_X1 U11839 ( .A1(n9675), .A2(n11932), .ZN(n9416) );
  INV_X1 U11840 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11719) );
  OR2_X1 U11841 ( .A1(n9695), .A2(n11719), .ZN(n9415) );
  NAND4_X1 U11842 ( .A1(n9418), .A2(n9417), .A3(n9416), .A4(n9415), .ZN(n13561) );
  OR2_X1 U11843 ( .A1(n10444), .A2(n9253), .ZN(n9423) );
  NAND2_X1 U11844 ( .A1(n9420), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9419) );
  MUX2_X1 U11845 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9419), .S(
        P1_IR_REG_13__SCAN_IN), .Z(n9421) );
  AOI22_X1 U11846 ( .A1(n9506), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n10162), 
        .B2(n14596), .ZN(n9422) );
  MUX2_X1 U11847 ( .A(n13561), .B(n11934), .S(n9289), .Z(n9427) );
  NAND2_X1 U11848 ( .A1(n9426), .A2(n9427), .ZN(n9425) );
  MUX2_X1 U11849 ( .A(n13561), .B(n11934), .S(n9725), .Z(n9424) );
  NAND2_X1 U11850 ( .A1(n9425), .A2(n9424), .ZN(n9443) );
  INV_X1 U11851 ( .A(n9426), .ZN(n9429) );
  INV_X1 U11852 ( .A(n9427), .ZN(n9428) );
  NAND2_X1 U11853 ( .A1(n9429), .A2(n9428), .ZN(n9442) );
  NAND2_X1 U11854 ( .A1(n10645), .A2(n9715), .ZN(n9433) );
  NAND2_X1 U11855 ( .A1(n9430), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9431) );
  XNOR2_X1 U11856 ( .A(n9431), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11342) );
  AOI22_X1 U11857 ( .A1(n9506), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n10162), 
        .B2(n11342), .ZN(n9432) );
  NAND2_X1 U11858 ( .A1(n9621), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n9441) );
  INV_X1 U11859 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11839) );
  OR2_X1 U11860 ( .A1(n9695), .A2(n11839), .ZN(n9440) );
  NAND2_X1 U11861 ( .A1(n9435), .A2(n9434), .ZN(n9436) );
  NAND2_X1 U11862 ( .A1(n9450), .A2(n9436), .ZN(n12011) );
  OR2_X1 U11863 ( .A1(n9675), .A2(n12011), .ZN(n9439) );
  INV_X1 U11864 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9437) );
  OR2_X1 U11865 ( .A1(n6424), .A2(n9437), .ZN(n9438) );
  NAND2_X1 U11866 ( .A1(n14528), .A2(n13992), .ZN(n9457) );
  NAND2_X1 U11867 ( .A1(n13733), .A2(n9457), .ZN(n11835) );
  NAND2_X1 U11868 ( .A1(n10893), .A2(n9715), .ZN(n9448) );
  OR2_X1 U11869 ( .A1(n9444), .A2(n9445), .ZN(n9446) );
  XNOR2_X1 U11870 ( .A(n9446), .B(P1_IR_REG_15__SCAN_IN), .ZN(n11607) );
  AOI22_X1 U11871 ( .A1(n9506), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n10162), 
        .B2(n11607), .ZN(n9447) );
  NAND2_X1 U11872 ( .A1(n9621), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n9456) );
  INV_X1 U11873 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9449) );
  OR2_X1 U11874 ( .A1(n9695), .A2(n9449), .ZN(n9455) );
  NAND2_X1 U11875 ( .A1(n9450), .A2(n14183), .ZN(n9451) );
  NAND2_X1 U11876 ( .A1(n9484), .A2(n9451), .ZN(n13999) );
  OR2_X1 U11877 ( .A1(n9675), .A2(n13999), .ZN(n9454) );
  INV_X1 U11878 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9452) );
  OR2_X1 U11879 ( .A1(n6425), .A2(n9452), .ZN(n9453) );
  NAND2_X1 U11880 ( .A1(n14522), .A2(n12051), .ZN(n9734) );
  NAND2_X1 U11881 ( .A1(n9734), .A2(n9457), .ZN(n9459) );
  NAND2_X1 U11882 ( .A1(n13735), .A2(n13733), .ZN(n9458) );
  MUX2_X1 U11883 ( .A(n9459), .B(n9458), .S(n9707), .Z(n9461) );
  MUX2_X1 U11884 ( .A(n9734), .B(n13735), .S(n9725), .Z(n9460) );
  NAND2_X1 U11885 ( .A1(n11206), .A2(n9715), .ZN(n9465) );
  INV_X1 U11886 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9462) );
  NAND2_X1 U11887 ( .A1(n9444), .A2(n9462), .ZN(n9491) );
  NAND2_X1 U11888 ( .A1(n9473), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9463) );
  XNOR2_X1 U11889 ( .A(n9463), .B(P1_IR_REG_18__SCAN_IN), .ZN(n13683) );
  AOI22_X1 U11890 ( .A1(n9506), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n10162), 
        .B2(n13683), .ZN(n9464) );
  NAND2_X1 U11891 ( .A1(n9486), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9478) );
  INV_X1 U11892 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9466) );
  NAND2_X1 U11893 ( .A1(n9478), .A2(n9466), .ZN(n9467) );
  AND2_X1 U11894 ( .A1(n9510), .A2(n9467), .ZN(n13945) );
  INV_X1 U11895 ( .A(n9675), .ZN(n9551) );
  NAND2_X1 U11896 ( .A1(n13945), .A2(n9551), .ZN(n9471) );
  AOI22_X1 U11897 ( .A1(n9672), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9621), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n9470) );
  INV_X1 U11898 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9468) );
  OR2_X1 U11899 ( .A1(n6425), .A2(n9468), .ZN(n9469) );
  NAND2_X1 U11900 ( .A1(n13946), .A2(n13955), .ZN(n9516) );
  NAND2_X1 U11901 ( .A1(n13741), .A2(n9516), .ZN(n13940) );
  NAND2_X1 U11902 ( .A1(n11104), .A2(n9715), .ZN(n9476) );
  NAND2_X1 U11903 ( .A1(n9493), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9472) );
  MUX2_X1 U11904 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9472), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n9474) );
  AND2_X1 U11905 ( .A1(n9474), .A2(n9473), .ZN(n11704) );
  AOI22_X1 U11906 ( .A1(n9506), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n10162), 
        .B2(n11704), .ZN(n9475) );
  OR2_X1 U11907 ( .A1(n9486), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9477) );
  NAND2_X1 U11908 ( .A1(n9478), .A2(n9477), .ZN(n13954) );
  INV_X1 U11909 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n13669) );
  OAI22_X1 U11910 ( .A1(n13954), .A2(n9675), .B1(n6424), .B2(n13669), .ZN(
        n9481) );
  INV_X1 U11911 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n13959) );
  NAND2_X1 U11912 ( .A1(n9621), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n9479) );
  OAI21_X1 U11913 ( .B1(n9695), .B2(n13959), .A(n9479), .ZN(n9480) );
  NAND2_X1 U11914 ( .A1(n14232), .A2(n13984), .ZN(n13714) );
  OR2_X1 U11915 ( .A1(n14232), .A2(n13984), .ZN(n9482) );
  NOR2_X1 U11916 ( .A1(n13940), .A2(n13713), .ZN(n9499) );
  AND2_X1 U11917 ( .A1(n9484), .A2(n9483), .ZN(n9485) );
  NOR2_X1 U11918 ( .A1(n9486), .A2(n9485), .ZN(n13975) );
  NAND2_X1 U11919 ( .A1(n13975), .A2(n9551), .ZN(n9490) );
  NAND2_X1 U11920 ( .A1(n9621), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n9489) );
  NAND2_X1 U11921 ( .A1(n9672), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9488) );
  NAND2_X1 U11922 ( .A1(n9512), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9487) );
  NAND2_X1 U11923 ( .A1(n10981), .A2(n9715), .ZN(n9496) );
  NAND2_X1 U11924 ( .A1(n9491), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9492) );
  MUX2_X1 U11925 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9492), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n9494) );
  AND2_X1 U11926 ( .A1(n9494), .A2(n9493), .ZN(n11610) );
  AOI22_X1 U11927 ( .A1(n9506), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n10162), 
        .B2(n11610), .ZN(n9495) );
  MUX2_X1 U11928 ( .A(n13994), .B(n13977), .S(n9707), .Z(n9501) );
  INV_X1 U11929 ( .A(n13994), .ZN(n13560) );
  MUX2_X1 U11930 ( .A(n13560), .B(n14240), .S(n9725), .Z(n9500) );
  NAND2_X1 U11931 ( .A1(n9501), .A2(n9500), .ZN(n9497) );
  INV_X1 U11932 ( .A(n9499), .ZN(n9502) );
  OR3_X1 U11933 ( .A1(n9502), .A2(n9501), .A3(n9500), .ZN(n9520) );
  NAND2_X1 U11934 ( .A1(n9725), .A2(n13984), .ZN(n9504) );
  INV_X1 U11935 ( .A(n13984), .ZN(n13739) );
  NAND3_X1 U11936 ( .A1(n14232), .A2(n13739), .A3(n9289), .ZN(n9503) );
  OAI21_X1 U11937 ( .B1(n14232), .B2(n9504), .A(n9503), .ZN(n9505) );
  NAND2_X1 U11938 ( .A1(n13935), .A2(n9505), .ZN(n9515) );
  NAND2_X1 U11939 ( .A1(n11264), .A2(n9715), .ZN(n9508) );
  INV_X1 U11940 ( .A(n11268), .ZN(n13691) );
  AOI22_X1 U11941 ( .A1(n9506), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n13691), 
        .B2(n10162), .ZN(n9507) );
  INV_X1 U11942 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9509) );
  AND2_X1 U11943 ( .A1(n9510), .A2(n9509), .ZN(n9511) );
  OR2_X1 U11944 ( .A1(n9511), .A2(n9524), .ZN(n13923) );
  AOI22_X1 U11945 ( .A1(n9512), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n9621), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n9514) );
  NAND2_X1 U11946 ( .A1(n9672), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n9513) );
  OAI211_X1 U11947 ( .C1(n13923), .C2(n9675), .A(n9514), .B(n9513), .ZN(n13903) );
  INV_X1 U11948 ( .A(n13903), .ZN(n9736) );
  NAND2_X1 U11949 ( .A1(n14221), .A2(n9736), .ZN(n13742) );
  OAI211_X1 U11950 ( .C1(n9725), .C2(n9516), .A(n9515), .B(n13742), .ZN(n9518)
         );
  OR2_X1 U11951 ( .A1(n14221), .A2(n9736), .ZN(n9521) );
  AOI21_X1 U11952 ( .B1(n9521), .B2(n13741), .A(n9289), .ZN(n9517) );
  NOR2_X1 U11953 ( .A1(n9518), .A2(n9517), .ZN(n9519) );
  MUX2_X1 U11954 ( .A(n13742), .B(n9521), .S(n9707), .Z(n9522) );
  NOR2_X1 U11955 ( .A1(n9524), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n9525) );
  OR2_X1 U11956 ( .A1(n9537), .A2(n9525), .ZN(n13912) );
  INV_X1 U11957 ( .A(n13912), .ZN(n9529) );
  INV_X1 U11958 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n14085) );
  NAND2_X1 U11959 ( .A1(n9621), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n9527) );
  NAND2_X1 U11960 ( .A1(n9672), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n9526) );
  OAI211_X1 U11961 ( .C1(n6425), .C2(n14085), .A(n9527), .B(n9526), .ZN(n9528)
         );
  AOI21_X1 U11962 ( .B1(n9529), .B2(n9551), .A(n9528), .ZN(n13743) );
  OR2_X1 U11963 ( .A1(n11534), .A2(n9253), .ZN(n9531) );
  OR2_X1 U11964 ( .A1(n9716), .A2(n11533), .ZN(n9530) );
  MUX2_X1 U11965 ( .A(n13743), .B(n14082), .S(n9289), .Z(n9533) );
  INV_X1 U11966 ( .A(n13743), .ZN(n13559) );
  MUX2_X1 U11967 ( .A(n13559), .B(n13915), .S(n9725), .Z(n9532) );
  OAI21_X1 U11968 ( .B1(n9534), .B2(n9533), .A(n9532), .ZN(n9536) );
  NAND2_X1 U11969 ( .A1(n9534), .A2(n9533), .ZN(n9535) );
  NOR2_X1 U11970 ( .A1(n9537), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9538) );
  OR2_X1 U11971 ( .A1(n9549), .A2(n9538), .ZN(n13890) );
  INV_X1 U11972 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9541) );
  NAND2_X1 U11973 ( .A1(n9672), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9540) );
  NAND2_X1 U11974 ( .A1(n9621), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9539) );
  OAI211_X1 U11975 ( .C1(n9541), .C2(n6424), .A(n9540), .B(n9539), .ZN(n9542)
         );
  INV_X1 U11976 ( .A(n9542), .ZN(n9543) );
  OAI21_X1 U11977 ( .B1(n13890), .B2(n9675), .A(n9543), .ZN(n13904) );
  OR2_X1 U11978 ( .A1(n11649), .A2(n9253), .ZN(n9545) );
  OR2_X1 U11979 ( .A1(n9716), .A2(n14126), .ZN(n9544) );
  MUX2_X1 U11980 ( .A(n13904), .B(n14073), .S(n9725), .Z(n9547) );
  MUX2_X1 U11981 ( .A(n13904), .B(n14073), .S(n9707), .Z(n9546) );
  INV_X1 U11982 ( .A(n9547), .ZN(n9548) );
  OR2_X1 U11983 ( .A1(n9549), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9550) );
  NAND2_X1 U11984 ( .A1(n9549), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9568) );
  AND2_X1 U11985 ( .A1(n9550), .A2(n9568), .ZN(n13878) );
  NAND2_X1 U11986 ( .A1(n13878), .A2(n9551), .ZN(n9556) );
  INV_X1 U11987 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n14124) );
  NAND2_X1 U11988 ( .A1(n9672), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9553) );
  NAND2_X1 U11989 ( .A1(n9621), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n9552) );
  OAI211_X1 U11990 ( .C1(n14124), .C2(n6425), .A(n9553), .B(n9552), .ZN(n9554)
         );
  INV_X1 U11991 ( .A(n9554), .ZN(n9555) );
  NAND2_X1 U11992 ( .A1(n9556), .A2(n9555), .ZN(n13745) );
  OR2_X1 U11993 ( .A1(n7853), .A2(n10049), .ZN(n9557) );
  XNOR2_X1 U11994 ( .A(n9557), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14283) );
  NAND2_X1 U11995 ( .A1(n9561), .A2(n9562), .ZN(n9560) );
  MUX2_X1 U11996 ( .A(n13745), .B(n13875), .S(n9725), .Z(n9559) );
  NAND2_X1 U11997 ( .A1(n9560), .A2(n9559), .ZN(n9566) );
  INV_X1 U11998 ( .A(n9561), .ZN(n9564) );
  INV_X1 U11999 ( .A(n9562), .ZN(n9563) );
  NAND2_X1 U12000 ( .A1(n9564), .A2(n9563), .ZN(n9565) );
  NAND2_X1 U12001 ( .A1(n9566), .A2(n9565), .ZN(n9579) );
  NAND2_X1 U12002 ( .A1(n9672), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9574) );
  INV_X1 U12003 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9567) );
  OR2_X1 U12004 ( .A1(n9697), .A2(n9567), .ZN(n9573) );
  NAND2_X1 U12005 ( .A1(n9569), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n9586) );
  OAI21_X1 U12006 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n9569), .A(n9586), .ZN(
        n13859) );
  OR2_X1 U12007 ( .A1(n9675), .A2(n13859), .ZN(n9572) );
  INV_X1 U12008 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9570) );
  OR2_X1 U12009 ( .A1(n6424), .A2(n9570), .ZN(n9571) );
  NAND4_X1 U12010 ( .A1(n9574), .A2(n9573), .A3(n9572), .A4(n9571), .ZN(n13721) );
  OR2_X1 U12011 ( .A1(n9716), .A2(n9575), .ZN(n9576) );
  NAND2_X1 U12012 ( .A1(n9579), .A2(n9580), .ZN(n9578) );
  MUX2_X1 U12013 ( .A(n13721), .B(n14058), .S(n9707), .Z(n9577) );
  NAND2_X1 U12014 ( .A1(n9578), .A2(n9577), .ZN(n9584) );
  INV_X1 U12015 ( .A(n9579), .ZN(n9582) );
  INV_X1 U12016 ( .A(n9580), .ZN(n9581) );
  NAND2_X1 U12017 ( .A1(n9582), .A2(n9581), .ZN(n9583) );
  NAND2_X1 U12018 ( .A1(n9672), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n9592) );
  INV_X1 U12019 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9585) );
  OR2_X1 U12020 ( .A1(n9697), .A2(n9585), .ZN(n9591) );
  NAND2_X1 U12021 ( .A1(n9587), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n9604) );
  OAI21_X1 U12022 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n9587), .A(n9604), .ZN(
        n13504) );
  OR2_X1 U12023 ( .A1(n9675), .A2(n13504), .ZN(n9590) );
  INV_X1 U12024 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9588) );
  OR2_X1 U12025 ( .A1(n6424), .A2(n9588), .ZN(n9589) );
  NAND4_X1 U12026 ( .A1(n9592), .A2(n9591), .A3(n9590), .A4(n9589), .ZN(n13725) );
  OR2_X1 U12027 ( .A1(n12019), .A2(n9253), .ZN(n9594) );
  INV_X1 U12028 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12018) );
  OR2_X1 U12029 ( .A1(n9716), .A2(n12018), .ZN(n9593) );
  NAND2_X2 U12030 ( .A1(n9594), .A2(n9593), .ZN(n14051) );
  NAND2_X1 U12031 ( .A1(n9597), .A2(n9598), .ZN(n9596) );
  MUX2_X1 U12032 ( .A(n14051), .B(n13725), .S(n9707), .Z(n9595) );
  NAND2_X1 U12033 ( .A1(n9596), .A2(n9595), .ZN(n9602) );
  INV_X1 U12034 ( .A(n9597), .ZN(n9600) );
  INV_X1 U12035 ( .A(n9598), .ZN(n9599) );
  NAND2_X1 U12036 ( .A1(n9600), .A2(n9599), .ZN(n9601) );
  NAND2_X1 U12037 ( .A1(n9602), .A2(n9601), .ZN(n9615) );
  NAND2_X1 U12038 ( .A1(n9672), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n9610) );
  INV_X1 U12039 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9603) );
  OR2_X1 U12040 ( .A1(n9697), .A2(n9603), .ZN(n9609) );
  NAND2_X1 U12041 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n9605), .ZN(n9624) );
  OAI21_X1 U12042 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n9605), .A(n9624), .ZN(
        n13827) );
  OR2_X1 U12043 ( .A1(n9675), .A2(n13827), .ZN(n9608) );
  INV_X1 U12044 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9606) );
  OR2_X1 U12045 ( .A1(n6425), .A2(n9606), .ZN(n9607) );
  NAND4_X1 U12046 ( .A1(n9610), .A2(n9609), .A3(n9608), .A4(n9607), .ZN(n13728) );
  NAND2_X1 U12047 ( .A1(n13436), .A2(n9715), .ZN(n9612) );
  OR2_X1 U12048 ( .A1(n9716), .A2(n14279), .ZN(n9611) );
  NAND2_X2 U12049 ( .A1(n9612), .A2(n9611), .ZN(n14045) );
  MUX2_X1 U12050 ( .A(n13728), .B(n14045), .S(n9725), .Z(n9616) );
  NAND2_X1 U12051 ( .A1(n9615), .A2(n9616), .ZN(n9614) );
  MUX2_X1 U12052 ( .A(n13728), .B(n14045), .S(n9289), .Z(n9613) );
  NAND2_X1 U12053 ( .A1(n9614), .A2(n9613), .ZN(n9620) );
  INV_X1 U12054 ( .A(n9615), .ZN(n9618) );
  INV_X1 U12055 ( .A(n9616), .ZN(n9617) );
  NAND2_X1 U12056 ( .A1(n9618), .A2(n9617), .ZN(n9619) );
  NAND2_X1 U12057 ( .A1(n9621), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n9630) );
  INV_X1 U12058 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9622) );
  OR2_X1 U12059 ( .A1(n9695), .A2(n9622), .ZN(n9629) );
  INV_X1 U12060 ( .A(n9624), .ZN(n9623) );
  NAND2_X1 U12061 ( .A1(n9623), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n9643) );
  INV_X1 U12062 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n13539) );
  NAND2_X1 U12063 ( .A1(n9624), .A2(n13539), .ZN(n9625) );
  NAND2_X1 U12064 ( .A1(n9643), .A2(n9625), .ZN(n13815) );
  OR2_X1 U12065 ( .A1(n9675), .A2(n13815), .ZN(n9628) );
  INV_X1 U12066 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9626) );
  OR2_X1 U12067 ( .A1(n6424), .A2(n9626), .ZN(n9627) );
  NAND4_X1 U12068 ( .A1(n9630), .A2(n9629), .A3(n9628), .A4(n9627), .ZN(n13749) );
  NAND2_X1 U12069 ( .A1(n13432), .A2(n9715), .ZN(n9632) );
  OR2_X1 U12070 ( .A1(n9716), .A2(n14275), .ZN(n9631) );
  NAND2_X1 U12071 ( .A1(n9635), .A2(n9636), .ZN(n9634) );
  MUX2_X1 U12072 ( .A(n13749), .B(n13817), .S(n9724), .Z(n9633) );
  NAND2_X1 U12073 ( .A1(n9634), .A2(n9633), .ZN(n9640) );
  INV_X1 U12074 ( .A(n9635), .ZN(n9638) );
  INV_X1 U12075 ( .A(n9636), .ZN(n9637) );
  NAND2_X1 U12076 ( .A1(n9638), .A2(n9637), .ZN(n9639) );
  NAND2_X1 U12077 ( .A1(n9672), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9649) );
  INV_X1 U12078 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9641) );
  OR2_X1 U12079 ( .A1(n9697), .A2(n9641), .ZN(n9648) );
  INV_X1 U12080 ( .A(n9643), .ZN(n9642) );
  NAND2_X1 U12081 ( .A1(n9642), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n9673) );
  INV_X1 U12082 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n13447) );
  NAND2_X1 U12083 ( .A1(n9643), .A2(n13447), .ZN(n9644) );
  NAND2_X1 U12084 ( .A1(n9673), .A2(n9644), .ZN(n13446) );
  OR2_X1 U12085 ( .A1(n9675), .A2(n13446), .ZN(n9647) );
  INV_X1 U12086 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9645) );
  OR2_X1 U12087 ( .A1(n6425), .A2(n9645), .ZN(n9646) );
  NAND4_X1 U12088 ( .A1(n9649), .A2(n9648), .A3(n9647), .A4(n9646), .ZN(n13774) );
  NAND2_X1 U12089 ( .A1(n12023), .A2(n9715), .ZN(n9651) );
  OR2_X1 U12090 ( .A1(n9716), .A2(n14273), .ZN(n9650) );
  MUX2_X1 U12091 ( .A(n13774), .B(n14034), .S(n9725), .Z(n9653) );
  MUX2_X1 U12092 ( .A(n13774), .B(n14034), .S(n9289), .Z(n9652) );
  INV_X1 U12093 ( .A(n9653), .ZN(n9654) );
  NAND2_X1 U12094 ( .A1(n9672), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9660) );
  INV_X1 U12095 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9655) );
  OR2_X1 U12096 ( .A1(n9697), .A2(n9655), .ZN(n9659) );
  INV_X1 U12097 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9656) );
  XNOR2_X1 U12098 ( .A(n9673), .B(n9656), .ZN(n13780) );
  OR2_X1 U12099 ( .A1(n9675), .A2(n13780), .ZN(n9658) );
  INV_X1 U12100 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n14195) );
  OR2_X1 U12101 ( .A1(n6424), .A2(n14195), .ZN(n9657) );
  NAND4_X1 U12102 ( .A1(n9660), .A2(n9659), .A3(n9658), .A4(n9657), .ZN(n13765) );
  NAND2_X1 U12103 ( .A1(n12021), .A2(n9715), .ZN(n9662) );
  OR2_X1 U12104 ( .A1(n9716), .A2(n12022), .ZN(n9661) );
  MUX2_X1 U12105 ( .A(n13765), .B(n14028), .S(n9707), .Z(n9666) );
  NAND2_X1 U12106 ( .A1(n9665), .A2(n9666), .ZN(n9664) );
  MUX2_X1 U12107 ( .A(n14028), .B(n13765), .S(n9289), .Z(n9663) );
  INV_X1 U12108 ( .A(n9665), .ZN(n9668) );
  INV_X1 U12109 ( .A(n9666), .ZN(n9667) );
  NAND2_X1 U12110 ( .A1(n9669), .A2(n9715), .ZN(n9671) );
  OR2_X1 U12111 ( .A1(n9716), .A2(n12030), .ZN(n9670) );
  NAND2_X1 U12112 ( .A1(n9672), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9680) );
  INV_X1 U12113 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n14199) );
  OR2_X1 U12114 ( .A1(n9697), .A2(n14199), .ZN(n9679) );
  INV_X1 U12115 ( .A(n9673), .ZN(n9674) );
  NAND2_X1 U12116 ( .A1(n9674), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n13764) );
  OR2_X1 U12117 ( .A1(n9675), .A2(n13764), .ZN(n9678) );
  INV_X1 U12118 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9676) );
  OR2_X1 U12119 ( .A1(n6425), .A2(n9676), .ZN(n9677) );
  MUX2_X1 U12120 ( .A(n14020), .B(n9681), .S(n9707), .Z(n9683) );
  MUX2_X1 U12121 ( .A(n13773), .B(n13758), .S(n9289), .Z(n9682) );
  INV_X1 U12122 ( .A(n9683), .ZN(n9684) );
  INV_X1 U12123 ( .A(n9711), .ZN(n9714) );
  OR2_X1 U12124 ( .A1(n9716), .A2(n14271), .ZN(n9685) );
  INV_X1 U12125 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9687) );
  OR2_X1 U12126 ( .A1(n6425), .A2(n9687), .ZN(n9691) );
  INV_X1 U12127 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n13705) );
  OR2_X1 U12128 ( .A1(n9695), .A2(n13705), .ZN(n9690) );
  INV_X1 U12129 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9688) );
  OR2_X1 U12130 ( .A1(n9697), .A2(n9688), .ZN(n9689) );
  AND3_X1 U12131 ( .A1(n9691), .A2(n9690), .A3(n9689), .ZN(n9705) );
  INV_X1 U12132 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9692) );
  NOR2_X1 U12133 ( .A1(n6424), .A2(n9692), .ZN(n9700) );
  INV_X1 U12134 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9694) );
  NOR2_X1 U12135 ( .A1(n9695), .A2(n9694), .ZN(n9699) );
  INV_X1 U12136 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9696) );
  NOR2_X1 U12137 ( .A1(n9697), .A2(n9696), .ZN(n9698) );
  INV_X1 U12138 ( .A(n9701), .ZN(n9702) );
  AOI21_X1 U12139 ( .B1(n9725), .B2(n13699), .A(n9702), .ZN(n9703) );
  OAI22_X1 U12140 ( .A1(n14016), .A2(n9725), .B1(n9705), .B2(n9703), .ZN(n9710) );
  INV_X1 U12141 ( .A(n9710), .ZN(n9713) );
  INV_X1 U12142 ( .A(n9704), .ZN(n9706) );
  INV_X1 U12143 ( .A(n9705), .ZN(n13760) );
  OAI21_X1 U12144 ( .B1(n13699), .B2(n9706), .A(n13760), .ZN(n9708) );
  MUX2_X1 U12145 ( .A(n14016), .B(n9708), .S(n9707), .Z(n9709) );
  NAND2_X1 U12146 ( .A1(n14268), .A2(n9715), .ZN(n9718) );
  INV_X1 U12147 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14264) );
  OR2_X1 U12148 ( .A1(n9716), .A2(n14264), .ZN(n9717) );
  XOR2_X1 U12149 ( .A(n13699), .B(n9755), .Z(n9746) );
  NAND2_X1 U12150 ( .A1(n9719), .A2(n11085), .ZN(n10604) );
  INV_X1 U12151 ( .A(n9719), .ZN(n9721) );
  NAND2_X1 U12152 ( .A1(n9721), .A2(n9720), .ZN(n11086) );
  NAND2_X1 U12153 ( .A1(n10604), .A2(n11086), .ZN(n9722) );
  INV_X1 U12154 ( .A(n10591), .ZN(n10595) );
  NAND2_X1 U12155 ( .A1(n10595), .A2(n13691), .ZN(n11137) );
  NAND2_X1 U12156 ( .A1(n9722), .A2(n11137), .ZN(n9752) );
  NOR2_X1 U12157 ( .A1(n9746), .A2(n9752), .ZN(n9723) );
  AND2_X1 U12158 ( .A1(n9766), .A2(n9723), .ZN(n9774) );
  NOR2_X1 U12159 ( .A1(n9755), .A2(n9724), .ZN(n9751) );
  NAND2_X1 U12160 ( .A1(n11650), .A2(n11257), .ZN(n11088) );
  NAND2_X1 U12161 ( .A1(n9752), .A2(n11088), .ZN(n9754) );
  NAND2_X1 U12162 ( .A1(n9755), .A2(n9725), .ZN(n9761) );
  NOR2_X1 U12163 ( .A1(n9761), .A2(n13699), .ZN(n9726) );
  AOI211_X1 U12164 ( .C1(n9751), .C2(n13699), .A(n9754), .B(n9726), .ZN(n9727)
         );
  INV_X1 U12165 ( .A(n9727), .ZN(n9765) );
  INV_X1 U12166 ( .A(n14016), .ZN(n13707) );
  XNOR2_X1 U12167 ( .A(n13707), .B(n13760), .ZN(n9744) );
  INV_X1 U12168 ( .A(n13749), .ZN(n12141) );
  XNOR2_X1 U12169 ( .A(n13817), .B(n12141), .ZN(n13811) );
  XNOR2_X1 U12170 ( .A(n14045), .B(n13728), .ZN(n13835) );
  INV_X1 U12171 ( .A(n13721), .ZN(n13746) );
  XNOR2_X1 U12172 ( .A(n14066), .B(n13745), .ZN(n13873) );
  XNOR2_X1 U12173 ( .A(n13915), .B(n13743), .ZN(n13717) );
  INV_X1 U12174 ( .A(n13904), .ZN(n13744) );
  XNOR2_X1 U12175 ( .A(n14073), .B(n13744), .ZN(n13897) );
  INV_X1 U12176 ( .A(n13561), .ZN(n11928) );
  XNOR2_X1 U12177 ( .A(n11934), .B(n11928), .ZN(n11846) );
  XNOR2_X1 U12178 ( .A(n11594), .B(n11582), .ZN(n11429) );
  INV_X1 U12179 ( .A(n13566), .ZN(n11467) );
  XNOR2_X1 U12180 ( .A(n11469), .B(n11467), .ZN(n11365) );
  XNOR2_X1 U12181 ( .A(n11517), .B(n13567), .ZN(n11509) );
  INV_X1 U12182 ( .A(n11258), .ZN(n9728) );
  INV_X1 U12183 ( .A(n11073), .ZN(n13572) );
  NAND4_X1 U12184 ( .A1(n9728), .A2(n11186), .A3(n11131), .A4(n14630), .ZN(
        n9729) );
  XNOR2_X1 U12185 ( .A(n11077), .B(n11274), .ZN(n11069) );
  NOR2_X1 U12186 ( .A1(n9729), .A2(n11069), .ZN(n9730) );
  XNOR2_X1 U12187 ( .A(n14616), .B(n13568), .ZN(n14611) );
  XNOR2_X1 U12188 ( .A(n11293), .B(n13569), .ZN(n11079) );
  NAND4_X1 U12189 ( .A1(n11509), .A2(n9730), .A3(n14611), .A4(n11079), .ZN(
        n9731) );
  OR4_X1 U12190 ( .A1(n11549), .A2(n11429), .A3(n11365), .A4(n9731), .ZN(n9732) );
  INV_X1 U12191 ( .A(n13562), .ZN(n11882) );
  XNOR2_X1 U12192 ( .A(n11884), .B(n11882), .ZN(n11714) );
  XNOR2_X1 U12193 ( .A(n11797), .B(n11781), .ZN(n11676) );
  OR4_X1 U12194 ( .A1(n11846), .A2(n9732), .A3(n11714), .A4(n11676), .ZN(n9735) );
  NAND2_X1 U12195 ( .A1(n14240), .A2(n13994), .ZN(n13738) );
  OR2_X1 U12196 ( .A1(n14240), .A2(n13994), .ZN(n9733) );
  NAND2_X1 U12197 ( .A1(n13738), .A2(n9733), .ZN(n13737) );
  NAND2_X1 U12198 ( .A1(n13735), .A2(n9734), .ZN(n13989) );
  OR4_X1 U12199 ( .A1(n9735), .A2(n13737), .A3(n13989), .A4(n11835), .ZN(n9737) );
  XNOR2_X1 U12200 ( .A(n14221), .B(n9736), .ZN(n13928) );
  OR4_X1 U12201 ( .A1(n9737), .A2(n13928), .A3(n13713), .A4(n13940), .ZN(n9738) );
  OR4_X1 U12202 ( .A1(n13873), .A2(n13717), .A3(n13897), .A4(n9738), .ZN(n9739) );
  NOR2_X1 U12203 ( .A1(n13863), .A2(n9739), .ZN(n9740) );
  XNOR2_X1 U12204 ( .A(n14051), .B(n13725), .ZN(n13851) );
  NAND3_X1 U12205 ( .A1(n13835), .A2(n9740), .A3(n13851), .ZN(n9741) );
  NOR2_X1 U12206 ( .A1(n13811), .A2(n9741), .ZN(n9743) );
  XNOR2_X1 U12207 ( .A(n14034), .B(n13774), .ZN(n13791) );
  NAND2_X1 U12208 ( .A1(n14028), .A2(n13765), .ZN(n13732) );
  OR2_X1 U12209 ( .A1(n14028), .A2(n13765), .ZN(n9742) );
  NAND2_X1 U12210 ( .A1(n13732), .A2(n9742), .ZN(n13784) );
  NAND4_X1 U12211 ( .A1(n9744), .A2(n9743), .A3(n13791), .A4(n13784), .ZN(
        n9745) );
  NOR3_X1 U12212 ( .A1(n9746), .A2(n13754), .A3(n9745), .ZN(n9747) );
  XNOR2_X1 U12213 ( .A(n9747), .B(n11268), .ZN(n9749) );
  INV_X1 U12214 ( .A(n11088), .ZN(n9748) );
  INV_X1 U12215 ( .A(n13699), .ZN(n9757) );
  INV_X1 U12216 ( .A(n9752), .ZN(n9750) );
  NAND2_X1 U12217 ( .A1(n9757), .A2(n9750), .ZN(n9760) );
  XOR2_X1 U12218 ( .A(n9752), .B(n9751), .Z(n9753) );
  NAND3_X1 U12219 ( .A1(n9753), .A2(n14013), .A3(n13699), .ZN(n9759) );
  INV_X1 U12220 ( .A(n9754), .ZN(n9756) );
  NAND4_X1 U12221 ( .A1(n9761), .A2(n9757), .A3(n9756), .A4(n9755), .ZN(n9758)
         );
  OAI211_X1 U12222 ( .C1(n9761), .C2(n9760), .A(n9759), .B(n9758), .ZN(n9762)
         );
  INV_X1 U12223 ( .A(n9762), .ZN(n9763) );
  OAI21_X1 U12224 ( .B1(n9766), .B2(n9765), .A(n7341), .ZN(n9773) );
  INV_X1 U12225 ( .A(n9767), .ZN(n9769) );
  NAND2_X1 U12226 ( .A1(n9769), .A2(n9768), .ZN(n9775) );
  NAND2_X1 U12227 ( .A1(n9775), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9771) );
  INV_X1 U12228 ( .A(n10163), .ZN(n10108) );
  NAND2_X1 U12229 ( .A1(n10108), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10161) );
  OAI21_X1 U12230 ( .B1(n9774), .B2(n9773), .A(n9772), .ZN(n9787) );
  INV_X1 U12231 ( .A(n9775), .ZN(n9776) );
  NAND2_X1 U12232 ( .A1(n9776), .A2(n9770), .ZN(n9778) );
  OAI21_X2 U12233 ( .B1(n9778), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9777) );
  NAND2_X1 U12234 ( .A1(n6506), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9780) );
  MUX2_X1 U12235 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9780), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n9782) );
  NAND2_X1 U12236 ( .A1(n9782), .A2(n9781), .ZN(n14277) );
  NAND3_X2 U12237 ( .A1(n10103), .A2(n10102), .A3(n10311), .ZN(n10596) );
  OR2_X1 U12238 ( .A1(n10604), .A2(n10592), .ZN(n10735) );
  INV_X1 U12239 ( .A(n6588), .ZN(n10277) );
  INV_X1 U12240 ( .A(n10604), .ZN(n10164) );
  NAND3_X1 U12241 ( .A1(n10747), .A2(n10277), .A3(n13981), .ZN(n9785) );
  OAI211_X1 U12242 ( .C1(n9719), .C2(n10161), .A(n9785), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9786) );
  NAND2_X1 U12243 ( .A1(n9787), .A2(n9786), .ZN(P1_U3242) );
  OAI21_X1 U12244 ( .B1(n9884), .B2(n9886), .A(n9885), .ZN(n9788) );
  NAND2_X1 U12245 ( .A1(n9788), .A2(n11360), .ZN(n9790) );
  OAI21_X1 U12246 ( .B1(n10832), .B2(n9886), .A(n9884), .ZN(n9789) );
  NAND2_X1 U12247 ( .A1(n9790), .A2(n9789), .ZN(n10568) );
  AND2_X1 U12248 ( .A1(n15130), .A2(n9791), .ZN(n9792) );
  NAND2_X1 U12249 ( .A1(n10568), .A2(n9792), .ZN(n9794) );
  AND2_X1 U12250 ( .A1(n10984), .A2(n9886), .ZN(n9793) );
  NAND2_X1 U12251 ( .A1(n11339), .A2(n9793), .ZN(n9882) );
  INV_X1 U12252 ( .A(n9795), .ZN(n12564) );
  NOR2_X1 U12253 ( .A1(n12564), .A2(n9796), .ZN(n9798) );
  XNOR2_X1 U12254 ( .A(n9798), .B(n9797), .ZN(n12560) );
  NAND2_X1 U12255 ( .A1(n9800), .A2(n9799), .ZN(n10547) );
  NAND2_X1 U12256 ( .A1(n9801), .A2(n15073), .ZN(n15072) );
  NAND2_X1 U12257 ( .A1(n15072), .A2(n10558), .ZN(n15058) );
  NAND2_X1 U12258 ( .A1(n15058), .A2(n9803), .ZN(n15057) );
  NAND2_X1 U12259 ( .A1(n10776), .A2(n9804), .ZN(n10837) );
  AND2_X1 U12260 ( .A1(n9805), .A2(n10837), .ZN(n9806) );
  NAND2_X1 U12261 ( .A1(n15057), .A2(n9806), .ZN(n10840) );
  NAND2_X1 U12262 ( .A1(n12451), .A2(n10845), .ZN(n9807) );
  NAND2_X1 U12263 ( .A1(n10840), .A2(n9807), .ZN(n10824) );
  NAND2_X1 U12264 ( .A1(n10824), .A2(n9808), .ZN(n9810) );
  NAND2_X1 U12265 ( .A1(n12450), .A2(n11005), .ZN(n9809) );
  NAND2_X1 U12266 ( .A1(n11377), .A2(n11177), .ZN(n11196) );
  AND2_X1 U12267 ( .A1(n11198), .A2(n11196), .ZN(n9812) );
  NAND2_X1 U12268 ( .A1(n12448), .A2(n11521), .ZN(n9813) );
  NAND2_X1 U12269 ( .A1(n11197), .A2(n9813), .ZN(n11248) );
  NAND2_X1 U12270 ( .A1(n11248), .A2(n11387), .ZN(n9816) );
  NAND2_X1 U12271 ( .A1(n11562), .A2(n9814), .ZN(n9815) );
  NAND2_X1 U12272 ( .A1(n9816), .A2(n9815), .ZN(n11315) );
  INV_X1 U12273 ( .A(n11315), .ZN(n9818) );
  INV_X1 U12274 ( .A(n11317), .ZN(n9817) );
  NAND2_X1 U12275 ( .A1(n11566), .A2(n15131), .ZN(n9819) );
  NAND2_X1 U12276 ( .A1(n15027), .A2(n9822), .ZN(n9824) );
  INV_X1 U12277 ( .A(n15039), .ZN(n11946) );
  OR2_X1 U12278 ( .A1(n11946), .A2(n15033), .ZN(n9823) );
  INV_X1 U12279 ( .A(n11818), .ZN(n11822) );
  NAND2_X1 U12280 ( .A1(n11982), .A2(n14452), .ZN(n9825) );
  NAND2_X1 U12281 ( .A1(n11821), .A2(n9825), .ZN(n11867) );
  NAND2_X1 U12282 ( .A1(n11867), .A2(n11868), .ZN(n11866) );
  INV_X1 U12283 ( .A(n12870), .ZN(n12396) );
  NAND2_X1 U12284 ( .A1(n12396), .A2(n12446), .ZN(n9826) );
  NAND2_X1 U12285 ( .A1(n11866), .A2(n9826), .ZN(n11911) );
  INV_X1 U12286 ( .A(n12445), .ZN(n12739) );
  OR2_X1 U12287 ( .A1(n12866), .A2(n12739), .ZN(n9827) );
  NAND2_X1 U12288 ( .A1(n12862), .A2(n12357), .ZN(n12720) );
  AND2_X1 U12289 ( .A1(n12732), .A2(n12738), .ZN(n9830) );
  INV_X1 U12290 ( .A(n9830), .ZN(n9828) );
  AND2_X1 U12291 ( .A1(n12720), .A2(n9828), .ZN(n12704) );
  AND2_X1 U12292 ( .A1(n12704), .A2(n12708), .ZN(n9832) );
  INV_X1 U12293 ( .A(n12708), .ZN(n9831) );
  OR2_X1 U12294 ( .A1(n12862), .A2(n12357), .ZN(n12721) );
  AND2_X1 U12295 ( .A1(n12721), .A2(n7321), .ZN(n9829) );
  OR2_X1 U12296 ( .A1(n9830), .A2(n9829), .ZN(n12705) );
  INV_X1 U12297 ( .A(n12725), .ZN(n12693) );
  NOR2_X1 U12298 ( .A1(n12788), .A2(n12691), .ZN(n9835) );
  OAI22_X2 U12299 ( .A1(n12674), .A2(n9835), .B1(n12411), .B2(n12683), .ZN(
        n12662) );
  INV_X1 U12300 ( .A(n12608), .ZN(n9841) );
  NAND2_X1 U12301 ( .A1(n12567), .A2(n12568), .ZN(n12566) );
  NAND2_X1 U12302 ( .A1(n12829), .A2(n12422), .ZN(n9843) );
  AND2_X1 U12303 ( .A1(n12566), .A2(n9843), .ZN(n9846) );
  NAND2_X1 U12304 ( .A1(n12566), .A2(n9844), .ZN(n9898) );
  NAND2_X1 U12305 ( .A1(n11339), .A2(n9885), .ZN(n9868) );
  OAI211_X1 U12306 ( .C1(n9846), .C2(n9797), .A(n9898), .B(n15074), .ZN(n9848)
         );
  INV_X1 U12307 ( .A(n12422), .ZN(n12584) );
  NAND2_X1 U12308 ( .A1(n12584), .A2(n15076), .ZN(n9847) );
  OAI211_X1 U12309 ( .C1(n12327), .C2(n15059), .A(n9848), .B(n9847), .ZN(
        n12555) );
  AOI21_X1 U12310 ( .B1(n15099), .B2(n12560), .A(n12555), .ZN(n9892) );
  XNOR2_X1 U12311 ( .A(n9849), .B(P3_B_REG_SCAN_IN), .ZN(n9850) );
  NAND2_X1 U12312 ( .A1(n9850), .A2(n11908), .ZN(n9852) );
  NAND2_X1 U12313 ( .A1(n9852), .A2(n9851), .ZN(n9855) );
  OR2_X1 U12314 ( .A1(n9855), .A2(P3_D_REG_1__SCAN_IN), .ZN(n9854) );
  NAND2_X1 U12315 ( .A1(n11908), .A2(n11955), .ZN(n9853) );
  NAND2_X1 U12316 ( .A1(n9849), .A2(n11955), .ZN(n9856) );
  INV_X1 U12317 ( .A(n9881), .ZN(n9867) );
  NOR2_X1 U12318 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_7__SCAN_IN), .ZN(
        n14185) );
  NOR4_X1 U12319 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_22__SCAN_IN), .A4(P3_D_REG_17__SCAN_IN), .ZN(n9859) );
  NOR4_X1 U12320 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_24__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_10__SCAN_IN), .ZN(n9858) );
  NOR4_X1 U12321 ( .A1(P3_D_REG_25__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n9857) );
  NAND4_X1 U12322 ( .A1(n14185), .A2(n9859), .A3(n9858), .A4(n9857), .ZN(n9865) );
  NOR4_X1 U12323 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_9__SCAN_IN), .A3(
        P3_D_REG_16__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n9863) );
  NOR4_X1 U12324 ( .A1(P3_D_REG_14__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_26__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n9862) );
  NOR4_X1 U12325 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_4__SCAN_IN), .ZN(n9861) );
  NOR4_X1 U12326 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_23__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n9860) );
  NAND4_X1 U12327 ( .A1(n9863), .A2(n9862), .A3(n9861), .A4(n9860), .ZN(n9864)
         );
  NOR2_X1 U12328 ( .A1(n9865), .A2(n9864), .ZN(n9866) );
  NAND2_X1 U12329 ( .A1(n9867), .A2(n9878), .ZN(n10572) );
  OR2_X1 U12330 ( .A1(n9868), .A2(n10554), .ZN(n10569) );
  AND2_X1 U12331 ( .A1(n10499), .A2(n10569), .ZN(n9871) );
  NAND2_X1 U12332 ( .A1(n10813), .A2(n10553), .ZN(n9880) );
  INV_X1 U12333 ( .A(n9878), .ZN(n9869) );
  INV_X1 U12334 ( .A(n10568), .ZN(n9870) );
  OAI22_X1 U12335 ( .A1(n10572), .A2(n9871), .B1(n10570), .B2(n9870), .ZN(
        n9872) );
  OR2_X1 U12336 ( .A1(n9892), .A2(n15144), .ZN(n9877) );
  INV_X1 U12337 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n9873) );
  OR2_X1 U12338 ( .A1(n15146), .A2(n9873), .ZN(n9874) );
  INV_X1 U12339 ( .A(n9875), .ZN(n9876) );
  NAND2_X1 U12340 ( .A1(n9877), .A2(n9876), .ZN(P3_U3455) );
  AND2_X1 U12341 ( .A1(n9878), .A2(n10573), .ZN(n9879) );
  NAND2_X1 U12342 ( .A1(n9887), .A2(n9888), .ZN(n10536) );
  NAND2_X1 U12343 ( .A1(n9883), .A2(n9882), .ZN(n10812) );
  AND2_X1 U12344 ( .A1(n10536), .A2(n10812), .ZN(n10814) );
  OAI22_X1 U12345 ( .A1(n15130), .A2(n9886), .B1(n9885), .B2(n9884), .ZN(n9889) );
  AOI21_X1 U12346 ( .B1(n9889), .B2(n9888), .A(n9887), .ZN(n9890) );
  MUX2_X1 U12347 ( .A(n10814), .B(n9890), .S(n10813), .Z(n9891) );
  OR2_X1 U12348 ( .A1(n9892), .A2(n15163), .ZN(n9897) );
  NOR2_X1 U12349 ( .A1(n15166), .A2(n9893), .ZN(n9894) );
  NAND2_X1 U12350 ( .A1(n9897), .A2(n9896), .ZN(P3_U3487) );
  NAND2_X1 U12351 ( .A1(n9898), .A2(n7340), .ZN(n9899) );
  XNOR2_X1 U12352 ( .A(n9899), .B(n9907), .ZN(n9905) );
  INV_X1 U12353 ( .A(P3_B_REG_SCAN_IN), .ZN(n9900) );
  OAI21_X1 U12354 ( .B1(n12029), .B2(n9900), .A(n15079), .ZN(n12539) );
  NOR2_X1 U12355 ( .A1(n9901), .A2(n12539), .ZN(n9902) );
  XOR2_X1 U12356 ( .A(n9907), .B(n9906), .Z(n12546) );
  AND2_X1 U12357 ( .A1(n12546), .A2(n15099), .ZN(n9908) );
  NOR2_X1 U12358 ( .A1(n12547), .A2(n9908), .ZN(n9912) );
  MUX2_X1 U12359 ( .A(n9909), .B(n9912), .S(n15166), .Z(n9911) );
  NAND2_X1 U12360 ( .A1(n9911), .A2(n7322), .ZN(P3_U3488) );
  INV_X1 U12361 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9913) );
  MUX2_X1 U12362 ( .A(n9913), .B(n9912), .S(n15146), .Z(n9914) );
  NAND2_X1 U12363 ( .A1(n9914), .A2(n7323), .ZN(P3_U3456) );
  INV_X1 U12364 ( .A(n9915), .ZN(n9916) );
  INV_X1 U12365 ( .A(n6429), .ZN(n9957) );
  NAND2_X1 U12366 ( .A1(n9957), .A2(n10694), .ZN(n9917) );
  NAND2_X1 U12367 ( .A1(n10479), .A2(n9917), .ZN(n10612) );
  NAND2_X1 U12368 ( .A1(n8272), .A2(n10956), .ZN(n9918) );
  NAND2_X1 U12369 ( .A1(n10610), .A2(n9918), .ZN(n10703) );
  NAND2_X1 U12370 ( .A1(n10703), .A2(n10702), .ZN(n10701) );
  INV_X1 U12371 ( .A(n13028), .ZN(n10660) );
  NAND2_X1 U12372 ( .A1(n10660), .A2(n11018), .ZN(n9919) );
  NAND2_X1 U12373 ( .A1(n10701), .A2(n9919), .ZN(n10755) );
  INV_X1 U12374 ( .A(n13027), .ZN(n10408) );
  NAND2_X1 U12375 ( .A1(n10408), .A2(n10887), .ZN(n9920) );
  NAND2_X1 U12376 ( .A1(n10754), .A2(n9920), .ZN(n10860) );
  INV_X1 U12377 ( .A(n10863), .ZN(n10859) );
  NAND2_X1 U12378 ( .A1(n10860), .A2(n10859), .ZN(n10858) );
  INV_X1 U12379 ( .A(n13026), .ZN(n9966) );
  NAND2_X1 U12380 ( .A1(n6758), .A2(n9966), .ZN(n9921) );
  NAND2_X1 U12381 ( .A1(n10858), .A2(n9921), .ZN(n10972) );
  INV_X1 U12382 ( .A(n9969), .ZN(n10974) );
  OR2_X1 U12383 ( .A1(n11096), .A2(n13025), .ZN(n9922) );
  NAND2_X1 U12384 ( .A1(n10971), .A2(n9922), .ZN(n11158) );
  INV_X1 U12385 ( .A(n11162), .ZN(n11157) );
  OR2_X1 U12386 ( .A1(n11168), .A2(n13024), .ZN(n9923) );
  INV_X1 U12387 ( .A(n11231), .ZN(n11226) );
  NAND2_X1 U12388 ( .A1(n14881), .A2(n13023), .ZN(n9924) );
  NAND2_X1 U12389 ( .A1(n11325), .A2(n11327), .ZN(n9926) );
  NAND2_X1 U12390 ( .A1(n11543), .A2(n13022), .ZN(n9925) );
  NAND2_X1 U12391 ( .A1(n9926), .A2(n9925), .ZN(n11490) );
  NAND2_X1 U12392 ( .A1(n11490), .A2(n11491), .ZN(n9928) );
  NAND2_X1 U12393 ( .A1(n11500), .A2(n13021), .ZN(n9927) );
  NAND2_X1 U12394 ( .A1(n9928), .A2(n9927), .ZN(n11621) );
  AND2_X1 U12395 ( .A1(n12208), .A2(n13020), .ZN(n9930) );
  OR2_X1 U12396 ( .A1(n12208), .A2(n13020), .ZN(n9929) );
  OR2_X1 U12397 ( .A1(n11643), .A2(n13019), .ZN(n9931) );
  NOR2_X1 U12398 ( .A1(n11666), .A2(n13018), .ZN(n9932) );
  NAND2_X1 U12399 ( .A1(n11666), .A2(n13018), .ZN(n9933) );
  INV_X1 U12400 ( .A(n11893), .ZN(n11902) );
  OR2_X1 U12401 ( .A1(n11860), .A2(n13016), .ZN(n9936) );
  INV_X1 U12402 ( .A(n13266), .ZN(n13258) );
  OR2_X1 U12403 ( .A1(n13359), .A2(n13013), .ZN(n9939) );
  NAND2_X1 U12404 ( .A1(n13229), .A2(n13012), .ZN(n9940) );
  AND2_X1 U12405 ( .A1(n13406), .A2(n13011), .ZN(n9941) );
  INV_X1 U12406 ( .A(n13181), .ZN(n13184) );
  OR2_X1 U12407 ( .A1(n13192), .A2(n12896), .ZN(n9942) );
  NOR2_X1 U12408 ( .A1(n13394), .A2(n12979), .ZN(n9945) );
  NAND2_X1 U12409 ( .A1(n13129), .A2(n12888), .ZN(n9947) );
  XNOR2_X1 U12410 ( .A(n9949), .B(n10006), .ZN(n13302) );
  NOR2_X1 U12411 ( .A1(n9950), .A2(n10490), .ZN(n9951) );
  NAND2_X1 U12412 ( .A1(n10290), .A2(n9952), .ZN(n9953) );
  NAND2_X1 U12413 ( .A1(n9955), .A2(n8022), .ZN(n11238) );
  NAND2_X1 U12414 ( .A1(n9954), .A2(n11238), .ZN(n9956) );
  INV_X1 U12415 ( .A(n13150), .ZN(n13155) );
  NAND2_X1 U12416 ( .A1(n9957), .A2(n10967), .ZN(n9958) );
  NAND2_X1 U12417 ( .A1(n10617), .A2(n10616), .ZN(n9960) );
  NAND2_X1 U12418 ( .A1(n8272), .A2(n10622), .ZN(n9959) );
  INV_X1 U12419 ( .A(n10702), .ZN(n10706) );
  NAND2_X1 U12420 ( .A1(n10705), .A2(n10706), .ZN(n9962) );
  NAND2_X1 U12421 ( .A1(n10660), .A2(n10712), .ZN(n9961) );
  INV_X1 U12422 ( .A(n10757), .ZN(n9963) );
  NAND2_X1 U12423 ( .A1(n10408), .A2(n10761), .ZN(n9964) );
  NAND2_X1 U12424 ( .A1(n9965), .A2(n9964), .ZN(n10864) );
  NAND2_X1 U12425 ( .A1(n10864), .A2(n10863), .ZN(n9968) );
  NAND2_X1 U12426 ( .A1(n12171), .A2(n9966), .ZN(n9967) );
  INV_X1 U12427 ( .A(n13025), .ZN(n9970) );
  NAND2_X1 U12428 ( .A1(n11096), .A2(n9970), .ZN(n9971) );
  INV_X1 U12429 ( .A(n13024), .ZN(n12215) );
  AND2_X1 U12430 ( .A1(n11168), .A2(n12215), .ZN(n9972) );
  OR2_X1 U12431 ( .A1(n14881), .A2(n11144), .ZN(n9973) );
  NAND2_X1 U12432 ( .A1(n9974), .A2(n9973), .ZN(n11326) );
  INV_X1 U12433 ( .A(n11327), .ZN(n9975) );
  NAND2_X1 U12434 ( .A1(n11326), .A2(n9975), .ZN(n9978) );
  OR2_X1 U12435 ( .A1(n11543), .A2(n9976), .ZN(n9977) );
  NAND2_X1 U12436 ( .A1(n9978), .A2(n9977), .ZN(n11492) );
  INV_X1 U12437 ( .A(n11491), .ZN(n11489) );
  OR2_X1 U12438 ( .A1(n11500), .A2(n12200), .ZN(n9979) );
  INV_X1 U12439 ( .A(n11620), .ZN(n11619) );
  INV_X1 U12440 ( .A(n13020), .ZN(n9980) );
  NAND2_X1 U12441 ( .A1(n12208), .A2(n9980), .ZN(n11637) );
  AND2_X1 U12442 ( .A1(n11636), .A2(n11637), .ZN(n9981) );
  NAND2_X1 U12443 ( .A1(n11616), .A2(n9981), .ZN(n11635) );
  NAND2_X1 U12444 ( .A1(n11745), .A2(n11748), .ZN(n9984) );
  INV_X1 U12445 ( .A(n13018), .ZN(n12189) );
  OR2_X1 U12446 ( .A1(n11666), .A2(n12189), .ZN(n9983) );
  NAND2_X2 U12447 ( .A1(n9984), .A2(n9983), .ZN(n14473) );
  NAND2_X1 U12448 ( .A1(n14473), .A2(n13017), .ZN(n9985) );
  INV_X1 U12449 ( .A(n13017), .ZN(n9986) );
  OR2_X1 U12450 ( .A1(n11860), .A2(n12188), .ZN(n9988) );
  INV_X1 U12451 ( .A(n13276), .ZN(n9990) );
  NAND2_X1 U12452 ( .A1(n9990), .A2(n9989), .ZN(n13274) );
  NAND2_X1 U12453 ( .A1(n13285), .A2(n11961), .ZN(n9991) );
  NAND2_X1 U12454 ( .A1(n13416), .A2(n13014), .ZN(n9992) );
  INV_X1 U12455 ( .A(n13242), .ZN(n9994) );
  INV_X1 U12456 ( .A(n13013), .ZN(n9993) );
  AOI21_X2 U12457 ( .B1(n9994), .B2(n7320), .A(n7319), .ZN(n13236) );
  INV_X1 U12458 ( .A(n13235), .ZN(n13225) );
  INV_X1 U12459 ( .A(n13012), .ZN(n12969) );
  OR2_X1 U12460 ( .A1(n13229), .A2(n12969), .ZN(n9995) );
  INV_X1 U12461 ( .A(n13209), .ZN(n13212) );
  NAND2_X1 U12462 ( .A1(n13406), .A2(n9996), .ZN(n9997) );
  OR2_X1 U12463 ( .A1(n13344), .A2(n12958), .ZN(n9998) );
  AND2_X1 U12464 ( .A1(n13192), .A2(n13009), .ZN(n9999) );
  NAND2_X1 U12465 ( .A1(n13174), .A2(n13008), .ZN(n10000) );
  INV_X1 U12466 ( .A(n13138), .ZN(n13135) );
  INV_X1 U12467 ( .A(n10002), .ZN(n10003) );
  INV_X1 U12468 ( .A(n13090), .ZN(n13093) );
  NAND2_X1 U12469 ( .A1(n13116), .A2(n12985), .ZN(n13094) );
  NAND3_X1 U12470 ( .A1(n13108), .A2(n13093), .A3(n13094), .ZN(n13092) );
  NAND2_X1 U12471 ( .A1(n13092), .A2(n10005), .ZN(n10008) );
  XNOR2_X1 U12472 ( .A(n10008), .B(n10007), .ZN(n10017) );
  NAND2_X1 U12473 ( .A1(n10009), .A2(n8022), .ZN(n10011) );
  NAND2_X1 U12474 ( .A1(n13003), .A2(n12986), .ZN(n10015) );
  NOR2_X1 U12475 ( .A1(n12024), .A2(n10012), .ZN(n10013) );
  NOR2_X1 U12476 ( .A1(n12984), .A2(n10013), .ZN(n13078) );
  INV_X2 U12477 ( .A(n14868), .ZN(n14478) );
  INV_X1 U12478 ( .A(n12208), .ZN(n11729) );
  INV_X1 U12479 ( .A(n11500), .ZN(n14890) );
  NAND2_X1 U12480 ( .A1(n10704), .A2(n11018), .ZN(n10756) );
  NOR2_X2 U12481 ( .A1(n11543), .A2(n11331), .ZN(n11497) );
  NAND2_X1 U12482 ( .A1(n14493), .A2(n14484), .ZN(n13284) );
  OR2_X2 U12483 ( .A1(n13285), .A2(n13284), .ZN(n13286) );
  INV_X1 U12484 ( .A(n13102), .ZN(n10021) );
  AOI211_X1 U12485 ( .C1(n8282), .C2(n10021), .A(n7779), .B(n13082), .ZN(
        n13299) );
  INV_X1 U12486 ( .A(n10022), .ZN(n10023) );
  INV_X1 U12487 ( .A(n10024), .ZN(n10025) );
  INV_X1 U12488 ( .A(n14863), .ZN(n14849) );
  AOI22_X1 U12489 ( .A1(n10025), .A2(n14849), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n14478), .ZN(n10026) );
  OAI21_X1 U12490 ( .B1(n10027), .B2(n14853), .A(n10026), .ZN(n10028) );
  NAND2_X1 U12491 ( .A1(n10112), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10032) );
  INV_X1 U12492 ( .A(n10033), .ZN(n10034) );
  NOR2_X1 U12493 ( .A1(n10049), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12872) );
  INV_X2 U12494 ( .A(n12872), .ZN(n12880) );
  OAI222_X1 U12495 ( .A1(n12880), .A2(n10037), .B1(n12040), .B2(n10036), .C1(
        n10035), .C2(P3_U3151), .ZN(P3_U3289) );
  INV_X1 U12496 ( .A(n10038), .ZN(n10041) );
  INV_X1 U12497 ( .A(SI_5_), .ZN(n10040) );
  OAI222_X1 U12498 ( .A1(n12880), .A2(n10041), .B1(n12040), .B2(n10040), .C1(
        n10039), .C2(P3_U3151), .ZN(P3_U3290) );
  INV_X1 U12499 ( .A(n10042), .ZN(n10044) );
  INV_X1 U12500 ( .A(SI_2_), .ZN(n10043) );
  OAI222_X1 U12501 ( .A1(n9121), .A2(P3_U3151), .B1(n12880), .B2(n10044), .C1(
        n10043), .C2(n12040), .ZN(P3_U3293) );
  INV_X1 U12502 ( .A(n10045), .ZN(n10047) );
  INV_X1 U12503 ( .A(SI_7_), .ZN(n10046) );
  OAI222_X1 U12504 ( .A1(n10799), .A2(P3_U3151), .B1(n12880), .B2(n10047), 
        .C1(n10046), .C2(n12040), .ZN(P3_U3288) );
  NAND2_X2 U12505 ( .A1(n10049), .A2(P2_U3088), .ZN(n13438) );
  AOI22_X1 U12506 ( .A1(n13433), .A2(P1_DATAO_REG_1__SCAN_IN), .B1(
        P2_STATE_REG_SCAN_IN), .B2(n14749), .ZN(n10048) );
  OAI21_X1 U12507 ( .B1(n10050), .B2(n13438), .A(n10048), .ZN(P2_U3326) );
  NAND2_X2 U12508 ( .A1(n10049), .A2(P1_U3086), .ZN(n14278) );
  NOR2_X1 U12509 ( .A1(n10049), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14267) );
  INV_X2 U12510 ( .A(n14267), .ZN(n14281) );
  OAI222_X1 U12511 ( .A1(n14278), .A2(n7367), .B1(n14281), .B2(n10050), .C1(
        P1_U3086), .C2(n13577), .ZN(P1_U3354) );
  INV_X1 U12512 ( .A(SI_3_), .ZN(n10053) );
  INV_X1 U12513 ( .A(n10051), .ZN(n10052) );
  OAI222_X1 U12514 ( .A1(P3_U3151), .A2(n10054), .B1(n12040), .B2(n10053), 
        .C1(n12880), .C2(n10052), .ZN(P3_U3292) );
  INV_X1 U12515 ( .A(n10055), .ZN(n10057) );
  INV_X1 U12516 ( .A(SI_4_), .ZN(n10056) );
  OAI222_X1 U12517 ( .A1(n12880), .A2(n10057), .B1(n12040), .B2(n10056), .C1(
        n10478), .C2(P3_U3151), .ZN(P3_U3291) );
  INV_X1 U12518 ( .A(n13607), .ZN(n10059) );
  INV_X1 U12519 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10058) );
  OAI222_X1 U12520 ( .A1(P1_U3086), .A2(n10059), .B1(n14281), .B2(n10077), 
        .C1(n10058), .C2(n14278), .ZN(P1_U3352) );
  OAI222_X1 U12521 ( .A1(P1_U3086), .A2(n13598), .B1(n14281), .B2(n10082), 
        .C1(n10060), .C2(n14278), .ZN(P1_U3353) );
  OAI222_X1 U12522 ( .A1(P1_U3086), .A2(n6613), .B1(n14281), .B2(n10080), .C1(
        n10061), .C2(n14278), .ZN(P1_U3350) );
  INV_X1 U12523 ( .A(n14579), .ZN(n10064) );
  INV_X1 U12524 ( .A(n10062), .ZN(n10085) );
  OAI222_X1 U12525 ( .A1(P1_U3086), .A2(n10064), .B1(n14281), .B2(n10085), 
        .C1(n10063), .C2(n14278), .ZN(P1_U3351) );
  OAI222_X1 U12526 ( .A1(P3_U3151), .A2(n10066), .B1(n12040), .B2(n7369), .C1(
        n12880), .C2(n10065), .ZN(P3_U3294) );
  OAI222_X1 U12527 ( .A1(n10993), .A2(P3_U3151), .B1(n12880), .B2(n10068), 
        .C1(n10067), .C2(n12040), .ZN(P3_U3287) );
  OAI222_X1 U12528 ( .A1(n10071), .A2(P3_U3151), .B1(n12880), .B2(n10070), 
        .C1(n10069), .C2(n12040), .ZN(P3_U3286) );
  OAI222_X1 U12529 ( .A1(n12880), .A2(n10073), .B1(n12040), .B2(n10072), .C1(
        n14973), .C2(P3_U3151), .ZN(P3_U3285) );
  INV_X1 U12530 ( .A(n10414), .ZN(n10419) );
  OAI222_X1 U12531 ( .A1(P1_U3086), .A2(n10419), .B1(n14281), .B2(n10075), 
        .C1(n10074), .C2(n14278), .ZN(P1_U3349) );
  INV_X1 U12532 ( .A(n10182), .ZN(n14774) );
  INV_X2 U12533 ( .A(n13433), .ZN(n13440) );
  OAI222_X1 U12534 ( .A1(n13438), .A2(n10075), .B1(n14774), .B2(P2_U3088), 
        .C1(n7139), .C2(n13440), .ZN(P2_U3321) );
  OAI222_X1 U12535 ( .A1(n13438), .A2(n10077), .B1(n10172), .B2(P2_U3088), 
        .C1(n10076), .C2(n13440), .ZN(P2_U3324) );
  INV_X1 U12536 ( .A(n13036), .ZN(n10079) );
  OAI222_X1 U12537 ( .A1(n13438), .A2(n10080), .B1(n10079), .B2(P2_U3088), 
        .C1(n10078), .C2(n13440), .ZN(P2_U3322) );
  INV_X1 U12538 ( .A(n10143), .ZN(n10157) );
  OAI222_X1 U12539 ( .A1(n13438), .A2(n10082), .B1(n10157), .B2(P2_U3088), 
        .C1(n10081), .C2(n13440), .ZN(P2_U3325) );
  INV_X1 U12540 ( .A(n14763), .ZN(n10084) );
  OAI222_X1 U12541 ( .A1(n13438), .A2(n10085), .B1(n10084), .B2(P2_U3088), 
        .C1(n10083), .C2(n13440), .ZN(P2_U3323) );
  NAND2_X1 U12542 ( .A1(n10208), .A2(P3_D_REG_0__SCAN_IN), .ZN(n10086) );
  OAI21_X1 U12543 ( .B1(n10553), .B2(n10208), .A(n10086), .ZN(P3_U3376) );
  NAND2_X1 U12544 ( .A1(n10208), .A2(P3_D_REG_1__SCAN_IN), .ZN(n10087) );
  OAI21_X1 U12545 ( .B1(n10813), .B2(n10208), .A(n10087), .ZN(P3_U3377) );
  OAI222_X1 U12546 ( .A1(n12880), .A2(n10089), .B1(n12040), .B2(n10088), .C1(
        n14989), .C2(P3_U3151), .ZN(P3_U3284) );
  INV_X1 U12547 ( .A(n13052), .ZN(n10091) );
  OAI222_X1 U12548 ( .A1(n13438), .A2(n10093), .B1(n10091), .B2(P2_U3088), 
        .C1(n10090), .C2(n13440), .ZN(P2_U3320) );
  INV_X1 U12549 ( .A(n13638), .ZN(n10330) );
  OAI222_X1 U12550 ( .A1(P1_U3086), .A2(n10330), .B1(n14281), .B2(n10093), 
        .C1(n10092), .C2(n14278), .ZN(P1_U3348) );
  INV_X1 U12551 ( .A(n10188), .ZN(n10251) );
  OAI222_X1 U12552 ( .A1(n13438), .A2(n10096), .B1(n10251), .B2(P2_U3088), 
        .C1(n10094), .C2(n13440), .ZN(P2_U3319) );
  INV_X1 U12553 ( .A(n10372), .ZN(n10097) );
  OAI222_X1 U12554 ( .A1(P1_U3086), .A2(n10097), .B1(n14281), .B2(n10096), 
        .C1(n10095), .C2(n14278), .ZN(P1_U3347) );
  INV_X1 U12555 ( .A(n10098), .ZN(n10101) );
  INV_X1 U12556 ( .A(SI_12_), .ZN(n10099) );
  OAI222_X1 U12557 ( .A1(n12880), .A2(n10101), .B1(n10100), .B2(P3_U3151), 
        .C1(n10099), .C2(n12040), .ZN(P3_U3283) );
  INV_X1 U12558 ( .A(n10102), .ZN(n12020) );
  NAND2_X1 U12559 ( .A1(n12020), .A2(P1_B_REG_SCAN_IN), .ZN(n10104) );
  OR2_X1 U12560 ( .A1(n10104), .A2(n10103), .ZN(n10106) );
  INV_X1 U12561 ( .A(P1_B_REG_SCAN_IN), .ZN(n13697) );
  AOI21_X1 U12562 ( .B1(n10102), .B2(n13697), .A(n14277), .ZN(n10105) );
  INV_X1 U12563 ( .A(n10310), .ZN(n10107) );
  INV_X1 U12564 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10308) );
  NOR3_X1 U12565 ( .A1(n10108), .A2(n10311), .A3(P1_U3086), .ZN(n10109) );
  AOI22_X1 U12566 ( .A1(n14651), .A2(n10308), .B1(n10109), .B2(n12020), .ZN(
        P1_U3445) );
  INV_X1 U12567 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10309) );
  INV_X1 U12568 ( .A(n10103), .ZN(n14282) );
  AOI22_X1 U12569 ( .A1(n14651), .A2(n10309), .B1(n10109), .B2(n14282), .ZN(
        P1_U3446) );
  INV_X1 U12570 ( .A(n10110), .ZN(n10159) );
  INV_X1 U12571 ( .A(n14278), .ZN(n12036) );
  AOI22_X1 U12572 ( .A1(n13656), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n12036), .ZN(n10111) );
  OAI21_X1 U12573 ( .B1(n10159), .B2(n14281), .A(n10111), .ZN(P1_U3346) );
  INV_X1 U12574 ( .A(n10112), .ZN(n10117) );
  NAND2_X1 U12575 ( .A1(n10113), .A2(n10112), .ZN(n10115) );
  NAND2_X1 U12576 ( .A1(n10115), .A2(n10114), .ZN(n10116) );
  OAI21_X1 U12577 ( .B1(n10118), .B2(n10117), .A(n10116), .ZN(n10133) );
  AND2_X1 U12578 ( .A1(n10133), .A2(n8032), .ZN(n14746) );
  INV_X1 U12579 ( .A(n14845), .ZN(n14818) );
  NOR2_X1 U12580 ( .A1(n8032), .A2(P2_U3088), .ZN(n13429) );
  AND2_X1 U12581 ( .A1(n13429), .A2(n12024), .ZN(n10119) );
  NAND2_X1 U12582 ( .A1(n10133), .A2(n10119), .ZN(n14836) );
  INV_X1 U12583 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10144) );
  MUX2_X1 U12584 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n10144), .S(n10143), .Z(
        n10122) );
  INV_X1 U12585 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10120) );
  MUX2_X1 U12586 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n10120), .S(n14749), .Z(
        n14755) );
  AND2_X1 U12587 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n14756) );
  NAND2_X1 U12588 ( .A1(n14755), .A2(n14756), .ZN(n14754) );
  NAND2_X1 U12589 ( .A1(n14749), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10145) );
  NAND2_X1 U12590 ( .A1(n14754), .A2(n10145), .ZN(n10121) );
  NAND2_X1 U12591 ( .A1(n10122), .A2(n10121), .ZN(n10148) );
  NAND2_X1 U12592 ( .A1(n10143), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10126) );
  NAND2_X1 U12593 ( .A1(n10148), .A2(n10126), .ZN(n10125) );
  INV_X1 U12594 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10123) );
  MUX2_X1 U12595 ( .A(n10123), .B(P2_REG1_REG_3__SCAN_IN), .S(n10172), .Z(
        n10124) );
  NAND2_X1 U12596 ( .A1(n10125), .A2(n10124), .ZN(n10175) );
  MUX2_X1 U12597 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n10123), .S(n10172), .Z(
        n10127) );
  NAND3_X1 U12598 ( .A1(n10127), .A2(n10148), .A3(n10126), .ZN(n10128) );
  NAND2_X1 U12599 ( .A1(n10175), .A2(n10128), .ZN(n10130) );
  OAI22_X1 U12600 ( .A1(n14836), .A2(n10130), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10129), .ZN(n10141) );
  INV_X1 U12601 ( .A(n12024), .ZN(n10131) );
  AND2_X1 U12602 ( .A1(n13429), .A2(n10131), .ZN(n10132) );
  INV_X1 U12603 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10134) );
  MUX2_X1 U12604 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n10134), .S(n14749), .Z(
        n14752) );
  NAND3_X1 U12605 ( .A1(n14752), .A2(P2_REG2_REG_0__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n14751) );
  NAND2_X1 U12606 ( .A1(n14749), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10150) );
  MUX2_X1 U12607 ( .A(n7414), .B(P2_REG2_REG_2__SCAN_IN), .S(n10143), .Z(
        n10151) );
  AOI21_X1 U12608 ( .B1(n14751), .B2(n10150), .A(n10151), .ZN(n10153) );
  NOR2_X1 U12609 ( .A1(n10157), .A2(n7414), .ZN(n10137) );
  INV_X1 U12610 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10135) );
  MUX2_X1 U12611 ( .A(n10135), .B(P2_REG2_REG_3__SCAN_IN), .S(n10172), .Z(
        n10136) );
  OAI21_X1 U12612 ( .B1(n10153), .B2(n10137), .A(n10136), .ZN(n10166) );
  INV_X1 U12613 ( .A(n10166), .ZN(n10139) );
  NOR3_X1 U12614 ( .A1(n10153), .A2(n10137), .A3(n10136), .ZN(n10138) );
  NOR3_X1 U12615 ( .A1(n14838), .A2(n10139), .A3(n10138), .ZN(n10140) );
  AOI211_X1 U12616 ( .C1(n14818), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n10141), .B(
        n10140), .ZN(n10142) );
  OAI21_X1 U12617 ( .B1(n10172), .B2(n10396), .A(n10142), .ZN(P2_U3217) );
  MUX2_X1 U12618 ( .A(n10144), .B(P2_REG1_REG_2__SCAN_IN), .S(n10143), .Z(
        n10146) );
  NAND3_X1 U12619 ( .A1(n10146), .A2(n14754), .A3(n10145), .ZN(n10147) );
  NAND2_X1 U12620 ( .A1(n10148), .A2(n10147), .ZN(n10149) );
  INV_X1 U12621 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10955) );
  OAI22_X1 U12622 ( .A1(n14836), .A2(n10149), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10955), .ZN(n10155) );
  AND3_X1 U12623 ( .A1(n10151), .A2(n14751), .A3(n10150), .ZN(n10152) );
  NOR3_X1 U12624 ( .A1(n14838), .A2(n10153), .A3(n10152), .ZN(n10154) );
  AOI211_X1 U12625 ( .C1(n14818), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n10155), .B(
        n10154), .ZN(n10156) );
  OAI21_X1 U12626 ( .B1(n10157), .B2(n10396), .A(n10156), .ZN(P2_U3216) );
  AOI22_X1 U12627 ( .A1(n10426), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n12036), .ZN(n10158) );
  OAI21_X1 U12628 ( .B1(n10207), .B2(n14281), .A(n10158), .ZN(P1_U3345) );
  INV_X1 U12629 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10160) );
  INV_X1 U12630 ( .A(n10266), .ZN(n10204) );
  OAI222_X1 U12631 ( .A1(n13440), .A2(n10160), .B1(n13438), .B2(n10159), .C1(
        P2_U3088), .C2(n10204), .ZN(P2_U3318) );
  INV_X1 U12632 ( .A(n10275), .ZN(n10165) );
  AOI21_X1 U12633 ( .B1(n10164), .B2(n10163), .A(n10162), .ZN(n10274) );
  NOR2_X2 U12634 ( .A1(n10165), .A2(n10274), .ZN(n14578) );
  NOR2_X1 U12635 ( .A1(n14578), .A2(P1_U4016), .ZN(P1_U3085) );
  OAI21_X1 U12636 ( .B1(n10135), .B2(n10172), .A(n10166), .ZN(n14766) );
  INV_X1 U12637 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10884) );
  MUX2_X1 U12638 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10884), .S(n14763), .Z(
        n14765) );
  NAND2_X1 U12639 ( .A1(n14766), .A2(n14765), .ZN(n14764) );
  NAND2_X1 U12640 ( .A1(n14763), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n13032) );
  INV_X1 U12641 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10167) );
  MUX2_X1 U12642 ( .A(n10167), .B(P2_REG2_REG_5__SCAN_IN), .S(n13036), .Z(
        n13031) );
  AOI21_X1 U12643 ( .B1(n14764), .B2(n13032), .A(n13031), .ZN(n13034) );
  AOI21_X1 U12644 ( .B1(n13036), .B2(P2_REG2_REG_5__SCAN_IN), .A(n13034), .ZN(
        n14782) );
  INV_X1 U12645 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10168) );
  MUX2_X1 U12646 ( .A(n10168), .B(P2_REG2_REG_6__SCAN_IN), .S(n10182), .Z(
        n14781) );
  NOR2_X1 U12647 ( .A1(n14782), .A2(n14781), .ZN(n14780) );
  NOR2_X1 U12648 ( .A1(n14774), .A2(n10168), .ZN(n13047) );
  INV_X1 U12649 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10169) );
  MUX2_X1 U12650 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10169), .S(n13052), .Z(
        n10170) );
  OAI21_X1 U12651 ( .B1(n14780), .B2(n13047), .A(n10170), .ZN(n13050) );
  NAND2_X1 U12652 ( .A1(n13052), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10241) );
  INV_X1 U12653 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10171) );
  MUX2_X1 U12654 ( .A(n10171), .B(P2_REG2_REG_8__SCAN_IN), .S(n10188), .Z(
        n10240) );
  AOI21_X1 U12655 ( .B1(n13050), .B2(n10241), .A(n10240), .ZN(n10239) );
  AOI21_X1 U12656 ( .B1(n10188), .B2(P2_REG2_REG_8__SCAN_IN), .A(n10239), .ZN(
        n10194) );
  INV_X1 U12657 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10192) );
  NOR3_X1 U12658 ( .A1(n10194), .A2(n10192), .A3(n14838), .ZN(n10191) );
  INV_X1 U12659 ( .A(n10172), .ZN(n10173) );
  NAND2_X1 U12660 ( .A1(n10173), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10174) );
  NAND2_X1 U12661 ( .A1(n10175), .A2(n10174), .ZN(n14769) );
  INV_X1 U12662 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10176) );
  MUX2_X1 U12663 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10176), .S(n14763), .Z(
        n14768) );
  NAND2_X1 U12664 ( .A1(n14769), .A2(n14768), .ZN(n14767) );
  NAND2_X1 U12665 ( .A1(n14763), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n13038) );
  NAND2_X1 U12666 ( .A1(n14767), .A2(n13038), .ZN(n10179) );
  INV_X1 U12667 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10177) );
  MUX2_X1 U12668 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n10177), .S(n13036), .Z(
        n10178) );
  NAND2_X1 U12669 ( .A1(n10179), .A2(n10178), .ZN(n13040) );
  NAND2_X1 U12670 ( .A1(n13036), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10180) );
  NAND2_X1 U12671 ( .A1(n13040), .A2(n10180), .ZN(n14779) );
  INV_X1 U12672 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10181) );
  MUX2_X1 U12673 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10181), .S(n10182), .Z(
        n14778) );
  NAND2_X1 U12674 ( .A1(n14779), .A2(n14778), .ZN(n14777) );
  NAND2_X1 U12675 ( .A1(n10182), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n13054) );
  NAND2_X1 U12676 ( .A1(n14777), .A2(n13054), .ZN(n10185) );
  INV_X1 U12677 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10183) );
  MUX2_X1 U12678 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10183), .S(n13052), .Z(
        n10184) );
  NAND2_X1 U12679 ( .A1(n10185), .A2(n10184), .ZN(n13056) );
  NAND2_X1 U12680 ( .A1(n13052), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10186) );
  NAND2_X1 U12681 ( .A1(n13056), .A2(n10186), .ZN(n10246) );
  INV_X1 U12682 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10187) );
  MUX2_X1 U12683 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n10187), .S(n10188), .Z(
        n10245) );
  NAND2_X1 U12684 ( .A1(n10246), .A2(n10245), .ZN(n10244) );
  NAND2_X1 U12685 ( .A1(n10188), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10189) );
  AND2_X1 U12686 ( .A1(n10244), .A2(n10189), .ZN(n10199) );
  INV_X1 U12687 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n14094) );
  NOR3_X1 U12688 ( .A1(n14836), .A2(n10199), .A3(n14094), .ZN(n10190) );
  NOR3_X1 U12689 ( .A1(n10191), .A2(n14841), .A3(n10190), .ZN(n10205) );
  NAND2_X1 U12690 ( .A1(n10204), .A2(n10192), .ZN(n10259) );
  MUX2_X1 U12691 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n10192), .S(n10266), .Z(
        n10193) );
  NAND2_X1 U12692 ( .A1(n10194), .A2(n10193), .ZN(n10260) );
  OAI21_X1 U12693 ( .B1(n10194), .B2(n10259), .A(n10260), .ZN(n10197) );
  INV_X1 U12694 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10195) );
  NAND2_X1 U12695 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n11145) );
  OAI21_X1 U12696 ( .B1(n14845), .B2(n10195), .A(n11145), .ZN(n10196) );
  AOI21_X1 U12697 ( .B1(n10197), .B2(n14820), .A(n10196), .ZN(n10203) );
  NOR3_X1 U12698 ( .A1(n10199), .A2(P2_REG1_REG_9__SCAN_IN), .A3(n10266), .ZN(
        n10201) );
  MUX2_X1 U12699 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n14094), .S(n10266), .Z(
        n10198) );
  NAND2_X1 U12700 ( .A1(n10199), .A2(n10198), .ZN(n10265) );
  INV_X1 U12701 ( .A(n10265), .ZN(n10200) );
  OAI21_X1 U12702 ( .B1(n10201), .B2(n10200), .A(n14825), .ZN(n10202) );
  OAI211_X1 U12703 ( .C1(n10205), .C2(n10204), .A(n10203), .B(n10202), .ZN(
        P2_U3223) );
  INV_X1 U12704 ( .A(n10386), .ZN(n10380) );
  INV_X1 U12705 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10206) );
  OAI222_X1 U12706 ( .A1(n13438), .A2(n10207), .B1(n10380), .B2(P2_U3088), 
        .C1(n10206), .C2(n13440), .ZN(P2_U3317) );
  INV_X1 U12707 ( .A(n9855), .ZN(n10209) );
  CLKBUF_X1 U12708 ( .A(n10213), .Z(n10237) );
  INV_X1 U12709 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10210) );
  NOR2_X1 U12710 ( .A1(n10237), .A2(n10210), .ZN(P3_U3252) );
  INV_X1 U12711 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10211) );
  NOR2_X1 U12712 ( .A1(n10237), .A2(n10211), .ZN(P3_U3254) );
  INV_X1 U12713 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10212) );
  NOR2_X1 U12714 ( .A1(n10237), .A2(n10212), .ZN(P3_U3250) );
  INV_X1 U12715 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10214) );
  NOR2_X1 U12716 ( .A1(n10237), .A2(n10214), .ZN(P3_U3260) );
  INV_X1 U12717 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10215) );
  NOR2_X1 U12718 ( .A1(n10237), .A2(n10215), .ZN(P3_U3256) );
  INV_X1 U12719 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10216) );
  NOR2_X1 U12720 ( .A1(n10237), .A2(n10216), .ZN(P3_U3247) );
  INV_X1 U12721 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10217) );
  NOR2_X1 U12722 ( .A1(n10237), .A2(n10217), .ZN(P3_U3246) );
  INV_X1 U12723 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10218) );
  NOR2_X1 U12724 ( .A1(n10237), .A2(n10218), .ZN(P3_U3249) );
  INV_X1 U12725 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10219) );
  NOR2_X1 U12726 ( .A1(n10213), .A2(n10219), .ZN(P3_U3244) );
  INV_X1 U12727 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10220) );
  NOR2_X1 U12728 ( .A1(n10237), .A2(n10220), .ZN(P3_U3248) );
  INV_X1 U12729 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10221) );
  NOR2_X1 U12730 ( .A1(n10237), .A2(n10221), .ZN(P3_U3253) );
  INV_X1 U12731 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10222) );
  NOR2_X1 U12732 ( .A1(n10213), .A2(n10222), .ZN(P3_U3242) );
  INV_X1 U12733 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10223) );
  NOR2_X1 U12734 ( .A1(n10213), .A2(n10223), .ZN(P3_U3245) );
  INV_X1 U12735 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10224) );
  NOR2_X1 U12736 ( .A1(n10213), .A2(n10224), .ZN(P3_U3241) );
  INV_X1 U12737 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n14128) );
  NOR2_X1 U12738 ( .A1(n10213), .A2(n14128), .ZN(P3_U3243) );
  INV_X1 U12739 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10225) );
  NOR2_X1 U12740 ( .A1(n10213), .A2(n10225), .ZN(P3_U3240) );
  INV_X1 U12741 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10226) );
  NOR2_X1 U12742 ( .A1(n10237), .A2(n10226), .ZN(P3_U3263) );
  INV_X1 U12743 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10227) );
  NOR2_X1 U12744 ( .A1(n10213), .A2(n10227), .ZN(P3_U3262) );
  INV_X1 U12745 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10228) );
  NOR2_X1 U12746 ( .A1(n10237), .A2(n10228), .ZN(P3_U3261) );
  INV_X1 U12747 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10229) );
  NOR2_X1 U12748 ( .A1(n10213), .A2(n10229), .ZN(P3_U3238) );
  INV_X1 U12749 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10230) );
  NOR2_X1 U12750 ( .A1(n10237), .A2(n10230), .ZN(P3_U3259) );
  INV_X1 U12751 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n14146) );
  NOR2_X1 U12752 ( .A1(n10213), .A2(n14146), .ZN(P3_U3258) );
  INV_X1 U12753 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10231) );
  NOR2_X1 U12754 ( .A1(n10237), .A2(n10231), .ZN(P3_U3257) );
  INV_X1 U12755 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10232) );
  NOR2_X1 U12756 ( .A1(n10213), .A2(n10232), .ZN(P3_U3237) );
  INV_X1 U12757 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10233) );
  NOR2_X1 U12758 ( .A1(n10237), .A2(n10233), .ZN(P3_U3255) );
  INV_X1 U12759 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10234) );
  NOR2_X1 U12760 ( .A1(n10213), .A2(n10234), .ZN(P3_U3236) );
  INV_X1 U12761 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10235) );
  NOR2_X1 U12762 ( .A1(n10237), .A2(n10235), .ZN(P3_U3235) );
  INV_X1 U12763 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n14173) );
  NOR2_X1 U12764 ( .A1(n10237), .A2(n14173), .ZN(P3_U3234) );
  INV_X1 U12765 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10236) );
  NOR2_X1 U12766 ( .A1(n10237), .A2(n10236), .ZN(P3_U3251) );
  INV_X1 U12767 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10238) );
  NOR2_X1 U12768 ( .A1(n10237), .A2(n10238), .ZN(P3_U3239) );
  INV_X1 U12769 ( .A(n10239), .ZN(n10243) );
  NAND3_X1 U12770 ( .A1(n13050), .A2(n10241), .A3(n10240), .ZN(n10242) );
  NAND3_X1 U12771 ( .A1(n10243), .A2(n14820), .A3(n10242), .ZN(n10250) );
  NAND2_X1 U12772 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n12212) );
  OAI211_X1 U12773 ( .C1(n10246), .C2(n10245), .A(n14825), .B(n10244), .ZN(
        n10247) );
  NAND2_X1 U12774 ( .A1(n12212), .A2(n10247), .ZN(n10248) );
  AOI21_X1 U12775 ( .B1(n14818), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n10248), .ZN(
        n10249) );
  OAI211_X1 U12776 ( .C1(n10396), .C2(n10251), .A(n10250), .B(n10249), .ZN(
        P2_U3222) );
  AOI22_X1 U12777 ( .A1(n14825), .A2(P2_REG1_REG_0__SCAN_IN), .B1(n14820), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n10254) );
  OAI22_X1 U12778 ( .A1(n14838), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n14836), .ZN(n10252) );
  NOR2_X1 U12779 ( .A1(n10252), .A2(n14841), .ZN(n10253) );
  MUX2_X1 U12780 ( .A(n10254), .B(n10253), .S(P2_IR_REG_0__SCAN_IN), .Z(n10256) );
  AOI22_X1 U12781 ( .A1(n14818), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n10255) );
  NAND2_X1 U12782 ( .A1(n10256), .A2(n10255), .ZN(P2_U3214) );
  OAI222_X1 U12783 ( .A1(n12880), .A2(n10258), .B1(n12040), .B2(n10257), .C1(
        n15007), .C2(P3_U3151), .ZN(P3_U3282) );
  NAND2_X1 U12784 ( .A1(n10260), .A2(n10259), .ZN(n10263) );
  INV_X1 U12785 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10261) );
  MUX2_X1 U12786 ( .A(n10261), .B(P2_REG2_REG_10__SCAN_IN), .S(n10386), .Z(
        n10262) );
  NOR2_X1 U12787 ( .A1(n10263), .A2(n10262), .ZN(n10385) );
  AOI211_X1 U12788 ( .C1(n10263), .C2(n10262), .A(n14838), .B(n10385), .ZN(
        n10264) );
  INV_X1 U12789 ( .A(n10264), .ZN(n10273) );
  NAND2_X1 U12790 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n11448)
         );
  INV_X1 U12791 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n14901) );
  MUX2_X1 U12792 ( .A(n14901), .B(P2_REG1_REG_10__SCAN_IN), .S(n10386), .Z(
        n10268) );
  OAI21_X1 U12793 ( .B1(n10266), .B2(P2_REG1_REG_9__SCAN_IN), .A(n10265), .ZN(
        n10267) );
  NOR2_X1 U12794 ( .A1(n10267), .A2(n10268), .ZN(n13073) );
  AOI211_X1 U12795 ( .C1(n10268), .C2(n10267), .A(n13073), .B(n14836), .ZN(
        n10269) );
  INV_X1 U12796 ( .A(n10269), .ZN(n10270) );
  NAND2_X1 U12797 ( .A1(n11448), .A2(n10270), .ZN(n10271) );
  AOI21_X1 U12798 ( .B1(n14818), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n10271), 
        .ZN(n10272) );
  OAI211_X1 U12799 ( .C1(n10396), .C2(n10380), .A(n10273), .B(n10272), .ZN(
        P2_U3224) );
  INV_X1 U12800 ( .A(n14578), .ZN(n14593) );
  NAND2_X1 U12801 ( .A1(n10275), .A2(n10274), .ZN(n10337) );
  INV_X1 U12802 ( .A(n10337), .ZN(n10332) );
  NOR2_X1 U12803 ( .A1(n6588), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10276) );
  NOR2_X1 U12804 ( .A1(n10276), .A2(n9784), .ZN(n13590) );
  OAI21_X1 U12805 ( .B1(n10277), .B2(P1_REG1_REG_0__SCAN_IN), .A(n13590), .ZN(
        n10278) );
  XNOR2_X1 U12806 ( .A(n10278), .B(n14284), .ZN(n10279) );
  AOI22_X1 U12807 ( .A1(n10332), .A2(n10279), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10280) );
  OAI21_X1 U12808 ( .B1(n14593), .B2(n6672), .A(n10280), .ZN(P1_U3243) );
  INV_X1 U12809 ( .A(P3_DATAO_REG_9__SCAN_IN), .ZN(n14186) );
  NAND2_X1 U12810 ( .A1(n11807), .A2(P3_U3897), .ZN(n10281) );
  OAI21_X1 U12811 ( .B1(P3_U3897), .B2(n14186), .A(n10281), .ZN(P3_U3500) );
  INV_X1 U12812 ( .A(n10282), .ZN(n10285) );
  INV_X1 U12813 ( .A(n13066), .ZN(n10388) );
  OAI222_X1 U12814 ( .A1(n13440), .A2(n10283), .B1(n13438), .B2(n10285), .C1(
        P2_U3088), .C2(n10388), .ZN(P2_U3316) );
  INV_X1 U12815 ( .A(n10519), .ZN(n10524) );
  OAI222_X1 U12816 ( .A1(n10524), .A2(P1_U3086), .B1(n14281), .B2(n10285), 
        .C1(n10284), .C2(n14278), .ZN(P1_U3344) );
  INV_X1 U12817 ( .A(P3_DATAO_REG_7__SCAN_IN), .ZN(n14152) );
  NAND2_X1 U12818 ( .A1(n11562), .A2(P3_U3897), .ZN(n10286) );
  OAI21_X1 U12819 ( .B1(P3_U3897), .B2(n14152), .A(n10286), .ZN(P3_U3498) );
  NAND3_X1 U12820 ( .A1(n14879), .A2(n10288), .A3(n10287), .ZN(n10491) );
  INV_X1 U12821 ( .A(n10491), .ZN(n10289) );
  INV_X1 U12822 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10296) );
  AND2_X1 U12823 ( .A1(n13279), .A2(n9954), .ZN(n10291) );
  OR2_X1 U12824 ( .A1(n14859), .A2(n10291), .ZN(n10292) );
  NAND2_X1 U12825 ( .A1(n6429), .A2(n12946), .ZN(n10672) );
  NAND2_X1 U12826 ( .A1(n10292), .A2(n10672), .ZN(n14864) );
  INV_X1 U12827 ( .A(n14864), .ZN(n10294) );
  NAND2_X1 U12828 ( .A1(n10668), .A2(n10293), .ZN(n14860) );
  OAI211_X1 U12829 ( .C1(n14859), .C2(n11535), .A(n10294), .B(n14860), .ZN(
        n13375) );
  NAND2_X1 U12830 ( .A1(n13375), .A2(n14898), .ZN(n10295) );
  OAI21_X1 U12831 ( .B1(n14898), .B2(n10296), .A(n10295), .ZN(P2_U3430) );
  NOR4_X1 U12832 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n10305) );
  NOR4_X1 U12833 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n10304) );
  NOR4_X1 U12834 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n10300) );
  NOR4_X1 U12835 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n10299) );
  NOR4_X1 U12836 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n10298) );
  NOR4_X1 U12837 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n10297) );
  NAND4_X1 U12838 ( .A1(n10300), .A2(n10299), .A3(n10298), .A4(n10297), .ZN(
        n10301) );
  NOR4_X1 U12839 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n10302), .A4(n10301), .ZN(n10303) );
  NAND3_X1 U12840 ( .A1(n10305), .A2(n10304), .A3(n10303), .ZN(n10306) );
  NAND2_X1 U12841 ( .A1(n10310), .A2(n10306), .ZN(n10746) );
  OR2_X1 U12842 ( .A1(n11086), .A2(n11268), .ZN(n14704) );
  AND2_X1 U12843 ( .A1(n10746), .A2(n11054), .ZN(n10314) );
  NOR2_X1 U12844 ( .A1(n10102), .A2(n10311), .ZN(n10307) );
  NAND2_X1 U12845 ( .A1(n10310), .A2(n10309), .ZN(n10313) );
  NAND2_X2 U12846 ( .A1(n10315), .A2(n10591), .ZN(n12160) );
  OR2_X1 U12847 ( .A1(n10315), .A2(n10591), .ZN(n10316) );
  NAND2_X1 U12848 ( .A1(n11058), .A2(n11268), .ZN(n14703) );
  NAND2_X1 U12849 ( .A1(n9719), .A2(n13691), .ZN(n10318) );
  OAI21_X1 U12850 ( .B1(n14729), .B2(n14708), .A(n11258), .ZN(n10319) );
  NOR2_X1 U12851 ( .A1(n11085), .A2(n9719), .ZN(n10593) );
  AOI22_X1 U12852 ( .A1(n10630), .A2(n13983), .B1(n10593), .B2(n11125), .ZN(
        n11261) );
  NAND2_X1 U12853 ( .A1(n10319), .A2(n11261), .ZN(n10751) );
  NAND2_X1 U12854 ( .A1(n14745), .A2(n10751), .ZN(n10320) );
  OAI21_X1 U12855 ( .B1(n14745), .B2(n10602), .A(n10320), .ZN(P1_U3528) );
  OAI222_X1 U12856 ( .A1(n12880), .A2(n10322), .B1(n12040), .B2(n10321), .C1(
        n12474), .C2(P3_U3151), .ZN(P3_U3281) );
  MUX2_X1 U12857 ( .A(n10323), .B(P1_REG1_REG_2__SCAN_IN), .S(n13598), .Z(
        n10327) );
  AND2_X1 U12858 ( .A1(n14284), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10325) );
  OR2_X1 U12859 ( .A1(n13577), .A2(n10324), .ZN(n13591) );
  NAND2_X1 U12860 ( .A1(n10327), .A2(n10326), .ZN(n13594) );
  INV_X1 U12861 ( .A(n13594), .ZN(n13613) );
  NOR2_X1 U12862 ( .A1(n13598), .A2(n10323), .ZN(n13612) );
  MUX2_X1 U12863 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10328), .S(n13607), .Z(
        n13614) );
  OAI21_X1 U12864 ( .B1(n13613), .B2(n13612), .A(n13614), .ZN(n14574) );
  NAND2_X1 U12865 ( .A1(n13607), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n14573) );
  INV_X1 U12866 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n14735) );
  MUX2_X1 U12867 ( .A(n14735), .B(P1_REG1_REG_4__SCAN_IN), .S(n14579), .Z(
        n14572) );
  AOI21_X1 U12868 ( .B1(n14574), .B2(n14573), .A(n14572), .ZN(n14571) );
  MUX2_X1 U12869 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6612), .S(n13621), .Z(
        n13628) );
  MUX2_X1 U12870 ( .A(n9305), .B(P1_REG1_REG_6__SCAN_IN), .S(n10414), .Z(
        n10412) );
  NOR2_X1 U12871 ( .A1(n10419), .A2(n9305), .ZN(n13634) );
  MUX2_X1 U12872 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n10329), .S(n13638), .Z(
        n13633) );
  OAI21_X1 U12873 ( .B1(n13635), .B2(n13634), .A(n13633), .ZN(n13637) );
  OAI21_X1 U12874 ( .B1(n10329), .B2(n10330), .A(n13637), .ZN(n10369) );
  MUX2_X1 U12875 ( .A(n10331), .B(P1_REG1_REG_8__SCAN_IN), .S(n10372), .Z(
        n10370) );
  NOR2_X1 U12876 ( .A1(n10369), .A2(n10370), .ZN(n13651) );
  NOR2_X1 U12877 ( .A1(n10372), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n13649) );
  MUX2_X1 U12878 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9349), .S(n13656), .Z(
        n13650) );
  OAI21_X1 U12879 ( .B1(n13651), .B2(n13649), .A(n13650), .ZN(n13648) );
  OAI21_X1 U12880 ( .B1(n13656), .B2(P1_REG1_REG_9__SCAN_IN), .A(n13648), .ZN(
        n10334) );
  INV_X1 U12881 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n14743) );
  MUX2_X1 U12882 ( .A(n14743), .B(P1_REG1_REG_10__SCAN_IN), .S(n10426), .Z(
        n10333) );
  NAND2_X1 U12883 ( .A1(n10332), .A2(n6588), .ZN(n13688) );
  NOR2_X1 U12884 ( .A1(n10334), .A2(n10333), .ZN(n10423) );
  AOI211_X1 U12885 ( .C1(n10334), .C2(n10333), .A(n13688), .B(n10423), .ZN(
        n10368) );
  NOR2_X2 U12886 ( .A1(n10337), .A2(n13587), .ZN(n14595) );
  INV_X1 U12887 ( .A(n10426), .ZN(n10366) );
  NOR2_X1 U12888 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10335), .ZN(n11756) );
  AOI21_X1 U12889 ( .B1(n14578), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n11756), 
        .ZN(n10365) );
  OR2_X1 U12890 ( .A1(n9784), .A2(n6588), .ZN(n10336) );
  NOR2_X2 U12891 ( .A1(n10337), .A2(n10336), .ZN(n14602) );
  MUX2_X1 U12892 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10338), .S(n13607), .Z(
        n10343) );
  MUX2_X1 U12893 ( .A(n10339), .B(P1_REG2_REG_2__SCAN_IN), .S(n13598), .Z(
        n10341) );
  MUX2_X1 U12894 ( .A(n14202), .B(P1_REG2_REG_1__SCAN_IN), .S(n13577), .Z(
        n13580) );
  AND2_X1 U12895 ( .A1(n14284), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n13586) );
  NAND2_X1 U12896 ( .A1(n13580), .A2(n13586), .ZN(n13600) );
  INV_X1 U12897 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n14202) );
  OR2_X1 U12898 ( .A1(n13577), .A2(n14202), .ZN(n13599) );
  NAND2_X1 U12899 ( .A1(n13600), .A2(n13599), .ZN(n10340) );
  NAND2_X1 U12900 ( .A1(n10341), .A2(n10340), .ZN(n13609) );
  INV_X1 U12901 ( .A(n13598), .ZN(n13596) );
  NAND2_X1 U12902 ( .A1(n13596), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n13608) );
  NAND2_X1 U12903 ( .A1(n13609), .A2(n13608), .ZN(n10342) );
  NAND2_X1 U12904 ( .A1(n10343), .A2(n10342), .ZN(n14582) );
  NAND2_X1 U12905 ( .A1(n13607), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n14581) );
  NAND2_X1 U12906 ( .A1(n14582), .A2(n14581), .ZN(n10346) );
  MUX2_X1 U12907 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10344), .S(n14579), .Z(
        n10345) );
  NAND2_X1 U12908 ( .A1(n10346), .A2(n10345), .ZN(n14584) );
  NAND2_X1 U12909 ( .A1(n14579), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n13623) );
  NAND2_X1 U12910 ( .A1(n14584), .A2(n13623), .ZN(n10348) );
  INV_X1 U12911 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n11083) );
  MUX2_X1 U12912 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n11083), .S(n13621), .Z(
        n10347) );
  NAND2_X1 U12913 ( .A1(n10348), .A2(n10347), .ZN(n13625) );
  NAND2_X1 U12914 ( .A1(n13621), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10416) );
  NAND2_X1 U12915 ( .A1(n13625), .A2(n10416), .ZN(n10351) );
  MUX2_X1 U12916 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10349), .S(n10414), .Z(
        n10350) );
  NAND2_X1 U12917 ( .A1(n10351), .A2(n10350), .ZN(n13641) );
  NAND2_X1 U12918 ( .A1(n10414), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n13640) );
  NAND2_X1 U12919 ( .A1(n13641), .A2(n13640), .ZN(n10353) );
  MUX2_X1 U12920 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n11513), .S(n13638), .Z(
        n10352) );
  NAND2_X1 U12921 ( .A1(n10353), .A2(n10352), .ZN(n13643) );
  NAND2_X1 U12922 ( .A1(n13638), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10374) );
  NAND2_X1 U12923 ( .A1(n13643), .A2(n10374), .ZN(n10356) );
  INV_X1 U12924 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10354) );
  MUX2_X1 U12925 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10354), .S(n10372), .Z(
        n10355) );
  NAND2_X1 U12926 ( .A1(n10356), .A2(n10355), .ZN(n13659) );
  NAND2_X1 U12927 ( .A1(n10372), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n13658) );
  NAND2_X1 U12928 ( .A1(n13659), .A2(n13658), .ZN(n10358) );
  MUX2_X1 U12929 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n11307), .S(n13656), .Z(
        n10357) );
  NAND2_X1 U12930 ( .A1(n10358), .A2(n10357), .ZN(n13661) );
  NAND2_X1 U12931 ( .A1(n13656), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10362) );
  NAND2_X1 U12932 ( .A1(n13661), .A2(n10362), .ZN(n10360) );
  MUX2_X1 U12933 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n11433), .S(n10426), .Z(
        n10359) );
  NAND2_X1 U12934 ( .A1(n10360), .A2(n10359), .ZN(n10431) );
  MUX2_X1 U12935 ( .A(n11433), .B(P1_REG2_REG_10__SCAN_IN), .S(n10426), .Z(
        n10361) );
  NAND3_X1 U12936 ( .A1(n13661), .A2(n10362), .A3(n10361), .ZN(n10363) );
  NAND3_X1 U12937 ( .A1(n14602), .A2(n10431), .A3(n10363), .ZN(n10364) );
  OAI211_X1 U12938 ( .C1(n13677), .C2(n10366), .A(n10365), .B(n10364), .ZN(
        n10367) );
  OR2_X1 U12939 ( .A1(n10368), .A2(n10367), .ZN(P1_U3253) );
  AOI21_X1 U12940 ( .B1(n10370), .B2(n10369), .A(n13651), .ZN(n10378) );
  NAND2_X1 U12941 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11484) );
  OAI21_X1 U12942 ( .B1(n14593), .B2(n14307), .A(n11484), .ZN(n10371) );
  AOI21_X1 U12943 ( .B1(n10372), .B2(n14595), .A(n10371), .ZN(n10377) );
  MUX2_X1 U12944 ( .A(n10354), .B(P1_REG2_REG_8__SCAN_IN), .S(n10372), .Z(
        n10373) );
  NAND3_X1 U12945 ( .A1(n13643), .A2(n10374), .A3(n10373), .ZN(n10375) );
  NAND3_X1 U12946 ( .A1(n14602), .A2(n13659), .A3(n10375), .ZN(n10376) );
  OAI211_X1 U12947 ( .C1(n10378), .C2(n13688), .A(n10377), .B(n10376), .ZN(
        P1_U3251) );
  INV_X1 U12948 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n14512) );
  NOR2_X1 U12949 ( .A1(n10390), .A2(n14512), .ZN(n10379) );
  AOI21_X1 U12950 ( .B1(n14512), .B2(n10390), .A(n10379), .ZN(n10384) );
  INV_X1 U12951 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n13067) );
  NOR2_X1 U12952 ( .A1(n10380), .A2(n14901), .ZN(n13068) );
  MUX2_X1 U12953 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n13067), .S(n13066), .Z(
        n10381) );
  OAI21_X1 U12954 ( .B1(n13073), .B2(n13068), .A(n10381), .ZN(n13071) );
  OAI21_X1 U12955 ( .B1(n13067), .B2(n10388), .A(n13071), .ZN(n10383) );
  INV_X1 U12956 ( .A(n10390), .ZN(n11411) );
  NOR2_X1 U12957 ( .A1(n11411), .A2(n14512), .ZN(n10382) );
  AOI211_X1 U12958 ( .C1(n11411), .C2(n14512), .A(n10382), .B(n10383), .ZN(
        n11397) );
  AOI21_X1 U12959 ( .B1(n10384), .B2(n10383), .A(n11397), .ZN(n10401) );
  AOI21_X1 U12960 ( .B1(n10386), .B2(P2_REG2_REG_10__SCAN_IN), .A(n10385), 
        .ZN(n13062) );
  INV_X1 U12961 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10387) );
  MUX2_X1 U12962 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n10387), .S(n13066), .Z(
        n13061) );
  NAND2_X1 U12963 ( .A1(n13062), .A2(n13061), .ZN(n13060) );
  NAND2_X1 U12964 ( .A1(n10388), .A2(n10387), .ZN(n10393) );
  INV_X1 U12965 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n10389) );
  OR2_X1 U12966 ( .A1(n10390), .A2(n10389), .ZN(n10392) );
  NAND2_X1 U12967 ( .A1(n10390), .A2(n10389), .ZN(n10391) );
  AND2_X1 U12968 ( .A1(n10392), .A2(n10391), .ZN(n10394) );
  AOI21_X1 U12969 ( .B1(n13060), .B2(n10393), .A(n10394), .ZN(n11410) );
  AND3_X1 U12970 ( .A1(n13060), .A2(n10394), .A3(n10393), .ZN(n10395) );
  OAI21_X1 U12971 ( .B1(n11410), .B2(n10395), .A(n14820), .ZN(n10400) );
  NOR2_X1 U12972 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11657), .ZN(n10398) );
  NOR2_X1 U12973 ( .A1(n10396), .A2(n11411), .ZN(n10397) );
  AOI211_X1 U12974 ( .C1(n14818), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n10398), 
        .B(n10397), .ZN(n10399) );
  OAI211_X1 U12975 ( .C1(n10401), .C2(n14836), .A(n10400), .B(n10399), .ZN(
        P2_U3226) );
  INV_X1 U12976 ( .A(n10407), .ZN(n10405) );
  INV_X1 U12977 ( .A(n10650), .ZN(n10403) );
  NAND2_X1 U12978 ( .A1(n10403), .A2(n10402), .ZN(n10406) );
  INV_X1 U12979 ( .A(n10406), .ZN(n10404) );
  OAI21_X1 U12980 ( .B1(n10405), .B2(n10404), .A(n12996), .ZN(n10411) );
  NOR2_X1 U12981 ( .A1(n10407), .A2(n10406), .ZN(n10651) );
  OAI22_X1 U12982 ( .A1(n8272), .A2(n12967), .B1(n10408), .B2(n12984), .ZN(
        n10707) );
  AOI22_X1 U12983 ( .A1(n10712), .A2(n12976), .B1(n12992), .B2(n10707), .ZN(
        n10410) );
  MUX2_X1 U12984 ( .A(n12990), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n10409) );
  OAI211_X1 U12985 ( .C1(n10411), .C2(n10651), .A(n10410), .B(n10409), .ZN(
        P2_U3190) );
  AOI211_X1 U12986 ( .C1(n10413), .C2(n10412), .A(n13635), .B(n13688), .ZN(
        n10422) );
  MUX2_X1 U12987 ( .A(n10349), .B(P1_REG2_REG_6__SCAN_IN), .S(n10414), .Z(
        n10415) );
  NAND3_X1 U12988 ( .A1(n13625), .A2(n10416), .A3(n10415), .ZN(n10417) );
  AND3_X1 U12989 ( .A1(n14602), .A2(n13641), .A3(n10417), .ZN(n10421) );
  NAND2_X1 U12990 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n11121) );
  NAND2_X1 U12991 ( .A1(n14578), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n10418) );
  OAI211_X1 U12992 ( .C1(n13677), .C2(n10419), .A(n11121), .B(n10418), .ZN(
        n10420) );
  OR3_X1 U12993 ( .A1(n10422), .A2(n10421), .A3(n10420), .ZN(P1_U3249) );
  MUX2_X1 U12994 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9382), .S(n10519), .Z(
        n10425) );
  OAI21_X1 U12995 ( .B1(n10425), .B2(n10424), .A(n10528), .ZN(n10436) );
  AND2_X1 U12996 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n11793) );
  AOI21_X1 U12997 ( .B1(n14578), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n11793), 
        .ZN(n10434) );
  NAND2_X1 U12998 ( .A1(n10426), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10430) );
  NAND2_X1 U12999 ( .A1(n10431), .A2(n10430), .ZN(n10428) );
  INV_X1 U13000 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11554) );
  MUX2_X1 U13001 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n11554), .S(n10519), .Z(
        n10427) );
  NAND2_X1 U13002 ( .A1(n10428), .A2(n10427), .ZN(n10521) );
  MUX2_X1 U13003 ( .A(n11554), .B(P1_REG2_REG_11__SCAN_IN), .S(n10519), .Z(
        n10429) );
  NAND3_X1 U13004 ( .A1(n10431), .A2(n10430), .A3(n10429), .ZN(n10432) );
  NAND3_X1 U13005 ( .A1(n14602), .A2(n10521), .A3(n10432), .ZN(n10433) );
  OAI211_X1 U13006 ( .C1(n13677), .C2(n10524), .A(n10434), .B(n10433), .ZN(
        n10435) );
  AOI21_X1 U13007 ( .B1(n10436), .B2(n14597), .A(n10435), .ZN(n10437) );
  INV_X1 U13008 ( .A(n10437), .ZN(P1_U3254) );
  OAI222_X1 U13009 ( .A1(n13438), .A2(n10444), .B1(n11412), .B2(P2_U3088), 
        .C1(n10438), .C2(n13440), .ZN(P2_U3314) );
  INV_X1 U13010 ( .A(n10439), .ZN(n10460) );
  OAI222_X1 U13011 ( .A1(n13438), .A2(n10460), .B1(n11411), .B2(P2_U3088), 
        .C1(n10440), .C2(n13440), .ZN(P2_U3315) );
  OAI222_X1 U13012 ( .A1(n12880), .A2(n10442), .B1(n12040), .B2(n10441), .C1(
        n14437), .C2(P3_U3151), .ZN(P3_U3280) );
  INV_X1 U13013 ( .A(n14596), .ZN(n10929) );
  OAI222_X1 U13014 ( .A1(P1_U3086), .A2(n10929), .B1(n14281), .B2(n10444), 
        .C1(n10443), .C2(n14278), .ZN(P1_U3342) );
  INV_X1 U13015 ( .A(n14960), .ZN(n15008) );
  INV_X1 U13016 ( .A(n15023), .ZN(n12472) );
  OAI21_X1 U13017 ( .B1(n10447), .B2(n9033), .A(n10446), .ZN(n10454) );
  INV_X1 U13018 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15055) );
  OAI22_X1 U13019 ( .A1(n15005), .A2(n14291), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15055), .ZN(n10453) );
  NAND2_X1 U13020 ( .A1(n10449), .A2(n10448), .ZN(n10450) );
  AOI21_X1 U13021 ( .B1(n10451), .B2(n10450), .A(n15017), .ZN(n10452) );
  AOI211_X1 U13022 ( .C1(n12472), .C2(n10454), .A(n10453), .B(n10452), .ZN(
        n10459) );
  XNOR2_X1 U13023 ( .A(n10456), .B(n10455), .ZN(n10457) );
  NAND2_X1 U13024 ( .A1(n10457), .A2(n14963), .ZN(n10458) );
  OAI211_X1 U13025 ( .C1(n15008), .C2(n9121), .A(n10459), .B(n10458), .ZN(
        P3_U3184) );
  INV_X1 U13026 ( .A(n10532), .ZN(n10931) );
  OAI222_X1 U13027 ( .A1(n14278), .A2(n10461), .B1(n14281), .B2(n10460), .C1(
        P1_U3086), .C2(n10931), .ZN(P1_U3343) );
  OAI21_X1 U13028 ( .B1(n10464), .B2(n10463), .A(n10462), .ZN(n10476) );
  AOI21_X1 U13029 ( .B1(n10467), .B2(n10466), .A(n10465), .ZN(n10474) );
  OAI21_X1 U13030 ( .B1(n10470), .B2(n10469), .A(n10468), .ZN(n10471) );
  NAND2_X1 U13031 ( .A1(n9160), .A2(n10471), .ZN(n10473) );
  INV_X1 U13032 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n14145) );
  NOR2_X1 U13033 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14145), .ZN(n11014) );
  AOI21_X1 U13034 ( .B1(n14983), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n11014), .ZN(
        n10472) );
  OAI211_X1 U13035 ( .C1(n10474), .C2(n15023), .A(n10473), .B(n10472), .ZN(
        n10475) );
  AOI21_X1 U13036 ( .B1(n14963), .B2(n10476), .A(n10475), .ZN(n10477) );
  OAI21_X1 U13037 ( .B1(n10478), .B2(n15008), .A(n10477), .ZN(P3_U3186) );
  INV_X1 U13038 ( .A(n10479), .ZN(n10480) );
  AOI21_X1 U13039 ( .B1(n10481), .B2(n9915), .A(n10480), .ZN(n10970) );
  INV_X1 U13040 ( .A(n10970), .ZN(n10489) );
  AOI21_X1 U13041 ( .B1(n10668), .B2(n10967), .A(n7779), .ZN(n10482) );
  AND2_X1 U13042 ( .A1(n10482), .A2(n10613), .ZN(n10965) );
  OAI21_X1 U13043 ( .B1(n10484), .B2(n9915), .A(n10483), .ZN(n10485) );
  NAND2_X1 U13044 ( .A1(n10485), .A2(n14475), .ZN(n10488) );
  NAND2_X1 U13045 ( .A1(n13029), .A2(n12946), .ZN(n10487) );
  NAND2_X1 U13046 ( .A1(n13030), .A2(n12986), .ZN(n10486) );
  AND2_X1 U13047 ( .A1(n10487), .A2(n10486), .ZN(n10693) );
  NAND2_X1 U13048 ( .A1(n10488), .A2(n10693), .ZN(n10964) );
  AOI211_X1 U13049 ( .C1(n10489), .C2(n14511), .A(n10965), .B(n10964), .ZN(
        n10498) );
  NOR2_X1 U13050 ( .A1(n10491), .A2(n10490), .ZN(n10493) );
  AOI22_X1 U13051 ( .A1(n13351), .A2(n10967), .B1(n14900), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n10494) );
  OAI21_X1 U13052 ( .B1(n10498), .B2(n14900), .A(n10494), .ZN(P2_U3500) );
  INV_X1 U13053 ( .A(n13407), .ZN(n13420) );
  INV_X1 U13054 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10495) );
  OAI22_X1 U13055 ( .A1(n13420), .A2(n10694), .B1(n14898), .B2(n10495), .ZN(
        n10496) );
  INV_X1 U13056 ( .A(n10496), .ZN(n10497) );
  OAI21_X1 U13057 ( .B1(n10498), .B2(n14896), .A(n10497), .ZN(P2_U3433) );
  NAND2_X1 U13058 ( .A1(n10499), .A2(n15130), .ZN(n10500) );
  OR2_X1 U13059 ( .A1(n10581), .A2(n10500), .ZN(n10502) );
  OR2_X1 U13060 ( .A1(n15062), .A2(n15059), .ZN(n10501) );
  AND2_X1 U13061 ( .A1(n10502), .A2(n10501), .ZN(n10821) );
  MUX2_X1 U13062 ( .A(n10503), .B(n10821), .S(n15166), .Z(n10504) );
  OAI21_X1 U13063 ( .B1(n10582), .B2(n12817), .A(n10504), .ZN(P3_U3459) );
  XOR2_X1 U13064 ( .A(n14907), .B(n10505), .Z(n10518) );
  AOI21_X1 U13065 ( .B1(n15147), .B2(n10507), .A(n10506), .ZN(n10515) );
  INV_X1 U13066 ( .A(n10508), .ZN(n10509) );
  NOR2_X1 U13067 ( .A1(n10509), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n10510) );
  OAI21_X1 U13068 ( .B1(n10511), .B2(n10510), .A(n12472), .ZN(n10514) );
  INV_X1 U13069 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10578) );
  NOR2_X1 U13070 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10578), .ZN(n10512) );
  AOI21_X1 U13071 ( .B1(n14983), .B2(P3_ADDR_REG_1__SCAN_IN), .A(n10512), .ZN(
        n10513) );
  OAI211_X1 U13072 ( .C1(n10515), .C2(n15017), .A(n10514), .B(n10513), .ZN(
        n10516) );
  AOI21_X1 U13073 ( .B1(n8437), .B2(n14960), .A(n10516), .ZN(n10517) );
  OAI21_X1 U13074 ( .B1(n15015), .B2(n10518), .A(n10517), .ZN(P3_U3183) );
  MUX2_X1 U13075 ( .A(n11687), .B(P1_REG2_REG_12__SCAN_IN), .S(n10532), .Z(
        n10523) );
  NAND2_X1 U13076 ( .A1(n10519), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10520) );
  NAND2_X1 U13077 ( .A1(n10521), .A2(n10520), .ZN(n10522) );
  NOR2_X1 U13078 ( .A1(n10522), .A2(n10523), .ZN(n10930) );
  AOI21_X1 U13079 ( .B1(n10523), .B2(n10522), .A(n10930), .ZN(n10535) );
  INV_X1 U13080 ( .A(n14602), .ZN(n11355) );
  NAND2_X1 U13081 ( .A1(n10524), .A2(n9382), .ZN(n10526) );
  MUX2_X1 U13082 ( .A(n10525), .B(P1_REG1_REG_12__SCAN_IN), .S(n10532), .Z(
        n10527) );
  AND3_X1 U13083 ( .A1(n10528), .A2(n10527), .A3(n10526), .ZN(n10529) );
  OAI21_X1 U13084 ( .B1(n10923), .B2(n10529), .A(n14597), .ZN(n10534) );
  INV_X1 U13085 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10530) );
  NAND2_X1 U13086 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n11888)
         );
  OAI21_X1 U13087 ( .B1(n14593), .B2(n10530), .A(n11888), .ZN(n10531) );
  AOI21_X1 U13088 ( .B1(n10532), .B2(n14595), .A(n10531), .ZN(n10533) );
  OAI211_X1 U13089 ( .C1(n10535), .C2(n11355), .A(n10534), .B(n10533), .ZN(
        P1_U3255) );
  INV_X1 U13090 ( .A(n10570), .ZN(n10538) );
  OAI211_X1 U13091 ( .C1(n10538), .C2(n10569), .A(n10537), .B(n10536), .ZN(
        n10539) );
  AOI21_X1 U13092 ( .B1(n10572), .B2(n10568), .A(n10539), .ZN(n10540) );
  NOR2_X1 U13093 ( .A1(n10540), .A2(P3_U3151), .ZN(n10541) );
  AOI21_X1 U13094 ( .B1(n10549), .B2(n10570), .A(n10541), .ZN(n10771) );
  AND2_X1 U13095 ( .A1(n10771), .A2(n10542), .ZN(n10807) );
  NAND2_X1 U13096 ( .A1(n10573), .A2(n15084), .ZN(n10543) );
  OR2_X1 U13097 ( .A1(n10572), .A2(n10543), .ZN(n10545) );
  NOR2_X1 U13098 ( .A1(n15130), .A2(n15086), .ZN(n10544) );
  NAND2_X1 U13099 ( .A1(n10549), .A2(n10547), .ZN(n10546) );
  INV_X1 U13100 ( .A(n10547), .ZN(n10548) );
  NAND2_X1 U13101 ( .A1(n10549), .A2(n10548), .ZN(n10550) );
  INV_X1 U13102 ( .A(n15077), .ZN(n10551) );
  OAI22_X1 U13103 ( .A1(n10776), .A2(n12421), .B1(n12433), .B2(n10551), .ZN(
        n10552) );
  AOI21_X1 U13104 ( .B1(n15085), .B2(n12424), .A(n10552), .ZN(n10577) );
  INV_X1 U13105 ( .A(n10554), .ZN(n10555) );
  OAI21_X1 U13106 ( .B1(n10832), .B2(n10984), .A(n11211), .ZN(n10556) );
  NAND2_X4 U13107 ( .A1(n10557), .A2(n10556), .ZN(n12284) );
  NAND3_X1 U13108 ( .A1(n11386), .A2(n15085), .A3(n12452), .ZN(n10562) );
  NAND2_X1 U13109 ( .A1(n10558), .A2(n11386), .ZN(n10561) );
  NAND2_X1 U13110 ( .A1(n10561), .A2(n10560), .ZN(n10774) );
  INV_X1 U13111 ( .A(n15073), .ZN(n10563) );
  AOI21_X1 U13112 ( .B1(n10564), .B2(n12284), .A(n10563), .ZN(n10565) );
  INV_X1 U13113 ( .A(n10566), .ZN(n15082) );
  NAND3_X1 U13114 ( .A1(n15082), .A2(n9801), .A3(n12284), .ZN(n10567) );
  OAI211_X1 U13115 ( .C1(n6572), .C2(n15073), .A(n10775), .B(n10567), .ZN(
        n10575) );
  NAND2_X1 U13116 ( .A1(n10568), .A2(n15130), .ZN(n10571) );
  OAI22_X1 U13117 ( .A1(n10572), .A2(n10571), .B1(n10570), .B2(n10569), .ZN(
        n10574) );
  INV_X1 U13118 ( .A(n12439), .ZN(n12381) );
  NAND2_X1 U13119 ( .A1(n10575), .A2(n12381), .ZN(n10576) );
  OAI211_X1 U13120 ( .C1(n10807), .C2(n10578), .A(n10577), .B(n10576), .ZN(
        P3_U3162) );
  INV_X1 U13121 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10579) );
  MUX2_X1 U13122 ( .A(n10579), .B(n10821), .S(n15146), .Z(n10580) );
  OAI21_X1 U13123 ( .B1(n10582), .B2(n12871), .A(n10580), .ZN(P3_U3390) );
  INV_X1 U13124 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10586) );
  INV_X1 U13125 ( .A(n10581), .ZN(n10584) );
  OAI22_X1 U13126 ( .A1(n12434), .A2(n10582), .B1(n15062), .B2(n12421), .ZN(
        n10583) );
  AOI21_X1 U13127 ( .B1(n12381), .B2(n10584), .A(n10583), .ZN(n10585) );
  OAI21_X1 U13128 ( .B1(n10807), .B2(n10586), .A(n10585), .ZN(P3_U3172) );
  OAI222_X1 U13129 ( .A1(n12880), .A2(n10588), .B1(n12497), .B2(P3_U3151), 
        .C1(n10587), .C2(n12040), .ZN(P3_U3279) );
  INV_X1 U13130 ( .A(n11125), .ZN(n11059) );
  INV_X1 U13131 ( .A(n13761), .ZN(n11052) );
  NAND3_X1 U13132 ( .A1(n11052), .A2(n10748), .A3(n10746), .ZN(n10606) );
  NAND2_X1 U13133 ( .A1(n10606), .A2(n11054), .ZN(n10737) );
  INV_X1 U13134 ( .A(n10592), .ZN(n10589) );
  INV_X1 U13135 ( .A(n10747), .ZN(n10590) );
  NOR2_X1 U13136 ( .A1(n13540), .A2(n13993), .ZN(n13511) );
  NAND2_X1 U13137 ( .A1(n10593), .A2(n10592), .ZN(n13958) );
  INV_X1 U13138 ( .A(n11060), .ZN(n13575) );
  NAND2_X1 U13139 ( .A1(n10634), .A2(n13575), .ZN(n10599) );
  NAND2_X1 U13140 ( .A1(n10596), .A2(n10595), .ZN(n10629) );
  INV_X1 U13141 ( .A(n10596), .ZN(n10597) );
  OR2_X1 U13142 ( .A1(n10900), .A2(n11059), .ZN(n10601) );
  OR2_X1 U13143 ( .A1(n6434), .A2(n11060), .ZN(n10600) );
  OAI21_X1 U13144 ( .B1(n6463), .B2(n10637), .A(n10638), .ZN(n10603) );
  INV_X1 U13145 ( .A(n10603), .ZN(n13585) );
  NAND3_X1 U13146 ( .A1(n11056), .A2(n10604), .A3(n14726), .ZN(n10605) );
  NAND2_X1 U13147 ( .A1(n10737), .A2(n10747), .ZN(n10716) );
  NAND2_X1 U13148 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n10716), .ZN(n10607) );
  OAI21_X1 U13149 ( .B1(n13585), .B2(n13557), .A(n10607), .ZN(n10608) );
  AOI21_X1 U13150 ( .B1(n13511), .B2(n10630), .A(n10608), .ZN(n10609) );
  OAI21_X1 U13151 ( .B1(n11059), .B2(n13526), .A(n10609), .ZN(P1_U3232) );
  OAI21_X1 U13152 ( .B1(n10612), .B2(n10611), .A(n10610), .ZN(n10960) );
  NAND2_X1 U13153 ( .A1(n10613), .A2(n10622), .ZN(n10614) );
  NAND2_X1 U13154 ( .A1(n10614), .A2(n13083), .ZN(n10615) );
  NOR2_X1 U13155 ( .A1(n10704), .A2(n10615), .ZN(n10959) );
  XNOR2_X1 U13156 ( .A(n10617), .B(n10616), .ZN(n10619) );
  AOI22_X1 U13157 ( .A1(n12986), .A2(n6429), .B1(n13028), .B2(n12946), .ZN(
        n10849) );
  INV_X1 U13158 ( .A(n10849), .ZN(n10618) );
  AOI21_X1 U13159 ( .B1(n10619), .B2(n14475), .A(n10618), .ZN(n10963) );
  INV_X1 U13160 ( .A(n10963), .ZN(n10620) );
  AOI211_X1 U13161 ( .C1(n14511), .C2(n10960), .A(n10959), .B(n10620), .ZN(
        n10624) );
  AOI22_X1 U13162 ( .A1(n13407), .A2(n10622), .B1(n14896), .B2(
        P2_REG0_REG_2__SCAN_IN), .ZN(n10621) );
  OAI21_X1 U13163 ( .B1(n10624), .B2(n14896), .A(n10621), .ZN(P2_U3436) );
  AOI22_X1 U13164 ( .A1(n13351), .A2(n10622), .B1(n14900), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n10623) );
  OAI21_X1 U13165 ( .B1(n10624), .B2(n14900), .A(n10623), .ZN(P2_U3501) );
  OR2_X1 U13166 ( .A1(n10900), .A2(n14661), .ZN(n10627) );
  INV_X4 U13167 ( .A(n12160), .ZN(n12122) );
  XNOR2_X1 U13168 ( .A(n10628), .B(n12122), .ZN(n10726) );
  OAI22_X1 U13169 ( .A1(n12159), .A2(n11073), .B1(n14661), .B2(n12071), .ZN(
        n10725) );
  XNOR2_X1 U13170 ( .A(n10726), .B(n10725), .ZN(n10641) );
  NOR2_X1 U13171 ( .A1(n6434), .A2(n10631), .ZN(n10633) );
  AOI21_X1 U13172 ( .B1(n10634), .B2(n10630), .A(n10633), .ZN(n10635) );
  INV_X1 U13173 ( .A(n10635), .ZN(n10636) );
  NAND2_X1 U13174 ( .A1(n10717), .A2(n10639), .ZN(n10640) );
  OAI21_X1 U13175 ( .B1(n10641), .B2(n10640), .A(n10734), .ZN(n10642) );
  NAND2_X1 U13176 ( .A1(n10642), .A2(n13537), .ZN(n10644) );
  INV_X1 U13177 ( .A(n13540), .ZN(n13475) );
  INV_X1 U13178 ( .A(n13981), .ZN(n13991) );
  OAI22_X1 U13179 ( .A1(n11067), .A2(n13993), .B1(n9224), .B2(n13991), .ZN(
        n14632) );
  AOI22_X1 U13180 ( .A1(P1_REG3_REG_2__SCAN_IN), .A2(n10716), .B1(n13475), 
        .B2(n14632), .ZN(n10643) );
  OAI211_X1 U13181 ( .C1(n14661), .C2(n13526), .A(n10644), .B(n10643), .ZN(
        P1_U3237) );
  INV_X1 U13182 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n14182) );
  INV_X1 U13183 ( .A(n10645), .ZN(n10647) );
  INV_X1 U13184 ( .A(n14801), .ZN(n11415) );
  OAI222_X1 U13185 ( .A1(n13440), .A2(n14182), .B1(n13438), .B2(n10647), .C1(
        P2_U3088), .C2(n11415), .ZN(P2_U3313) );
  INV_X1 U13186 ( .A(n11342), .ZN(n11347) );
  OAI222_X1 U13187 ( .A1(n11347), .A2(P1_U3086), .B1(n14281), .B2(n10647), 
        .C1(n10646), .C2(n14278), .ZN(P1_U3341) );
  XNOR2_X1 U13188 ( .A(n10649), .B(n10648), .ZN(n10657) );
  NOR3_X1 U13189 ( .A1(n10651), .A2(n10650), .A3(n10657), .ZN(n12179) );
  AOI21_X1 U13190 ( .B1(n10657), .B2(n10651), .A(n12179), .ZN(n10664) );
  INV_X1 U13191 ( .A(n12990), .ZN(n12964) );
  NAND2_X1 U13192 ( .A1(n12976), .A2(n10761), .ZN(n10656) );
  NAND2_X1 U13193 ( .A1(n13026), .A2(n12946), .ZN(n10653) );
  NAND2_X1 U13194 ( .A1(n13028), .A2(n12986), .ZN(n10652) );
  AND2_X1 U13195 ( .A1(n10653), .A2(n10652), .ZN(n10758) );
  INV_X1 U13196 ( .A(n10758), .ZN(n10654) );
  NAND2_X1 U13197 ( .A1(n12992), .A2(n10654), .ZN(n10655) );
  OAI211_X1 U13198 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n14761), .A(n10656), .B(
        n10655), .ZN(n10662) );
  NAND2_X1 U13199 ( .A1(n12996), .A2(n7779), .ZN(n12978) );
  INV_X1 U13200 ( .A(n10657), .ZN(n10658) );
  NOR4_X1 U13201 ( .A1(n12978), .A2(n10660), .A3(n10659), .A4(n10658), .ZN(
        n10661) );
  AOI211_X1 U13202 ( .C1(n12964), .C2(n10885), .A(n10662), .B(n10661), .ZN(
        n10663) );
  OAI21_X1 U13203 ( .B1(n10664), .B2(n12971), .A(n10663), .ZN(P2_U3202) );
  INV_X1 U13204 ( .A(n10665), .ZN(n10666) );
  OAI21_X1 U13205 ( .B1(n10666), .B2(n12971), .A(n12994), .ZN(n10669) );
  OR2_X1 U13206 ( .A1(n10667), .A2(P2_U3088), .ZN(n10855) );
  AOI22_X1 U13207 ( .A1(n10669), .A2(n10668), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n10855), .ZN(n10671) );
  NAND3_X1 U13208 ( .A1(n12953), .A2(n13030), .A3(n10696), .ZN(n10670) );
  OAI211_X1 U13209 ( .C1(n12961), .C2(n10672), .A(n10671), .B(n10670), .ZN(
        P2_U3204) );
  AOI21_X1 U13210 ( .B1(n10675), .B2(n10674), .A(n10673), .ZN(n10688) );
  NAND2_X1 U13211 ( .A1(n14932), .A2(n10676), .ZN(n10677) );
  XNOR2_X1 U13212 ( .A(n10678), .B(n10677), .ZN(n10681) );
  NOR2_X1 U13213 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10679), .ZN(n11179) );
  AOI21_X1 U13214 ( .B1(n14983), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n11179), .ZN(
        n10680) );
  OAI21_X1 U13215 ( .B1(n15015), .B2(n10681), .A(n10680), .ZN(n10686) );
  AOI21_X1 U13216 ( .B1(n15155), .B2(n10683), .A(n10682), .ZN(n10684) );
  NOR2_X1 U13217 ( .A1(n10684), .A2(n15017), .ZN(n10685) );
  AOI211_X1 U13218 ( .C1(n14960), .C2(n7079), .A(n10686), .B(n10685), .ZN(
        n10687) );
  OAI21_X1 U13219 ( .B1(n10688), .B2(n15023), .A(n10687), .ZN(P3_U3187) );
  INV_X1 U13220 ( .A(n10689), .ZN(n10692) );
  INV_X1 U13221 ( .A(n10695), .ZN(n10691) );
  INV_X1 U13222 ( .A(n10690), .ZN(n10851) );
  AOI21_X1 U13223 ( .B1(n10692), .B2(n10691), .A(n10851), .ZN(n10700) );
  OAI22_X1 U13224 ( .A1(n10694), .A2(n12994), .B1(n12961), .B2(n10693), .ZN(
        n10698) );
  NOR3_X1 U13225 ( .A1(n12978), .A2(n10696), .A3(n10695), .ZN(n10697) );
  AOI211_X1 U13226 ( .C1(P2_REG3_REG_1__SCAN_IN), .C2(n10855), .A(n10698), .B(
        n10697), .ZN(n10699) );
  OAI21_X1 U13227 ( .B1(n10700), .B2(n12971), .A(n10699), .ZN(P2_U3194) );
  OAI21_X1 U13228 ( .B1(n10703), .B2(n10702), .A(n10701), .ZN(n11024) );
  OAI211_X1 U13229 ( .C1(n10704), .C2(n11018), .A(n10756), .B(n13083), .ZN(
        n11019) );
  INV_X1 U13230 ( .A(n11019), .ZN(n10710) );
  XNOR2_X1 U13231 ( .A(n10706), .B(n10705), .ZN(n10708) );
  AOI21_X1 U13232 ( .B1(n10708), .B2(n14475), .A(n10707), .ZN(n11020) );
  INV_X1 U13233 ( .A(n11020), .ZN(n10709) );
  AOI211_X1 U13234 ( .C1(n14511), .C2(n11024), .A(n10710), .B(n10709), .ZN(
        n10714) );
  AOI22_X1 U13235 ( .A1(n13407), .A2(n10712), .B1(n14896), .B2(
        P2_REG0_REG_3__SCAN_IN), .ZN(n10711) );
  OAI21_X1 U13236 ( .B1(n10714), .B2(n14896), .A(n10711), .ZN(P2_U3439) );
  AOI22_X1 U13237 ( .A1(n13351), .A2(n10712), .B1(n14900), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n10713) );
  OAI21_X1 U13238 ( .B1(n10714), .B2(n14900), .A(n10713), .ZN(P2_U3502) );
  INV_X1 U13239 ( .A(n13551), .ZN(n10950) );
  INV_X1 U13240 ( .A(n13511), .ZN(n13549) );
  OAI22_X1 U13241 ( .A1(n11060), .A2(n10950), .B1(n13549), .B2(n11073), .ZN(
        n10715) );
  AOI21_X1 U13242 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n10716), .A(n10715), .ZN(
        n10721) );
  OAI21_X1 U13243 ( .B1(n7344), .B2(n10718), .A(n10717), .ZN(n10719) );
  NAND2_X1 U13244 ( .A1(n10719), .A2(n13537), .ZN(n10720) );
  OAI211_X1 U13245 ( .C1(n10631), .C2(n13526), .A(n10721), .B(n10720), .ZN(
        P1_U3222) );
  OAI222_X1 U13246 ( .A1(n12880), .A2(n10724), .B1(n12040), .B2(n10723), .C1(
        n10722), .C2(P3_U3151), .ZN(P3_U3278) );
  INV_X1 U13247 ( .A(n10725), .ZN(n10727) );
  NAND2_X1 U13248 ( .A1(n10727), .A2(n10726), .ZN(n10731) );
  OR2_X1 U13249 ( .A1(n6434), .A2(n11067), .ZN(n10729) );
  NAND2_X1 U13250 ( .A1(n6435), .A2(n14668), .ZN(n10728) );
  XNOR2_X1 U13251 ( .A(n10730), .B(n12122), .ZN(n10895) );
  XNOR2_X1 U13252 ( .A(n10895), .B(n10896), .ZN(n10732) );
  AOI21_X1 U13253 ( .B1(n10734), .B2(n10731), .A(n10732), .ZN(n10745) );
  AND2_X1 U13254 ( .A1(n10732), .A2(n10731), .ZN(n10733) );
  AND2_X1 U13255 ( .A1(n10596), .A2(n10735), .ZN(n10736) );
  NAND2_X1 U13256 ( .A1(n10737), .A2(n10736), .ZN(n10738) );
  AOI21_X2 U13257 ( .B1(n10738), .B2(P1_STATE_REG_SCAN_IN), .A(n9772), .ZN(
        n13553) );
  INV_X1 U13258 ( .A(n13553), .ZN(n13543) );
  OR2_X1 U13259 ( .A1(n11073), .A2(n13991), .ZN(n10740) );
  OR2_X1 U13260 ( .A1(n11077), .A2(n13993), .ZN(n10739) );
  NAND2_X1 U13261 ( .A1(n10740), .A2(n10739), .ZN(n11187) );
  AOI22_X1 U13262 ( .A1(n13475), .A2(n11187), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10741) );
  OAI21_X1 U13263 ( .B1(n13526), .B2(n11190), .A(n10741), .ZN(n10742) );
  AOI21_X1 U13264 ( .B1(n9266), .B2(n13543), .A(n10742), .ZN(n10743) );
  OAI21_X1 U13265 ( .B1(n10745), .B2(n10744), .A(n10743), .ZN(P1_U3218) );
  NAND2_X1 U13266 ( .A1(n10747), .A2(n10746), .ZN(n10749) );
  NAND2_X1 U13267 ( .A1(n13761), .A2(n11054), .ZN(n10750) );
  INV_X2 U13268 ( .A(n14731), .ZN(n14260) );
  INV_X1 U13269 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10753) );
  NAND2_X1 U13270 ( .A1(n14260), .A2(n10751), .ZN(n10752) );
  OAI21_X1 U13271 ( .B1(n14260), .B2(n10753), .A(n10752), .ZN(P1_U3459) );
  OAI21_X1 U13272 ( .B1(n10755), .B2(n10757), .A(n10754), .ZN(n10881) );
  AOI211_X1 U13273 ( .C1(n10761), .C2(n10756), .A(n7779), .B(n6759), .ZN(
        n10889) );
  OAI21_X1 U13274 ( .B1(n10759), .B2(n13279), .A(n10758), .ZN(n10882) );
  AOI211_X1 U13275 ( .C1(n14511), .C2(n10881), .A(n10889), .B(n10882), .ZN(
        n10763) );
  AOI22_X1 U13276 ( .A1(n13407), .A2(n10761), .B1(n14896), .B2(
        P2_REG0_REG_4__SCAN_IN), .ZN(n10760) );
  OAI21_X1 U13277 ( .B1(n10763), .B2(n14896), .A(n10760), .ZN(P2_U3442) );
  AOI22_X1 U13278 ( .A1(n13351), .A2(n10761), .B1(n14900), .B2(
        P2_REG1_REG_4__SCAN_IN), .ZN(n10762) );
  OAI21_X1 U13279 ( .B1(n10763), .B2(n14900), .A(n10762), .ZN(P2_U3503) );
  INV_X1 U13280 ( .A(n11095), .ZN(n10770) );
  OAI211_X1 U13281 ( .C1(n10765), .C2(n6568), .A(n11043), .B(n12996), .ZN(
        n10769) );
  AOI22_X1 U13282 ( .A1(n12986), .A2(n13026), .B1(n13024), .B2(n12946), .ZN(
        n10976) );
  OAI22_X1 U13283 ( .A1(n12961), .A2(n10976), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10766), .ZN(n10767) );
  AOI21_X1 U13284 ( .B1(n11096), .B2(n12976), .A(n10767), .ZN(n10768) );
  OAI211_X1 U13285 ( .C1(n12990), .C2(n10770), .A(n10769), .B(n10768), .ZN(
        P2_U3211) );
  NOR2_X1 U13286 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8456), .ZN(n14919) );
  OAI22_X1 U13287 ( .A1(n12434), .A2(n10772), .B1(n11176), .B2(n12421), .ZN(
        n10773) );
  AOI211_X1 U13288 ( .C1(n12418), .C2(n15078), .A(n14919), .B(n10773), .ZN(
        n10787) );
  XNOR2_X1 U13289 ( .A(n12284), .B(n15053), .ZN(n10777) );
  XNOR2_X1 U13290 ( .A(n10777), .B(n15078), .ZN(n10806) );
  NAND2_X1 U13291 ( .A1(n10777), .A2(n10776), .ZN(n10778) );
  NAND2_X1 U13292 ( .A1(n10779), .A2(n10778), .ZN(n10781) );
  XNOR2_X1 U13293 ( .A(n12284), .B(n10845), .ZN(n11006) );
  XNOR2_X1 U13294 ( .A(n11006), .B(n15060), .ZN(n10782) );
  AOI21_X1 U13295 ( .B1(n10781), .B2(n10782), .A(n12439), .ZN(n10785) );
  INV_X1 U13296 ( .A(n10781), .ZN(n10784) );
  NAND2_X1 U13297 ( .A1(n10785), .A2(n11009), .ZN(n10786) );
  OAI211_X1 U13298 ( .C1(n11810), .C2(P3_REG3_REG_3__SCAN_IN), .A(n10787), .B(
        n10786), .ZN(P3_U3158) );
  AOI21_X1 U13299 ( .B1(n11253), .B2(n10789), .A(n10788), .ZN(n10804) );
  AOI21_X1 U13300 ( .B1(n9082), .B2(n10791), .A(n10790), .ZN(n10792) );
  NOR2_X1 U13301 ( .A1(n10792), .A2(n15017), .ZN(n10802) );
  OR3_X1 U13302 ( .A1(n14930), .A2(n10794), .A3(n10793), .ZN(n10795) );
  AOI21_X1 U13303 ( .B1(n10796), .B2(n10795), .A(n15015), .ZN(n10801) );
  INV_X1 U13304 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n10797) );
  NOR2_X1 U13305 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10797), .ZN(n11391) );
  AOI21_X1 U13306 ( .B1(n14983), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n11391), .ZN(
        n10798) );
  OAI21_X1 U13307 ( .B1(n15008), .B2(n10799), .A(n10798), .ZN(n10800) );
  NOR3_X1 U13308 ( .A1(n10802), .A2(n10801), .A3(n10800), .ZN(n10803) );
  OAI21_X1 U13309 ( .B1(n10804), .B2(n15023), .A(n10803), .ZN(P3_U3189) );
  XOR2_X1 U13310 ( .A(n10805), .B(n10806), .Z(n10811) );
  OAI22_X1 U13311 ( .A1(n15062), .A2(n12433), .B1(n12421), .B2(n15060), .ZN(
        n10809) );
  NOR2_X1 U13312 ( .A1(n10807), .A2(n15055), .ZN(n10808) );
  AOI211_X1 U13313 ( .C1(n15053), .C2(n12424), .A(n10809), .B(n10808), .ZN(
        n10810) );
  OAI21_X1 U13314 ( .B1(n12439), .B2(n10811), .A(n10810), .ZN(P3_U3177) );
  INV_X1 U13315 ( .A(n10812), .ZN(n10815) );
  MUX2_X1 U13316 ( .A(n10815), .B(n10814), .S(n10813), .Z(n10816) );
  INV_X1 U13317 ( .A(n12744), .ZN(n12635) );
  AOI22_X1 U13318 ( .A1(n12635), .A2(n10818), .B1(n15090), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n10823) );
  MUX2_X1 U13319 ( .A(n10821), .B(n10820), .S(n15071), .Z(n10822) );
  NAND2_X1 U13320 ( .A1(n10823), .A2(n10822), .ZN(P3_U3233) );
  XNOR2_X1 U13321 ( .A(n10824), .B(n10828), .ZN(n10826) );
  OAI22_X1 U13322 ( .A1(n11377), .A2(n15059), .B1(n15060), .B2(n15061), .ZN(
        n10825) );
  AOI21_X1 U13323 ( .B1(n10826), .B2(n15074), .A(n10825), .ZN(n10831) );
  XNOR2_X1 U13325 ( .A(n10827), .B(n10828), .ZN(n15112) );
  NAND2_X1 U13326 ( .A1(n15112), .A2(n15083), .ZN(n10830) );
  AND2_X1 U13327 ( .A1(n10831), .A2(n10830), .ZN(n15114) );
  AND2_X1 U13328 ( .A1(n15054), .A2(n10832), .ZN(n15069) );
  AND2_X1 U13329 ( .A1(n11005), .A2(n15084), .ZN(n15111) );
  AOI22_X1 U13330 ( .A1(n15048), .A2(n15111), .B1(n15090), .B2(n11004), .ZN(
        n10833) );
  OAI21_X1 U13331 ( .B1(n9037), .B2(n15094), .A(n10833), .ZN(n10834) );
  AOI21_X1 U13332 ( .B1(n15091), .B2(n15112), .A(n10834), .ZN(n10835) );
  OAI21_X1 U13333 ( .B1(n15114), .B2(n15071), .A(n10835), .ZN(P3_U3229) );
  XNOR2_X1 U13334 ( .A(n10836), .B(n10838), .ZN(n15107) );
  INV_X1 U13335 ( .A(n15107), .ZN(n10848) );
  INV_X1 U13336 ( .A(n15091), .ZN(n11205) );
  NAND2_X1 U13337 ( .A1(n15107), .A2(n15083), .ZN(n10844) );
  AOI22_X1 U13338 ( .A1(n12450), .A2(n15079), .B1(n15076), .B2(n15078), .ZN(
        n10843) );
  NAND2_X1 U13339 ( .A1(n15057), .A2(n10837), .ZN(n10839) );
  NAND2_X1 U13340 ( .A1(n10839), .A2(n10838), .ZN(n10841) );
  NAND3_X1 U13341 ( .A1(n10841), .A2(n15074), .A3(n10840), .ZN(n10842) );
  AND3_X1 U13342 ( .A1(n10844), .A2(n10843), .A3(n10842), .ZN(n15109) );
  MUX2_X1 U13343 ( .A(n15109), .B(n14912), .S(n15071), .Z(n10847) );
  AND2_X1 U13344 ( .A1(n10845), .A2(n15084), .ZN(n15106) );
  AOI22_X1 U13345 ( .A1(n15048), .A2(n15106), .B1(n15090), .B2(n8456), .ZN(
        n10846) );
  OAI211_X1 U13346 ( .C1(n10848), .C2(n11205), .A(n10847), .B(n10846), .ZN(
        P3_U3230) );
  OAI22_X1 U13347 ( .A1(n10956), .A2(n12994), .B1(n12961), .B2(n10849), .ZN(
        n10854) );
  AOI22_X1 U13348 ( .A1(n12953), .A2(n6429), .B1(n12996), .B2(n7410), .ZN(
        n10852) );
  NOR3_X1 U13349 ( .A1(n10852), .A2(n10851), .A3(n10850), .ZN(n10853) );
  AOI211_X1 U13350 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(n10855), .A(n10854), .B(
        n10853), .ZN(n10856) );
  OAI21_X1 U13351 ( .B1(n10857), .B2(n12971), .A(n10856), .ZN(P2_U3209) );
  OAI21_X1 U13352 ( .B1(n10860), .B2(n10859), .A(n10858), .ZN(n10872) );
  AOI21_X1 U13353 ( .B1(n10861), .B2(n12171), .A(n7799), .ZN(n10862) );
  AND2_X1 U13354 ( .A1(n10973), .A2(n10862), .ZN(n10877) );
  XNOR2_X1 U13355 ( .A(n10864), .B(n10863), .ZN(n10865) );
  NAND2_X1 U13356 ( .A1(n10865), .A2(n14475), .ZN(n10868) );
  NAND2_X1 U13357 ( .A1(n13025), .A2(n12946), .ZN(n10867) );
  NAND2_X1 U13358 ( .A1(n13027), .A2(n12986), .ZN(n10866) );
  AND2_X1 U13359 ( .A1(n10867), .A2(n10866), .ZN(n12172) );
  NAND2_X1 U13360 ( .A1(n10868), .A2(n12172), .ZN(n10873) );
  AOI211_X1 U13361 ( .C1(n14511), .C2(n10872), .A(n10877), .B(n10873), .ZN(
        n10871) );
  AOI22_X1 U13362 ( .A1(n13351), .A2(n12171), .B1(n14900), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n10869) );
  OAI21_X1 U13363 ( .B1(n10871), .B2(n14900), .A(n10869), .ZN(P2_U3504) );
  AOI22_X1 U13364 ( .A1(n13407), .A2(n12171), .B1(n14896), .B2(
        P2_REG0_REG_5__SCAN_IN), .ZN(n10870) );
  OAI21_X1 U13365 ( .B1(n10871), .B2(n14896), .A(n10870), .ZN(P2_U3445) );
  INV_X1 U13366 ( .A(n10872), .ZN(n10880) );
  INV_X1 U13367 ( .A(n10873), .ZN(n10874) );
  MUX2_X1 U13368 ( .A(n10167), .B(n10874), .S(n14868), .Z(n10879) );
  INV_X1 U13369 ( .A(n12182), .ZN(n10875) );
  OAI22_X1 U13370 ( .A1(n14853), .A2(n6758), .B1(n10875), .B2(n14863), .ZN(
        n10876) );
  AOI21_X1 U13371 ( .B1(n14847), .B2(n10877), .A(n10876), .ZN(n10878) );
  OAI211_X1 U13372 ( .C1(n13254), .C2(n10880), .A(n10879), .B(n10878), .ZN(
        P2_U3260) );
  INV_X1 U13373 ( .A(n10881), .ZN(n10892) );
  INV_X1 U13374 ( .A(n10882), .ZN(n10883) );
  MUX2_X1 U13375 ( .A(n10884), .B(n10883), .S(n14868), .Z(n10891) );
  INV_X1 U13376 ( .A(n10885), .ZN(n10886) );
  OAI22_X1 U13377 ( .A1(n14853), .A2(n10887), .B1(n14863), .B2(n10886), .ZN(
        n10888) );
  AOI21_X1 U13378 ( .B1(n10889), .B2(n14847), .A(n10888), .ZN(n10890) );
  OAI211_X1 U13379 ( .C1(n13254), .C2(n10892), .A(n10891), .B(n10890), .ZN(
        P2_U3261) );
  INV_X1 U13380 ( .A(n11607), .ZN(n11350) );
  INV_X1 U13381 ( .A(n10893), .ZN(n10939) );
  OAI222_X1 U13382 ( .A1(P1_U3086), .A2(n11350), .B1(n14281), .B2(n10939), 
        .C1(n10894), .C2(n14278), .ZN(P1_U3340) );
  INV_X1 U13383 ( .A(n10895), .ZN(n10897) );
  NAND2_X1 U13384 ( .A1(n10897), .A2(n10896), .ZN(n10903) );
  NOR2_X1 U13385 ( .A1(n12162), .A2(n14680), .ZN(n10898) );
  AOI21_X1 U13386 ( .B1(n6594), .B2(n13570), .A(n10898), .ZN(n10904) );
  AND2_X1 U13387 ( .A1(n10903), .A2(n10904), .ZN(n10899) );
  OR2_X1 U13388 ( .A1(n12071), .A2(n11077), .ZN(n10901) );
  OAI21_X1 U13389 ( .B1(n10900), .B2(n14680), .A(n10901), .ZN(n10902) );
  XNOR2_X1 U13390 ( .A(n10902), .B(n12160), .ZN(n10948) );
  NAND2_X1 U13391 ( .A1(n10946), .A2(n10948), .ZN(n10907) );
  INV_X1 U13392 ( .A(n10904), .ZN(n10905) );
  INV_X1 U13393 ( .A(n13569), .ZN(n11292) );
  NAND2_X1 U13394 ( .A1(n10625), .A2(n11293), .ZN(n10908) );
  OAI21_X1 U13395 ( .B1(n12159), .B2(n11292), .A(n10908), .ZN(n10914) );
  INV_X1 U13396 ( .A(n10914), .ZN(n10913) );
  NAND2_X1 U13397 ( .A1(n6435), .A2(n11293), .ZN(n10910) );
  OR2_X1 U13398 ( .A1(n12071), .A2(n11292), .ZN(n10909) );
  NAND2_X1 U13399 ( .A1(n10910), .A2(n10909), .ZN(n10911) );
  XNOR2_X1 U13400 ( .A(n10911), .B(n12160), .ZN(n10915) );
  INV_X1 U13401 ( .A(n10915), .ZN(n10912) );
  NAND2_X1 U13402 ( .A1(n10913), .A2(n10912), .ZN(n11105) );
  AND2_X1 U13403 ( .A1(n10915), .A2(n10914), .ZN(n11106) );
  NOR2_X1 U13404 ( .A1(n6989), .A2(n11106), .ZN(n10916) );
  XNOR2_X1 U13405 ( .A(n11107), .B(n10916), .ZN(n10922) );
  NOR2_X1 U13406 ( .A1(n6819), .A2(n14726), .ZN(n14687) );
  OR2_X1 U13407 ( .A1(n11077), .A2(n13991), .ZN(n10918) );
  NAND2_X1 U13408 ( .A1(n13568), .A2(n13983), .ZN(n10917) );
  AND2_X1 U13409 ( .A1(n10918), .A2(n10917), .ZN(n11081) );
  NAND2_X1 U13410 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n13619) );
  OAI21_X1 U13411 ( .B1(n13540), .B2(n11081), .A(n13619), .ZN(n10920) );
  NOR2_X1 U13412 ( .A1(n13553), .A2(n11090), .ZN(n10919) );
  AOI211_X1 U13413 ( .C1(n13529), .C2(n14687), .A(n10920), .B(n10919), .ZN(
        n10921) );
  OAI21_X1 U13414 ( .B1(n10922), .B2(n13557), .A(n10921), .ZN(P1_U3227) );
  NOR2_X1 U13415 ( .A1(n10929), .A2(n10924), .ZN(n10925) );
  AOI21_X1 U13416 ( .B1(n10924), .B2(n10929), .A(n10925), .ZN(n14599) );
  NAND2_X1 U13417 ( .A1(n14600), .A2(n14599), .ZN(n14598) );
  OAI21_X1 U13418 ( .B1(n10924), .B2(n10929), .A(n14598), .ZN(n10927) );
  AOI22_X1 U13419 ( .A1(n11342), .A2(n9437), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n11347), .ZN(n10926) );
  NOR2_X1 U13420 ( .A1(n10926), .A2(n10927), .ZN(n11346) );
  AOI21_X1 U13421 ( .B1(n10927), .B2(n10926), .A(n11346), .ZN(n10938) );
  AOI22_X1 U13422 ( .A1(n11342), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n11839), 
        .B2(n11347), .ZN(n10934) );
  NAND2_X1 U13423 ( .A1(n14596), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n10932) );
  INV_X1 U13424 ( .A(n10932), .ZN(n10928) );
  AOI21_X1 U13425 ( .B1(n11719), .B2(n10929), .A(n10928), .ZN(n14604) );
  AOI21_X1 U13426 ( .B1(n10931), .B2(n11687), .A(n10930), .ZN(n14603) );
  NAND2_X1 U13427 ( .A1(n14604), .A2(n14603), .ZN(n14601) );
  NAND2_X1 U13428 ( .A1(n10932), .A2(n14601), .ZN(n10933) );
  NAND2_X1 U13429 ( .A1(n10934), .A2(n10933), .ZN(n11343) );
  OAI211_X1 U13430 ( .C1(n10934), .C2(n10933), .A(n14602), .B(n11343), .ZN(
        n10937) );
  INV_X1 U13431 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14316) );
  NAND2_X1 U13432 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n12008)
         );
  OAI21_X1 U13433 ( .B1(n14593), .B2(n14316), .A(n12008), .ZN(n10935) );
  AOI21_X1 U13434 ( .B1(n11342), .B2(n14595), .A(n10935), .ZN(n10936) );
  OAI211_X1 U13435 ( .C1(n10938), .C2(n13688), .A(n10937), .B(n10936), .ZN(
        P1_U3257) );
  INV_X1 U13436 ( .A(n14809), .ZN(n11400) );
  OAI222_X1 U13437 ( .A1(n13440), .A2(n10940), .B1(n11400), .B2(P2_U3088), 
        .C1(n13438), .C2(n10939), .ZN(P2_U3312) );
  INV_X1 U13438 ( .A(n10941), .ZN(n10944) );
  INV_X1 U13439 ( .A(SI_18_), .ZN(n10943) );
  OAI222_X1 U13440 ( .A1(n12880), .A2(n10944), .B1(n12040), .B2(n10943), .C1(
        n10942), .C2(P3_U3151), .ZN(P3_U3277) );
  NAND2_X1 U13441 ( .A1(n10945), .A2(n10946), .ZN(n10947) );
  XOR2_X1 U13442 ( .A(n10948), .B(n10947), .Z(n10954) );
  OAI22_X1 U13443 ( .A1(n10950), .A2(n11067), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10949), .ZN(n10952) );
  OAI22_X1 U13444 ( .A1(n13526), .A2(n14680), .B1(n13553), .B2(n11272), .ZN(
        n10951) );
  AOI211_X1 U13445 ( .C1(n13511), .C2(n13569), .A(n10952), .B(n10951), .ZN(
        n10953) );
  OAI21_X1 U13446 ( .B1(n10954), .B2(n13557), .A(n10953), .ZN(P1_U3230) );
  OAI22_X1 U13447 ( .A1(n14868), .A2(n7414), .B1(n10955), .B2(n14863), .ZN(
        n10958) );
  NOR2_X1 U13448 ( .A1(n14853), .A2(n10956), .ZN(n10957) );
  AOI211_X1 U13449 ( .C1(n10959), .C2(n14847), .A(n10958), .B(n10957), .ZN(
        n10962) );
  NAND2_X1 U13450 ( .A1(n14856), .A2(n10960), .ZN(n10961) );
  OAI211_X1 U13451 ( .C1(n14478), .C2(n10963), .A(n10962), .B(n10961), .ZN(
        P2_U3263) );
  AOI22_X1 U13452 ( .A1(n14847), .A2(n10965), .B1(n14868), .B2(n10964), .ZN(
        n10969) );
  INV_X1 U13453 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n14747) );
  OAI22_X1 U13454 ( .A1(n14868), .A2(n10134), .B1(n14747), .B2(n14863), .ZN(
        n10966) );
  AOI21_X1 U13455 ( .B1(n14479), .B2(n10967), .A(n10966), .ZN(n10968) );
  OAI211_X1 U13456 ( .C1(n13254), .C2(n10970), .A(n10969), .B(n10968), .ZN(
        P2_U3264) );
  OAI21_X1 U13457 ( .B1(n10972), .B2(n10974), .A(n10971), .ZN(n11102) );
  AOI211_X1 U13458 ( .C1(n11096), .C2(n10973), .A(n7779), .B(n11159), .ZN(
        n11094) );
  XNOR2_X1 U13459 ( .A(n10975), .B(n10974), .ZN(n10977) );
  OAI21_X1 U13460 ( .B1(n10977), .B2(n13279), .A(n10976), .ZN(n11099) );
  AOI211_X1 U13461 ( .C1(n14511), .C2(n11102), .A(n11094), .B(n11099), .ZN(
        n10980) );
  AOI22_X1 U13462 ( .A1(n13351), .A2(n11096), .B1(n14900), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n10978) );
  OAI21_X1 U13463 ( .B1(n10980), .B2(n14900), .A(n10978), .ZN(P2_U3505) );
  AOI22_X1 U13464 ( .A1(n13407), .A2(n11096), .B1(n14896), .B2(
        P2_REG0_REG_6__SCAN_IN), .ZN(n10979) );
  OAI21_X1 U13465 ( .B1(n10980), .B2(n14896), .A(n10979), .ZN(P2_U3448) );
  INV_X1 U13466 ( .A(n10981), .ZN(n11003) );
  INV_X1 U13467 ( .A(n14823), .ZN(n11406) );
  OAI222_X1 U13468 ( .A1(n13438), .A2(n11003), .B1(n11406), .B2(P2_U3088), 
        .C1(n10982), .C2(n13440), .ZN(P2_U3311) );
  INV_X1 U13469 ( .A(SI_19_), .ZN(n10983) );
  OAI222_X1 U13470 ( .A1(n12880), .A2(n10985), .B1(n10984), .B2(P3_U3151), 
        .C1(n10983), .C2(n12040), .ZN(P3_U3276) );
  AOI21_X1 U13471 ( .B1(n10988), .B2(n10987), .A(n10986), .ZN(n11002) );
  OAI21_X1 U13472 ( .B1(n10991), .B2(n10990), .A(n10989), .ZN(n11000) );
  AND2_X1 U13473 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n11571) );
  AOI21_X1 U13474 ( .B1(n14983), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n11571), .ZN(
        n10992) );
  OAI21_X1 U13475 ( .B1(n15008), .B2(n10993), .A(n10992), .ZN(n10999) );
  AOI21_X1 U13476 ( .B1(n10996), .B2(n10995), .A(n10994), .ZN(n10997) );
  NOR2_X1 U13477 ( .A1(n10997), .A2(n15017), .ZN(n10998) );
  AOI211_X1 U13478 ( .C1(n14963), .C2(n11000), .A(n10999), .B(n10998), .ZN(
        n11001) );
  OAI21_X1 U13479 ( .B1(n11002), .B2(n15023), .A(n11001), .ZN(P3_U3190) );
  INV_X1 U13480 ( .A(n11610), .ZN(n11696) );
  OAI222_X1 U13481 ( .A1(P1_U3086), .A2(n11696), .B1(n14281), .B2(n11003), 
        .C1(n14181), .C2(n14278), .ZN(P1_U3339) );
  INV_X1 U13482 ( .A(n11004), .ZN(n11017) );
  XNOR2_X1 U13483 ( .A(n12284), .B(n11005), .ZN(n11173) );
  XNOR2_X1 U13484 ( .A(n11173), .B(n12450), .ZN(n11010) );
  INV_X1 U13485 ( .A(n11006), .ZN(n11007) );
  NAND2_X1 U13486 ( .A1(n11007), .A2(n12451), .ZN(n11008) );
  OAI21_X1 U13487 ( .B1(n11010), .B2(n6574), .A(n11174), .ZN(n11011) );
  NAND2_X1 U13488 ( .A1(n11011), .A2(n12381), .ZN(n11016) );
  INV_X1 U13489 ( .A(n12421), .ZN(n12431) );
  OAI22_X1 U13490 ( .A1(n12434), .A2(n11012), .B1(n15060), .B2(n12433), .ZN(
        n11013) );
  AOI211_X1 U13491 ( .C1(n12431), .C2(n12449), .A(n11014), .B(n11013), .ZN(
        n11015) );
  OAI211_X1 U13492 ( .C1(n11017), .C2(n11810), .A(n11016), .B(n11015), .ZN(
        P3_U3170) );
  OAI22_X1 U13493 ( .A1(n13221), .A2(n11019), .B1(n11018), .B2(n14853), .ZN(
        n11023) );
  OAI21_X1 U13494 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n14863), .A(n11020), .ZN(
        n11021) );
  MUX2_X1 U13495 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n11021), .S(n14868), .Z(
        n11022) );
  AOI211_X1 U13496 ( .C1(n14856), .C2(n11024), .A(n11023), .B(n11022), .ZN(
        n11025) );
  INV_X1 U13497 ( .A(n11025), .ZN(P2_U3262) );
  INV_X1 U13498 ( .A(n11026), .ZN(n11027) );
  AOI21_X1 U13499 ( .B1(n11030), .B2(n11028), .A(n11027), .ZN(n11033) );
  AOI22_X1 U13500 ( .A1(n15076), .A2(n12450), .B1(n12448), .B2(n15079), .ZN(
        n11032) );
  XNOR2_X1 U13501 ( .A(n11029), .B(n11030), .ZN(n15118) );
  NAND2_X1 U13502 ( .A1(n15118), .A2(n15083), .ZN(n11031) );
  OAI211_X1 U13503 ( .C1(n11033), .C2(n12736), .A(n11032), .B(n11031), .ZN(
        n15116) );
  INV_X1 U13504 ( .A(n15116), .ZN(n11037) );
  NOR2_X1 U13505 ( .A1(n11177), .A2(n15130), .ZN(n15117) );
  AOI22_X1 U13506 ( .A1(n15048), .A2(n15117), .B1(n15090), .B2(n11180), .ZN(
        n11034) );
  OAI21_X1 U13507 ( .B1(n10675), .B2(n15094), .A(n11034), .ZN(n11035) );
  AOI21_X1 U13508 ( .B1(n15118), .B2(n15091), .A(n11035), .ZN(n11036) );
  OAI21_X1 U13509 ( .B1(n11037), .B2(n15071), .A(n11036), .ZN(P3_U3228) );
  INV_X1 U13510 ( .A(n14850), .ZN(n11041) );
  NAND2_X1 U13511 ( .A1(n13023), .A2(n12946), .ZN(n11039) );
  NAND2_X1 U13512 ( .A1(n13025), .A2(n12986), .ZN(n11038) );
  NAND2_X1 U13513 ( .A1(n11039), .A2(n11038), .ZN(n11164) );
  NAND2_X1 U13514 ( .A1(n12992), .A2(n11164), .ZN(n11040) );
  NAND2_X1 U13515 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n13045) );
  OAI211_X1 U13516 ( .C1(n12990), .C2(n11041), .A(n11040), .B(n13045), .ZN(
        n11050) );
  NAND3_X1 U13517 ( .A1(n12953), .A2(n13025), .A3(n11042), .ZN(n11048) );
  INV_X1 U13518 ( .A(n11043), .ZN(n11045) );
  OAI21_X1 U13519 ( .B1(n11045), .B2(n11044), .A(n12996), .ZN(n11047) );
  INV_X1 U13520 ( .A(n11046), .ZN(n12218) );
  AOI21_X1 U13521 ( .B1(n11048), .B2(n11047), .A(n12218), .ZN(n11049) );
  AOI211_X1 U13522 ( .C1(n11168), .C2(n12976), .A(n11050), .B(n11049), .ZN(
        n11051) );
  INV_X1 U13523 ( .A(n11051), .ZN(P2_U3185) );
  INV_X1 U13524 ( .A(n13762), .ZN(n11053) );
  NAND2_X1 U13525 ( .A1(n11053), .A2(n11052), .ZN(n11057) );
  INV_X1 U13526 ( .A(n11054), .ZN(n11055) );
  INV_X1 U13527 ( .A(n11131), .ZN(n11128) );
  INV_X1 U13528 ( .A(n11132), .ZN(n11061) );
  NAND2_X1 U13529 ( .A1(n9224), .A2(n10631), .ZN(n11062) );
  NAND2_X1 U13530 ( .A1(n14629), .A2(n11063), .ZN(n11065) );
  NAND2_X1 U13531 ( .A1(n11065), .A2(n11064), .ZN(n11184) );
  NAND2_X1 U13532 ( .A1(n11067), .A2(n11190), .ZN(n11068) );
  INV_X1 U13533 ( .A(n11069), .ZN(n11279) );
  NAND2_X1 U13534 ( .A1(n11274), .A2(n13570), .ZN(n11070) );
  NAND2_X1 U13535 ( .A1(n11275), .A2(n11070), .ZN(n11288) );
  XOR2_X1 U13536 ( .A(n11079), .B(n11288), .Z(n14684) );
  NAND2_X1 U13537 ( .A1(n9224), .A2(n11141), .ZN(n11072) );
  NAND2_X1 U13538 ( .A1(n11073), .A2(n14638), .ZN(n11074) );
  NAND2_X1 U13539 ( .A1(n11185), .A2(n11186), .ZN(n11076) );
  NOR2_X1 U13540 ( .A1(n13570), .A2(n14680), .ZN(n11078) );
  XNOR2_X1 U13541 ( .A(n11296), .B(n11079), .ZN(n11080) );
  NOR2_X1 U13542 ( .A1(n11080), .A2(n14077), .ZN(n14688) );
  INV_X1 U13543 ( .A(n11081), .ZN(n14685) );
  NOR2_X1 U13544 ( .A1(n14688), .A2(n14685), .ZN(n11082) );
  MUX2_X1 U13545 ( .A(n11083), .B(n11082), .S(n13962), .Z(n11093) );
  NAND2_X1 U13546 ( .A1(n13962), .A2(n11268), .ZN(n14643) );
  INV_X1 U13547 ( .A(n14637), .ZN(n11084) );
  INV_X1 U13548 ( .A(n14617), .ZN(n11087) );
  AOI211_X1 U13549 ( .C1(n11293), .C2(n11271), .A(n14636), .B(n11087), .ZN(
        n14686) );
  NOR2_X1 U13550 ( .A1(n9719), .A2(n11088), .ZN(n11089) );
  OAI22_X1 U13551 ( .A1(n14002), .A2(n6819), .B1(n13913), .B2(n11090), .ZN(
        n11091) );
  AOI21_X1 U13552 ( .B1(n14623), .B2(n14686), .A(n11091), .ZN(n11092) );
  OAI211_X1 U13553 ( .C1(n14008), .C2(n14684), .A(n11093), .B(n11092), .ZN(
        P1_U3288) );
  INV_X1 U13554 ( .A(n11094), .ZN(n11098) );
  AOI22_X1 U13555 ( .A1(n14479), .A2(n11096), .B1(n14849), .B2(n11095), .ZN(
        n11097) );
  OAI21_X1 U13556 ( .B1(n11098), .B2(n13221), .A(n11097), .ZN(n11101) );
  MUX2_X1 U13557 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11099), .S(n14868), .Z(
        n11100) );
  AOI211_X1 U13558 ( .C1(n14856), .C2(n11102), .A(n11101), .B(n11100), .ZN(
        n11103) );
  INV_X1 U13559 ( .A(n11103), .ZN(P2_U3259) );
  INV_X1 U13560 ( .A(n11104), .ZN(n11172) );
  INV_X1 U13561 ( .A(n11425), .ZN(n12231) );
  OAI222_X1 U13562 ( .A1(n13438), .A2(n11172), .B1(n12231), .B2(P2_U3088), 
        .C1(n14123), .C2(n13440), .ZN(P2_U3310) );
  NAND2_X1 U13563 ( .A1(n14616), .A2(n6435), .ZN(n11109) );
  INV_X1 U13564 ( .A(n13568), .ZN(n11297) );
  OR2_X1 U13565 ( .A1(n12162), .A2(n11297), .ZN(n11108) );
  NAND2_X1 U13566 ( .A1(n11109), .A2(n11108), .ZN(n11110) );
  XNOR2_X1 U13567 ( .A(n11110), .B(n12160), .ZN(n11116) );
  INV_X1 U13568 ( .A(n11116), .ZN(n11114) );
  NAND2_X1 U13569 ( .A1(n14616), .A2(n10625), .ZN(n11112) );
  NAND2_X1 U13570 ( .A1(n6594), .A2(n13568), .ZN(n11111) );
  NAND2_X1 U13571 ( .A1(n11112), .A2(n11111), .ZN(n11115) );
  INV_X1 U13572 ( .A(n11115), .ZN(n11113) );
  NAND2_X1 U13573 ( .A1(n11114), .A2(n11113), .ZN(n11214) );
  NAND2_X1 U13574 ( .A1(n11116), .A2(n11115), .ZN(n11212) );
  NAND2_X1 U13575 ( .A1(n11214), .A2(n11212), .ZN(n11117) );
  XNOR2_X1 U13576 ( .A(n11213), .B(n11117), .ZN(n11124) );
  AND2_X1 U13577 ( .A1(n14616), .A2(n14669), .ZN(n14692) );
  NAND2_X1 U13578 ( .A1(n13569), .A2(n13981), .ZN(n11119) );
  NAND2_X1 U13579 ( .A1(n13567), .A2(n13983), .ZN(n11118) );
  NAND2_X1 U13580 ( .A1(n11119), .A2(n11118), .ZN(n14691) );
  NAND2_X1 U13581 ( .A1(n13475), .A2(n14691), .ZN(n11120) );
  OAI211_X1 U13582 ( .C1(n13553), .C2(n14614), .A(n11121), .B(n11120), .ZN(
        n11122) );
  AOI21_X1 U13583 ( .B1(n13529), .B2(n14692), .A(n11122), .ZN(n11123) );
  OAI21_X1 U13584 ( .B1(n11124), .B2(n13557), .A(n11123), .ZN(P1_U3239) );
  NAND2_X1 U13585 ( .A1(n11141), .A2(n11125), .ZN(n11126) );
  NAND2_X1 U13586 ( .A1(n14637), .A2(n11126), .ZN(n11136) );
  XNOR2_X1 U13587 ( .A(n9224), .B(n11136), .ZN(n11127) );
  OAI21_X1 U13588 ( .B1(n11127), .B2(n14077), .A(n11060), .ZN(n11135) );
  OAI21_X1 U13589 ( .B1(n11128), .B2(n11060), .A(n14708), .ZN(n11129) );
  NAND2_X1 U13590 ( .A1(n11129), .A2(n13991), .ZN(n11134) );
  NAND2_X1 U13591 ( .A1(n11132), .A2(n11131), .ZN(n11133) );
  NAND2_X1 U13592 ( .A1(n11130), .A2(n11133), .ZN(n14657) );
  INV_X1 U13593 ( .A(n14703), .ZN(n14675) );
  AOI222_X1 U13594 ( .A1(n11135), .A2(n11134), .B1(n13572), .B2(n13983), .C1(
        n14657), .C2(n14675), .ZN(n14654) );
  NOR2_X1 U13595 ( .A1(n11136), .A2(n14636), .ZN(n14652) );
  INV_X1 U13596 ( .A(n11137), .ZN(n11138) );
  NAND2_X1 U13597 ( .A1(n13962), .A2(n11138), .ZN(n14641) );
  INV_X1 U13598 ( .A(n14641), .ZN(n14624) );
  AOI22_X1 U13599 ( .A1(n14623), .A2(n14652), .B1(n14624), .B2(n14657), .ZN(
        n11143) );
  OAI22_X1 U13600 ( .A1(n13962), .A2(n14202), .B1(n11139), .B2(n13913), .ZN(
        n11140) );
  AOI21_X1 U13601 ( .B1(n14634), .B2(n11141), .A(n11140), .ZN(n11142) );
  OAI211_X1 U13602 ( .C1(n14647), .C2(n14654), .A(n11143), .B(n11142), .ZN(
        P1_U3292) );
  INV_X1 U13603 ( .A(n11332), .ZN(n11147) );
  OAI22_X1 U13604 ( .A1(n11144), .A2(n12967), .B1(n12200), .B2(n12984), .ZN(
        n11328) );
  NAND2_X1 U13605 ( .A1(n12992), .A2(n11328), .ZN(n11146) );
  OAI211_X1 U13606 ( .C1(n12990), .C2(n11147), .A(n11146), .B(n11145), .ZN(
        n11153) );
  INV_X1 U13607 ( .A(n12224), .ZN(n11151) );
  AOI22_X1 U13608 ( .A1(n11148), .A2(n12996), .B1(n12953), .B2(n13023), .ZN(
        n11150) );
  NOR3_X1 U13609 ( .A1(n11151), .A2(n11150), .A3(n11149), .ZN(n11152) );
  AOI211_X1 U13610 ( .C1(n11543), .C2(n12976), .A(n11153), .B(n11152), .ZN(
        n11154) );
  OAI21_X1 U13611 ( .B1(n11155), .B2(n12971), .A(n11154), .ZN(P2_U3203) );
  OAI21_X1 U13612 ( .B1(n11158), .B2(n11157), .A(n11156), .ZN(n14855) );
  INV_X1 U13613 ( .A(n11159), .ZN(n11161) );
  INV_X1 U13614 ( .A(n11239), .ZN(n11160) );
  AOI211_X1 U13615 ( .C1(n11168), .C2(n11161), .A(n7779), .B(n11160), .ZN(
        n14848) );
  XNOR2_X1 U13616 ( .A(n11163), .B(n11162), .ZN(n11165) );
  AOI21_X1 U13617 ( .B1(n11165), .B2(n14475), .A(n11164), .ZN(n14858) );
  INV_X1 U13618 ( .A(n14858), .ZN(n11166) );
  AOI211_X1 U13619 ( .C1(n14511), .C2(n14855), .A(n14848), .B(n11166), .ZN(
        n11170) );
  AOI22_X1 U13620 ( .A1(n13351), .A2(n11168), .B1(n14900), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n11167) );
  OAI21_X1 U13621 ( .B1(n11170), .B2(n14900), .A(n11167), .ZN(P2_U3506) );
  AOI22_X1 U13622 ( .A1(n13407), .A2(n11168), .B1(n14896), .B2(
        P2_REG0_REG_7__SCAN_IN), .ZN(n11169) );
  OAI21_X1 U13623 ( .B1(n11170), .B2(n14896), .A(n11169), .ZN(P2_U3451) );
  INV_X1 U13624 ( .A(n11704), .ZN(n13668) );
  OAI222_X1 U13625 ( .A1(P1_U3086), .A2(n13668), .B1(n14281), .B2(n11172), 
        .C1(n11171), .C2(n14278), .ZN(P1_U3338) );
  XNOR2_X1 U13626 ( .A(n12284), .B(n11175), .ZN(n11378) );
  XOR2_X1 U13627 ( .A(n11376), .B(n11375), .Z(n11183) );
  OAI22_X1 U13628 ( .A1(n12434), .A2(n11177), .B1(n11176), .B2(n12433), .ZN(
        n11178) );
  AOI211_X1 U13629 ( .C1(n12431), .C2(n12448), .A(n11179), .B(n11178), .ZN(
        n11182) );
  NAND2_X1 U13630 ( .A1(n12437), .A2(n11180), .ZN(n11181) );
  OAI211_X1 U13631 ( .C1(n11183), .C2(n12439), .A(n11182), .B(n11181), .ZN(
        P3_U3167) );
  XNOR2_X1 U13632 ( .A(n11186), .B(n11184), .ZN(n14672) );
  AOI211_X1 U13633 ( .C1(n14668), .C2(n14639), .A(n14636), .B(n6571), .ZN(
        n14667) );
  XNOR2_X1 U13634 ( .A(n11186), .B(n11185), .ZN(n11188) );
  AOI21_X1 U13635 ( .B1(n11188), .B2(n14708), .A(n11187), .ZN(n14670) );
  NOR2_X1 U13636 ( .A1(n14670), .A2(n14647), .ZN(n11192) );
  INV_X1 U13637 ( .A(n13913), .ZN(n14635) );
  AOI22_X1 U13638 ( .A1(n14647), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n14635), 
        .B2(n9266), .ZN(n11189) );
  OAI21_X1 U13639 ( .B1(n14002), .B2(n11190), .A(n11189), .ZN(n11191) );
  AOI211_X1 U13640 ( .C1(n14667), .C2(n14623), .A(n11192), .B(n11191), .ZN(
        n11193) );
  OAI21_X1 U13641 ( .B1(n14008), .B2(n14672), .A(n11193), .ZN(P1_U3290) );
  XNOR2_X1 U13642 ( .A(n11194), .B(n11198), .ZN(n15120) );
  OAI22_X1 U13643 ( .A1(n11377), .A2(n15061), .B1(n11569), .B2(n15059), .ZN(
        n11195) );
  INV_X1 U13644 ( .A(n11195), .ZN(n11201) );
  AND2_X1 U13645 ( .A1(n11026), .A2(n11196), .ZN(n11199) );
  OAI211_X1 U13646 ( .C1(n11199), .C2(n11198), .A(n11197), .B(n15074), .ZN(
        n11200) );
  OAI211_X1 U13647 ( .C1(n15120), .C2(n15067), .A(n11201), .B(n11200), .ZN(
        n15121) );
  INV_X1 U13648 ( .A(n15121), .ZN(n11202) );
  MUX2_X1 U13649 ( .A(n9042), .B(n11202), .S(n15094), .Z(n11204) );
  AND2_X1 U13650 ( .A1(n11521), .A2(n15084), .ZN(n15122) );
  AOI22_X1 U13651 ( .A1(n15048), .A2(n15122), .B1(n15090), .B2(n11529), .ZN(
        n11203) );
  OAI211_X1 U13652 ( .C1(n15120), .C2(n11205), .A(n11204), .B(n11203), .ZN(
        P3_U3227) );
  INV_X1 U13653 ( .A(n13683), .ZN(n13676) );
  INV_X1 U13654 ( .A(n11206), .ZN(n11224) );
  OAI222_X1 U13655 ( .A1(P1_U3086), .A2(n13676), .B1(n14281), .B2(n11224), 
        .C1(n11207), .C2(n14278), .ZN(P1_U3337) );
  INV_X1 U13656 ( .A(n11208), .ZN(n11209) );
  OAI222_X1 U13657 ( .A1(P3_U3151), .A2(n11211), .B1(n12040), .B2(n11210), 
        .C1(n12880), .C2(n11209), .ZN(P3_U3275) );
  NAND2_X1 U13658 ( .A1(n11517), .A2(n6435), .ZN(n11216) );
  INV_X1 U13659 ( .A(n13567), .ZN(n11300) );
  OR2_X1 U13660 ( .A1(n12071), .A2(n11300), .ZN(n11215) );
  NAND2_X1 U13661 ( .A1(n11216), .A2(n11215), .ZN(n11217) );
  XNOR2_X1 U13662 ( .A(n11217), .B(n12122), .ZN(n11457) );
  NOR2_X1 U13663 ( .A1(n12159), .A2(n11300), .ZN(n11218) );
  AOI21_X1 U13664 ( .B1(n11517), .B2(n10625), .A(n11218), .ZN(n11458) );
  XNOR2_X1 U13665 ( .A(n11457), .B(n11458), .ZN(n11462) );
  XNOR2_X1 U13666 ( .A(n11463), .B(n11462), .ZN(n11223) );
  AOI22_X1 U13667 ( .A1(n13981), .A2(n13568), .B1(n13566), .B2(n13983), .ZN(
        n14699) );
  INV_X1 U13668 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n11219) );
  OAI22_X1 U13669 ( .A1(n13540), .A2(n14699), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11219), .ZN(n11221) );
  NOR2_X1 U13670 ( .A1(n13553), .A2(n11515), .ZN(n11220) );
  AOI211_X1 U13671 ( .C1(n13555), .C2(n11517), .A(n11221), .B(n11220), .ZN(
        n11222) );
  OAI21_X1 U13672 ( .B1(n11223), .B2(n13557), .A(n11222), .ZN(P1_U3213) );
  INV_X1 U13673 ( .A(n14842), .ZN(n11225) );
  OAI222_X1 U13674 ( .A1(n13440), .A2(n14112), .B1(n11225), .B2(P2_U3088), 
        .C1(n13438), .C2(n11224), .ZN(P2_U3309) );
  NAND2_X1 U13675 ( .A1(n11227), .A2(n11226), .ZN(n11228) );
  NAND2_X1 U13676 ( .A1(n11229), .A2(n11228), .ZN(n11237) );
  OR2_X1 U13677 ( .A1(n11237), .A2(n9954), .ZN(n11236) );
  XNOR2_X1 U13678 ( .A(n11230), .B(n11231), .ZN(n11234) );
  NAND2_X1 U13679 ( .A1(n13022), .A2(n12946), .ZN(n11233) );
  NAND2_X1 U13680 ( .A1(n13024), .A2(n12986), .ZN(n11232) );
  NAND2_X1 U13681 ( .A1(n11233), .A2(n11232), .ZN(n12211) );
  AOI21_X1 U13682 ( .B1(n11234), .B2(n14475), .A(n12211), .ZN(n11235) );
  INV_X1 U13683 ( .A(n11237), .ZN(n14885) );
  INV_X1 U13684 ( .A(n11238), .ZN(n14866) );
  AND2_X1 U13685 ( .A1(n14868), .A2(n14866), .ZN(n11630) );
  AOI21_X1 U13686 ( .B1(n11239), .B2(n14881), .A(n7799), .ZN(n11240) );
  NAND2_X1 U13687 ( .A1(n11240), .A2(n11331), .ZN(n14882) );
  AOI22_X1 U13688 ( .A1(n14478), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n11241), 
        .B2(n14849), .ZN(n11243) );
  NAND2_X1 U13689 ( .A1(n14479), .A2(n14881), .ZN(n11242) );
  OAI211_X1 U13690 ( .C1(n14882), .C2(n13221), .A(n11243), .B(n11242), .ZN(
        n11244) );
  AOI21_X1 U13691 ( .B1(n14885), .B2(n11630), .A(n11244), .ZN(n11245) );
  OAI21_X1 U13692 ( .B1(n14887), .B2(n14478), .A(n11245), .ZN(P2_U3257) );
  XNOR2_X1 U13693 ( .A(n11246), .B(n11387), .ZN(n11252) );
  XNOR2_X1 U13694 ( .A(n11248), .B(n11247), .ZN(n11250) );
  OAI22_X1 U13695 ( .A1(n11389), .A2(n15061), .B1(n11566), .B2(n15059), .ZN(
        n11249) );
  AOI21_X1 U13696 ( .B1(n11250), .B2(n15074), .A(n11249), .ZN(n11251) );
  OAI21_X1 U13697 ( .B1(n11252), .B2(n15067), .A(n11251), .ZN(n15126) );
  AOI21_X1 U13698 ( .B1(n15090), .B2(n11374), .A(n15126), .ZN(n11256) );
  INV_X1 U13699 ( .A(n11252), .ZN(n15128) );
  OAI22_X1 U13700 ( .A1(n12744), .A2(n15125), .B1(n11253), .B2(n15094), .ZN(
        n11254) );
  AOI21_X1 U13701 ( .B1(n15128), .B2(n15091), .A(n11254), .ZN(n11255) );
  OAI21_X1 U13702 ( .B1(n11256), .B2(n15071), .A(n11255), .ZN(P3_U3226) );
  AOI21_X1 U13703 ( .B1(n11257), .B2(n13962), .A(n14623), .ZN(n11262) );
  AOI22_X1 U13704 ( .A1(n14647), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n14635), .ZN(n11260) );
  NOR2_X1 U13705 ( .A1(n14647), .A2(n14077), .ZN(n13869) );
  OAI21_X1 U13706 ( .B1(n13967), .B2(n13869), .A(n11258), .ZN(n11259) );
  OAI211_X1 U13707 ( .C1(n11262), .C2(n11261), .A(n11260), .B(n11259), .ZN(
        P1_U3293) );
  NAND2_X1 U13708 ( .A1(n12443), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n11263) );
  OAI21_X1 U13709 ( .B1(n12327), .B2(n12443), .A(n11263), .ZN(P3_U3520) );
  INV_X1 U13710 ( .A(n11264), .ZN(n11267) );
  OAI222_X1 U13711 ( .A1(n13440), .A2(n11265), .B1(n13438), .B2(n11267), .C1(
        P2_U3088), .C2(n12239), .ZN(P2_U3308) );
  OAI222_X1 U13712 ( .A1(P1_U3086), .A2(n11268), .B1(n14281), .B2(n11267), 
        .C1(n11266), .C2(n14278), .ZN(P1_U3336) );
  INV_X1 U13713 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n14163) );
  NAND2_X1 U13714 ( .A1(n11269), .A2(P3_U3897), .ZN(n11270) );
  OAI21_X1 U13715 ( .B1(P3_U3897), .B2(n14163), .A(n11270), .ZN(P3_U3522) );
  OAI211_X1 U13716 ( .C1(n6571), .C2(n14680), .A(n11271), .B(n14618), .ZN(
        n14678) );
  INV_X1 U13717 ( .A(n11272), .ZN(n11273) );
  AOI22_X1 U13718 ( .A1(n14634), .A2(n11274), .B1(n14635), .B2(n11273), .ZN(
        n11278) );
  NAND2_X1 U13719 ( .A1(n11276), .A2(n11279), .ZN(n14677) );
  NAND3_X1 U13720 ( .A1(n13967), .A2(n11275), .A3(n14677), .ZN(n11277) );
  OAI211_X1 U13721 ( .C1(n14643), .C2(n14678), .A(n11278), .B(n11277), .ZN(
        n11285) );
  XNOR2_X1 U13722 ( .A(n11280), .B(n11279), .ZN(n11281) );
  NAND2_X1 U13723 ( .A1(n11281), .A2(n14708), .ZN(n11283) );
  AOI22_X1 U13724 ( .A1(n13981), .A2(n13571), .B1(n13569), .B2(n13983), .ZN(
        n11282) );
  NAND2_X1 U13725 ( .A1(n11283), .A2(n11282), .ZN(n14681) );
  MUX2_X1 U13726 ( .A(n14681), .B(P1_REG2_REG_4__SCAN_IN), .S(n14647), .Z(
        n11284) );
  OR2_X1 U13727 ( .A1(n11285), .A2(n11284), .ZN(P1_U3289) );
  NAND2_X1 U13728 ( .A1(n6819), .A2(n11292), .ZN(n11287) );
  AND2_X1 U13729 ( .A1(n11293), .A2(n13569), .ZN(n11286) );
  AOI21_X1 U13730 ( .B1(n11288), .B2(n11287), .A(n11286), .ZN(n14610) );
  INV_X1 U13731 ( .A(n14611), .ZN(n14609) );
  NAND2_X1 U13732 ( .A1(n14610), .A2(n14609), .ZN(n14608) );
  OR2_X1 U13733 ( .A1(n14616), .A2(n13568), .ZN(n11289) );
  NAND2_X1 U13734 ( .A1(n14608), .A2(n11289), .ZN(n11507) );
  INV_X1 U13735 ( .A(n11509), .ZN(n11506) );
  OR2_X1 U13736 ( .A1(n11517), .A2(n13567), .ZN(n11290) );
  NAND2_X1 U13737 ( .A1(n11469), .A2(n13566), .ZN(n11291) );
  XNOR2_X1 U13738 ( .A(n11430), .B(n11438), .ZN(n14717) );
  NOR2_X1 U13739 ( .A1(n11293), .A2(n11292), .ZN(n11295) );
  NAND2_X1 U13740 ( .A1(n11293), .A2(n11292), .ZN(n11294) );
  NAND2_X1 U13741 ( .A1(n14616), .A2(n11297), .ZN(n11298) );
  AND2_X1 U13742 ( .A1(n11517), .A2(n11300), .ZN(n11302) );
  OR2_X1 U13743 ( .A1(n11517), .A2(n11300), .ZN(n11301) );
  INV_X1 U13744 ( .A(n11365), .ZN(n11303) );
  XNOR2_X1 U13745 ( .A(n11439), .B(n11438), .ZN(n11305) );
  OAI22_X1 U13746 ( .A1(n11763), .A2(n13993), .B1(n11467), .B2(n13991), .ZN(
        n11304) );
  AOI21_X1 U13747 ( .B1(n11305), .B2(n14708), .A(n11304), .ZN(n11306) );
  OAI21_X1 U13748 ( .B1(n14717), .B2(n14703), .A(n11306), .ZN(n14719) );
  NAND2_X1 U13749 ( .A1(n14719), .A2(n13962), .ZN(n11312) );
  OAI22_X1 U13750 ( .A1(n13962), .A2(n11307), .B1(n11592), .B2(n13913), .ZN(
        n11310) );
  INV_X1 U13751 ( .A(n11469), .ZN(n11481) );
  INV_X1 U13752 ( .A(n11517), .ZN(n14701) );
  NOR2_X1 U13753 ( .A1(n14617), .A2(n14616), .ZN(n14620) );
  INV_X1 U13754 ( .A(n11362), .ZN(n11308) );
  OAI211_X1 U13755 ( .C1(n6828), .C2(n11308), .A(n14618), .B(n11434), .ZN(
        n14718) );
  NOR2_X1 U13756 ( .A1(n14718), .A2(n14643), .ZN(n11309) );
  AOI211_X1 U13757 ( .C1(n14634), .C2(n11594), .A(n11310), .B(n11309), .ZN(
        n11311) );
  OAI211_X1 U13758 ( .C1(n14717), .C2(n14641), .A(n11312), .B(n11311), .ZN(
        P1_U3284) );
  INV_X1 U13759 ( .A(n11313), .ZN(n11314) );
  AOI21_X1 U13760 ( .B1(n11317), .B2(n11315), .A(n11314), .ZN(n11320) );
  AOI22_X1 U13761 ( .A1(n11562), .A2(n15076), .B1(n15079), .B2(n11807), .ZN(
        n11319) );
  XNOR2_X1 U13762 ( .A(n11316), .B(n11317), .ZN(n15134) );
  NAND2_X1 U13763 ( .A1(n15134), .A2(n15083), .ZN(n11318) );
  OAI211_X1 U13764 ( .C1(n11320), .C2(n12736), .A(n11319), .B(n11318), .ZN(
        n15132) );
  INV_X1 U13765 ( .A(n15132), .ZN(n11324) );
  AOI22_X1 U13766 ( .A1(n15071), .A2(P3_REG2_REG_8__SCAN_IN), .B1(n15090), 
        .B2(n11560), .ZN(n11321) );
  OAI21_X1 U13767 ( .B1(n12744), .B2(n15131), .A(n11321), .ZN(n11322) );
  AOI21_X1 U13768 ( .B1(n15134), .B2(n15091), .A(n11322), .ZN(n11323) );
  OAI21_X1 U13769 ( .B1(n11324), .B2(n15071), .A(n11323), .ZN(P3_U3225) );
  XNOR2_X1 U13770 ( .A(n11325), .B(n11327), .ZN(n11536) );
  INV_X1 U13771 ( .A(n11630), .ZN(n11338) );
  XNOR2_X1 U13772 ( .A(n11326), .B(n11327), .ZN(n11329) );
  AOI21_X1 U13773 ( .B1(n11329), .B2(n14475), .A(n11328), .ZN(n11330) );
  OAI21_X1 U13774 ( .B1(n11536), .B2(n9954), .A(n11330), .ZN(n11537) );
  NAND2_X1 U13775 ( .A1(n11537), .A2(n14868), .ZN(n11337) );
  AOI211_X1 U13776 ( .C1(n11543), .C2(n11331), .A(n7799), .B(n11497), .ZN(
        n11538) );
  INV_X1 U13777 ( .A(n11543), .ZN(n11334) );
  AOI22_X1 U13778 ( .A1(n14478), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n11332), 
        .B2(n14849), .ZN(n11333) );
  OAI21_X1 U13779 ( .B1(n11334), .B2(n14853), .A(n11333), .ZN(n11335) );
  AOI21_X1 U13780 ( .B1(n11538), .B2(n14847), .A(n11335), .ZN(n11336) );
  OAI211_X1 U13781 ( .C1(n11536), .C2(n11338), .A(n11337), .B(n11336), .ZN(
        P2_U3256) );
  OAI22_X1 U13782 ( .A1(n11339), .A2(P3_U3151), .B1(SI_22_), .B2(n12040), .ZN(
        n11340) );
  AOI21_X1 U13783 ( .B1(n11341), .B2(n12872), .A(n11340), .ZN(P3_U3273) );
  NAND2_X1 U13784 ( .A1(n11342), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11344) );
  NAND2_X1 U13785 ( .A1(n11344), .A2(n11343), .ZN(n11599) );
  XOR2_X1 U13786 ( .A(n11599), .B(n11350), .Z(n11345) );
  NOR2_X1 U13787 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n11345), .ZN(n11600) );
  AOI21_X1 U13788 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n11345), .A(n11600), 
        .ZN(n11356) );
  AOI21_X1 U13789 ( .B1(n11347), .B2(n9437), .A(n11346), .ZN(n11606) );
  XOR2_X1 U13790 ( .A(n11350), .B(n11606), .Z(n11348) );
  NOR2_X1 U13791 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n11348), .ZN(n11608) );
  AOI21_X1 U13792 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n11348), .A(n11608), 
        .ZN(n11349) );
  OR2_X1 U13793 ( .A1(n11349), .A2(n13688), .ZN(n11354) );
  NOR2_X1 U13794 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14183), .ZN(n11352) );
  NOR2_X1 U13795 ( .A1(n13677), .A2(n11350), .ZN(n11351) );
  AOI211_X1 U13796 ( .C1(n14578), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n11352), 
        .B(n11351), .ZN(n11353) );
  OAI211_X1 U13797 ( .C1(n11356), .C2(n11355), .A(n11354), .B(n11353), .ZN(
        P1_U3258) );
  INV_X1 U13798 ( .A(n11357), .ZN(n11358) );
  OAI222_X1 U13799 ( .A1(P3_U3151), .A2(n11360), .B1(n12040), .B2(n11359), 
        .C1(n12880), .C2(n11358), .ZN(P3_U3274) );
  XNOR2_X1 U13800 ( .A(n11361), .B(n11365), .ZN(n14716) );
  OAI211_X1 U13801 ( .C1(n11481), .C2(n11511), .A(n14618), .B(n11362), .ZN(
        n14712) );
  INV_X1 U13802 ( .A(n11485), .ZN(n11363) );
  AOI22_X1 U13803 ( .A1(n14634), .A2(n11469), .B1(n14635), .B2(n11363), .ZN(
        n11364) );
  OAI21_X1 U13804 ( .B1(n14643), .B2(n14712), .A(n11364), .ZN(n11372) );
  XNOR2_X1 U13805 ( .A(n11366), .B(n11365), .ZN(n11367) );
  NAND2_X1 U13806 ( .A1(n11367), .A2(n14708), .ZN(n14714) );
  NAND2_X1 U13807 ( .A1(n13567), .A2(n13981), .ZN(n11369) );
  NAND2_X1 U13808 ( .A1(n13565), .A2(n13983), .ZN(n11368) );
  NAND2_X1 U13809 ( .A1(n11369), .A2(n11368), .ZN(n11482) );
  INV_X1 U13810 ( .A(n11482), .ZN(n14713) );
  NAND2_X1 U13811 ( .A1(n14714), .A2(n14713), .ZN(n11370) );
  MUX2_X1 U13812 ( .A(n11370), .B(P1_REG2_REG_8__SCAN_IN), .S(n14647), .Z(
        n11371) );
  AOI211_X1 U13813 ( .C1(n13967), .C2(n14716), .A(n11372), .B(n11371), .ZN(
        n11373) );
  INV_X1 U13814 ( .A(n11373), .ZN(P1_U3285) );
  INV_X1 U13815 ( .A(n11374), .ZN(n11394) );
  NAND2_X1 U13816 ( .A1(n11376), .A2(n11375), .ZN(n11380) );
  NAND2_X1 U13817 ( .A1(n11378), .A2(n11377), .ZN(n11379) );
  NAND2_X1 U13818 ( .A1(n11380), .A2(n11379), .ZN(n11525) );
  INV_X1 U13819 ( .A(n11525), .ZN(n11383) );
  XNOR2_X1 U13820 ( .A(n12284), .B(n11381), .ZN(n11384) );
  XNOR2_X1 U13821 ( .A(n11384), .B(n12448), .ZN(n11526) );
  NAND2_X1 U13822 ( .A1(n11383), .A2(n11382), .ZN(n11523) );
  NAND2_X1 U13823 ( .A1(n11384), .A2(n12448), .ZN(n11385) );
  NAND2_X1 U13824 ( .A1(n11523), .A2(n11385), .ZN(n11388) );
  XNOR2_X1 U13825 ( .A(n11387), .B(n11386), .ZN(n11561) );
  NAND2_X1 U13826 ( .A1(n11388), .A2(n11561), .ZN(n11565) );
  OAI211_X1 U13827 ( .C1(n11388), .C2(n11561), .A(n11565), .B(n12381), .ZN(
        n11393) );
  OAI22_X1 U13828 ( .A1(n12434), .A2(n15125), .B1(n11389), .B2(n12433), .ZN(
        n11390) );
  AOI211_X1 U13829 ( .C1(n12431), .C2(n15040), .A(n11391), .B(n11390), .ZN(
        n11392) );
  OAI211_X1 U13830 ( .C1(n11394), .C2(n11810), .A(n11393), .B(n11392), .ZN(
        P3_U3153) );
  INV_X1 U13831 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13367) );
  AOI22_X1 U13832 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n11425), .B1(n12231), 
        .B2(n13367), .ZN(n11404) );
  INV_X1 U13833 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n13372) );
  XNOR2_X1 U13834 ( .A(n14823), .B(n13372), .ZN(n14827) );
  INV_X1 U13835 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n14500) );
  OR2_X1 U13836 ( .A1(n14801), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n11396) );
  NAND2_X1 U13837 ( .A1(n14801), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n11395) );
  AND2_X1 U13838 ( .A1(n11396), .A2(n11395), .ZN(n14804) );
  INV_X1 U13839 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n14505) );
  AOI21_X1 U13840 ( .B1(n14512), .B2(n11411), .A(n11397), .ZN(n14790) );
  NOR2_X1 U13841 ( .A1(n11412), .A2(n14505), .ZN(n11398) );
  AOI21_X1 U13842 ( .B1(n14505), .B2(n11412), .A(n11398), .ZN(n14789) );
  NAND2_X1 U13843 ( .A1(n14790), .A2(n14789), .ZN(n14788) );
  OAI21_X1 U13844 ( .B1(n11412), .B2(n14505), .A(n14788), .ZN(n14803) );
  NAND2_X1 U13845 ( .A1(n14804), .A2(n14803), .ZN(n14802) );
  OAI21_X1 U13846 ( .B1(n11415), .B2(n14500), .A(n14802), .ZN(n11399) );
  XNOR2_X1 U13847 ( .A(n11399), .B(n14809), .ZN(n14812) );
  INV_X1 U13848 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n11402) );
  INV_X1 U13849 ( .A(n11399), .ZN(n11401) );
  OAI22_X1 U13850 ( .A1(n14812), .A2(n11402), .B1(n11401), .B2(n11400), .ZN(
        n14826) );
  NAND2_X1 U13851 ( .A1(n14827), .A2(n14826), .ZN(n14824) );
  OAI21_X1 U13852 ( .B1(n11406), .B2(n13372), .A(n14824), .ZN(n11403) );
  NAND2_X1 U13853 ( .A1(n11404), .A2(n11403), .ZN(n12230) );
  OAI21_X1 U13854 ( .B1(n11404), .B2(n11403), .A(n12230), .ZN(n11428) );
  NAND2_X1 U13855 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n14823), .ZN(n11419) );
  INV_X1 U13856 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11407) );
  INV_X1 U13857 ( .A(n11419), .ZN(n11405) );
  AOI21_X1 U13858 ( .B1(n11407), .B2(n11406), .A(n11405), .ZN(n14821) );
  INV_X1 U13859 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11413) );
  OR2_X1 U13860 ( .A1(n11412), .A2(n11413), .ZN(n11409) );
  NAND2_X1 U13861 ( .A1(n11412), .A2(n11413), .ZN(n11408) );
  AND2_X1 U13862 ( .A1(n11409), .A2(n11408), .ZN(n14792) );
  AOI21_X1 U13863 ( .B1(n10389), .B2(n11411), .A(n11410), .ZN(n14793) );
  NAND2_X1 U13864 ( .A1(n14792), .A2(n14793), .ZN(n14791) );
  OAI21_X1 U13865 ( .B1(n11413), .B2(n11412), .A(n14791), .ZN(n11414) );
  NAND2_X1 U13866 ( .A1(n14801), .A2(n11414), .ZN(n11416) );
  XNOR2_X1 U13867 ( .A(n11415), .B(n11414), .ZN(n14800) );
  NAND2_X1 U13868 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n14800), .ZN(n14799) );
  NAND2_X1 U13869 ( .A1(n11416), .A2(n14799), .ZN(n11417) );
  XOR2_X1 U13870 ( .A(n14809), .B(n11417), .Z(n14810) );
  AOI22_X1 U13871 ( .A1(n14810), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n14809), 
        .B2(n11417), .ZN(n11418) );
  INV_X1 U13872 ( .A(n11418), .ZN(n14822) );
  NAND2_X1 U13873 ( .A1(n14821), .A2(n14822), .ZN(n14819) );
  NAND2_X1 U13874 ( .A1(n11419), .A2(n14819), .ZN(n11422) );
  NAND2_X1 U13875 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n11425), .ZN(n12226) );
  INV_X1 U13876 ( .A(n12226), .ZN(n11420) );
  AOI21_X1 U13877 ( .B1(n13263), .B2(n12231), .A(n11420), .ZN(n11421) );
  NAND2_X1 U13878 ( .A1(n11421), .A2(n11422), .ZN(n12225) );
  OAI211_X1 U13879 ( .C1(n11422), .C2(n11421), .A(n14820), .B(n12225), .ZN(
        n11427) );
  INV_X1 U13880 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n11423) );
  NAND2_X1 U13881 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n11956)
         );
  OAI21_X1 U13882 ( .B1(n14845), .B2(n11423), .A(n11956), .ZN(n11424) );
  AOI21_X1 U13883 ( .B1(n11425), .B2(n14841), .A(n11424), .ZN(n11426) );
  OAI211_X1 U13884 ( .C1(n11428), .C2(n14836), .A(n11427), .B(n11426), .ZN(
        P2_U3231) );
  OR2_X1 U13885 ( .A1(n11594), .A2(n13565), .ZN(n11431) );
  NAND2_X1 U13886 ( .A1(n11432), .A2(n11431), .ZN(n11550) );
  XNOR2_X1 U13887 ( .A(n11550), .B(n11549), .ZN(n14730) );
  INV_X1 U13888 ( .A(n14730), .ZN(n11445) );
  OAI22_X1 U13889 ( .A1(n13962), .A2(n11433), .B1(n11759), .B2(n13913), .ZN(
        n11437) );
  INV_X1 U13890 ( .A(n11434), .ZN(n11435) );
  OAI211_X1 U13891 ( .C1(n6827), .C2(n11435), .A(n6829), .B(n14618), .ZN(
        n14725) );
  NAND2_X1 U13892 ( .A1(n13563), .A2(n13983), .ZN(n14724) );
  AOI21_X1 U13893 ( .B1(n14725), .B2(n14724), .A(n14643), .ZN(n11436) );
  AOI211_X1 U13894 ( .C1(n14634), .C2(n11776), .A(n11437), .B(n11436), .ZN(
        n11444) );
  INV_X1 U13895 ( .A(n11549), .ZN(n11440) );
  OAI211_X1 U13896 ( .C1(n11441), .C2(n11440), .A(n14708), .B(n11547), .ZN(
        n11442) );
  OAI21_X1 U13897 ( .B1(n11582), .B2(n13991), .A(n11442), .ZN(n14727) );
  NAND2_X1 U13898 ( .A1(n14727), .A2(n13962), .ZN(n11443) );
  OAI211_X1 U13899 ( .C1(n11445), .C2(n14008), .A(n11444), .B(n11443), .ZN(
        P1_U3283) );
  INV_X1 U13900 ( .A(n11499), .ZN(n11450) );
  NAND2_X1 U13901 ( .A1(n13020), .A2(n12946), .ZN(n11447) );
  NAND2_X1 U13902 ( .A1(n13022), .A2(n12986), .ZN(n11446) );
  NAND2_X1 U13903 ( .A1(n11447), .A2(n11446), .ZN(n11493) );
  NAND2_X1 U13904 ( .A1(n12992), .A2(n11493), .ZN(n11449) );
  OAI211_X1 U13905 ( .C1(n12990), .C2(n11450), .A(n11449), .B(n11448), .ZN(
        n11455) );
  INV_X1 U13906 ( .A(n11451), .ZN(n12203) );
  AOI211_X1 U13907 ( .C1(n11453), .C2(n11452), .A(n12971), .B(n12203), .ZN(
        n11454) );
  AOI211_X1 U13908 ( .C1(n11500), .C2(n12976), .A(n11455), .B(n11454), .ZN(
        n11456) );
  INV_X1 U13909 ( .A(n11456), .ZN(P2_U3189) );
  INV_X1 U13910 ( .A(n11457), .ZN(n11460) );
  INV_X1 U13911 ( .A(n11458), .ZN(n11459) );
  NAND2_X1 U13912 ( .A1(n11460), .A2(n11459), .ZN(n11461) );
  NAND2_X1 U13913 ( .A1(n11469), .A2(n6435), .ZN(n11465) );
  OR2_X1 U13914 ( .A1(n12162), .A2(n11467), .ZN(n11464) );
  NAND2_X1 U13915 ( .A1(n11465), .A2(n11464), .ZN(n11466) );
  XNOR2_X1 U13916 ( .A(n11466), .B(n12122), .ZN(n11470) );
  NOR2_X1 U13917 ( .A1(n12159), .A2(n11467), .ZN(n11468) );
  AOI21_X1 U13918 ( .B1(n11469), .B2(n10625), .A(n11468), .ZN(n11471) );
  NAND2_X1 U13919 ( .A1(n11470), .A2(n11471), .ZN(n11584) );
  INV_X1 U13920 ( .A(n11470), .ZN(n11473) );
  INV_X1 U13921 ( .A(n11471), .ZN(n11472) );
  NAND2_X1 U13922 ( .A1(n11473), .A2(n11472), .ZN(n11474) );
  NAND2_X1 U13923 ( .A1(n11584), .A2(n11474), .ZN(n11479) );
  INV_X1 U13924 ( .A(n11475), .ZN(n11477) );
  INV_X1 U13925 ( .A(n11479), .ZN(n11476) );
  INV_X1 U13926 ( .A(n11585), .ZN(n11478) );
  AOI21_X1 U13927 ( .B1(n11480), .B2(n11479), .A(n11478), .ZN(n11488) );
  NOR2_X1 U13928 ( .A1(n11481), .A2(n14726), .ZN(n14710) );
  NAND2_X1 U13929 ( .A1(n13475), .A2(n11482), .ZN(n11483) );
  OAI211_X1 U13930 ( .C1(n13553), .C2(n11485), .A(n11484), .B(n11483), .ZN(
        n11486) );
  AOI21_X1 U13931 ( .B1(n13529), .B2(n14710), .A(n11486), .ZN(n11487) );
  OAI21_X1 U13932 ( .B1(n11488), .B2(n13557), .A(n11487), .ZN(P1_U3221) );
  XNOR2_X1 U13933 ( .A(n11490), .B(n11489), .ZN(n14893) );
  INV_X1 U13934 ( .A(n9954), .ZN(n11622) );
  NAND2_X1 U13935 ( .A1(n14893), .A2(n11622), .ZN(n11496) );
  XNOR2_X1 U13936 ( .A(n11492), .B(n11491), .ZN(n11494) );
  AOI21_X1 U13937 ( .B1(n11494), .B2(n14475), .A(n11493), .ZN(n11495) );
  OAI21_X1 U13938 ( .B1(n14890), .B2(n11497), .A(n13083), .ZN(n11498) );
  OR2_X1 U13939 ( .A1(n11498), .A2(n11625), .ZN(n14889) );
  AOI22_X1 U13940 ( .A1(n14478), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n11499), 
        .B2(n14849), .ZN(n11502) );
  NAND2_X1 U13941 ( .A1(n11500), .A2(n14479), .ZN(n11501) );
  OAI211_X1 U13942 ( .C1(n14889), .C2(n13221), .A(n11502), .B(n11501), .ZN(
        n11503) );
  AOI21_X1 U13943 ( .B1(n14893), .B2(n11630), .A(n11503), .ZN(n11504) );
  OAI21_X1 U13944 ( .B1(n14895), .B2(n14478), .A(n11504), .ZN(P2_U3255) );
  OAI21_X1 U13945 ( .B1(n11507), .B2(n11506), .A(n11505), .ZN(n11508) );
  INV_X1 U13946 ( .A(n11508), .ZN(n14702) );
  XNOR2_X1 U13947 ( .A(n11510), .B(n11509), .ZN(n14707) );
  INV_X1 U13948 ( .A(n11511), .ZN(n11512) );
  OAI211_X1 U13949 ( .C1(n14701), .C2(n14620), .A(n11512), .B(n14618), .ZN(
        n14700) );
  MUX2_X1 U13950 ( .A(n14699), .B(n11513), .S(n14647), .Z(n11514) );
  OAI21_X1 U13951 ( .B1(n13913), .B2(n11515), .A(n11514), .ZN(n11516) );
  AOI21_X1 U13952 ( .B1(n14634), .B2(n11517), .A(n11516), .ZN(n11518) );
  OAI21_X1 U13953 ( .B1(n14643), .B2(n14700), .A(n11518), .ZN(n11519) );
  AOI21_X1 U13954 ( .B1(n13869), .B2(n14707), .A(n11519), .ZN(n11520) );
  OAI21_X1 U13955 ( .B1(n14702), .B2(n14008), .A(n11520), .ZN(P1_U3286) );
  AOI22_X1 U13956 ( .A1(n12424), .A2(n11521), .B1(n12418), .B2(n12449), .ZN(
        n11522) );
  NAND2_X1 U13957 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n14946) );
  OAI211_X1 U13958 ( .C1(n11569), .C2(n12421), .A(n11522), .B(n14946), .ZN(
        n11528) );
  INV_X1 U13959 ( .A(n11523), .ZN(n11524) );
  AOI211_X1 U13960 ( .C1(n11526), .C2(n11525), .A(n12439), .B(n11524), .ZN(
        n11527) );
  AOI211_X1 U13961 ( .C1(n11529), .C2(n12437), .A(n11528), .B(n11527), .ZN(
        n11530) );
  INV_X1 U13962 ( .A(n11530), .ZN(P3_U3179) );
  OAI222_X1 U13963 ( .A1(n13438), .A2(n11534), .B1(n11532), .B2(P2_U3088), 
        .C1(n11531), .C2(n13440), .ZN(P2_U3307) );
  OAI222_X1 U13964 ( .A1(n9720), .A2(P1_U3086), .B1(n14281), .B2(n11534), .C1(
        n11533), .C2(n14278), .ZN(P1_U3335) );
  INV_X1 U13965 ( .A(n11535), .ZN(n14892) );
  INV_X1 U13966 ( .A(n11536), .ZN(n11539) );
  AOI211_X1 U13967 ( .C1(n14892), .C2(n11539), .A(n11538), .B(n11537), .ZN(
        n11545) );
  AOI22_X1 U13968 ( .A1(n11543), .A2(n13351), .B1(n14900), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n11540) );
  OAI21_X1 U13969 ( .B1(n11545), .B2(n14900), .A(n11540), .ZN(P2_U3508) );
  INV_X1 U13970 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11541) );
  NOR2_X1 U13971 ( .A1(n14898), .A2(n11541), .ZN(n11542) );
  AOI21_X1 U13972 ( .B1(n11543), .B2(n13407), .A(n11542), .ZN(n11544) );
  OAI21_X1 U13973 ( .B1(n11545), .B2(n14896), .A(n11544), .ZN(P2_U3457) );
  OR2_X1 U13974 ( .A1(n11776), .A2(n11763), .ZN(n11546) );
  NAND2_X1 U13975 ( .A1(n11547), .A2(n11546), .ZN(n11681) );
  INV_X1 U13976 ( .A(n11676), .ZN(n11680) );
  XNOR2_X1 U13977 ( .A(n11681), .B(n11680), .ZN(n11548) );
  OAI222_X1 U13978 ( .A1(n13993), .A2(n11882), .B1(n11548), .B2(n14077), .C1(
        n13991), .C2(n11763), .ZN(n14542) );
  INV_X1 U13979 ( .A(n14542), .ZN(n11559) );
  NAND2_X1 U13980 ( .A1(n11550), .A2(n11549), .ZN(n11552) );
  OR2_X1 U13981 ( .A1(n11776), .A2(n13564), .ZN(n11551) );
  NAND2_X1 U13982 ( .A1(n11552), .A2(n11551), .ZN(n11677) );
  XNOR2_X1 U13983 ( .A(n11677), .B(n11676), .ZN(n14544) );
  INV_X1 U13984 ( .A(n11797), .ZN(n14541) );
  OAI211_X1 U13985 ( .C1(n14541), .C2(n11553), .A(n14618), .B(n11688), .ZN(
        n14540) );
  OAI22_X1 U13986 ( .A1(n13962), .A2(n11554), .B1(n11795), .B2(n13913), .ZN(
        n11555) );
  AOI21_X1 U13987 ( .B1(n11797), .B2(n14634), .A(n11555), .ZN(n11556) );
  OAI21_X1 U13988 ( .B1(n14540), .B2(n14643), .A(n11556), .ZN(n11557) );
  AOI21_X1 U13989 ( .B1(n14544), .B2(n13967), .A(n11557), .ZN(n11558) );
  OAI21_X1 U13990 ( .B1(n11559), .B2(n14647), .A(n11558), .ZN(P1_U3282) );
  INV_X1 U13991 ( .A(n11560), .ZN(n11574) );
  INV_X1 U13992 ( .A(n11561), .ZN(n11563) );
  NAND2_X1 U13993 ( .A1(n11563), .A2(n11562), .ZN(n11564) );
  NAND2_X1 U13994 ( .A1(n11565), .A2(n11564), .ZN(n11568) );
  XNOR2_X1 U13995 ( .A(n12284), .B(n15131), .ZN(n11734) );
  XNOR2_X1 U13996 ( .A(n11734), .B(n11566), .ZN(n11567) );
  NAND2_X1 U13997 ( .A1(n11568), .A2(n11567), .ZN(n11736) );
  OAI211_X1 U13998 ( .C1(n11568), .C2(n11567), .A(n11736), .B(n12381), .ZN(
        n11573) );
  OAI22_X1 U13999 ( .A1(n12434), .A2(n15131), .B1(n11569), .B2(n12433), .ZN(
        n11570) );
  AOI211_X1 U14000 ( .C1(n12431), .C2(n11807), .A(n11571), .B(n11570), .ZN(
        n11572) );
  OAI211_X1 U14001 ( .C1(n11574), .C2(n11810), .A(n11573), .B(n11572), .ZN(
        P3_U3161) );
  NAND2_X1 U14002 ( .A1(n11575), .A2(n12872), .ZN(n11577) );
  OAI211_X1 U14003 ( .C1(n11578), .C2(n12040), .A(n11577), .B(n11576), .ZN(
        P3_U3272) );
  NAND2_X1 U14004 ( .A1(n11594), .A2(n6435), .ZN(n11580) );
  OR2_X1 U14005 ( .A1(n12071), .A2(n11582), .ZN(n11579) );
  NAND2_X1 U14006 ( .A1(n11580), .A2(n11579), .ZN(n11581) );
  XNOR2_X1 U14007 ( .A(n11581), .B(n12160), .ZN(n11765) );
  NOR2_X1 U14008 ( .A1(n12159), .A2(n11582), .ZN(n11583) );
  AOI21_X1 U14009 ( .B1(n11594), .B2(n10625), .A(n11583), .ZN(n11766) );
  XNOR2_X1 U14010 ( .A(n11765), .B(n11766), .ZN(n11587) );
  OAI21_X1 U14011 ( .B1(n11587), .B2(n11586), .A(n11769), .ZN(n11588) );
  NAND2_X1 U14012 ( .A1(n11588), .A2(n13537), .ZN(n11596) );
  NAND2_X1 U14013 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n13654) );
  INV_X1 U14014 ( .A(n13654), .ZN(n11589) );
  AOI21_X1 U14015 ( .B1(n13511), .B2(n13564), .A(n11589), .ZN(n11591) );
  NAND2_X1 U14016 ( .A1(n13551), .A2(n13566), .ZN(n11590) );
  OAI211_X1 U14017 ( .C1(n13553), .C2(n11592), .A(n11591), .B(n11590), .ZN(
        n11593) );
  AOI21_X1 U14018 ( .B1(n13555), .B2(n11594), .A(n11593), .ZN(n11595) );
  NAND2_X1 U14019 ( .A1(n11596), .A2(n11595), .ZN(P1_U3231) );
  OAI222_X1 U14020 ( .A1(n13438), .A2(n11649), .B1(n11598), .B2(P2_U3088), 
        .C1(n11597), .C2(n13440), .ZN(P2_U3306) );
  NOR2_X1 U14021 ( .A1(n11607), .A2(n11599), .ZN(n11601) );
  NOR2_X1 U14022 ( .A1(n11601), .A2(n11600), .ZN(n11605) );
  INV_X1 U14023 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11603) );
  NAND2_X1 U14024 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n11610), .ZN(n11703) );
  INV_X1 U14025 ( .A(n11703), .ZN(n11602) );
  AOI21_X1 U14026 ( .B1(n11603), .B2(n11696), .A(n11602), .ZN(n11604) );
  NAND2_X1 U14027 ( .A1(n11604), .A2(n11605), .ZN(n11702) );
  OAI211_X1 U14028 ( .C1(n11605), .C2(n11604), .A(n14602), .B(n11702), .ZN(
        n11615) );
  NAND2_X1 U14029 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13486)
         );
  NOR2_X1 U14030 ( .A1(n11607), .A2(n11606), .ZN(n11609) );
  XNOR2_X1 U14031 ( .A(n11610), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n11695) );
  XNOR2_X1 U14032 ( .A(n11694), .B(n11695), .ZN(n11611) );
  NAND2_X1 U14033 ( .A1(n14597), .A2(n11611), .ZN(n11612) );
  NAND2_X1 U14034 ( .A1(n13486), .A2(n11612), .ZN(n11613) );
  AOI21_X1 U14035 ( .B1(n14578), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n11613), 
        .ZN(n11614) );
  OAI211_X1 U14036 ( .C1(n13677), .C2(n11696), .A(n11615), .B(n11614), .ZN(
        P1_U3259) );
  INV_X1 U14037 ( .A(n11616), .ZN(n11617) );
  AOI21_X1 U14038 ( .B1(n11619), .B2(n11618), .A(n11617), .ZN(n11624) );
  AOI22_X1 U14039 ( .A1(n12986), .A2(n13021), .B1(n13019), .B2(n12946), .ZN(
        n12199) );
  XNOR2_X1 U14040 ( .A(n11621), .B(n11620), .ZN(n11727) );
  NAND2_X1 U14041 ( .A1(n11727), .A2(n11622), .ZN(n11623) );
  OAI211_X1 U14042 ( .C1(n11624), .C2(n13279), .A(n12199), .B(n11623), .ZN(
        n11725) );
  INV_X1 U14043 ( .A(n11725), .ZN(n11632) );
  INV_X1 U14044 ( .A(n11625), .ZN(n11626) );
  AOI211_X1 U14045 ( .C1(n12208), .C2(n11626), .A(n7779), .B(n6560), .ZN(
        n11726) );
  NAND2_X1 U14046 ( .A1(n11726), .A2(n14847), .ZN(n11628) );
  AOI22_X1 U14047 ( .A1(n14478), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n12197), 
        .B2(n14849), .ZN(n11627) );
  OAI211_X1 U14048 ( .C1(n11729), .C2(n14853), .A(n11628), .B(n11627), .ZN(
        n11629) );
  AOI21_X1 U14049 ( .B1(n11727), .B2(n11630), .A(n11629), .ZN(n11631) );
  OAI21_X1 U14050 ( .B1(n11632), .B2(n14478), .A(n11631), .ZN(P2_U3254) );
  XNOR2_X1 U14051 ( .A(n11634), .B(n11633), .ZN(n14510) );
  INV_X1 U14052 ( .A(n14510), .ZN(n11648) );
  NAND2_X1 U14053 ( .A1(n11635), .A2(n14475), .ZN(n11641) );
  AOI21_X1 U14054 ( .B1(n11616), .B2(n11637), .A(n11636), .ZN(n11640) );
  NAND2_X1 U14055 ( .A1(n13018), .A2(n12946), .ZN(n11639) );
  NAND2_X1 U14056 ( .A1(n13020), .A2(n12986), .ZN(n11638) );
  AND2_X1 U14057 ( .A1(n11639), .A2(n11638), .ZN(n11658) );
  OAI21_X1 U14058 ( .B1(n11641), .B2(n11640), .A(n11658), .ZN(n14508) );
  INV_X1 U14059 ( .A(n11643), .ZN(n14507) );
  OAI211_X1 U14060 ( .C1(n6560), .C2(n14507), .A(n13083), .B(n6774), .ZN(
        n14506) );
  AOI22_X1 U14061 ( .A1(n14478), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n11661), 
        .B2(n14849), .ZN(n11645) );
  NAND2_X1 U14062 ( .A1(n11643), .A2(n14479), .ZN(n11644) );
  OAI211_X1 U14063 ( .C1(n14506), .C2(n13221), .A(n11645), .B(n11644), .ZN(
        n11646) );
  AOI21_X1 U14064 ( .B1(n14508), .B2(n14868), .A(n11646), .ZN(n11647) );
  OAI21_X1 U14065 ( .B1(n11648), .B2(n13254), .A(n11647), .ZN(P2_U3253) );
  OAI222_X1 U14066 ( .A1(n11650), .A2(P1_U3086), .B1(n14281), .B2(n11649), 
        .C1(n14126), .C2(n14278), .ZN(P1_U3334) );
  INV_X1 U14067 ( .A(n11668), .ZN(n11662) );
  INV_X1 U14068 ( .A(n11651), .ZN(n11654) );
  AOI21_X1 U14069 ( .B1(n11654), .B2(n11653), .A(n11652), .ZN(n11655) );
  AOI21_X1 U14070 ( .B1(n11662), .B2(n11656), .A(n11655), .ZN(n11665) );
  OAI22_X1 U14071 ( .A1(n12961), .A2(n11658), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11657), .ZN(n11660) );
  NOR2_X1 U14072 ( .A1(n14507), .A2(n12994), .ZN(n11659) );
  AOI211_X1 U14073 ( .C1(n12964), .C2(n11661), .A(n11660), .B(n11659), .ZN(
        n11664) );
  NAND3_X1 U14074 ( .A1(n11662), .A2(n12953), .A3(n13019), .ZN(n11663) );
  OAI211_X1 U14075 ( .C1(n11665), .C2(n12971), .A(n11664), .B(n11663), .ZN(
        P2_U3196) );
  OAI211_X1 U14076 ( .C1(n11669), .C2(n11668), .A(n11667), .B(n12996), .ZN(
        n11675) );
  NAND2_X1 U14077 ( .A1(n13017), .A2(n12946), .ZN(n11671) );
  NAND2_X1 U14078 ( .A1(n13019), .A2(n12986), .ZN(n11670) );
  NAND2_X1 U14079 ( .A1(n11671), .A2(n11670), .ZN(n11746) );
  INV_X1 U14080 ( .A(n11746), .ZN(n11672) );
  OAI22_X1 U14081 ( .A1(n12961), .A2(n11672), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7687), .ZN(n11673) );
  AOI21_X1 U14082 ( .B1(n11750), .B2(n12964), .A(n11673), .ZN(n11674) );
  OAI211_X1 U14083 ( .C1(n10019), .C2(n12994), .A(n11675), .B(n11674), .ZN(
        P2_U3206) );
  NAND2_X1 U14084 ( .A1(n11677), .A2(n11676), .ZN(n11679) );
  OR2_X1 U14085 ( .A1(n11797), .A2(n13563), .ZN(n11678) );
  NAND2_X1 U14086 ( .A1(n11679), .A2(n11678), .ZN(n11715) );
  INV_X1 U14087 ( .A(n11714), .ZN(n11709) );
  XNOR2_X1 U14088 ( .A(n11715), .B(n11709), .ZN(n14411) );
  NAND2_X1 U14089 ( .A1(n11681), .A2(n11680), .ZN(n11683) );
  OR2_X1 U14090 ( .A1(n11797), .A2(n11781), .ZN(n11682) );
  NAND2_X1 U14091 ( .A1(n11683), .A2(n11682), .ZN(n11710) );
  XNOR2_X1 U14092 ( .A(n11710), .B(n11714), .ZN(n11685) );
  OAI22_X1 U14093 ( .A1(n11928), .A2(n13993), .B1(n11781), .B2(n13991), .ZN(
        n11684) );
  AOI21_X1 U14094 ( .B1(n11685), .B2(n14708), .A(n11684), .ZN(n11686) );
  OAI21_X1 U14095 ( .B1(n14411), .B2(n14703), .A(n11686), .ZN(n14414) );
  NAND2_X1 U14096 ( .A1(n14414), .A2(n13962), .ZN(n11693) );
  OAI22_X1 U14097 ( .A1(n13962), .A2(n11687), .B1(n11887), .B2(n13913), .ZN(
        n11691) );
  INV_X1 U14098 ( .A(n11688), .ZN(n11689) );
  INV_X1 U14099 ( .A(n11884), .ZN(n14413) );
  OAI211_X1 U14100 ( .C1(n11689), .C2(n14413), .A(n14618), .B(n11717), .ZN(
        n14412) );
  NOR2_X1 U14101 ( .A1(n14412), .A2(n14643), .ZN(n11690) );
  AOI211_X1 U14102 ( .C1(n14634), .C2(n11884), .A(n11691), .B(n11690), .ZN(
        n11692) );
  OAI211_X1 U14103 ( .C1(n14411), .C2(n14641), .A(n11693), .B(n11692), .ZN(
        P1_U3281) );
  NAND2_X1 U14104 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13494)
         );
  XNOR2_X1 U14105 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n13668), .ZN(n11699) );
  INV_X1 U14106 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n11697) );
  OAI211_X1 U14107 ( .C1(n11699), .C2(n11698), .A(n14597), .B(n13667), .ZN(
        n11700) );
  NAND2_X1 U14108 ( .A1(n13494), .A2(n11700), .ZN(n11701) );
  AOI21_X1 U14109 ( .B1(n14578), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n11701), 
        .ZN(n11708) );
  NAND2_X1 U14110 ( .A1(n11703), .A2(n11702), .ZN(n11706) );
  AOI22_X1 U14111 ( .A1(n11704), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n13959), 
        .B2(n13668), .ZN(n11705) );
  NAND2_X1 U14112 ( .A1(n11705), .A2(n11706), .ZN(n13665) );
  OAI211_X1 U14113 ( .C1(n11706), .C2(n11705), .A(n14602), .B(n13665), .ZN(
        n11707) );
  OAI211_X1 U14114 ( .C1(n13677), .C2(n13668), .A(n11708), .B(n11707), .ZN(
        P1_U3260) );
  NAND2_X1 U14115 ( .A1(n11710), .A2(n11709), .ZN(n11712) );
  OR2_X1 U14116 ( .A1(n11884), .A2(n11882), .ZN(n11711) );
  NAND2_X1 U14117 ( .A1(n11712), .A2(n11711), .ZN(n11833) );
  INV_X1 U14118 ( .A(n11846), .ZN(n11832) );
  XNOR2_X1 U14119 ( .A(n11833), .B(n11832), .ZN(n11713) );
  OAI222_X1 U14120 ( .A1(n13993), .A2(n13992), .B1(n11713), .B2(n14077), .C1(
        n13991), .C2(n11882), .ZN(n14537) );
  INV_X1 U14121 ( .A(n14537), .ZN(n11724) );
  OR2_X1 U14122 ( .A1(n11884), .A2(n13562), .ZN(n11716) );
  XNOR2_X1 U14123 ( .A(n11847), .B(n11846), .ZN(n14539) );
  INV_X1 U14124 ( .A(n11934), .ZN(n14536) );
  INV_X1 U14125 ( .A(n11717), .ZN(n11718) );
  INV_X1 U14126 ( .A(n11842), .ZN(n11840) );
  OAI211_X1 U14127 ( .C1(n14536), .C2(n11718), .A(n14618), .B(n11840), .ZN(
        n14535) );
  OAI22_X1 U14128 ( .A1(n13962), .A2(n11719), .B1(n11932), .B2(n13913), .ZN(
        n11720) );
  AOI21_X1 U14129 ( .B1(n11934), .B2(n14634), .A(n11720), .ZN(n11721) );
  OAI21_X1 U14130 ( .B1(n14535), .B2(n14643), .A(n11721), .ZN(n11722) );
  AOI21_X1 U14131 ( .B1(n14539), .B2(n13967), .A(n11722), .ZN(n11723) );
  OAI21_X1 U14132 ( .B1(n11724), .B2(n14647), .A(n11723), .ZN(P1_U3280) );
  AOI211_X1 U14133 ( .C1(n14892), .C2(n11727), .A(n11726), .B(n11725), .ZN(
        n11733) );
  INV_X1 U14134 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n11728) );
  OAI22_X1 U14135 ( .A1(n11729), .A2(n13420), .B1(n14898), .B2(n11728), .ZN(
        n11730) );
  INV_X1 U14136 ( .A(n11730), .ZN(n11731) );
  OAI21_X1 U14137 ( .B1(n11733), .B2(n14896), .A(n11731), .ZN(P2_U3463) );
  AOI22_X1 U14138 ( .A1(n12208), .A2(n13351), .B1(n14900), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n11732) );
  OAI21_X1 U14139 ( .B1(n11733), .B2(n14900), .A(n11732), .ZN(P2_U3510) );
  XNOR2_X1 U14140 ( .A(n12284), .B(n15046), .ZN(n11800) );
  XNOR2_X1 U14141 ( .A(n11800), .B(n11807), .ZN(n11739) );
  NAND2_X1 U14142 ( .A1(n11734), .A2(n15040), .ZN(n11735) );
  INV_X1 U14143 ( .A(n11803), .ZN(n11737) );
  AOI21_X1 U14144 ( .B1(n11739), .B2(n11738), .A(n11737), .ZN(n11744) );
  NOR2_X1 U14145 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11740), .ZN(n14951) );
  OAI22_X1 U14146 ( .A1(n12434), .A2(n15046), .B1(n11946), .B2(n12421), .ZN(
        n11741) );
  AOI211_X1 U14147 ( .C1(n12418), .C2(n15040), .A(n14951), .B(n11741), .ZN(
        n11743) );
  NAND2_X1 U14148 ( .A1(n12437), .A2(n15047), .ZN(n11742) );
  OAI211_X1 U14149 ( .C1(n11744), .C2(n12439), .A(n11743), .B(n11742), .ZN(
        P3_U3171) );
  XOR2_X1 U14150 ( .A(n11745), .B(n11748), .Z(n11747) );
  AOI21_X1 U14151 ( .B1(n11747), .B2(n14475), .A(n11746), .ZN(n14502) );
  XOR2_X1 U14152 ( .A(n11749), .B(n11748), .Z(n14504) );
  NAND2_X1 U14153 ( .A1(n14504), .A2(n14856), .ZN(n11755) );
  OAI211_X1 U14154 ( .C1(n10019), .C2(n11642), .A(n13083), .B(n14483), .ZN(
        n14501) );
  INV_X1 U14155 ( .A(n14501), .ZN(n11753) );
  AOI22_X1 U14156 ( .A1(n14478), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n11750), 
        .B2(n14849), .ZN(n11751) );
  OAI21_X1 U14157 ( .B1(n10019), .B2(n14853), .A(n11751), .ZN(n11752) );
  AOI21_X1 U14158 ( .B1(n11753), .B2(n14847), .A(n11752), .ZN(n11754) );
  OAI211_X1 U14159 ( .C1(n14478), .C2(n14502), .A(n11755), .B(n11754), .ZN(
        P2_U3252) );
  AOI21_X1 U14160 ( .B1(n13511), .B2(n13563), .A(n11756), .ZN(n11758) );
  NAND2_X1 U14161 ( .A1(n13551), .A2(n13565), .ZN(n11757) );
  OAI211_X1 U14162 ( .C1(n13553), .C2(n11759), .A(n11758), .B(n11757), .ZN(
        n11775) );
  NAND2_X1 U14163 ( .A1(n11776), .A2(n6435), .ZN(n11761) );
  OR2_X1 U14164 ( .A1(n12071), .A2(n11763), .ZN(n11760) );
  NAND2_X1 U14165 ( .A1(n11761), .A2(n11760), .ZN(n11762) );
  XNOR2_X1 U14166 ( .A(n11762), .B(n12160), .ZN(n11785) );
  NOR2_X1 U14167 ( .A1(n12159), .A2(n11763), .ZN(n11764) );
  AOI21_X1 U14168 ( .B1(n11776), .B2(n10625), .A(n11764), .ZN(n11783) );
  XNOR2_X1 U14169 ( .A(n11785), .B(n11783), .ZN(n11770) );
  INV_X1 U14170 ( .A(n11765), .ZN(n11767) );
  NAND2_X1 U14171 ( .A1(n11767), .A2(n11766), .ZN(n11771) );
  AND2_X1 U14172 ( .A1(n11770), .A2(n11771), .ZN(n11768) );
  INV_X1 U14173 ( .A(n11787), .ZN(n11773) );
  AOI21_X1 U14174 ( .B1(n11769), .B2(n11771), .A(n11770), .ZN(n11772) );
  NOR3_X1 U14175 ( .A1(n11773), .A2(n11772), .A3(n13557), .ZN(n11774) );
  AOI211_X1 U14176 ( .C1(n13555), .C2(n11776), .A(n11775), .B(n11774), .ZN(
        n11777) );
  INV_X1 U14177 ( .A(n11777), .ZN(P1_U3217) );
  NAND2_X1 U14178 ( .A1(n11797), .A2(n6435), .ZN(n11779) );
  OR2_X1 U14179 ( .A1(n12162), .A2(n11781), .ZN(n11778) );
  NAND2_X1 U14180 ( .A1(n11779), .A2(n11778), .ZN(n11780) );
  XNOR2_X1 U14181 ( .A(n11780), .B(n12122), .ZN(n11876) );
  NOR2_X1 U14182 ( .A1(n12159), .A2(n11781), .ZN(n11782) );
  AOI21_X1 U14183 ( .B1(n11797), .B2(n10625), .A(n11782), .ZN(n11875) );
  XNOR2_X1 U14184 ( .A(n11876), .B(n11875), .ZN(n11791) );
  INV_X1 U14185 ( .A(n11783), .ZN(n11784) );
  NAND2_X1 U14186 ( .A1(n11785), .A2(n11784), .ZN(n11786) );
  INV_X1 U14187 ( .A(n11878), .ZN(n11789) );
  AOI21_X1 U14188 ( .B1(n11791), .B2(n11790), .A(n11789), .ZN(n11799) );
  NOR2_X1 U14189 ( .A1(n13549), .A2(n11882), .ZN(n11792) );
  AOI211_X1 U14190 ( .C1(n13551), .C2(n13564), .A(n11793), .B(n11792), .ZN(
        n11794) );
  OAI21_X1 U14191 ( .B1(n13553), .B2(n11795), .A(n11794), .ZN(n11796) );
  AOI21_X1 U14192 ( .B1(n13555), .B2(n11797), .A(n11796), .ZN(n11798) );
  OAI21_X1 U14193 ( .B1(n11799), .B2(n13557), .A(n11798), .ZN(P1_U3236) );
  INV_X1 U14194 ( .A(n15034), .ZN(n11811) );
  INV_X1 U14195 ( .A(n11800), .ZN(n11801) );
  INV_X1 U14196 ( .A(n11807), .ZN(n15028) );
  NAND2_X1 U14197 ( .A1(n11801), .A2(n15028), .ZN(n11802) );
  XNOR2_X1 U14198 ( .A(n12284), .B(n15033), .ZN(n11937) );
  XNOR2_X1 U14199 ( .A(n11937), .B(n11946), .ZN(n11804) );
  OAI211_X1 U14200 ( .C1(n6569), .C2(n11804), .A(n11939), .B(n12381), .ZN(
        n11809) );
  NAND2_X1 U14201 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_U3151), .ZN(n14972)
         );
  OAI21_X1 U14202 ( .B1(n12421), .B2(n6892), .A(n14972), .ZN(n11806) );
  NOR2_X1 U14203 ( .A1(n12434), .A2(n15033), .ZN(n11805) );
  AOI211_X1 U14204 ( .C1(n12418), .C2(n11807), .A(n11806), .B(n11805), .ZN(
        n11808) );
  OAI211_X1 U14205 ( .C1(n11811), .C2(n11810), .A(n11809), .B(n11808), .ZN(
        P3_U3157) );
  INV_X1 U14206 ( .A(n11812), .ZN(n11813) );
  OAI222_X1 U14207 ( .A1(n9849), .A2(P3_U3151), .B1(n12040), .B2(n14087), .C1(
        n12880), .C2(n11813), .ZN(P3_U3271) );
  OAI222_X1 U14208 ( .A1(n13438), .A2(n11816), .B1(n11815), .B2(P2_U3088), 
        .C1(n11814), .C2(n13440), .ZN(P2_U3305) );
  XNOR2_X1 U14209 ( .A(n11817), .B(n11818), .ZN(n14463) );
  INV_X1 U14210 ( .A(n14463), .ZN(n11831) );
  OR2_X1 U14211 ( .A1(n15083), .A2(n15069), .ZN(n11819) );
  NAND2_X1 U14212 ( .A1(n15094), .A2(n11819), .ZN(n12553) );
  OAI211_X1 U14213 ( .C1(n11820), .C2(n11822), .A(n15074), .B(n11821), .ZN(
        n11824) );
  AOI22_X1 U14214 ( .A1(n15076), .A2(n12447), .B1(n12446), .B2(n15079), .ZN(
        n11823) );
  NAND2_X1 U14215 ( .A1(n11824), .A2(n11823), .ZN(n14461) );
  NAND2_X1 U14216 ( .A1(n14461), .A2(n15094), .ZN(n11830) );
  INV_X1 U14217 ( .A(n11982), .ZN(n11825) );
  NOR2_X1 U14218 ( .A1(n11825), .A2(n15130), .ZN(n14462) );
  INV_X1 U14219 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11827) );
  INV_X1 U14220 ( .A(n11986), .ZN(n11826) );
  OAI22_X1 U14221 ( .A1(n15094), .A2(n11827), .B1(n11826), .B2(n15056), .ZN(
        n11828) );
  AOI21_X1 U14222 ( .B1(n14462), .B2(n15048), .A(n11828), .ZN(n11829) );
  OAI211_X1 U14223 ( .C1(n11831), .C2(n12553), .A(n11830), .B(n11829), .ZN(
        P3_U3221) );
  OR2_X1 U14224 ( .A1(n11934), .A2(n11928), .ZN(n11834) );
  OAI211_X1 U14225 ( .C1(n11836), .C2(n11850), .A(n13734), .B(n14708), .ZN(
        n11838) );
  AOI22_X1 U14226 ( .A1(n13982), .A2(n13983), .B1(n13981), .B2(n13561), .ZN(
        n11837) );
  OAI22_X1 U14227 ( .A1(n13962), .A2(n11839), .B1(n12011), .B2(n13913), .ZN(
        n11845) );
  AOI21_X1 U14228 ( .B1(n14528), .B2(n11840), .A(n14636), .ZN(n11843) );
  NAND2_X1 U14229 ( .A1(n11843), .A2(n13998), .ZN(n14530) );
  NOR2_X1 U14230 ( .A1(n14530), .A2(n14643), .ZN(n11844) );
  AOI211_X1 U14231 ( .C1(n14634), .C2(n14528), .A(n11845), .B(n11844), .ZN(
        n11852) );
  OR2_X1 U14232 ( .A1(n11934), .A2(n13561), .ZN(n11848) );
  NAND2_X1 U14233 ( .A1(n11849), .A2(n11850), .ZN(n14531) );
  NAND3_X1 U14234 ( .A1(n6539), .A2(n14531), .A3(n13967), .ZN(n11851) );
  OAI211_X1 U14235 ( .C1(n14534), .C2(n14647), .A(n11852), .B(n11851), .ZN(
        P1_U3279) );
  AOI22_X1 U14236 ( .A1(n11853), .A2(n12996), .B1(n12953), .B2(n13016), .ZN(
        n11863) );
  INV_X1 U14237 ( .A(n11854), .ZN(n11862) );
  INV_X1 U14238 ( .A(n11898), .ZN(n11858) );
  NAND2_X1 U14239 ( .A1(n13015), .A2(n12946), .ZN(n11856) );
  NAND2_X1 U14240 ( .A1(n13017), .A2(n12986), .ZN(n11855) );
  NAND2_X1 U14241 ( .A1(n11856), .A2(n11855), .ZN(n11895) );
  AOI22_X1 U14242 ( .A1(n12992), .A2(n11895), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11857) );
  OAI21_X1 U14243 ( .B1(n11858), .B2(n12990), .A(n11857), .ZN(n11859) );
  AOI21_X1 U14244 ( .B1(n11860), .B2(n12976), .A(n11859), .ZN(n11861) );
  OAI21_X1 U14245 ( .B1(n11863), .B2(n11862), .A(n11861), .ZN(P2_U3213) );
  XNOR2_X1 U14246 ( .A(n11865), .B(n11864), .ZN(n12815) );
  INV_X1 U14247 ( .A(n12815), .ZN(n11874) );
  OAI211_X1 U14248 ( .C1(n11868), .C2(n11867), .A(n11866), .B(n15074), .ZN(
        n11870) );
  AOI22_X1 U14249 ( .A1(n14452), .A2(n15076), .B1(n15079), .B2(n12445), .ZN(
        n11869) );
  NAND2_X1 U14250 ( .A1(n11870), .A2(n11869), .ZN(n12814) );
  AOI22_X1 U14251 ( .A1(n15071), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n15090), 
        .B2(n12392), .ZN(n11871) );
  OAI21_X1 U14252 ( .B1(n12870), .B2(n12744), .A(n11871), .ZN(n11872) );
  AOI21_X1 U14253 ( .B1(n12814), .B2(n15094), .A(n11872), .ZN(n11873) );
  OAI21_X1 U14254 ( .B1(n12553), .B2(n11874), .A(n11873), .ZN(P3_U3220) );
  NAND2_X1 U14255 ( .A1(n11876), .A2(n11875), .ZN(n11877) );
  AND2_X2 U14256 ( .A1(n11878), .A2(n11877), .ZN(n11886) );
  NAND2_X1 U14257 ( .A1(n11884), .A2(n6435), .ZN(n11880) );
  OR2_X1 U14258 ( .A1(n12162), .A2(n11882), .ZN(n11879) );
  NAND2_X1 U14259 ( .A1(n11880), .A2(n11879), .ZN(n11881) );
  XNOR2_X1 U14260 ( .A(n11881), .B(n12160), .ZN(n11922) );
  NOR2_X1 U14261 ( .A1(n12159), .A2(n11882), .ZN(n11883) );
  AOI21_X1 U14262 ( .B1(n11884), .B2(n10625), .A(n11883), .ZN(n11920) );
  XNOR2_X1 U14263 ( .A(n11922), .B(n11920), .ZN(n11885) );
  OAI211_X1 U14264 ( .C1(n11886), .C2(n11885), .A(n11924), .B(n13537), .ZN(
        n11892) );
  NOR2_X1 U14265 ( .A1(n13553), .A2(n11887), .ZN(n11890) );
  OAI21_X1 U14266 ( .B1(n13549), .B2(n11928), .A(n11888), .ZN(n11889) );
  AOI211_X1 U14267 ( .C1(n13551), .C2(n13563), .A(n11890), .B(n11889), .ZN(
        n11891) );
  OAI211_X1 U14268 ( .C1(n14413), .C2(n13526), .A(n11892), .B(n11891), .ZN(
        P1_U3224) );
  AOI21_X1 U14269 ( .B1(n11894), .B2(n11893), .A(n13279), .ZN(n11897) );
  AOI21_X1 U14270 ( .B1(n11897), .B2(n11896), .A(n11895), .ZN(n14492) );
  OAI211_X1 U14271 ( .C1(n14493), .C2(n14484), .A(n13083), .B(n13284), .ZN(
        n14491) );
  INV_X1 U14272 ( .A(n14491), .ZN(n11901) );
  AOI22_X1 U14273 ( .A1(n14478), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n11898), 
        .B2(n14849), .ZN(n11899) );
  OAI21_X1 U14274 ( .B1(n14493), .B2(n14853), .A(n11899), .ZN(n11900) );
  AOI21_X1 U14275 ( .B1(n11901), .B2(n14847), .A(n11900), .ZN(n11905) );
  XNOR2_X1 U14276 ( .A(n11903), .B(n11902), .ZN(n14495) );
  NAND2_X1 U14277 ( .A1(n14495), .A2(n14856), .ZN(n11904) );
  OAI211_X1 U14278 ( .C1(n14492), .C2(n14478), .A(n11905), .B(n11904), .ZN(
        P2_U3250) );
  INV_X1 U14279 ( .A(n11906), .ZN(n11909) );
  OAI222_X1 U14280 ( .A1(n12880), .A2(n11909), .B1(P3_U3151), .B2(n11908), 
        .C1(n11907), .C2(n12040), .ZN(P3_U3270) );
  OAI211_X1 U14281 ( .C1(n11911), .C2(n11914), .A(n11910), .B(n15074), .ZN(
        n11913) );
  AOI22_X1 U14282 ( .A1(n12724), .A2(n15079), .B1(n15076), .B2(n12446), .ZN(
        n11912) );
  NAND2_X1 U14283 ( .A1(n11913), .A2(n11912), .ZN(n12810) );
  INV_X1 U14284 ( .A(n12810), .ZN(n11919) );
  XNOR2_X1 U14285 ( .A(n11915), .B(n11914), .ZN(n12811) );
  AOI22_X1 U14286 ( .A1(n15071), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15090), 
        .B2(n12298), .ZN(n11916) );
  OAI21_X1 U14287 ( .B1(n12866), .B2(n12744), .A(n11916), .ZN(n11917) );
  AOI21_X1 U14288 ( .B1(n12811), .B2(n14458), .A(n11917), .ZN(n11918) );
  OAI21_X1 U14289 ( .B1(n11919), .B2(n15071), .A(n11918), .ZN(P3_U3219) );
  INV_X1 U14290 ( .A(n11920), .ZN(n11921) );
  NAND2_X1 U14291 ( .A1(n11922), .A2(n11921), .ZN(n11923) );
  NAND2_X1 U14292 ( .A1(n11934), .A2(n6435), .ZN(n11926) );
  OR2_X1 U14293 ( .A1(n12162), .A2(n11928), .ZN(n11925) );
  NAND2_X1 U14294 ( .A1(n11926), .A2(n11925), .ZN(n11927) );
  XNOR2_X1 U14295 ( .A(n11927), .B(n12160), .ZN(n12002) );
  NOR2_X1 U14296 ( .A1(n12159), .A2(n11928), .ZN(n11929) );
  AOI21_X1 U14297 ( .B1(n11934), .B2(n10625), .A(n11929), .ZN(n12000) );
  XNOR2_X1 U14298 ( .A(n12002), .B(n12000), .ZN(n11998) );
  XNOR2_X1 U14299 ( .A(n11999), .B(n11998), .ZN(n11936) );
  NAND2_X1 U14300 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n14591)
         );
  OAI21_X1 U14301 ( .B1(n13549), .B2(n13992), .A(n14591), .ZN(n11930) );
  AOI21_X1 U14302 ( .B1(n13551), .B2(n13562), .A(n11930), .ZN(n11931) );
  OAI21_X1 U14303 ( .B1(n13553), .B2(n11932), .A(n11931), .ZN(n11933) );
  AOI21_X1 U14304 ( .B1(n11934), .B2(n13555), .A(n11933), .ZN(n11935) );
  OAI21_X1 U14305 ( .B1(n11936), .B2(n13557), .A(n11935), .ZN(P1_U3234) );
  NAND2_X1 U14306 ( .A1(n11937), .A2(n15039), .ZN(n11938) );
  XNOR2_X1 U14307 ( .A(n14457), .B(n11386), .ZN(n11941) );
  NAND2_X1 U14308 ( .A1(n11940), .A2(n11941), .ZN(n11976) );
  INV_X1 U14309 ( .A(n11940), .ZN(n11943) );
  INV_X1 U14310 ( .A(n11941), .ZN(n11942) );
  NAND2_X1 U14311 ( .A1(n11943), .A2(n11942), .ZN(n11977) );
  NAND2_X1 U14312 ( .A1(n11976), .A2(n11977), .ZN(n11944) );
  XNOR2_X1 U14313 ( .A(n11944), .B(n6892), .ZN(n11951) );
  NOR2_X1 U14314 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11945), .ZN(n14999) );
  NOR2_X1 U14315 ( .A1(n12433), .A2(n11946), .ZN(n11947) );
  AOI211_X1 U14316 ( .C1(n12431), .C2(n14452), .A(n14999), .B(n11947), .ZN(
        n11948) );
  OAI21_X1 U14317 ( .B1(n12434), .B2(n14457), .A(n11948), .ZN(n11949) );
  AOI21_X1 U14318 ( .B1(n12437), .B2(n14454), .A(n11949), .ZN(n11950) );
  OAI21_X1 U14319 ( .B1(n11951), .B2(n12439), .A(n11950), .ZN(P3_U3176) );
  INV_X1 U14320 ( .A(n11952), .ZN(n11954) );
  OAI222_X1 U14321 ( .A1(P3_U3151), .A2(n11955), .B1(n12880), .B2(n11954), 
        .C1(n11953), .C2(n12040), .ZN(P3_U3269) );
  NOR2_X1 U14322 ( .A1(n12990), .A2(n13262), .ZN(n11958) );
  AOI22_X1 U14323 ( .A1(n13013), .A2(n12946), .B1(n12986), .B2(n13015), .ZN(
        n13260) );
  OAI21_X1 U14324 ( .B1(n12961), .B2(n13260), .A(n11956), .ZN(n11957) );
  AOI211_X1 U14325 ( .C1(n13265), .C2(n12976), .A(n11958), .B(n11957), .ZN(
        n11965) );
  OAI22_X1 U14326 ( .A1(n11962), .A2(n12971), .B1(n11961), .B2(n12978), .ZN(
        n11963) );
  NAND3_X1 U14327 ( .A1(n11959), .A2(n6686), .A3(n11963), .ZN(n11964) );
  OAI211_X1 U14328 ( .C1(n11966), .C2(n12971), .A(n11965), .B(n11964), .ZN(
        P2_U3200) );
  INV_X1 U14329 ( .A(n11959), .ZN(n11967) );
  AOI21_X1 U14330 ( .B1(n11969), .B2(n11968), .A(n11967), .ZN(n11975) );
  INV_X1 U14331 ( .A(n11970), .ZN(n13281) );
  NOR2_X1 U14332 ( .A1(n12990), .A2(n13281), .ZN(n11973) );
  AOI22_X1 U14333 ( .A1(n13014), .A2(n12946), .B1(n12986), .B2(n13016), .ZN(
        n13278) );
  OAI22_X1 U14334 ( .A1(n12961), .A2(n13278), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11971), .ZN(n11972) );
  AOI211_X1 U14335 ( .C1(n13285), .C2(n12976), .A(n11973), .B(n11972), .ZN(
        n11974) );
  OAI21_X1 U14336 ( .B1(n11975), .B2(n12971), .A(n11974), .ZN(P2_U3198) );
  XNOR2_X1 U14337 ( .A(n11982), .B(n12284), .ZN(n12248) );
  XNOR2_X1 U14338 ( .A(n12248), .B(n12247), .ZN(n11980) );
  NAND2_X1 U14339 ( .A1(n11976), .A2(n12447), .ZN(n11978) );
  AOI21_X1 U14340 ( .B1(n11980), .B2(n11979), .A(n7209), .ZN(n11988) );
  NOR2_X1 U14341 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11981), .ZN(n12458) );
  AOI21_X1 U14342 ( .B1(n12431), .B2(n12446), .A(n12458), .ZN(n11984) );
  NAND2_X1 U14343 ( .A1(n11982), .A2(n12424), .ZN(n11983) );
  OAI211_X1 U14344 ( .C1(n6892), .C2(n12433), .A(n11984), .B(n11983), .ZN(
        n11985) );
  AOI21_X1 U14345 ( .B1(n12437), .B2(n11986), .A(n11985), .ZN(n11987) );
  OAI21_X1 U14346 ( .B1(n11988), .B2(n12439), .A(n11987), .ZN(P3_U3164) );
  NAND2_X1 U14347 ( .A1(n14528), .A2(n6435), .ZN(n11990) );
  OR2_X1 U14348 ( .A1(n12071), .A2(n13992), .ZN(n11989) );
  NAND2_X1 U14349 ( .A1(n11990), .A2(n11989), .ZN(n11991) );
  XNOR2_X1 U14350 ( .A(n11991), .B(n12122), .ZN(n11993) );
  NOR2_X1 U14351 ( .A1(n12159), .A2(n13992), .ZN(n11992) );
  AOI21_X1 U14352 ( .B1(n14528), .B2(n10625), .A(n11992), .ZN(n11994) );
  NAND2_X1 U14353 ( .A1(n11993), .A2(n11994), .ZN(n12048) );
  INV_X1 U14354 ( .A(n11993), .ZN(n11996) );
  INV_X1 U14355 ( .A(n11994), .ZN(n11995) );
  NAND2_X1 U14356 ( .A1(n11996), .A2(n11995), .ZN(n11997) );
  NAND2_X1 U14357 ( .A1(n12048), .A2(n11997), .ZN(n12007) );
  INV_X1 U14358 ( .A(n12000), .ZN(n12001) );
  NAND2_X1 U14359 ( .A1(n12002), .A2(n12001), .ZN(n12003) );
  INV_X1 U14360 ( .A(n12007), .ZN(n12004) );
  INV_X1 U14361 ( .A(n12049), .ZN(n12005) );
  AOI21_X1 U14362 ( .B1(n12007), .B2(n12006), .A(n12005), .ZN(n12014) );
  OAI21_X1 U14363 ( .B1(n13549), .B2(n12051), .A(n12008), .ZN(n12009) );
  AOI21_X1 U14364 ( .B1(n13551), .B2(n13561), .A(n12009), .ZN(n12010) );
  OAI21_X1 U14365 ( .B1(n13553), .B2(n12011), .A(n12010), .ZN(n12012) );
  AOI21_X1 U14366 ( .B1(n14528), .B2(n13555), .A(n12012), .ZN(n12013) );
  OAI21_X1 U14367 ( .B1(n12014), .B2(n13557), .A(n12013), .ZN(P1_U3215) );
  INV_X1 U14368 ( .A(n12015), .ZN(n12017) );
  OAI222_X1 U14369 ( .A1(n13438), .A2(n12019), .B1(n12017), .B2(P2_U3088), 
        .C1(n12016), .C2(n13440), .ZN(P2_U3303) );
  OAI222_X1 U14370 ( .A1(n12020), .A2(P1_U3086), .B1(n14281), .B2(n12019), 
        .C1(n12018), .C2(n14278), .ZN(P1_U3331) );
  INV_X1 U14371 ( .A(n12021), .ZN(n13431) );
  OAI222_X1 U14372 ( .A1(P1_U3086), .A2(n9784), .B1(n14281), .B2(n13431), .C1(
        n12022), .C2(n14278), .ZN(P1_U3327) );
  INV_X1 U14373 ( .A(n12023), .ZN(n14274) );
  OAI222_X1 U14374 ( .A1(n13440), .A2(n12025), .B1(n13438), .B2(n14274), .C1(
        P2_U3088), .C2(n12024), .ZN(P2_U3300) );
  INV_X1 U14375 ( .A(n12026), .ZN(n12028) );
  OAI222_X1 U14376 ( .A1(n12029), .A2(P3_U3151), .B1(n12880), .B2(n12028), 
        .C1(n12027), .C2(n12040), .ZN(P3_U3267) );
  INV_X1 U14377 ( .A(n9669), .ZN(n13428) );
  OAI222_X1 U14378 ( .A1(P1_U3086), .A2(n12031), .B1(n14281), .B2(n13428), 
        .C1(n12030), .C2(n14278), .ZN(P1_U3326) );
  OAI222_X1 U14379 ( .A1(n13438), .A2(n14272), .B1(n12033), .B2(P2_U3088), 
        .C1(n12032), .C2(n13440), .ZN(P2_U3297) );
  AOI21_X1 U14380 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n13433), .A(n12034), 
        .ZN(n12035) );
  OAI21_X1 U14381 ( .B1(n12038), .B2(n13438), .A(n12035), .ZN(P2_U3304) );
  AOI21_X1 U14382 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n12036), .A(n9772), 
        .ZN(n12037) );
  OAI21_X1 U14383 ( .B1(n12038), .B2(n14281), .A(n12037), .ZN(P1_U3332) );
  INV_X1 U14384 ( .A(n12039), .ZN(n12043) );
  OAI222_X1 U14385 ( .A1(n12880), .A2(n12043), .B1(n12042), .B2(P3_U3151), 
        .C1(n12041), .C2(n12040), .ZN(P3_U3266) );
  INV_X1 U14386 ( .A(n14058), .ZN(n13860) );
  AND2_X1 U14387 ( .A1(n6594), .A2(n13903), .ZN(n12044) );
  AOI21_X1 U14388 ( .B1(n14221), .B2(n10625), .A(n12044), .ZN(n12075) );
  INV_X1 U14389 ( .A(n12075), .ZN(n12081) );
  NAND2_X1 U14390 ( .A1(n14221), .A2(n6435), .ZN(n12046) );
  NAND2_X1 U14391 ( .A1(n13903), .A2(n10625), .ZN(n12045) );
  NAND2_X1 U14392 ( .A1(n12046), .A2(n12045), .ZN(n12047) );
  XNOR2_X1 U14393 ( .A(n12047), .B(n12122), .ZN(n12076) );
  INV_X1 U14394 ( .A(n12076), .ZN(n12080) );
  AOI22_X1 U14395 ( .A1(n14522), .A2(n6435), .B1(n10625), .B2(n13982), .ZN(
        n12050) );
  XOR2_X1 U14396 ( .A(n12160), .B(n12050), .Z(n12054) );
  INV_X1 U14397 ( .A(n14522), .ZN(n14003) );
  OAI22_X1 U14398 ( .A1(n14003), .A2(n12162), .B1(n12051), .B2(n12159), .ZN(
        n13547) );
  INV_X1 U14399 ( .A(n12052), .ZN(n12053) );
  AOI22_X2 U14400 ( .A1(n13548), .A2(n13547), .B1(n12054), .B2(n12053), .ZN(
        n13482) );
  OAI22_X1 U14401 ( .A1(n13977), .A2(n10900), .B1(n13994), .B2(n12071), .ZN(
        n12055) );
  XNOR2_X1 U14402 ( .A(n12055), .B(n12122), .ZN(n12059) );
  INV_X1 U14403 ( .A(n12059), .ZN(n12061) );
  OR2_X1 U14404 ( .A1(n13977), .A2(n12162), .ZN(n12057) );
  NAND2_X1 U14405 ( .A1(n6594), .A2(n13560), .ZN(n12056) );
  AND2_X1 U14406 ( .A1(n12057), .A2(n12056), .ZN(n12058) );
  INV_X1 U14407 ( .A(n12058), .ZN(n12060) );
  AOI21_X1 U14408 ( .B1(n12061), .B2(n12060), .A(n12062), .ZN(n13483) );
  INV_X1 U14409 ( .A(n12062), .ZN(n13491) );
  NAND2_X1 U14410 ( .A1(n14232), .A2(n6435), .ZN(n12064) );
  NAND2_X1 U14411 ( .A1(n10625), .A2(n13984), .ZN(n12063) );
  NAND2_X1 U14412 ( .A1(n12064), .A2(n12063), .ZN(n12065) );
  XNOR2_X1 U14413 ( .A(n12065), .B(n12122), .ZN(n12068) );
  NOR2_X1 U14414 ( .A1(n12159), .A2(n13739), .ZN(n12066) );
  AOI21_X1 U14415 ( .B1(n14232), .B2(n10625), .A(n12066), .ZN(n12067) );
  NAND2_X1 U14416 ( .A1(n12068), .A2(n12067), .ZN(n12069) );
  OAI21_X1 U14417 ( .B1(n12068), .B2(n12067), .A(n12069), .ZN(n13490) );
  INV_X1 U14418 ( .A(n12069), .ZN(n12070) );
  INV_X1 U14419 ( .A(n13955), .ZN(n13715) );
  AOI22_X1 U14420 ( .A1(n13946), .A2(n10625), .B1(n6594), .B2(n13715), .ZN(
        n12077) );
  NAND2_X1 U14421 ( .A1(n13946), .A2(n6435), .ZN(n12073) );
  OR2_X1 U14422 ( .A1(n13955), .A2(n12071), .ZN(n12072) );
  NAND2_X1 U14423 ( .A1(n12073), .A2(n12072), .ZN(n12074) );
  XNOR2_X1 U14424 ( .A(n12074), .B(n12160), .ZN(n12079) );
  XOR2_X1 U14425 ( .A(n12077), .B(n12079), .Z(n13527) );
  XNOR2_X1 U14426 ( .A(n12076), .B(n12075), .ZN(n13452) );
  INV_X1 U14427 ( .A(n12077), .ZN(n12078) );
  NOR2_X1 U14428 ( .A1(n12079), .A2(n12078), .ZN(n13453) );
  OAI22_X1 U14429 ( .A1(n14082), .A2(n10900), .B1(n13743), .B2(n12162), .ZN(
        n12082) );
  XNOR2_X1 U14430 ( .A(n12082), .B(n12160), .ZN(n12084) );
  OAI22_X1 U14431 ( .A1(n14082), .A2(n12071), .B1(n13743), .B2(n12159), .ZN(
        n12083) );
  XNOR2_X1 U14432 ( .A(n12084), .B(n12083), .ZN(n13509) );
  NAND2_X1 U14433 ( .A1(n14073), .A2(n6435), .ZN(n12086) );
  NAND2_X1 U14434 ( .A1(n13904), .A2(n10625), .ZN(n12085) );
  NAND2_X1 U14435 ( .A1(n12086), .A2(n12085), .ZN(n12087) );
  XNOR2_X1 U14436 ( .A(n12087), .B(n12122), .ZN(n12090) );
  AND2_X1 U14437 ( .A1(n13904), .A2(n6594), .ZN(n12088) );
  AOI21_X1 U14438 ( .B1(n14073), .B2(n10625), .A(n12088), .ZN(n12089) );
  NAND2_X1 U14439 ( .A1(n12090), .A2(n12089), .ZN(n12091) );
  OAI21_X1 U14440 ( .B1(n12090), .B2(n12089), .A(n12091), .ZN(n13462) );
  INV_X1 U14441 ( .A(n12091), .ZN(n13519) );
  NAND2_X1 U14442 ( .A1(n13875), .A2(n6435), .ZN(n12093) );
  NAND2_X1 U14443 ( .A1(n13745), .A2(n10625), .ZN(n12092) );
  NAND2_X1 U14444 ( .A1(n12093), .A2(n12092), .ZN(n12094) );
  XNOR2_X1 U14445 ( .A(n12094), .B(n12122), .ZN(n12096) );
  AND2_X1 U14446 ( .A1(n13745), .A2(n6594), .ZN(n12095) );
  AOI21_X1 U14447 ( .B1(n13875), .B2(n10625), .A(n12095), .ZN(n12097) );
  NAND2_X1 U14448 ( .A1(n12096), .A2(n12097), .ZN(n12111) );
  INV_X1 U14449 ( .A(n12096), .ZN(n12099) );
  INV_X1 U14450 ( .A(n12097), .ZN(n12098) );
  NAND2_X1 U14451 ( .A1(n12099), .A2(n12098), .ZN(n12100) );
  AND2_X1 U14452 ( .A1(n12111), .A2(n12100), .ZN(n13518) );
  NAND2_X1 U14453 ( .A1(n14058), .A2(n6435), .ZN(n12102) );
  OR2_X1 U14454 ( .A1(n12071), .A2(n13746), .ZN(n12101) );
  NAND2_X1 U14455 ( .A1(n12102), .A2(n12101), .ZN(n12103) );
  XNOR2_X1 U14456 ( .A(n12103), .B(n12122), .ZN(n12105) );
  NOR2_X1 U14457 ( .A1(n12159), .A2(n13746), .ZN(n12104) );
  AOI21_X1 U14458 ( .B1(n14058), .B2(n10625), .A(n12104), .ZN(n12106) );
  NAND2_X1 U14459 ( .A1(n12105), .A2(n12106), .ZN(n12119) );
  INV_X1 U14460 ( .A(n12105), .ZN(n12108) );
  INV_X1 U14461 ( .A(n12106), .ZN(n12107) );
  NAND2_X1 U14462 ( .A1(n12108), .A2(n12107), .ZN(n12109) );
  NAND2_X1 U14463 ( .A1(n12119), .A2(n12109), .ZN(n12110) );
  AND3_X1 U14464 ( .A1(n13517), .A2(n12111), .A3(n12110), .ZN(n12112) );
  OAI21_X1 U14465 ( .B1(n12130), .B2(n12112), .A(n13537), .ZN(n12118) );
  INV_X1 U14466 ( .A(n13859), .ZN(n12116) );
  AND2_X1 U14467 ( .A1(n13725), .A2(n13983), .ZN(n12113) );
  AOI21_X1 U14468 ( .B1(n13745), .B2(n13981), .A(n12113), .ZN(n14056) );
  INV_X1 U14469 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n12114) );
  OAI22_X1 U14470 ( .A1(n14056), .A2(n13540), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12114), .ZN(n12115) );
  AOI21_X1 U14471 ( .B1(n12116), .B2(n13543), .A(n12115), .ZN(n12117) );
  OAI211_X1 U14472 ( .C1(n13860), .C2(n13526), .A(n12118), .B(n12117), .ZN(
        P1_U3216) );
  INV_X1 U14473 ( .A(n12119), .ZN(n13501) );
  NAND2_X1 U14474 ( .A1(n14051), .A2(n6435), .ZN(n12121) );
  INV_X1 U14475 ( .A(n13725), .ZN(n13747) );
  OR2_X1 U14476 ( .A1(n12162), .A2(n13747), .ZN(n12120) );
  NAND2_X1 U14477 ( .A1(n12121), .A2(n12120), .ZN(n12123) );
  XNOR2_X1 U14478 ( .A(n12123), .B(n12122), .ZN(n12125) );
  NOR2_X1 U14479 ( .A1(n12159), .A2(n13747), .ZN(n12124) );
  AOI21_X1 U14480 ( .B1(n14051), .B2(n10625), .A(n12124), .ZN(n12126) );
  NAND2_X1 U14481 ( .A1(n12125), .A2(n12126), .ZN(n12131) );
  INV_X1 U14482 ( .A(n12125), .ZN(n12128) );
  INV_X1 U14483 ( .A(n12126), .ZN(n12127) );
  NAND2_X1 U14484 ( .A1(n12128), .A2(n12127), .ZN(n12129) );
  AND2_X1 U14485 ( .A1(n12131), .A2(n12129), .ZN(n13500) );
  NAND2_X1 U14486 ( .A1(n14045), .A2(n6435), .ZN(n12133) );
  INV_X1 U14487 ( .A(n13728), .ZN(n13748) );
  OR2_X1 U14488 ( .A1(n12071), .A2(n13748), .ZN(n12132) );
  NAND2_X1 U14489 ( .A1(n12133), .A2(n12132), .ZN(n12134) );
  XNOR2_X1 U14490 ( .A(n12134), .B(n12160), .ZN(n12138) );
  NAND2_X1 U14491 ( .A1(n14045), .A2(n10625), .ZN(n12136) );
  NAND2_X1 U14492 ( .A1(n6594), .A2(n13728), .ZN(n12135) );
  NAND2_X1 U14493 ( .A1(n12136), .A2(n12135), .ZN(n12137) );
  NOR2_X1 U14494 ( .A1(n12138), .A2(n12137), .ZN(n12139) );
  AOI21_X1 U14495 ( .B1(n12138), .B2(n12137), .A(n12139), .ZN(n13472) );
  NAND2_X1 U14496 ( .A1(n13470), .A2(n13472), .ZN(n13471) );
  INV_X1 U14497 ( .A(n12139), .ZN(n12140) );
  NAND2_X1 U14498 ( .A1(n13817), .A2(n6435), .ZN(n12143) );
  OR2_X1 U14499 ( .A1(n12071), .A2(n12141), .ZN(n12142) );
  NAND2_X1 U14500 ( .A1(n12143), .A2(n12142), .ZN(n12144) );
  XNOR2_X1 U14501 ( .A(n12144), .B(n12160), .ZN(n12148) );
  NAND2_X1 U14502 ( .A1(n13817), .A2(n10625), .ZN(n12146) );
  NAND2_X1 U14503 ( .A1(n6594), .A2(n13749), .ZN(n12145) );
  NAND2_X1 U14504 ( .A1(n12146), .A2(n12145), .ZN(n12147) );
  NOR2_X1 U14505 ( .A1(n12148), .A2(n12147), .ZN(n12149) );
  AOI21_X1 U14506 ( .B1(n12148), .B2(n12147), .A(n12149), .ZN(n13536) );
  INV_X1 U14507 ( .A(n12149), .ZN(n12150) );
  INV_X1 U14508 ( .A(n13774), .ZN(n13751) );
  NOR2_X1 U14509 ( .A1(n12162), .A2(n13751), .ZN(n12151) );
  AOI21_X1 U14510 ( .B1(n14034), .B2(n6435), .A(n12151), .ZN(n12153) );
  XNOR2_X1 U14511 ( .A(n12153), .B(n12160), .ZN(n12156) );
  NOR2_X1 U14512 ( .A1(n12159), .A2(n13751), .ZN(n12154) );
  AOI21_X1 U14513 ( .B1(n14034), .B2(n10625), .A(n12154), .ZN(n12155) );
  NAND2_X1 U14514 ( .A1(n12156), .A2(n12155), .ZN(n12158) );
  OAI21_X1 U14515 ( .B1(n12156), .B2(n12155), .A(n12158), .ZN(n12157) );
  INV_X1 U14516 ( .A(n12157), .ZN(n13444) );
  INV_X1 U14517 ( .A(n14028), .ZN(n13783) );
  INV_X1 U14518 ( .A(n13765), .ZN(n13752) );
  OAI22_X1 U14519 ( .A1(n13783), .A2(n12162), .B1(n13752), .B2(n12159), .ZN(
        n12161) );
  XNOR2_X1 U14520 ( .A(n12161), .B(n12160), .ZN(n12164) );
  OAI22_X1 U14521 ( .A1(n13783), .A2(n10900), .B1(n13752), .B2(n12071), .ZN(
        n12163) );
  XNOR2_X1 U14522 ( .A(n12164), .B(n12163), .ZN(n12165) );
  AOI22_X1 U14523 ( .A1(n13551), .A2(n13774), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12167) );
  NAND2_X1 U14524 ( .A1(n13511), .A2(n13773), .ZN(n12166) );
  OAI211_X1 U14525 ( .C1(n13553), .C2(n13780), .A(n12167), .B(n12166), .ZN(
        n12168) );
  AOI21_X1 U14526 ( .B1(n14028), .B2(n13555), .A(n12168), .ZN(n12169) );
  OAI21_X1 U14527 ( .B1(n12170), .B2(n13557), .A(n12169), .ZN(P1_U3220) );
  NAND2_X1 U14528 ( .A1(n12976), .A2(n12171), .ZN(n12175) );
  INV_X1 U14529 ( .A(n12172), .ZN(n12173) );
  NAND2_X1 U14530 ( .A1(n12992), .A2(n12173), .ZN(n12174) );
  NAND2_X1 U14531 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n13043) );
  NAND3_X1 U14532 ( .A1(n12175), .A2(n12174), .A3(n13043), .ZN(n12181) );
  AOI22_X1 U14533 ( .A1(n12953), .A2(n13027), .B1(n12996), .B2(n12176), .ZN(
        n12178) );
  NOR3_X1 U14534 ( .A1(n12179), .A2(n12178), .A3(n12177), .ZN(n12180) );
  AOI211_X1 U14535 ( .C1(n12964), .C2(n12182), .A(n12181), .B(n12180), .ZN(
        n12183) );
  OAI21_X1 U14536 ( .B1(n12184), .B2(n12971), .A(n12183), .ZN(P2_U3199) );
  NAND3_X1 U14537 ( .A1(n12185), .A2(n12953), .A3(n13018), .ZN(n12186) );
  OAI21_X1 U14538 ( .B1(n11667), .B2(n12971), .A(n12186), .ZN(n12194) );
  INV_X1 U14539 ( .A(n12187), .ZN(n12193) );
  OAI22_X1 U14540 ( .A1(n12189), .A2(n12967), .B1(n12188), .B2(n12984), .ZN(
        n14474) );
  AOI22_X1 U14541 ( .A1(n12992), .A2(n14474), .B1(P2_REG3_REG_14__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12191) );
  NAND2_X1 U14542 ( .A1(n12964), .A2(n14477), .ZN(n12190) );
  OAI211_X1 U14543 ( .C1(n6771), .C2(n12994), .A(n12191), .B(n12190), .ZN(
        n12192) );
  AOI21_X1 U14544 ( .B1(n12194), .B2(n12193), .A(n12192), .ZN(n12195) );
  OAI21_X1 U14545 ( .B1(n12196), .B2(n12971), .A(n12195), .ZN(P2_U3187) );
  NAND2_X1 U14546 ( .A1(n12964), .A2(n12197), .ZN(n12198) );
  NAND2_X1 U14547 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n13064)
         );
  OAI211_X1 U14548 ( .C1(n12961), .C2(n12199), .A(n12198), .B(n13064), .ZN(
        n12207) );
  NOR3_X1 U14549 ( .A1(n12201), .A2(n12200), .A3(n12978), .ZN(n12202) );
  AOI21_X1 U14550 ( .B1(n12203), .B2(n12996), .A(n12202), .ZN(n12205) );
  NOR2_X1 U14551 ( .A1(n12205), .A2(n12204), .ZN(n12206) );
  AOI211_X1 U14552 ( .C1(n12208), .C2(n12976), .A(n12207), .B(n12206), .ZN(
        n12209) );
  OAI21_X1 U14553 ( .B1(n12210), .B2(n12971), .A(n12209), .ZN(P2_U3208) );
  NAND2_X1 U14554 ( .A1(n12992), .A2(n12211), .ZN(n12213) );
  OAI211_X1 U14555 ( .C1(n12990), .C2(n12214), .A(n12213), .B(n12212), .ZN(
        n12222) );
  NOR3_X1 U14556 ( .A1(n12216), .A2(n12978), .A3(n12215), .ZN(n12217) );
  AOI21_X1 U14557 ( .B1(n12218), .B2(n12996), .A(n12217), .ZN(n12220) );
  NOR2_X1 U14558 ( .A1(n12220), .A2(n12219), .ZN(n12221) );
  AOI211_X1 U14559 ( .C1(n14881), .C2(n12976), .A(n12222), .B(n12221), .ZN(
        n12223) );
  OAI21_X1 U14560 ( .B1(n12224), .B2(n12971), .A(n12223), .ZN(P2_U3193) );
  NAND2_X1 U14561 ( .A1(n12226), .A2(n12225), .ZN(n12227) );
  NOR2_X1 U14562 ( .A1(n14842), .A2(n12227), .ZN(n12228) );
  XNOR2_X1 U14563 ( .A(n14842), .B(n12227), .ZN(n14833) );
  NOR2_X1 U14564 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n14833), .ZN(n14832) );
  NOR2_X1 U14565 ( .A1(n12228), .A2(n14832), .ZN(n12229) );
  XOR2_X1 U14566 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n12229), .Z(n12238) );
  INV_X1 U14567 ( .A(n12238), .ZN(n12236) );
  OAI21_X1 U14568 ( .B1(n12231), .B2(n13367), .A(n12230), .ZN(n12232) );
  NAND2_X1 U14569 ( .A1(n14842), .A2(n12232), .ZN(n12233) );
  XOR2_X1 U14570 ( .A(n14842), .B(n12232), .Z(n14835) );
  NAND2_X1 U14571 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n14835), .ZN(n14834) );
  NAND2_X1 U14572 ( .A1(n12233), .A2(n14834), .ZN(n12234) );
  XOR2_X1 U14573 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n12234), .Z(n12237) );
  NOR2_X1 U14574 ( .A1(n12237), .A2(n14836), .ZN(n12235) );
  AOI211_X1 U14575 ( .C1(n12236), .C2(n14820), .A(n14841), .B(n12235), .ZN(
        n12241) );
  AOI22_X1 U14576 ( .A1(n12238), .A2(n14820), .B1(n14825), .B2(n12237), .ZN(
        n12240) );
  MUX2_X1 U14577 ( .A(n12241), .B(n12240), .S(n12239), .Z(n12242) );
  NAND2_X1 U14578 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n12909)
         );
  OAI211_X1 U14579 ( .C1(n12243), .C2(n14845), .A(n12242), .B(n12909), .ZN(
        P2_U3233) );
  INV_X1 U14580 ( .A(n12244), .ZN(n12245) );
  OAI222_X1 U14581 ( .A1(P3_U3151), .A2(n8408), .B1(n12040), .B2(n12246), .C1(
        n12880), .C2(n12245), .ZN(P3_U3265) );
  XNOR2_X1 U14582 ( .A(n12289), .B(n11386), .ZN(n12320) );
  XNOR2_X1 U14583 ( .A(n12320), .B(n12422), .ZN(n12322) );
  XNOR2_X1 U14584 ( .A(n12870), .B(n11386), .ZN(n12390) );
  INV_X1 U14585 ( .A(n12446), .ZN(n12389) );
  AND2_X1 U14586 ( .A1(n12390), .A2(n12389), .ZN(n12249) );
  XNOR2_X1 U14587 ( .A(n12866), .B(n12284), .ZN(n12250) );
  XNOR2_X1 U14588 ( .A(n12250), .B(n12739), .ZN(n12292) );
  NAND2_X1 U14589 ( .A1(n12250), .A2(n12445), .ZN(n12251) );
  NAND2_X1 U14590 ( .A1(n12252), .A2(n12251), .ZN(n12427) );
  INV_X1 U14591 ( .A(n12427), .ZN(n12257) );
  XNOR2_X1 U14592 ( .A(n12862), .B(n11386), .ZN(n12253) );
  NAND2_X1 U14593 ( .A1(n12253), .A2(n12357), .ZN(n12258) );
  INV_X1 U14594 ( .A(n12253), .ZN(n12254) );
  NAND2_X1 U14595 ( .A1(n12254), .A2(n12724), .ZN(n12255) );
  NAND2_X1 U14596 ( .A1(n12258), .A2(n12255), .ZN(n12430) );
  NAND2_X1 U14597 ( .A1(n12257), .A2(n12256), .ZN(n12428) );
  NAND2_X1 U14598 ( .A1(n12428), .A2(n12258), .ZN(n12351) );
  XNOR2_X1 U14599 ( .A(n12803), .B(n11386), .ZN(n12352) );
  NAND2_X1 U14600 ( .A1(n12352), .A2(n12710), .ZN(n12259) );
  NAND2_X1 U14601 ( .A1(n12351), .A2(n12259), .ZN(n12262) );
  INV_X1 U14602 ( .A(n12352), .ZN(n12260) );
  NAND2_X1 U14603 ( .A1(n12260), .A2(n12738), .ZN(n12261) );
  NAND2_X1 U14604 ( .A1(n12262), .A2(n12261), .ZN(n12361) );
  XNOR2_X1 U14605 ( .A(n12857), .B(n12284), .ZN(n12263) );
  XNOR2_X1 U14606 ( .A(n12263), .B(n12725), .ZN(n12362) );
  NAND2_X1 U14607 ( .A1(n12263), .A2(n12725), .ZN(n12264) );
  XNOR2_X1 U14608 ( .A(n12793), .B(n12284), .ZN(n12408) );
  XNOR2_X1 U14609 ( .A(n12788), .B(n12284), .ZN(n12265) );
  NAND2_X1 U14610 ( .A1(n12265), .A2(n12411), .ZN(n12310) );
  NAND2_X1 U14611 ( .A1(n12312), .A2(n12310), .ZN(n12267) );
  INV_X1 U14612 ( .A(n12265), .ZN(n12266) );
  NAND2_X1 U14613 ( .A1(n12266), .A2(n12691), .ZN(n12311) );
  NAND2_X1 U14614 ( .A1(n12267), .A2(n12311), .ZN(n12383) );
  XNOR2_X1 U14615 ( .A(n12784), .B(n12284), .ZN(n12268) );
  XNOR2_X1 U14616 ( .A(n12268), .B(n12675), .ZN(n12382) );
  INV_X1 U14617 ( .A(n12268), .ZN(n12269) );
  NAND2_X1 U14618 ( .A1(n12269), .A2(n12675), .ZN(n12270) );
  XNOR2_X1 U14619 ( .A(n12341), .B(n12284), .ZN(n12272) );
  XNOR2_X1 U14620 ( .A(n12272), .B(n12642), .ZN(n12337) );
  NAND2_X1 U14621 ( .A1(n12272), .A2(n12642), .ZN(n12273) );
  XNOR2_X1 U14622 ( .A(n12838), .B(n12284), .ZN(n12371) );
  AOI22_X1 U14623 ( .A1(n12371), .A2(n12630), .B1(n6538), .B2(n12444), .ZN(
        n12274) );
  XNOR2_X1 U14624 ( .A(n12403), .B(n11386), .ZN(n12301) );
  INV_X1 U14625 ( .A(n12301), .ZN(n12302) );
  NAND3_X1 U14626 ( .A1(n12274), .A2(n12654), .A3(n12302), .ZN(n12279) );
  INV_X1 U14627 ( .A(n12371), .ZN(n12277) );
  OAI21_X1 U14628 ( .B1(n6538), .B2(n12444), .A(n12630), .ZN(n12276) );
  NOR3_X1 U14629 ( .A1(n6538), .A2(n12444), .A3(n12630), .ZN(n12275) );
  AOI21_X1 U14630 ( .B1(n12277), .B2(n12276), .A(n12275), .ZN(n12278) );
  XNOR2_X1 U14631 ( .A(n12602), .B(n11386), .ZN(n12282) );
  XNOR2_X1 U14632 ( .A(n12282), .B(n12614), .ZN(n12345) );
  INV_X1 U14633 ( .A(n12282), .ZN(n12283) );
  XNOR2_X1 U14634 ( .A(n12591), .B(n12284), .ZN(n12285) );
  XNOR2_X1 U14635 ( .A(n12285), .B(n12570), .ZN(n12417) );
  OAI22_X1 U14636 ( .A1(n12416), .A2(n12417), .B1(n12285), .B2(n12570), .ZN(
        n12323) );
  XOR2_X1 U14637 ( .A(n12322), .B(n12323), .Z(n12291) );
  AOI22_X1 U14638 ( .A1(n12570), .A2(n12418), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12287) );
  NAND2_X1 U14639 ( .A1(n12437), .A2(n12575), .ZN(n12286) );
  OAI211_X1 U14640 ( .C1(n12442), .C2(n12421), .A(n12287), .B(n12286), .ZN(
        n12288) );
  AOI21_X1 U14641 ( .B1(n12289), .B2(n12424), .A(n12288), .ZN(n12290) );
  OAI21_X1 U14642 ( .B1(n12291), .B2(n12439), .A(n12290), .ZN(P3_U3154) );
  XNOR2_X1 U14643 ( .A(n12293), .B(n12292), .ZN(n12300) );
  NOR2_X1 U14644 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12294), .ZN(n12479) );
  AOI21_X1 U14645 ( .B1(n12418), .B2(n12446), .A(n12479), .ZN(n12295) );
  OAI21_X1 U14646 ( .B1(n12357), .B2(n12421), .A(n12295), .ZN(n12297) );
  NOR2_X1 U14647 ( .A1(n12866), .A2(n12434), .ZN(n12296) );
  AOI211_X1 U14648 ( .C1(n12298), .C2(n12437), .A(n12297), .B(n12296), .ZN(
        n12299) );
  OAI21_X1 U14649 ( .B1(n12300), .B2(n12439), .A(n12299), .ZN(P3_U3155) );
  XNOR2_X1 U14650 ( .A(n12303), .B(n12301), .ZN(n12399) );
  AND2_X1 U14651 ( .A1(n12303), .A2(n12302), .ZN(n12304) );
  XNOR2_X1 U14652 ( .A(n12370), .B(n12643), .ZN(n12309) );
  NAND2_X1 U14653 ( .A1(n12437), .A2(n12633), .ZN(n12306) );
  AOI22_X1 U14654 ( .A1(n12630), .A2(n12431), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12305) );
  OAI211_X1 U14655 ( .C1(n12654), .C2(n12433), .A(n12306), .B(n12305), .ZN(
        n12307) );
  AOI21_X1 U14656 ( .B1(n12771), .B2(n12424), .A(n12307), .ZN(n12308) );
  OAI21_X1 U14657 ( .B1(n12309), .B2(n12439), .A(n12308), .ZN(P3_U3156) );
  NAND2_X1 U14658 ( .A1(n12311), .A2(n12310), .ZN(n12313) );
  XOR2_X1 U14659 ( .A(n12313), .B(n12312), .Z(n12319) );
  NAND2_X1 U14660 ( .A1(n12418), .A2(n12711), .ZN(n12315) );
  OAI211_X1 U14661 ( .C1(n12653), .C2(n12421), .A(n12315), .B(n12314), .ZN(
        n12317) );
  NOR2_X1 U14662 ( .A1(n12683), .A2(n12434), .ZN(n12316) );
  AOI211_X1 U14663 ( .C1(n12681), .C2(n12437), .A(n12317), .B(n12316), .ZN(
        n12318) );
  OAI21_X1 U14664 ( .B1(n12319), .B2(n12439), .A(n12318), .ZN(P3_U3159) );
  INV_X1 U14665 ( .A(n12320), .ZN(n12321) );
  AOI22_X1 U14666 ( .A1(n12323), .A2(n12322), .B1(n12422), .B2(n12321), .ZN(
        n12325) );
  XNOR2_X1 U14667 ( .A(n9797), .B(n11386), .ZN(n12324) );
  XNOR2_X1 U14668 ( .A(n12325), .B(n12324), .ZN(n12333) );
  OAI22_X1 U14669 ( .A1(n12422), .A2(n12433), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12326), .ZN(n12329) );
  NOR2_X1 U14670 ( .A1(n12327), .A2(n12421), .ZN(n12328) );
  AOI211_X1 U14671 ( .C1(n12437), .C2(n12556), .A(n12329), .B(n12328), .ZN(
        n12332) );
  NAND2_X1 U14672 ( .A1(n12330), .A2(n12424), .ZN(n12331) );
  OAI211_X1 U14673 ( .C1(n12333), .C2(n12439), .A(n12332), .B(n12331), .ZN(
        P3_U3160) );
  INV_X1 U14674 ( .A(n12334), .ZN(n12335) );
  AOI21_X1 U14675 ( .B1(n12337), .B2(n12336), .A(n12335), .ZN(n12343) );
  NAND2_X1 U14676 ( .A1(n12437), .A2(n12657), .ZN(n12339) );
  AOI22_X1 U14677 ( .A1(n12675), .A2(n12418), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12338) );
  OAI211_X1 U14678 ( .C1(n12654), .C2(n12421), .A(n12339), .B(n12338), .ZN(
        n12340) );
  AOI21_X1 U14679 ( .B1(n12341), .B2(n12424), .A(n12340), .ZN(n12342) );
  OAI21_X1 U14680 ( .B1(n12343), .B2(n12439), .A(n12342), .ZN(P3_U3163) );
  XOR2_X1 U14681 ( .A(n12345), .B(n12344), .Z(n12350) );
  NAND2_X1 U14682 ( .A1(n12437), .A2(n12603), .ZN(n12347) );
  AOI22_X1 U14683 ( .A1(n12630), .A2(n12418), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12346) );
  OAI211_X1 U14684 ( .C1(n12596), .C2(n12421), .A(n12347), .B(n12346), .ZN(
        n12348) );
  AOI21_X1 U14685 ( .B1(n12602), .B2(n12424), .A(n12348), .ZN(n12349) );
  OAI21_X1 U14686 ( .B1(n12350), .B2(n12439), .A(n12349), .ZN(P3_U3165) );
  XNOR2_X1 U14687 ( .A(n12352), .B(n12710), .ZN(n12353) );
  XNOR2_X1 U14688 ( .A(n12351), .B(n12353), .ZN(n12360) );
  NAND2_X1 U14689 ( .A1(n12437), .A2(n12730), .ZN(n12356) );
  NOR2_X1 U14690 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12354), .ZN(n12495) );
  AOI21_X1 U14691 ( .B1(n12431), .B2(n12725), .A(n12495), .ZN(n12355) );
  OAI211_X1 U14692 ( .C1(n12357), .C2(n12433), .A(n12356), .B(n12355), .ZN(
        n12358) );
  AOI21_X1 U14693 ( .B1(n12803), .B2(n12424), .A(n12358), .ZN(n12359) );
  OAI21_X1 U14694 ( .B1(n12360), .B2(n12439), .A(n12359), .ZN(P3_U3166) );
  AOI21_X1 U14695 ( .B1(n12361), .B2(n12362), .A(n12439), .ZN(n12364) );
  NAND2_X1 U14696 ( .A1(n12364), .A2(n12363), .ZN(n12368) );
  NAND2_X1 U14697 ( .A1(n12418), .A2(n12710), .ZN(n12365) );
  NAND2_X1 U14698 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12509)
         );
  OAI211_X1 U14699 ( .C1(n12407), .C2(n12421), .A(n12365), .B(n12509), .ZN(
        n12366) );
  AOI21_X1 U14700 ( .B1(n12437), .B2(n12716), .A(n12366), .ZN(n12367) );
  OAI211_X1 U14701 ( .C1(n12434), .C2(n12857), .A(n12368), .B(n12367), .ZN(
        P3_U3168) );
  XNOR2_X1 U14702 ( .A(n12371), .B(n12630), .ZN(n12372) );
  XNOR2_X1 U14703 ( .A(n12373), .B(n12372), .ZN(n12379) );
  NAND2_X1 U14704 ( .A1(n12437), .A2(n12618), .ZN(n12375) );
  AOI22_X1 U14705 ( .A1(n12583), .A2(n12431), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12374) );
  OAI211_X1 U14706 ( .C1(n12643), .C2(n12433), .A(n12375), .B(n12374), .ZN(
        n12376) );
  AOI21_X1 U14707 ( .B1(n12377), .B2(n12424), .A(n12376), .ZN(n12378) );
  OAI21_X1 U14708 ( .B1(n12379), .B2(n12439), .A(n12378), .ZN(P3_U3169) );
  INV_X1 U14709 ( .A(n12784), .ZN(n12671) );
  OAI211_X1 U14710 ( .C1(n12383), .C2(n12382), .A(n12380), .B(n12381), .ZN(
        n12387) );
  AOI22_X1 U14711 ( .A1(n12431), .A2(n12663), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12384) );
  OAI21_X1 U14712 ( .B1(n12411), .B2(n12433), .A(n12384), .ZN(n12385) );
  AOI21_X1 U14713 ( .B1(n12437), .B2(n12669), .A(n12385), .ZN(n12386) );
  OAI211_X1 U14714 ( .C1(n12671), .C2(n12434), .A(n12387), .B(n12386), .ZN(
        P3_U3173) );
  XNOR2_X1 U14715 ( .A(n12390), .B(n12389), .ZN(n12391) );
  XNOR2_X1 U14716 ( .A(n12388), .B(n12391), .ZN(n12398) );
  NAND2_X1 U14717 ( .A1(n12437), .A2(n12392), .ZN(n12394) );
  AND2_X1 U14718 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n15021) );
  AOI21_X1 U14719 ( .B1(n12418), .B2(n14452), .A(n15021), .ZN(n12393) );
  OAI211_X1 U14720 ( .C1(n12739), .C2(n12421), .A(n12394), .B(n12393), .ZN(
        n12395) );
  AOI21_X1 U14721 ( .B1(n12396), .B2(n12424), .A(n12395), .ZN(n12397) );
  OAI21_X1 U14722 ( .B1(n12398), .B2(n12439), .A(n12397), .ZN(P3_U3174) );
  XNOR2_X1 U14723 ( .A(n12399), .B(n12629), .ZN(n12405) );
  NAND2_X1 U14724 ( .A1(n12437), .A2(n12646), .ZN(n12401) );
  AOI22_X1 U14725 ( .A1(n12418), .A2(n12663), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12400) );
  OAI211_X1 U14726 ( .C1(n12643), .C2(n12421), .A(n12401), .B(n12400), .ZN(
        n12402) );
  AOI21_X1 U14727 ( .B1(n12403), .B2(n12424), .A(n12402), .ZN(n12404) );
  OAI21_X1 U14728 ( .B1(n12405), .B2(n12439), .A(n12404), .ZN(P3_U3175) );
  XNOR2_X1 U14729 ( .A(n12408), .B(n12407), .ZN(n12409) );
  XNOR2_X1 U14730 ( .A(n12406), .B(n12409), .ZN(n12415) );
  NAND2_X1 U14731 ( .A1(n12418), .A2(n12725), .ZN(n12410) );
  NAND2_X1 U14732 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12531)
         );
  OAI211_X1 U14733 ( .C1(n12411), .C2(n12421), .A(n12410), .B(n12531), .ZN(
        n12413) );
  NOR2_X1 U14734 ( .A1(n12793), .A2(n12434), .ZN(n12412) );
  AOI211_X1 U14735 ( .C1(n12700), .C2(n12437), .A(n12413), .B(n12412), .ZN(
        n12414) );
  OAI21_X1 U14736 ( .B1(n12415), .B2(n12439), .A(n12414), .ZN(P3_U3178) );
  XOR2_X1 U14737 ( .A(n12417), .B(n12416), .Z(n12426) );
  NAND2_X1 U14738 ( .A1(n12437), .A2(n12589), .ZN(n12420) );
  AOI22_X1 U14739 ( .A1(n12583), .A2(n12418), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12419) );
  OAI211_X1 U14740 ( .C1(n12422), .C2(n12421), .A(n12420), .B(n12419), .ZN(
        n12423) );
  AOI21_X1 U14741 ( .B1(n12758), .B2(n12424), .A(n12423), .ZN(n12425) );
  OAI21_X1 U14742 ( .B1(n12426), .B2(n12439), .A(n12425), .ZN(P3_U3180) );
  INV_X1 U14743 ( .A(n12428), .ZN(n12429) );
  AOI21_X1 U14744 ( .B1(n12427), .B2(n12430), .A(n12429), .ZN(n12440) );
  AND2_X1 U14745 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n14448) );
  AOI21_X1 U14746 ( .B1(n12431), .B2(n12710), .A(n14448), .ZN(n12432) );
  OAI21_X1 U14747 ( .B1(n12739), .B2(n12433), .A(n12432), .ZN(n12436) );
  NOR2_X1 U14748 ( .A1(n12862), .A2(n12434), .ZN(n12435) );
  AOI211_X1 U14749 ( .C1(n12742), .C2(n12437), .A(n12436), .B(n12435), .ZN(
        n12438) );
  OAI21_X1 U14750 ( .B1(n12440), .B2(n12439), .A(n12438), .ZN(P3_U3181) );
  MUX2_X1 U14751 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(n12441), .S(P3_U3897), .Z(
        P3_U3521) );
  INV_X1 U14752 ( .A(n12442), .ZN(n12571) );
  MUX2_X1 U14753 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12571), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14754 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12584), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14755 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12570), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14756 ( .A(n12583), .B(P3_DATAO_REG_25__SCAN_IN), .S(n12443), .Z(
        P3_U3516) );
  MUX2_X1 U14757 ( .A(n12630), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12443), .Z(
        P3_U3515) );
  MUX2_X1 U14758 ( .A(n12444), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12443), .Z(
        P3_U3514) );
  MUX2_X1 U14759 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12629), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14760 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12663), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14761 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12675), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14762 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n12691), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14763 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12711), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14764 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12725), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14765 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12710), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14766 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12724), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14767 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12445), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14768 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12446), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14769 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n14452), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14770 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12447), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14771 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n15039), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14772 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n15040), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14773 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12448), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14774 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12449), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14775 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12450), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14776 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12451), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14777 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n15078), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14778 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n12452), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U14779 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n15077), .S(P3_U3897), .Z(
        P3_U3491) );
  XNOR2_X1 U14780 ( .A(n12454), .B(n12453), .ZN(n12467) );
  XNOR2_X1 U14781 ( .A(n12456), .B(n12455), .ZN(n12461) );
  NAND2_X1 U14782 ( .A1(n14960), .A2(n12457), .ZN(n12460) );
  AOI21_X1 U14783 ( .B1(n14983), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n12458), 
        .ZN(n12459) );
  OAI211_X1 U14784 ( .C1(n12461), .C2(n15015), .A(n12460), .B(n12459), .ZN(
        n12466) );
  AOI21_X1 U14785 ( .B1(n6547), .B2(n12463), .A(n12462), .ZN(n12464) );
  NOR2_X1 U14786 ( .A1(n12464), .A2(n15017), .ZN(n12465) );
  AOI211_X1 U14787 ( .C1(n12467), .C2(n12472), .A(n12466), .B(n12465), .ZN(
        n12468) );
  INV_X1 U14788 ( .A(n12468), .ZN(P3_U3194) );
  AOI21_X1 U14789 ( .B1(n6548), .B2(n12470), .A(n12469), .ZN(n12487) );
  XNOR2_X1 U14790 ( .A(n6541), .B(n12471), .ZN(n12473) );
  NAND2_X1 U14791 ( .A1(n12473), .A2(n12472), .ZN(n12486) );
  INV_X1 U14792 ( .A(n12474), .ZN(n12484) );
  NAND2_X1 U14793 ( .A1(n14983), .A2(P3_ADDR_REG_14__SCAN_IN), .ZN(n12482) );
  INV_X1 U14794 ( .A(n12475), .ZN(n12476) );
  OAI211_X1 U14795 ( .C1(n12478), .C2(n12477), .A(n14963), .B(n12476), .ZN(
        n12481) );
  INV_X1 U14796 ( .A(n12479), .ZN(n12480) );
  NAND3_X1 U14797 ( .A1(n12482), .A2(n12481), .A3(n12480), .ZN(n12483) );
  AOI21_X1 U14798 ( .B1(n14960), .B2(n12484), .A(n12483), .ZN(n12485) );
  OAI211_X1 U14799 ( .C1(n12487), .C2(n15017), .A(n12486), .B(n12485), .ZN(
        P3_U3196) );
  AOI21_X1 U14800 ( .B1(n6531), .B2(n12489), .A(n12488), .ZN(n12505) );
  INV_X1 U14801 ( .A(n12490), .ZN(n12491) );
  NAND2_X1 U14802 ( .A1(n12492), .A2(n12491), .ZN(n12493) );
  XNOR2_X1 U14803 ( .A(n12494), .B(n12493), .ZN(n12503) );
  AOI21_X1 U14804 ( .B1(n14983), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n12495), 
        .ZN(n12496) );
  OAI21_X1 U14805 ( .B1(n15008), .B2(n12497), .A(n12496), .ZN(n12502) );
  AOI21_X1 U14806 ( .B1(n6484), .B2(n12499), .A(n12498), .ZN(n12500) );
  NOR2_X1 U14807 ( .A1(n12500), .A2(n15017), .ZN(n12501) );
  AOI211_X1 U14808 ( .C1(n14963), .C2(n12503), .A(n12502), .B(n12501), .ZN(
        n12504) );
  OAI21_X1 U14809 ( .B1(n12505), .B2(n15023), .A(n12504), .ZN(P3_U3198) );
  AOI21_X1 U14810 ( .B1(n12508), .B2(n12507), .A(n12506), .ZN(n12522) );
  INV_X1 U14811 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n12510) );
  OAI21_X1 U14812 ( .B1(n15005), .B2(n12510), .A(n12509), .ZN(n12515) );
  AOI211_X1 U14813 ( .C1(n12513), .C2(n12512), .A(n12511), .B(n15015), .ZN(
        n12514) );
  AOI211_X1 U14814 ( .C1(n14960), .C2(n12516), .A(n12515), .B(n12514), .ZN(
        n12521) );
  AOI21_X1 U14815 ( .B1(n12801), .B2(n12518), .A(n12517), .ZN(n12519) );
  OR2_X1 U14816 ( .A1(n12519), .A2(n15017), .ZN(n12520) );
  OAI211_X1 U14817 ( .C1(n12522), .C2(n15023), .A(n12521), .B(n12520), .ZN(
        P3_U3199) );
  AOI21_X1 U14818 ( .B1(n12525), .B2(n12524), .A(n12523), .ZN(n12538) );
  INV_X1 U14819 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n14429) );
  OAI21_X1 U14820 ( .B1(n12528), .B2(n12527), .A(n12526), .ZN(n12529) );
  NAND2_X1 U14821 ( .A1(n14963), .A2(n12529), .ZN(n12530) );
  OAI211_X1 U14822 ( .C1(n15005), .C2(n14429), .A(n12531), .B(n12530), .ZN(
        n12535) );
  OAI21_X1 U14823 ( .B1(n12538), .B2(n15023), .A(n12537), .ZN(P3_U3200) );
  NOR2_X1 U14824 ( .A1(n12540), .A2(n12539), .ZN(n12819) );
  NOR2_X1 U14825 ( .A1(n12541), .A2(n15056), .ZN(n12550) );
  AOI21_X1 U14826 ( .B1(n12819), .B2(n15094), .A(n12550), .ZN(n12545) );
  NAND2_X1 U14827 ( .A1(n15071), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12542) );
  OAI211_X1 U14828 ( .C1(n12543), .C2(n12744), .A(n12545), .B(n12542), .ZN(
        P3_U3202) );
  NAND2_X1 U14829 ( .A1(n15071), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n12544) );
  OAI211_X1 U14830 ( .C1(n12753), .C2(n12744), .A(n12545), .B(n12544), .ZN(
        P3_U3203) );
  INV_X1 U14831 ( .A(n12546), .ZN(n12554) );
  NAND2_X1 U14832 ( .A1(n12547), .A2(n15094), .ZN(n12552) );
  NOR2_X1 U14833 ( .A1(n12548), .A2(n12744), .ZN(n12549) );
  AOI211_X1 U14834 ( .C1(n15071), .C2(P3_REG2_REG_29__SCAN_IN), .A(n12550), 
        .B(n12549), .ZN(n12551) );
  OAI211_X1 U14835 ( .C1(n12554), .C2(n12553), .A(n12552), .B(n12551), .ZN(
        P3_U3204) );
  INV_X1 U14836 ( .A(n12555), .ZN(n12562) );
  AOI22_X1 U14837 ( .A1(n12556), .A2(n15090), .B1(P3_REG2_REG_28__SCAN_IN), 
        .B2(n15071), .ZN(n12557) );
  OAI21_X1 U14838 ( .B1(n12558), .B2(n12744), .A(n12557), .ZN(n12559) );
  AOI21_X1 U14839 ( .B1(n12560), .B2(n14458), .A(n12559), .ZN(n12561) );
  OAI21_X1 U14840 ( .B1(n12562), .B2(n15071), .A(n12561), .ZN(P3_U3205) );
  INV_X1 U14841 ( .A(n12563), .ZN(n12565) );
  OAI21_X1 U14842 ( .B1(n12568), .B2(n12567), .A(n12566), .ZN(n12569) );
  NAND2_X1 U14843 ( .A1(n12569), .A2(n15074), .ZN(n12573) );
  AOI22_X1 U14844 ( .A1(n12571), .A2(n15079), .B1(n15076), .B2(n12570), .ZN(
        n12572) );
  OAI211_X1 U14845 ( .C1(n15067), .C2(n12574), .A(n12573), .B(n12572), .ZN(
        n12754) );
  INV_X1 U14846 ( .A(n12754), .ZN(n12579) );
  INV_X1 U14847 ( .A(n12574), .ZN(n12755) );
  AOI22_X1 U14848 ( .A1(n12575), .A2(n15090), .B1(P3_REG2_REG_27__SCAN_IN), 
        .B2(n15071), .ZN(n12576) );
  OAI21_X1 U14849 ( .B1(n12829), .B2(n12744), .A(n12576), .ZN(n12577) );
  AOI21_X1 U14850 ( .B1(n12755), .B2(n15091), .A(n12577), .ZN(n12578) );
  OAI21_X1 U14851 ( .B1(n12579), .B2(n15071), .A(n12578), .ZN(P3_U3206) );
  XNOR2_X1 U14852 ( .A(n6476), .B(n12580), .ZN(n12587) );
  XNOR2_X1 U14853 ( .A(n12582), .B(n12581), .ZN(n12588) );
  AOI22_X1 U14854 ( .A1(n12584), .A2(n15079), .B1(n15076), .B2(n12583), .ZN(
        n12585) );
  OAI21_X1 U14855 ( .B1(n12588), .B2(n15067), .A(n12585), .ZN(n12586) );
  AOI21_X1 U14856 ( .B1(n12587), .B2(n15074), .A(n12586), .ZN(n12761) );
  INV_X1 U14857 ( .A(n12588), .ZN(n12759) );
  AOI22_X1 U14858 ( .A1(n12589), .A2(n15090), .B1(P3_REG2_REG_26__SCAN_IN), 
        .B2(n15071), .ZN(n12590) );
  OAI21_X1 U14859 ( .B1(n12591), .B2(n12744), .A(n12590), .ZN(n12592) );
  AOI21_X1 U14860 ( .B1(n12759), .B2(n15091), .A(n12592), .ZN(n12593) );
  OAI21_X1 U14861 ( .B1(n12761), .B2(n15071), .A(n12593), .ZN(P3_U3207) );
  XNOR2_X1 U14862 ( .A(n12594), .B(n12599), .ZN(n12764) );
  OAI22_X1 U14863 ( .A1(n12596), .A2(n15059), .B1(n12595), .B2(n15061), .ZN(
        n12601) );
  AOI211_X1 U14864 ( .C1(n12599), .C2(n12598), .A(n12736), .B(n12597), .ZN(
        n12600) );
  AOI211_X1 U14865 ( .C1(n15083), .C2(n12764), .A(n12601), .B(n12600), .ZN(
        n12762) );
  INV_X1 U14866 ( .A(n12602), .ZN(n12834) );
  AOI22_X1 U14867 ( .A1(n12603), .A2(n15090), .B1(P3_REG2_REG_25__SCAN_IN), 
        .B2(n15071), .ZN(n12604) );
  OAI21_X1 U14868 ( .B1(n12834), .B2(n12744), .A(n12604), .ZN(n12605) );
  AOI21_X1 U14869 ( .B1(n12764), .B2(n15091), .A(n12605), .ZN(n12606) );
  OAI21_X1 U14870 ( .B1(n12762), .B2(n15071), .A(n12606), .ZN(P3_U3208) );
  XNOR2_X1 U14871 ( .A(n12608), .B(n12607), .ZN(n12617) );
  INV_X1 U14872 ( .A(n12625), .ZN(n12611) );
  OAI21_X1 U14873 ( .B1(n12611), .B2(n12610), .A(n12609), .ZN(n12613) );
  NAND2_X1 U14874 ( .A1(n12613), .A2(n12612), .ZN(n12768) );
  OAI22_X1 U14875 ( .A1(n12614), .A2(n15059), .B1(n12643), .B2(n15061), .ZN(
        n12615) );
  AOI21_X1 U14876 ( .B1(n12768), .B2(n15083), .A(n12615), .ZN(n12616) );
  OAI21_X1 U14877 ( .B1(n12617), .B2(n12736), .A(n12616), .ZN(n12767) );
  INV_X1 U14878 ( .A(n12767), .ZN(n12622) );
  AOI22_X1 U14879 ( .A1(n15071), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n12618), 
        .B2(n15090), .ZN(n12619) );
  OAI21_X1 U14880 ( .B1(n12838), .B2(n12744), .A(n12619), .ZN(n12620) );
  AOI21_X1 U14881 ( .B1(n12768), .B2(n15091), .A(n12620), .ZN(n12621) );
  OAI21_X1 U14882 ( .B1(n12622), .B2(n15071), .A(n12621), .ZN(P3_U3209) );
  OR2_X1 U14883 ( .A1(n12623), .A2(n12626), .ZN(n12624) );
  NAND2_X1 U14884 ( .A1(n12625), .A2(n12624), .ZN(n12634) );
  XNOR2_X1 U14885 ( .A(n12627), .B(n12626), .ZN(n12628) );
  NAND2_X1 U14886 ( .A1(n12628), .A2(n15074), .ZN(n12632) );
  AOI22_X1 U14887 ( .A1(n12630), .A2(n15079), .B1(n15076), .B2(n12629), .ZN(
        n12631) );
  OAI211_X1 U14888 ( .C1(n15067), .C2(n12634), .A(n12632), .B(n12631), .ZN(
        n12772) );
  NAND2_X1 U14889 ( .A1(n12772), .A2(n15094), .ZN(n12639) );
  AOI22_X1 U14890 ( .A1(n15071), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n15090), 
        .B2(n12633), .ZN(n12638) );
  INV_X1 U14891 ( .A(n12634), .ZN(n12773) );
  NAND2_X1 U14892 ( .A1(n12773), .A2(n15091), .ZN(n12637) );
  NAND2_X1 U14893 ( .A1(n12771), .A2(n12635), .ZN(n12636) );
  NAND4_X1 U14894 ( .A1(n12639), .A2(n12638), .A3(n12637), .A4(n12636), .ZN(
        P3_U3210) );
  XOR2_X1 U14895 ( .A(n12640), .B(n12645), .Z(n12641) );
  OAI222_X1 U14896 ( .A1(n15059), .A2(n12643), .B1(n15061), .B2(n12642), .C1(
        n12736), .C2(n12641), .ZN(n12776) );
  INV_X1 U14897 ( .A(n12776), .ZN(n12650) );
  XOR2_X1 U14898 ( .A(n12645), .B(n12644), .Z(n12777) );
  AOI22_X1 U14899 ( .A1(n15071), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15090), 
        .B2(n12646), .ZN(n12647) );
  OAI21_X1 U14900 ( .B1(n12846), .B2(n12744), .A(n12647), .ZN(n12648) );
  AOI21_X1 U14901 ( .B1(n12777), .B2(n14458), .A(n12648), .ZN(n12649) );
  OAI21_X1 U14902 ( .B1(n12650), .B2(n15071), .A(n12649), .ZN(P3_U3211) );
  XNOR2_X1 U14903 ( .A(n12651), .B(n12655), .ZN(n12652) );
  OAI222_X1 U14904 ( .A1(n15059), .A2(n12654), .B1(n15061), .B2(n12653), .C1(
        n12736), .C2(n12652), .ZN(n12780) );
  INV_X1 U14905 ( .A(n12780), .ZN(n12661) );
  XOR2_X1 U14906 ( .A(n12656), .B(n12655), .Z(n12781) );
  AOI22_X1 U14907 ( .A1(n15071), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15090), 
        .B2(n12657), .ZN(n12658) );
  OAI21_X1 U14908 ( .B1(n12850), .B2(n12744), .A(n12658), .ZN(n12659) );
  AOI21_X1 U14909 ( .B1(n12781), .B2(n14458), .A(n12659), .ZN(n12660) );
  OAI21_X1 U14910 ( .B1(n12661), .B2(n15071), .A(n12660), .ZN(P3_U3212) );
  XNOR2_X1 U14911 ( .A(n12662), .B(n8718), .ZN(n12664) );
  AOI222_X1 U14912 ( .A1(n15074), .A2(n12664), .B1(n12663), .B2(n15079), .C1(
        n12691), .C2(n15076), .ZN(n12787) );
  INV_X1 U14913 ( .A(n12665), .ZN(n12666) );
  AOI21_X1 U14914 ( .B1(n12668), .B2(n12667), .A(n12666), .ZN(n12785) );
  AOI22_X1 U14915 ( .A1(n15071), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15090), 
        .B2(n12669), .ZN(n12670) );
  OAI21_X1 U14916 ( .B1(n12671), .B2(n12744), .A(n12670), .ZN(n12672) );
  AOI21_X1 U14917 ( .B1(n12785), .B2(n14458), .A(n12672), .ZN(n12673) );
  OAI21_X1 U14918 ( .B1(n12787), .B2(n15071), .A(n12673), .ZN(P3_U3213) );
  XNOR2_X1 U14919 ( .A(n12674), .B(n12680), .ZN(n12676) );
  AOI222_X1 U14920 ( .A1(n15074), .A2(n12676), .B1(n12675), .B2(n15079), .C1(
        n12711), .C2(n15076), .ZN(n12790) );
  INV_X1 U14921 ( .A(n12677), .ZN(n12678) );
  AOI21_X1 U14922 ( .B1(n12680), .B2(n12679), .A(n12678), .ZN(n12791) );
  INV_X1 U14923 ( .A(n12791), .ZN(n12685) );
  AOI22_X1 U14924 ( .A1(n15071), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15090), 
        .B2(n12681), .ZN(n12682) );
  OAI21_X1 U14925 ( .B1(n12683), .B2(n12744), .A(n12682), .ZN(n12684) );
  AOI21_X1 U14926 ( .B1(n12685), .B2(n14458), .A(n12684), .ZN(n12686) );
  OAI21_X1 U14927 ( .B1(n12790), .B2(n15071), .A(n12686), .ZN(P3_U3214) );
  NAND2_X1 U14928 ( .A1(n12688), .A2(n12687), .ZN(n12689) );
  NAND2_X1 U14929 ( .A1(n12690), .A2(n12689), .ZN(n12695) );
  NAND2_X1 U14930 ( .A1(n12691), .A2(n15079), .ZN(n12692) );
  OAI21_X1 U14931 ( .B1(n12693), .B2(n15061), .A(n12692), .ZN(n12694) );
  AOI21_X1 U14932 ( .B1(n12695), .B2(n15074), .A(n12694), .ZN(n12797) );
  NAND2_X1 U14933 ( .A1(n12697), .A2(n12696), .ZN(n12698) );
  AOI22_X1 U14934 ( .A1(n15071), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n15090), 
        .B2(n12700), .ZN(n12701) );
  OAI21_X1 U14935 ( .B1(n12793), .B2(n12744), .A(n12701), .ZN(n12702) );
  AOI21_X1 U14936 ( .B1(n12795), .B2(n14458), .A(n12702), .ZN(n12703) );
  OAI21_X1 U14937 ( .B1(n12797), .B2(n15071), .A(n12703), .ZN(P3_U3215) );
  NAND2_X1 U14938 ( .A1(n12735), .A2(n12704), .ZN(n12706) );
  NAND2_X1 U14939 ( .A1(n12706), .A2(n12705), .ZN(n12709) );
  OAI211_X1 U14940 ( .C1(n12709), .C2(n12708), .A(n12707), .B(n15074), .ZN(
        n12713) );
  AOI22_X1 U14941 ( .A1(n12711), .A2(n15079), .B1(n12710), .B2(n15076), .ZN(
        n12712) );
  AND2_X1 U14942 ( .A1(n12713), .A2(n12712), .ZN(n12800) );
  XNOR2_X1 U14943 ( .A(n12715), .B(n9831), .ZN(n12798) );
  AOI22_X1 U14944 ( .A1(n15071), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15090), 
        .B2(n12716), .ZN(n12717) );
  OAI21_X1 U14945 ( .B1(n12857), .B2(n12744), .A(n12717), .ZN(n12718) );
  AOI21_X1 U14946 ( .B1(n12798), .B2(n14458), .A(n12718), .ZN(n12719) );
  OAI21_X1 U14947 ( .B1(n12800), .B2(n15071), .A(n12719), .ZN(P3_U3216) );
  NAND2_X1 U14948 ( .A1(n12735), .A2(n12720), .ZN(n12722) );
  NAND2_X1 U14949 ( .A1(n12722), .A2(n12721), .ZN(n12723) );
  XNOR2_X1 U14950 ( .A(n12723), .B(n12728), .ZN(n12726) );
  AOI222_X1 U14951 ( .A1(n15074), .A2(n12726), .B1(n12725), .B2(n15079), .C1(
        n12724), .C2(n15076), .ZN(n12806) );
  XNOR2_X1 U14952 ( .A(n12729), .B(n12728), .ZN(n12804) );
  AOI22_X1 U14953 ( .A1(n15071), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15090), 
        .B2(n12730), .ZN(n12731) );
  OAI21_X1 U14954 ( .B1(n12732), .B2(n12744), .A(n12731), .ZN(n12733) );
  AOI21_X1 U14955 ( .B1(n12804), .B2(n14458), .A(n12733), .ZN(n12734) );
  OAI21_X1 U14956 ( .B1(n12806), .B2(n15071), .A(n12734), .ZN(P3_U3217) );
  XOR2_X1 U14957 ( .A(n12735), .B(n12740), .Z(n12737) );
  OAI222_X1 U14958 ( .A1(n15061), .A2(n12739), .B1(n15059), .B2(n12738), .C1(
        n12737), .C2(n12736), .ZN(n12807) );
  INV_X1 U14959 ( .A(n12807), .ZN(n12747) );
  XNOR2_X1 U14960 ( .A(n12741), .B(n12740), .ZN(n12808) );
  AOI22_X1 U14961 ( .A1(n15071), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15090), 
        .B2(n12742), .ZN(n12743) );
  OAI21_X1 U14962 ( .B1(n12862), .B2(n12744), .A(n12743), .ZN(n12745) );
  AOI21_X1 U14963 ( .B1(n12808), .B2(n14458), .A(n12745), .ZN(n12746) );
  OAI21_X1 U14964 ( .B1(n12747), .B2(n15071), .A(n12746), .ZN(P3_U3218) );
  INV_X1 U14965 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n12750) );
  INV_X1 U14966 ( .A(n12817), .ZN(n12748) );
  NAND2_X1 U14967 ( .A1(n12818), .A2(n12748), .ZN(n12749) );
  NAND2_X1 U14968 ( .A1(n12819), .A2(n15166), .ZN(n12751) );
  OAI211_X1 U14969 ( .C1(n15166), .C2(n12750), .A(n12749), .B(n12751), .ZN(
        P3_U3490) );
  NAND2_X1 U14970 ( .A1(n15163), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n12752) );
  OAI211_X1 U14971 ( .C1(n12753), .C2(n12817), .A(n12752), .B(n12751), .ZN(
        P3_U3489) );
  MUX2_X1 U14972 ( .A(n12756), .B(n12826), .S(n15166), .Z(n12757) );
  AOI22_X1 U14973 ( .A1(n12759), .A2(n15143), .B1(n15084), .B2(n12758), .ZN(
        n12760) );
  NAND2_X1 U14974 ( .A1(n12761), .A2(n12760), .ZN(n12830) );
  MUX2_X1 U14975 ( .A(P3_REG1_REG_26__SCAN_IN), .B(n12830), .S(n15166), .Z(
        P3_U3485) );
  INV_X1 U14976 ( .A(n12762), .ZN(n12763) );
  AOI21_X1 U14977 ( .B1(n15143), .B2(n12764), .A(n12763), .ZN(n12831) );
  MUX2_X1 U14978 ( .A(n12765), .B(n12831), .S(n15166), .Z(n12766) );
  OAI21_X1 U14979 ( .B1(n12834), .B2(n12817), .A(n12766), .ZN(P3_U3484) );
  AOI21_X1 U14980 ( .B1(n15143), .B2(n12768), .A(n12767), .ZN(n12835) );
  MUX2_X1 U14981 ( .A(n12769), .B(n12835), .S(n15166), .Z(n12770) );
  OAI21_X1 U14982 ( .B1(n12838), .B2(n12817), .A(n12770), .ZN(P3_U3483) );
  INV_X1 U14983 ( .A(n12771), .ZN(n12842) );
  AOI21_X1 U14984 ( .B1(n15143), .B2(n12773), .A(n12772), .ZN(n12839) );
  MUX2_X1 U14985 ( .A(n12774), .B(n12839), .S(n15166), .Z(n12775) );
  OAI21_X1 U14986 ( .B1(n12842), .B2(n12817), .A(n12775), .ZN(P3_U3482) );
  AOI21_X1 U14987 ( .B1(n15099), .B2(n12777), .A(n12776), .ZN(n12843) );
  MUX2_X1 U14988 ( .A(n12778), .B(n12843), .S(n15166), .Z(n12779) );
  OAI21_X1 U14989 ( .B1(n12846), .B2(n12817), .A(n12779), .ZN(P3_U3481) );
  AOI21_X1 U14990 ( .B1(n12781), .B2(n15099), .A(n12780), .ZN(n12847) );
  MUX2_X1 U14991 ( .A(n12782), .B(n12847), .S(n15166), .Z(n12783) );
  OAI21_X1 U14992 ( .B1(n12850), .B2(n12817), .A(n12783), .ZN(P3_U3480) );
  AOI22_X1 U14993 ( .A1(n12785), .A2(n15099), .B1(n15084), .B2(n12784), .ZN(
        n12786) );
  NAND2_X1 U14994 ( .A1(n12787), .A2(n12786), .ZN(n12851) );
  MUX2_X1 U14995 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n12851), .S(n15166), .Z(
        P3_U3479) );
  INV_X1 U14996 ( .A(n15099), .ZN(n12792) );
  NAND2_X1 U14997 ( .A1(n12788), .A2(n15084), .ZN(n12789) );
  OAI211_X1 U14998 ( .C1(n12792), .C2(n12791), .A(n12790), .B(n12789), .ZN(
        n12852) );
  MUX2_X1 U14999 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n12852), .S(n15166), .Z(
        P3_U3478) );
  NOR2_X1 U15000 ( .A1(n12793), .A2(n15130), .ZN(n12794) );
  AOI21_X1 U15001 ( .B1(n12795), .B2(n15099), .A(n12794), .ZN(n12796) );
  NAND2_X1 U15002 ( .A1(n12797), .A2(n12796), .ZN(n12853) );
  MUX2_X1 U15003 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n12853), .S(n15166), .Z(
        P3_U3477) );
  NAND2_X1 U15004 ( .A1(n12798), .A2(n15099), .ZN(n12799) );
  MUX2_X1 U15005 ( .A(n12801), .B(n12854), .S(n15166), .Z(n12802) );
  OAI21_X1 U15006 ( .B1(n12817), .B2(n12857), .A(n12802), .ZN(P3_U3476) );
  AOI22_X1 U15007 ( .A1(n12804), .A2(n15099), .B1(n15084), .B2(n12803), .ZN(
        n12805) );
  NAND2_X1 U15008 ( .A1(n12806), .A2(n12805), .ZN(n12858) );
  MUX2_X1 U15009 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n12858), .S(n15166), .Z(
        P3_U3475) );
  AOI21_X1 U15010 ( .B1(n12808), .B2(n15099), .A(n12807), .ZN(n12859) );
  MUX2_X1 U15011 ( .A(n14440), .B(n12859), .S(n15166), .Z(n12809) );
  OAI21_X1 U15012 ( .B1(n12817), .B2(n12862), .A(n12809), .ZN(P3_U3474) );
  INV_X1 U15013 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12812) );
  AOI21_X1 U15014 ( .B1(n15099), .B2(n12811), .A(n12810), .ZN(n12863) );
  MUX2_X1 U15015 ( .A(n12812), .B(n12863), .S(n15166), .Z(n12813) );
  OAI21_X1 U15016 ( .B1(n12817), .B2(n12866), .A(n12813), .ZN(P3_U3473) );
  AOI21_X1 U15017 ( .B1(n12815), .B2(n15099), .A(n12814), .ZN(n12867) );
  MUX2_X1 U15018 ( .A(n15011), .B(n12867), .S(n15166), .Z(n12816) );
  OAI21_X1 U15019 ( .B1(n12817), .B2(n12870), .A(n12816), .ZN(P3_U3472) );
  INV_X1 U15020 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n14148) );
  INV_X1 U15021 ( .A(n12871), .ZN(n12821) );
  NAND2_X1 U15022 ( .A1(n12818), .A2(n12821), .ZN(n12820) );
  NAND2_X1 U15023 ( .A1(n12819), .A2(n15146), .ZN(n12823) );
  OAI211_X1 U15024 ( .C1(n15146), .C2(n14148), .A(n12820), .B(n12823), .ZN(
        P3_U3458) );
  INV_X1 U15025 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n12825) );
  NAND2_X1 U15026 ( .A1(n12822), .A2(n12821), .ZN(n12824) );
  OAI211_X1 U15027 ( .C1(n15146), .C2(n12825), .A(n12824), .B(n12823), .ZN(
        P3_U3457) );
  INV_X1 U15028 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n12827) );
  MUX2_X1 U15029 ( .A(n12827), .B(n12826), .S(n15146), .Z(n12828) );
  MUX2_X1 U15030 ( .A(P3_REG0_REG_26__SCAN_IN), .B(n12830), .S(n15146), .Z(
        P3_U3453) );
  INV_X1 U15031 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n12832) );
  MUX2_X1 U15032 ( .A(n12832), .B(n12831), .S(n15146), .Z(n12833) );
  OAI21_X1 U15033 ( .B1(n12834), .B2(n12871), .A(n12833), .ZN(P3_U3452) );
  INV_X1 U15034 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12836) );
  MUX2_X1 U15035 ( .A(n12836), .B(n12835), .S(n15146), .Z(n12837) );
  OAI21_X1 U15036 ( .B1(n12838), .B2(n12871), .A(n12837), .ZN(P3_U3451) );
  INV_X1 U15037 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12840) );
  MUX2_X1 U15038 ( .A(n12840), .B(n12839), .S(n15146), .Z(n12841) );
  OAI21_X1 U15039 ( .B1(n12842), .B2(n12871), .A(n12841), .ZN(P3_U3450) );
  INV_X1 U15040 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12844) );
  MUX2_X1 U15041 ( .A(n12844), .B(n12843), .S(n15146), .Z(n12845) );
  OAI21_X1 U15042 ( .B1(n12846), .B2(n12871), .A(n12845), .ZN(P3_U3449) );
  INV_X1 U15043 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12848) );
  MUX2_X1 U15044 ( .A(n12848), .B(n12847), .S(n15146), .Z(n12849) );
  OAI21_X1 U15045 ( .B1(n12850), .B2(n12871), .A(n12849), .ZN(P3_U3448) );
  MUX2_X1 U15046 ( .A(P3_REG0_REG_20__SCAN_IN), .B(n12851), .S(n15146), .Z(
        P3_U3447) );
  MUX2_X1 U15047 ( .A(P3_REG0_REG_19__SCAN_IN), .B(n12852), .S(n15146), .Z(
        P3_U3446) );
  MUX2_X1 U15048 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n12853), .S(n15146), .Z(
        P3_U3444) );
  INV_X1 U15049 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n12855) );
  MUX2_X1 U15050 ( .A(n12855), .B(n12854), .S(n15146), .Z(n12856) );
  OAI21_X1 U15051 ( .B1(n12871), .B2(n12857), .A(n12856), .ZN(P3_U3441) );
  MUX2_X1 U15052 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n12858), .S(n15146), .Z(
        P3_U3438) );
  INV_X1 U15053 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12860) );
  MUX2_X1 U15054 ( .A(n12860), .B(n12859), .S(n15146), .Z(n12861) );
  OAI21_X1 U15055 ( .B1(n12871), .B2(n12862), .A(n12861), .ZN(P3_U3435) );
  INV_X1 U15056 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12864) );
  MUX2_X1 U15057 ( .A(n12864), .B(n12863), .S(n15146), .Z(n12865) );
  OAI21_X1 U15058 ( .B1(n12871), .B2(n12866), .A(n12865), .ZN(P3_U3432) );
  INV_X1 U15059 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n12868) );
  MUX2_X1 U15060 ( .A(n12868), .B(n12867), .S(n15146), .Z(n12869) );
  OAI21_X1 U15061 ( .B1(n12871), .B2(n12870), .A(n12869), .ZN(P3_U3429) );
  NAND2_X1 U15062 ( .A1(n12873), .A2(n12872), .ZN(n12876) );
  NOR2_X1 U15063 ( .A1(n8479), .A2(P3_IR_REG_30__SCAN_IN), .ZN(n12874) );
  NAND3_X1 U15064 ( .A1(n8404), .A2(P3_STATE_REG_SCAN_IN), .A3(n12874), .ZN(
        n12875) );
  OAI211_X1 U15065 ( .C1(n12877), .C2(n12040), .A(n12876), .B(n12875), .ZN(
        P3_U3264) );
  INV_X1 U15066 ( .A(n12878), .ZN(n12879) );
  OAI222_X1 U15067 ( .A1(P3_U3151), .A2(n12882), .B1(n12040), .B2(n12881), 
        .C1(n12880), .C2(n12879), .ZN(P3_U3268) );
  MUX2_X1 U15068 ( .A(n12884), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  OAI211_X1 U15069 ( .C1(n12887), .C2(n12886), .A(n12885), .B(n12996), .ZN(
        n12893) );
  AOI22_X1 U15070 ( .A1(n13115), .A2(n12964), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12892) );
  OR2_X1 U15071 ( .A1(n13389), .A2(n12994), .ZN(n12891) );
  OAI22_X1 U15072 ( .A1(n12889), .A2(n12984), .B1(n12888), .B2(n12967), .ZN(
        n13111) );
  NAND2_X1 U15073 ( .A1(n13111), .A2(n12992), .ZN(n12890) );
  NAND4_X1 U15074 ( .A1(n12893), .A2(n12892), .A3(n12891), .A4(n12890), .ZN(
        P2_U3186) );
  INV_X1 U15075 ( .A(n12894), .ZN(n12901) );
  AOI22_X1 U15076 ( .A1(n12895), .A2(n12996), .B1(n12953), .B2(n13008), .ZN(
        n12900) );
  OAI22_X1 U15077 ( .A1(n12924), .A2(n12984), .B1(n12896), .B2(n12967), .ZN(
        n13167) );
  AOI22_X1 U15078 ( .A1(n13167), .A2(n12992), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12897) );
  OAI21_X1 U15079 ( .B1(n13171), .B2(n12990), .A(n12897), .ZN(n12898) );
  AOI21_X1 U15080 ( .B1(n6769), .B2(n12976), .A(n12898), .ZN(n12899) );
  OAI21_X1 U15081 ( .B1(n12901), .B2(n12900), .A(n12899), .ZN(P2_U3188) );
  INV_X1 U15082 ( .A(n12944), .ZN(n12912) );
  INV_X1 U15083 ( .A(n12902), .ZN(n12904) );
  NAND2_X1 U15084 ( .A1(n12904), .A2(n12903), .ZN(n12906) );
  AOI22_X1 U15085 ( .A1(n12912), .A2(n12907), .B1(n12906), .B2(n12905), .ZN(
        n12915) );
  NOR2_X1 U15086 ( .A1(n12990), .A2(n13230), .ZN(n12911) );
  AND2_X1 U15087 ( .A1(n13013), .A2(n12986), .ZN(n12908) );
  AOI21_X1 U15088 ( .B1(n13011), .B2(n12946), .A(n12908), .ZN(n13237) );
  OAI21_X1 U15089 ( .B1(n12961), .B2(n13237), .A(n12909), .ZN(n12910) );
  AOI211_X1 U15090 ( .C1(n13229), .C2(n12976), .A(n12911), .B(n12910), .ZN(
        n12914) );
  NAND3_X1 U15091 ( .A1(n12912), .A2(n12953), .A3(n13012), .ZN(n12913) );
  OAI211_X1 U15092 ( .C1(n12915), .C2(n12971), .A(n12914), .B(n12913), .ZN(
        P2_U3191) );
  OAI211_X1 U15093 ( .C1(n12918), .C2(n12917), .A(n12916), .B(n12996), .ZN(
        n12923) );
  INV_X1 U15094 ( .A(n13199), .ZN(n12921) );
  AOI22_X1 U15095 ( .A1(n13009), .A2(n12946), .B1(n12986), .B2(n13011), .ZN(
        n13205) );
  OAI22_X1 U15096 ( .A1(n13205), .A2(n12961), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12919), .ZN(n12920) );
  AOI21_X1 U15097 ( .B1(n12921), .B2(n12964), .A(n12920), .ZN(n12922) );
  OAI211_X1 U15098 ( .C1(n6767), .C2(n12994), .A(n12923), .B(n12922), .ZN(
        P2_U3195) );
  NOR3_X1 U15099 ( .A1(n12925), .A2(n12924), .A3(n12978), .ZN(n12930) );
  AOI21_X1 U15100 ( .B1(n12935), .B2(n12926), .A(n12971), .ZN(n12929) );
  INV_X1 U15101 ( .A(n12927), .ZN(n12928) );
  OAI21_X1 U15102 ( .B1(n12930), .B2(n12929), .A(n12928), .ZN(n12934) );
  AOI22_X1 U15103 ( .A1(n13005), .A2(n12946), .B1(n12986), .B2(n13007), .ZN(
        n13139) );
  OAI22_X1 U15104 ( .A1(n13139), .A2(n12961), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12931), .ZN(n12932) );
  AOI21_X1 U15105 ( .B1(n13143), .B2(n12964), .A(n12932), .ZN(n12933) );
  OAI211_X1 U15106 ( .C1(n13394), .C2(n12994), .A(n12934), .B(n12933), .ZN(
        P2_U3197) );
  OAI211_X1 U15107 ( .C1(n12937), .C2(n12936), .A(n12935), .B(n12996), .ZN(
        n12941) );
  OAI22_X1 U15108 ( .A1(n12979), .A2(n12984), .B1(n12959), .B2(n12967), .ZN(
        n13152) );
  AOI22_X1 U15109 ( .A1(n13152), .A2(n12992), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12938) );
  OAI21_X1 U15110 ( .B1(n13159), .B2(n12990), .A(n12938), .ZN(n12939) );
  AOI21_X1 U15111 ( .B1(n13162), .B2(n12976), .A(n12939), .ZN(n12940) );
  NAND2_X1 U15112 ( .A1(n12941), .A2(n12940), .ZN(P2_U3201) );
  INV_X1 U15113 ( .A(n12942), .ZN(n12943) );
  AOI21_X1 U15114 ( .B1(n12945), .B2(n12944), .A(n12943), .ZN(n12952) );
  NAND2_X1 U15115 ( .A1(n13010), .A2(n12946), .ZN(n12948) );
  NAND2_X1 U15116 ( .A1(n13012), .A2(n12986), .ZN(n12947) );
  NAND2_X1 U15117 ( .A1(n12948), .A2(n12947), .ZN(n13213) );
  AOI22_X1 U15118 ( .A1(n12992), .A2(n13213), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12949) );
  OAI21_X1 U15119 ( .B1(n13217), .B2(n12990), .A(n12949), .ZN(n12950) );
  AOI21_X1 U15120 ( .B1(n13406), .B2(n12976), .A(n12950), .ZN(n12951) );
  OAI21_X1 U15121 ( .B1(n12952), .B2(n12971), .A(n12951), .ZN(P2_U3205) );
  NAND2_X1 U15122 ( .A1(n12953), .A2(n13009), .ZN(n12957) );
  NAND2_X1 U15123 ( .A1(n12954), .A2(n12996), .ZN(n12956) );
  MUX2_X1 U15124 ( .A(n12957), .B(n12956), .S(n12955), .Z(n12966) );
  OAI22_X1 U15125 ( .A1(n12959), .A2(n12984), .B1(n12958), .B2(n12967), .ZN(
        n13182) );
  INV_X1 U15126 ( .A(n13182), .ZN(n12962) );
  OAI22_X1 U15127 ( .A1(n12962), .A2(n12961), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12960), .ZN(n12963) );
  AOI21_X1 U15128 ( .B1(n13190), .B2(n12964), .A(n12963), .ZN(n12965) );
  OAI211_X1 U15129 ( .C1(n13192), .C2(n12994), .A(n12966), .B(n12965), .ZN(
        P2_U3207) );
  OAI22_X1 U15130 ( .A1(n12969), .A2(n12984), .B1(n12968), .B2(n12967), .ZN(
        n13244) );
  NAND2_X1 U15131 ( .A1(n12992), .A2(n13244), .ZN(n12970) );
  NAND2_X1 U15132 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n14843)
         );
  OAI211_X1 U15133 ( .C1(n12990), .C2(n13247), .A(n12970), .B(n14843), .ZN(
        n12975) );
  AOI211_X1 U15134 ( .C1(n12973), .C2(n12972), .A(n12971), .B(n6550), .ZN(
        n12974) );
  AOI211_X1 U15135 ( .C1(n13359), .C2(n12976), .A(n12975), .B(n12974), .ZN(
        n12977) );
  INV_X1 U15136 ( .A(n12977), .ZN(P2_U3210) );
  NOR3_X1 U15137 ( .A1(n12980), .A2(n12979), .A3(n12978), .ZN(n12981) );
  AOI21_X1 U15138 ( .B1(n12927), .B2(n12996), .A(n12981), .ZN(n13000) );
  INV_X1 U15139 ( .A(n12982), .ZN(n12999) );
  OR2_X1 U15140 ( .A1(n12985), .A2(n12984), .ZN(n12988) );
  NAND2_X1 U15141 ( .A1(n13006), .A2(n12986), .ZN(n12987) );
  NAND2_X1 U15142 ( .A1(n12988), .A2(n12987), .ZN(n13122) );
  OAI22_X1 U15143 ( .A1(n13126), .A2(n12990), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12989), .ZN(n12991) );
  AOI21_X1 U15144 ( .B1(n13122), .B2(n12992), .A(n12991), .ZN(n12993) );
  OAI21_X1 U15145 ( .B1(n13129), .B2(n12994), .A(n12993), .ZN(n12995) );
  AOI21_X1 U15146 ( .B1(n12997), .B2(n12996), .A(n12995), .ZN(n12998) );
  OAI21_X1 U15147 ( .B1(n13000), .B2(n12999), .A(n12998), .ZN(P2_U3212) );
  MUX2_X1 U15148 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13079), .S(n6427), .Z(
        P2_U3562) );
  MUX2_X1 U15149 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13001), .S(n6427), .Z(
        P2_U3561) );
  MUX2_X1 U15150 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13002), .S(n6427), .Z(
        P2_U3560) );
  MUX2_X1 U15151 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13003), .S(P2_U3947), .Z(
        P2_U3559) );
  MUX2_X1 U15152 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13004), .S(P2_U3947), .Z(
        P2_U3558) );
  MUX2_X1 U15153 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13005), .S(P2_U3947), .Z(
        P2_U3557) );
  MUX2_X1 U15154 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13006), .S(P2_U3947), .Z(
        P2_U3556) );
  MUX2_X1 U15155 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13007), .S(P2_U3947), .Z(
        P2_U3555) );
  MUX2_X1 U15156 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13008), .S(P2_U3947), .Z(
        P2_U3554) );
  MUX2_X1 U15157 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13009), .S(n6427), .Z(
        P2_U3553) );
  MUX2_X1 U15158 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13010), .S(n6427), .Z(
        P2_U3552) );
  MUX2_X1 U15159 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13011), .S(n6427), .Z(
        P2_U3551) );
  MUX2_X1 U15160 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13012), .S(n6427), .Z(
        P2_U3550) );
  MUX2_X1 U15161 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13013), .S(n6427), .Z(
        P2_U3549) );
  MUX2_X1 U15162 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13014), .S(n6427), .Z(
        P2_U3548) );
  MUX2_X1 U15163 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13015), .S(n6427), .Z(
        P2_U3547) );
  MUX2_X1 U15164 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13016), .S(n6427), .Z(
        P2_U3546) );
  MUX2_X1 U15165 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13017), .S(n6427), .Z(
        P2_U3545) );
  MUX2_X1 U15166 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n13018), .S(n6427), .Z(
        P2_U3544) );
  MUX2_X1 U15167 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13019), .S(n6427), .Z(
        P2_U3543) );
  MUX2_X1 U15168 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13020), .S(n6427), .Z(
        P2_U3542) );
  MUX2_X1 U15169 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13021), .S(n6427), .Z(
        P2_U3541) );
  MUX2_X1 U15170 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13022), .S(n6427), .Z(
        P2_U3540) );
  MUX2_X1 U15171 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13023), .S(n6427), .Z(
        P2_U3539) );
  MUX2_X1 U15172 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13024), .S(n6427), .Z(
        P2_U3538) );
  MUX2_X1 U15173 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13025), .S(n6427), .Z(
        P2_U3537) );
  MUX2_X1 U15174 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13026), .S(n6427), .Z(
        P2_U3536) );
  MUX2_X1 U15175 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13027), .S(n6427), .Z(
        P2_U3535) );
  MUX2_X1 U15176 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13028), .S(n6427), .Z(
        P2_U3534) );
  MUX2_X1 U15177 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n13029), .S(n6427), .Z(
        P2_U3533) );
  MUX2_X1 U15178 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n6429), .S(n6427), .Z(
        P2_U3532) );
  MUX2_X1 U15179 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n13030), .S(n6427), .Z(
        P2_U3531) );
  AND3_X1 U15180 ( .A1(n14764), .A2(n13032), .A3(n13031), .ZN(n13033) );
  NOR3_X1 U15181 ( .A1(n14838), .A2(n13034), .A3(n13033), .ZN(n13035) );
  AOI21_X1 U15182 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(n14818), .A(n13035), .ZN(
        n13044) );
  NAND2_X1 U15183 ( .A1(n14841), .A2(n13036), .ZN(n13042) );
  MUX2_X1 U15184 ( .A(n10177), .B(P2_REG1_REG_5__SCAN_IN), .S(n13036), .Z(
        n13037) );
  NAND3_X1 U15185 ( .A1(n14767), .A2(n13038), .A3(n13037), .ZN(n13039) );
  NAND3_X1 U15186 ( .A1(n14825), .A2(n13040), .A3(n13039), .ZN(n13041) );
  NAND4_X1 U15187 ( .A1(n13044), .A2(n13043), .A3(n13042), .A4(n13041), .ZN(
        P2_U3219) );
  OAI21_X1 U15188 ( .B1(n14845), .B2(n7057), .A(n13045), .ZN(n13046) );
  AOI21_X1 U15189 ( .B1(n13052), .B2(n14841), .A(n13046), .ZN(n13059) );
  MUX2_X1 U15190 ( .A(n10169), .B(P2_REG2_REG_7__SCAN_IN), .S(n13052), .Z(
        n13049) );
  INV_X1 U15191 ( .A(n13047), .ZN(n13048) );
  NAND2_X1 U15192 ( .A1(n13049), .A2(n13048), .ZN(n13051) );
  OAI211_X1 U15193 ( .C1(n14780), .C2(n13051), .A(n13050), .B(n14820), .ZN(
        n13058) );
  MUX2_X1 U15194 ( .A(n10183), .B(P2_REG1_REG_7__SCAN_IN), .S(n13052), .Z(
        n13053) );
  NAND3_X1 U15195 ( .A1(n14777), .A2(n13054), .A3(n13053), .ZN(n13055) );
  NAND3_X1 U15196 ( .A1(n14825), .A2(n13056), .A3(n13055), .ZN(n13057) );
  NAND3_X1 U15197 ( .A1(n13059), .A2(n13058), .A3(n13057), .ZN(P2_U3221) );
  OAI21_X1 U15198 ( .B1(n13062), .B2(n13061), .A(n13060), .ZN(n13063) );
  NAND2_X1 U15199 ( .A1(n13063), .A2(n14820), .ZN(n13076) );
  INV_X1 U15200 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14365) );
  OAI21_X1 U15201 ( .B1(n14845), .B2(n14365), .A(n13064), .ZN(n13065) );
  AOI21_X1 U15202 ( .B1(n13066), .B2(n14841), .A(n13065), .ZN(n13075) );
  MUX2_X1 U15203 ( .A(n13067), .B(P2_REG1_REG_11__SCAN_IN), .S(n13066), .Z(
        n13070) );
  INV_X1 U15204 ( .A(n13068), .ZN(n13069) );
  NAND2_X1 U15205 ( .A1(n13070), .A2(n13069), .ZN(n13072) );
  OAI211_X1 U15206 ( .C1(n13073), .C2(n13072), .A(n13071), .B(n14825), .ZN(
        n13074) );
  NAND3_X1 U15207 ( .A1(n13076), .A2(n13075), .A3(n13074), .ZN(P2_U3225) );
  NAND2_X1 U15208 ( .A1(n13082), .A2(n13086), .ZN(n13085) );
  XNOR2_X1 U15209 ( .A(n13378), .B(n13085), .ZN(n13077) );
  NOR2_X1 U15210 ( .A1(n14868), .A2(n14205), .ZN(n13080) );
  NAND2_X1 U15211 ( .A1(n13079), .A2(n13078), .ZN(n13295) );
  NOR2_X1 U15212 ( .A1(n14478), .A2(n13295), .ZN(n13088) );
  AOI211_X1 U15213 ( .C1(n13378), .C2(n14479), .A(n13080), .B(n13088), .ZN(
        n13081) );
  OAI21_X1 U15214 ( .B1(n13292), .B2(n13221), .A(n13081), .ZN(P2_U3234) );
  OR2_X1 U15215 ( .A1(n13082), .A2(n13086), .ZN(n13084) );
  NAND3_X1 U15216 ( .A1(n13085), .A2(n13084), .A3(n13083), .ZN(n13296) );
  NOR2_X1 U15217 ( .A1(n13086), .A2(n14853), .ZN(n13087) );
  AOI211_X1 U15218 ( .C1(n14478), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13088), 
        .B(n13087), .ZN(n13089) );
  OAI21_X1 U15219 ( .B1(n13221), .B2(n13296), .A(n13089), .ZN(P2_U3235) );
  NAND2_X1 U15220 ( .A1(n13092), .A2(n14475), .ZN(n13098) );
  AOI21_X1 U15221 ( .B1(n13108), .B2(n13094), .A(n13093), .ZN(n13097) );
  INV_X1 U15222 ( .A(n13095), .ZN(n13096) );
  OAI21_X1 U15223 ( .B1(n13098), .B2(n13097), .A(n13096), .ZN(n13304) );
  NOR2_X1 U15224 ( .A1(n13099), .A2(n14863), .ZN(n13100) );
  OAI21_X1 U15225 ( .B1(n13304), .B2(n13100), .A(n14868), .ZN(n13106) );
  NOR2_X1 U15226 ( .A1(n13306), .A2(n13114), .ZN(n13101) );
  NOR3_X1 U15227 ( .A1(n13102), .A2(n13101), .A3(n7799), .ZN(n13307) );
  OAI22_X1 U15228 ( .A1(n13306), .A2(n14853), .B1(n14868), .B2(n13103), .ZN(
        n13104) );
  AOI21_X1 U15229 ( .B1(n13307), .B2(n14847), .A(n13104), .ZN(n13105) );
  OAI211_X1 U15230 ( .C1(n13254), .C2(n13303), .A(n13106), .B(n13105), .ZN(
        P2_U3237) );
  XNOR2_X1 U15231 ( .A(n13107), .B(n13109), .ZN(n13314) );
  OAI21_X1 U15232 ( .B1(n13110), .B2(n13109), .A(n13108), .ZN(n13112) );
  AOI21_X1 U15233 ( .B1(n13112), .B2(n14475), .A(n13111), .ZN(n13313) );
  NOR2_X1 U15234 ( .A1(n13389), .A2(n13124), .ZN(n13113) );
  AOI22_X1 U15235 ( .A1(n13115), .A2(n14849), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n14478), .ZN(n13118) );
  NAND2_X1 U15236 ( .A1(n13116), .A2(n14479), .ZN(n13117) );
  OAI211_X1 U15237 ( .C1(n13312), .C2(n13221), .A(n13118), .B(n13117), .ZN(
        n13119) );
  AOI21_X1 U15238 ( .B1(n6609), .B2(n14868), .A(n13119), .ZN(n13120) );
  OAI21_X1 U15239 ( .B1(n13314), .B2(n13254), .A(n13120), .ZN(P2_U3238) );
  XOR2_X1 U15240 ( .A(n13131), .B(n13121), .Z(n13123) );
  AOI21_X1 U15241 ( .B1(n13123), .B2(n14475), .A(n13122), .ZN(n13320) );
  INV_X1 U15242 ( .A(n13142), .ZN(n13125) );
  AOI211_X1 U15243 ( .C1(n13318), .C2(n13125), .A(n7779), .B(n13124), .ZN(
        n13317) );
  INV_X1 U15244 ( .A(n13126), .ZN(n13127) );
  AOI22_X1 U15245 ( .A1(n13127), .A2(n14849), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n14478), .ZN(n13128) );
  OAI21_X1 U15246 ( .B1(n13129), .B2(n14853), .A(n13128), .ZN(n13133) );
  XNOR2_X1 U15247 ( .A(n13131), .B(n13130), .ZN(n13321) );
  NOR2_X1 U15248 ( .A1(n13321), .A2(n13254), .ZN(n13132) );
  AOI211_X1 U15249 ( .C1(n13317), .C2(n14847), .A(n13133), .B(n13132), .ZN(
        n13134) );
  OAI21_X1 U15250 ( .B1(n14478), .B2(n13320), .A(n13134), .ZN(P2_U3239) );
  XNOR2_X1 U15251 ( .A(n13135), .B(n13136), .ZN(n13323) );
  INV_X1 U15252 ( .A(n13323), .ZN(n13148) );
  XNOR2_X1 U15253 ( .A(n13138), .B(n13137), .ZN(n13140) );
  OAI21_X1 U15254 ( .B1(n13140), .B2(n13279), .A(n13139), .ZN(n13322) );
  NAND2_X1 U15255 ( .A1(n13322), .A2(n14868), .ZN(n13147) );
  OAI21_X1 U15256 ( .B1(n13394), .B2(n13158), .A(n13083), .ZN(n13141) );
  AOI22_X1 U15257 ( .A1(P2_REG2_REG_25__SCAN_IN), .A2(n14478), .B1(n13143), 
        .B2(n14849), .ZN(n13144) );
  OAI21_X1 U15258 ( .B1(n13394), .B2(n14853), .A(n13144), .ZN(n13145) );
  AOI21_X1 U15259 ( .B1(n6466), .B2(n14847), .A(n13145), .ZN(n13146) );
  OAI211_X1 U15260 ( .C1(n13148), .C2(n13254), .A(n13147), .B(n13146), .ZN(
        P2_U3240) );
  XNOR2_X1 U15261 ( .A(n13150), .B(n13149), .ZN(n13151) );
  INV_X1 U15262 ( .A(n13152), .ZN(n13153) );
  XNOR2_X1 U15263 ( .A(n13156), .B(n13155), .ZN(n13328) );
  OAI21_X1 U15264 ( .B1(n13398), .B2(n13169), .A(n13083), .ZN(n13157) );
  OR2_X1 U15265 ( .A1(n13158), .A2(n13157), .ZN(n13326) );
  INV_X1 U15266 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13160) );
  OAI22_X1 U15267 ( .A1(n14868), .A2(n13160), .B1(n13159), .B2(n14863), .ZN(
        n13161) );
  AOI21_X1 U15268 ( .B1(n13162), .B2(n14479), .A(n13161), .ZN(n13163) );
  OAI21_X1 U15269 ( .B1(n13326), .B2(n13221), .A(n13163), .ZN(n13164) );
  AOI21_X1 U15270 ( .B1(n13328), .B2(n14856), .A(n13164), .ZN(n13165) );
  OAI21_X1 U15271 ( .B1(n13329), .B2(n14478), .A(n13165), .ZN(P2_U3241) );
  XNOR2_X1 U15272 ( .A(n13166), .B(n13176), .ZN(n13168) );
  AOI21_X1 U15273 ( .B1(n13168), .B2(n14475), .A(n13167), .ZN(n13334) );
  INV_X1 U15274 ( .A(n13189), .ZN(n13170) );
  AOI211_X1 U15275 ( .C1(n6769), .C2(n13170), .A(n7779), .B(n13169), .ZN(
        n13333) );
  INV_X1 U15276 ( .A(n13171), .ZN(n13172) );
  AOI22_X1 U15277 ( .A1(n14478), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n13172), 
        .B2(n14849), .ZN(n13173) );
  OAI21_X1 U15278 ( .B1(n13174), .B2(n14853), .A(n13173), .ZN(n13178) );
  XOR2_X1 U15279 ( .A(n13175), .B(n13176), .Z(n13336) );
  NOR2_X1 U15280 ( .A1(n13336), .A2(n13254), .ZN(n13177) );
  AOI211_X1 U15281 ( .C1(n13333), .C2(n14847), .A(n13178), .B(n13177), .ZN(
        n13179) );
  OAI21_X1 U15282 ( .B1(n14478), .B2(n13334), .A(n13179), .ZN(P2_U3242) );
  XNOR2_X1 U15283 ( .A(n13180), .B(n13181), .ZN(n13183) );
  AOI21_X1 U15284 ( .B1(n13183), .B2(n14475), .A(n13182), .ZN(n13338) );
  NAND2_X1 U15285 ( .A1(n13185), .A2(n13184), .ZN(n13186) );
  NAND2_X1 U15286 ( .A1(n13187), .A2(n13186), .ZN(n13339) );
  INV_X1 U15287 ( .A(n13339), .ZN(n13195) );
  NOR2_X1 U15288 ( .A1(n13192), .A2(n13198), .ZN(n13188) );
  OR3_X1 U15289 ( .A1(n13189), .A2(n13188), .A3(n7799), .ZN(n13337) );
  NOR2_X1 U15290 ( .A1(n13337), .A2(n13221), .ZN(n13194) );
  AOI22_X1 U15291 ( .A1(n14478), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n13190), 
        .B2(n14849), .ZN(n13191) );
  OAI21_X1 U15292 ( .B1(n13192), .B2(n14853), .A(n13191), .ZN(n13193) );
  AOI211_X1 U15293 ( .C1(n13195), .C2(n14856), .A(n13194), .B(n13193), .ZN(
        n13196) );
  OAI21_X1 U15294 ( .B1(n14478), .B2(n13338), .A(n13196), .ZN(P2_U3243) );
  XOR2_X1 U15295 ( .A(n13197), .B(n13203), .Z(n13346) );
  AOI211_X1 U15296 ( .C1(n13344), .C2(n13215), .A(n7779), .B(n13198), .ZN(
        n13343) );
  NOR2_X1 U15297 ( .A1(n6767), .A2(n14853), .ZN(n13202) );
  INV_X1 U15298 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n13200) );
  OAI22_X1 U15299 ( .A1(n14868), .A2(n13200), .B1(n13199), .B2(n14863), .ZN(
        n13201) );
  AOI211_X1 U15300 ( .C1(n13343), .C2(n14847), .A(n13202), .B(n13201), .ZN(
        n13208) );
  XNOR2_X1 U15301 ( .A(n13204), .B(n13203), .ZN(n13206) );
  OAI21_X1 U15302 ( .B1(n13206), .B2(n13279), .A(n13205), .ZN(n13342) );
  NAND2_X1 U15303 ( .A1(n13342), .A2(n14868), .ZN(n13207) );
  OAI211_X1 U15304 ( .C1(n13346), .C2(n13254), .A(n13208), .B(n13207), .ZN(
        P2_U3244) );
  XNOR2_X1 U15305 ( .A(n13210), .B(n13209), .ZN(n13349) );
  OAI21_X1 U15306 ( .B1(n6525), .B2(n13212), .A(n13211), .ZN(n13214) );
  AOI21_X1 U15307 ( .B1(n13214), .B2(n14475), .A(n13213), .ZN(n13348) );
  INV_X1 U15308 ( .A(n13348), .ZN(n13223) );
  AOI21_X1 U15309 ( .B1(n13406), .B2(n13228), .A(n7799), .ZN(n13216) );
  NAND2_X1 U15310 ( .A1(n13216), .A2(n13215), .ZN(n13347) );
  INV_X1 U15311 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n13218) );
  OAI22_X1 U15312 ( .A1(n14868), .A2(n13218), .B1(n13217), .B2(n14863), .ZN(
        n13219) );
  AOI21_X1 U15313 ( .B1(n13406), .B2(n14479), .A(n13219), .ZN(n13220) );
  OAI21_X1 U15314 ( .B1(n13347), .B2(n13221), .A(n13220), .ZN(n13222) );
  AOI21_X1 U15315 ( .B1(n13223), .B2(n14868), .A(n13222), .ZN(n13224) );
  OAI21_X1 U15316 ( .B1(n13349), .B2(n13254), .A(n13224), .ZN(P2_U3245) );
  XNOR2_X1 U15317 ( .A(n13226), .B(n13225), .ZN(n13355) );
  INV_X1 U15318 ( .A(n13355), .ZN(n13241) );
  AOI211_X1 U15319 ( .C1(n13229), .C2(n13246), .A(n7779), .B(n6761), .ZN(
        n13354) );
  NOR2_X1 U15320 ( .A1(n10020), .A2(n14853), .ZN(n13233) );
  OAI22_X1 U15321 ( .A1(n14868), .A2(n13231), .B1(n13230), .B2(n14863), .ZN(
        n13232) );
  AOI211_X1 U15322 ( .C1(n13354), .C2(n14847), .A(n13233), .B(n13232), .ZN(
        n13240) );
  OAI211_X1 U15323 ( .C1(n13236), .C2(n13235), .A(n14475), .B(n6593), .ZN(
        n13238) );
  NAND2_X1 U15324 ( .A1(n13238), .A2(n13237), .ZN(n13353) );
  NAND2_X1 U15325 ( .A1(n13353), .A2(n14868), .ZN(n13239) );
  OAI211_X1 U15326 ( .C1(n13241), .C2(n13254), .A(n13240), .B(n13239), .ZN(
        P2_U3246) );
  XNOR2_X1 U15327 ( .A(n13243), .B(n13251), .ZN(n13245) );
  AOI21_X1 U15328 ( .B1(n13245), .B2(n14475), .A(n13244), .ZN(n13361) );
  AOI211_X1 U15329 ( .C1(n13359), .C2(n6558), .A(n7779), .B(n13227), .ZN(
        n13358) );
  INV_X1 U15330 ( .A(n13247), .ZN(n13248) );
  AOI22_X1 U15331 ( .A1(n14478), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13248), 
        .B2(n14849), .ZN(n13249) );
  OAI21_X1 U15332 ( .B1(n6763), .B2(n14853), .A(n13249), .ZN(n13256) );
  OAI21_X1 U15333 ( .B1(n13252), .B2(n13251), .A(n13250), .ZN(n13253) );
  INV_X1 U15334 ( .A(n13253), .ZN(n13363) );
  NOR2_X1 U15335 ( .A1(n13363), .A2(n13254), .ZN(n13255) );
  AOI211_X1 U15336 ( .C1(n13358), .C2(n14847), .A(n13256), .B(n13255), .ZN(
        n13257) );
  OAI21_X1 U15337 ( .B1(n14478), .B2(n13361), .A(n13257), .ZN(P2_U3247) );
  XNOR2_X1 U15338 ( .A(n13259), .B(n13258), .ZN(n13261) );
  OAI21_X1 U15339 ( .B1(n13261), .B2(n13279), .A(n13260), .ZN(n13364) );
  NAND2_X1 U15340 ( .A1(n13364), .A2(n14868), .ZN(n13273) );
  OAI22_X1 U15341 ( .A1(n14868), .A2(n13263), .B1(n13262), .B2(n14863), .ZN(
        n13264) );
  AOI21_X1 U15342 ( .B1(n13265), .B2(n14479), .A(n13264), .ZN(n13272) );
  XNOR2_X1 U15343 ( .A(n13267), .B(n13266), .ZN(n13366) );
  NAND2_X1 U15344 ( .A1(n13366), .A2(n14856), .ZN(n13271) );
  OR2_X1 U15345 ( .A1(n13416), .A2(n13268), .ZN(n13269) );
  AND3_X1 U15346 ( .A1(n6558), .A2(n13269), .A3(n13083), .ZN(n13365) );
  NAND2_X1 U15347 ( .A1(n13365), .A2(n14847), .ZN(n13270) );
  NAND4_X1 U15348 ( .A1(n13273), .A2(n13272), .A3(n13271), .A4(n13270), .ZN(
        P2_U3248) );
  INV_X1 U15349 ( .A(n13274), .ZN(n13275) );
  AOI21_X1 U15350 ( .B1(n13277), .B2(n13276), .A(n13275), .ZN(n13280) );
  OAI21_X1 U15351 ( .B1(n13280), .B2(n13279), .A(n13278), .ZN(n13369) );
  NAND2_X1 U15352 ( .A1(n13369), .A2(n14868), .ZN(n13291) );
  OAI22_X1 U15353 ( .A1(n14868), .A2(n11407), .B1(n13281), .B2(n14863), .ZN(
        n13282) );
  AOI21_X1 U15354 ( .B1(n13285), .B2(n14479), .A(n13282), .ZN(n13290) );
  AOI21_X1 U15355 ( .B1(n9989), .B2(n13283), .A(n6555), .ZN(n13371) );
  NAND2_X1 U15356 ( .A1(n13371), .A2(n14856), .ZN(n13289) );
  AOI21_X1 U15357 ( .B1(n13285), .B2(n13284), .A(n7799), .ZN(n13287) );
  AND2_X1 U15358 ( .A1(n13287), .A2(n13286), .ZN(n13370) );
  NAND2_X1 U15359 ( .A1(n13370), .A2(n14847), .ZN(n13288) );
  NAND4_X1 U15360 ( .A1(n13291), .A2(n13290), .A3(n13289), .A4(n13288), .ZN(
        P2_U3249) );
  NAND2_X1 U15361 ( .A1(n13292), .A2(n13295), .ZN(n13376) );
  MUX2_X1 U15362 ( .A(n13376), .B(P2_REG1_REG_31__SCAN_IN), .S(n14900), .Z(
        n13293) );
  AOI21_X1 U15363 ( .B1(n13351), .B2(n13378), .A(n13293), .ZN(n13294) );
  INV_X1 U15364 ( .A(n13294), .ZN(P2_U3530) );
  NAND2_X1 U15365 ( .A1(n13296), .A2(n13295), .ZN(n13380) );
  MUX2_X1 U15366 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13380), .S(n14903), .Z(
        n13297) );
  AOI21_X1 U15367 ( .B1(n13351), .B2(n13382), .A(n13297), .ZN(n13298) );
  INV_X1 U15368 ( .A(n13298), .ZN(P2_U3529) );
  AOI21_X1 U15369 ( .B1(n14490), .B2(n8282), .A(n13299), .ZN(n13300) );
  OAI211_X1 U15370 ( .C1(n13302), .C2(n13362), .A(n13301), .B(n13300), .ZN(
        n13384) );
  MUX2_X1 U15371 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13384), .S(n14903), .Z(
        P2_U3528) );
  INV_X1 U15372 ( .A(n13304), .ZN(n13310) );
  INV_X1 U15373 ( .A(n14490), .ZN(n13305) );
  NOR2_X1 U15374 ( .A1(n13308), .A2(n13307), .ZN(n13309) );
  NAND3_X1 U15375 ( .A1(n13311), .A2(n13310), .A3(n13309), .ZN(n13385) );
  MUX2_X1 U15376 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13385), .S(n14903), .Z(
        P2_U3527) );
  MUX2_X1 U15377 ( .A(n13315), .B(n13386), .S(n14903), .Z(n13316) );
  AOI21_X1 U15378 ( .B1(n14490), .B2(n13318), .A(n13317), .ZN(n13319) );
  OAI211_X1 U15379 ( .C1(n13362), .C2(n13321), .A(n13320), .B(n13319), .ZN(
        n13390) );
  MUX2_X1 U15380 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13390), .S(n14903), .Z(
        P2_U3525) );
  AOI211_X1 U15381 ( .C1(n14511), .C2(n13323), .A(n6466), .B(n13322), .ZN(
        n13391) );
  MUX2_X1 U15382 ( .A(n13324), .B(n13391), .S(n14903), .Z(n13325) );
  OAI21_X1 U15383 ( .B1(n13394), .B2(n13374), .A(n13325), .ZN(P2_U3524) );
  INV_X1 U15384 ( .A(n13326), .ZN(n13327) );
  AOI21_X1 U15385 ( .B1(n13328), .B2(n14511), .A(n13327), .ZN(n13330) );
  MUX2_X1 U15386 ( .A(n13396), .B(n13331), .S(n14900), .Z(n13332) );
  OAI21_X1 U15387 ( .B1(n13398), .B2(n13374), .A(n13332), .ZN(P2_U3523) );
  AOI21_X1 U15388 ( .B1(n14490), .B2(n6769), .A(n13333), .ZN(n13335) );
  OAI211_X1 U15389 ( .C1(n13362), .C2(n13336), .A(n13335), .B(n13334), .ZN(
        n13399) );
  MUX2_X1 U15390 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13399), .S(n14903), .Z(
        P2_U3522) );
  OAI211_X1 U15391 ( .C1(n13339), .C2(n13362), .A(n13338), .B(n13337), .ZN(
        n13400) );
  MUX2_X1 U15392 ( .A(n13400), .B(P2_REG1_REG_22__SCAN_IN), .S(n14900), .Z(
        n13340) );
  AOI21_X1 U15393 ( .B1(n13351), .B2(n6770), .A(n13340), .ZN(n13341) );
  INV_X1 U15394 ( .A(n13341), .ZN(P2_U3521) );
  AOI211_X1 U15395 ( .C1(n14490), .C2(n13344), .A(n13343), .B(n13342), .ZN(
        n13345) );
  OAI21_X1 U15396 ( .B1(n13362), .B2(n13346), .A(n13345), .ZN(n13403) );
  MUX2_X1 U15397 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13403), .S(n14903), .Z(
        P2_U3520) );
  OAI211_X1 U15398 ( .C1(n13349), .C2(n13362), .A(n13348), .B(n13347), .ZN(
        n13404) );
  MUX2_X1 U15399 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13404), .S(n14903), .Z(
        n13350) );
  AOI21_X1 U15400 ( .B1(n13351), .B2(n13406), .A(n13350), .ZN(n13352) );
  INV_X1 U15401 ( .A(n13352), .ZN(P2_U3519) );
  INV_X1 U15402 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13356) );
  AOI211_X1 U15403 ( .C1(n13355), .C2(n14511), .A(n13354), .B(n13353), .ZN(
        n13409) );
  MUX2_X1 U15404 ( .A(n13356), .B(n13409), .S(n14903), .Z(n13357) );
  OAI21_X1 U15405 ( .B1(n10020), .B2(n13374), .A(n13357), .ZN(P2_U3518) );
  AOI21_X1 U15406 ( .B1(n14490), .B2(n13359), .A(n13358), .ZN(n13360) );
  OAI211_X1 U15407 ( .C1(n13363), .C2(n13362), .A(n13361), .B(n13360), .ZN(
        n13412) );
  MUX2_X1 U15408 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13412), .S(n14903), .Z(
        P2_U3517) );
  AOI211_X1 U15409 ( .C1(n14511), .C2(n13366), .A(n13365), .B(n13364), .ZN(
        n13413) );
  MUX2_X1 U15410 ( .A(n13367), .B(n13413), .S(n14903), .Z(n13368) );
  OAI21_X1 U15411 ( .B1(n13416), .B2(n13374), .A(n13368), .ZN(P2_U3516) );
  AOI211_X1 U15412 ( .C1(n13371), .C2(n14511), .A(n13370), .B(n13369), .ZN(
        n13417) );
  MUX2_X1 U15413 ( .A(n13372), .B(n13417), .S(n14903), .Z(n13373) );
  OAI21_X1 U15414 ( .B1(n13421), .B2(n13374), .A(n13373), .ZN(P2_U3515) );
  MUX2_X1 U15415 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n13375), .S(n14903), .Z(
        P2_U3499) );
  MUX2_X1 U15416 ( .A(n13376), .B(P2_REG0_REG_31__SCAN_IN), .S(n14896), .Z(
        n13377) );
  AOI21_X1 U15417 ( .B1(n13407), .B2(n13378), .A(n13377), .ZN(n13379) );
  INV_X1 U15418 ( .A(n13379), .ZN(P2_U3498) );
  MUX2_X1 U15419 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13380), .S(n14898), .Z(
        n13381) );
  AOI21_X1 U15420 ( .B1(n13407), .B2(n13382), .A(n13381), .ZN(n13383) );
  INV_X1 U15421 ( .A(n13383), .ZN(P2_U3497) );
  MUX2_X1 U15422 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13384), .S(n14898), .Z(
        P2_U3496) );
  MUX2_X1 U15423 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13385), .S(n14898), .Z(
        P2_U3495) );
  INV_X1 U15424 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n13387) );
  MUX2_X1 U15425 ( .A(n13387), .B(n13386), .S(n14898), .Z(n13388) );
  MUX2_X1 U15426 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13390), .S(n14898), .Z(
        P2_U3493) );
  INV_X1 U15427 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n13392) );
  MUX2_X1 U15428 ( .A(n13392), .B(n13391), .S(n14898), .Z(n13393) );
  OAI21_X1 U15429 ( .B1(n13394), .B2(n13420), .A(n13393), .ZN(P2_U3492) );
  INV_X1 U15430 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n13395) );
  MUX2_X1 U15431 ( .A(n13396), .B(n13395), .S(n14896), .Z(n13397) );
  OAI21_X1 U15432 ( .B1(n13398), .B2(n13420), .A(n13397), .ZN(P2_U3491) );
  MUX2_X1 U15433 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13399), .S(n14898), .Z(
        P2_U3490) );
  MUX2_X1 U15434 ( .A(n13400), .B(P2_REG0_REG_22__SCAN_IN), .S(n14896), .Z(
        n13401) );
  AOI21_X1 U15435 ( .B1(n13407), .B2(n6770), .A(n13401), .ZN(n13402) );
  INV_X1 U15436 ( .A(n13402), .ZN(P2_U3489) );
  MUX2_X1 U15437 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13403), .S(n14898), .Z(
        P2_U3488) );
  MUX2_X1 U15438 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13404), .S(n14898), .Z(
        n13405) );
  AOI21_X1 U15439 ( .B1(n13407), .B2(n13406), .A(n13405), .ZN(n13408) );
  INV_X1 U15440 ( .A(n13408), .ZN(P2_U3487) );
  INV_X1 U15441 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n13410) );
  MUX2_X1 U15442 ( .A(n13410), .B(n13409), .S(n14898), .Z(n13411) );
  OAI21_X1 U15443 ( .B1(n10020), .B2(n13420), .A(n13411), .ZN(P2_U3486) );
  MUX2_X1 U15444 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13412), .S(n14898), .Z(
        P2_U3484) );
  INV_X1 U15445 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n13414) );
  MUX2_X1 U15446 ( .A(n13414), .B(n13413), .S(n14898), .Z(n13415) );
  OAI21_X1 U15447 ( .B1(n13416), .B2(n13420), .A(n13415), .ZN(P2_U3481) );
  INV_X1 U15448 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n13418) );
  MUX2_X1 U15449 ( .A(n13418), .B(n13417), .S(n14898), .Z(n13419) );
  OAI21_X1 U15450 ( .B1(n13421), .B2(n13420), .A(n13419), .ZN(P2_U3478) );
  INV_X1 U15451 ( .A(n14268), .ZN(n13425) );
  NOR4_X1 U15452 ( .A1(n13422), .A2(P2_IR_REG_30__SCAN_IN), .A3(n7677), .A4(
        P2_U3088), .ZN(n13423) );
  AOI21_X1 U15453 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n13433), .A(n13423), 
        .ZN(n13424) );
  OAI21_X1 U15454 ( .B1(n13425), .B2(n13438), .A(n13424), .ZN(P2_U3296) );
  OAI222_X1 U15455 ( .A1(n13438), .A2(n13428), .B1(n13427), .B2(P2_U3088), 
        .C1(n13426), .C2(n13440), .ZN(P2_U3298) );
  AOI21_X1 U15456 ( .B1(n13433), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13429), 
        .ZN(n13430) );
  OAI21_X1 U15457 ( .B1(n13431), .B2(n13438), .A(n13430), .ZN(P2_U3299) );
  INV_X1 U15458 ( .A(n13432), .ZN(n14276) );
  AOI22_X1 U15459 ( .A1(n13434), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n13433), .ZN(n13435) );
  OAI21_X1 U15460 ( .B1(n14276), .B2(n13438), .A(n13435), .ZN(P2_U3301) );
  INV_X1 U15461 ( .A(n13436), .ZN(n14280) );
  OAI222_X1 U15462 ( .A1(n13440), .A2(n13439), .B1(n13438), .B2(n14280), .C1(
        P2_U3088), .C2(n13437), .ZN(P2_U3302) );
  INV_X1 U15463 ( .A(n13441), .ZN(n13442) );
  MUX2_X1 U15464 ( .A(n13442), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  INV_X1 U15465 ( .A(n14034), .ZN(n13804) );
  NAND2_X1 U15466 ( .A1(n13445), .A2(n13537), .ZN(n13450) );
  INV_X1 U15467 ( .A(n13446), .ZN(n13801) );
  AOI22_X1 U15468 ( .A1(n13981), .A2(n13749), .B1(n13765), .B2(n13983), .ZN(
        n13793) );
  OAI22_X1 U15469 ( .A1(n13540), .A2(n13793), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13447), .ZN(n13448) );
  AOI21_X1 U15470 ( .B1(n13543), .B2(n13801), .A(n13448), .ZN(n13449) );
  OAI211_X1 U15471 ( .C1(n13804), .C2(n13526), .A(n13450), .B(n13449), .ZN(
        P1_U3214) );
  INV_X1 U15472 ( .A(n13451), .ZN(n13455) );
  OAI21_X1 U15473 ( .B1(n6465), .B2(n13453), .A(n13452), .ZN(n13454) );
  NAND3_X1 U15474 ( .A1(n13455), .A2(n13537), .A3(n13454), .ZN(n13460) );
  OR2_X1 U15475 ( .A1(n13743), .A2(n13993), .ZN(n13457) );
  OR2_X1 U15476 ( .A1(n13955), .A2(n13991), .ZN(n13456) );
  NAND2_X1 U15477 ( .A1(n13457), .A2(n13456), .ZN(n14220) );
  AND2_X1 U15478 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13693) );
  NOR2_X1 U15479 ( .A1(n13553), .A2(n13923), .ZN(n13458) );
  AOI211_X1 U15480 ( .C1(n13475), .C2(n14220), .A(n13693), .B(n13458), .ZN(
        n13459) );
  OAI211_X1 U15481 ( .C1(n6826), .C2(n13526), .A(n13460), .B(n13459), .ZN(
        P1_U3219) );
  AOI21_X1 U15482 ( .B1(n13463), .B2(n13462), .A(n13461), .ZN(n13469) );
  NAND2_X1 U15483 ( .A1(n13745), .A2(n13983), .ZN(n13465) );
  OR2_X1 U15484 ( .A1(n13743), .A2(n13991), .ZN(n13464) );
  NAND2_X1 U15485 ( .A1(n13465), .A2(n13464), .ZN(n14072) );
  AOI22_X1 U15486 ( .A1(n14072), .A2(n13475), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13466) );
  OAI21_X1 U15487 ( .B1(n13553), .B2(n13890), .A(n13466), .ZN(n13467) );
  AOI21_X1 U15488 ( .B1(n14073), .B2(n13555), .A(n13467), .ZN(n13468) );
  OAI21_X1 U15489 ( .B1(n13469), .B2(n13557), .A(n13468), .ZN(P1_U3223) );
  OAI21_X1 U15490 ( .B1(n13472), .B2(n13470), .A(n13471), .ZN(n13479) );
  NAND2_X1 U15491 ( .A1(n14045), .A2(n13555), .ZN(n13477) );
  NAND2_X1 U15492 ( .A1(n13725), .A2(n13981), .ZN(n13474) );
  NAND2_X1 U15493 ( .A1(n13749), .A2(n13983), .ZN(n13473) );
  NAND2_X1 U15494 ( .A1(n13474), .A2(n13473), .ZN(n14044) );
  AOI22_X1 U15495 ( .A1(n13475), .A2(n14044), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13476) );
  OAI211_X1 U15496 ( .C1(n13553), .C2(n13827), .A(n13477), .B(n13476), .ZN(
        n13478) );
  AOI21_X1 U15497 ( .B1(n13479), .B2(n13537), .A(n13478), .ZN(n13480) );
  INV_X1 U15498 ( .A(n13480), .ZN(P1_U3225) );
  OAI21_X1 U15499 ( .B1(n13483), .B2(n13482), .A(n13481), .ZN(n13484) );
  NAND2_X1 U15500 ( .A1(n13484), .A2(n13537), .ZN(n13489) );
  NAND2_X1 U15501 ( .A1(n13551), .A2(n13982), .ZN(n13485) );
  OAI211_X1 U15502 ( .C1(n13549), .C2(n13739), .A(n13486), .B(n13485), .ZN(
        n13487) );
  AOI21_X1 U15503 ( .B1(n13975), .B2(n13543), .A(n13487), .ZN(n13488) );
  OAI211_X1 U15504 ( .C1(n13977), .C2(n13526), .A(n13489), .B(n13488), .ZN(
        P1_U3226) );
  INV_X1 U15505 ( .A(n14232), .ZN(n13960) );
  AND3_X1 U15506 ( .A1(n13481), .A2(n13491), .A3(n13490), .ZN(n13492) );
  OAI21_X1 U15507 ( .B1(n13493), .B2(n13492), .A(n13537), .ZN(n13498) );
  NOR2_X1 U15508 ( .A1(n13553), .A2(n13954), .ZN(n13496) );
  OAI21_X1 U15509 ( .B1(n13549), .B2(n13955), .A(n13494), .ZN(n13495) );
  AOI211_X1 U15510 ( .C1(n13551), .C2(n13560), .A(n13496), .B(n13495), .ZN(
        n13497) );
  OAI211_X1 U15511 ( .C1(n13960), .C2(n13526), .A(n13498), .B(n13497), .ZN(
        P1_U3228) );
  INV_X1 U15512 ( .A(n13499), .ZN(n13503) );
  NOR3_X1 U15513 ( .A1(n12130), .A2(n13501), .A3(n13500), .ZN(n13502) );
  OAI21_X1 U15514 ( .B1(n13503), .B2(n13502), .A(n13537), .ZN(n13508) );
  INV_X1 U15515 ( .A(n13504), .ZN(n13846) );
  AOI22_X1 U15516 ( .A1(n13981), .A2(n13721), .B1(n13728), .B2(n13983), .ZN(
        n13841) );
  INV_X1 U15517 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n13505) );
  OAI22_X1 U15518 ( .A1(n13540), .A2(n13841), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13505), .ZN(n13506) );
  AOI21_X1 U15519 ( .B1(n13543), .B2(n13846), .A(n13506), .ZN(n13507) );
  OAI211_X1 U15520 ( .C1(n6830), .C2(n13526), .A(n13508), .B(n13507), .ZN(
        P1_U3229) );
  XNOR2_X1 U15521 ( .A(n13510), .B(n13509), .ZN(n13516) );
  AOI22_X1 U15522 ( .A1(n13511), .A2(n13904), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13513) );
  NAND2_X1 U15523 ( .A1(n13551), .A2(n13903), .ZN(n13512) );
  OAI211_X1 U15524 ( .C1(n13553), .C2(n13912), .A(n13513), .B(n13512), .ZN(
        n13514) );
  AOI21_X1 U15525 ( .B1(n13915), .B2(n13555), .A(n13514), .ZN(n13515) );
  OAI21_X1 U15526 ( .B1(n13516), .B2(n13557), .A(n13515), .ZN(P1_U3233) );
  INV_X1 U15527 ( .A(n13517), .ZN(n13521) );
  NOR3_X1 U15528 ( .A1(n13461), .A2(n13519), .A3(n13518), .ZN(n13520) );
  OAI21_X1 U15529 ( .B1(n13521), .B2(n13520), .A(n13537), .ZN(n13525) );
  AOI22_X1 U15530 ( .A1(n13904), .A2(n13981), .B1(n13983), .B2(n13721), .ZN(
        n14064) );
  INV_X1 U15531 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13522) );
  OAI22_X1 U15532 ( .A1(n14064), .A2(n13540), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13522), .ZN(n13523) );
  AOI21_X1 U15533 ( .B1(n13543), .B2(n13878), .A(n13523), .ZN(n13524) );
  OAI211_X1 U15534 ( .C1(n13526), .C2(n14066), .A(n13525), .B(n13524), .ZN(
        P1_U3235) );
  AOI21_X1 U15535 ( .B1(n13528), .B2(n13527), .A(n6465), .ZN(n13533) );
  AOI22_X1 U15536 ( .A1(n13903), .A2(n13983), .B1(n13981), .B2(n13984), .ZN(
        n13937) );
  NAND2_X1 U15537 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13672)
         );
  OAI21_X1 U15538 ( .B1(n13540), .B2(n13937), .A(n13672), .ZN(n13531) );
  NAND2_X1 U15539 ( .A1(n13946), .A2(n14669), .ZN(n14227) );
  INV_X1 U15540 ( .A(n13529), .ZN(n13546) );
  NOR2_X1 U15541 ( .A1(n14227), .A2(n13546), .ZN(n13530) );
  AOI211_X1 U15542 ( .C1(n13945), .C2(n13543), .A(n13531), .B(n13530), .ZN(
        n13532) );
  OAI21_X1 U15543 ( .B1(n13533), .B2(n13557), .A(n13532), .ZN(P1_U3238) );
  NAND2_X1 U15544 ( .A1(n13817), .A2(n14669), .ZN(n14038) );
  OAI21_X1 U15545 ( .B1(n13536), .B2(n13535), .A(n13534), .ZN(n13538) );
  NAND2_X1 U15546 ( .A1(n13538), .A2(n13537), .ZN(n13545) );
  INV_X1 U15547 ( .A(n13815), .ZN(n13542) );
  AOI22_X1 U15548 ( .A1(n13981), .A2(n13728), .B1(n13774), .B2(n13983), .ZN(
        n13808) );
  OAI22_X1 U15549 ( .A1(n13540), .A2(n13808), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13539), .ZN(n13541) );
  AOI21_X1 U15550 ( .B1(n13543), .B2(n13542), .A(n13541), .ZN(n13544) );
  OAI211_X1 U15551 ( .C1(n14038), .C2(n13546), .A(n13545), .B(n13544), .ZN(
        P1_U3240) );
  XNOR2_X1 U15552 ( .A(n13548), .B(n13547), .ZN(n13558) );
  INV_X1 U15553 ( .A(n13992), .ZN(n13709) );
  OAI22_X1 U15554 ( .A1(n13549), .A2(n13994), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14183), .ZN(n13550) );
  AOI21_X1 U15555 ( .B1(n13551), .B2(n13709), .A(n13550), .ZN(n13552) );
  OAI21_X1 U15556 ( .B1(n13553), .B2(n13999), .A(n13552), .ZN(n13554) );
  AOI21_X1 U15557 ( .B1(n14522), .B2(n13555), .A(n13554), .ZN(n13556) );
  OAI21_X1 U15558 ( .B1(n13558), .B2(n13557), .A(n13556), .ZN(P1_U3241) );
  INV_X1 U15559 ( .A(P1_U4016), .ZN(n13574) );
  MUX2_X1 U15560 ( .A(n13699), .B(P1_DATAO_REG_31__SCAN_IN), .S(n13574), .Z(
        P1_U3591) );
  MUX2_X1 U15561 ( .A(n13760), .B(P1_DATAO_REG_30__SCAN_IN), .S(n13573), .Z(
        P1_U3590) );
  MUX2_X1 U15562 ( .A(n13773), .B(P1_DATAO_REG_29__SCAN_IN), .S(n13574), .Z(
        P1_U3589) );
  MUX2_X1 U15563 ( .A(n13765), .B(P1_DATAO_REG_28__SCAN_IN), .S(n13574), .Z(
        P1_U3588) );
  MUX2_X1 U15564 ( .A(n13774), .B(P1_DATAO_REG_27__SCAN_IN), .S(n13574), .Z(
        P1_U3587) );
  MUX2_X1 U15565 ( .A(n13749), .B(P1_DATAO_REG_26__SCAN_IN), .S(n13574), .Z(
        P1_U3586) );
  MUX2_X1 U15566 ( .A(n13728), .B(P1_DATAO_REG_25__SCAN_IN), .S(n13573), .Z(
        P1_U3585) );
  MUX2_X1 U15567 ( .A(n13725), .B(P1_DATAO_REG_24__SCAN_IN), .S(n13574), .Z(
        P1_U3584) );
  MUX2_X1 U15568 ( .A(n13721), .B(P1_DATAO_REG_23__SCAN_IN), .S(n13573), .Z(
        P1_U3583) );
  MUX2_X1 U15569 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n13745), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U15570 ( .A(n13904), .B(P1_DATAO_REG_21__SCAN_IN), .S(n13573), .Z(
        P1_U3581) );
  MUX2_X1 U15571 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13559), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15572 ( .A(n13903), .B(P1_DATAO_REG_19__SCAN_IN), .S(n13573), .Z(
        P1_U3579) );
  MUX2_X1 U15573 ( .A(n13715), .B(P1_DATAO_REG_18__SCAN_IN), .S(n13574), .Z(
        P1_U3578) );
  MUX2_X1 U15574 ( .A(n13984), .B(P1_DATAO_REG_17__SCAN_IN), .S(n13573), .Z(
        P1_U3577) );
  MUX2_X1 U15575 ( .A(n13560), .B(P1_DATAO_REG_16__SCAN_IN), .S(n13573), .Z(
        P1_U3576) );
  MUX2_X1 U15576 ( .A(n13982), .B(P1_DATAO_REG_15__SCAN_IN), .S(n13573), .Z(
        P1_U3575) );
  MUX2_X1 U15577 ( .A(n13709), .B(P1_DATAO_REG_14__SCAN_IN), .S(n13574), .Z(
        P1_U3574) );
  MUX2_X1 U15578 ( .A(n13561), .B(P1_DATAO_REG_13__SCAN_IN), .S(n13573), .Z(
        P1_U3573) );
  MUX2_X1 U15579 ( .A(n13562), .B(P1_DATAO_REG_12__SCAN_IN), .S(n13573), .Z(
        P1_U3572) );
  MUX2_X1 U15580 ( .A(n13563), .B(P1_DATAO_REG_11__SCAN_IN), .S(n13573), .Z(
        P1_U3571) );
  MUX2_X1 U15581 ( .A(n13564), .B(P1_DATAO_REG_10__SCAN_IN), .S(n13574), .Z(
        P1_U3570) );
  MUX2_X1 U15582 ( .A(n13565), .B(P1_DATAO_REG_9__SCAN_IN), .S(n13573), .Z(
        P1_U3569) );
  MUX2_X1 U15583 ( .A(n13566), .B(P1_DATAO_REG_8__SCAN_IN), .S(n13574), .Z(
        P1_U3568) );
  MUX2_X1 U15584 ( .A(n13567), .B(P1_DATAO_REG_7__SCAN_IN), .S(n13573), .Z(
        P1_U3567) );
  MUX2_X1 U15585 ( .A(n13568), .B(P1_DATAO_REG_6__SCAN_IN), .S(n13574), .Z(
        P1_U3566) );
  MUX2_X1 U15586 ( .A(n13569), .B(P1_DATAO_REG_5__SCAN_IN), .S(n13573), .Z(
        P1_U3565) );
  MUX2_X1 U15587 ( .A(n13570), .B(P1_DATAO_REG_4__SCAN_IN), .S(n13574), .Z(
        P1_U3564) );
  MUX2_X1 U15588 ( .A(n13571), .B(P1_DATAO_REG_3__SCAN_IN), .S(n13573), .Z(
        P1_U3563) );
  MUX2_X1 U15589 ( .A(n13572), .B(P1_DATAO_REG_2__SCAN_IN), .S(n13574), .Z(
        P1_U3562) );
  MUX2_X1 U15590 ( .A(n10630), .B(P1_DATAO_REG_1__SCAN_IN), .S(n13573), .Z(
        P1_U3561) );
  MUX2_X1 U15591 ( .A(n13575), .B(P1_DATAO_REG_0__SCAN_IN), .S(n13574), .Z(
        P1_U3560) );
  AOI22_X1 U15592 ( .A1(n14578), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n13584) );
  INV_X1 U15593 ( .A(n13577), .ZN(n13576) );
  NAND2_X1 U15594 ( .A1(n14595), .A2(n13576), .ZN(n13583) );
  MUX2_X1 U15595 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10324), .S(n13577), .Z(
        n13578) );
  OAI21_X1 U15596 ( .B1(n10602), .B2(n7294), .A(n13578), .ZN(n13579) );
  NAND3_X1 U15597 ( .A1(n14597), .A2(n13592), .A3(n13579), .ZN(n13582) );
  OAI211_X1 U15598 ( .C1(n13586), .C2(n13580), .A(n14602), .B(n13600), .ZN(
        n13581) );
  NAND4_X1 U15599 ( .A1(n13584), .A2(n13583), .A3(n13582), .A4(n13581), .ZN(
        P1_U3244) );
  MUX2_X1 U15600 ( .A(n13586), .B(n13585), .S(n6588), .Z(n13588) );
  NAND2_X1 U15601 ( .A1(n13588), .A2(n13587), .ZN(n13589) );
  OAI211_X1 U15602 ( .C1(n14284), .C2(n13590), .A(n13589), .B(P1_U4016), .ZN(
        n14589) );
  AOI22_X1 U15603 ( .A1(n14578), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n13605) );
  MUX2_X1 U15604 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10323), .S(n13598), .Z(
        n13593) );
  NAND3_X1 U15605 ( .A1(n13593), .A2(n13592), .A3(n13591), .ZN(n13595) );
  AND2_X1 U15606 ( .A1(n13595), .A2(n13594), .ZN(n13597) );
  AOI22_X1 U15607 ( .A1(n14597), .A2(n13597), .B1(n14595), .B2(n13596), .ZN(
        n13604) );
  MUX2_X1 U15608 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10339), .S(n13598), .Z(
        n13601) );
  NAND3_X1 U15609 ( .A1(n13601), .A2(n13600), .A3(n13599), .ZN(n13602) );
  NAND3_X1 U15610 ( .A1(n14602), .A2(n13609), .A3(n13602), .ZN(n13603) );
  NAND4_X1 U15611 ( .A1(n14589), .A2(n13605), .A3(n13604), .A4(n13603), .ZN(
        P1_U3245) );
  OAI22_X1 U15612 ( .A1(n14593), .A2(n14293), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9266), .ZN(n13606) );
  AOI21_X1 U15613 ( .B1(n13607), .B2(n14595), .A(n13606), .ZN(n13618) );
  MUX2_X1 U15614 ( .A(n10338), .B(P1_REG2_REG_3__SCAN_IN), .S(n13607), .Z(
        n13610) );
  NAND3_X1 U15615 ( .A1(n13610), .A2(n13609), .A3(n13608), .ZN(n13611) );
  NAND3_X1 U15616 ( .A1(n14602), .A2(n14582), .A3(n13611), .ZN(n13617) );
  OR3_X1 U15617 ( .A1(n13614), .A2(n13613), .A3(n13612), .ZN(n13615) );
  NAND3_X1 U15618 ( .A1(n14597), .A2(n14574), .A3(n13615), .ZN(n13616) );
  NAND3_X1 U15619 ( .A1(n13618), .A2(n13617), .A3(n13616), .ZN(P1_U3246) );
  OAI21_X1 U15620 ( .B1(n14593), .B2(n14341), .A(n13619), .ZN(n13620) );
  AOI21_X1 U15621 ( .B1(n13621), .B2(n14595), .A(n13620), .ZN(n13632) );
  MUX2_X1 U15622 ( .A(n11083), .B(P1_REG2_REG_5__SCAN_IN), .S(n13621), .Z(
        n13622) );
  NAND3_X1 U15623 ( .A1(n14584), .A2(n13623), .A3(n13622), .ZN(n13624) );
  NAND3_X1 U15624 ( .A1(n14602), .A2(n13625), .A3(n13624), .ZN(n13631) );
  OAI21_X1 U15625 ( .B1(n13628), .B2(n13627), .A(n13626), .ZN(n13629) );
  NAND2_X1 U15626 ( .A1(n14597), .A2(n13629), .ZN(n13630) );
  NAND3_X1 U15627 ( .A1(n13632), .A2(n13631), .A3(n13630), .ZN(P1_U3248) );
  AOI22_X1 U15628 ( .A1(n14578), .A2(P1_ADDR_REG_7__SCAN_IN), .B1(
        P1_REG3_REG_7__SCAN_IN), .B2(P1_U3086), .ZN(n13647) );
  NAND2_X1 U15629 ( .A1(n14595), .A2(n13638), .ZN(n13646) );
  OR3_X1 U15630 ( .A1(n13635), .A2(n13634), .A3(n13633), .ZN(n13636) );
  NAND3_X1 U15631 ( .A1(n14597), .A2(n13637), .A3(n13636), .ZN(n13645) );
  MUX2_X1 U15632 ( .A(n11513), .B(P1_REG2_REG_7__SCAN_IN), .S(n13638), .Z(
        n13639) );
  NAND3_X1 U15633 ( .A1(n13641), .A2(n13640), .A3(n13639), .ZN(n13642) );
  NAND3_X1 U15634 ( .A1(n14602), .A2(n13643), .A3(n13642), .ZN(n13644) );
  NAND4_X1 U15635 ( .A1(n13647), .A2(n13646), .A3(n13645), .A4(n13644), .ZN(
        P1_U3250) );
  INV_X1 U15636 ( .A(n13648), .ZN(n13653) );
  NOR3_X1 U15637 ( .A1(n13651), .A2(n13650), .A3(n13649), .ZN(n13652) );
  OAI21_X1 U15638 ( .B1(n13653), .B2(n13652), .A(n14597), .ZN(n13664) );
  OAI21_X1 U15639 ( .B1(n14593), .B2(n14309), .A(n13654), .ZN(n13655) );
  AOI21_X1 U15640 ( .B1(n13656), .B2(n14595), .A(n13655), .ZN(n13663) );
  MUX2_X1 U15641 ( .A(n11307), .B(P1_REG2_REG_9__SCAN_IN), .S(n13656), .Z(
        n13657) );
  NAND3_X1 U15642 ( .A1(n13659), .A2(n13658), .A3(n13657), .ZN(n13660) );
  NAND3_X1 U15643 ( .A1(n14602), .A2(n13661), .A3(n13660), .ZN(n13662) );
  NAND3_X1 U15644 ( .A1(n13664), .A2(n13663), .A3(n13662), .ZN(P1_U3252) );
  OAI21_X1 U15645 ( .B1(n13959), .B2(n13668), .A(n13665), .ZN(n13682) );
  XOR2_X1 U15646 ( .A(n13683), .B(n13682), .Z(n13666) );
  NAND2_X1 U15647 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n13666), .ZN(n13685) );
  OAI211_X1 U15648 ( .C1(n13666), .C2(P1_REG2_REG_18__SCAN_IN), .A(n14602), 
        .B(n13685), .ZN(n13675) );
  OAI21_X1 U15649 ( .B1(n13669), .B2(n13668), .A(n13667), .ZN(n13678) );
  XNOR2_X1 U15650 ( .A(n13678), .B(n13676), .ZN(n13670) );
  NAND2_X1 U15651 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n13670), .ZN(n13680) );
  OAI211_X1 U15652 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n13670), .A(n14597), 
        .B(n13680), .ZN(n13671) );
  NAND2_X1 U15653 ( .A1(n13672), .A2(n13671), .ZN(n13673) );
  AOI21_X1 U15654 ( .B1(n14578), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n13673), 
        .ZN(n13674) );
  OAI211_X1 U15655 ( .C1(n13677), .C2(n13676), .A(n13675), .B(n13674), .ZN(
        P1_U3261) );
  NAND2_X1 U15656 ( .A1(n13683), .A2(n13678), .ZN(n13679) );
  NAND2_X1 U15657 ( .A1(n13680), .A2(n13679), .ZN(n13681) );
  XOR2_X1 U15658 ( .A(n13681), .B(P1_REG1_REG_19__SCAN_IN), .Z(n13689) );
  NAND2_X1 U15659 ( .A1(n13683), .A2(n13682), .ZN(n13684) );
  NAND2_X1 U15660 ( .A1(n13685), .A2(n13684), .ZN(n13686) );
  XOR2_X1 U15661 ( .A(n13686), .B(P1_REG2_REG_19__SCAN_IN), .Z(n13687) );
  AOI22_X1 U15662 ( .A1(n13689), .A2(n14597), .B1(n14602), .B2(n13687), .ZN(
        n13692) );
  INV_X1 U15663 ( .A(n13687), .ZN(n13690) );
  AOI21_X1 U15664 ( .B1(n14578), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n13693), 
        .ZN(n13694) );
  INV_X1 U15665 ( .A(n13946), .ZN(n13695) );
  INV_X1 U15666 ( .A(n13817), .ZN(n13750) );
  NAND2_X1 U15667 ( .A1(n13696), .A2(n14618), .ZN(n14012) );
  NOR2_X1 U15668 ( .A1(n6588), .A2(n13697), .ZN(n13698) );
  NOR2_X1 U15669 ( .A1(n13993), .A2(n13698), .ZN(n13759) );
  NAND2_X1 U15670 ( .A1(n13759), .A2(n13699), .ZN(n14014) );
  NOR2_X1 U15671 ( .A1(n14647), .A2(n14014), .ZN(n13703) );
  NOR2_X1 U15672 ( .A1(n14013), .A2(n14002), .ZN(n13700) );
  AOI211_X1 U15673 ( .C1(n14647), .C2(P1_REG2_REG_31__SCAN_IN), .A(n13703), 
        .B(n13700), .ZN(n13701) );
  OAI21_X1 U15674 ( .B1(n14012), .B2(n14643), .A(n13701), .ZN(P1_U3263) );
  OAI211_X1 U15675 ( .C1(n14016), .C2(n13756), .A(n13702), .B(n14618), .ZN(
        n14015) );
  INV_X1 U15676 ( .A(n13703), .ZN(n13704) );
  OAI21_X1 U15677 ( .B1(n13962), .B2(n13705), .A(n13704), .ZN(n13706) );
  AOI21_X1 U15678 ( .B1(n13707), .B2(n14634), .A(n13706), .ZN(n13708) );
  OAI21_X1 U15679 ( .B1(n14015), .B2(n14643), .A(n13708), .ZN(P1_U3264) );
  NAND2_X1 U15680 ( .A1(n14528), .A2(n13709), .ZN(n13710) );
  INV_X1 U15681 ( .A(n13989), .ZN(n14007) );
  OR2_X1 U15682 ( .A1(n14522), .A2(n13982), .ZN(n13711) );
  NAND2_X1 U15683 ( .A1(n14004), .A2(n13711), .ZN(n13972) );
  NAND2_X1 U15684 ( .A1(n13977), .A2(n13994), .ZN(n13712) );
  OR2_X1 U15685 ( .A1(n13946), .A2(n13715), .ZN(n13716) );
  OR2_X1 U15686 ( .A1(n14082), .A2(n13743), .ZN(n13718) );
  INV_X1 U15687 ( .A(n13897), .ZN(n13886) );
  OR2_X1 U15688 ( .A1(n14073), .A2(n13904), .ZN(n13719) );
  NOR2_X1 U15689 ( .A1(n13875), .A2(n13745), .ZN(n13720) );
  NAND2_X1 U15690 ( .A1(n13864), .A2(n13863), .ZN(n13865) );
  NAND2_X1 U15691 ( .A1(n14058), .A2(n13721), .ZN(n13722) );
  NAND2_X1 U15692 ( .A1(n13865), .A2(n13722), .ZN(n13850) );
  INV_X1 U15693 ( .A(n13850), .ZN(n13724) );
  OR2_X1 U15694 ( .A1(n14051), .A2(n13725), .ZN(n13726) );
  NAND2_X1 U15695 ( .A1(n13817), .A2(n13749), .ZN(n13729) );
  OR2_X1 U15696 ( .A1(n14034), .A2(n13774), .ZN(n13730) );
  INV_X1 U15697 ( .A(n13784), .ZN(n13731) );
  INV_X1 U15698 ( .A(n13735), .ZN(n13736) );
  NAND2_X1 U15699 ( .A1(n13979), .A2(n13980), .ZN(n13978) );
  NAND2_X1 U15700 ( .A1(n13978), .A2(n13738), .ZN(n13951) );
  NAND2_X1 U15701 ( .A1(n13960), .A2(n13984), .ZN(n13740) );
  NAND2_X1 U15702 ( .A1(n13936), .A2(n13935), .ZN(n13934) );
  INV_X1 U15703 ( .A(n13863), .ZN(n13855) );
  OAI22_X1 U15704 ( .A1(n6694), .A2(n13753), .B1(n13752), .B2(n14028), .ZN(
        n13755) );
  XNOR2_X1 U15705 ( .A(n13755), .B(n13754), .ZN(n14024) );
  INV_X1 U15706 ( .A(n13779), .ZN(n13757) );
  AOI211_X1 U15707 ( .C1(n13758), .C2(n13757), .A(n14636), .B(n13756), .ZN(
        n14017) );
  NAND2_X1 U15708 ( .A1(n14017), .A2(n14623), .ZN(n13769) );
  NAND2_X1 U15709 ( .A1(n13760), .A2(n13759), .ZN(n14018) );
  OR3_X1 U15710 ( .A1(n13762), .A2(n14018), .A3(n13761), .ZN(n13763) );
  OAI21_X1 U15711 ( .B1(n13913), .B2(n13764), .A(n13763), .ZN(n13767) );
  NAND2_X1 U15712 ( .A1(n13765), .A2(n13981), .ZN(n14019) );
  NOR2_X1 U15713 ( .A1(n14647), .A2(n14019), .ZN(n13766) );
  AOI211_X1 U15714 ( .C1(n14647), .C2(P1_REG2_REG_29__SCAN_IN), .A(n13767), 
        .B(n13766), .ZN(n13768) );
  OAI211_X1 U15715 ( .C1(n14020), .C2(n14002), .A(n13769), .B(n13768), .ZN(
        n13770) );
  AOI21_X1 U15716 ( .B1(n14024), .B2(n13869), .A(n13770), .ZN(n13771) );
  OAI21_X1 U15717 ( .B1(n14026), .B2(n14008), .A(n13771), .ZN(P1_U3356) );
  XNOR2_X1 U15718 ( .A(n13772), .B(n13731), .ZN(n13778) );
  NAND2_X1 U15719 ( .A1(n13773), .A2(n13983), .ZN(n13776) );
  NAND2_X1 U15720 ( .A1(n13774), .A2(n13981), .ZN(n13775) );
  AOI211_X1 U15721 ( .C1(n14028), .C2(n13798), .A(n14636), .B(n13779), .ZN(
        n14027) );
  INV_X1 U15722 ( .A(n13780), .ZN(n13781) );
  AOI22_X1 U15723 ( .A1(n14647), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n13781), 
        .B2(n14635), .ZN(n13782) );
  OAI21_X1 U15724 ( .B1(n13783), .B2(n14002), .A(n13782), .ZN(n13789) );
  NAND2_X1 U15725 ( .A1(n13785), .A2(n13784), .ZN(n13786) );
  NAND2_X1 U15726 ( .A1(n13787), .A2(n13786), .ZN(n14031) );
  NOR2_X1 U15727 ( .A1(n14031), .A2(n14008), .ZN(n13788) );
  OAI21_X1 U15728 ( .B1(n14030), .B2(n14647), .A(n13790), .ZN(P1_U3265) );
  XNOR2_X1 U15729 ( .A(n13792), .B(n13791), .ZN(n13795) );
  INV_X1 U15730 ( .A(n13793), .ZN(n13794) );
  AOI21_X1 U15731 ( .B1(n13795), .B2(n14708), .A(n13794), .ZN(n14036) );
  OAI21_X1 U15732 ( .B1(n6699), .B2(n13797), .A(n13796), .ZN(n14032) );
  INV_X1 U15733 ( .A(n13798), .ZN(n13799) );
  AOI211_X1 U15734 ( .C1(n14034), .C2(n13800), .A(n14636), .B(n13799), .ZN(
        n14033) );
  NAND2_X1 U15735 ( .A1(n14033), .A2(n14623), .ZN(n13803) );
  AOI22_X1 U15736 ( .A1(n14647), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n13801), 
        .B2(n14635), .ZN(n13802) );
  OAI211_X1 U15737 ( .C1(n13804), .C2(n14002), .A(n13803), .B(n13802), .ZN(
        n13805) );
  AOI21_X1 U15738 ( .B1(n14032), .B2(n13967), .A(n13805), .ZN(n13806) );
  OAI21_X1 U15739 ( .B1(n14036), .B2(n14647), .A(n13806), .ZN(P1_U3266) );
  XOR2_X1 U15740 ( .A(n13811), .B(n13807), .Z(n13809) );
  OAI21_X1 U15741 ( .B1(n13809), .B2(n14077), .A(n13808), .ZN(n14042) );
  OAI21_X1 U15742 ( .B1(n13812), .B2(n13811), .A(n13810), .ZN(n14040) );
  NOR2_X1 U15743 ( .A1(n14040), .A2(n14008), .ZN(n13820) );
  XNOR2_X1 U15744 ( .A(n13826), .B(n13817), .ZN(n13813) );
  NAND2_X1 U15745 ( .A1(n13813), .A2(n14618), .ZN(n14039) );
  NAND2_X1 U15746 ( .A1(n14647), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n13814) );
  OAI21_X1 U15747 ( .B1(n13913), .B2(n13815), .A(n13814), .ZN(n13816) );
  AOI21_X1 U15748 ( .B1(n13817), .B2(n14634), .A(n13816), .ZN(n13818) );
  OAI21_X1 U15749 ( .B1(n14039), .B2(n14643), .A(n13818), .ZN(n13819) );
  AOI211_X1 U15750 ( .C1(n14042), .C2(n13962), .A(n13820), .B(n13819), .ZN(
        n13821) );
  INV_X1 U15751 ( .A(n13821), .ZN(P1_U3267) );
  AOI21_X1 U15752 ( .B1(n13727), .B2(n13823), .A(n13822), .ZN(n14049) );
  INV_X1 U15753 ( .A(n13869), .ZN(n13970) );
  NAND2_X1 U15754 ( .A1(n14045), .A2(n13843), .ZN(n13824) );
  NAND2_X1 U15755 ( .A1(n13824), .A2(n14618), .ZN(n13825) );
  NOR2_X1 U15756 ( .A1(n13826), .A2(n13825), .ZN(n14043) );
  NAND2_X1 U15757 ( .A1(n14045), .A2(n14634), .ZN(n13832) );
  INV_X1 U15758 ( .A(n14044), .ZN(n13828) );
  OAI22_X1 U15759 ( .A1(n14647), .A2(n13828), .B1(n13827), .B2(n13913), .ZN(
        n13829) );
  INV_X1 U15760 ( .A(n13829), .ZN(n13831) );
  NAND2_X1 U15761 ( .A1(n14647), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n13830) );
  NAND3_X1 U15762 ( .A1(n13832), .A2(n13831), .A3(n13830), .ZN(n13833) );
  AOI21_X1 U15763 ( .B1(n14043), .B2(n14623), .A(n13833), .ZN(n13838) );
  NAND2_X1 U15764 ( .A1(n13836), .A2(n13835), .ZN(n14046) );
  NAND3_X1 U15765 ( .A1(n13834), .A2(n13967), .A3(n14046), .ZN(n13837) );
  OAI211_X1 U15766 ( .C1(n14049), .C2(n13970), .A(n13838), .B(n13837), .ZN(
        P1_U3268) );
  OAI211_X1 U15767 ( .C1(n13840), .C2(n13851), .A(n13839), .B(n14708), .ZN(
        n13842) );
  INV_X1 U15768 ( .A(n13843), .ZN(n13844) );
  AOI211_X1 U15769 ( .C1(n14051), .C2(n13845), .A(n14636), .B(n13844), .ZN(
        n14050) );
  AOI22_X1 U15770 ( .A1(n14647), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n13846), 
        .B2(n14635), .ZN(n13847) );
  OAI21_X1 U15771 ( .B1(n6830), .B2(n14002), .A(n13847), .ZN(n13853) );
  INV_X1 U15772 ( .A(n13848), .ZN(n13849) );
  AOI21_X1 U15773 ( .B1(n13851), .B2(n13850), .A(n13849), .ZN(n14054) );
  NOR2_X1 U15774 ( .A1(n14054), .A2(n14008), .ZN(n13852) );
  AOI211_X1 U15775 ( .C1(n14050), .C2(n14623), .A(n13853), .B(n13852), .ZN(
        n13854) );
  OAI21_X1 U15776 ( .B1(n14647), .B2(n14052), .A(n13854), .ZN(P1_U3269) );
  XNOR2_X1 U15777 ( .A(n13856), .B(n13855), .ZN(n14055) );
  INV_X1 U15778 ( .A(n13876), .ZN(n13857) );
  XNOR2_X1 U15779 ( .A(n14058), .B(n13857), .ZN(n13858) );
  NAND2_X1 U15780 ( .A1(n13858), .A2(n14618), .ZN(n14060) );
  OAI22_X1 U15781 ( .A1(n14056), .A2(n14647), .B1(n13859), .B2(n13913), .ZN(
        n13862) );
  NOR2_X1 U15782 ( .A1(n13860), .A2(n14002), .ZN(n13861) );
  AOI211_X1 U15783 ( .C1(n14647), .C2(P1_REG2_REG_23__SCAN_IN), .A(n13862), 
        .B(n13861), .ZN(n13867) );
  OR2_X1 U15784 ( .A1(n13864), .A2(n13863), .ZN(n14059) );
  NAND3_X1 U15785 ( .A1(n14059), .A2(n13865), .A3(n13967), .ZN(n13866) );
  OAI211_X1 U15786 ( .C1(n14060), .C2(n14643), .A(n13867), .B(n13866), .ZN(
        n13868) );
  AOI21_X1 U15787 ( .B1(n13869), .B2(n14055), .A(n13868), .ZN(n13870) );
  INV_X1 U15788 ( .A(n13870), .ZN(P1_U3270) );
  XOR2_X1 U15789 ( .A(n13873), .B(n13871), .Z(n14070) );
  XNOR2_X1 U15790 ( .A(n13872), .B(n13873), .ZN(n14068) );
  INV_X1 U15791 ( .A(n13874), .ZN(n13888) );
  AOI21_X1 U15792 ( .B1(n13875), .B2(n13888), .A(n14636), .ZN(n13877) );
  NAND2_X1 U15793 ( .A1(n13877), .A2(n13876), .ZN(n14065) );
  INV_X1 U15794 ( .A(n13878), .ZN(n13879) );
  OAI22_X1 U15795 ( .A1(n14064), .A2(n14647), .B1(n13879), .B2(n13913), .ZN(
        n13881) );
  NOR2_X1 U15796 ( .A1(n14066), .A2(n14002), .ZN(n13880) );
  AOI211_X1 U15797 ( .C1(n14647), .C2(P1_REG2_REG_22__SCAN_IN), .A(n13881), 
        .B(n13880), .ZN(n13882) );
  OAI21_X1 U15798 ( .B1(n14643), .B2(n14065), .A(n13882), .ZN(n13883) );
  AOI21_X1 U15799 ( .B1(n13967), .B2(n14068), .A(n13883), .ZN(n13884) );
  OAI21_X1 U15800 ( .B1(n14070), .B2(n13970), .A(n13884), .ZN(P1_U3271) );
  OAI21_X1 U15801 ( .B1(n13887), .B2(n13886), .A(n13885), .ZN(n14078) );
  AOI21_X1 U15802 ( .B1(n14073), .B2(n13907), .A(n14636), .ZN(n13889) );
  AND2_X1 U15803 ( .A1(n13889), .A2(n13888), .ZN(n14071) );
  NAND2_X1 U15804 ( .A1(n14073), .A2(n14634), .ZN(n13894) );
  NOR2_X1 U15805 ( .A1(n13890), .A2(n13913), .ZN(n13891) );
  AOI21_X1 U15806 ( .B1(n13962), .B2(n14072), .A(n13891), .ZN(n13893) );
  NAND2_X1 U15807 ( .A1(n14647), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n13892) );
  NAND3_X1 U15808 ( .A1(n13894), .A2(n13893), .A3(n13892), .ZN(n13895) );
  AOI21_X1 U15809 ( .B1(n14071), .B2(n14623), .A(n13895), .ZN(n13900) );
  OAI21_X1 U15810 ( .B1(n13898), .B2(n13897), .A(n13896), .ZN(n14074) );
  NAND2_X1 U15811 ( .A1(n14074), .A2(n13967), .ZN(n13899) );
  OAI211_X1 U15812 ( .C1(n14078), .C2(n13970), .A(n13900), .B(n13899), .ZN(
        P1_U3272) );
  OAI211_X1 U15813 ( .C1(n13902), .C2(n13909), .A(n13901), .B(n14708), .ZN(
        n13906) );
  AOI22_X1 U15814 ( .A1(n13904), .A2(n13983), .B1(n13981), .B2(n13903), .ZN(
        n13905) );
  NAND2_X1 U15815 ( .A1(n13906), .A2(n13905), .ZN(n14084) );
  OAI211_X1 U15816 ( .C1(n14082), .C2(n6540), .A(n14618), .B(n13907), .ZN(
        n14080) );
  NAND2_X1 U15817 ( .A1(n13910), .A2(n13909), .ZN(n14079) );
  NAND3_X1 U15818 ( .A1(n13908), .A2(n14079), .A3(n13967), .ZN(n13917) );
  NAND2_X1 U15819 ( .A1(n14647), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n13911) );
  OAI21_X1 U15820 ( .B1(n13913), .B2(n13912), .A(n13911), .ZN(n13914) );
  AOI21_X1 U15821 ( .B1(n13915), .B2(n14634), .A(n13914), .ZN(n13916) );
  OAI211_X1 U15822 ( .C1(n14080), .C2(n14643), .A(n13917), .B(n13916), .ZN(
        n13918) );
  AOI21_X1 U15823 ( .B1(n14084), .B2(n13962), .A(n13918), .ZN(n13919) );
  INV_X1 U15824 ( .A(n13919), .ZN(P1_U3273) );
  XOR2_X1 U15825 ( .A(n13920), .B(n13928), .Z(n14224) );
  NAND2_X1 U15826 ( .A1(n13943), .A2(n14221), .ZN(n13921) );
  NAND2_X1 U15827 ( .A1(n13921), .A2(n14618), .ZN(n13922) );
  NOR2_X1 U15828 ( .A1(n6540), .A2(n13922), .ZN(n14219) );
  INV_X1 U15829 ( .A(n13923), .ZN(n13924) );
  AOI22_X1 U15830 ( .A1(n14647), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n13924), 
        .B2(n14635), .ZN(n13925) );
  OAI21_X1 U15831 ( .B1(n6826), .B2(n14002), .A(n13925), .ZN(n13932) );
  AOI21_X1 U15832 ( .B1(n13928), .B2(n13927), .A(n13926), .ZN(n13929) );
  OR2_X1 U15833 ( .A1(n13929), .A2(n14077), .ZN(n14222) );
  INV_X1 U15834 ( .A(n14220), .ZN(n13930) );
  AOI21_X1 U15835 ( .B1(n14222), .B2(n13930), .A(n14647), .ZN(n13931) );
  AOI211_X1 U15836 ( .C1(n14219), .C2(n14623), .A(n13932), .B(n13931), .ZN(
        n13933) );
  OAI21_X1 U15837 ( .B1(n14008), .B2(n14224), .A(n13933), .ZN(P1_U3274) );
  OAI211_X1 U15838 ( .C1(n13936), .C2(n13935), .A(n13934), .B(n14708), .ZN(
        n13938) );
  AND2_X1 U15839 ( .A1(n13938), .A2(n13937), .ZN(n14228) );
  INV_X1 U15840 ( .A(n13939), .ZN(n13941) );
  OAI21_X1 U15841 ( .B1(n13941), .B2(n13940), .A(n6446), .ZN(n14225) );
  INV_X1 U15842 ( .A(n13942), .ZN(n13953) );
  AOI21_X1 U15843 ( .B1(n13946), .B2(n13953), .A(n14636), .ZN(n13944) );
  NAND2_X1 U15844 ( .A1(n13944), .A2(n13943), .ZN(n14226) );
  AOI22_X1 U15845 ( .A1(n14647), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n13945), 
        .B2(n14635), .ZN(n13948) );
  NAND2_X1 U15846 ( .A1(n13946), .A2(n14634), .ZN(n13947) );
  OAI211_X1 U15847 ( .C1(n14226), .C2(n14643), .A(n13948), .B(n13947), .ZN(
        n13949) );
  AOI21_X1 U15848 ( .B1(n14225), .B2(n13967), .A(n13949), .ZN(n13950) );
  OAI21_X1 U15849 ( .B1(n14647), .B2(n14228), .A(n13950), .ZN(P1_U3275) );
  XNOR2_X1 U15850 ( .A(n13951), .B(n13966), .ZN(n14237) );
  INV_X1 U15851 ( .A(n14237), .ZN(n13971) );
  NAND2_X1 U15852 ( .A1(n14232), .A2(n13974), .ZN(n13952) );
  NAND2_X1 U15853 ( .A1(n13953), .A2(n13952), .ZN(n14235) );
  INV_X1 U15854 ( .A(n13954), .ZN(n13956) );
  OAI22_X1 U15855 ( .A1(n13955), .A2(n13993), .B1(n13994), .B2(n13991), .ZN(
        n14231) );
  AOI21_X1 U15856 ( .B1(n13956), .B2(n14635), .A(n14231), .ZN(n13957) );
  OAI21_X1 U15857 ( .B1(n14235), .B2(n13958), .A(n13957), .ZN(n13963) );
  OAI22_X1 U15858 ( .A1(n13960), .A2(n14002), .B1(n13959), .B2(n13962), .ZN(
        n13961) );
  AOI21_X1 U15859 ( .B1(n13963), .B2(n13962), .A(n13961), .ZN(n13969) );
  NAND2_X1 U15860 ( .A1(n13965), .A2(n13966), .ZN(n14230) );
  NAND3_X1 U15861 ( .A1(n13964), .A2(n14230), .A3(n13967), .ZN(n13968) );
  OAI211_X1 U15862 ( .C1(n13971), .C2(n13970), .A(n13969), .B(n13968), .ZN(
        P1_U3276) );
  XNOR2_X1 U15863 ( .A(n13972), .B(n13980), .ZN(n14243) );
  OR2_X1 U15864 ( .A1(n13977), .A2(n13997), .ZN(n13973) );
  AND3_X1 U15865 ( .A1(n13974), .A2(n13973), .A3(n14618), .ZN(n14239) );
  AOI22_X1 U15866 ( .A1(n14647), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n13975), 
        .B2(n14635), .ZN(n13976) );
  OAI21_X1 U15867 ( .B1(n13977), .B2(n14002), .A(n13976), .ZN(n13987) );
  OAI21_X1 U15868 ( .B1(n13980), .B2(n13979), .A(n13978), .ZN(n13985) );
  AOI222_X1 U15869 ( .A1(n14708), .A2(n13985), .B1(n13984), .B2(n13983), .C1(
        n13982), .C2(n13981), .ZN(n14242) );
  NOR2_X1 U15870 ( .A1(n14242), .A2(n14647), .ZN(n13986) );
  AOI211_X1 U15871 ( .C1(n14239), .C2(n14623), .A(n13987), .B(n13986), .ZN(
        n13988) );
  OAI21_X1 U15872 ( .B1(n14243), .B2(n14008), .A(n13988), .ZN(P1_U3277) );
  XNOR2_X1 U15873 ( .A(n13990), .B(n13989), .ZN(n13996) );
  OAI22_X1 U15874 ( .A1(n13994), .A2(n13993), .B1(n13992), .B2(n13991), .ZN(
        n13995) );
  AOI21_X1 U15875 ( .B1(n13996), .B2(n14708), .A(n13995), .ZN(n14524) );
  AOI211_X1 U15876 ( .C1(n14522), .C2(n13998), .A(n14636), .B(n13997), .ZN(
        n14521) );
  INV_X1 U15877 ( .A(n13999), .ZN(n14000) );
  AOI22_X1 U15878 ( .A1(n14647), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n14000), 
        .B2(n14635), .ZN(n14001) );
  OAI21_X1 U15879 ( .B1(n14003), .B2(n14002), .A(n14001), .ZN(n14010) );
  INV_X1 U15880 ( .A(n14004), .ZN(n14005) );
  AOI21_X1 U15881 ( .B1(n14007), .B2(n14006), .A(n14005), .ZN(n14526) );
  NOR2_X1 U15882 ( .A1(n14526), .A2(n14008), .ZN(n14009) );
  AOI211_X1 U15883 ( .C1(n14623), .C2(n14521), .A(n14010), .B(n14009), .ZN(
        n14011) );
  OAI21_X1 U15884 ( .B1(n14647), .B2(n14524), .A(n14011), .ZN(P1_U3278) );
  OAI211_X1 U15885 ( .C1(n14013), .C2(n14726), .A(n14012), .B(n14014), .ZN(
        n14244) );
  MUX2_X1 U15886 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14244), .S(n14745), .Z(
        P1_U3559) );
  OAI211_X1 U15887 ( .C1(n14016), .C2(n14726), .A(n14015), .B(n14014), .ZN(
        n14245) );
  MUX2_X1 U15888 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14245), .S(n14745), .Z(
        P1_U3558) );
  OAI211_X1 U15889 ( .C1(n14020), .C2(n14726), .A(n14019), .B(n14018), .ZN(
        n14021) );
  INV_X1 U15890 ( .A(n14021), .ZN(n14022) );
  NAND2_X1 U15891 ( .A1(n14024), .A2(n14708), .ZN(n14025) );
  MUX2_X1 U15892 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14246), .S(n14745), .Z(
        P1_U3557) );
  AOI21_X1 U15893 ( .B1(n14669), .B2(n14028), .A(n14027), .ZN(n14029) );
  OAI211_X1 U15894 ( .C1(n14525), .C2(n14031), .A(n14030), .B(n14029), .ZN(
        n14247) );
  MUX2_X1 U15895 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14247), .S(n14745), .Z(
        P1_U3556) );
  INV_X1 U15896 ( .A(n14032), .ZN(n14037) );
  AOI21_X1 U15897 ( .B1(n14669), .B2(n14034), .A(n14033), .ZN(n14035) );
  OAI211_X1 U15898 ( .C1(n14525), .C2(n14037), .A(n14036), .B(n14035), .ZN(
        n14248) );
  MUX2_X1 U15899 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14248), .S(n14745), .Z(
        P1_U3555) );
  OAI211_X1 U15900 ( .C1(n14040), .C2(n14525), .A(n14039), .B(n14038), .ZN(
        n14041) );
  MUX2_X1 U15901 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14249), .S(n14745), .Z(
        P1_U3554) );
  AOI211_X1 U15902 ( .C1(n14669), .C2(n14045), .A(n14044), .B(n14043), .ZN(
        n14048) );
  NAND3_X1 U15903 ( .A1(n13834), .A2(n14729), .A3(n14046), .ZN(n14047) );
  OAI211_X1 U15904 ( .C1(n14049), .C2(n14077), .A(n14048), .B(n14047), .ZN(
        n14250) );
  MUX2_X1 U15905 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14250), .S(n14745), .Z(
        P1_U3553) );
  AOI21_X1 U15906 ( .B1(n14669), .B2(n14051), .A(n14050), .ZN(n14053) );
  OAI211_X1 U15907 ( .C1(n14525), .C2(n14054), .A(n14053), .B(n14052), .ZN(
        n14251) );
  MUX2_X1 U15908 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14251), .S(n14745), .Z(
        P1_U3552) );
  NAND2_X1 U15909 ( .A1(n14055), .A2(n14708), .ZN(n14063) );
  INV_X1 U15910 ( .A(n14056), .ZN(n14057) );
  AOI21_X1 U15911 ( .B1(n14058), .B2(n14669), .A(n14057), .ZN(n14062) );
  NAND3_X1 U15912 ( .A1(n13865), .A2(n14059), .A3(n14729), .ZN(n14061) );
  NAND4_X1 U15913 ( .A1(n14063), .A2(n14062), .A3(n14061), .A4(n14060), .ZN(
        n14252) );
  MUX2_X1 U15914 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14252), .S(n14745), .Z(
        P1_U3551) );
  OAI211_X1 U15915 ( .C1(n14726), .C2(n14066), .A(n14065), .B(n14064), .ZN(
        n14067) );
  AOI21_X1 U15916 ( .B1(n14068), .B2(n14729), .A(n14067), .ZN(n14069) );
  OAI21_X1 U15917 ( .B1(n14070), .B2(n14077), .A(n14069), .ZN(n14253) );
  MUX2_X1 U15918 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14253), .S(n14745), .Z(
        P1_U3550) );
  AOI211_X1 U15919 ( .C1(n14669), .C2(n14073), .A(n14072), .B(n14071), .ZN(
        n14076) );
  NAND2_X1 U15920 ( .A1(n14074), .A2(n14729), .ZN(n14075) );
  OAI211_X1 U15921 ( .C1(n14078), .C2(n14077), .A(n14076), .B(n14075), .ZN(
        n14254) );
  MUX2_X1 U15922 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14254), .S(n14745), .Z(
        P1_U3549) );
  NAND3_X1 U15923 ( .A1(n13908), .A2(n14079), .A3(n14729), .ZN(n14081) );
  OAI211_X1 U15924 ( .C1(n14082), .C2(n14726), .A(n14081), .B(n14080), .ZN(
        n14083) );
  NOR2_X1 U15925 ( .A1(n14084), .A2(n14083), .ZN(n14256) );
  MUX2_X1 U15926 ( .A(n14085), .B(n14256), .S(n14745), .Z(n14218) );
  INV_X1 U15927 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14384) );
  AOI22_X1 U15928 ( .A1(n14087), .A2(keyinput27), .B1(keyinput9), .B2(n14384), 
        .ZN(n14086) );
  OAI221_X1 U15929 ( .B1(n14087), .B2(keyinput27), .C1(n14384), .C2(keyinput9), 
        .A(n14086), .ZN(n14092) );
  AOI22_X1 U15930 ( .A1(n14085), .A2(keyinput21), .B1(n14182), .B2(keyinput48), 
        .ZN(n14088) );
  OAI221_X1 U15931 ( .B1(n14085), .B2(keyinput21), .C1(n14182), .C2(keyinput48), .A(n14088), .ZN(n14091) );
  INV_X1 U15932 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n14872) );
  XNOR2_X1 U15933 ( .A(keyinput10), .B(n14872), .ZN(n14090) );
  XNOR2_X1 U15934 ( .A(keyinput51), .B(n15055), .ZN(n14089) );
  OR4_X1 U15935 ( .A1(n14092), .A2(n14091), .A3(n14090), .A4(n14089), .ZN(
        n14110) );
  AOI22_X1 U15936 ( .A1(n14094), .A2(keyinput41), .B1(n14273), .B2(keyinput2), 
        .ZN(n14093) );
  OAI221_X1 U15937 ( .B1(n14094), .B2(keyinput41), .C1(n14273), .C2(keyinput2), 
        .A(n14093), .ZN(n14109) );
  XOR2_X1 U15938 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput19), .Z(n14098) );
  XOR2_X1 U15939 ( .A(P1_REG0_REG_29__SCAN_IN), .B(keyinput13), .Z(n14097) );
  XNOR2_X1 U15940 ( .A(n14750), .B(keyinput31), .ZN(n14096) );
  XNOR2_X1 U15941 ( .A(n14183), .B(keyinput4), .ZN(n14095) );
  NOR4_X1 U15942 ( .A1(n14098), .A2(n14097), .A3(n14096), .A4(n14095), .ZN(
        n14102) );
  XOR2_X1 U15943 ( .A(n10120), .B(keyinput22), .Z(n14101) );
  XNOR2_X1 U15944 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput29), .ZN(n14100) );
  XNOR2_X1 U15945 ( .A(n14284), .B(keyinput18), .ZN(n14099) );
  NAND4_X1 U15946 ( .A1(n14102), .A2(n14101), .A3(n14100), .A4(n14099), .ZN(
        n14108) );
  XNOR2_X1 U15947 ( .A(P2_IR_REG_3__SCAN_IN), .B(keyinput5), .ZN(n14106) );
  XNOR2_X1 U15948 ( .A(P3_IR_REG_4__SCAN_IN), .B(keyinput20), .ZN(n14105) );
  XNOR2_X1 U15949 ( .A(P2_REG2_REG_28__SCAN_IN), .B(keyinput46), .ZN(n14104)
         );
  XNOR2_X1 U15950 ( .A(P3_IR_REG_22__SCAN_IN), .B(keyinput57), .ZN(n14103) );
  NAND4_X1 U15951 ( .A1(n14106), .A2(n14105), .A3(n14104), .A4(n14103), .ZN(
        n14107) );
  OR4_X1 U15952 ( .A1(n14110), .A2(n14109), .A3(n14108), .A4(n14107), .ZN(
        n14180) );
  AOI22_X1 U15953 ( .A1(n14112), .A2(keyinput49), .B1(keyinput55), .B2(n14202), 
        .ZN(n14111) );
  OAI221_X1 U15954 ( .B1(n14112), .B2(keyinput49), .C1(n14202), .C2(keyinput55), .A(n14111), .ZN(n14121) );
  INV_X1 U15955 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n14114) );
  AOI22_X1 U15956 ( .A1(n14114), .A2(keyinput15), .B1(P3_U3151), .B2(
        keyinput38), .ZN(n14113) );
  OAI221_X1 U15957 ( .B1(n14114), .B2(keyinput15), .C1(P3_U3151), .C2(
        keyinput38), .A(n14113), .ZN(n14120) );
  XNOR2_X1 U15958 ( .A(P3_REG3_REG_22__SCAN_IN), .B(keyinput54), .ZN(n14118)
         );
  XNOR2_X1 U15959 ( .A(P3_IR_REG_21__SCAN_IN), .B(keyinput32), .ZN(n14117) );
  XNOR2_X1 U15960 ( .A(P2_REG1_REG_21__SCAN_IN), .B(keyinput36), .ZN(n14116)
         );
  XNOR2_X1 U15961 ( .A(P2_IR_REG_15__SCAN_IN), .B(keyinput63), .ZN(n14115) );
  NAND4_X1 U15962 ( .A1(n14118), .A2(n14117), .A3(n14116), .A4(n14115), .ZN(
        n14119) );
  NOR3_X1 U15963 ( .A1(n14121), .A2(n14120), .A3(n14119), .ZN(n14160) );
  AOI22_X1 U15964 ( .A1(n14124), .A2(keyinput35), .B1(n14123), .B2(keyinput39), 
        .ZN(n14122) );
  OAI221_X1 U15965 ( .B1(n14124), .B2(keyinput35), .C1(n14123), .C2(keyinput39), .A(n14122), .ZN(n14133) );
  AOI22_X1 U15966 ( .A1(n15149), .A2(keyinput45), .B1(n14126), .B2(keyinput60), 
        .ZN(n14125) );
  OAI221_X1 U15967 ( .B1(n15149), .B2(keyinput45), .C1(n14126), .C2(keyinput60), .A(n14125), .ZN(n14132) );
  AOI22_X1 U15968 ( .A1(n14128), .A2(keyinput7), .B1(keyinput8), .B2(n14365), 
        .ZN(n14127) );
  OAI221_X1 U15969 ( .B1(n14128), .B2(keyinput7), .C1(n14365), .C2(keyinput8), 
        .A(n14127), .ZN(n14131) );
  AOI22_X1 U15970 ( .A1(n14195), .A2(keyinput62), .B1(n14196), .B2(keyinput24), 
        .ZN(n14129) );
  OAI221_X1 U15971 ( .B1(n14195), .B2(keyinput62), .C1(n14196), .C2(keyinput24), .A(n14129), .ZN(n14130) );
  NOR4_X1 U15972 ( .A1(n14133), .A2(n14132), .A3(n14131), .A4(n14130), .ZN(
        n14159) );
  INV_X1 U15973 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n14135) );
  INV_X1 U15974 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n14649) );
  AOI22_X1 U15975 ( .A1(n14135), .A2(keyinput6), .B1(keyinput1), .B2(n14649), 
        .ZN(n14134) );
  OAI221_X1 U15976 ( .B1(n14135), .B2(keyinput6), .C1(n14649), .C2(keyinput1), 
        .A(n14134), .ZN(n14143) );
  INV_X1 U15977 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n14871) );
  AOI22_X1 U15978 ( .A1(n9332), .A2(keyinput59), .B1(n14871), .B2(keyinput23), 
        .ZN(n14136) );
  OAI221_X1 U15979 ( .B1(n9332), .B2(keyinput59), .C1(n14871), .C2(keyinput23), 
        .A(n14136), .ZN(n14142) );
  XNOR2_X1 U15980 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(keyinput34), .ZN(n14139)
         );
  XNOR2_X1 U15981 ( .A(P3_IR_REG_29__SCAN_IN), .B(keyinput26), .ZN(n14138) );
  XNOR2_X1 U15982 ( .A(SI_2_), .B(keyinput25), .ZN(n14137) );
  NAND3_X1 U15983 ( .A1(n14139), .A2(n14138), .A3(n14137), .ZN(n14141) );
  XNOR2_X1 U15984 ( .A(n14186), .B(keyinput53), .ZN(n14140) );
  NOR4_X1 U15985 ( .A1(n14143), .A2(n14142), .A3(n14141), .A4(n14140), .ZN(
        n14158) );
  AOI22_X1 U15986 ( .A1(n14146), .A2(keyinput37), .B1(keyinput47), .B2(n14145), 
        .ZN(n14144) );
  OAI221_X1 U15987 ( .B1(n14146), .B2(keyinput37), .C1(n14145), .C2(keyinput47), .A(n14144), .ZN(n14156) );
  AOI22_X1 U15988 ( .A1(n14181), .A2(keyinput44), .B1(keyinput12), .B2(n14148), 
        .ZN(n14147) );
  OAI221_X1 U15989 ( .B1(n14181), .B2(keyinput44), .C1(n14148), .C2(keyinput12), .A(n14147), .ZN(n14155) );
  XOR2_X1 U15990 ( .A(n13200), .B(keyinput3), .Z(n14151) );
  XNOR2_X1 U15991 ( .A(P1_REG3_REG_8__SCAN_IN), .B(keyinput42), .ZN(n14150) );
  XNOR2_X1 U15992 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput58), .ZN(n14149) );
  NAND3_X1 U15993 ( .A1(n14151), .A2(n14150), .A3(n14149), .ZN(n14154) );
  XNOR2_X1 U15994 ( .A(n14152), .B(keyinput33), .ZN(n14153) );
  NOR4_X1 U15995 ( .A1(n14156), .A2(n14155), .A3(n14154), .A4(n14153), .ZN(
        n14157) );
  NAND4_X1 U15996 ( .A1(n14160), .A2(n14159), .A3(n14158), .A4(n14157), .ZN(
        n14179) );
  AOI22_X1 U15997 ( .A1(n14287), .A2(keyinput30), .B1(n15036), .B2(keyinput40), 
        .ZN(n14161) );
  OAI221_X1 U15998 ( .B1(n14287), .B2(keyinput30), .C1(n15036), .C2(keyinput40), .A(n14161), .ZN(n14168) );
  AOI22_X1 U15999 ( .A1(n14200), .A2(keyinput52), .B1(keyinput11), .B2(n14163), 
        .ZN(n14162) );
  OAI221_X1 U16000 ( .B1(n14200), .B2(keyinput52), .C1(n14163), .C2(keyinput11), .A(n14162), .ZN(n14167) );
  INV_X1 U16001 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15124) );
  AOI22_X1 U16002 ( .A1(n14206), .A2(keyinput0), .B1(n15124), .B2(keyinput17), 
        .ZN(n14164) );
  OAI221_X1 U16003 ( .B1(n14206), .B2(keyinput0), .C1(n15124), .C2(keyinput17), 
        .A(n14164), .ZN(n14166) );
  INV_X1 U16004 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14464) );
  XNOR2_X1 U16005 ( .A(n14464), .B(keyinput14), .ZN(n14165) );
  NOR4_X1 U16006 ( .A1(n14168), .A2(n14167), .A3(n14166), .A4(n14165), .ZN(
        n14177) );
  INV_X1 U16007 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n14205) );
  AOI22_X1 U16008 ( .A1(n14440), .A2(keyinput43), .B1(keyinput50), .B2(n14205), 
        .ZN(n14169) );
  OAI221_X1 U16009 ( .B1(n14440), .B2(keyinput43), .C1(n14205), .C2(keyinput50), .A(n14169), .ZN(n14172) );
  INV_X1 U16010 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n14648) );
  INV_X1 U16011 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14547) );
  AOI22_X1 U16012 ( .A1(n14648), .A2(keyinput56), .B1(keyinput28), .B2(n14547), 
        .ZN(n14170) );
  OAI221_X1 U16013 ( .B1(n14648), .B2(keyinput56), .C1(n14547), .C2(keyinput28), .A(n14170), .ZN(n14171) );
  NOR2_X1 U16014 ( .A1(n14172), .A2(n14171), .ZN(n14176) );
  XOR2_X1 U16015 ( .A(keyinput16), .B(n14173), .Z(n14175) );
  INV_X1 U16016 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14375) );
  XOR2_X1 U16017 ( .A(keyinput61), .B(n14375), .Z(n14174) );
  NAND4_X1 U16018 ( .A1(n14177), .A2(n14176), .A3(n14175), .A4(n14174), .ZN(
        n14178) );
  NOR3_X1 U16019 ( .A1(n14180), .A2(n14179), .A3(n14178), .ZN(n14216) );
  NAND4_X1 U16020 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), 
        .A3(P1_REG1_REG_20__SCAN_IN), .A4(n14649), .ZN(n14194) );
  NAND4_X1 U16021 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(P1_DATAO_REG_9__SCAN_IN), .A3(n14182), .A4(n14181), .ZN(n14193) );
  NOR4_X1 U16022 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(n14284), .A3(
        P1_REG3_REG_8__SCAN_IN), .A4(n14183), .ZN(n14184) );
  NAND4_X1 U16023 ( .A1(n14185), .A2(P2_ADDR_REG_4__SCAN_IN), .A3(
        P1_ADDR_REG_4__SCAN_IN), .A4(n14184), .ZN(n14192) );
  NOR4_X1 U16024 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_REG1_REG_12__SCAN_IN), 
        .A3(P2_IR_REG_3__SCAN_IN), .A4(n10120), .ZN(n14190) );
  NOR4_X1 U16025 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(SI_24_), .A3(
        P3_ADDR_REG_16__SCAN_IN), .A4(n14375), .ZN(n14189) );
  NOR4_X1 U16026 ( .A1(P3_REG0_REG_31__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), 
        .A3(P2_REG2_REG_21__SCAN_IN), .A4(P3_DATAO_REG_7__SCAN_IN), .ZN(n14188) );
  NOR4_X1 U16027 ( .A1(P3_IR_REG_29__SCAN_IN), .A2(P3_REG2_REG_14__SCAN_IN), 
        .A3(P2_D_REG_14__SCAN_IN), .A4(n14186), .ZN(n14187) );
  NAND4_X1 U16028 ( .A1(n14190), .A2(n14189), .A3(n14188), .A4(n14187), .ZN(
        n14191) );
  NOR4_X1 U16029 ( .A1(n14194), .A2(n14193), .A3(n14192), .A4(n14191), .ZN(
        n14214) );
  NAND4_X1 U16030 ( .A1(P3_STATE_REG_SCAN_IN), .A2(P3_REG3_REG_22__SCAN_IN), 
        .A3(P3_REG2_REG_10__SCAN_IN), .A4(P2_REG2_REG_28__SCAN_IN), .ZN(n14198) );
  NAND4_X1 U16031 ( .A1(P1_REG1_REG_22__SCAN_IN), .A2(n14196), .A3(n14195), 
        .A4(n14365), .ZN(n14197) );
  NOR2_X1 U16032 ( .A1(n14198), .A2(n14197), .ZN(n14203) );
  AND3_X1 U16033 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(n14200), .A3(n14199), .ZN(
        n14201) );
  NAND4_X1 U16034 ( .A1(SI_2_), .A2(n14203), .A3(n14202), .A4(n14201), .ZN(
        n14204) );
  NOR4_X1 U16035 ( .A1(n14204), .A2(n14872), .A3(P2_IR_REG_0__SCAN_IN), .A4(
        P3_DATAO_REG_31__SCAN_IN), .ZN(n14213) );
  NAND4_X1 U16036 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(P2_DATAO_REG_27__SCAN_IN), .A3(P3_REG0_REG_6__SCAN_IN), .A4(n14205), .ZN(n14210) );
  NAND4_X1 U16037 ( .A1(n14206), .A2(n14547), .A3(P2_DATAO_REG_21__SCAN_IN), 
        .A4(P1_REG0_REG_8__SCAN_IN), .ZN(n14209) );
  NAND4_X1 U16038 ( .A1(n14207), .A2(n15149), .A3(P1_DATAO_REG_18__SCAN_IN), 
        .A4(P3_REG3_REG_2__SCAN_IN), .ZN(n14208) );
  NOR3_X1 U16039 ( .A1(n14210), .A2(n14209), .A3(n14208), .ZN(n14212) );
  AND4_X1 U16040 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P2_IR_REG_15__SCAN_IN), .A4(P2_REG1_REG_21__SCAN_IN), .ZN(n14211) );
  NAND4_X1 U16041 ( .A1(n14214), .A2(n14213), .A3(n14212), .A4(n14211), .ZN(
        n14215) );
  XNOR2_X1 U16042 ( .A(n14216), .B(n14215), .ZN(n14217) );
  XNOR2_X1 U16043 ( .A(n14218), .B(n14217), .ZN(P1_U3548) );
  AOI211_X1 U16044 ( .C1(n14669), .C2(n14221), .A(n14220), .B(n14219), .ZN(
        n14223) );
  OAI211_X1 U16045 ( .C1(n14224), .C2(n14525), .A(n14223), .B(n14222), .ZN(
        n14257) );
  MUX2_X1 U16046 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14257), .S(n14745), .Z(
        P1_U3547) );
  NAND2_X1 U16047 ( .A1(n14225), .A2(n14729), .ZN(n14229) );
  NAND4_X1 U16048 ( .A1(n14229), .A2(n14228), .A3(n14227), .A4(n14226), .ZN(
        n14258) );
  MUX2_X1 U16049 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14258), .S(n14745), .Z(
        P1_U3546) );
  NAND3_X1 U16050 ( .A1(n13964), .A2(n14230), .A3(n14729), .ZN(n14234) );
  AOI21_X1 U16051 ( .B1(n14232), .B2(n14669), .A(n14231), .ZN(n14233) );
  OAI211_X1 U16052 ( .C1(n14636), .C2(n14235), .A(n14234), .B(n14233), .ZN(
        n14236) );
  AOI21_X1 U16053 ( .B1(n14708), .B2(n14237), .A(n14236), .ZN(n14238) );
  INV_X1 U16054 ( .A(n14238), .ZN(n14259) );
  MUX2_X1 U16055 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14259), .S(n14745), .Z(
        P1_U3545) );
  AOI21_X1 U16056 ( .B1(n14669), .B2(n14240), .A(n14239), .ZN(n14241) );
  OAI211_X1 U16057 ( .C1(n14525), .C2(n14243), .A(n14242), .B(n14241), .ZN(
        n14261) );
  MUX2_X1 U16058 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14261), .S(n14745), .Z(
        P1_U3544) );
  MUX2_X1 U16059 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14244), .S(n14260), .Z(
        P1_U3527) );
  MUX2_X1 U16060 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14245), .S(n14260), .Z(
        P1_U3526) );
  MUX2_X1 U16061 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14246), .S(n14260), .Z(
        P1_U3525) );
  MUX2_X1 U16062 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14247), .S(n14260), .Z(
        P1_U3524) );
  MUX2_X1 U16063 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14248), .S(n14260), .Z(
        P1_U3523) );
  MUX2_X1 U16064 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14249), .S(n14260), .Z(
        P1_U3522) );
  MUX2_X1 U16065 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14250), .S(n14260), .Z(
        P1_U3521) );
  MUX2_X1 U16066 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14251), .S(n14260), .Z(
        P1_U3520) );
  MUX2_X1 U16067 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14252), .S(n14260), .Z(
        P1_U3519) );
  MUX2_X1 U16068 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14253), .S(n14260), .Z(
        P1_U3518) );
  MUX2_X1 U16069 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14254), .S(n14260), .Z(
        P1_U3517) );
  NAND2_X1 U16070 ( .A1(n14731), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n14255) );
  OAI21_X1 U16071 ( .B1(n14256), .B2(n14731), .A(n14255), .ZN(P1_U3516) );
  MUX2_X1 U16072 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14257), .S(n14260), .Z(
        P1_U3515) );
  MUX2_X1 U16073 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14258), .S(n14260), .Z(
        P1_U3513) );
  MUX2_X1 U16074 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14259), .S(n14260), .Z(
        P1_U3510) );
  MUX2_X1 U16075 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14261), .S(n14260), .Z(
        P1_U3507) );
  NAND3_X1 U16076 ( .A1(n14263), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n14265) );
  OAI22_X1 U16077 ( .A1(n14262), .A2(n14265), .B1(n14264), .B2(n14278), .ZN(
        n14266) );
  AOI21_X1 U16078 ( .B1(n14268), .B2(n14267), .A(n14266), .ZN(n14269) );
  INV_X1 U16079 ( .A(n14269), .ZN(P1_U3324) );
  OAI222_X1 U16080 ( .A1(P1_U3086), .A2(n14270), .B1(n14281), .B2(n14272), 
        .C1(n14271), .C2(n14278), .ZN(P1_U3325) );
  OAI222_X1 U16081 ( .A1(n6588), .A2(P1_U3086), .B1(n14281), .B2(n14274), .C1(
        n14273), .C2(n14278), .ZN(P1_U3328) );
  OAI222_X1 U16082 ( .A1(n14277), .A2(P1_U3086), .B1(n14281), .B2(n14276), 
        .C1(n14275), .C2(n14278), .ZN(P1_U3329) );
  OAI222_X1 U16083 ( .A1(P1_U3086), .A2(n14282), .B1(n14281), .B2(n14280), 
        .C1(n14279), .C2(n14278), .ZN(P1_U3330) );
  MUX2_X1 U16084 ( .A(n9719), .B(n14283), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16085 ( .A(n14285), .B(n14284), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3355) );
  INV_X1 U16086 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n14846) );
  INV_X1 U16087 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14383) );
  NAND2_X1 U16088 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14384), .ZN(n14286) );
  OAI21_X1 U16089 ( .B1(n14384), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n14286), 
        .ZN(n14319) );
  INV_X1 U16090 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n14592) );
  INV_X1 U16091 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14314) );
  XOR2_X1 U16092 ( .A(n14314), .B(P1_ADDR_REG_12__SCAN_IN), .Z(n14367) );
  AND2_X1 U16093 ( .A1(n14988), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n14312) );
  XNOR2_X1 U16094 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(n14309), .ZN(n14357) );
  XOR2_X1 U16095 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(n14307), .Z(n14322) );
  INV_X1 U16096 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14301) );
  NAND2_X1 U16097 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n14287), .ZN(n14296) );
  INV_X1 U16098 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n14288) );
  AOI22_X1 U16099 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n14288), .B1(
        P3_ADDR_REG_4__SCAN_IN), .B2(n14287), .ZN(n14324) );
  XOR2_X1 U16100 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n14291), .Z(n14327) );
  NAND2_X1 U16101 ( .A1(n14330), .A2(n14329), .ZN(n14289) );
  NAND2_X1 U16102 ( .A1(n14327), .A2(n14328), .ZN(n14290) );
  NAND2_X1 U16103 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n14292), .ZN(n14295) );
  NAND2_X1 U16104 ( .A1(n14336), .A2(n14293), .ZN(n14294) );
  NAND2_X1 U16105 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n14297), .ZN(n14299) );
  NAND2_X1 U16106 ( .A1(n14340), .A2(n14341), .ZN(n14298) );
  NAND2_X1 U16107 ( .A1(n14299), .A2(n14298), .ZN(n14348) );
  NAND2_X1 U16108 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n14948), .ZN(n14300) );
  INV_X1 U16109 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n14302) );
  NAND2_X1 U16110 ( .A1(n14303), .A2(n14302), .ZN(n14305) );
  XNOR2_X1 U16111 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n14303), .ZN(n14350) );
  NAND2_X1 U16112 ( .A1(n14350), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n14304) );
  NAND2_X1 U16113 ( .A1(n14305), .A2(n14304), .ZN(n14323) );
  NAND2_X1 U16114 ( .A1(n14322), .A2(n14323), .ZN(n14306) );
  NAND2_X1 U16115 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n14358), .ZN(n14311) );
  NOR2_X1 U16116 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n14358), .ZN(n14310) );
  NAND2_X1 U16117 ( .A1(n14367), .A2(n14366), .ZN(n14313) );
  INV_X1 U16118 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n15006) );
  NAND2_X1 U16119 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n15006), .ZN(n14315) );
  AOI22_X1 U16120 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n14592), .B1(n14320), 
        .B2(n14315), .ZN(n14374) );
  NAND2_X1 U16121 ( .A1(P3_ADDR_REG_14__SCAN_IN), .A2(n14316), .ZN(n14317) );
  INV_X1 U16122 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14372) );
  AOI22_X1 U16123 ( .A1(n14374), .A2(n14317), .B1(P1_ADDR_REG_14__SCAN_IN), 
        .B2(n14372), .ZN(n14378) );
  INV_X1 U16124 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14436) );
  NAND2_X1 U16125 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n14436), .ZN(n14318) );
  INV_X1 U16126 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14377) );
  AOI22_X1 U16127 ( .A1(n14378), .A2(n14318), .B1(P3_ADDR_REG_15__SCAN_IN), 
        .B2(n14377), .ZN(n14386) );
  XNOR2_X1 U16128 ( .A(n14319), .B(n14386), .ZN(n14568) );
  INV_X1 U16129 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14371) );
  XOR2_X1 U16130 ( .A(n15006), .B(P1_ADDR_REG_13__SCAN_IN), .Z(n14321) );
  XNOR2_X1 U16131 ( .A(n14321), .B(n14320), .ZN(n14557) );
  INV_X1 U16132 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14361) );
  XOR2_X1 U16133 ( .A(n14323), .B(n14322), .Z(n14355) );
  XNOR2_X1 U16134 ( .A(n14325), .B(n14324), .ZN(n14326) );
  NAND2_X1 U16135 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14326), .ZN(n14339) );
  XOR2_X1 U16136 ( .A(P2_ADDR_REG_4__SCAN_IN), .B(n14326), .Z(n15168) );
  INV_X1 U16137 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14335) );
  XNOR2_X1 U16138 ( .A(n14328), .B(n14327), .ZN(n14397) );
  NAND2_X1 U16139 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14331), .ZN(n14333) );
  AOI21_X1 U16140 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14910), .A(n14330), .ZN(
        n15171) );
  INV_X1 U16141 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15170) );
  NOR2_X1 U16142 ( .A1(n15171), .A2(n15170), .ZN(n15180) );
  NAND2_X1 U16143 ( .A1(n15180), .A2(n15179), .ZN(n14332) );
  NAND2_X1 U16144 ( .A1(n14333), .A2(n14332), .ZN(n14398) );
  NAND2_X1 U16145 ( .A1(n14397), .A2(n14398), .ZN(n14334) );
  NOR2_X1 U16146 ( .A1(n14397), .A2(n14398), .ZN(n14396) );
  AOI21_X1 U16147 ( .B1(n14335), .B2(n14334), .A(n14396), .ZN(n15175) );
  XOR2_X1 U16148 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n14336), .Z(n15176) );
  NOR2_X1 U16149 ( .A1(n15175), .A2(n15176), .ZN(n14337) );
  INV_X1 U16150 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15177) );
  NAND2_X1 U16151 ( .A1(n15175), .A2(n15176), .ZN(n15174) );
  OAI21_X1 U16152 ( .B1(n14337), .B2(n15177), .A(n15174), .ZN(n15167) );
  NAND2_X1 U16153 ( .A1(n15168), .A2(n15167), .ZN(n14338) );
  NAND2_X1 U16154 ( .A1(n14339), .A2(n14338), .ZN(n14343) );
  XNOR2_X1 U16155 ( .A(n14341), .B(n14340), .ZN(n14342) );
  NOR2_X1 U16156 ( .A1(n14343), .A2(n14342), .ZN(n14345) );
  XNOR2_X1 U16157 ( .A(n14343), .B(n14342), .ZN(n15169) );
  NOR2_X1 U16158 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n15169), .ZN(n14344) );
  NAND2_X1 U16159 ( .A1(n14346), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14349) );
  XNOR2_X1 U16160 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n14948), .ZN(n14347) );
  XOR2_X1 U16161 ( .A(n14348), .B(n14347), .Z(n14400) );
  XOR2_X1 U16162 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n14350), .Z(n15173) );
  NAND2_X1 U16163 ( .A1(n15172), .A2(n15173), .ZN(n14353) );
  NAND2_X1 U16164 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14351), .ZN(n14352) );
  XNOR2_X1 U16165 ( .A(n14355), .B(n14354), .ZN(n14402) );
  XNOR2_X1 U16166 ( .A(n14357), .B(n14356), .ZN(n14404) );
  XNOR2_X1 U16167 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(P3_ADDR_REG_10__SCAN_IN), 
        .ZN(n14359) );
  XOR2_X1 U16168 ( .A(n14359), .B(n14358), .Z(n14408) );
  NAND2_X1 U16169 ( .A1(n14409), .A2(n14408), .ZN(n14360) );
  NOR2_X1 U16170 ( .A1(n14409), .A2(n14408), .ZN(n14407) );
  XNOR2_X1 U16171 ( .A(n14988), .B(P1_ADDR_REG_11__SCAN_IN), .ZN(n14362) );
  XNOR2_X1 U16172 ( .A(n14363), .B(n14362), .ZN(n14553) );
  NAND2_X1 U16173 ( .A1(n14554), .A2(n14553), .ZN(n14364) );
  NOR2_X1 U16174 ( .A1(n14554), .A2(n14553), .ZN(n14552) );
  XNOR2_X1 U16175 ( .A(n14367), .B(n14366), .ZN(n14369) );
  NOR2_X1 U16176 ( .A1(n14368), .A2(n14369), .ZN(n14370) );
  XNOR2_X1 U16177 ( .A(n14372), .B(P1_ADDR_REG_14__SCAN_IN), .ZN(n14373) );
  XNOR2_X1 U16178 ( .A(n14374), .B(n14373), .ZN(n14561) );
  XOR2_X1 U16179 ( .A(n14377), .B(P3_ADDR_REG_15__SCAN_IN), .Z(n14379) );
  XOR2_X1 U16180 ( .A(n14379), .B(n14378), .Z(n14381) );
  NAND2_X1 U16181 ( .A1(n14568), .A2(n14569), .ZN(n14382) );
  NOR2_X1 U16182 ( .A1(n14568), .A2(n14569), .ZN(n14567) );
  INV_X1 U16183 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14388) );
  OR2_X1 U16184 ( .A1(n14384), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n14385) );
  AOI22_X1 U16185 ( .A1(n14386), .A2(n14385), .B1(P1_ADDR_REG_16__SCAN_IN), 
        .B2(n14384), .ZN(n14389) );
  XOR2_X1 U16186 ( .A(n14388), .B(n14389), .Z(n14390) );
  XNOR2_X1 U16187 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14390), .ZN(n14421) );
  NOR2_X1 U16188 ( .A1(n14420), .A2(n14421), .ZN(n14387) );
  NAND2_X1 U16189 ( .A1(n14420), .A2(n14421), .ZN(n14419) );
  NAND2_X1 U16190 ( .A1(n14389), .A2(n14388), .ZN(n14392) );
  NAND2_X1 U16191 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n14390), .ZN(n14391) );
  NAND2_X1 U16192 ( .A1(n14392), .A2(n14391), .ZN(n14426) );
  NOR2_X1 U16193 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n14429), .ZN(n14393) );
  AOI21_X1 U16194 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n14429), .A(n14393), 
        .ZN(n14427) );
  XNOR2_X1 U16195 ( .A(n14426), .B(n14427), .ZN(n14424) );
  XOR2_X1 U16196 ( .A(n14846), .B(n14423), .Z(SUB_1596_U62) );
  AOI21_X1 U16197 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14394) );
  OAI21_X1 U16198 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14394), 
        .ZN(U28) );
  AOI21_X1 U16199 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14395) );
  OAI21_X1 U16200 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14395), 
        .ZN(U29) );
  AOI21_X1 U16201 ( .B1(n14398), .B2(n14397), .A(n14396), .ZN(n14399) );
  XOR2_X1 U16202 ( .A(n14399), .B(P2_ADDR_REG_2__SCAN_IN), .Z(SUB_1596_U61) );
  XOR2_X1 U16203 ( .A(n14401), .B(n14400), .Z(SUB_1596_U57) );
  XNOR2_X1 U16204 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n14402), .ZN(SUB_1596_U55)
         );
  AOI21_X1 U16205 ( .B1(n14405), .B2(n14404), .A(n14403), .ZN(n14406) );
  XOR2_X1 U16206 ( .A(n14406), .B(P2_ADDR_REG_9__SCAN_IN), .Z(SUB_1596_U54) );
  AOI21_X1 U16207 ( .B1(n14409), .B2(n14408), .A(n14407), .ZN(n14410) );
  XOR2_X1 U16208 ( .A(n14410), .B(P2_ADDR_REG_10__SCAN_IN), .Z(SUB_1596_U70)
         );
  INV_X1 U16209 ( .A(n14704), .ZN(n14722) );
  INV_X1 U16210 ( .A(n14411), .ZN(n14416) );
  OAI21_X1 U16211 ( .B1(n14413), .B2(n14726), .A(n14412), .ZN(n14415) );
  AOI211_X1 U16212 ( .C1(n14722), .C2(n14416), .A(n14415), .B(n14414), .ZN(
        n14418) );
  INV_X1 U16213 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14417) );
  AOI22_X1 U16214 ( .A1(n14260), .A2(n14418), .B1(n14417), .B2(n14731), .ZN(
        P1_U3495) );
  AOI22_X1 U16215 ( .A1(n14745), .A2(n14418), .B1(n10525), .B2(n14742), .ZN(
        P1_U3540) );
  OAI21_X1 U16216 ( .B1(n14421), .B2(n14420), .A(n14419), .ZN(n14422) );
  XOR2_X1 U16217 ( .A(n14422), .B(n11423), .Z(SUB_1596_U63) );
  NAND2_X1 U16218 ( .A1(n14427), .A2(n14426), .ZN(n14428) );
  OAI21_X1 U16219 ( .B1(n14429), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n14428), 
        .ZN(n14430) );
  XNOR2_X1 U16220 ( .A(n14430), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n14432) );
  XNOR2_X1 U16221 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n14431) );
  AOI21_X1 U16222 ( .B1(n14435), .B2(n14434), .A(n14433), .ZN(n14450) );
  OAI22_X1 U16223 ( .A1(n15008), .A2(n14437), .B1(n14436), .B2(n15005), .ZN(
        n14447) );
  AOI21_X1 U16224 ( .B1(n14440), .B2(n14439), .A(n14438), .ZN(n14445) );
  AOI21_X1 U16225 ( .B1(n14443), .B2(n14442), .A(n14441), .ZN(n14444) );
  OAI22_X1 U16226 ( .A1(n14445), .A2(n15017), .B1(n14444), .B2(n15015), .ZN(
        n14446) );
  NOR3_X1 U16227 ( .A1(n14448), .A2(n14447), .A3(n14446), .ZN(n14449) );
  OAI21_X1 U16228 ( .B1(n14450), .B2(n15023), .A(n14449), .ZN(P3_U3197) );
  XNOR2_X1 U16229 ( .A(n14451), .B(n14455), .ZN(n14453) );
  AOI222_X1 U16230 ( .A1(n15074), .A2(n14453), .B1(n14452), .B2(n15079), .C1(
        n15039), .C2(n15076), .ZN(n14465) );
  AOI22_X1 U16231 ( .A1(n15071), .A2(P3_REG2_REG_11__SCAN_IN), .B1(n15090), 
        .B2(n14454), .ZN(n14460) );
  XNOR2_X1 U16232 ( .A(n14456), .B(n14455), .ZN(n14468) );
  NOR2_X1 U16233 ( .A1(n14457), .A2(n15130), .ZN(n14467) );
  AOI22_X1 U16234 ( .A1(n14468), .A2(n14458), .B1(n15048), .B2(n14467), .ZN(
        n14459) );
  OAI211_X1 U16235 ( .C1(n15071), .C2(n14465), .A(n14460), .B(n14459), .ZN(
        P3_U3222) );
  AOI211_X1 U16236 ( .C1(n14463), .C2(n15099), .A(n14462), .B(n14461), .ZN(
        n14470) );
  AOI22_X1 U16237 ( .A1(n15166), .A2(n14470), .B1(n14464), .B2(n15163), .ZN(
        P3_U3471) );
  INV_X1 U16238 ( .A(n14465), .ZN(n14466) );
  AOI211_X1 U16239 ( .C1(n14468), .C2(n15099), .A(n14467), .B(n14466), .ZN(
        n14472) );
  AOI22_X1 U16240 ( .A1(n15166), .A2(n14472), .B1(n9067), .B2(n15163), .ZN(
        P3_U3470) );
  INV_X1 U16241 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14469) );
  AOI22_X1 U16242 ( .A1(n15146), .A2(n14470), .B1(n14469), .B2(n15144), .ZN(
        P3_U3426) );
  INV_X1 U16243 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14471) );
  AOI22_X1 U16244 ( .A1(n15146), .A2(n14472), .B1(n14471), .B2(n15144), .ZN(
        P3_U3423) );
  XNOR2_X1 U16245 ( .A(n14473), .B(n14481), .ZN(n14476) );
  AOI21_X1 U16246 ( .B1(n14476), .B2(n14475), .A(n14474), .ZN(n14497) );
  AOI222_X1 U16247 ( .A1(n14480), .A2(n14479), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(n14478), .C1(n14849), .C2(n14477), .ZN(n14489) );
  XOR2_X1 U16248 ( .A(n14482), .B(n14481), .Z(n14499) );
  INV_X1 U16249 ( .A(n14483), .ZN(n14486) );
  INV_X1 U16250 ( .A(n14484), .ZN(n14485) );
  OAI211_X1 U16251 ( .C1(n6771), .C2(n14486), .A(n14485), .B(n13083), .ZN(
        n14496) );
  INV_X1 U16252 ( .A(n14496), .ZN(n14487) );
  AOI22_X1 U16253 ( .A1(n14499), .A2(n14856), .B1(n14847), .B2(n14487), .ZN(
        n14488) );
  OAI211_X1 U16254 ( .C1(n14478), .C2(n14497), .A(n14489), .B(n14488), .ZN(
        P2_U3251) );
  OAI211_X1 U16255 ( .C1(n14493), .C2(n13305), .A(n14492), .B(n14491), .ZN(
        n14494) );
  AOI21_X1 U16256 ( .B1(n14511), .B2(n14495), .A(n14494), .ZN(n14514) );
  AOI22_X1 U16257 ( .A1(n14903), .A2(n14514), .B1(n11402), .B2(n14900), .ZN(
        P2_U3514) );
  OAI211_X1 U16258 ( .C1(n6771), .C2(n13305), .A(n14497), .B(n14496), .ZN(
        n14498) );
  AOI21_X1 U16259 ( .B1(n14499), .B2(n14511), .A(n14498), .ZN(n14516) );
  AOI22_X1 U16260 ( .A1(n14903), .A2(n14516), .B1(n14500), .B2(n14900), .ZN(
        P2_U3513) );
  OAI211_X1 U16261 ( .C1(n10019), .C2(n13305), .A(n14502), .B(n14501), .ZN(
        n14503) );
  AOI21_X1 U16262 ( .B1(n14504), .B2(n14511), .A(n14503), .ZN(n14518) );
  AOI22_X1 U16263 ( .A1(n14903), .A2(n14518), .B1(n14505), .B2(n14900), .ZN(
        P2_U3512) );
  OAI21_X1 U16264 ( .B1(n14507), .B2(n13305), .A(n14506), .ZN(n14509) );
  AOI211_X1 U16265 ( .C1(n14511), .C2(n14510), .A(n14509), .B(n14508), .ZN(
        n14520) );
  AOI22_X1 U16266 ( .A1(n14903), .A2(n14520), .B1(n14512), .B2(n14900), .ZN(
        P2_U3511) );
  INV_X1 U16267 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n14513) );
  AOI22_X1 U16268 ( .A1(n14898), .A2(n14514), .B1(n14513), .B2(n14896), .ZN(
        P2_U3475) );
  INV_X1 U16269 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14515) );
  AOI22_X1 U16270 ( .A1(n14898), .A2(n14516), .B1(n14515), .B2(n14896), .ZN(
        P2_U3472) );
  INV_X1 U16271 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n14517) );
  AOI22_X1 U16272 ( .A1(n14898), .A2(n14518), .B1(n14517), .B2(n14896), .ZN(
        P2_U3469) );
  INV_X1 U16273 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14519) );
  AOI22_X1 U16274 ( .A1(n14898), .A2(n14520), .B1(n14519), .B2(n14896), .ZN(
        P2_U3466) );
  AOI21_X1 U16275 ( .B1(n14669), .B2(n14522), .A(n14521), .ZN(n14523) );
  OAI211_X1 U16276 ( .C1(n14526), .C2(n14525), .A(n14524), .B(n14523), .ZN(
        n14527) );
  INV_X1 U16277 ( .A(n14527), .ZN(n14546) );
  AOI22_X1 U16278 ( .A1(n14745), .A2(n14546), .B1(n9452), .B2(n14742), .ZN(
        P1_U3543) );
  NAND2_X1 U16279 ( .A1(n14528), .A2(n14669), .ZN(n14529) );
  AND2_X1 U16280 ( .A1(n14530), .A2(n14529), .ZN(n14533) );
  NAND3_X1 U16281 ( .A1(n6539), .A2(n14531), .A3(n14729), .ZN(n14532) );
  AOI22_X1 U16282 ( .A1(n14745), .A2(n14548), .B1(n9437), .B2(n14742), .ZN(
        P1_U3542) );
  OAI21_X1 U16283 ( .B1(n14536), .B2(n14726), .A(n14535), .ZN(n14538) );
  AOI211_X1 U16284 ( .C1(n14539), .C2(n14729), .A(n14538), .B(n14537), .ZN(
        n14550) );
  AOI22_X1 U16285 ( .A1(n14745), .A2(n14550), .B1(n10924), .B2(n14742), .ZN(
        P1_U3541) );
  OAI21_X1 U16286 ( .B1(n14541), .B2(n14726), .A(n14540), .ZN(n14543) );
  AOI211_X1 U16287 ( .C1(n14544), .C2(n14729), .A(n14543), .B(n14542), .ZN(
        n14551) );
  AOI22_X1 U16288 ( .A1(n14745), .A2(n14551), .B1(n9382), .B2(n14742), .ZN(
        P1_U3539) );
  INV_X1 U16289 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n14545) );
  AOI22_X1 U16290 ( .A1(n14260), .A2(n14546), .B1(n14545), .B2(n14731), .ZN(
        P1_U3504) );
  AOI22_X1 U16291 ( .A1(n14260), .A2(n14548), .B1(n14547), .B2(n14731), .ZN(
        P1_U3501) );
  INV_X1 U16292 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14549) );
  AOI22_X1 U16293 ( .A1(n14260), .A2(n14550), .B1(n14549), .B2(n14731), .ZN(
        P1_U3498) );
  AOI22_X1 U16294 ( .A1(n14260), .A2(n14551), .B1(n9381), .B2(n14731), .ZN(
        P1_U3492) );
  AOI21_X1 U16295 ( .B1(n14554), .B2(n14553), .A(n14552), .ZN(n14555) );
  XOR2_X1 U16296 ( .A(n14555), .B(P2_ADDR_REG_11__SCAN_IN), .Z(SUB_1596_U69)
         );
  XNOR2_X1 U16297 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n14556), .ZN(SUB_1596_U68)
         );
  AOI21_X1 U16298 ( .B1(n14558), .B2(n14557), .A(n6551), .ZN(n14559) );
  XOR2_X1 U16299 ( .A(n14559), .B(P2_ADDR_REG_13__SCAN_IN), .Z(SUB_1596_U67)
         );
  AOI21_X1 U16300 ( .B1(n14562), .B2(n14561), .A(n14560), .ZN(n14563) );
  XOR2_X1 U16301 ( .A(n14563), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  NOR2_X1 U16302 ( .A1(n14565), .A2(n14564), .ZN(n14566) );
  XOR2_X1 U16303 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n14566), .Z(SUB_1596_U65)
         );
  AOI21_X1 U16304 ( .B1(n14569), .B2(n14568), .A(n14567), .ZN(n14570) );
  XOR2_X1 U16305 ( .A(n14570), .B(P2_ADDR_REG_16__SCAN_IN), .Z(SUB_1596_U64)
         );
  INV_X1 U16306 ( .A(n14571), .ZN(n14576) );
  NAND3_X1 U16307 ( .A1(n14574), .A2(n14573), .A3(n14572), .ZN(n14575) );
  NAND3_X1 U16308 ( .A1(n14597), .A2(n14576), .A3(n14575), .ZN(n14588) );
  AND2_X1 U16309 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n14577) );
  AOI21_X1 U16310 ( .B1(n14578), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n14577), .ZN(
        n14587) );
  NAND2_X1 U16311 ( .A1(n14595), .A2(n14579), .ZN(n14586) );
  MUX2_X1 U16312 ( .A(n10344), .B(P1_REG2_REG_4__SCAN_IN), .S(n14579), .Z(
        n14580) );
  NAND3_X1 U16313 ( .A1(n14582), .A2(n14581), .A3(n14580), .ZN(n14583) );
  NAND3_X1 U16314 ( .A1(n14602), .A2(n14584), .A3(n14583), .ZN(n14585) );
  AND4_X1 U16315 ( .A1(n14588), .A2(n14587), .A3(n14586), .A4(n14585), .ZN(
        n14590) );
  NAND2_X1 U16316 ( .A1(n14590), .A2(n14589), .ZN(P1_U3247) );
  OAI21_X1 U16317 ( .B1(n14593), .B2(n14592), .A(n14591), .ZN(n14594) );
  AOI21_X1 U16318 ( .B1(n14596), .B2(n14595), .A(n14594), .ZN(n14607) );
  OAI211_X1 U16319 ( .C1(n14600), .C2(n14599), .A(n14598), .B(n14597), .ZN(
        n14606) );
  OAI211_X1 U16320 ( .C1(n14604), .C2(n14603), .A(n14602), .B(n14601), .ZN(
        n14605) );
  NAND3_X1 U16321 ( .A1(n14607), .A2(n14606), .A3(n14605), .ZN(P1_U3256) );
  OAI21_X1 U16322 ( .B1(n14610), .B2(n14609), .A(n14608), .ZN(n14697) );
  XNOR2_X1 U16323 ( .A(n14612), .B(n14611), .ZN(n14613) );
  AND2_X1 U16324 ( .A1(n14613), .A2(n14708), .ZN(n14695) );
  AOI211_X1 U16325 ( .C1(n14675), .C2(n14697), .A(n14691), .B(n14695), .ZN(
        n14627) );
  INV_X1 U16326 ( .A(n14614), .ZN(n14615) );
  AOI222_X1 U16327 ( .A1(n14616), .A2(n14634), .B1(P1_REG2_REG_6__SCAN_IN), 
        .B2(n14647), .C1(n14635), .C2(n14615), .ZN(n14626) );
  NAND2_X1 U16328 ( .A1(n14617), .A2(n14616), .ZN(n14619) );
  NAND2_X1 U16329 ( .A1(n14619), .A2(n14618), .ZN(n14621) );
  OR2_X1 U16330 ( .A1(n14621), .A2(n14620), .ZN(n14694) );
  INV_X1 U16331 ( .A(n14694), .ZN(n14622) );
  AOI22_X1 U16332 ( .A1(n14697), .A2(n14624), .B1(n14623), .B2(n14622), .ZN(
        n14625) );
  OAI211_X1 U16333 ( .C1(n14647), .C2(n14627), .A(n14626), .B(n14625), .ZN(
        P1_U3287) );
  XNOR2_X1 U16334 ( .A(n14630), .B(n14628), .ZN(n14633) );
  XNOR2_X1 U16335 ( .A(n14630), .B(n14629), .ZN(n14659) );
  NOR2_X1 U16336 ( .A1(n14659), .A2(n14703), .ZN(n14631) );
  AOI211_X1 U16337 ( .C1(n14708), .C2(n14633), .A(n14632), .B(n14631), .ZN(
        n14662) );
  AOI222_X1 U16338 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(n14647), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n14635), .C1(n14638), .C2(n14634), .ZN(
        n14646) );
  AOI21_X1 U16339 ( .B1(n14638), .B2(n14637), .A(n14636), .ZN(n14640) );
  NAND2_X1 U16340 ( .A1(n14640), .A2(n14639), .ZN(n14660) );
  OR2_X1 U16341 ( .A1(n14641), .A2(n14659), .ZN(n14642) );
  OAI21_X1 U16342 ( .B1(n14643), .B2(n14660), .A(n14642), .ZN(n14644) );
  INV_X1 U16343 ( .A(n14644), .ZN(n14645) );
  OAI211_X1 U16344 ( .C1(n14647), .C2(n14662), .A(n14646), .B(n14645), .ZN(
        P1_U3291) );
  AND2_X1 U16345 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14651), .ZN(P1_U3294) );
  AND2_X1 U16346 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14651), .ZN(P1_U3295) );
  AND2_X1 U16347 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14651), .ZN(P1_U3296) );
  AND2_X1 U16348 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14651), .ZN(P1_U3297) );
  AND2_X1 U16349 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14651), .ZN(P1_U3298) );
  AND2_X1 U16350 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14651), .ZN(P1_U3299) );
  AND2_X1 U16351 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14651), .ZN(P1_U3300) );
  AND2_X1 U16352 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14651), .ZN(P1_U3301) );
  AND2_X1 U16353 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14651), .ZN(P1_U3302) );
  AND2_X1 U16354 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14651), .ZN(P1_U3303) );
  AND2_X1 U16355 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14651), .ZN(P1_U3304) );
  AND2_X1 U16356 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14651), .ZN(P1_U3305) );
  AND2_X1 U16357 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14651), .ZN(P1_U3306) );
  AND2_X1 U16358 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14651), .ZN(P1_U3307) );
  AND2_X1 U16359 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14651), .ZN(P1_U3308) );
  AND2_X1 U16360 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14651), .ZN(P1_U3309) );
  AND2_X1 U16361 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14651), .ZN(P1_U3310) );
  AND2_X1 U16362 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14651), .ZN(P1_U3311) );
  AND2_X1 U16363 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14651), .ZN(P1_U3312) );
  INV_X1 U16364 ( .A(n14651), .ZN(n14650) );
  NOR2_X1 U16365 ( .A1(n14650), .A2(n14648), .ZN(P1_U3313) );
  AND2_X1 U16366 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14651), .ZN(P1_U3314) );
  AND2_X1 U16367 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14651), .ZN(P1_U3315) );
  AND2_X1 U16368 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14651), .ZN(P1_U3316) );
  AND2_X1 U16369 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14651), .ZN(P1_U3317) );
  AND2_X1 U16370 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14651), .ZN(P1_U3318) );
  AND2_X1 U16371 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14651), .ZN(P1_U3319) );
  AND2_X1 U16372 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14651), .ZN(P1_U3320) );
  AND2_X1 U16373 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14651), .ZN(P1_U3321) );
  NOR2_X1 U16374 ( .A1(n14650), .A2(n14649), .ZN(P1_U3322) );
  AND2_X1 U16375 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14651), .ZN(P1_U3323) );
  INV_X1 U16376 ( .A(n14652), .ZN(n14653) );
  OAI21_X1 U16377 ( .B1(n10631), .B2(n14726), .A(n14653), .ZN(n14656) );
  INV_X1 U16378 ( .A(n14654), .ZN(n14655) );
  AOI211_X1 U16379 ( .C1(n14722), .C2(n14657), .A(n14656), .B(n14655), .ZN(
        n14732) );
  INV_X1 U16380 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14658) );
  AOI22_X1 U16381 ( .A1(n14260), .A2(n14732), .B1(n14658), .B2(n14731), .ZN(
        P1_U3462) );
  INV_X1 U16382 ( .A(n14659), .ZN(n14665) );
  OAI21_X1 U16383 ( .B1(n14661), .B2(n14726), .A(n14660), .ZN(n14664) );
  INV_X1 U16384 ( .A(n14662), .ZN(n14663) );
  AOI211_X1 U16385 ( .C1(n14722), .C2(n14665), .A(n14664), .B(n14663), .ZN(
        n14733) );
  INV_X1 U16386 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n14666) );
  AOI22_X1 U16387 ( .A1(n14260), .A2(n14733), .B1(n14666), .B2(n14731), .ZN(
        P1_U3465) );
  INV_X1 U16388 ( .A(n14672), .ZN(n14674) );
  AOI21_X1 U16389 ( .B1(n14669), .B2(n14668), .A(n14667), .ZN(n14671) );
  OAI211_X1 U16390 ( .C1(n14704), .C2(n14672), .A(n14671), .B(n14670), .ZN(
        n14673) );
  AOI21_X1 U16391 ( .B1(n14675), .B2(n14674), .A(n14673), .ZN(n14734) );
  INV_X1 U16392 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n14676) );
  AOI22_X1 U16393 ( .A1(n14260), .A2(n14734), .B1(n14676), .B2(n14731), .ZN(
        P1_U3468) );
  NAND3_X1 U16394 ( .A1(n11275), .A2(n14677), .A3(n14729), .ZN(n14679) );
  OAI211_X1 U16395 ( .C1(n14680), .C2(n14726), .A(n14679), .B(n14678), .ZN(
        n14682) );
  NOR2_X1 U16396 ( .A1(n14682), .A2(n14681), .ZN(n14736) );
  INV_X1 U16397 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14683) );
  AOI22_X1 U16398 ( .A1(n14260), .A2(n14736), .B1(n14683), .B2(n14731), .ZN(
        P1_U3471) );
  INV_X1 U16399 ( .A(n14684), .ZN(n14690) );
  OR4_X1 U16400 ( .A1(n14688), .A2(n14687), .A3(n14686), .A4(n14685), .ZN(
        n14689) );
  AOI21_X1 U16401 ( .B1(n14690), .B2(n14729), .A(n14689), .ZN(n14737) );
  AOI22_X1 U16402 ( .A1(n14260), .A2(n14737), .B1(n9278), .B2(n14731), .ZN(
        P1_U3474) );
  NOR2_X1 U16403 ( .A1(n14692), .A2(n14691), .ZN(n14693) );
  NAND2_X1 U16404 ( .A1(n14694), .A2(n14693), .ZN(n14696) );
  AOI211_X1 U16405 ( .C1(n14729), .C2(n14697), .A(n14696), .B(n14695), .ZN(
        n14738) );
  INV_X1 U16406 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14698) );
  AOI22_X1 U16407 ( .A1(n14260), .A2(n14738), .B1(n14698), .B2(n14731), .ZN(
        P1_U3477) );
  OAI211_X1 U16408 ( .C1(n14701), .C2(n14726), .A(n14700), .B(n14699), .ZN(
        n14706) );
  AOI21_X1 U16409 ( .B1(n14704), .B2(n14703), .A(n14702), .ZN(n14705) );
  AOI211_X1 U16410 ( .C1(n14708), .C2(n14707), .A(n14706), .B(n14705), .ZN(
        n14739) );
  INV_X1 U16411 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n14709) );
  AOI22_X1 U16412 ( .A1(n14260), .A2(n14739), .B1(n14709), .B2(n14731), .ZN(
        P1_U3480) );
  INV_X1 U16413 ( .A(n14710), .ZN(n14711) );
  NAND4_X1 U16414 ( .A1(n14714), .A2(n14713), .A3(n14712), .A4(n14711), .ZN(
        n14715) );
  AOI21_X1 U16415 ( .B1(n14716), .B2(n14729), .A(n14715), .ZN(n14740) );
  AOI22_X1 U16416 ( .A1(n14260), .A2(n14740), .B1(n9332), .B2(n14731), .ZN(
        P1_U3483) );
  INV_X1 U16417 ( .A(n14717), .ZN(n14721) );
  OAI21_X1 U16418 ( .B1(n6828), .B2(n14726), .A(n14718), .ZN(n14720) );
  AOI211_X1 U16419 ( .C1(n14722), .C2(n14721), .A(n14720), .B(n14719), .ZN(
        n14741) );
  INV_X1 U16420 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14723) );
  AOI22_X1 U16421 ( .A1(n14260), .A2(n14741), .B1(n14723), .B2(n14731), .ZN(
        P1_U3486) );
  OAI211_X1 U16422 ( .C1(n6827), .C2(n14726), .A(n14725), .B(n14724), .ZN(
        n14728) );
  AOI211_X1 U16423 ( .C1(n14730), .C2(n14729), .A(n14728), .B(n14727), .ZN(
        n14744) );
  AOI22_X1 U16424 ( .A1(n14260), .A2(n14744), .B1(n14206), .B2(n14731), .ZN(
        P1_U3489) );
  AOI22_X1 U16425 ( .A1(n14745), .A2(n14732), .B1(n10324), .B2(n14742), .ZN(
        P1_U3529) );
  AOI22_X1 U16426 ( .A1(n14745), .A2(n14733), .B1(n10323), .B2(n14742), .ZN(
        P1_U3530) );
  AOI22_X1 U16427 ( .A1(n14745), .A2(n14734), .B1(n10328), .B2(n14742), .ZN(
        P1_U3531) );
  AOI22_X1 U16428 ( .A1(n14745), .A2(n14736), .B1(n14735), .B2(n14742), .ZN(
        P1_U3532) );
  AOI22_X1 U16429 ( .A1(n14745), .A2(n14737), .B1(n6612), .B2(n14742), .ZN(
        P1_U3533) );
  AOI22_X1 U16430 ( .A1(n14745), .A2(n14738), .B1(n9305), .B2(n14742), .ZN(
        P1_U3534) );
  AOI22_X1 U16431 ( .A1(n14745), .A2(n14739), .B1(n10329), .B2(n14742), .ZN(
        P1_U3535) );
  AOI22_X1 U16432 ( .A1(n14745), .A2(n14740), .B1(n10331), .B2(n14742), .ZN(
        P1_U3536) );
  AOI22_X1 U16433 ( .A1(n14745), .A2(n14741), .B1(n9349), .B2(n14742), .ZN(
        P1_U3537) );
  AOI22_X1 U16434 ( .A1(n14745), .A2(n14744), .B1(n14743), .B2(n14742), .ZN(
        P1_U3538) );
  NOR2_X1 U16435 ( .A1(n14818), .A2(P2_U3947), .ZN(P2_U3087) );
  OR2_X1 U16436 ( .A1(n14746), .A2(P2_U3088), .ZN(n14776) );
  NAND2_X1 U16437 ( .A1(P2_U3088), .A2(n14747), .ZN(n14748) );
  OAI211_X1 U16438 ( .C1(n14749), .C2(P2_U3088), .A(n14776), .B(n14748), .ZN(
        n14760) );
  NOR2_X1 U16439 ( .A1(n14750), .A2(n7405), .ZN(n14753) );
  OAI211_X1 U16440 ( .C1(n14753), .C2(n14752), .A(n14820), .B(n14751), .ZN(
        n14759) );
  OAI211_X1 U16441 ( .C1(n14756), .C2(n14755), .A(n14825), .B(n14754), .ZN(
        n14758) );
  NAND2_X1 U16442 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14818), .ZN(n14757) );
  NAND4_X1 U16443 ( .A1(n14760), .A2(n14759), .A3(n14758), .A4(n14757), .ZN(
        P2_U3215) );
  NAND2_X1 U16444 ( .A1(P2_U3088), .A2(n14761), .ZN(n14762) );
  OAI211_X1 U16445 ( .C1(n14763), .C2(P2_U3088), .A(n14776), .B(n14762), .ZN(
        n14773) );
  OAI211_X1 U16446 ( .C1(n14766), .C2(n14765), .A(n14820), .B(n14764), .ZN(
        n14772) );
  NAND2_X1 U16447 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14818), .ZN(n14771) );
  OAI211_X1 U16448 ( .C1(n14769), .C2(n14768), .A(n14825), .B(n14767), .ZN(
        n14770) );
  NAND4_X1 U16449 ( .A1(n14773), .A2(n14772), .A3(n14771), .A4(n14770), .ZN(
        P2_U3218) );
  NAND2_X1 U16450 ( .A1(n14774), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14775) );
  OAI211_X1 U16451 ( .C1(P2_STATE_REG_SCAN_IN), .C2(P2_REG3_REG_6__SCAN_IN), 
        .A(n14776), .B(n14775), .ZN(n14787) );
  OAI211_X1 U16452 ( .C1(n14779), .C2(n14778), .A(n14825), .B(n14777), .ZN(
        n14786) );
  AOI211_X1 U16453 ( .C1(n14782), .C2(n14781), .A(n14780), .B(n14838), .ZN(
        n14783) );
  INV_X1 U16454 ( .A(n14783), .ZN(n14785) );
  NAND2_X1 U16455 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n14818), .ZN(n14784) );
  NAND4_X1 U16456 ( .A1(n14787), .A2(n14786), .A3(n14785), .A4(n14784), .ZN(
        P2_U3220) );
  AOI22_X1 U16457 ( .A1(n14818), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3088), .ZN(n14798) );
  OAI211_X1 U16458 ( .C1(n14790), .C2(n14789), .A(n14825), .B(n14788), .ZN(
        n14797) );
  OAI211_X1 U16459 ( .C1(n14793), .C2(n14792), .A(n14820), .B(n14791), .ZN(
        n14796) );
  NAND2_X1 U16460 ( .A1(n14841), .A2(n14794), .ZN(n14795) );
  NAND4_X1 U16461 ( .A1(n14798), .A2(n14797), .A3(n14796), .A4(n14795), .ZN(
        P2_U3227) );
  AOI22_X1 U16462 ( .A1(n14818), .A2(P2_ADDR_REG_14__SCAN_IN), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(P2_U3088), .ZN(n14808) );
  OAI211_X1 U16463 ( .C1(P2_REG2_REG_14__SCAN_IN), .C2(n14800), .A(n14820), 
        .B(n14799), .ZN(n14807) );
  NAND2_X1 U16464 ( .A1(n14841), .A2(n14801), .ZN(n14806) );
  OAI211_X1 U16465 ( .C1(n14804), .C2(n14803), .A(n14825), .B(n14802), .ZN(
        n14805) );
  NAND4_X1 U16466 ( .A1(n14808), .A2(n14807), .A3(n14806), .A4(n14805), .ZN(
        P2_U3228) );
  AOI22_X1 U16467 ( .A1(n14818), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n14817) );
  NAND2_X1 U16468 ( .A1(n14841), .A2(n14809), .ZN(n14816) );
  XOR2_X1 U16469 ( .A(P2_REG2_REG_15__SCAN_IN), .B(n14810), .Z(n14811) );
  NAND2_X1 U16470 ( .A1(n14811), .A2(n14820), .ZN(n14815) );
  XNOR2_X1 U16471 ( .A(n14812), .B(P2_REG1_REG_15__SCAN_IN), .ZN(n14813) );
  NAND2_X1 U16472 ( .A1(n14825), .A2(n14813), .ZN(n14814) );
  NAND4_X1 U16473 ( .A1(n14817), .A2(n14816), .A3(n14815), .A4(n14814), .ZN(
        P2_U3229) );
  AOI22_X1 U16474 ( .A1(n14818), .A2(P2_ADDR_REG_16__SCAN_IN), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(P2_U3088), .ZN(n14831) );
  OAI211_X1 U16475 ( .C1(n14822), .C2(n14821), .A(n14820), .B(n14819), .ZN(
        n14830) );
  NAND2_X1 U16476 ( .A1(n14823), .A2(n14841), .ZN(n14829) );
  OAI211_X1 U16477 ( .C1(n14827), .C2(n14826), .A(n14825), .B(n14824), .ZN(
        n14828) );
  NAND4_X1 U16478 ( .A1(n14831), .A2(n14830), .A3(n14829), .A4(n14828), .ZN(
        P2_U3230) );
  AOI21_X1 U16479 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n14833), .A(n14832), 
        .ZN(n14839) );
  OAI21_X1 U16480 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(n14835), .A(n14834), 
        .ZN(n14837) );
  OAI22_X1 U16481 ( .A1(n14839), .A2(n14838), .B1(n14837), .B2(n14836), .ZN(
        n14840) );
  AOI21_X1 U16482 ( .B1(n14842), .B2(n14841), .A(n14840), .ZN(n14844) );
  OAI211_X1 U16483 ( .C1(n14846), .C2(n14845), .A(n14844), .B(n14843), .ZN(
        P2_U3232) );
  NAND2_X1 U16484 ( .A1(n14848), .A2(n14847), .ZN(n14852) );
  AOI22_X1 U16485 ( .A1(n14478), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n14850), 
        .B2(n14849), .ZN(n14851) );
  OAI211_X1 U16486 ( .C1(n6839), .C2(n14853), .A(n14852), .B(n14851), .ZN(
        n14854) );
  AOI21_X1 U16487 ( .B1(n14856), .B2(n14855), .A(n14854), .ZN(n14857) );
  OAI21_X1 U16488 ( .B1(n14478), .B2(n14858), .A(n14857), .ZN(P2_U3258) );
  INV_X1 U16489 ( .A(n14859), .ZN(n14867) );
  INV_X1 U16490 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n14862) );
  OAI22_X1 U16491 ( .A1(n14863), .A2(n14862), .B1(n14861), .B2(n14860), .ZN(
        n14865) );
  AOI211_X1 U16492 ( .C1(n14867), .C2(n14866), .A(n14865), .B(n14864), .ZN(
        n14869) );
  AOI22_X1 U16493 ( .A1(n14478), .A2(n7405), .B1(n14869), .B2(n14868), .ZN(
        P2_U3265) );
  AND2_X1 U16494 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14874), .ZN(P2_U3266) );
  AND2_X1 U16495 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14874), .ZN(P2_U3267) );
  AND2_X1 U16496 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14874), .ZN(P2_U3268) );
  AND2_X1 U16497 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14874), .ZN(P2_U3269) );
  AND2_X1 U16498 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14874), .ZN(P2_U3270) );
  AND2_X1 U16499 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14874), .ZN(P2_U3271) );
  AND2_X1 U16500 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14874), .ZN(P2_U3272) );
  AND2_X1 U16501 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14874), .ZN(P2_U3273) );
  AND2_X1 U16502 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14874), .ZN(P2_U3274) );
  AND2_X1 U16503 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14874), .ZN(P2_U3275) );
  AND2_X1 U16504 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14874), .ZN(P2_U3276) );
  AND2_X1 U16505 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14874), .ZN(P2_U3277) );
  AND2_X1 U16506 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14874), .ZN(P2_U3278) );
  AND2_X1 U16507 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14874), .ZN(P2_U3279) );
  AND2_X1 U16508 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14874), .ZN(P2_U3280) );
  AND2_X1 U16509 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14874), .ZN(P2_U3281) );
  AND2_X1 U16510 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14874), .ZN(P2_U3282) );
  NOR2_X1 U16511 ( .A1(n14873), .A2(n14871), .ZN(P2_U3283) );
  AND2_X1 U16512 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14874), .ZN(P2_U3284) );
  AND2_X1 U16513 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14874), .ZN(P2_U3285) );
  AND2_X1 U16514 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14874), .ZN(P2_U3286) );
  AND2_X1 U16515 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14874), .ZN(P2_U3287) );
  AND2_X1 U16516 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14874), .ZN(P2_U3288) );
  NOR2_X1 U16517 ( .A1(n14873), .A2(n14872), .ZN(P2_U3289) );
  AND2_X1 U16518 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14874), .ZN(P2_U3290) );
  AND2_X1 U16519 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14874), .ZN(P2_U3291) );
  AND2_X1 U16520 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14874), .ZN(P2_U3292) );
  AND2_X1 U16521 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14874), .ZN(P2_U3293) );
  AND2_X1 U16522 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14874), .ZN(P2_U3294) );
  AND2_X1 U16523 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14874), .ZN(P2_U3295) );
  OAI21_X1 U16524 ( .B1(n14880), .B2(n14876), .A(n14875), .ZN(P2_U3416) );
  AOI22_X1 U16525 ( .A1(n14880), .A2(n14879), .B1(n14878), .B2(n14877), .ZN(
        P2_U3417) );
  INV_X1 U16526 ( .A(n14881), .ZN(n14883) );
  OAI21_X1 U16527 ( .B1(n14883), .B2(n13305), .A(n14882), .ZN(n14884) );
  AOI21_X1 U16528 ( .B1(n14885), .B2(n14892), .A(n14884), .ZN(n14886) );
  AND2_X1 U16529 ( .A1(n14887), .A2(n14886), .ZN(n14899) );
  INV_X1 U16530 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n14888) );
  AOI22_X1 U16531 ( .A1(n14898), .A2(n14899), .B1(n14888), .B2(n14896), .ZN(
        P2_U3454) );
  OAI21_X1 U16532 ( .B1(n14890), .B2(n13305), .A(n14889), .ZN(n14891) );
  AOI21_X1 U16533 ( .B1(n14893), .B2(n14892), .A(n14891), .ZN(n14894) );
  INV_X1 U16534 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n14897) );
  AOI22_X1 U16535 ( .A1(n14898), .A2(n14902), .B1(n14897), .B2(n14896), .ZN(
        P2_U3460) );
  AOI22_X1 U16536 ( .A1(n14903), .A2(n14899), .B1(n10187), .B2(n14900), .ZN(
        P2_U3507) );
  AOI22_X1 U16537 ( .A1(n14903), .A2(n14902), .B1(n14901), .B2(n14900), .ZN(
        P2_U3509) );
  NOR2_X1 U16538 ( .A1(P3_U3897), .A2(n14983), .ZN(P3_U3150) );
  AOI22_X1 U16539 ( .A1(n14960), .A2(P3_IR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n14909) );
  NOR2_X1 U16540 ( .A1(n14904), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n14906) );
  NAND3_X1 U16541 ( .A1(n15023), .A2(n15017), .A3(n15015), .ZN(n14905) );
  OAI21_X1 U16542 ( .B1(n14907), .B2(n14906), .A(n14905), .ZN(n14908) );
  OAI211_X1 U16543 ( .C1(n14910), .C2(n15005), .A(n14909), .B(n14908), .ZN(
        P3_U3182) );
  AOI21_X1 U16544 ( .B1(n14913), .B2(n14912), .A(n14911), .ZN(n14917) );
  AOI21_X1 U16545 ( .B1(n14915), .B2(n15151), .A(n14914), .ZN(n14916) );
  OAI22_X1 U16546 ( .A1(n14917), .A2(n15023), .B1(n15017), .B2(n14916), .ZN(
        n14918) );
  AOI211_X1 U16547 ( .C1(P3_ADDR_REG_3__SCAN_IN), .C2(n14983), .A(n14919), .B(
        n14918), .ZN(n14926) );
  OAI21_X1 U16548 ( .B1(n14922), .B2(n14921), .A(n14920), .ZN(n14924) );
  AOI22_X1 U16549 ( .A1(n14924), .A2(n14963), .B1(n14960), .B2(n14923), .ZN(
        n14925) );
  NAND2_X1 U16550 ( .A1(n14926), .A2(n14925), .ZN(P3_U3185) );
  AOI21_X1 U16551 ( .B1(n14929), .B2(n14928), .A(n14927), .ZN(n14944) );
  INV_X1 U16552 ( .A(n14930), .ZN(n14935) );
  NAND3_X1 U16553 ( .A1(n14933), .A2(n14932), .A3(n14931), .ZN(n14934) );
  AOI21_X1 U16554 ( .B1(n14935), .B2(n14934), .A(n15015), .ZN(n14941) );
  AOI21_X1 U16555 ( .B1(n14938), .B2(n14937), .A(n14936), .ZN(n14939) );
  NOR2_X1 U16556 ( .A1(n14939), .A2(n15017), .ZN(n14940) );
  AOI211_X1 U16557 ( .C1(n14960), .C2(n14942), .A(n14941), .B(n14940), .ZN(
        n14943) );
  OAI21_X1 U16558 ( .B1(n14944), .B2(n15023), .A(n14943), .ZN(n14945) );
  INV_X1 U16559 ( .A(n14945), .ZN(n14947) );
  OAI211_X1 U16560 ( .C1(n14948), .C2(n15005), .A(n14947), .B(n14946), .ZN(
        P3_U3188) );
  AOI21_X1 U16561 ( .B1(n15050), .B2(n14950), .A(n14949), .ZN(n14968) );
  INV_X1 U16562 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n14953) );
  INV_X1 U16563 ( .A(n14951), .ZN(n14952) );
  OAI21_X1 U16564 ( .B1(n15005), .B2(n14953), .A(n14952), .ZN(n14958) );
  AOI21_X1 U16565 ( .B1(n15161), .B2(n14955), .A(n14954), .ZN(n14956) );
  NOR2_X1 U16566 ( .A1(n14956), .A2(n15017), .ZN(n14957) );
  AOI211_X1 U16567 ( .C1(n14960), .C2(n14959), .A(n14958), .B(n14957), .ZN(
        n14967) );
  NOR2_X1 U16568 ( .A1(n14962), .A2(n14961), .ZN(n14964) );
  OAI21_X1 U16569 ( .B1(n14965), .B2(n14964), .A(n14963), .ZN(n14966) );
  OAI211_X1 U16570 ( .C1(n14968), .C2(n15023), .A(n14967), .B(n14966), .ZN(
        P3_U3191) );
  AOI21_X1 U16571 ( .B1(n14971), .B2(n14970), .A(n14969), .ZN(n14985) );
  OAI21_X1 U16572 ( .B1(n15008), .B2(n14973), .A(n14972), .ZN(n14982) );
  AOI21_X1 U16573 ( .B1(n6561), .B2(n14975), .A(n14974), .ZN(n14980) );
  AOI21_X1 U16574 ( .B1(n14978), .B2(n14977), .A(n14976), .ZN(n14979) );
  OAI22_X1 U16575 ( .A1(n14980), .A2(n15017), .B1(n14979), .B2(n15015), .ZN(
        n14981) );
  AOI211_X1 U16576 ( .C1(n14983), .C2(P3_ADDR_REG_10__SCAN_IN), .A(n14982), 
        .B(n14981), .ZN(n14984) );
  OAI21_X1 U16577 ( .B1(n14985), .B2(n15023), .A(n14984), .ZN(P3_U3192) );
  AOI21_X1 U16578 ( .B1(n9068), .B2(n14987), .A(n14986), .ZN(n15001) );
  OAI22_X1 U16579 ( .A1(n15008), .A2(n14989), .B1(n14988), .B2(n15005), .ZN(
        n14998) );
  AOI21_X1 U16580 ( .B1(n9067), .B2(n14991), .A(n14990), .ZN(n14996) );
  AOI21_X1 U16581 ( .B1(n14994), .B2(n14993), .A(n14992), .ZN(n14995) );
  OAI22_X1 U16582 ( .A1(n14996), .A2(n15017), .B1(n14995), .B2(n15015), .ZN(
        n14997) );
  NOR3_X1 U16583 ( .A1(n14999), .A2(n14998), .A3(n14997), .ZN(n15000) );
  OAI21_X1 U16584 ( .B1(n15001), .B2(n15023), .A(n15000), .ZN(P3_U3193) );
  AOI21_X1 U16585 ( .B1(n15004), .B2(n15003), .A(n15002), .ZN(n15024) );
  OAI22_X1 U16586 ( .A1(n15008), .A2(n15007), .B1(n15006), .B2(n15005), .ZN(
        n15020) );
  AOI21_X1 U16587 ( .B1(n15011), .B2(n15010), .A(n15009), .ZN(n15018) );
  AOI21_X1 U16588 ( .B1(n15014), .B2(n15013), .A(n15012), .ZN(n15016) );
  OAI22_X1 U16589 ( .A1(n15018), .A2(n15017), .B1(n15016), .B2(n15015), .ZN(
        n15019) );
  NOR3_X1 U16590 ( .A1(n15021), .A2(n15020), .A3(n15019), .ZN(n15022) );
  OAI21_X1 U16591 ( .B1(n15024), .B2(n15023), .A(n15022), .ZN(P3_U3195) );
  XNOR2_X1 U16592 ( .A(n15025), .B(n15026), .ZN(n15032) );
  INV_X1 U16593 ( .A(n15032), .ZN(n15142) );
  XNOR2_X1 U16594 ( .A(n15027), .B(n15026), .ZN(n15030) );
  OAI22_X1 U16595 ( .A1(n15028), .A2(n15061), .B1(n6892), .B2(n15059), .ZN(
        n15029) );
  AOI21_X1 U16596 ( .B1(n15030), .B2(n15074), .A(n15029), .ZN(n15031) );
  OAI21_X1 U16597 ( .B1(n15067), .B2(n15032), .A(n15031), .ZN(n15140) );
  AOI21_X1 U16598 ( .B1(n15069), .B2(n15142), .A(n15140), .ZN(n15037) );
  NOR2_X1 U16599 ( .A1(n15033), .A2(n15130), .ZN(n15141) );
  AOI22_X1 U16600 ( .A1(n15048), .A2(n15141), .B1(n15090), .B2(n15034), .ZN(
        n15035) );
  OAI221_X1 U16601 ( .B1(n15071), .B2(n15037), .C1(n15094), .C2(n15036), .A(
        n15035), .ZN(P3_U3223) );
  XOR2_X1 U16602 ( .A(n15041), .B(n15038), .Z(n15045) );
  INV_X1 U16603 ( .A(n15045), .ZN(n15138) );
  AOI22_X1 U16604 ( .A1(n15040), .A2(n15076), .B1(n15079), .B2(n15039), .ZN(
        n15044) );
  OAI211_X1 U16605 ( .C1(n6570), .C2(n9820), .A(n15074), .B(n15042), .ZN(
        n15043) );
  OAI211_X1 U16606 ( .C1(n15045), .C2(n15067), .A(n15044), .B(n15043), .ZN(
        n15136) );
  AOI21_X1 U16607 ( .B1(n15069), .B2(n15138), .A(n15136), .ZN(n15051) );
  NOR2_X1 U16608 ( .A1(n15046), .A2(n15130), .ZN(n15137) );
  AOI22_X1 U16609 ( .A1(n15048), .A2(n15137), .B1(n15090), .B2(n15047), .ZN(
        n15049) );
  OAI221_X1 U16610 ( .B1(n15071), .B2(n15051), .C1(n15094), .C2(n15050), .A(
        n15049), .ZN(P3_U3224) );
  XNOR2_X1 U16611 ( .A(n9803), .B(n15052), .ZN(n15066) );
  INV_X1 U16612 ( .A(n15066), .ZN(n15104) );
  NAND2_X1 U16613 ( .A1(n15053), .A2(n15084), .ZN(n15101) );
  OAI22_X1 U16614 ( .A1(n15056), .A2(n15055), .B1(n15054), .B2(n15101), .ZN(
        n15068) );
  OAI21_X1 U16615 ( .B1(n15058), .B2(n9803), .A(n15057), .ZN(n15064) );
  OAI22_X1 U16616 ( .A1(n15062), .A2(n15061), .B1(n15060), .B2(n15059), .ZN(
        n15063) );
  AOI21_X1 U16617 ( .B1(n15064), .B2(n15074), .A(n15063), .ZN(n15065) );
  OAI21_X1 U16618 ( .B1(n15067), .B2(n15066), .A(n15065), .ZN(n15102) );
  AOI211_X1 U16619 ( .C1(n15069), .C2(n15104), .A(n15068), .B(n15102), .ZN(
        n15070) );
  AOI22_X1 U16620 ( .A1(n15071), .A2(n7005), .B1(n15070), .B2(n15094), .ZN(
        P3_U3231) );
  OAI21_X1 U16621 ( .B1(n9801), .B2(n15073), .A(n15072), .ZN(n15075) );
  NAND2_X1 U16622 ( .A1(n15075), .A2(n15074), .ZN(n15081) );
  AOI22_X1 U16623 ( .A1(n15079), .A2(n15078), .B1(n15077), .B2(n15076), .ZN(
        n15080) );
  NAND2_X1 U16624 ( .A1(n15081), .A2(n15080), .ZN(n15096) );
  INV_X1 U16625 ( .A(n15096), .ZN(n15089) );
  XNOR2_X1 U16626 ( .A(n15082), .B(n9801), .ZN(n15098) );
  NAND2_X1 U16627 ( .A1(n15098), .A2(n15083), .ZN(n15088) );
  AND2_X1 U16628 ( .A1(n15085), .A2(n15084), .ZN(n15097) );
  NAND2_X1 U16629 ( .A1(n15097), .A2(n15086), .ZN(n15087) );
  AND3_X1 U16630 ( .A1(n15089), .A2(n15088), .A3(n15087), .ZN(n15095) );
  AOI22_X1 U16631 ( .A1(n15091), .A2(n15098), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15090), .ZN(n15092) );
  OAI221_X1 U16632 ( .B1(n15071), .B2(n15095), .C1(n15094), .C2(n15093), .A(
        n15092), .ZN(P3_U3232) );
  AOI211_X1 U16633 ( .C1(n15099), .C2(n15098), .A(n15097), .B(n15096), .ZN(
        n15148) );
  INV_X1 U16634 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15100) );
  AOI22_X1 U16635 ( .A1(n15146), .A2(n15148), .B1(n15100), .B2(n15144), .ZN(
        P3_U3393) );
  INV_X1 U16636 ( .A(n15101), .ZN(n15103) );
  AOI211_X1 U16637 ( .C1(n15104), .C2(n15143), .A(n15103), .B(n15102), .ZN(
        n15150) );
  INV_X1 U16638 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15105) );
  AOI22_X1 U16639 ( .A1(n15146), .A2(n15150), .B1(n15105), .B2(n15144), .ZN(
        P3_U3396) );
  AOI21_X1 U16640 ( .B1(n15107), .B2(n15143), .A(n15106), .ZN(n15108) );
  AND2_X1 U16641 ( .A1(n15109), .A2(n15108), .ZN(n15152) );
  INV_X1 U16642 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15110) );
  AOI22_X1 U16643 ( .A1(n15146), .A2(n15152), .B1(n15110), .B2(n15144), .ZN(
        P3_U3399) );
  AOI21_X1 U16644 ( .B1(n15112), .B2(n15143), .A(n15111), .ZN(n15113) );
  AND2_X1 U16645 ( .A1(n15114), .A2(n15113), .ZN(n15154) );
  INV_X1 U16646 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15115) );
  AOI22_X1 U16647 ( .A1(n15146), .A2(n15154), .B1(n15115), .B2(n15144), .ZN(
        P3_U3402) );
  AOI211_X1 U16648 ( .C1(n15118), .C2(n15143), .A(n15117), .B(n15116), .ZN(
        n15156) );
  INV_X1 U16649 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15119) );
  AOI22_X1 U16650 ( .A1(n15146), .A2(n15156), .B1(n15119), .B2(n15144), .ZN(
        P3_U3405) );
  INV_X1 U16651 ( .A(n15120), .ZN(n15123) );
  AOI211_X1 U16652 ( .C1(n15123), .C2(n15143), .A(n15122), .B(n15121), .ZN(
        n15157) );
  AOI22_X1 U16653 ( .A1(n15146), .A2(n15157), .B1(n15124), .B2(n15144), .ZN(
        P3_U3408) );
  NOR2_X1 U16654 ( .A1(n15125), .A2(n15130), .ZN(n15127) );
  AOI211_X1 U16655 ( .C1(n15128), .C2(n15143), .A(n15127), .B(n15126), .ZN(
        n15158) );
  INV_X1 U16656 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15129) );
  AOI22_X1 U16657 ( .A1(n15146), .A2(n15158), .B1(n15129), .B2(n15144), .ZN(
        P3_U3411) );
  NOR2_X1 U16658 ( .A1(n15131), .A2(n15130), .ZN(n15133) );
  AOI211_X1 U16659 ( .C1(n15134), .C2(n15143), .A(n15133), .B(n15132), .ZN(
        n15160) );
  INV_X1 U16660 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15135) );
  AOI22_X1 U16661 ( .A1(n15146), .A2(n15160), .B1(n15135), .B2(n15144), .ZN(
        P3_U3414) );
  AOI211_X1 U16662 ( .C1(n15138), .C2(n15143), .A(n15137), .B(n15136), .ZN(
        n15162) );
  INV_X1 U16663 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15139) );
  AOI22_X1 U16664 ( .A1(n15146), .A2(n15162), .B1(n15139), .B2(n15144), .ZN(
        P3_U3417) );
  AOI211_X1 U16665 ( .C1(n15143), .C2(n15142), .A(n15141), .B(n15140), .ZN(
        n15165) );
  INV_X1 U16666 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15145) );
  AOI22_X1 U16667 ( .A1(n15146), .A2(n15165), .B1(n15145), .B2(n15144), .ZN(
        P3_U3420) );
  AOI22_X1 U16668 ( .A1(n15166), .A2(n15148), .B1(n15147), .B2(n15163), .ZN(
        P3_U3460) );
  AOI22_X1 U16669 ( .A1(n15166), .A2(n15150), .B1(n15149), .B2(n15163), .ZN(
        P3_U3461) );
  AOI22_X1 U16670 ( .A1(n15166), .A2(n15152), .B1(n15151), .B2(n15163), .ZN(
        P3_U3462) );
  AOI22_X1 U16671 ( .A1(n15166), .A2(n15154), .B1(n15153), .B2(n15163), .ZN(
        P3_U3463) );
  AOI22_X1 U16672 ( .A1(n15166), .A2(n15156), .B1(n15155), .B2(n15163), .ZN(
        P3_U3464) );
  AOI22_X1 U16673 ( .A1(n15166), .A2(n15157), .B1(n9077), .B2(n15163), .ZN(
        P3_U3465) );
  AOI22_X1 U16674 ( .A1(n15166), .A2(n15158), .B1(n9082), .B2(n15163), .ZN(
        P3_U3466) );
  AOI22_X1 U16675 ( .A1(n15166), .A2(n15160), .B1(n15159), .B2(n15163), .ZN(
        P3_U3467) );
  AOI22_X1 U16676 ( .A1(n15166), .A2(n15162), .B1(n15161), .B2(n15163), .ZN(
        P3_U3468) );
  AOI22_X1 U16677 ( .A1(n15166), .A2(n15165), .B1(n15164), .B2(n15163), .ZN(
        P3_U3469) );
  XOR2_X1 U16678 ( .A(n15168), .B(n15167), .Z(SUB_1596_U59) );
  XNOR2_X1 U16679 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n15169), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U16680 ( .B1(n15171), .B2(n15170), .A(n15180), .ZN(SUB_1596_U53) );
  XOR2_X1 U16681 ( .A(n15173), .B(n15172), .Z(SUB_1596_U56) );
  OAI21_X1 U16682 ( .B1(n15176), .B2(n15175), .A(n15174), .ZN(n15178) );
  XOR2_X1 U16683 ( .A(n15178), .B(n15177), .Z(SUB_1596_U60) );
  XOR2_X1 U16684 ( .A(n15180), .B(n15179), .Z(SUB_1596_U5) );
  CLKBUF_X1 U7198 ( .A(n6849), .Z(n6843) );
  CLKBUF_X1 U7220 ( .A(n13234), .Z(n6593) );
  CLKBUF_X2 U7249 ( .A(n9693), .Z(n6424) );
  CLKBUF_X3 U7785 ( .A(n9693), .Z(n6425) );
  CLKBUF_X1 U8256 ( .A(n9193), .Z(n9194) );
  INV_X2 U9407 ( .A(n7799), .ZN(n13083) );
endmodule

