

module b20_C_AntiSAT_k_256_7 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, ADD_1068_U4, ADD_1068_U55, 
        ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, 
        ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, 
        ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, 
        ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, 
        P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, 
        P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, 
        P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, 
        P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, 
        P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, 
        P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, 
        P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, 
        P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, 
        P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, 
        P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, 
        P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, 
        P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, 
        P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, 
        P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, 
        P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, 
        P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, 
        P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, 
        P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, 
        P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, 
        P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, 
        P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, 
        P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503;

  AND2_X1 U4998 ( .A1(n4660), .A2(n8122), .ZN(n4659) );
  CLKBUF_X2 U4999 ( .A(n8627), .Z(n8728) );
  INV_X1 U5000 ( .A(n5166), .ZN(n5434) );
  CLKBUF_X2 U5001 ( .A(n8735), .Z(n4503) );
  CLKBUF_X3 U5002 ( .A(n8587), .Z(n4493) );
  NAND2_X1 U5003 ( .A1(n4726), .A2(n4725), .ZN(n5210) );
  INV_X1 U5004 ( .A(n7900), .ZN(n5982) );
  INV_X1 U5005 ( .A(n8553), .ZN(n5974) );
  CLKBUF_X2 U5006 ( .A(n4497), .Z(n4499) );
  NAND2_X1 U5007 ( .A1(n4939), .A2(n4937), .ZN(n5442) );
  NOR3_X1 U5008 ( .A1(n5736), .A2(n5735), .A3(n5734), .ZN(n9232) );
  AOI21_X1 U5009 ( .B1(n7182), .B2(n6110), .A(n4534), .ZN(n7254) );
  INV_X1 U5010 ( .A(n9381), .ZN(n5726) );
  INV_X1 U5011 ( .A(n5151), .ZN(n5330) );
  INV_X1 U5012 ( .A(n6314), .ZN(n6050) );
  NAND2_X1 U5013 ( .A1(n7959), .A2(n7966), .ZN(n6711) );
  NAND2_X1 U5014 ( .A1(n6307), .A2(n8067), .ZN(n8376) );
  INV_X1 U5015 ( .A(n8286), .ZN(n6043) );
  INV_X1 U5016 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n4674) );
  CLKBUF_X3 U5017 ( .A(n4493), .Z(n7517) );
  OAI21_X1 U5018 ( .B1(n6771), .B2(n6773), .A(n6772), .ZN(n6923) );
  NOR2_X1 U5019 ( .A1(n7744), .A2(n7621), .ZN(n4915) );
  INV_X1 U5021 ( .A(n5173), .ZN(n5406) );
  AOI211_X1 U5022 ( .C1(n7653), .C2(n7441), .A(n9794), .B(n7503), .ZN(n7579)
         );
  INV_X1 U5023 ( .A(n7361), .ZN(n10138) );
  NAND2_X1 U5024 ( .A1(n5886), .A2(n5889), .ZN(n6322) );
  CLKBUF_X2 U5025 ( .A(n5889), .Z(n5948) );
  INV_X1 U5026 ( .A(n5455), .ZN(n9365) );
  XNOR2_X1 U5027 ( .A(n5239), .B(n5238), .ZN(n6480) );
  NAND2_X1 U5028 ( .A1(n5172), .A2(n5171), .ZN(n5179) );
  MUX2_X1 U5029 ( .A(n8449), .B(n8502), .S(n10446), .Z(n8450) );
  MUX2_X1 U5030 ( .A(n8503), .B(n8502), .S(n10430), .Z(n8504) );
  NOR2_X1 U5031 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5922) );
  BUF_X4 U5032 ( .A(n4497), .Z(n4500) );
  INV_X2 U5034 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5108) );
  AOI211_X1 U5035 ( .C1(n7304), .C2(n9385), .A(n7305), .B(n5733), .ZN(n5736)
         );
  NAND2_X1 U5036 ( .A1(n9137), .A2(n8595), .ZN(n9183) );
  INV_X4 U5037 ( .A(n8627), .ZN(n8733) );
  NAND2_X2 U5038 ( .A1(n5245), .A2(n5244), .ZN(n7653) );
  OAI21_X2 U5039 ( .B1(n8719), .B2(n8717), .A(n8715), .ZN(n9160) );
  OAI21_X2 U5040 ( .B1(n5210), .B2(n5209), .A(n5211), .ZN(n5221) );
  NAND2_X1 U5041 ( .A1(n6530), .A2(n6529), .ZN(n8587) );
  OAI222_X1 U5042 ( .A1(n8555), .A2(n8554), .B1(P2_U3151), .B2(n8553), .C1(
        n8552), .C2(n8551), .ZN(P2_U3266) );
  XNOR2_X2 U5043 ( .A(n5972), .B(n5971), .ZN(n8553) );
  AOI21_X2 U5044 ( .B1(n7636), .B2(n7635), .A(n4543), .ZN(n4927) );
  OR2_X1 U5045 ( .A1(n7647), .A2(n7646), .ZN(n4543) );
  AOI21_X2 U5046 ( .B1(n7634), .B2(n7633), .A(n7632), .ZN(n7635) );
  AND2_X1 U5047 ( .A1(n4659), .A2(n4658), .ZN(n4654) );
  NAND2_X1 U5048 ( .A1(n8735), .A2(n8587), .ZN(n7040) );
  INV_X1 U5049 ( .A(n8735), .ZN(n8653) );
  INV_X1 U5050 ( .A(n6763), .ZN(n5507) );
  INV_X2 U5051 ( .A(n4493), .ZN(n8731) );
  AND2_X1 U5053 ( .A1(n9720), .A2(n7225), .ZN(n6545) );
  AOI21_X1 U5054 ( .B1(n5191), .B2(n4991), .A(n4548), .ZN(n4990) );
  BUF_X4 U5055 ( .A(n5527), .Z(n4494) );
  CLKBUF_X1 U5056 ( .A(n6031), .Z(n7893) );
  NAND2_X1 U5058 ( .A1(n7873), .A2(n4731), .ZN(n5958) );
  OR2_X1 U5059 ( .A1(n8739), .A2(n4590), .ZN(n8751) );
  OAI21_X1 U5060 ( .B1(n7881), .B2(n9815), .A(n7874), .ZN(n4732) );
  AND2_X1 U5061 ( .A1(n8696), .A2(n8695), .ZN(n9151) );
  NOR2_X1 U5062 ( .A1(n9813), .A2(n9812), .ZN(n9814) );
  NAND2_X1 U5063 ( .A1(n7792), .A2(n7791), .ZN(n9813) );
  OAI22_X1 U5064 ( .A1(n8635), .A2(n8636), .B1(n8690), .B2(n8632), .ZN(n4930)
         );
  MUX2_X1 U5065 ( .A(n9325), .B(n9324), .S(n9458), .Z(n9326) );
  OR2_X1 U5066 ( .A1(n8495), .A2(n8293), .ZN(n8119) );
  NAND2_X1 U5067 ( .A1(n5695), .A2(n5694), .ZN(n9632) );
  OAI21_X1 U5068 ( .B1(n9618), .B2(n4717), .A(n4715), .ZN(n7782) );
  NAND2_X1 U5069 ( .A1(n5685), .A2(n5098), .ZN(n4789) );
  OAI21_X1 U5070 ( .B1(n8324), .B2(n6261), .A(n4512), .ZN(n8313) );
  OR2_X1 U5071 ( .A1(n5425), .A2(n5424), .ZN(n5430) );
  OAI21_X1 U5072 ( .B1(n5419), .B2(n9107), .A(n5418), .ZN(n5425) );
  AOI211_X1 U5073 ( .C1(n9308), .C2(n9307), .A(n9303), .B(n9448), .ZN(n9304)
         );
  OR2_X1 U5074 ( .A1(n5765), .A2(n8745), .ZN(n7793) );
  XNOR2_X1 U5075 ( .A(n5417), .B(n5416), .ZN(n5419) );
  NAND2_X1 U5076 ( .A1(n6274), .A2(n6273), .ZN(n8303) );
  NAND2_X1 U5077 ( .A1(n5408), .A2(n5407), .ZN(n8745) );
  OR2_X1 U5078 ( .A1(n8448), .A2(n8327), .ZN(n8094) );
  NAND2_X1 U5079 ( .A1(n5402), .A2(n5401), .ZN(n9628) );
  NAND2_X1 U5080 ( .A1(n6263), .A2(n6262), .ZN(n8448) );
  NOR2_X1 U5081 ( .A1(n4788), .A2(n4574), .ZN(n4787) );
  NAND2_X1 U5082 ( .A1(n8421), .A2(n8420), .ZN(n8477) );
  NAND2_X1 U5083 ( .A1(n8486), .A2(n7928), .ZN(n8421) );
  AOI21_X1 U5084 ( .B1(n4764), .B2(n4762), .A(n4761), .ZN(n4760) );
  NAND2_X1 U5085 ( .A1(n7733), .A2(n4769), .ZN(n8486) );
  NAND2_X1 U5086 ( .A1(n5373), .A2(n5372), .ZN(n9671) );
  NAND2_X1 U5087 ( .A1(n6130), .A2(n5061), .ZN(n5060) );
  NAND2_X1 U5088 ( .A1(n5343), .A2(n5342), .ZN(n9715) );
  NAND2_X1 U5089 ( .A1(n6210), .A2(n6209), .ZN(n8463) );
  NAND2_X1 U5090 ( .A1(n4702), .A2(n4700), .ZN(n9789) );
  AND2_X1 U5091 ( .A1(n5338), .A2(n5337), .ZN(n9913) );
  NAND2_X1 U5092 ( .A1(n6178), .A2(n6177), .ZN(n8435) );
  NAND2_X1 U5093 ( .A1(n5315), .A2(n5314), .ZN(n9765) );
  NAND2_X1 U5094 ( .A1(n4839), .A2(n4840), .ZN(n5356) );
  NAND2_X1 U5095 ( .A1(n7386), .A2(n4729), .ZN(n7496) );
  OAI21_X1 U5096 ( .B1(n5320), .B2(n5319), .A(n5318), .ZN(n5335) );
  NAND2_X1 U5097 ( .A1(n7324), .A2(n7238), .ZN(n7515) );
  NAND2_X1 U5098 ( .A1(n5280), .A2(n5279), .ZN(n9218) );
  NAND2_X1 U5099 ( .A1(n7234), .A2(n7233), .ZN(n7324) );
  OR2_X1 U5100 ( .A1(n7351), .A2(n9396), .ZN(n7385) );
  AND2_X1 U5101 ( .A1(n7406), .A2(n10169), .ZN(n7442) );
  NAND2_X1 U5102 ( .A1(n7290), .A2(n9394), .ZN(n7351) );
  AND2_X1 U5103 ( .A1(n7640), .A2(n7639), .ZN(n7684) );
  NOR2_X1 U5104 ( .A1(n6959), .A2(n6960), .ZN(n7057) );
  NAND2_X2 U5105 ( .A1(n5237), .A2(n5236), .ZN(n7693) );
  AND2_X1 U5106 ( .A1(n6091), .A2(n6090), .ZN(n10419) );
  NAND2_X1 U5107 ( .A1(n4593), .A2(n5224), .ZN(n8713) );
  NAND2_X1 U5108 ( .A1(n6604), .A2(n10373), .ZN(n8237) );
  INV_X1 U5109 ( .A(n10398), .ZN(n7008) );
  INV_X1 U5110 ( .A(n7510), .ZN(n5006) );
  INV_X1 U5111 ( .A(n10044), .ZN(n10145) );
  OAI211_X1 U5112 ( .C1(n5151), .C2(n6440), .A(n5185), .B(n5184), .ZN(n7361)
         );
  AND2_X1 U5113 ( .A1(n6074), .A2(n6073), .ZN(n7114) );
  INV_X2 U5114 ( .A(n10381), .ZN(n4495) );
  OAI21_X2 U5115 ( .B1(n6458), .B2(n6080), .A(n6079), .ZN(n10416) );
  AND2_X1 U5116 ( .A1(n7983), .A2(n7992), .ZN(n7911) );
  OAI211_X1 U5117 ( .C1(n5151), .C2(n6435), .A(n5175), .B(n5174), .ZN(n7298)
         );
  NAND2_X2 U5119 ( .A1(n6613), .A2(n10383), .ZN(n7959) );
  INV_X1 U5120 ( .A(n7279), .ZN(n10104) );
  INV_X1 U5121 ( .A(n8282), .ZN(n7152) );
  INV_X1 U5122 ( .A(n7314), .ZN(n10125) );
  XNOR2_X1 U5123 ( .A(n8289), .B(n6658), .ZN(n7971) );
  INV_X2 U5124 ( .A(n6467), .ZN(n6501) );
  NAND3_X1 U5125 ( .A1(n5493), .A2(n5492), .A3(n5491), .ZN(n7279) );
  NAND3_X1 U5126 ( .A1(n5093), .A2(n6000), .A3(n5999), .ZN(n8289) );
  AND4_X1 U5127 ( .A1(n5992), .A2(n5993), .A3(n5991), .A4(n5990), .ZN(n6717)
         );
  OR2_X1 U5128 ( .A1(n5166), .A2(n6444), .ZN(n5492) );
  NAND2_X2 U5129 ( .A1(n4915), .A2(n5468), .ZN(n6530) );
  MUX2_X1 U5130 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9937), .S(n5127), .Z(n7172) );
  NOR2_X2 U5131 ( .A1(n8106), .A2(n6656), .ZN(n6321) );
  AOI21_X1 U5132 ( .B1(n4858), .B2(n4520), .A(n4857), .ZN(n4856) );
  AOI21_X1 U5133 ( .B1(n4728), .B2(n5199), .A(n4547), .ZN(n4725) );
  NAND2_X1 U5135 ( .A1(n5462), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U5136 ( .A1(n5462), .A2(n5461), .ZN(n7744) );
  XNOR2_X1 U5137 ( .A(n5470), .B(n5469), .ZN(n5455) );
  NOR2_X1 U5138 ( .A1(n4992), .A2(n4989), .ZN(n4988) );
  XNOR2_X1 U5139 ( .A(n5464), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5467) );
  OR2_X1 U5140 ( .A1(n8547), .A2(n4674), .ZN(n5969) );
  XNOR2_X1 U5141 ( .A(n5445), .B(n5444), .ZN(n7884) );
  OR2_X1 U5142 ( .A1(n5118), .A2(n5117), .ZN(n5123) );
  OR2_X1 U5143 ( .A1(n5463), .A2(n9931), .ZN(n5464) );
  NAND2_X1 U5144 ( .A1(n5448), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5450) );
  NAND2_X1 U5145 ( .A1(n9932), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5445) );
  XNOR2_X1 U5146 ( .A(n5439), .B(n5438), .ZN(n9381) );
  NAND2_X1 U5147 ( .A1(n5441), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U5148 ( .A1(n4526), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5439) );
  NAND2_X1 U5149 ( .A1(n4527), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5312) );
  NAND2_X2 U5150 ( .A1(n4835), .A2(P1_U3086), .ZN(n7819) );
  INV_X2 U5151 ( .A(n7574), .ZN(n4496) );
  AND2_X1 U5152 ( .A1(n5163), .A2(n5164), .ZN(n5177) );
  AND2_X1 U5153 ( .A1(n4776), .A2(n5056), .ZN(n4775) );
  AND2_X1 U5154 ( .A1(n5021), .A2(n5113), .ZN(n5020) );
  INV_X2 U5155 ( .A(n5124), .ZN(n4497) );
  NOR2_X1 U5156 ( .A1(n5152), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5163) );
  AND4_X1 U5157 ( .A1(n5277), .A2(n8789), .A3(n5241), .A4(n5110), .ZN(n4778)
         );
  NOR2_X1 U5158 ( .A1(n5078), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n5021) );
  INV_X1 U5159 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5444) );
  INV_X1 U5160 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5832) );
  INV_X1 U5161 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5277) );
  INV_X1 U5162 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5241) );
  INV_X1 U5163 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5779) );
  NOR2_X1 U5164 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5107) );
  INV_X1 U5165 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5164) );
  NOR2_X1 U5166 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4916) );
  NOR2_X2 U5167 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5129) );
  INV_X1 U5168 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5968) );
  INV_X1 U5169 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5825) );
  INV_X1 U5170 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8789) );
  INV_X4 U5171 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  AOI21_X2 U5172 ( .B1(n8770), .B2(n8591), .A(n5086), .ZN(n9137) );
  BUF_X1 U5173 ( .A(n4497), .Z(n4498) );
  NAND2_X1 U5174 ( .A1(n6923), .A2(n6922), .ZN(n6924) );
  AND2_X4 U5176 ( .A1(n5495), .A2(n5494), .ZN(n5518) );
  NAND3_X1 U5177 ( .A1(n6526), .A2(n6530), .A3(n10045), .ZN(n8735) );
  NAND2_X1 U5178 ( .A1(n8577), .A2(n8576), .ZN(n8581) );
  AND2_X1 U5179 ( .A1(n7884), .A2(n5494), .ZN(n5527) );
  OAI21_X2 U5180 ( .B1(n6458), .B2(n5166), .A(n4733), .ZN(n7605) );
  XNOR2_X2 U5181 ( .A(n5225), .B(n5226), .ZN(n6460) );
  NOR2_X2 U5182 ( .A1(n5442), .A2(n4829), .ZN(n5440) );
  OAI21_X2 U5183 ( .B1(n9183), .B2(n9179), .A(n9180), .ZN(n8719) );
  NAND2_X1 U5184 ( .A1(n6639), .A2(n6638), .ZN(n6761) );
  NAND2_X2 U5185 ( .A1(n5454), .A2(n5456), .ZN(n5127) );
  XNOR2_X2 U5186 ( .A(n5116), .B(n5115), .ZN(n5454) );
  AOI211_X1 U5187 ( .C1(n6763), .C2(n7274), .A(n9794), .B(n10064), .ZN(n10110)
         );
  NOR2_X1 U5188 ( .A1(n7274), .A2(n6763), .ZN(n10064) );
  NOR2_X2 U5189 ( .A1(n6641), .A2(n6640), .ZN(n6771) );
  AND2_X1 U5190 ( .A1(n4995), .A2(n4994), .ZN(n4504) );
  AOI21_X1 U5191 ( .B1(n4867), .B2(n4868), .A(n5255), .ZN(n4865) );
  INV_X1 U5192 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5003) );
  NAND2_X1 U5193 ( .A1(n8128), .A2(n7957), .ZN(n8106) );
  NAND2_X1 U5194 ( .A1(n9253), .A2(n9258), .ZN(n4597) );
  INV_X1 U5195 ( .A(n5344), .ZN(n5345) );
  XNOR2_X1 U5196 ( .A(n6681), .B(n4697), .ZN(n7108) );
  INV_X1 U5197 ( .A(n10406), .ZN(n4697) );
  NAND2_X1 U5198 ( .A1(n4974), .A2(n4542), .ZN(n6651) );
  XNOR2_X1 U5199 ( .A(n6681), .B(n10394), .ZN(n4980) );
  NAND2_X1 U5200 ( .A1(n4986), .A2(n4985), .ZN(n4984) );
  AOI21_X1 U5201 ( .B1(n8495), .B2(n8105), .A(n7963), .ZN(n4985) );
  OAI211_X1 U5202 ( .C1(n7898), .C2(n7897), .A(n4545), .B(n8119), .ZN(n4986)
         );
  INV_X1 U5203 ( .A(n5973), .ZN(n5975) );
  AND2_X1 U5204 ( .A1(n5042), .A2(n5041), .ZN(n5040) );
  NAND2_X1 U5205 ( .A1(n4521), .A2(n6261), .ZN(n5041) );
  NAND2_X1 U5206 ( .A1(n6309), .A2(n5043), .ZN(n5042) );
  OR2_X1 U5207 ( .A1(n8181), .A2(n8187), .ZN(n8041) );
  INV_X1 U5208 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5785) );
  NOR2_X1 U5209 ( .A1(n5780), .A2(n5781), .ZN(n5782) );
  AND2_X1 U5210 ( .A1(n4775), .A2(n4777), .ZN(n4881) );
  XNOR2_X1 U5211 ( .A(n5450), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5494) );
  NAND2_X1 U5212 ( .A1(n9237), .A2(n9233), .ZN(n4699) );
  INV_X1 U5213 ( .A(n5127), .ZN(n5140) );
  AND2_X1 U5214 ( .A1(n5440), .A2(n5113), .ZN(n5463) );
  AND2_X1 U5215 ( .A1(n5308), .A2(n5303), .ZN(n5306) );
  INV_X1 U5216 ( .A(n4859), .ZN(n4858) );
  OAI21_X1 U5217 ( .B1(n4862), .B2(n4520), .A(n5296), .ZN(n4859) );
  INV_X1 U5218 ( .A(n5240), .ZN(n4870) );
  OAI21_X1 U5219 ( .B1(n4500), .B2(P1_DATAO_REG_5__SCAN_IN), .A(n4594), .ZN(
        n5180) );
  NAND2_X1 U5220 ( .A1(n4499), .A2(n6436), .ZN(n4594) );
  XNOR2_X1 U5221 ( .A(n5811), .B(n5810), .ZN(n5889) );
  OR2_X1 U5222 ( .A1(n5795), .A2(n4674), .ZN(n5811) );
  NAND2_X1 U5223 ( .A1(n4695), .A2(n4571), .ZN(n4693) );
  INV_X1 U5224 ( .A(n7902), .ZN(n6316) );
  XNOR2_X1 U5225 ( .A(n4980), .B(n8286), .ZN(n6957) );
  NAND2_X1 U5226 ( .A1(n6322), .A2(n4499), .ZN(n6031) );
  INV_X1 U5227 ( .A(n4680), .ZN(n4679) );
  AOI21_X1 U5228 ( .B1(n4680), .B2(n4678), .A(n4550), .ZN(n4677) );
  INV_X1 U5229 ( .A(n7826), .ZN(n4678) );
  OR2_X1 U5230 ( .A1(n7748), .A2(n7749), .ZN(n4696) );
  INV_X1 U5232 ( .A(n8130), .ZN(n4657) );
  OR2_X1 U5233 ( .A1(n8117), .A2(n8116), .ZN(n8120) );
  INV_X1 U5234 ( .A(n6285), .ZN(n6266) );
  NOR2_X1 U5235 ( .A1(n4530), .A2(n10235), .ZN(n10234) );
  NAND2_X1 U5236 ( .A1(n4906), .A2(n5920), .ZN(n4905) );
  AOI21_X1 U5237 ( .B1(n5055), .B2(n4505), .A(n4549), .ZN(n5054) );
  NAND2_X1 U5238 ( .A1(n8399), .A2(n6198), .ZN(n8385) );
  NAND2_X1 U5239 ( .A1(n7837), .A2(n8390), .ZN(n6198) );
  NAND2_X1 U5240 ( .A1(n6322), .A2(n4835), .ZN(n6080) );
  INV_X1 U5241 ( .A(n7963), .ZN(n7957) );
  OR2_X1 U5242 ( .A1(n8513), .A2(n8350), .ZN(n5044) );
  NAND2_X1 U5243 ( .A1(n5070), .A2(n5069), .ZN(n8399) );
  AND2_X1 U5244 ( .A1(n8400), .A2(n4569), .ZN(n5069) );
  NOR2_X1 U5245 ( .A1(n4533), .A2(n5059), .ZN(n5058) );
  AND4_X1 U5246 ( .A1(n6139), .A2(n6138), .A3(n6137), .A4(n6136), .ZN(n8259)
         );
  INV_X1 U5247 ( .A(n8427), .ZN(n8391) );
  INV_X1 U5248 ( .A(n6080), .ZN(n7891) );
  INV_X1 U5249 ( .A(n6031), .ZN(n6176) );
  INV_X1 U5250 ( .A(n6322), .ZN(n6175) );
  AND2_X1 U5251 ( .A1(n8112), .A2(n6656), .ZN(n8427) );
  XNOR2_X1 U5252 ( .A(n5809), .B(n5967), .ZN(n5886) );
  NAND2_X1 U5253 ( .A1(n5966), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5809) );
  AND2_X1 U5254 ( .A1(n4777), .A2(n4559), .ZN(n4774) );
  NOR2_X1 U5255 ( .A1(n9998), .A2(n9997), .ZN(n9996) );
  NAND2_X1 U5256 ( .A1(n9880), .A2(n5012), .ZN(n5016) );
  NAND2_X1 U5257 ( .A1(n4820), .A2(n4509), .ZN(n4817) );
  NAND2_X1 U5258 ( .A1(n4553), .A2(n4509), .ZN(n4816) );
  NAND2_X1 U5259 ( .A1(n4823), .A2(n4820), .ZN(n4819) );
  INV_X1 U5260 ( .A(n4811), .ZN(n4810) );
  OAI21_X1 U5261 ( .B1(n4812), .B2(n9347), .A(n5607), .ZN(n4811) );
  AND2_X1 U5262 ( .A1(n5741), .A2(n9402), .ZN(n4729) );
  OR2_X1 U5263 ( .A1(n7164), .A2(n9467), .ZN(n9794) );
  AOI21_X1 U5264 ( .B1(n5764), .B2(n10054), .A(n8741), .ZN(n7873) );
  XNOR2_X1 U5265 ( .A(n7782), .B(n5722), .ZN(n5764) );
  AND2_X1 U5266 ( .A1(n10031), .A2(n10143), .ZN(n9815) );
  NAND2_X1 U5267 ( .A1(n5020), .A2(n4828), .ZN(n4827) );
  NOR2_X1 U5268 ( .A1(n6977), .A2(n4878), .ZN(n6838) );
  NOR2_X1 U5269 ( .A1(n4879), .A2(n4609), .ZN(n4878) );
  INV_X1 U5270 ( .A(n5895), .ZN(n4879) );
  OR2_X1 U5271 ( .A1(n6855), .A2(n6856), .ZN(n4876) );
  INV_X1 U5272 ( .A(n9720), .ZN(n9598) );
  NAND2_X1 U5273 ( .A1(n4624), .A2(n8106), .ZN(n4623) );
  NAND2_X1 U5274 ( .A1(n4625), .A2(n7997), .ZN(n4624) );
  NAND2_X1 U5275 ( .A1(n7999), .A2(n7998), .ZN(n4625) );
  AND2_X1 U5276 ( .A1(n8002), .A2(n8001), .ZN(n4621) );
  NAND2_X1 U5277 ( .A1(n4643), .A2(n8106), .ZN(n4642) );
  NAND2_X1 U5278 ( .A1(n8011), .A2(n8010), .ZN(n4643) );
  NAND2_X1 U5279 ( .A1(n4641), .A2(n4640), .ZN(n4639) );
  NOR2_X1 U5280 ( .A1(n8005), .A2(n8106), .ZN(n4640) );
  NAND2_X1 U5281 ( .A1(n8007), .A2(n8006), .ZN(n4641) );
  NAND2_X1 U5282 ( .A1(n4555), .A2(n8039), .ZN(n4634) );
  NAND2_X1 U5283 ( .A1(n4508), .A2(n7527), .ZN(n4633) );
  NAND2_X1 U5284 ( .A1(n4516), .A2(n4632), .ZN(n4631) );
  NAND2_X1 U5285 ( .A1(n8034), .A2(n4508), .ZN(n4632) );
  NAND2_X1 U5286 ( .A1(n8420), .A2(n8046), .ZN(n4636) );
  AND2_X1 U5287 ( .A1(n5333), .A2(SI_20_), .ZN(n4853) );
  INV_X1 U5288 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5778) );
  INV_X1 U5289 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5777) );
  INV_X1 U5290 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5775) );
  NOR2_X1 U5291 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5776) );
  NAND2_X1 U5292 ( .A1(n9313), .A2(n9309), .ZN(n9448) );
  NOR2_X1 U5293 ( .A1(n9765), .A2(n9333), .ZN(n5009) );
  INV_X1 U5294 ( .A(n4846), .ZN(n4843) );
  INV_X1 U5295 ( .A(n4523), .ZN(n4841) );
  AOI21_X1 U5296 ( .B1(n5334), .B2(n4853), .A(n4852), .ZN(n4851) );
  INV_X1 U5297 ( .A(n5339), .ZN(n4852) );
  AOI21_X1 U5298 ( .B1(n5334), .B2(n5333), .A(SI_20_), .ZN(n4854) );
  NAND2_X1 U5299 ( .A1(n7750), .A2(n8277), .ZN(n4695) );
  NAND2_X1 U5300 ( .A1(n4967), .A2(n7059), .ZN(n4966) );
  INV_X1 U5301 ( .A(n7056), .ZN(n4967) );
  INV_X1 U5302 ( .A(n4693), .ZN(n4692) );
  NAND2_X1 U5303 ( .A1(n6312), .A2(n7963), .ZN(n4983) );
  OR2_X1 U5304 ( .A1(n6966), .A2(n4608), .ZN(n4607) );
  NOR2_X1 U5305 ( .A1(n4609), .A2(n10369), .ZN(n4608) );
  NAND2_X1 U5306 ( .A1(n6857), .A2(n4739), .ZN(n5930) );
  OR2_X1 U5307 ( .A1(n6869), .A2(n6023), .ZN(n4739) );
  NAND2_X1 U5308 ( .A1(n5864), .A2(n5095), .ZN(n5865) );
  NAND2_X1 U5309 ( .A1(n6878), .A2(n4568), .ZN(n5932) );
  NAND2_X1 U5310 ( .A1(n10226), .A2(n4606), .ZN(n5872) );
  OR2_X1 U5311 ( .A1(n10225), .A2(n5867), .ZN(n4606) );
  AOI21_X1 U5312 ( .B1(n10250), .B2(n4888), .A(n10267), .ZN(n4887) );
  NAND2_X1 U5313 ( .A1(n10258), .A2(n4602), .ZN(n5875) );
  OR2_X1 U5314 ( .A1(n10257), .A2(n5874), .ZN(n4602) );
  NAND2_X1 U5315 ( .A1(n10261), .A2(n4740), .ZN(n5936) );
  OR2_X1 U5316 ( .A1(n10257), .A2(n9052), .ZN(n4740) );
  NAND2_X1 U5317 ( .A1(n10294), .A2(n4742), .ZN(n5938) );
  NAND2_X1 U5318 ( .A1(n6522), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4742) );
  NAND2_X1 U5319 ( .A1(n5913), .A2(n10307), .ZN(n4899) );
  NOR2_X1 U5320 ( .A1(n4900), .A2(n4896), .ZN(n4895) );
  INV_X1 U5321 ( .A(n4899), .ZN(n4896) );
  NOR2_X1 U5322 ( .A1(n7936), .A2(n4521), .ZN(n5037) );
  NOR2_X1 U5323 ( .A1(n8114), .A2(n8315), .ZN(n5036) );
  INV_X1 U5324 ( .A(n7936), .ZN(n5039) );
  NOR2_X1 U5325 ( .A1(n6231), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6244) );
  NAND2_X1 U5326 ( .A1(n6154), .A2(n5964), .ZN(n6179) );
  NAND2_X1 U5327 ( .A1(n6940), .A2(n5995), .ZN(n7966) );
  AND2_X1 U5328 ( .A1(n6349), .A2(n6348), .ZN(n6378) );
  NOR2_X1 U5329 ( .A1(n7908), .A2(n4764), .ZN(n4758) );
  OR2_X1 U5330 ( .A1(n8518), .A2(n8361), .ZN(n8083) );
  OR2_X1 U5331 ( .A1(n8469), .A2(n8222), .ZN(n8067) );
  NOR2_X1 U5332 ( .A1(n5089), .A2(n4536), .ZN(n6048) );
  AND2_X1 U5333 ( .A1(n7261), .A2(n7138), .ZN(n6649) );
  INV_X1 U5334 ( .A(n7776), .ZN(n6333) );
  NAND2_X1 U5335 ( .A1(n4972), .A2(n6332), .ZN(n4974) );
  AND2_X1 U5336 ( .A1(n5784), .A2(n5057), .ZN(n5056) );
  INV_X1 U5337 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5784) );
  INV_X1 U5338 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5057) );
  NOR2_X1 U5339 ( .A1(n5798), .A2(n4674), .ZN(n4671) );
  AND4_X1 U5340 ( .A1(n5840), .A2(n5848), .A3(n5854), .A4(n5772), .ZN(n5773)
         );
  INV_X1 U5341 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5772) );
  AND2_X1 U5342 ( .A1(n4969), .A2(n5056), .ZN(n4968) );
  INV_X1 U5343 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4969) );
  NOR2_X1 U5344 ( .A1(n7660), .A2(n7659), .ZN(n5077) );
  NAND2_X1 U5345 ( .A1(n4796), .A2(n5704), .ZN(n4793) );
  NOR2_X1 U5346 ( .A1(n9624), .A2(n4797), .ZN(n4795) );
  NOR2_X1 U5347 ( .A1(n5025), .A2(n9656), .ZN(n5024) );
  INV_X1 U5348 ( .A(n5026), .ZN(n5025) );
  AND2_X1 U5349 ( .A1(n9687), .A2(n4722), .ZN(n4721) );
  NAND2_X1 U5350 ( .A1(n4723), .A2(n9296), .ZN(n4722) );
  INV_X1 U5351 ( .A(n9372), .ZN(n4720) );
  NAND2_X1 U5352 ( .A1(n9690), .A2(n9171), .ZN(n9372) );
  NOR2_X1 U5353 ( .A1(n4519), .A2(n9715), .ZN(n9702) );
  AND2_X1 U5354 ( .A1(n9421), .A2(n4712), .ZN(n4711) );
  NAND2_X1 U5355 ( .A1(n9270), .A2(n9276), .ZN(n4712) );
  INV_X1 U5356 ( .A(n9276), .ZN(n4713) );
  INV_X1 U5357 ( .A(n7719), .ZN(n4805) );
  INV_X1 U5358 ( .A(n9347), .ZN(n5746) );
  INV_X1 U5359 ( .A(n9349), .ZN(n4705) );
  NOR2_X1 U5360 ( .A1(n4783), .A2(n4781), .ZN(n4780) );
  NAND2_X1 U5361 ( .A1(n9515), .A2(n10125), .ZN(n9391) );
  NAND2_X1 U5362 ( .A1(n5507), .A2(n9517), .ZN(n9385) );
  AOI21_X1 U5363 ( .B1(n9624), .B2(n9616), .A(n4716), .ZN(n4715) );
  INV_X1 U5364 ( .A(n9310), .ZN(n4716) );
  NAND2_X1 U5365 ( .A1(n5438), .A2(n4830), .ZN(n4829) );
  INV_X1 U5366 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4830) );
  NOR2_X1 U5367 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n5446) );
  NAND2_X1 U5368 ( .A1(n4834), .A2(n5405), .ZN(n5410) );
  AND2_X1 U5369 ( .A1(n5395), .A2(n5390), .ZN(n5393) );
  NAND2_X1 U5370 ( .A1(n4832), .A2(n5376), .ZN(n5384) );
  AND2_X1 U5371 ( .A1(n5385), .A2(n5380), .ZN(n5383) );
  AND2_X1 U5372 ( .A1(n4849), .A2(n4847), .ZN(n4846) );
  NAND2_X1 U5373 ( .A1(n4854), .A2(n4850), .ZN(n4849) );
  NAND2_X1 U5374 ( .A1(n4851), .A2(n4848), .ZN(n4847) );
  INV_X1 U5375 ( .A(n5333), .ZN(n4850) );
  INV_X1 U5376 ( .A(n5335), .ZN(n4845) );
  INV_X1 U5377 ( .A(n4867), .ZN(n4866) );
  OAI21_X1 U5378 ( .B1(n4504), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n4698), .ZN(
        n5133) );
  NAND2_X1 U5379 ( .A1(n4504), .A2(n4836), .ZN(n4698) );
  XNOR2_X1 U5380 ( .A(n7108), .B(n8284), .ZN(n7059) );
  AND2_X1 U5381 ( .A1(n4695), .A2(n4696), .ZN(n4694) );
  OR2_X1 U5382 ( .A1(n7057), .A2(n4966), .ZN(n7110) );
  OR2_X1 U5383 ( .A1(n6080), .A2(n6433), .ZN(n4627) );
  INV_X1 U5384 ( .A(n4966), .ZN(n4965) );
  AOI21_X1 U5385 ( .B1(n7154), .B2(n4964), .A(n5076), .ZN(n4963) );
  INV_X1 U5386 ( .A(n7109), .ZN(n4964) );
  NOR2_X1 U5387 ( .A1(n4956), .A2(n4953), .ZN(n4952) );
  NAND2_X1 U5388 ( .A1(n4677), .A2(n4679), .ZN(n4675) );
  INV_X1 U5389 ( .A(n8199), .ZN(n4953) );
  INV_X1 U5390 ( .A(n7840), .ZN(n4955) );
  NAND2_X1 U5391 ( .A1(n7424), .A2(n4682), .ZN(n7455) );
  OR2_X1 U5392 ( .A1(n7425), .A2(n7426), .ZN(n4682) );
  OAI21_X1 U5393 ( .B1(n6690), .B2(n4979), .A(n4978), .ZN(n6959) );
  NAND2_X1 U5394 ( .A1(n4977), .A2(n4976), .ZN(n4978) );
  NAND2_X1 U5395 ( .A1(n6703), .A2(n8286), .ZN(n4976) );
  AOI21_X1 U5396 ( .B1(n4960), .B2(n4962), .A(n4573), .ZN(n4958) );
  INV_X1 U5397 ( .A(n7821), .ZN(n4971) );
  INV_X1 U5398 ( .A(n4691), .ZN(n4690) );
  OAI21_X1 U5399 ( .B1(n4694), .B2(n4692), .A(n7752), .ZN(n4691) );
  NAND2_X1 U5400 ( .A1(n4690), .A2(n4692), .ZN(n4687) );
  OAI21_X1 U5401 ( .B1(n7747), .B2(n4692), .A(n4690), .ZN(n7822) );
  XNOR2_X1 U5402 ( .A(n5851), .B(n5850), .ZN(n6992) );
  AOI21_X1 U5403 ( .B1(n6992), .B2(P2_REG2_REG_3__SCAN_IN), .A(n5852), .ZN(
        n6967) );
  AND2_X1 U5404 ( .A1(n5851), .A2(n6999), .ZN(n5852) );
  XNOR2_X1 U5405 ( .A(n5865), .B(n10209), .ZN(n10211) );
  NAND2_X1 U5406 ( .A1(n10211), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n10210) );
  XNOR2_X1 U5407 ( .A(n5932), .B(n10209), .ZN(n10213) );
  NAND2_X1 U5408 ( .A1(n10213), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n10212) );
  NOR2_X1 U5409 ( .A1(n6875), .A2(n4872), .ZN(n10219) );
  NOR2_X1 U5410 ( .A1(n4874), .A2(n4873), .ZN(n4872) );
  INV_X1 U5411 ( .A(n5902), .ZN(n4874) );
  NOR2_X1 U5412 ( .A1(n10219), .A2(n10218), .ZN(n10217) );
  NAND2_X1 U5413 ( .A1(n10227), .A2(n10228), .ZN(n10226) );
  NAND2_X1 U5414 ( .A1(n10243), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n10242) );
  NAND2_X1 U5415 ( .A1(n10259), .A2(n10260), .ZN(n10258) );
  NAND2_X1 U5416 ( .A1(n10262), .A2(n10263), .ZN(n10261) );
  INV_X1 U5417 ( .A(n5906), .ZN(n4890) );
  INV_X1 U5418 ( .A(n4887), .ZN(n4886) );
  AOI21_X1 U5419 ( .B1(n10225), .B2(n5905), .A(n10234), .ZN(n10251) );
  NOR2_X1 U5420 ( .A1(n10251), .A2(n10250), .ZN(n10249) );
  XNOR2_X1 U5421 ( .A(n5936), .B(n10274), .ZN(n10278) );
  NAND2_X1 U5422 ( .A1(n10295), .A2(n10296), .ZN(n10294) );
  AOI21_X1 U5423 ( .B1(n4898), .B2(n10300), .A(n10315), .ZN(n4897) );
  AOI21_X1 U5424 ( .B1(n10274), .B2(n5910), .A(n10282), .ZN(n10301) );
  NOR2_X1 U5425 ( .A1(n10301), .A2(n10300), .ZN(n10299) );
  XNOR2_X1 U5426 ( .A(n5938), .B(n10307), .ZN(n10311) );
  NAND2_X1 U5427 ( .A1(n9948), .A2(n9949), .ZN(n9947) );
  NOR2_X1 U5428 ( .A1(n4908), .A2(n5920), .ZN(n4902) );
  OAI22_X1 U5429 ( .A1(n4905), .A2(n4907), .B1(n4906), .B2(n5920), .ZN(n4904)
         );
  OR2_X1 U5430 ( .A1(n10353), .A2(n10352), .ZN(n10350) );
  NOR2_X1 U5431 ( .A1(n5048), .A2(n8375), .ZN(n5055) );
  NOR2_X1 U5432 ( .A1(n8382), .A2(n4505), .ZN(n5048) );
  AND2_X1 U5433 ( .A1(n6220), .A2(n6219), .ZN(n7845) );
  AND2_X1 U5434 ( .A1(n8067), .A2(n8066), .ZN(n8384) );
  AND2_X1 U5435 ( .A1(n7941), .A2(n8055), .ZN(n8420) );
  AND4_X1 U5436 ( .A1(n6128), .A2(n6127), .A3(n6126), .A4(n6125), .ZN(n8020)
         );
  AND4_X1 U5437 ( .A1(n6119), .A2(n6118), .A3(n6117), .A4(n6116), .ZN(n7749)
         );
  INV_X1 U5438 ( .A(n8280), .ZN(n7457) );
  NOR2_X1 U5439 ( .A1(n7918), .A2(n5002), .ZN(n7191) );
  INV_X1 U5440 ( .A(n7949), .ZN(n5002) );
  OR2_X1 U5441 ( .A1(n6037), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6053) );
  INV_X1 U5442 ( .A(n4753), .ZN(n4752) );
  OAI21_X1 U5443 ( .B1(n7981), .B2(n4754), .A(n7984), .ZN(n4753) );
  INV_X1 U5444 ( .A(n7993), .ZN(n4754) );
  NAND2_X1 U5445 ( .A1(n6715), .A2(n5996), .ZN(n6584) );
  NOR2_X1 U5446 ( .A1(n7907), .A2(n4999), .ZN(n4998) );
  INV_X1 U5447 ( .A(n8082), .ZN(n4999) );
  OR2_X1 U5448 ( .A1(n8513), .A2(n8326), .ZN(n8082) );
  NAND2_X1 U5449 ( .A1(n8518), .A2(n8338), .ZN(n6239) );
  NOR2_X1 U5450 ( .A1(n8518), .A2(n8338), .ZN(n6238) );
  INV_X1 U5451 ( .A(n8348), .ZN(n6240) );
  INV_X1 U5452 ( .A(n8078), .ZN(n4761) );
  AND2_X1 U5453 ( .A1(n8084), .A2(n8078), .ZN(n8358) );
  INV_X1 U5454 ( .A(n8384), .ZN(n8382) );
  NOR2_X1 U5455 ( .A1(n6140), .A2(n5062), .ZN(n5061) );
  AND2_X1 U5456 ( .A1(n6303), .A2(n8029), .ZN(n8025) );
  INV_X1 U5457 ( .A(n8387), .ZN(n8430) );
  INV_X1 U5458 ( .A(n4987), .ZN(n4767) );
  NAND2_X1 U5459 ( .A1(n7098), .A2(n4768), .ZN(n4766) );
  INV_X1 U5460 ( .A(n6940), .ZN(n10383) );
  AND2_X1 U5461 ( .A1(n4559), .A2(n5967), .ZN(n5066) );
  AND3_X1 U5462 ( .A1(n5783), .A2(n4511), .A3(n4661), .ZN(n5795) );
  AND2_X1 U5463 ( .A1(n5782), .A2(n4880), .ZN(n4661) );
  AND2_X1 U5464 ( .A1(n5056), .A2(n5068), .ZN(n4880) );
  INV_X1 U5465 ( .A(n4671), .ZN(n4670) );
  AOI21_X1 U5466 ( .B1(n4949), .B2(n4674), .A(n4674), .ZN(n4947) );
  INV_X1 U5467 ( .A(n4950), .ZN(n4949) );
  INV_X1 U5468 ( .A(n4673), .ZN(n4672) );
  OAI21_X1 U5469 ( .B1(n5801), .B2(n4674), .A(n5798), .ZN(n4673) );
  INV_X1 U5470 ( .A(n5805), .ZN(n6293) );
  INV_X1 U5471 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5840) );
  INV_X1 U5472 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5848) );
  INV_X1 U5473 ( .A(n9517), .ZN(n6930) );
  XNOR2_X1 U5474 ( .A(n4598), .B(n8731), .ZN(n6639) );
  NAND2_X1 U5475 ( .A1(n4924), .A2(n7652), .ZN(n4920) );
  NAND2_X1 U5476 ( .A1(n4930), .A2(n9149), .ZN(n9152) );
  OR2_X1 U5477 ( .A1(n8620), .A2(n8619), .ZN(n8621) );
  NOR2_X1 U5478 ( .A1(n6543), .A2(n6850), .ZN(n6546) );
  AND4_X1 U5479 ( .A1(n5599), .A2(n5598), .A3(n5597), .A4(n5596), .ZN(n7708)
         );
  AND4_X1 U5480 ( .A1(n5573), .A2(n5572), .A3(n5571), .A4(n5570), .ZN(n7638)
         );
  AND4_X1 U5481 ( .A1(n5557), .A2(n5556), .A3(n5555), .A4(n5554), .ZN(n7516)
         );
  AND4_X1 U5482 ( .A1(n5550), .A2(n5549), .A3(n5548), .A4(n5547), .ZN(n7339)
         );
  NOR2_X1 U5483 ( .A1(n9996), .A2(n4525), .ZN(n9520) );
  OR2_X1 U5484 ( .A1(n9520), .A2(n9519), .ZN(n4929) );
  AND2_X1 U5485 ( .A1(n4929), .A2(n4928), .ZN(n10021) );
  NAND2_X1 U5486 ( .A1(n9525), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4928) );
  OR2_X1 U5487 ( .A1(n6796), .A2(n6795), .ZN(n4932) );
  NOR2_X1 U5488 ( .A1(n7766), .A2(n4581), .ZN(n9532) );
  OR2_X1 U5489 ( .A1(n9548), .A2(n9547), .ZN(n9555) );
  INV_X1 U5490 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4831) );
  AND2_X1 U5491 ( .A1(n9297), .A2(n9372), .ZN(n9687) );
  INV_X1 U5492 ( .A(n9694), .ZN(n4802) );
  NAND2_X1 U5493 ( .A1(n9696), .A2(n9697), .ZN(n9695) );
  INV_X1 U5494 ( .A(n9728), .ZN(n5650) );
  INV_X1 U5495 ( .A(n4824), .ZN(n4821) );
  AOI21_X1 U5496 ( .B1(n4513), .B2(n5630), .A(n4539), .ZN(n4824) );
  INV_X1 U5497 ( .A(n5600), .ZN(n4813) );
  NAND2_X1 U5498 ( .A1(n4707), .A2(n5746), .ZN(n4706) );
  INV_X1 U5499 ( .A(n7587), .ZN(n4707) );
  NAND2_X1 U5500 ( .A1(n9409), .A2(n9258), .ZN(n9347) );
  NAND2_X1 U5501 ( .A1(n7385), .A2(n5740), .ZN(n7386) );
  NOR2_X1 U5502 ( .A1(n5080), .A2(n7605), .ZN(n7406) );
  INV_X1 U5503 ( .A(n5140), .ZN(n5151) );
  INV_X1 U5504 ( .A(n9794), .ZN(n10063) );
  NAND2_X1 U5505 ( .A1(n5428), .A2(n5427), .ZN(n9458) );
  OR2_X1 U5506 ( .A1(n7164), .A2(n6545), .ZN(n10168) );
  INV_X1 U5507 ( .A(n4829), .ZN(n4828) );
  INV_X1 U5508 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5449) );
  NOR2_X1 U5509 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5120) );
  AND2_X1 U5510 ( .A1(n5112), .A2(n5164), .ZN(n4938) );
  NOR3_X1 U5511 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .A3(
        P1_IR_REG_18__SCAN_IN), .ZN(n5112) );
  OAI21_X1 U5512 ( .B1(n5275), .B2(n4520), .A(n4858), .ZN(n5307) );
  NAND2_X1 U5513 ( .A1(n4861), .A2(n5284), .ZN(n5298) );
  NAND2_X1 U5514 ( .A1(n5275), .A2(n4862), .ZN(n4861) );
  NAND2_X1 U5515 ( .A1(n5275), .A2(n5274), .ZN(n5286) );
  NAND2_X1 U5516 ( .A1(n4864), .A2(n4867), .ZN(n5256) );
  NAND2_X1 U5517 ( .A1(n5239), .A2(n4869), .ZN(n4864) );
  INV_X1 U5518 ( .A(n5182), .ZN(n4991) );
  INV_X1 U5519 ( .A(n5191), .ZN(n4992) );
  XNOR2_X1 U5520 ( .A(n5133), .B(SI_1_), .ZN(n5132) );
  OR3_X1 U5521 ( .A1(n6332), .A2(n7776), .A3(n6331), .ZN(n6374) );
  INV_X1 U5522 ( .A(n8289), .ZN(n6942) );
  AND4_X1 U5523 ( .A1(n6149), .A2(n6148), .A3(n6147), .A4(n6146), .ZN(n8179)
         );
  AND4_X1 U5524 ( .A1(n6160), .A2(n6159), .A3(n6158), .A4(n6157), .ZN(n8187)
         );
  NAND2_X1 U5525 ( .A1(n7157), .A2(n7156), .ZN(n7424) );
  AND3_X1 U5526 ( .A1(n5978), .A2(n5977), .A3(n5976), .ZN(n8202) );
  AND2_X1 U5527 ( .A1(n6609), .A2(n6608), .ZN(n8251) );
  INV_X1 U5528 ( .A(n8129), .ZN(n4649) );
  NOR2_X1 U5529 ( .A1(n4653), .A2(n4510), .ZN(n4647) );
  NAND2_X1 U5530 ( .A1(n4655), .A2(n4658), .ZN(n4653) );
  NAND2_X1 U5531 ( .A1(n6227), .A2(n6226), .ZN(n8369) );
  NAND2_X1 U5532 ( .A1(n6218), .A2(n6217), .ZN(n8273) );
  INV_X1 U5533 ( .A(n8179), .ZN(n8275) );
  INV_X1 U5534 ( .A(n7063), .ZN(n8285) );
  OAI21_X1 U5535 ( .B1(n6838), .B2(n6837), .A(n4877), .ZN(n6855) );
  OR2_X1 U5536 ( .A1(n5897), .A2(n6845), .ZN(n4877) );
  NOR2_X1 U5537 ( .A1(n5817), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5815) );
  OAI21_X1 U5538 ( .B1(n9949), .B2(n9948), .A(n9947), .ZN(n4605) );
  INV_X1 U5539 ( .A(n6993), .ZN(n10348) );
  NAND2_X1 U5540 ( .A1(n9951), .A2(n9950), .ZN(n4603) );
  OAI21_X1 U5541 ( .B1(n6326), .B2(n8387), .A(n6324), .ZN(n4770) );
  NAND2_X1 U5542 ( .A1(n6284), .A2(n6283), .ZN(n7815) );
  OAI21_X1 U5543 ( .B1(n6364), .B2(n8387), .A(n6363), .ZN(n8299) );
  NOR2_X1 U5544 ( .A1(n6362), .A2(n6361), .ZN(n6363) );
  NOR2_X1 U5545 ( .A1(n8327), .A2(n8391), .ZN(n6362) );
  NAND2_X1 U5546 ( .A1(n5980), .A2(n5979), .ZN(n8476) );
  AND2_X1 U5547 ( .A1(n6306), .A2(n8051), .ZN(n4769) );
  NAND2_X1 U5548 ( .A1(n7807), .A2(n6330), .ZN(n5047) );
  NAND2_X1 U5549 ( .A1(n5353), .A2(n5352), .ZN(n9703) );
  NOR2_X1 U5550 ( .A1(n7485), .A2(n7484), .ZN(n7766) );
  XNOR2_X1 U5551 ( .A(n9532), .B(n9542), .ZN(n7768) );
  NOR2_X1 U5552 ( .A1(n9991), .A2(n9987), .ZN(n10017) );
  OAI21_X1 U5553 ( .B1(n9596), .B2(n9595), .A(n4945), .ZN(n4944) );
  AOI21_X1 U5554 ( .B1(n9597), .B2(n10017), .A(n10025), .ZN(n4945) );
  AND3_X1 U5555 ( .A1(n5017), .A2(n5014), .A3(n5013), .ZN(n9602) );
  AOI21_X1 U5556 ( .B1(n5016), .B2(n9327), .A(n9794), .ZN(n5013) );
  NAND2_X1 U5557 ( .A1(n7793), .A2(n9327), .ZN(n5017) );
  NAND2_X1 U5558 ( .A1(n7784), .A2(n10054), .ZN(n7792) );
  OR2_X1 U5559 ( .A1(n7876), .A2(n8736), .ZN(n5083) );
  NAND2_X1 U5560 ( .A1(n9381), .A2(n5455), .ZN(n7164) );
  NOR2_X1 U5561 ( .A1(n7876), .A2(n9875), .ZN(n5769) );
  INV_X1 U5562 ( .A(n4732), .ZN(n4731) );
  INV_X1 U5563 ( .A(n6387), .ZN(n9929) );
  INV_X1 U5564 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5115) );
  INV_X1 U5565 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5328) );
  NAND2_X1 U5566 ( .A1(n4620), .A2(n8003), .ZN(n8009) );
  NAND2_X1 U5567 ( .A1(n4623), .A2(n4538), .ZN(n4620) );
  NAND2_X1 U5568 ( .A1(n4638), .A2(n8017), .ZN(n8024) );
  NAND2_X1 U5569 ( .A1(n8024), .A2(n5062), .ZN(n8027) );
  NOR2_X1 U5570 ( .A1(n4636), .A2(n4630), .ZN(n4629) );
  NAND2_X1 U5571 ( .A1(n4634), .A2(n4633), .ZN(n4630) );
  NAND2_X1 U5572 ( .A1(n9260), .A2(n9325), .ZN(n4595) );
  NAND2_X1 U5573 ( .A1(n4597), .A2(n9321), .ZN(n4596) );
  INV_X1 U5574 ( .A(n6711), .ZN(n6297) );
  OAI211_X1 U5575 ( .C1(n9277), .C2(n9274), .A(n9423), .B(n9330), .ZN(n9275)
         );
  NAND2_X1 U5576 ( .A1(n8443), .A2(n8498), .ZN(n7896) );
  OR2_X1 U5577 ( .A1(n8100), .A2(n8099), .ZN(n8103) );
  INV_X1 U5578 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5820) );
  INV_X1 U5579 ( .A(n4913), .ZN(n4912) );
  OAI21_X1 U5580 ( .B1(n5918), .B2(n5919), .A(n4914), .ZN(n4913) );
  NAND2_X1 U5581 ( .A1(n8448), .A2(n8272), .ZN(n5043) );
  INV_X1 U5582 ( .A(SI_16_), .ZN(n9064) );
  NOR2_X1 U5583 ( .A1(n9690), .A2(n9671), .ZN(n5026) );
  NOR2_X1 U5584 ( .A1(n7653), .A2(n7693), .ZN(n5032) );
  NAND2_X1 U5585 ( .A1(n4833), .A2(n5413), .ZN(n5417) );
  INV_X1 U5586 ( .A(n4853), .ZN(n4848) );
  INV_X1 U5587 ( .A(n5306), .ZN(n4857) );
  INV_X1 U5588 ( .A(SI_17_), .ZN(n5300) );
  INV_X1 U5589 ( .A(SI_11_), .ZN(n9066) );
  AND2_X1 U5590 ( .A1(n7829), .A2(n4681), .ZN(n4680) );
  NAND2_X1 U5591 ( .A1(n4514), .A2(n7826), .ZN(n4681) );
  INV_X1 U5592 ( .A(n8159), .ZN(n4956) );
  INV_X1 U5593 ( .A(n6957), .ZN(n4975) );
  OAI21_X1 U5594 ( .B1(n6703), .B2(n8286), .A(n4980), .ZN(n4977) );
  INV_X1 U5595 ( .A(n4961), .ZN(n4960) );
  OAI21_X1 U5596 ( .B1(n8192), .B2(n4962), .A(n8166), .ZN(n4961) );
  INV_X1 U5597 ( .A(n7851), .ZN(n4962) );
  OR2_X1 U5598 ( .A1(n8103), .A2(n8102), .ZN(n8113) );
  NAND2_X1 U5599 ( .A1(n4744), .A2(n4743), .ZN(n5928) );
  NAND2_X1 U5600 ( .A1(n6973), .A2(n4748), .ZN(n4743) );
  INV_X1 U5601 ( .A(n4607), .ZN(n5856) );
  NAND2_X1 U5602 ( .A1(n7087), .A2(n5931), .ZN(n6880) );
  NAND2_X1 U5603 ( .A1(n10291), .A2(n5877), .ZN(n5878) );
  NAND2_X1 U5604 ( .A1(n10326), .A2(n4734), .ZN(n5940) );
  OR2_X1 U5605 ( .A1(n10322), .A2(n7680), .ZN(n4734) );
  NOR2_X1 U5606 ( .A1(n4911), .A2(n4910), .ZN(n4909) );
  INV_X1 U5607 ( .A(n5919), .ZN(n4910) );
  INV_X1 U5608 ( .A(n5918), .ZN(n4911) );
  NAND2_X1 U5609 ( .A1(n4912), .A2(n5919), .ZN(n4906) );
  NOR2_X1 U5610 ( .A1(n6181), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6190) );
  OR2_X1 U5611 ( .A1(n6179), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6181) );
  OR2_X1 U5612 ( .A1(n8435), .A2(n8154), .ZN(n7928) );
  NOR2_X1 U5613 ( .A1(n6144), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6143) );
  AND2_X1 U5614 ( .A1(n6052), .A2(n5962), .ZN(n6066) );
  NOR2_X1 U5615 ( .A1(n8420), .A2(n5072), .ZN(n5071) );
  INV_X1 U5616 ( .A(n5063), .ZN(n5059) );
  NOR2_X1 U5617 ( .A1(n6373), .A2(n6378), .ZN(n6615) );
  INV_X1 U5618 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5967) );
  INV_X1 U5619 ( .A(n5780), .ZN(n4776) );
  OAI21_X1 U5620 ( .B1(n5785), .B2(n4674), .A(n5786), .ZN(n4950) );
  NOR2_X1 U5621 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(n5780), .ZN(n4685) );
  AND2_X1 U5622 ( .A1(n4777), .A2(n5773), .ZN(n4686) );
  INV_X1 U5623 ( .A(n7635), .ZN(n4925) );
  INV_X1 U5624 ( .A(n9441), .ZN(n9454) );
  NAND2_X1 U5625 ( .A1(n9367), .A2(n4837), .ZN(n9441) );
  NAND2_X1 U5626 ( .A1(n9458), .A2(n9371), .ZN(n4837) );
  AND2_X1 U5627 ( .A1(n5455), .A2(n9598), .ZN(n9321) );
  INV_X1 U5628 ( .A(n6538), .ZN(n9463) );
  INV_X1 U5629 ( .A(n5686), .ZN(n4788) );
  NAND2_X1 U5630 ( .A1(n4552), .A2(n10034), .ZN(n9396) );
  NAND2_X1 U5631 ( .A1(n9678), .A2(n5026), .ZN(n9669) );
  NOR2_X1 U5632 ( .A1(n9748), .A2(n5008), .ZN(n5007) );
  INV_X1 U5633 ( .A(n5009), .ZN(n5008) );
  NAND2_X1 U5634 ( .A1(n7442), .A2(n5032), .ZN(n7589) );
  NAND2_X1 U5635 ( .A1(n5468), .A2(n5466), .ZN(n5475) );
  AND2_X1 U5636 ( .A1(n5405), .A2(n5400), .ZN(n5403) );
  NAND2_X1 U5637 ( .A1(n5367), .A2(n5366), .ZN(n5375) );
  AND2_X1 U5638 ( .A1(n5376), .A2(n5371), .ZN(n5374) );
  AOI21_X1 U5639 ( .B1(n4841), .B2(n4842), .A(n4578), .ZN(n4840) );
  NAND2_X1 U5640 ( .A1(n5335), .A2(n4842), .ZN(n4839) );
  INV_X1 U5641 ( .A(SI_19_), .ZN(n5321) );
  INV_X1 U5642 ( .A(n5284), .ZN(n4860) );
  INV_X1 U5643 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5109) );
  NOR2_X1 U5644 ( .A1(n5285), .A2(n4863), .ZN(n4862) );
  INV_X1 U5645 ( .A(n5274), .ZN(n4863) );
  AOI21_X1 U5646 ( .B1(n4869), .B2(n5238), .A(n4546), .ZN(n4867) );
  OAI21_X1 U5647 ( .B1(n4500), .B2(P1_DATAO_REG_3__SCAN_IN), .A(n5148), .ZN(
        n5156) );
  NAND2_X1 U5648 ( .A1(n4500), .A2(n6427), .ZN(n5148) );
  OAI21_X1 U5649 ( .B1(n4498), .B2(n4589), .A(n4588), .ZN(n5145) );
  NAND2_X1 U5650 ( .A1(n4497), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4588) );
  NAND2_X1 U5651 ( .A1(n4665), .A2(n6650), .ZN(n4664) );
  NAND2_X1 U5652 ( .A1(n6647), .A2(n6648), .ZN(n4665) );
  OR2_X1 U5653 ( .A1(n6211), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6221) );
  AND2_X1 U5654 ( .A1(n8010), .A2(n8006), .ZN(n7922) );
  XNOR2_X1 U5655 ( .A(n6653), .B(n10383), .ZN(n6655) );
  AND2_X1 U5656 ( .A1(n6626), .A2(n6625), .ZN(n6696) );
  INV_X1 U5657 ( .A(n7138), .ZN(n4658) );
  AND4_X1 U5658 ( .A1(n7906), .A2(n6289), .A3(n6288), .A4(n6287), .ZN(n7861)
         );
  INV_X1 U5659 ( .A(n5995), .ZN(n6613) );
  OAI22_X1 U5660 ( .A1(n7030), .A2(n7031), .B1(n5893), .B2(n5892), .ZN(n6990)
         );
  NOR2_X1 U5661 ( .A1(n6967), .A2(n6968), .ZN(n6966) );
  NOR2_X1 U5662 ( .A1(n6990), .A2(n6991), .ZN(n6989) );
  INV_X1 U5663 ( .A(n6973), .ZN(n4747) );
  NAND2_X1 U5664 ( .A1(n4745), .A2(n4749), .ZN(n4746) );
  XNOR2_X1 U5665 ( .A(n5928), .B(n6845), .ZN(n6839) );
  XNOR2_X1 U5666 ( .A(n4607), .B(n6437), .ZN(n6840) );
  NOR3_X1 U5667 ( .A1(n6989), .A2(n6979), .A3(n6978), .ZN(n6977) );
  XNOR2_X1 U5668 ( .A(n5930), .B(n6060), .ZN(n7088) );
  NAND2_X1 U5669 ( .A1(n7088), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7087) );
  NOR2_X1 U5670 ( .A1(n6876), .A2(n6877), .ZN(n6875) );
  NOR2_X1 U5671 ( .A1(n5901), .A2(n7081), .ZN(n6876) );
  OAI21_X1 U5672 ( .B1(n6869), .B2(n7006), .A(n6860), .ZN(n5860) );
  NAND2_X1 U5673 ( .A1(n7090), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7089) );
  INV_X1 U5674 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7158) );
  AND2_X1 U5675 ( .A1(n5903), .A2(n10209), .ZN(n4871) );
  NAND2_X1 U5676 ( .A1(n10210), .A2(n5866), .ZN(n10227) );
  NAND2_X1 U5677 ( .A1(n10212), .A2(n5933), .ZN(n10230) );
  NAND2_X1 U5678 ( .A1(n10242), .A2(n5873), .ZN(n10259) );
  NAND2_X1 U5679 ( .A1(n10244), .A2(n5935), .ZN(n10262) );
  INV_X1 U5680 ( .A(n4885), .ZN(n4882) );
  NOR2_X1 U5681 ( .A1(n10251), .A2(n4886), .ZN(n4883) );
  AOI21_X1 U5682 ( .B1(n4887), .B2(n4889), .A(n4583), .ZN(n4885) );
  INV_X1 U5683 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8206) );
  NAND2_X1 U5684 ( .A1(n10275), .A2(n5876), .ZN(n10292) );
  NAND2_X1 U5685 ( .A1(n10292), .A2(n10293), .ZN(n10291) );
  NAND2_X1 U5686 ( .A1(n10277), .A2(n5937), .ZN(n10295) );
  XNOR2_X1 U5687 ( .A(n5878), .B(n10307), .ZN(n10309) );
  NAND2_X1 U5688 ( .A1(n10310), .A2(n5939), .ZN(n10327) );
  NAND2_X1 U5689 ( .A1(n10327), .A2(n10328), .ZN(n10326) );
  NAND2_X1 U5690 ( .A1(n4894), .A2(n4899), .ZN(n4893) );
  INV_X1 U5691 ( .A(n4897), .ZN(n4894) );
  XNOR2_X1 U5692 ( .A(n5940), .B(n10341), .ZN(n10345) );
  NAND2_X1 U5693 ( .A1(n10343), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n10342) );
  OR2_X1 U5694 ( .A1(n8293), .A2(n8292), .ZN(n8441) );
  NAND2_X1 U5695 ( .A1(n6367), .A2(n6311), .ZN(n7898) );
  OAI21_X1 U5696 ( .B1(n8324), .B2(n5038), .A(n5035), .ZN(n6290) );
  NAND2_X1 U5697 ( .A1(n5040), .A2(n5039), .ZN(n5038) );
  AOI21_X1 U5698 ( .B1(n5040), .B2(n5037), .A(n5036), .ZN(n5035) );
  NAND2_X1 U5699 ( .A1(n5034), .A2(n5040), .ZN(n6360) );
  NAND2_X1 U5700 ( .A1(n8324), .A2(n4521), .ZN(n5034) );
  NOR2_X1 U5701 ( .A1(n7861), .A2(n8389), .ZN(n6361) );
  AND2_X1 U5702 ( .A1(n6244), .A2(n6243), .ZN(n6256) );
  OR2_X1 U5703 ( .A1(n6133), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6144) );
  AND4_X1 U5704 ( .A1(n6107), .A2(n6106), .A3(n6105), .A4(n6104), .ZN(n7558)
         );
  OR2_X1 U5705 ( .A1(n6102), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6114) );
  INV_X1 U5706 ( .A(n7922), .ZN(n7183) );
  AND2_X1 U5707 ( .A1(n5090), .A2(n6089), .ZN(n5064) );
  AND2_X1 U5708 ( .A1(n8004), .A2(n7950), .ZN(n7921) );
  NAND2_X1 U5709 ( .A1(n5065), .A2(n6089), .ZN(n7144) );
  NAND2_X1 U5710 ( .A1(n6078), .A2(n6077), .ZN(n7196) );
  NAND2_X1 U5711 ( .A1(n4752), .A2(n4754), .ZN(n4750) );
  OR2_X1 U5712 ( .A1(n6692), .A2(n7017), .ZN(n6579) );
  NAND2_X1 U5713 ( .A1(n6374), .A2(n6627), .ZN(n6623) );
  NAND2_X1 U5714 ( .A1(n6584), .A2(n6585), .ZN(n7013) );
  NOR2_X1 U5715 ( .A1(n8118), .A2(n7138), .ZN(n6714) );
  NAND2_X1 U5716 ( .A1(n6711), .A2(n6716), .ZN(n6715) );
  OR2_X1 U5717 ( .A1(n6717), .A2(n6654), .ZN(n6716) );
  OR2_X1 U5718 ( .A1(n6378), .A2(n6351), .ZN(n6663) );
  OR2_X1 U5719 ( .A1(n6667), .A2(n6665), .ZN(n6373) );
  AND2_X1 U5720 ( .A1(n6252), .A2(n6251), .ZN(n8326) );
  AND2_X1 U5721 ( .A1(n6375), .A2(n6295), .ZN(n8387) );
  INV_X1 U5722 ( .A(n8089), .ZN(n8323) );
  AOI21_X1 U5723 ( .B1(n4760), .B2(n4758), .A(n4757), .ZN(n4756) );
  INV_X1 U5724 ( .A(n8083), .ZN(n4757) );
  AND2_X1 U5725 ( .A1(n8082), .A2(n8091), .ZN(n8335) );
  INV_X1 U5726 ( .A(n6228), .ZN(n5053) );
  NAND2_X1 U5727 ( .A1(n8477), .A2(n5000), .ZN(n8381) );
  NOR2_X1 U5728 ( .A1(n5001), .A2(n7942), .ZN(n5000) );
  INV_X1 U5729 ( .A(n4567), .ZN(n5001) );
  AND2_X1 U5730 ( .A1(n8041), .A2(n8038), .ZN(n8037) );
  AND2_X1 U5731 ( .A1(n8022), .A2(n8023), .ZN(n7925) );
  OAI211_X1 U5732 ( .C1(n6322), .C2(n7036), .A(n6002), .B(n6001), .ZN(n6658)
         );
  NAND2_X1 U5733 ( .A1(n8112), .A2(n6649), .ZN(n6675) );
  NOR2_X1 U5734 ( .A1(n6624), .A2(n6623), .ZN(n6610) );
  NAND2_X1 U5735 ( .A1(n4974), .A2(n6333), .ZN(n6452) );
  XNOR2_X1 U5736 ( .A(n5803), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8128) );
  XNOR2_X1 U5737 ( .A(n5884), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8124) );
  INV_X1 U5738 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5854) );
  NOR2_X1 U5739 ( .A1(n5601), .A2(n8683), .ZN(n5609) );
  OR2_X1 U5740 ( .A1(n5552), .A2(n7521), .ZN(n5559) );
  INV_X1 U5741 ( .A(n7040), .ZN(n6531) );
  INV_X1 U5742 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5584) );
  OR2_X1 U5743 ( .A1(n5615), .A2(n8773), .ZN(n5624) );
  XNOR2_X1 U5744 ( .A(n7518), .B(n7517), .ZN(n7631) );
  AOI222_X1 U5745 ( .A1(n6533), .A2(n8653), .B1(n7172), .B2(n8655), .C1(
        P1_IR_REG_0__SCAN_IN), .C2(n6532), .ZN(n6631) );
  AND2_X1 U5746 ( .A1(n5454), .A2(n9463), .ZN(n9184) );
  OAI21_X1 U5747 ( .B1(n7637), .B2(n4921), .A(n4919), .ZN(n4922) );
  OR2_X1 U5748 ( .A1(n5585), .A2(n5584), .ZN(n5594) );
  INV_X1 U5749 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5593) );
  OR2_X1 U5750 ( .A1(n5594), .A2(n5593), .ZN(n5601) );
  AND2_X1 U5751 ( .A1(n6770), .A2(n6922), .ZN(n6772) );
  AND2_X1 U5752 ( .A1(n5631), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5637) );
  NOR2_X1 U5753 ( .A1(n8590), .A2(n9135), .ZN(n5086) );
  AND2_X1 U5754 ( .A1(n10005), .A2(n9463), .ZN(n9197) );
  AND4_X1 U5755 ( .A1(n5712), .A2(n5711), .A3(n5710), .A4(n5709), .ZN(n9196)
         );
  AND4_X1 U5756 ( .A1(n5590), .A2(n5589), .A3(n5588), .A4(n5587), .ZN(n7655)
         );
  AND4_X1 U5757 ( .A1(n5564), .A2(n5563), .A3(n5562), .A4(n5561), .ZN(n7597)
         );
  AND4_X1 U5758 ( .A1(n5542), .A2(n5541), .A3(n5540), .A4(n5539), .ZN(n7246)
         );
  AND4_X1 U5759 ( .A1(n5533), .A2(n5532), .A3(n5531), .A4(n5530), .ZN(n7326)
         );
  AND4_X1 U5760 ( .A1(n5523), .A2(n5522), .A3(n5521), .A4(n5520), .ZN(n5524)
         );
  AND4_X1 U5761 ( .A1(n5514), .A2(n5513), .A3(n5512), .A4(n5511), .ZN(n6919)
         );
  NOR2_X1 U5762 ( .A1(n10001), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4615) );
  NAND2_X1 U5763 ( .A1(n10001), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4616) );
  NAND2_X1 U5764 ( .A1(n10013), .A2(n10014), .ZN(n10012) );
  OR2_X1 U5765 ( .A1(n6811), .A2(n6810), .ZN(n4613) );
  AND2_X1 U5766 ( .A1(n4613), .A2(n4612), .ZN(n6562) );
  NAND2_X1 U5767 ( .A1(n6812), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n4612) );
  NAND2_X1 U5768 ( .A1(n6562), .A2(n6563), .ZN(n6784) );
  NOR2_X1 U5769 ( .A1(n7125), .A2(n7124), .ZN(n7127) );
  NAND2_X1 U5770 ( .A1(n7127), .A2(n7126), .ZN(n7373) );
  NOR2_X1 U5771 ( .A1(n7763), .A2(n4582), .ZN(n9543) );
  AND2_X1 U5772 ( .A1(n9555), .A2(n9554), .ZN(n9556) );
  NAND2_X1 U5773 ( .A1(n9560), .A2(n4584), .ZN(n9562) );
  NAND2_X1 U5774 ( .A1(n9562), .A2(n9563), .ZN(n9573) );
  NAND2_X1 U5775 ( .A1(n9556), .A2(n9557), .ZN(n9580) );
  NOR2_X1 U5776 ( .A1(n9327), .A2(n5016), .ZN(n5015) );
  INV_X1 U5777 ( .A(n7793), .ZN(n5019) );
  INV_X1 U5778 ( .A(n9197), .ZN(n9141) );
  INV_X1 U5779 ( .A(n4792), .ZN(n4791) );
  OAI21_X1 U5780 ( .B1(n9624), .B2(n4793), .A(n5713), .ZN(n4792) );
  NAND2_X1 U5781 ( .A1(n4714), .A2(n9624), .ZN(n9615) );
  NOR2_X1 U5782 ( .A1(n9639), .A2(n5023), .ZN(n5022) );
  INV_X1 U5783 ( .A(n5024), .ZN(n5023) );
  AND2_X1 U5784 ( .A1(n9309), .A2(n9222), .ZN(n9633) );
  AOI21_X1 U5785 ( .B1(n4507), .B2(n4800), .A(n4540), .ZN(n4799) );
  INV_X1 U5786 ( .A(n5094), .ZN(n4800) );
  INV_X1 U5787 ( .A(n9663), .ZN(n5752) );
  AOI21_X1 U5788 ( .B1(n4721), .B2(n4724), .A(n4720), .ZN(n4719) );
  INV_X1 U5789 ( .A(n9296), .ZN(n4724) );
  NAND2_X1 U5790 ( .A1(n4815), .A2(n4541), .ZN(n9726) );
  NAND2_X1 U5791 ( .A1(n4816), .A2(n4817), .ZN(n4814) );
  AND2_X1 U5792 ( .A1(n9288), .A2(n9286), .ZN(n9728) );
  AOI21_X1 U5793 ( .B1(n4711), .B2(n4713), .A(n4709), .ZN(n4708) );
  INV_X1 U5794 ( .A(n9330), .ZN(n4709) );
  NAND2_X1 U5795 ( .A1(n9772), .A2(n9276), .ZN(n9757) );
  NAND2_X1 U5796 ( .A1(n9791), .A2(n9416), .ZN(n9772) );
  NAND2_X1 U5797 ( .A1(n5295), .A2(n5011), .ZN(n9778) );
  AOI21_X1 U5798 ( .B1(n4506), .B2(n4812), .A(n4579), .ZN(n4804) );
  INV_X1 U5799 ( .A(n4701), .ZN(n4700) );
  NAND2_X1 U5800 ( .A1(n7587), .A2(n4704), .ZN(n4702) );
  AND2_X1 U5801 ( .A1(n7442), .A2(n5028), .ZN(n7726) );
  NOR2_X1 U5802 ( .A1(n9263), .A2(n5030), .ZN(n5028) );
  OR2_X1 U5803 ( .A1(n9794), .A2(n9720), .ZN(n6548) );
  NAND2_X1 U5804 ( .A1(n9402), .A2(n9399), .ZN(n9342) );
  AND2_X1 U5805 ( .A1(n5216), .A2(n4561), .ZN(n4733) );
  AOI21_X1 U5806 ( .B1(n7344), .B2(n4785), .A(n4544), .ZN(n4784) );
  INV_X1 U5807 ( .A(n5551), .ZN(n4785) );
  AND2_X1 U5808 ( .A1(n5176), .A2(n5006), .ZN(n5005) );
  NAND2_X1 U5809 ( .A1(n4570), .A2(n5176), .ZN(n10046) );
  AND2_X1 U5810 ( .A1(n5176), .A2(n4515), .ZN(n10047) );
  NAND2_X1 U5811 ( .A1(n10034), .A2(n9223), .ZN(n7356) );
  NAND2_X1 U5812 ( .A1(n5176), .A2(n10132), .ZN(n7357) );
  NAND2_X1 U5813 ( .A1(n9394), .A2(n9397), .ZN(n9335) );
  NAND2_X1 U5814 ( .A1(n9393), .A2(n9391), .ZN(n9334) );
  NAND2_X1 U5815 ( .A1(n5382), .A2(n5381), .ZN(n9656) );
  NAND2_X1 U5816 ( .A1(n5294), .A2(n5293), .ZN(n9796) );
  INV_X1 U5817 ( .A(n7605), .ZN(n10161) );
  AND2_X1 U5818 ( .A1(n6537), .A2(n6540), .ZN(n7168) );
  AND3_X1 U5819 ( .A1(n6534), .A2(n6535), .A3(n6548), .ZN(n5957) );
  INV_X1 U5820 ( .A(n7172), .ZN(n7275) );
  INV_X1 U5821 ( .A(n9815), .ZN(n10172) );
  NAND2_X1 U5822 ( .A1(n4946), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5460) );
  NAND2_X1 U5823 ( .A1(n5463), .A2(n5114), .ZN(n4946) );
  OAI21_X1 U5824 ( .B1(n5356), .B2(n5355), .A(n5354), .ZN(n5362) );
  XNOR2_X1 U5825 ( .A(n5473), .B(n5472), .ZN(n7576) );
  INV_X1 U5826 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U5827 ( .A1(n4844), .A2(n4846), .ZN(n5347) );
  NAND2_X1 U5828 ( .A1(n4845), .A2(n4523), .ZN(n4844) );
  INV_X1 U5829 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5325) );
  OR2_X1 U5830 ( .A1(n5217), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5234) );
  INV_X1 U5831 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5105) );
  NAND2_X1 U5832 ( .A1(n5136), .A2(n5135), .ZN(n5144) );
  XNOR2_X1 U5833 ( .A(n5128), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6422) );
  NOR2_X1 U5834 ( .A1(n7057), .A2(n7056), .ZN(n7060) );
  AOI21_X1 U5835 ( .B1(n8330), .B2(n6266), .A(n6260), .ZN(n8316) );
  NAND2_X1 U5836 ( .A1(n4689), .A2(n4693), .ZN(n7753) );
  NAND2_X1 U5837 ( .A1(n7747), .A2(n4694), .ZN(n4689) );
  OR2_X1 U5838 ( .A1(n8132), .A2(n8131), .ZN(n8133) );
  NAND2_X1 U5839 ( .A1(n7110), .A2(n7109), .ZN(n7155) );
  XNOR2_X1 U5840 ( .A(n6655), .B(n6652), .ZN(n6938) );
  NAND2_X1 U5841 ( .A1(n8198), .A2(n8199), .ZN(n4957) );
  NAND2_X1 U5842 ( .A1(n8191), .A2(n8192), .ZN(n4959) );
  AND4_X1 U5843 ( .A1(n6028), .A2(n6027), .A3(n6026), .A4(n6025), .ZN(n7063)
         );
  AND2_X1 U5844 ( .A1(n6704), .A2(n6703), .ZN(n6958) );
  INV_X1 U5845 ( .A(n8369), .ZN(n8221) );
  NAND2_X1 U5846 ( .A1(n6020), .A2(n4626), .ZN(n6694) );
  AND2_X1 U5847 ( .A1(n4627), .A2(n4531), .ZN(n4626) );
  AOI21_X1 U5848 ( .B1(n4535), .B2(n4684), .A(n4683), .ZN(n7157) );
  INV_X1 U5849 ( .A(n4963), .ZN(n4683) );
  INV_X1 U5850 ( .A(n7057), .ZN(n4684) );
  AND2_X1 U5851 ( .A1(n6657), .A2(n6612), .ZN(n8257) );
  NAND2_X1 U5852 ( .A1(n7747), .A2(n4696), .ZN(n8213) );
  NAND2_X1 U5853 ( .A1(n4951), .A2(n4954), .ZN(n8219) );
  AOI21_X1 U5854 ( .B1(n8159), .B2(n4955), .A(n4572), .ZN(n4954) );
  NAND2_X1 U5855 ( .A1(n4676), .A2(n4537), .ZN(n4951) );
  AOI22_X1 U5856 ( .A1(n7459), .A2(n7458), .B1(n7457), .B2(n7456), .ZN(n7460)
         );
  AND3_X1 U5857 ( .A1(n6172), .A2(n6171), .A3(n6170), .ZN(n8235) );
  INV_X1 U5858 ( .A(n8244), .ZN(n8260) );
  AND2_X1 U5859 ( .A1(n6696), .A2(n8130), .ZN(n8210) );
  INV_X1 U5860 ( .A(n8257), .ZN(n8246) );
  NAND2_X1 U5861 ( .A1(n4688), .A2(n4575), .ZN(n8254) );
  NOR2_X1 U5862 ( .A1(n8252), .A2(n4971), .ZN(n4970) );
  NAND2_X1 U5863 ( .A1(n7822), .A2(n7821), .ZN(n8253) );
  INV_X1 U5864 ( .A(n8210), .ZN(n8262) );
  INV_X1 U5865 ( .A(n8326), .ZN(n8350) );
  INV_X1 U5866 ( .A(P2_U3893), .ZN(n9946) );
  INV_X1 U5867 ( .A(n8154), .ZN(n8412) );
  INV_X1 U5868 ( .A(n8235), .ZN(n8428) );
  INV_X1 U5869 ( .A(n9946), .ZN(n8283) );
  NAND4_X1 U5870 ( .A1(n6019), .A2(n6018), .A3(n6017), .A4(n6016), .ZN(n8287)
         );
  AND2_X1 U5871 ( .A1(n5998), .A2(n5997), .ZN(n5999) );
  CLKBUF_X1 U5872 ( .A(n6613), .Z(n6652) );
  INV_X1 U5873 ( .A(n10340), .ZN(n9945) );
  INV_X1 U5874 ( .A(n4746), .ZN(n6972) );
  AND2_X1 U5875 ( .A1(n4876), .A2(n4875), .ZN(n7083) );
  NAND2_X1 U5876 ( .A1(n5898), .A2(n6869), .ZN(n4875) );
  NOR2_X1 U5877 ( .A1(n6873), .A2(n6874), .ZN(n6872) );
  AND2_X1 U5878 ( .A1(n7089), .A2(n4610), .ZN(n6873) );
  NAND2_X1 U5879 ( .A1(n5860), .A2(n7084), .ZN(n4610) );
  NOR2_X1 U5880 ( .A1(n10249), .A2(n4889), .ZN(n10268) );
  NOR2_X1 U5881 ( .A1(n10299), .A2(n4900), .ZN(n10316) );
  NAND2_X1 U5882 ( .A1(n10301), .A2(n4898), .ZN(n4892) );
  INV_X1 U5883 ( .A(n10200), .ZN(n10339) );
  NAND2_X1 U5884 ( .A1(n9947), .A2(n4586), .ZN(n4738) );
  AND2_X1 U5885 ( .A1(n5946), .A2(n5948), .ZN(n10347) );
  INV_X1 U5886 ( .A(n4904), .ZN(n4903) );
  OR2_X1 U5887 ( .A1(n6890), .A2(n5948), .ZN(n6993) );
  XNOR2_X1 U5888 ( .A(n7898), .B(n6312), .ZN(n7812) );
  NAND2_X1 U5889 ( .A1(n6254), .A2(n6253), .ZN(n8331) );
  INV_X1 U5890 ( .A(n7845), .ZN(n8460) );
  AOI21_X1 U5891 ( .B1(n8385), .B2(n8382), .A(n4505), .ZN(n8368) );
  NAND2_X1 U5892 ( .A1(n6165), .A2(n6164), .ZN(n8491) );
  INV_X1 U5893 ( .A(n10419), .ZN(n7432) );
  INV_X1 U5894 ( .A(n7918), .ZN(n7194) );
  OAI21_X1 U5895 ( .B1(n6576), .B2(n4754), .A(n4752), .ZN(n7004) );
  INV_X1 U5896 ( .A(n10390), .ZN(n7017) );
  INV_X1 U5897 ( .A(n8407), .ZN(n8438) );
  INV_X1 U5898 ( .A(n6658), .ZN(n10371) );
  OR2_X1 U5899 ( .A1(n10418), .A2(n6714), .ZN(n10370) );
  AND2_X1 U5900 ( .A1(n6672), .A2(n10373), .ZN(n10381) );
  NAND2_X1 U5901 ( .A1(n5097), .A2(n4772), .ZN(n6940) );
  OR2_X1 U5902 ( .A1(n6322), .A2(n10193), .ZN(n5097) );
  NOR2_X1 U5903 ( .A1(n6672), .A2(n10370), .ZN(n8419) );
  INV_X1 U5904 ( .A(n10373), .ZN(n8404) );
  CLKBUF_X1 U5905 ( .A(n8419), .Z(n8434) );
  AND2_X1 U5906 ( .A1(n8303), .A2(n10429), .ZN(n6365) );
  NAND2_X1 U5907 ( .A1(n6242), .A2(n6241), .ZN(n8513) );
  OAI21_X1 U5908 ( .B1(n8376), .B2(n4763), .A(n4760), .ZN(n8347) );
  NAND2_X1 U5909 ( .A1(n8377), .A2(n8071), .ZN(n8357) );
  NAND2_X1 U5910 ( .A1(n8477), .A2(n7941), .ZN(n8398) );
  NAND2_X1 U5911 ( .A1(n6153), .A2(n6152), .ZN(n8181) );
  NAND2_X1 U5912 ( .A1(n6142), .A2(n6141), .ZN(n8250) );
  NAND2_X1 U5913 ( .A1(n5060), .A2(n5063), .ZN(n7529) );
  NAND2_X1 U5914 ( .A1(n6132), .A2(n6131), .ZN(n7751) );
  NAND2_X1 U5915 ( .A1(n6130), .A2(n8023), .ZN(n7545) );
  NAND2_X1 U5916 ( .A1(n6122), .A2(n6121), .ZN(n8217) );
  INV_X1 U5917 ( .A(n8507), .ZN(n8533) );
  AND2_X1 U5918 ( .A1(n4767), .A2(n4766), .ZN(n7251) );
  OR2_X1 U5919 ( .A1(n10432), .A2(n10418), .ZN(n8507) );
  AND2_X1 U5920 ( .A1(n5951), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6627) );
  INV_X1 U5921 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5971) );
  NAND2_X1 U5922 ( .A1(n5797), .A2(n5796), .ZN(n7776) );
  INV_X1 U5923 ( .A(n5795), .ZN(n5796) );
  NAND2_X1 U5924 ( .A1(n5799), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5788) );
  NAND2_X1 U5925 ( .A1(n4668), .A2(n4672), .ZN(n5799) );
  INV_X1 U5926 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7673) );
  AOI21_X1 U5927 ( .B1(n4672), .B2(n4674), .A(n4577), .ZN(n4669) );
  OR2_X1 U5928 ( .A1(n5800), .A2(n4670), .ZN(n4667) );
  INV_X1 U5929 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7384) );
  NAND2_X1 U5930 ( .A1(n5804), .A2(n5807), .ZN(n7963) );
  INV_X1 U5931 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8894) );
  INV_X1 U5932 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8883) );
  INV_X1 U5933 ( .A(n8124), .ZN(n7138) );
  INV_X1 U5934 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6836) );
  INV_X1 U5935 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6833) );
  INV_X1 U5936 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n9103) );
  INV_X1 U5937 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6524) );
  INV_X1 U5938 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6484) );
  INV_X1 U5939 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9062) );
  NAND2_X1 U5940 ( .A1(n5836), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5849) );
  NAND2_X1 U5941 ( .A1(n4551), .A2(n4591), .ZN(n4590) );
  INV_X1 U5942 ( .A(n8746), .ZN(n4591) );
  INV_X1 U5943 ( .A(n4920), .ZN(n4923) );
  NAND2_X1 U5944 ( .A1(n7044), .A2(n7043), .ZN(n7212) );
  OAI211_X1 U5945 ( .C1(n5151), .C2(n6428), .A(n5161), .B(n5160), .ZN(n7314)
         );
  INV_X1 U5946 ( .A(n9970), .ZN(n9211) );
  INV_X1 U5947 ( .A(n8623), .ZN(n4599) );
  AND2_X1 U5948 ( .A1(n7322), .A2(n7232), .ZN(n7233) );
  AND2_X1 U5949 ( .A1(n6546), .A2(n6539), .ZN(n9966) );
  INV_X1 U5950 ( .A(n9960), .ZN(n9214) );
  NAND2_X1 U5951 ( .A1(n6550), .A2(n10056), .ZN(n9217) );
  INV_X1 U5952 ( .A(n9966), .ZN(n9220) );
  XNOR2_X1 U5953 ( .A(n5443), .B(P1_IR_REG_20__SCAN_IN), .ZN(n9467) );
  INV_X1 U5954 ( .A(n9196), .ZN(n9491) );
  INV_X1 U5955 ( .A(n6919), .ZN(n9516) );
  NOR2_X1 U5956 ( .A1(n5074), .A2(n5073), .ZN(n5506) );
  NAND2_X1 U5957 ( .A1(n5518), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U5958 ( .A1(n4616), .A2(n4614), .ZN(n9994) );
  INV_X1 U5959 ( .A(n4615), .ZN(n4614) );
  INV_X1 U5960 ( .A(n4929), .ZN(n9518) );
  NOR2_X1 U5961 ( .A1(n10019), .A2(n4528), .ZN(n6796) );
  INV_X1 U5962 ( .A(n4932), .ZN(n6794) );
  NOR2_X1 U5963 ( .A1(n6799), .A2(n6798), .ZN(n6797) );
  AND2_X1 U5964 ( .A1(n10012), .A2(n4619), .ZN(n6799) );
  NAND2_X1 U5965 ( .A1(n10024), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n4619) );
  NOR2_X1 U5966 ( .A1(n6821), .A2(n6820), .ZN(n6819) );
  AND2_X1 U5967 ( .A1(n4932), .A2(n4931), .ZN(n6821) );
  NAND2_X1 U5968 ( .A1(n6800), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4931) );
  NOR2_X1 U5969 ( .A1(n6555), .A2(n4934), .ZN(n6808) );
  NOR2_X1 U5970 ( .A1(n6554), .A2(n4935), .ZN(n4934) );
  NOR2_X1 U5971 ( .A1(n6808), .A2(n6807), .ZN(n6806) );
  INV_X1 U5972 ( .A(n4613), .ZN(n6809) );
  NOR2_X1 U5973 ( .A1(n6806), .A2(n4933), .ZN(n6557) );
  AND2_X1 U5974 ( .A1(n6812), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4933) );
  NAND2_X1 U5975 ( .A1(n6557), .A2(n6558), .ZN(n6781) );
  NAND2_X1 U5976 ( .A1(n6784), .A2(n4611), .ZN(n6788) );
  OR2_X1 U5977 ( .A1(n6785), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n4611) );
  NOR2_X1 U5978 ( .A1(n7068), .A2(n7069), .ZN(n7119) );
  NOR2_X1 U5979 ( .A1(n7067), .A2(n4941), .ZN(n7069) );
  AND2_X1 U5980 ( .A1(n7071), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4941) );
  NOR2_X1 U5981 ( .A1(n7070), .A2(n4617), .ZN(n7074) );
  AND2_X1 U5982 ( .A1(n7071), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n4617) );
  NOR2_X1 U5983 ( .A1(n7074), .A2(n7073), .ZN(n7125) );
  NOR2_X1 U5984 ( .A1(n7119), .A2(n4940), .ZN(n7122) );
  AND2_X1 U5985 ( .A1(n7123), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4940) );
  NAND2_X1 U5986 ( .A1(n7122), .A2(n7121), .ZN(n7369) );
  NOR2_X1 U5987 ( .A1(n7477), .A2(n4936), .ZN(n7480) );
  AND2_X1 U5988 ( .A1(n7482), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4936) );
  NOR2_X1 U5989 ( .A1(n7480), .A2(n7479), .ZN(n7763) );
  NOR2_X1 U5990 ( .A1(n7481), .A2(n4618), .ZN(n7485) );
  AND2_X1 U5991 ( .A1(n7482), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n4618) );
  XNOR2_X1 U5992 ( .A(n9543), .B(n9542), .ZN(n7765) );
  INV_X1 U5993 ( .A(n9593), .ZN(n10018) );
  NOR2_X1 U5994 ( .A1(n9533), .A2(n9534), .ZN(n9538) );
  NAND2_X1 U5995 ( .A1(n9538), .A2(n9537), .ZN(n9560) );
  OR2_X1 U5996 ( .A1(n7793), .A2(n5016), .ZN(n9606) );
  NAND2_X1 U5997 ( .A1(n4789), .A2(n5686), .ZN(n9646) );
  NAND2_X1 U5998 ( .A1(n9695), .A2(n9296), .ZN(n9683) );
  NAND2_X1 U5999 ( .A1(n4801), .A2(n4507), .ZN(n9688) );
  AND2_X1 U6000 ( .A1(n4801), .A2(n4529), .ZN(n9689) );
  NAND2_X1 U6001 ( .A1(n4802), .A2(n5094), .ZN(n4801) );
  NAND2_X1 U6002 ( .A1(n4818), .A2(n4820), .ZN(n9741) );
  NAND2_X1 U6003 ( .A1(n9776), .A2(n4822), .ZN(n4818) );
  NAND2_X1 U6004 ( .A1(n4808), .A2(n4807), .ZN(n4806) );
  NAND2_X1 U6005 ( .A1(n7586), .A2(n9347), .ZN(n4809) );
  AND2_X1 U6006 ( .A1(n4706), .A2(n9409), .ZN(n7706) );
  NAND2_X1 U6007 ( .A1(n7386), .A2(n9402), .ZN(n7437) );
  NAND2_X1 U6008 ( .A1(n9475), .A2(n6549), .ZN(n10056) );
  INV_X1 U6009 ( .A(n6548), .ZN(n6549) );
  NAND2_X1 U6010 ( .A1(n10032), .A2(n10033), .ZN(n4786) );
  INV_X1 U6011 ( .A(n9611), .ZN(n10066) );
  OR2_X1 U6012 ( .A1(n7170), .A2(n9598), .ZN(n9611) );
  INV_X1 U6013 ( .A(n9800), .ZN(n10060) );
  INV_X1 U6014 ( .A(n9458), .ZN(n9880) );
  OR2_X1 U6015 ( .A1(n10168), .A2(n5012), .ZN(n5084) );
  INV_X1 U6016 ( .A(n9628), .ZN(n9885) );
  INV_X1 U6017 ( .A(n9656), .ZN(n9893) );
  INV_X1 U6018 ( .A(n9671), .ZN(n9897) );
  INV_X1 U6019 ( .A(n9715), .ZN(n9909) );
  INV_X1 U6020 ( .A(n9796), .ZN(n9925) );
  INV_X1 U6021 ( .A(n7653), .ZN(n9964) );
  NOR2_X1 U6022 ( .A1(n6926), .A2(P1_U3086), .ZN(n9475) );
  INV_X1 U6023 ( .A(n9475), .ZN(n6850) );
  AND2_X1 U6024 ( .A1(n5020), .A2(n4566), .ZN(n4826) );
  INV_X1 U6025 ( .A(n5442), .ZN(n4825) );
  XNOR2_X1 U6026 ( .A(n5450), .B(n5449), .ZN(n7800) );
  NOR2_X1 U6027 ( .A1(n5121), .A2(n5120), .ZN(n5122) );
  INV_X1 U6028 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8913) );
  NOR2_X1 U6029 ( .A1(n4835), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7574) );
  INV_X1 U6030 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9041) );
  INV_X1 U6031 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7368) );
  INV_X1 U6032 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7224) );
  INV_X1 U6033 ( .A(n9467), .ZN(n7225) );
  INV_X1 U6034 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6600) );
  INV_X1 U6035 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6459) );
  NAND2_X1 U6036 ( .A1(n5179), .A2(n4988), .ZN(n4727) );
  NAND2_X1 U6037 ( .A1(n4993), .A2(n5182), .ZN(n5192) );
  NAND2_X1 U6038 ( .A1(n5179), .A2(n5178), .ZN(n4993) );
  INV_X1 U6039 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6436) );
  AOI21_X1 U6040 ( .B1(n4652), .B2(n4510), .A(n4649), .ZN(n4648) );
  NAND2_X1 U6041 ( .A1(n4651), .A2(n4652), .ZN(n4650) );
  INV_X1 U6042 ( .A(n4876), .ZN(n6854) );
  NAND2_X1 U6043 ( .A1(n4604), .A2(n4532), .ZN(P2_U3200) );
  NAND2_X1 U6044 ( .A1(n4605), .A2(n10348), .ZN(n4604) );
  OAI211_X1 U6045 ( .C1(n6993), .C2(n4737), .A(n4736), .B(n4735), .ZN(P2_U3201) );
  NOR2_X1 U6046 ( .A1(n5956), .A2(n5955), .ZN(n4735) );
  NAND2_X1 U6047 ( .A1(n5947), .A2(n10347), .ZN(n4736) );
  XNOR2_X1 U6048 ( .A(n4738), .B(n5887), .ZN(n4737) );
  INV_X1 U6049 ( .A(n6357), .ZN(n6358) );
  OAI21_X1 U6050 ( .B1(n6390), .B2(n8451), .A(n6356), .ZN(n6357) );
  OAI21_X1 U6051 ( .B1(n9599), .B2(n9598), .A(n4942), .ZN(P1_U3262) );
  AOI21_X1 U6052 ( .B1(n4944), .B2(n9598), .A(n4943), .ZN(n4942) );
  NOR2_X1 U6053 ( .A1(n5018), .A2(n9875), .ZN(n5488) );
  NOR2_X1 U6054 ( .A1(n5769), .A2(n5768), .ZN(n5770) );
  OR2_X1 U6055 ( .A1(n5018), .A2(n9929), .ZN(n5082) );
  OAI21_X1 U6056 ( .B1(n5958), .B2(n10173), .A(n4730), .ZN(n5961) );
  OR2_X1 U6057 ( .A1(n10175), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n4730) );
  NOR2_X1 U6058 ( .A1(n8469), .A2(n6208), .ZN(n4505) );
  AND2_X1 U6059 ( .A1(n4810), .A2(n4805), .ZN(n4506) );
  AND2_X1 U6060 ( .A1(n5677), .A2(n4529), .ZN(n4507) );
  AND2_X2 U6061 ( .A1(n4995), .A2(n4994), .ZN(n5124) );
  INV_X1 U6062 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9931) );
  AND2_X1 U6063 ( .A1(n8041), .A2(n8106), .ZN(n4508) );
  NAND2_X1 U6064 ( .A1(n9748), .A2(n9499), .ZN(n4509) );
  NAND2_X1 U6065 ( .A1(n8119), .A2(n7261), .ZN(n4510) );
  NAND2_X1 U6066 ( .A1(n6200), .A2(n6199), .ZN(n8469) );
  NAND2_X1 U6067 ( .A1(n6230), .A2(n6229), .ZN(n8518) );
  AND4_X1 U6068 ( .A1(n5792), .A2(n5791), .A3(n5790), .A4(n5789), .ZN(n4511)
         );
  OR2_X1 U6069 ( .A1(n8508), .A2(n8316), .ZN(n4512) );
  AND2_X1 U6070 ( .A1(n9333), .A2(n9501), .ZN(n4513) );
  NOR2_X1 U6071 ( .A1(n8172), .A2(n8187), .ZN(n4514) );
  INV_X1 U6072 ( .A(n8039), .ZN(n4637) );
  AND2_X1 U6073 ( .A1(n10132), .A2(n10138), .ZN(n4515) );
  OR2_X1 U6074 ( .A1(n8476), .A2(n8202), .ZN(n7941) );
  INV_X1 U6075 ( .A(n4812), .ZN(n4807) );
  OR2_X1 U6076 ( .A1(n4813), .A2(n5608), .ZN(n4812) );
  INV_X1 U6077 ( .A(n5030), .ZN(n5029) );
  NAND2_X1 U6078 ( .A1(n5032), .A2(n5031), .ZN(n5030) );
  AND2_X1 U6079 ( .A1(n9678), .A2(n5022), .ZN(n9612) );
  OR2_X1 U6080 ( .A1(n4637), .A2(n4635), .ZN(n4516) );
  INV_X1 U6081 ( .A(n8105), .ZN(n4982) );
  AND2_X1 U6082 ( .A1(n5113), .A2(n5117), .ZN(n4517) );
  AND2_X1 U6083 ( .A1(n5070), .A2(n4569), .ZN(n4518) );
  AOI21_X1 U6084 ( .B1(n10251), .B2(n4888), .A(n4886), .ZN(n4884) );
  XNOR2_X1 U6085 ( .A(n5788), .B(n5787), .ZN(n6332) );
  OR2_X1 U6086 ( .A1(n6690), .A2(n6691), .ZN(n6704) );
  AND2_X1 U6087 ( .A1(n5828), .A2(n5827), .ZN(n10290) );
  OR2_X1 U6088 ( .A1(n9732), .A2(n9734), .ZN(n4519) );
  NAND2_X1 U6089 ( .A1(n5127), .A2(n4500), .ZN(n5166) );
  OR2_X1 U6091 ( .A1(n5297), .A2(n4860), .ZN(n4520) );
  INV_X1 U6092 ( .A(n5783), .ZN(n5819) );
  AND2_X1 U6093 ( .A1(n4512), .A2(n5043), .ZN(n4521) );
  NAND4_X1 U6094 ( .A1(n5499), .A2(n5498), .A3(n5497), .A4(n5496), .ZN(n6633)
         );
  NAND2_X1 U6095 ( .A1(n5804), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5803) );
  XNOR2_X1 U6096 ( .A(n8463), .B(n8273), .ZN(n8375) );
  INV_X1 U6097 ( .A(n8375), .ZN(n4762) );
  AND2_X1 U6098 ( .A1(n4718), .A2(n4719), .ZN(n4522) );
  OR2_X1 U6099 ( .A1(n4854), .A2(n4851), .ZN(n4523) );
  NAND2_X1 U6100 ( .A1(n6651), .A2(n4664), .ZN(n6681) );
  INV_X1 U6101 ( .A(n6681), .ZN(n6653) );
  OR2_X1 U6102 ( .A1(n9765), .A2(n9500), .ZN(n4524) );
  NAND2_X1 U6103 ( .A1(n5805), .A2(n5785), .ZN(n5804) );
  NAND2_X1 U6104 ( .A1(n5177), .A2(n5107), .ZN(n5197) );
  NAND4_X2 U6105 ( .A1(n6042), .A2(n6041), .A3(n6040), .A4(n6039), .ZN(n8286)
         );
  AND2_X1 U6106 ( .A1(n10001), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4525) );
  OR2_X1 U6107 ( .A1(n5442), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n4526) );
  NAND2_X1 U6108 ( .A1(n4939), .A2(n5177), .ZN(n4527) );
  AND2_X1 U6109 ( .A1(n10024), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4528) );
  NAND2_X1 U6110 ( .A1(n4663), .A2(n7849), .ZN(n8191) );
  NAND2_X1 U6111 ( .A1(n4959), .A2(n7851), .ZN(n8165) );
  NAND2_X1 U6112 ( .A1(n9703), .A2(n9496), .ZN(n4529) );
  NOR2_X1 U6113 ( .A1(n10217), .A2(n4871), .ZN(n4530) );
  NAND2_X1 U6114 ( .A1(n6308), .A2(n8082), .ZN(n8322) );
  NAND2_X1 U6115 ( .A1(n4790), .A2(n4796), .ZN(n9623) );
  NAND2_X1 U6116 ( .A1(n4957), .A2(n7840), .ZN(n8158) );
  AND2_X1 U6117 ( .A1(n7895), .A2(n7894), .ZN(n8443) );
  OR2_X1 U6118 ( .A1(n6322), .A2(n6984), .ZN(n4531) );
  AND2_X1 U6119 ( .A1(n7884), .A2(n7800), .ZN(n5503) );
  AND4_X1 U6120 ( .A1(n6059), .A2(n6058), .A3(n6057), .A4(n6056), .ZN(n7058)
         );
  INV_X1 U6121 ( .A(n7058), .ZN(n8284) );
  AND3_X1 U6122 ( .A1(n6034), .A2(n6033), .A3(n6032), .ZN(n6736) );
  AND4_X1 U6123 ( .A1(n4603), .A2(n9955), .A3(n9953), .A4(n9954), .ZN(n4532)
         );
  INV_X1 U6124 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5842) );
  NOR2_X1 U6125 ( .A1(n6325), .A2(n4770), .ZN(n7807) );
  AND4_X1 U6126 ( .A1(n5986), .A2(n5985), .A3(n5984), .A4(n5983), .ZN(n5995)
         );
  INV_X1 U6127 ( .A(n8071), .ZN(n4765) );
  NOR2_X1 U6128 ( .A1(n6291), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n5805) );
  AND4_X1 U6129 ( .A1(n6087), .A2(n6086), .A3(n6085), .A4(n6084), .ZN(n7426)
         );
  INV_X1 U6130 ( .A(n9690), .ZN(n9901) );
  NAND2_X1 U6131 ( .A1(n5365), .A2(n5364), .ZN(n9690) );
  NAND2_X1 U6132 ( .A1(n5129), .A2(n5105), .ZN(n5141) );
  NOR2_X1 U6133 ( .A1(n8250), .A2(n8275), .ZN(n4533) );
  NAND2_X2 U6134 ( .A1(n5973), .A2(n5974), .ZN(n7900) );
  INV_X1 U6135 ( .A(n9639), .ZN(n9889) );
  NAND2_X1 U6136 ( .A1(n5392), .A2(n5391), .ZN(n9639) );
  NOR2_X1 U6137 ( .A1(n6109), .A2(n7183), .ZN(n4534) );
  NAND2_X1 U6138 ( .A1(n5437), .A2(n5436), .ZN(n9327) );
  INV_X1 U6139 ( .A(n4704), .ZN(n4703) );
  NOR2_X1 U6140 ( .A1(n4705), .A2(n5745), .ZN(n4704) );
  INV_X1 U6141 ( .A(n4869), .ZN(n4868) );
  NOR2_X1 U6142 ( .A1(n5248), .A2(n4870), .ZN(n4869) );
  AND2_X1 U6143 ( .A1(n4965), .A2(n7154), .ZN(n4535) );
  NOR2_X1 U6144 ( .A1(n7063), .A2(n7008), .ZN(n4536) );
  NOR2_X1 U6145 ( .A1(n4843), .A2(n5346), .ZN(n4842) );
  AND2_X1 U6146 ( .A1(n8518), .A2(n8361), .ZN(n7908) );
  INV_X1 U6147 ( .A(n7908), .ZN(n4759) );
  AND2_X1 U6148 ( .A1(n4952), .A2(n4675), .ZN(n4537) );
  INV_X1 U6149 ( .A(n4797), .ZN(n4796) );
  AOI21_X1 U6150 ( .B1(n7177), .B2(n8008), .A(n8005), .ZN(n4987) );
  AND2_X1 U6151 ( .A1(n4622), .A2(n4621), .ZN(n4538) );
  AND2_X1 U6152 ( .A1(n9765), .A2(n9500), .ZN(n4539) );
  AND2_X1 U6153 ( .A1(n9313), .A2(n9310), .ZN(n9624) );
  INV_X1 U6154 ( .A(n9624), .ZN(n4717) );
  INV_X1 U6155 ( .A(n5075), .ZN(n4918) );
  AND2_X1 U6156 ( .A1(n9901), .A2(n9171), .ZN(n4540) );
  INV_X1 U6157 ( .A(n4764), .ZN(n4763) );
  NOR2_X1 U6158 ( .A1(n4765), .A2(n7909), .ZN(n4764) );
  AND2_X1 U6159 ( .A1(n5650), .A2(n4814), .ZN(n4541) );
  AND2_X1 U6160 ( .A1(n6333), .A2(n4973), .ZN(n4542) );
  AND4_X1 U6161 ( .A1(n6008), .A2(n6007), .A3(n6006), .A4(n6005), .ZN(n6692)
         );
  AND2_X1 U6162 ( .A1(n7516), .A2(n5006), .ZN(n4544) );
  AND2_X1 U6163 ( .A1(n5092), .A2(n7896), .ZN(n4545) );
  NAND2_X1 U6164 ( .A1(n4794), .A2(n4791), .ZN(n5724) );
  INV_X1 U6165 ( .A(n4601), .ZN(n5839) );
  NOR2_X1 U6166 ( .A1(n5836), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n4601) );
  AND2_X1 U6167 ( .A1(n5247), .A2(SI_12_), .ZN(n4546) );
  AND2_X1 U6168 ( .A1(n5201), .A2(SI_7_), .ZN(n4547) );
  AND2_X1 U6169 ( .A1(n5193), .A2(SI_6_), .ZN(n4548) );
  NOR2_X1 U6170 ( .A1(n8463), .A2(n8273), .ZN(n4549) );
  OR2_X1 U6171 ( .A1(n5087), .A2(n5096), .ZN(n4550) );
  INV_X1 U6172 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5114) );
  NOR2_X1 U6173 ( .A1(n8747), .A2(n9220), .ZN(n4551) );
  AND2_X1 U6174 ( .A1(n4699), .A2(n9243), .ZN(n4552) );
  AND2_X1 U6175 ( .A1(n9295), .A2(n9296), .ZN(n9697) );
  INV_X1 U6176 ( .A(n9697), .ZN(n4723) );
  INV_X1 U6177 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6439) );
  NAND2_X1 U6178 ( .A1(n4821), .A2(n4524), .ZN(n4820) );
  NAND2_X1 U6179 ( .A1(n4819), .A2(n5643), .ZN(n4553) );
  INV_X1 U6180 ( .A(n4823), .ZN(n4822) );
  NAND2_X1 U6181 ( .A1(n4524), .A2(n5630), .ZN(n4823) );
  AND2_X1 U6182 ( .A1(n5446), .A2(n5449), .ZN(n4554) );
  NAND2_X1 U6183 ( .A1(n8037), .A2(n8036), .ZN(n4555) );
  AND2_X1 U6184 ( .A1(n5226), .A2(n5222), .ZN(n4556) );
  AND2_X1 U6185 ( .A1(n4760), .A2(n4759), .ZN(n4557) );
  INV_X1 U6186 ( .A(n4927), .ZN(n4926) );
  NOR2_X1 U6187 ( .A1(n7176), .A2(n8005), .ZN(n4558) );
  AND2_X1 U6188 ( .A1(n5810), .A2(n5068), .ZN(n4559) );
  AND2_X1 U6189 ( .A1(n5021), .A2(n4517), .ZN(n4560) );
  OR2_X1 U6190 ( .A1(n5151), .A2(n6567), .ZN(n4561) );
  NOR2_X1 U6191 ( .A1(n7938), .A2(n4983), .ZN(n4562) );
  AND2_X1 U6192 ( .A1(n4749), .A2(n4748), .ZN(n4563) );
  OAI22_X1 U6193 ( .A1(n6444), .A2(n4500), .B1(n4836), .B2(n4835), .ZN(n4773)
         );
  NOR2_X1 U6194 ( .A1(n7845), .A2(n8221), .ZN(n4564) );
  NAND2_X1 U6195 ( .A1(n10416), .A2(n8281), .ZN(n4565) );
  AND2_X1 U6196 ( .A1(n4554), .A2(n4828), .ZN(n4566) );
  AND2_X1 U6197 ( .A1(n8013), .A2(n8012), .ZN(n7923) );
  NAND2_X1 U6198 ( .A1(n7837), .A2(n8413), .ZN(n4567) );
  INV_X1 U6199 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5068) );
  NAND2_X1 U6200 ( .A1(n7098), .A2(n7944), .ZN(n6950) );
  INV_X1 U6201 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4836) );
  NAND2_X1 U6202 ( .A1(n9678), .A2(n9901), .ZN(n9668) );
  INV_X1 U6203 ( .A(n8023), .ZN(n5062) );
  NAND2_X1 U6204 ( .A1(n4706), .A2(n4704), .ZN(n7705) );
  NAND2_X1 U6205 ( .A1(n8376), .A2(n8375), .ZN(n8377) );
  OAI21_X1 U6206 ( .B1(n7637), .B2(n4926), .A(n4923), .ZN(n7662) );
  NAND2_X1 U6207 ( .A1(n5415), .A2(n5414), .ZN(n9810) );
  INV_X1 U6208 ( .A(n9810), .ZN(n5012) );
  NOR2_X1 U6209 ( .A1(n9795), .A2(n9796), .ZN(n5295) );
  OR2_X1 U6210 ( .A1(n6886), .A2(n6065), .ZN(n4568) );
  INV_X1 U6211 ( .A(n10209), .ZN(n6456) );
  INV_X1 U6212 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4589) );
  AND4_X1 U6213 ( .A1(n6493), .A2(n6492), .A3(n6491), .A4(n6490), .ZN(n6642)
         );
  INV_X1 U6214 ( .A(n8106), .ZN(n8112) );
  NAND2_X1 U6215 ( .A1(n8476), .A2(n8426), .ZN(n4569) );
  NAND2_X1 U6216 ( .A1(n4710), .A2(n4708), .ZN(n9742) );
  NAND2_X1 U6217 ( .A1(n4806), .A2(n4810), .ZN(n7725) );
  OAI21_X1 U6218 ( .B1(n9776), .B2(n4513), .A(n5630), .ZN(n9755) );
  NAND2_X1 U6219 ( .A1(n4809), .A2(n5600), .ZN(n7704) );
  AND2_X1 U6220 ( .A1(n4515), .A2(n10145), .ZN(n4570) );
  AND2_X1 U6221 ( .A1(n8211), .A2(n8020), .ZN(n4571) );
  NAND2_X1 U6222 ( .A1(n5269), .A2(n5268), .ZN(n9263) );
  NAND2_X1 U6223 ( .A1(n4881), .A2(n5783), .ZN(n5813) );
  AND2_X1 U6224 ( .A1(n7841), .A2(n8222), .ZN(n4572) );
  AND2_X1 U6225 ( .A1(n7852), .A2(n8326), .ZN(n4573) );
  NAND2_X1 U6226 ( .A1(n5783), .A2(n5782), .ZN(n5817) );
  NAND2_X1 U6227 ( .A1(n7733), .A2(n8051), .ZN(n8436) );
  AND2_X1 U6228 ( .A1(n9656), .A2(n9493), .ZN(n4574) );
  INV_X1 U6229 ( .A(n9748), .ZN(n9917) );
  NAND2_X1 U6230 ( .A1(n5332), .A2(n5331), .ZN(n9748) );
  AND2_X1 U6231 ( .A1(n6237), .A2(n6236), .ZN(n8361) );
  NAND2_X1 U6232 ( .A1(n9678), .A2(n5024), .ZN(n5027) );
  NAND2_X1 U6233 ( .A1(n5295), .A2(n5009), .ZN(n5010) );
  AND2_X1 U6234 ( .A1(n4970), .A2(n4687), .ZN(n4575) );
  AND2_X1 U6235 ( .A1(n4892), .A2(n4897), .ZN(n4576) );
  AND2_X1 U6236 ( .A1(n9702), .A2(n9905), .ZN(n9678) );
  AND2_X1 U6237 ( .A1(n4671), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n4577) );
  AND2_X1 U6238 ( .A1(n5345), .A2(SI_21_), .ZN(n4578) );
  AND2_X1 U6239 ( .A1(n9218), .A2(n9503), .ZN(n4579) );
  INV_X1 U6240 ( .A(n10058), .ZN(n10070) );
  NAND2_X1 U6241 ( .A1(n5305), .A2(n5304), .ZN(n9333) );
  AOI21_X1 U6242 ( .B1(n8392), .B2(n6266), .A(n6207), .ZN(n8222) );
  INV_X1 U6243 ( .A(n8222), .ZN(n6208) );
  AND2_X1 U6244 ( .A1(n5871), .A2(n5870), .ZN(n10241) );
  NAND2_X1 U6245 ( .A1(n7442), .A2(n7645), .ZN(n7441) );
  AND2_X1 U6246 ( .A1(n7212), .A2(n5075), .ZN(n4580) );
  INV_X1 U6247 ( .A(n10307), .ZN(n6601) );
  AND2_X1 U6248 ( .A1(n7767), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n4581) );
  AND2_X1 U6249 ( .A1(n7767), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4582) );
  INV_X1 U6250 ( .A(n10033), .ZN(n4783) );
  NAND2_X1 U6251 ( .A1(n6577), .A2(n7993), .ZN(n6735) );
  NAND2_X1 U6252 ( .A1(n4948), .A2(n4947), .ZN(n5800) );
  NAND2_X1 U6253 ( .A1(n4782), .A2(n4784), .ZN(n7403) );
  NAND2_X1 U6254 ( .A1(n4786), .A2(n5551), .ZN(n7343) );
  NAND2_X1 U6255 ( .A1(n4997), .A2(n6302), .ZN(n7544) );
  AND2_X1 U6256 ( .A1(n5908), .A2(n10257), .ZN(n4583) );
  NAND2_X1 U6257 ( .A1(n6576), .A2(n7981), .ZN(n6577) );
  NAND2_X1 U6258 ( .A1(n7442), .A2(n5029), .ZN(n5033) );
  INV_X1 U6259 ( .A(n4900), .ZN(n4898) );
  AND2_X1 U6260 ( .A1(n5912), .A2(n10290), .ZN(n4900) );
  INV_X2 U6261 ( .A(n10432), .ZN(n10430) );
  INV_X1 U6262 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n4935) );
  INV_X1 U6263 ( .A(n9950), .ZN(n4914) );
  NAND2_X1 U6264 ( .A1(n5254), .A2(n5253), .ZN(n7625) );
  INV_X1 U6265 ( .A(n7625), .ZN(n5031) );
  NOR2_X1 U6266 ( .A1(n4890), .A2(n6482), .ZN(n4889) );
  INV_X1 U6267 ( .A(n4889), .ZN(n4888) );
  OAI22_X1 U6268 ( .A1(n6938), .A2(n6939), .B1(n6655), .B2(n6652), .ZN(n6685)
         );
  OR2_X1 U6269 ( .A1(n9561), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n4584) );
  INV_X1 U6270 ( .A(n5728), .ZN(n9337) );
  XNOR2_X1 U6271 ( .A(n5500), .B(n6633), .ZN(n5728) );
  NAND2_X1 U6272 ( .A1(n5123), .A2(n5122), .ZN(n5456) );
  INV_X1 U6273 ( .A(n4908), .ZN(n4907) );
  NOR2_X1 U6274 ( .A1(n4912), .A2(n4909), .ZN(n4908) );
  AND2_X1 U6275 ( .A1(n4747), .A2(n4746), .ZN(n4585) );
  INV_X1 U6276 ( .A(n6886), .ZN(n4873) );
  AND2_X1 U6277 ( .A1(n6294), .A2(n6293), .ZN(n8118) );
  OR2_X1 U6278 ( .A1(n9950), .A2(n9114), .ZN(n4586) );
  NOR2_X1 U6279 ( .A1(n5970), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n8547) );
  NOR2_X1 U6280 ( .A1(n9995), .A2(n9994), .ZN(n4587) );
  INV_X1 U6281 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n6915) );
  INV_X1 U6282 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n4973) );
  NAND2_X1 U6283 ( .A1(n6984), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4748) );
  INV_X1 U6284 ( .A(n6984), .ZN(n4609) );
  NAND2_X1 U6285 ( .A1(n8752), .A2(n8621), .ZN(n8624) );
  NAND2_X1 U6286 ( .A1(n4600), .A2(n4599), .ZN(n8625) );
  AND2_X2 U6287 ( .A1(n9192), .A2(n8670), .ZN(n8739) );
  XNOR2_X2 U6288 ( .A(n4592), .B(n8731), .ZN(n7685) );
  OAI22_X2 U6289 ( .A1(n10169), .A2(n6531), .B1(n7638), .B2(n8728), .ZN(n4592)
         );
  NAND2_X1 U6290 ( .A1(n6460), .A2(n5434), .ZN(n4593) );
  OAI21_X1 U6291 ( .B1(n9259), .B2(n9406), .A(n9409), .ZN(n9260) );
  NAND2_X1 U6292 ( .A1(n4596), .A2(n4595), .ZN(n9261) );
  MUX2_X1 U6293 ( .A(n9324), .B(n9321), .S(n9458), .Z(n9323) );
  AOI21_X1 U6294 ( .B1(n9242), .B2(n9241), .A(n9240), .ZN(n9248) );
  NOR2_X1 U6295 ( .A1(n9273), .A2(n9272), .ZN(n9277) );
  AOI211_X1 U6296 ( .C1(n9616), .C2(n9313), .A(n9439), .B(n9304), .ZN(n9306)
         );
  NAND3_X1 U6297 ( .A1(n6915), .A2(n4831), .A3(n5099), .ZN(n4995) );
  INV_X1 U6298 ( .A(n5111), .ZN(n4779) );
  INV_X1 U6299 ( .A(n8624), .ZN(n4600) );
  INV_X1 U6300 ( .A(n5178), .ZN(n4989) );
  NAND2_X2 U6301 ( .A1(n5229), .A2(n5228), .ZN(n5239) );
  NAND2_X1 U6302 ( .A1(n4984), .A2(n4981), .ZN(n8123) );
  INV_X1 U6303 ( .A(n4656), .ZN(n4655) );
  AND2_X1 U6304 ( .A1(n6296), .A2(n7966), .ZN(n4771) );
  NAND2_X1 U6305 ( .A1(n5731), .A2(n5730), .ZN(n7304) );
  NAND3_X1 U6306 ( .A1(n6924), .A2(n6925), .A3(n5075), .ZN(n4917) );
  NAND2_X1 U6307 ( .A1(n6634), .A2(n6635), .ZN(n4598) );
  OAI21_X4 U6308 ( .B1(n7515), .B2(n7514), .A(n7513), .ZN(n7637) );
  NAND2_X1 U6309 ( .A1(n5327), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5329) );
  OAI21_X1 U6310 ( .B1(n9995), .B2(n4615), .A(n4616), .ZN(n9527) );
  NAND3_X1 U6311 ( .A1(n7991), .A2(n7990), .A3(n8112), .ZN(n4622) );
  NAND2_X1 U6312 ( .A1(n7982), .A2(n7981), .ZN(n7996) );
  XNOR2_X1 U6313 ( .A(n8287), .B(n6694), .ZN(n7981) );
  NAND2_X1 U6314 ( .A1(n4628), .A2(n4629), .ZN(n8059) );
  NAND2_X1 U6315 ( .A1(n8035), .A2(n4631), .ZN(n4628) );
  INV_X1 U6316 ( .A(n8034), .ZN(n4635) );
  NAND3_X1 U6317 ( .A1(n4642), .A2(n4639), .A3(n7923), .ZN(n4638) );
  OR2_X2 U6318 ( .A1(n8123), .A2(n7261), .ZN(n4660) );
  INV_X1 U6319 ( .A(n8121), .ZN(n4644) );
  NAND2_X1 U6320 ( .A1(n4644), .A2(n4652), .ZN(n4645) );
  NOR2_X2 U6321 ( .A1(n4656), .A2(n4654), .ZN(n4652) );
  INV_X1 U6322 ( .A(n8120), .ZN(n4651) );
  NAND4_X1 U6323 ( .A1(n4646), .A2(n4648), .A3(n4650), .A4(n4645), .ZN(
        P2_U3296) );
  NAND3_X1 U6324 ( .A1(n8120), .A2(n8121), .A3(n4647), .ZN(n4646) );
  OAI21_X2 U6325 ( .B1(n4659), .B2(n4658), .A(n4657), .ZN(n4656) );
  AND2_X2 U6326 ( .A1(n5774), .A2(n5773), .ZN(n5783) );
  NAND2_X1 U6327 ( .A1(n4662), .A2(n4958), .ZN(n8240) );
  NAND2_X1 U6328 ( .A1(n8191), .A2(n4960), .ZN(n4662) );
  NAND2_X1 U6329 ( .A1(n8140), .A2(n8221), .ZN(n4663) );
  OR2_X1 U6330 ( .A1(n5800), .A2(n4674), .ZN(n4668) );
  NAND3_X1 U6331 ( .A1(n4667), .A2(n4666), .A3(n4669), .ZN(n6331) );
  NAND2_X1 U6332 ( .A1(n5800), .A2(n4672), .ZN(n4666) );
  OAI21_X1 U6333 ( .B1(n8174), .B2(n4679), .A(n4677), .ZN(n8198) );
  NAND2_X1 U6334 ( .A1(n8174), .A2(n4677), .ZN(n4676) );
  OAI21_X1 U6335 ( .B1(n8174), .B2(n4514), .A(n7826), .ZN(n8146) );
  NAND4_X1 U6336 ( .A1(n5774), .A2(n4686), .A3(n4968), .A4(n4685), .ZN(n6291)
         );
  NAND4_X1 U6337 ( .A1(n5782), .A2(n5774), .A3(n4968), .A4(n5773), .ZN(n5883)
         );
  NAND2_X1 U6338 ( .A1(n7747), .A2(n4690), .ZN(n4688) );
  INV_X2 U6339 ( .A(n6681), .ZN(n7856) );
  AND2_X1 U6340 ( .A1(n9246), .A2(n5739), .ZN(n9237) );
  OAI21_X1 U6341 ( .B1(n4703), .B2(n5746), .A(n9414), .ZN(n4701) );
  NAND2_X1 U6342 ( .A1(n9791), .A2(n4711), .ZN(n4710) );
  NAND2_X1 U6343 ( .A1(n9618), .A2(n9222), .ZN(n4714) );
  NAND2_X1 U6344 ( .A1(n9696), .A2(n4721), .ZN(n4718) );
  NAND3_X1 U6345 ( .A1(n5179), .A2(n4988), .A3(n5199), .ZN(n4726) );
  NAND2_X1 U6346 ( .A1(n4727), .A2(n4990), .ZN(n5200) );
  INV_X1 U6347 ( .A(n4990), .ZN(n4728) );
  XNOR2_X2 U6348 ( .A(n5221), .B(n5219), .ZN(n6458) );
  XNOR2_X2 U6349 ( .A(n4741), .B(P2_IR_REG_2__SCAN_IN), .ZN(n7036) );
  NOR2_X1 U6350 ( .A1(n4492), .A2(n4674), .ZN(n4741) );
  NAND2_X1 U6351 ( .A1(n6985), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4745) );
  NAND2_X1 U6352 ( .A1(n4563), .A2(n4745), .ZN(n4744) );
  NAND2_X1 U6353 ( .A1(n5927), .A2(n6999), .ZN(n4749) );
  NAND2_X1 U6354 ( .A1(n4752), .A2(n6576), .ZN(n4751) );
  NAND3_X1 U6355 ( .A1(n4751), .A2(n4750), .A3(n7987), .ZN(n6299) );
  NAND2_X1 U6356 ( .A1(n8376), .A2(n4557), .ZN(n4755) );
  NAND2_X1 U6357 ( .A1(n4755), .A2(n4756), .ZN(n8334) );
  NAND3_X1 U6358 ( .A1(n4767), .A2(n7923), .A3(n4766), .ZN(n7252) );
  AND2_X1 U6359 ( .A1(n4558), .A2(n7944), .ZN(n4768) );
  OR2_X2 U6360 ( .A1(n7732), .A2(n8043), .ZN(n7733) );
  NAND2_X1 U6361 ( .A1(n6710), .A2(n7966), .ZN(n6589) );
  NAND2_X1 U6362 ( .A1(n4771), .A2(n7959), .ZN(n6710) );
  NAND2_X1 U6363 ( .A1(n6322), .A2(n4773), .ZN(n4772) );
  INV_X1 U6364 ( .A(n5781), .ZN(n4777) );
  NAND3_X1 U6365 ( .A1(n4881), .A2(n5783), .A3(n4511), .ZN(n5794) );
  NAND4_X1 U6366 ( .A1(n4511), .A2(n4774), .A3(n4775), .A4(n5783), .ZN(n5966)
         );
  AND2_X2 U6367 ( .A1(n5004), .A2(n5003), .ZN(n4939) );
  AND3_X2 U6368 ( .A1(n4779), .A2(n4778), .A3(n5107), .ZN(n5004) );
  NAND2_X1 U6369 ( .A1(n10032), .A2(n4780), .ZN(n4782) );
  INV_X1 U6370 ( .A(n7344), .ZN(n4781) );
  NAND2_X1 U6371 ( .A1(n4789), .A2(n4787), .ZN(n5695) );
  OR2_X1 U6372 ( .A1(n9632), .A2(n5704), .ZN(n4790) );
  NAND2_X1 U6373 ( .A1(n9632), .A2(n4795), .ZN(n4794) );
  NOR2_X1 U6374 ( .A1(n8673), .A2(n9889), .ZN(n4797) );
  NAND2_X1 U6375 ( .A1(n9694), .A2(n4507), .ZN(n4798) );
  NAND2_X1 U6376 ( .A1(n4798), .A2(n4799), .ZN(n9664) );
  INV_X1 U6377 ( .A(n7586), .ZN(n4808) );
  NAND2_X1 U6378 ( .A1(n4803), .A2(n4804), .ZN(n9785) );
  NAND2_X1 U6379 ( .A1(n7586), .A2(n4506), .ZN(n4803) );
  NAND2_X1 U6380 ( .A1(n9776), .A2(n4816), .ZN(n4815) );
  OAI21_X1 U6381 ( .B1(n9776), .B2(n4817), .A(n4816), .ZN(n9727) );
  NAND2_X1 U6382 ( .A1(n4825), .A2(n4826), .ZN(n9932) );
  NOR2_X1 U6383 ( .A1(n5442), .A2(n4827), .ZN(n5447) );
  NAND2_X1 U6384 ( .A1(n5502), .A2(n5501), .ZN(n7266) );
  NAND2_X1 U6385 ( .A1(n9152), .A2(n8646), .ZN(n8761) );
  NAND2_X1 U6386 ( .A1(n4838), .A2(n5222), .ZN(n5225) );
  OAI21_X2 U6387 ( .B1(n8680), .B2(n8681), .A(n8678), .ZN(n8577) );
  NAND2_X1 U6388 ( .A1(n9206), .A2(n8581), .ZN(n8770) );
  NAND2_X1 U6389 ( .A1(n4927), .A2(n4925), .ZN(n4924) );
  NAND2_X1 U6390 ( .A1(n5728), .A2(n7280), .ZN(n5502) );
  NAND2_X1 U6391 ( .A1(n6589), .A2(n7971), .ZN(n6588) );
  NAND2_X1 U6392 ( .A1(n8311), .A2(n8094), .ZN(n6368) );
  OAI21_X1 U6393 ( .B1(n7528), .B2(n7527), .A(n8036), .ZN(n7674) );
  NAND2_X1 U6394 ( .A1(n7417), .A2(n6301), .ZN(n4997) );
  OAI21_X1 U6395 ( .B1(n7435), .B2(n5583), .A(n5582), .ZN(n7495) );
  NAND2_X1 U6396 ( .A1(n10276), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n10275) );
  XNOR2_X1 U6397 ( .A(n5881), .B(n10341), .ZN(n10343) );
  NAND2_X1 U6398 ( .A1(n5622), .A2(n5621), .ZN(n9776) );
  NAND2_X1 U6399 ( .A1(n6368), .A2(n7936), .ZN(n6367) );
  OAI21_X1 U6400 ( .B1(n9601), .B2(n4831), .A(n9600), .ZN(n4943) );
  NAND2_X1 U6401 ( .A1(n5375), .A2(n5374), .ZN(n4832) );
  NAND2_X1 U6402 ( .A1(n5362), .A2(n5361), .ZN(n5367) );
  NAND2_X1 U6403 ( .A1(n5410), .A2(n5409), .ZN(n4833) );
  NAND2_X1 U6404 ( .A1(n5404), .A2(n5403), .ZN(n4834) );
  MUX2_X1 U6405 ( .A(n7137), .B(n8883), .S(n4835), .Z(n5322) );
  MUX2_X1 U6406 ( .A(n7368), .B(n7384), .S(n4835), .Z(n5344) );
  MUX2_X1 U6407 ( .A(n8913), .B(n7573), .S(n4835), .Z(n5358) );
  MUX2_X1 U6408 ( .A(n7804), .B(n7777), .S(n4835), .Z(n5388) );
  MUX2_X1 U6409 ( .A(n7818), .B(n6272), .S(n4835), .Z(n5412) );
  NAND2_X1 U6410 ( .A1(n5221), .A2(n5220), .ZN(n4838) );
  NAND2_X1 U6411 ( .A1(n4838), .A2(n4556), .ZN(n5229) );
  OAI21_X1 U6412 ( .B1(n5335), .B2(n5334), .A(n5333), .ZN(n5340) );
  NAND2_X1 U6413 ( .A1(n4855), .A2(n4856), .ZN(n5309) );
  NAND2_X1 U6414 ( .A1(n5275), .A2(n4858), .ZN(n4855) );
  OAI21_X1 U6415 ( .B1(n5239), .B2(n5238), .A(n5240), .ZN(n5249) );
  OAI21_X1 U6416 ( .B1(n5239), .B2(n4866), .A(n4865), .ZN(n5259) );
  NOR2_X1 U6417 ( .A1(n4883), .A2(n4882), .ZN(n10284) );
  NAND2_X1 U6418 ( .A1(n10301), .A2(n4895), .ZN(n4891) );
  NAND2_X1 U6419 ( .A1(n4891), .A2(n4893), .ZN(n10333) );
  NAND2_X1 U6420 ( .A1(n10350), .A2(n4902), .ZN(n4901) );
  OAI211_X1 U6421 ( .C1(n10350), .C2(n4905), .A(n4903), .B(n4901), .ZN(n5921)
         );
  NAND2_X1 U6422 ( .A1(n10350), .A2(n4909), .ZN(n9943) );
  AOI21_X1 U6423 ( .B1(n10350), .B2(n5918), .A(n5919), .ZN(n9942) );
  INV_X2 U6424 ( .A(n8627), .ZN(n8655) );
  NAND2_X4 U6425 ( .A1(n6530), .A2(n6525), .ZN(n8627) );
  XNOR2_X2 U6426 ( .A(n5458), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5468) );
  NOR2_X1 U6427 ( .A1(n9544), .A2(n9545), .ZN(n9548) );
  NAND2_X1 U6428 ( .A1(n5129), .A2(n4916), .ZN(n5152) );
  NAND2_X1 U6429 ( .A1(n6924), .A2(n6925), .ZN(n7044) );
  OAI211_X1 U6430 ( .C1(n7043), .C2(n4918), .A(n4917), .B(n7226), .ZN(n7234)
         );
  AOI21_X1 U6431 ( .B1(n7661), .B2(n4920), .A(n5077), .ZN(n4919) );
  NAND2_X1 U6432 ( .A1(n7661), .A2(n4927), .ZN(n4921) );
  INV_X1 U6433 ( .A(n4922), .ZN(n8569) );
  OAI21_X1 U6434 ( .B1(n7637), .B2(n7636), .A(n7635), .ZN(n7683) );
  AND2_X1 U6435 ( .A1(n5163), .A2(n4938), .ZN(n4937) );
  NAND3_X1 U6436 ( .A1(n8578), .A2(n8581), .A3(n8580), .ZN(n9206) );
  NAND2_X1 U6437 ( .A1(n8578), .A2(n8581), .ZN(n9208) );
  NAND2_X1 U6438 ( .A1(n5805), .A2(n4949), .ZN(n4948) );
  XNOR2_X1 U6439 ( .A(n6331), .B(P2_B_REG_SCAN_IN), .ZN(n4972) );
  NAND2_X1 U6440 ( .A1(n4975), .A2(n6688), .ZN(n4979) );
  NAND3_X1 U6441 ( .A1(n4562), .A2(n8119), .A3(n4982), .ZN(n4981) );
  NAND3_X1 U6442 ( .A1(n5100), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4994) );
  NAND2_X1 U6443 ( .A1(n4997), .A2(n4996), .ZN(n6304) );
  AND2_X1 U6444 ( .A1(n6303), .A2(n6302), .ZN(n4996) );
  NAND2_X1 U6445 ( .A1(n6308), .A2(n4998), .ZN(n8308) );
  NAND2_X1 U6446 ( .A1(n8308), .A2(n6310), .ZN(n8311) );
  NAND2_X1 U6447 ( .A1(n8381), .A2(n7939), .ZN(n6307) );
  OR2_X1 U6448 ( .A1(n7191), .A2(n6300), .ZN(n7140) );
  NAND2_X1 U6449 ( .A1(n7946), .A2(n7951), .ZN(n7918) );
  NAND2_X1 U6450 ( .A1(n5177), .A2(n5004), .ZN(n5291) );
  NAND2_X1 U6451 ( .A1(n4570), .A2(n5005), .ZN(n5080) );
  NAND2_X1 U6452 ( .A1(n5295), .A2(n5007), .ZN(n9732) );
  INV_X1 U6453 ( .A(n5010), .ZN(n9764) );
  INV_X1 U6454 ( .A(n9333), .ZN(n5011) );
  INV_X1 U6455 ( .A(n9327), .ZN(n5018) );
  NAND2_X1 U6456 ( .A1(n5019), .A2(n5015), .ZN(n5014) );
  NOR2_X1 U6457 ( .A1(n7793), .A2(n9810), .ZN(n9607) );
  NAND2_X1 U6458 ( .A1(n5440), .A2(n4560), .ZN(n5119) );
  INV_X1 U6459 ( .A(n5027), .ZN(n9655) );
  INV_X1 U6460 ( .A(n5033), .ZN(n7712) );
  OAI21_X2 U6461 ( .B1(n8336), .B2(n8335), .A(n5044), .ZN(n8324) );
  NAND2_X1 U6462 ( .A1(n5045), .A2(n6389), .ZN(n6391) );
  NAND2_X1 U6463 ( .A1(n7807), .A2(n5046), .ZN(n5045) );
  AND2_X1 U6464 ( .A1(n6330), .A2(n10430), .ZN(n5046) );
  NAND2_X1 U6465 ( .A1(n5047), .A2(n10446), .ZN(n6359) );
  OAI21_X2 U6466 ( .B1(n8385), .B2(n5052), .A(n5050), .ZN(n8348) );
  NAND2_X1 U6467 ( .A1(n5049), .A2(n5054), .ZN(n8359) );
  NAND2_X1 U6468 ( .A1(n8385), .A2(n5055), .ZN(n5049) );
  AOI21_X1 U6469 ( .B1(n5054), .B2(n5051), .A(n4564), .ZN(n5050) );
  NOR2_X1 U6470 ( .A1(n5055), .A2(n6228), .ZN(n5051) );
  NAND2_X1 U6471 ( .A1(n5054), .A2(n5053), .ZN(n5052) );
  NAND2_X1 U6472 ( .A1(n5060), .A2(n5058), .ZN(n6151) );
  OR2_X1 U6473 ( .A1(n7751), .A2(n8276), .ZN(n5063) );
  NAND2_X1 U6474 ( .A1(n5065), .A2(n5064), .ZN(n7182) );
  NAND3_X1 U6475 ( .A1(n6078), .A2(n6077), .A3(n4565), .ZN(n5065) );
  NAND2_X1 U6476 ( .A1(n5067), .A2(n5066), .ZN(n5970) );
  INV_X1 U6477 ( .A(n5794), .ZN(n5067) );
  NAND2_X1 U6478 ( .A1(n6187), .A2(n5071), .ZN(n5070) );
  NAND2_X1 U6479 ( .A1(n6187), .A2(n6186), .ZN(n8408) );
  INV_X1 U6480 ( .A(n5070), .ZN(n8411) );
  INV_X1 U6481 ( .A(n6186), .ZN(n5072) );
  AND2_X1 U6482 ( .A1(n6710), .A2(n6713), .ZN(n10384) );
  INV_X1 U6483 ( .A(n5515), .ZN(n10118) );
  NAND2_X1 U6484 ( .A1(n5732), .A2(n9385), .ZN(n7262) );
  NOR2_X1 U6485 ( .A1(n8299), .A2(n6365), .ZN(n6381) );
  NAND2_X1 U6486 ( .A1(n7778), .A2(n5725), .ZN(n7881) );
  NAND2_X1 U6487 ( .A1(n6651), .A2(n6648), .ZN(n6667) );
  INV_X1 U6488 ( .A(n7312), .ZN(n5176) );
  NAND2_X1 U6489 ( .A1(n6452), .A2(n6451), .ZN(n6467) );
  OR2_X1 U6490 ( .A1(n6452), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6335) );
  NAND2_X1 U6491 ( .A1(n5162), .A2(n10125), .ZN(n7312) );
  INV_X1 U6492 ( .A(n7311), .ZN(n5162) );
  INV_X1 U6493 ( .A(n10416), .ZN(n6088) );
  INV_X1 U6494 ( .A(n5119), .ZN(n5121) );
  NAND2_X1 U6495 ( .A1(n5119), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5116) );
  NAND2_X1 U6496 ( .A1(n6717), .A2(n6673), .ZN(n6712) );
  NAND2_X1 U6497 ( .A1(n5975), .A2(n8553), .ZN(n6013) );
  NAND2_X1 U6498 ( .A1(n6304), .A2(n8029), .ZN(n7528) );
  OR2_X1 U6499 ( .A1(n5447), .A2(n9931), .ZN(n5118) );
  NAND2_X1 U6500 ( .A1(n5970), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5972) );
  AOI21_X2 U6501 ( .B1(n6240), .B2(n6239), .A(n6238), .ZN(n8336) );
  AND3_X2 U6502 ( .A1(n6355), .A2(n6354), .A3(n6353), .ZN(n10446) );
  INV_X1 U6503 ( .A(n8493), .ZN(n6369) );
  AND2_X1 U6504 ( .A1(n5503), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5073) );
  AND2_X1 U6505 ( .A1(n5527), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5074) );
  OR2_X1 U6506 ( .A1(n7211), .A2(n7210), .ZN(n5075) );
  AND2_X1 U6507 ( .A1(n7153), .A2(n7152), .ZN(n5076) );
  AND4_X1 U6508 ( .A1(n7906), .A2(n7905), .A3(n7904), .A4(n7903), .ZN(n8293)
         );
  OR2_X1 U6509 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5078) );
  AND2_X2 U6510 ( .A1(n5495), .A2(n7800), .ZN(n5079) );
  INV_X1 U6511 ( .A(n10341), .ZN(n6834) );
  INV_X1 U6512 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5798) );
  OR2_X1 U6513 ( .A1(n6327), .A2(n8128), .ZN(n10420) );
  OR2_X1 U6514 ( .A1(n6390), .A2(n8507), .ZN(n5081) );
  AND2_X1 U6515 ( .A1(n6683), .A2(n6942), .ZN(n5085) );
  NOR2_X1 U6516 ( .A1(n7835), .A2(n8148), .ZN(n5087) );
  AND2_X1 U6517 ( .A1(n6309), .A2(n8093), .ZN(n5088) );
  NOR2_X1 U6518 ( .A1(n6047), .A2(n7000), .ZN(n5089) );
  NAND2_X1 U6519 ( .A1(n10419), .A2(n7457), .ZN(n5090) );
  OR2_X1 U6520 ( .A1(n9462), .A2(n9325), .ZN(n5091) );
  INV_X1 U6521 ( .A(n6712), .ZN(n6296) );
  AND2_X1 U6522 ( .A1(n8107), .A2(n7890), .ZN(n5092) );
  INV_X1 U6523 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5786) );
  NAND2_X1 U6524 ( .A1(n6314), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5093) );
  INV_X1 U6525 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5106) );
  INV_X1 U6526 ( .A(SI_18_), .ZN(n5310) );
  INV_X1 U6527 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U6528 ( .A1(n5756), .A2(n9364), .ZN(n10054) );
  INV_X1 U6529 ( .A(n10192), .ZN(n5490) );
  OR2_X1 U6530 ( .A1(n9703), .A2(n9496), .ZN(n5094) );
  OR2_X1 U6531 ( .A1(n6886), .A2(n5863), .ZN(n5095) );
  INV_X1 U6532 ( .A(n10274), .ZN(n6497) );
  AND2_X1 U6533 ( .A1(n7836), .A2(n8202), .ZN(n5096) );
  INV_X1 U6534 ( .A(n8306), .ZN(n6370) );
  OR2_X1 U6535 ( .A1(n9671), .A2(n9494), .ZN(n5098) );
  NAND2_X1 U6536 ( .A1(n4765), .A2(n8112), .ZN(n8072) );
  AND2_X1 U6537 ( .A1(n8084), .A2(n8072), .ZN(n8073) );
  INV_X1 U6538 ( .A(n8075), .ZN(n8076) );
  NAND2_X1 U6539 ( .A1(n8077), .A2(n8076), .ZN(n8085) );
  INV_X1 U6540 ( .A(n8096), .ZN(n8097) );
  INV_X1 U6541 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5110) );
  AOI21_X1 U6542 ( .B1(n8098), .B2(n5088), .A(n8097), .ZN(n8099) );
  INV_X1 U6543 ( .A(n7686), .ZN(n7646) );
  NOR2_X1 U6544 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5113) );
  INV_X1 U6545 ( .A(n6649), .ZN(n6650) );
  OR2_X1 U6546 ( .A1(n8425), .A2(n6185), .ZN(n6187) );
  INV_X1 U6547 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9044) );
  AND2_X1 U6548 ( .A1(n8693), .A2(n9148), .ZN(n8635) );
  OAI22_X1 U6549 ( .A1(n8609), .A2(n5507), .B1(n6930), .B2(n8627), .ZN(n6762)
         );
  INV_X1 U6550 ( .A(n9409), .ZN(n5745) );
  AND3_X1 U6551 ( .A1(n5493), .A2(n5492), .A3(n5491), .ZN(n5500) );
  INV_X1 U6552 ( .A(n6691), .ZN(n6688) );
  INV_X1 U6553 ( .A(n6999), .ZN(n5850) );
  NOR2_X1 U6554 ( .A1(n6114), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6113) );
  OR2_X1 U6555 ( .A1(n8567), .A2(n8566), .ZN(n8568) );
  AND2_X1 U6556 ( .A1(n6528), .A2(n6527), .ZN(n6529) );
  OR2_X1 U6557 ( .A1(n5166), .A2(n6430), .ZN(n5138) );
  INV_X1 U6558 ( .A(n7436), .ZN(n5741) );
  INV_X1 U6559 ( .A(SI_29_), .ZN(n9107) );
  INV_X1 U6560 ( .A(SI_26_), .ZN(n5387) );
  INV_X1 U6561 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5311) );
  INV_X1 U6562 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5250) );
  INV_X1 U6563 ( .A(SI_8_), .ZN(n9092) );
  INV_X1 U6564 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5810) );
  NAND2_X1 U6565 ( .A1(n6702), .A2(n6754), .ZN(n6703) );
  AND2_X1 U6566 ( .A1(n6657), .A2(n6656), .ZN(n8244) );
  NAND2_X1 U6567 ( .A1(n6202), .A2(n6201), .ZN(n6211) );
  INV_X1 U6568 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n6272) );
  OR2_X1 U6569 ( .A1(n6221), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6231) );
  AND2_X1 U6570 ( .A1(n6190), .A2(n6189), .ZN(n6202) );
  AND2_X1 U6571 ( .A1(n6143), .A2(n5963), .ZN(n6154) );
  OR2_X1 U6572 ( .A1(n6093), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6102) );
  INV_X1 U6573 ( .A(n10420), .ZN(n6328) );
  OR2_X1 U6574 ( .A1(n6670), .A2(n6378), .ZN(n6624) );
  INV_X1 U6575 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8773) );
  AND2_X1 U6576 ( .A1(n5637), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5644) );
  OAI22_X1 U6577 ( .A1(n8736), .A2(n9141), .B1(n7789), .B2(n9371), .ZN(n7790)
         );
  INV_X1 U6578 ( .A(n9687), .ZN(n5677) );
  AND2_X1 U6579 ( .A1(n5567), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5576) );
  INV_X1 U6580 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5117) );
  AND2_X1 U6581 ( .A1(n5366), .A2(n5360), .ZN(n5361) );
  INV_X1 U6582 ( .A(SI_12_), .ZN(n9026) );
  NAND2_X1 U6583 ( .A1(n7108), .A2(n7058), .ZN(n7109) );
  OR2_X1 U6584 ( .A1(n6285), .A2(n7808), .ZN(n7906) );
  INV_X1 U6585 ( .A(n10350), .ZN(n10351) );
  AND2_X1 U6586 ( .A1(n5949), .A2(n8556), .ZN(n5946) );
  AND2_X1 U6587 ( .A1(n7808), .A2(n6278), .ZN(n8300) );
  AND2_X1 U6588 ( .A1(n6256), .A2(n6255), .ZN(n6264) );
  INV_X1 U6589 ( .A(n8413), .ZN(n8390) );
  INV_X1 U6590 ( .A(n8437), .ZN(n6306) );
  AND2_X1 U6591 ( .A1(n7944), .A2(n7948), .ZN(n8001) );
  AND2_X1 U6592 ( .A1(n6320), .A2(n6322), .ZN(n6656) );
  NAND2_X1 U6593 ( .A1(n6335), .A2(n6334), .ZN(n6665) );
  NAND2_X1 U6594 ( .A1(n6329), .A2(n6328), .ZN(n6330) );
  INV_X1 U6595 ( .A(n6321), .ZN(n8389) );
  INV_X1 U6596 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5801) );
  INV_X1 U6597 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5787) );
  OR2_X1 U6598 ( .A1(n5868), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5870) );
  INV_X1 U6599 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8683) );
  INV_X1 U6600 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7521) );
  NOR2_X1 U6601 ( .A1(n5624), .A2(n5623), .ZN(n5631) );
  AND2_X1 U6602 ( .A1(n5644), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5652) );
  NAND2_X1 U6603 ( .A1(n8625), .A2(n8693), .ZN(n8690) );
  OR2_X1 U6604 ( .A1(n8594), .A2(n8593), .ZN(n8595) );
  AND2_X1 U6605 ( .A1(n9193), .A2(n9194), .ZN(n8659) );
  AND2_X1 U6606 ( .A1(n5757), .A2(n5717), .ZN(n8740) );
  INV_X1 U6607 ( .A(n7790), .ZN(n7791) );
  AND2_X1 U6608 ( .A1(n9284), .A2(n9423), .ZN(n9743) );
  NAND2_X1 U6609 ( .A1(n9236), .A2(n5739), .ZN(n7344) );
  OR2_X1 U6610 ( .A1(n6527), .A2(n9720), .ZN(n10045) );
  INV_X1 U6611 ( .A(n9184), .ZN(n9195) );
  NAND2_X1 U6612 ( .A1(n9811), .A2(n5084), .ZN(n9812) );
  INV_X1 U6613 ( .A(n9218), .ZN(n9978) );
  INV_X1 U6614 ( .A(n7693), .ZN(n7645) );
  INV_X1 U6615 ( .A(n8713), .ZN(n10169) );
  INV_X1 U6616 ( .A(n10054), .ZN(n10036) );
  INV_X1 U6617 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5459) );
  AOI21_X1 U6618 ( .B1(n6685), .B2(n6684), .A(n5085), .ZN(n6758) );
  INV_X1 U6619 ( .A(n6704), .ZN(n6689) );
  INV_X1 U6620 ( .A(n8251), .ZN(n8242) );
  AND2_X1 U6621 ( .A1(n6271), .A2(n6270), .ZN(n8327) );
  AND3_X1 U6622 ( .A1(n6184), .A2(n6183), .A3(n6182), .ZN(n8154) );
  MUX2_X1 U6623 ( .A(n8283), .B(n5950), .S(n5886), .Z(n10340) );
  OR2_X1 U6624 ( .A1(n6264), .A2(n6257), .ZN(n8330) );
  INV_X1 U6625 ( .A(n6736), .ZN(n10394) );
  OR2_X1 U6626 ( .A1(n6623), .A2(n6603), .ZN(n10373) );
  INV_X1 U6627 ( .A(n8451), .ZN(n8473) );
  NOR2_X1 U6628 ( .A1(n6663), .A2(n6352), .ZN(n6354) );
  INV_X1 U6629 ( .A(n8441), .ZN(n8496) );
  NAND2_X1 U6630 ( .A1(n7493), .A2(n7963), .ZN(n10418) );
  AND2_X1 U6631 ( .A1(n8036), .A2(n8040), .ZN(n8034) );
  AND2_X1 U6632 ( .A1(n7252), .A2(n7253), .ZN(n7285) );
  INV_X1 U6633 ( .A(n10418), .ZN(n10429) );
  NAND2_X1 U6634 ( .A1(n7200), .A2(n10420), .ZN(n10408) );
  XNOR2_X1 U6635 ( .A(n5800), .B(n5801), .ZN(n5951) );
  AOI21_X1 U6636 ( .B1(P1_REG1_REG_0__SCAN_IN), .B2(n6532), .A(n6630), .ZN(
        n6632) );
  AND2_X1 U6637 ( .A1(n6546), .A2(n6545), .ZN(n9960) );
  AND4_X1 U6638 ( .A1(n5676), .A2(n5675), .A3(n5674), .A4(n5673), .ZN(n9171)
         );
  AND4_X1 U6639 ( .A1(n5620), .A2(n5619), .A3(n5618), .A4(n5617), .ZN(n9142)
         );
  INV_X1 U6640 ( .A(n10017), .ZN(n9993) );
  INV_X1 U6641 ( .A(n10043), .ZN(n10058) );
  INV_X1 U6642 ( .A(n9803), .ZN(n10067) );
  INV_X1 U6643 ( .A(n10168), .ZN(n5959) );
  OR2_X1 U6644 ( .A1(n6538), .A2(n6545), .ZN(n6540) );
  INV_X1 U6645 ( .A(n5475), .ZN(n6849) );
  NAND2_X1 U6646 ( .A1(n6530), .A2(n7576), .ZN(n6926) );
  INV_X1 U6647 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5438) );
  INV_X1 U6648 ( .A(n6627), .ZN(n5802) );
  INV_X1 U6649 ( .A(n6673), .ZN(n6654) );
  INV_X1 U6650 ( .A(n8331), .ZN(n8508) );
  INV_X1 U6651 ( .A(n8327), .ZN(n8272) );
  INV_X1 U6652 ( .A(n8202), .ZN(n8426) );
  INV_X1 U6653 ( .A(n8020), .ZN(n8277) );
  OR2_X1 U6654 ( .A1(P2_U3150), .A2(n5952), .ZN(n10200) );
  NAND2_X1 U6655 ( .A1(P2_U3893), .A2(n5886), .ZN(n10354) );
  NAND2_X1 U6656 ( .A1(n4495), .A2(n10362), .ZN(n8407) );
  NAND2_X1 U6657 ( .A1(n10446), .A2(n10408), .ZN(n8493) );
  INV_X1 U6658 ( .A(n10446), .ZN(n10444) );
  OR2_X1 U6659 ( .A1(n10432), .A2(n10424), .ZN(n8544) );
  AND2_X1 U6660 ( .A1(n6380), .A2(n6379), .ZN(n10432) );
  INV_X1 U6661 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7886) );
  INV_X1 U6662 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n9038) );
  INV_X1 U6663 ( .A(n10290), .ZN(n6522) );
  AND2_X1 U6664 ( .A1(n6929), .A2(n6928), .ZN(n9970) );
  INV_X1 U6665 ( .A(n9217), .ZN(n9963) );
  AND4_X1 U6666 ( .A1(n5721), .A2(n5720), .A3(n5719), .A4(n5718), .ZN(n8736)
         );
  OR2_X1 U6667 ( .A1(n6530), .A2(n6392), .ZN(n9504) );
  OR2_X1 U6668 ( .A1(n6415), .A2(n6414), .ZN(n9601) );
  OR2_X1 U6669 ( .A1(n10070), .A2(n7171), .ZN(n9800) );
  OR2_X1 U6670 ( .A1(n10070), .A2(n7265), .ZN(n9803) );
  AND2_X1 U6671 ( .A1(n7170), .A2(n10056), .ZN(n10043) );
  NAND2_X1 U6672 ( .A1(n10192), .A2(n5959), .ZN(n9875) );
  AND3_X2 U6673 ( .A1(n6465), .A2(n5957), .A3(n6540), .ZN(n10192) );
  NAND2_X1 U6674 ( .A1(n8745), .A2(n6387), .ZN(n5960) );
  INV_X1 U6675 ( .A(n9703), .ZN(n9905) );
  INV_X1 U6676 ( .A(n9263), .ZN(n9930) );
  INV_X1 U6677 ( .A(n10175), .ZN(n10173) );
  AND3_X2 U6678 ( .A1(n5957), .A2(n9475), .A3(n7168), .ZN(n10175) );
  NOR2_X1 U6679 ( .A1(n6850), .A2(n6849), .ZN(n10084) );
  CLKBUF_X1 U6680 ( .A(n10084), .Z(n10102) );
  INV_X1 U6681 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7801) );
  INV_X1 U6682 ( .A(n5467), .ZN(n7621) );
  INV_X1 U6683 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7137) );
  NOR2_X2 U6684 ( .A1(n6374), .A2(n5802), .ZN(P2_U3893) );
  NAND2_X1 U6685 ( .A1(n5961), .A2(n5960), .ZN(P1_U3518) );
  INV_X1 U6686 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5099) );
  INV_X1 U6687 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5100) );
  INV_X1 U6688 ( .A(SI_0_), .ZN(n5102) );
  INV_X1 U6689 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5101) );
  OAI21_X1 U6690 ( .B1(n4835), .B2(n5102), .A(n5101), .ZN(n5104) );
  AND2_X1 U6691 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5103) );
  NAND2_X1 U6692 ( .A1(n4498), .A2(n5103), .ZN(n5126) );
  AND2_X1 U6693 ( .A1(n5104), .A2(n5126), .ZN(n9937) );
  INV_X2 U6694 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5267) );
  NAND4_X1 U6695 ( .A1(n5250), .A2(n5109), .A3(n5267), .A4(n5108), .ZN(n5111)
         );
  INV_X1 U6696 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6423) );
  OR2_X1 U6697 ( .A1(n5173), .A2(n6423), .ZN(n5493) );
  NAND3_X1 U6698 ( .A1(n5124), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n5125) );
  NAND2_X1 U6699 ( .A1(n5126), .A2(n5125), .ZN(n5131) );
  XNOR2_X1 U6700 ( .A(n5132), .B(n5131), .ZN(n6444) );
  NAND2_X1 U6701 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5128) );
  NAND2_X1 U6702 ( .A1(n5140), .A2(n6422), .ZN(n5491) );
  NAND2_X1 U6703 ( .A1(n7275), .A2(n10104), .ZN(n7274) );
  OR2_X1 U6704 ( .A1(n5129), .A2(n9931), .ZN(n5130) );
  XNOR2_X1 U6705 ( .A(n5130), .B(P1_IR_REG_2__SCAN_IN), .ZN(n10001) );
  INV_X1 U6706 ( .A(n10001), .ZN(n6424) );
  INV_X1 U6707 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6425) );
  OR2_X1 U6708 ( .A1(n5173), .A2(n6425), .ZN(n5139) );
  NAND2_X1 U6709 ( .A1(n5132), .A2(n5131), .ZN(n5136) );
  INV_X1 U6710 ( .A(n5133), .ZN(n5134) );
  NAND2_X1 U6711 ( .A1(n5134), .A2(SI_1_), .ZN(n5135) );
  INV_X1 U6712 ( .A(SI_2_), .ZN(n5137) );
  XNOR2_X1 U6713 ( .A(n5145), .B(n5137), .ZN(n5143) );
  XNOR2_X1 U6714 ( .A(n5144), .B(n5143), .ZN(n6430) );
  OAI211_X1 U6715 ( .C1(n5127), .C2(n6424), .A(n5139), .B(n5138), .ZN(n6763)
         );
  NAND2_X1 U6716 ( .A1(n5141), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5142) );
  XNOR2_X1 U6717 ( .A(n5142), .B(n5106), .ZN(n6426) );
  INV_X1 U6718 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6427) );
  OR2_X1 U6719 ( .A1(n5173), .A2(n6427), .ZN(n5150) );
  NAND2_X1 U6720 ( .A1(n5144), .A2(n5143), .ZN(n5147) );
  NAND2_X1 U6721 ( .A1(n5145), .A2(SI_2_), .ZN(n5146) );
  NAND2_X1 U6722 ( .A1(n5147), .A2(n5146), .ZN(n5155) );
  INV_X1 U6723 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6432) );
  XNOR2_X1 U6724 ( .A(n5156), .B(SI_3_), .ZN(n5154) );
  XNOR2_X1 U6725 ( .A(n5155), .B(n5154), .ZN(n6431) );
  OR2_X1 U6726 ( .A1(n5166), .A2(n6431), .ZN(n5149) );
  OAI211_X1 U6727 ( .C1(n5151), .C2(n6426), .A(n5150), .B(n5149), .ZN(n5515)
         );
  NAND2_X1 U6728 ( .A1(n10064), .A2(n10118), .ZN(n7311) );
  NAND2_X1 U6729 ( .A1(n5152), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5153) );
  XNOR2_X1 U6730 ( .A(n5153), .B(P1_IR_REG_4__SCAN_IN), .ZN(n10024) );
  INV_X1 U6731 ( .A(n10024), .ZN(n6428) );
  INV_X1 U6732 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6429) );
  OR2_X1 U6733 ( .A1(n5173), .A2(n6429), .ZN(n5161) );
  NAND2_X1 U6734 ( .A1(n5155), .A2(n5154), .ZN(n5159) );
  INV_X1 U6735 ( .A(n5156), .ZN(n5157) );
  NAND2_X1 U6736 ( .A1(n5157), .A2(SI_3_), .ZN(n5158) );
  NAND2_X1 U6737 ( .A1(n5159), .A2(n5158), .ZN(n5168) );
  INV_X1 U6738 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6434) );
  MUX2_X1 U6739 ( .A(n6434), .B(n6429), .S(n4500), .Z(n5169) );
  XNOR2_X1 U6740 ( .A(n5169), .B(SI_4_), .ZN(n5167) );
  XNOR2_X1 U6741 ( .A(n5168), .B(n5167), .ZN(n6433) );
  OR2_X1 U6742 ( .A1(n5166), .A2(n6433), .ZN(n5160) );
  OR2_X1 U6743 ( .A1(n5163), .A2(n9931), .ZN(n5165) );
  XNOR2_X1 U6744 ( .A(n5165), .B(n5164), .ZN(n6435) );
  NAND2_X1 U6745 ( .A1(n5168), .A2(n5167), .ZN(n5172) );
  INV_X1 U6746 ( .A(n5169), .ZN(n5170) );
  NAND2_X1 U6747 ( .A1(n5170), .A2(SI_4_), .ZN(n5171) );
  XNOR2_X1 U6748 ( .A(n5180), .B(SI_5_), .ZN(n5178) );
  XNOR2_X1 U6749 ( .A(n5179), .B(n5178), .ZN(n6438) );
  OR2_X1 U6750 ( .A1(n5166), .A2(n6438), .ZN(n5175) );
  OR2_X1 U6751 ( .A1(n5173), .A2(n6436), .ZN(n5174) );
  OR2_X1 U6752 ( .A1(n5177), .A2(n9931), .ZN(n5187) );
  XNOR2_X1 U6753 ( .A(n5187), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6825) );
  INV_X1 U6754 ( .A(n6825), .ZN(n6440) );
  INV_X1 U6755 ( .A(n5180), .ZN(n5181) );
  NAND2_X1 U6756 ( .A1(n5181), .A2(SI_5_), .ZN(n5182) );
  MUX2_X1 U6757 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n4498), .Z(n5193) );
  INV_X1 U6758 ( .A(SI_6_), .ZN(n5183) );
  XNOR2_X1 U6759 ( .A(n5193), .B(n5183), .ZN(n5191) );
  XNOR2_X1 U6760 ( .A(n5192), .B(n5191), .ZN(n6443) );
  OR2_X1 U6761 ( .A1(n5166), .A2(n6443), .ZN(n5185) );
  INV_X1 U6762 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6441) );
  OR2_X1 U6763 ( .A1(n5173), .A2(n6441), .ZN(n5184) );
  INV_X1 U6764 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U6765 ( .A1(n5187), .A2(n5186), .ZN(n5188) );
  NAND2_X1 U6766 ( .A1(n5188), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5190) );
  INV_X1 U6767 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5189) );
  XNOR2_X1 U6768 ( .A(n5190), .B(n5189), .ZN(n6554) );
  MUX2_X1 U6769 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n4500), .Z(n5201) );
  INV_X1 U6770 ( .A(SI_7_), .ZN(n5194) );
  XNOR2_X1 U6771 ( .A(n5201), .B(n5194), .ZN(n5199) );
  XNOR2_X1 U6772 ( .A(n5200), .B(n5199), .ZN(n6446) );
  OR2_X1 U6773 ( .A1(n5166), .A2(n6446), .ZN(n5196) );
  INV_X1 U6774 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6447) );
  OR2_X1 U6775 ( .A1(n5173), .A2(n6447), .ZN(n5195) );
  OAI211_X1 U6776 ( .C1(n5151), .C2(n6554), .A(n5196), .B(n5195), .ZN(n10044)
         );
  NAND2_X1 U6777 ( .A1(n5197), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5198) );
  XNOR2_X1 U6778 ( .A(n5198), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6812) );
  INV_X1 U6779 ( .A(n6812), .ZN(n6448) );
  INV_X1 U6780 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6450) );
  MUX2_X1 U6781 ( .A(n9062), .B(n6450), .S(n4499), .Z(n5202) );
  NAND2_X1 U6782 ( .A1(n5202), .A2(n9092), .ZN(n5211) );
  INV_X1 U6783 ( .A(n5202), .ZN(n5203) );
  NAND2_X1 U6784 ( .A1(n5203), .A2(SI_8_), .ZN(n5204) );
  NAND2_X1 U6785 ( .A1(n5211), .A2(n5204), .ZN(n5209) );
  INV_X1 U6786 ( .A(n5209), .ZN(n5205) );
  XNOR2_X1 U6787 ( .A(n5210), .B(n5205), .ZN(n6449) );
  OR2_X1 U6788 ( .A1(n5166), .A2(n6449), .ZN(n5207) );
  OR2_X1 U6789 ( .A1(n5173), .A2(n6450), .ZN(n5206) );
  OAI211_X1 U6790 ( .C1(n5151), .C2(n6448), .A(n5207), .B(n5206), .ZN(n7510)
         );
  OR2_X1 U6791 ( .A1(n5197), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5217) );
  NAND2_X1 U6792 ( .A1(n5217), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5208) );
  XNOR2_X1 U6793 ( .A(n5208), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6785) );
  INV_X1 U6794 ( .A(n6785), .ZN(n6567) );
  INV_X1 U6795 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6457) );
  MUX2_X1 U6796 ( .A(n6457), .B(n6459), .S(n4499), .Z(n5213) );
  INV_X1 U6797 ( .A(SI_9_), .ZN(n5212) );
  NAND2_X1 U6798 ( .A1(n5213), .A2(n5212), .ZN(n5222) );
  INV_X1 U6799 ( .A(n5213), .ZN(n5214) );
  NAND2_X1 U6800 ( .A1(n5214), .A2(SI_9_), .ZN(n5215) );
  NAND2_X1 U6801 ( .A1(n5222), .A2(n5215), .ZN(n5219) );
  OR2_X1 U6802 ( .A1(n5173), .A2(n6459), .ZN(n5216) );
  NAND2_X1 U6803 ( .A1(n5234), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5218) );
  XNOR2_X1 U6804 ( .A(n5218), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7071) );
  AOI22_X1 U6805 ( .A1(n5406), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5330), .B2(
        n7071), .ZN(n5224) );
  INV_X1 U6806 ( .A(n5219), .ZN(n5220) );
  MUX2_X1 U6807 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n4499), .Z(n5227) );
  INV_X1 U6808 ( .A(SI_10_), .ZN(n5223) );
  XNOR2_X1 U6809 ( .A(n5227), .B(n5223), .ZN(n5226) );
  NAND2_X1 U6810 ( .A1(n5227), .A2(SI_10_), .ZN(n5228) );
  INV_X1 U6811 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5230) );
  MUX2_X1 U6812 ( .A(n6484), .B(n5230), .S(n4500), .Z(n5231) );
  NAND2_X1 U6813 ( .A1(n5231), .A2(n9066), .ZN(n5240) );
  INV_X1 U6814 ( .A(n5231), .ZN(n5232) );
  NAND2_X1 U6815 ( .A1(n5232), .A2(SI_11_), .ZN(n5233) );
  NAND2_X1 U6816 ( .A1(n5240), .A2(n5233), .ZN(n5238) );
  NAND2_X1 U6817 ( .A1(n6480), .A2(n5434), .ZN(n5237) );
  NOR2_X1 U6818 ( .A1(n5234), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5242) );
  OR2_X1 U6819 ( .A1(n5242), .A2(n9931), .ZN(n5235) );
  XNOR2_X1 U6820 ( .A(n5235), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7123) );
  AOI22_X1 U6821 ( .A1(n5406), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5330), .B2(
        n7123), .ZN(n5236) );
  MUX2_X1 U6822 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n4500), .Z(n5247) );
  XNOR2_X1 U6823 ( .A(n5247), .B(n9026), .ZN(n5246) );
  XNOR2_X1 U6824 ( .A(n5249), .B(n5246), .ZN(n6486) );
  NAND2_X1 U6825 ( .A1(n6486), .A2(n5434), .ZN(n5245) );
  NAND2_X1 U6826 ( .A1(n5242), .A2(n5241), .ZN(n5243) );
  NAND2_X1 U6827 ( .A1(n5243), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5266) );
  XNOR2_X1 U6828 ( .A(n5266), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7374) );
  AOI22_X1 U6829 ( .A1(n5406), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5330), .B2(
        n7374), .ZN(n5244) );
  INV_X1 U6830 ( .A(n5246), .ZN(n5248) );
  MUX2_X1 U6831 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n4500), .Z(n5257) );
  XNOR2_X1 U6832 ( .A(n5257), .B(SI_13_), .ZN(n5255) );
  XNOR2_X1 U6833 ( .A(n5256), .B(n5255), .ZN(n6496) );
  NAND2_X1 U6834 ( .A1(n6496), .A2(n5434), .ZN(n5254) );
  NAND2_X1 U6835 ( .A1(n5266), .A2(n5250), .ZN(n5251) );
  NAND2_X1 U6836 ( .A1(n5251), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5252) );
  XNOR2_X1 U6837 ( .A(n5252), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7482) );
  AOI22_X1 U6838 ( .A1(n5406), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5330), .B2(
        n7482), .ZN(n5253) );
  NAND2_X1 U6839 ( .A1(n5257), .A2(SI_13_), .ZN(n5258) );
  NAND2_X1 U6840 ( .A1(n5259), .A2(n5258), .ZN(n5270) );
  INV_X1 U6841 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n5260) );
  MUX2_X1 U6842 ( .A(n6524), .B(n5260), .S(n4499), .Z(n5262) );
  INV_X1 U6843 ( .A(SI_14_), .ZN(n5261) );
  NAND2_X1 U6844 ( .A1(n5262), .A2(n5261), .ZN(n5274) );
  INV_X1 U6845 ( .A(n5262), .ZN(n5263) );
  NAND2_X1 U6846 ( .A1(n5263), .A2(SI_14_), .ZN(n5264) );
  NAND2_X1 U6847 ( .A1(n5274), .A2(n5264), .ZN(n5271) );
  XNOR2_X1 U6848 ( .A(n5270), .B(n5271), .ZN(n6516) );
  NAND2_X1 U6849 ( .A1(n6516), .A2(n5434), .ZN(n5269) );
  OAI21_X1 U6850 ( .B1(P1_IR_REG_12__SCAN_IN), .B2(P1_IR_REG_13__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5265) );
  NAND2_X1 U6851 ( .A1(n5266), .A2(n5265), .ZN(n5276) );
  XNOR2_X1 U6852 ( .A(n5276), .B(n5267), .ZN(n7767) );
  AOI22_X1 U6853 ( .A1(n5406), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5330), .B2(
        n7767), .ZN(n5268) );
  INV_X1 U6854 ( .A(n5270), .ZN(n5273) );
  INV_X1 U6855 ( .A(n5271), .ZN(n5272) );
  NAND2_X1 U6856 ( .A1(n5273), .A2(n5272), .ZN(n5275) );
  MUX2_X1 U6857 ( .A(n9103), .B(n6600), .S(n4500), .Z(n5282) );
  XNOR2_X1 U6858 ( .A(n5282), .B(SI_15_), .ZN(n5281) );
  XNOR2_X1 U6859 ( .A(n5286), .B(n5281), .ZN(n6599) );
  NAND2_X1 U6860 ( .A1(n6599), .A2(n5434), .ZN(n5280) );
  OAI21_X1 U6861 ( .B1(n5276), .B2(P1_IR_REG_14__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5278) );
  XNOR2_X1 U6862 ( .A(n5278), .B(n5277), .ZN(n9542) );
  INV_X1 U6863 ( .A(n9542), .ZN(n7769) );
  AOI22_X1 U6864 ( .A1(n5406), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5330), .B2(
        n7769), .ZN(n5279) );
  NAND2_X1 U6865 ( .A1(n7726), .A2(n9978), .ZN(n9795) );
  INV_X1 U6866 ( .A(n5281), .ZN(n5285) );
  INV_X1 U6867 ( .A(n5282), .ZN(n5283) );
  NAND2_X1 U6868 ( .A1(n5283), .A2(SI_15_), .ZN(n5284) );
  INV_X1 U6869 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5287) );
  MUX2_X1 U6870 ( .A(n6833), .B(n5287), .S(n4499), .Z(n5288) );
  NAND2_X1 U6871 ( .A1(n5288), .A2(n9064), .ZN(n5296) );
  INV_X1 U6872 ( .A(n5288), .ZN(n5289) );
  NAND2_X1 U6873 ( .A1(n5289), .A2(SI_16_), .ZN(n5290) );
  NAND2_X1 U6874 ( .A1(n5296), .A2(n5290), .ZN(n5297) );
  XNOR2_X1 U6875 ( .A(n5298), .B(n5297), .ZN(n6723) );
  NAND2_X1 U6876 ( .A1(n6723), .A2(n5434), .ZN(n5294) );
  NAND2_X1 U6877 ( .A1(n5291), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5292) );
  XNOR2_X1 U6878 ( .A(n5292), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9561) );
  AOI22_X1 U6879 ( .A1(n5406), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5330), .B2(
        n9561), .ZN(n5293) );
  INV_X1 U6880 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5299) );
  MUX2_X1 U6881 ( .A(n6836), .B(n5299), .S(n4500), .Z(n5301) );
  NAND2_X1 U6882 ( .A1(n5301), .A2(n5300), .ZN(n5308) );
  INV_X1 U6883 ( .A(n5301), .ZN(n5302) );
  NAND2_X1 U6884 ( .A1(n5302), .A2(SI_17_), .ZN(n5303) );
  XNOR2_X1 U6885 ( .A(n5307), .B(n5306), .ZN(n6779) );
  NAND2_X1 U6886 ( .A1(n6779), .A2(n5434), .ZN(n5305) );
  XNOR2_X1 U6887 ( .A(n5312), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9578) );
  AOI22_X1 U6888 ( .A1(n5406), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5330), .B2(
        n9578), .ZN(n5304) );
  NAND2_X1 U6889 ( .A1(n5309), .A2(n5308), .ZN(n5320) );
  MUX2_X1 U6890 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4500), .Z(n5317) );
  XNOR2_X1 U6891 ( .A(n5317), .B(n5310), .ZN(n5316) );
  XNOR2_X1 U6892 ( .A(n5320), .B(n5316), .ZN(n7051) );
  NAND2_X1 U6893 ( .A1(n7051), .A2(n5434), .ZN(n5315) );
  NAND2_X1 U6894 ( .A1(n5312), .A2(n5311), .ZN(n5313) );
  NAND2_X1 U6895 ( .A1(n5313), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5326) );
  XNOR2_X1 U6896 ( .A(n5326), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9587) );
  AOI22_X1 U6897 ( .A1(n5406), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5330), .B2(
        n9587), .ZN(n5314) );
  INV_X1 U6898 ( .A(n5316), .ZN(n5319) );
  NAND2_X1 U6899 ( .A1(n5317), .A2(SI_18_), .ZN(n5318) );
  NAND2_X1 U6900 ( .A1(n5322), .A2(n5321), .ZN(n5333) );
  INV_X1 U6901 ( .A(n5322), .ZN(n5323) );
  NAND2_X1 U6902 ( .A1(n5323), .A2(SI_19_), .ZN(n5324) );
  NAND2_X1 U6903 ( .A1(n5333), .A2(n5324), .ZN(n5334) );
  XNOR2_X1 U6904 ( .A(n5335), .B(n5334), .ZN(n7136) );
  NAND2_X1 U6905 ( .A1(n7136), .A2(n5434), .ZN(n5332) );
  NAND2_X1 U6906 ( .A1(n5326), .A2(n5325), .ZN(n5327) );
  XNOR2_X2 U6907 ( .A(n5329), .B(n5328), .ZN(n9720) );
  AOI22_X1 U6908 ( .A1(n5406), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5330), .B2(
        n9598), .ZN(n5331) );
  MUX2_X1 U6909 ( .A(n8894), .B(n7224), .S(n4499), .Z(n5339) );
  XNOR2_X1 U6910 ( .A(n5339), .B(SI_20_), .ZN(n5336) );
  XNOR2_X1 U6911 ( .A(n5340), .B(n5336), .ZN(n7223) );
  NAND2_X1 U6912 ( .A1(n7223), .A2(n5434), .ZN(n5338) );
  NAND2_X1 U6913 ( .A1(n5406), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5337) );
  INV_X1 U6914 ( .A(n9913), .ZN(n9734) );
  XNOR2_X1 U6915 ( .A(n5344), .B(SI_21_), .ZN(n5341) );
  XNOR2_X1 U6916 ( .A(n5347), .B(n5341), .ZN(n7367) );
  NAND2_X1 U6917 ( .A1(n7367), .A2(n5434), .ZN(n5343) );
  NAND2_X1 U6918 ( .A1(n5406), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5342) );
  NOR2_X1 U6919 ( .A1(n5345), .A2(SI_21_), .ZN(n5346) );
  MUX2_X1 U6920 ( .A(n9038), .B(n9041), .S(n4500), .Z(n5349) );
  INV_X1 U6921 ( .A(SI_22_), .ZN(n5348) );
  NAND2_X1 U6922 ( .A1(n5349), .A2(n5348), .ZN(n5354) );
  INV_X1 U6923 ( .A(n5349), .ZN(n5350) );
  NAND2_X1 U6924 ( .A1(n5350), .A2(SI_22_), .ZN(n5351) );
  NAND2_X1 U6925 ( .A1(n5354), .A2(n5351), .ZN(n5355) );
  XNOR2_X1 U6926 ( .A(n5356), .B(n5355), .ZN(n7492) );
  NAND2_X1 U6927 ( .A1(n7492), .A2(n5434), .ZN(n5353) );
  OR2_X1 U6928 ( .A1(n5173), .A2(n9041), .ZN(n5352) );
  INV_X1 U6929 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7573) );
  INV_X1 U6930 ( .A(SI_23_), .ZN(n5357) );
  NAND2_X1 U6931 ( .A1(n5358), .A2(n5357), .ZN(n5366) );
  INV_X1 U6932 ( .A(n5358), .ZN(n5359) );
  NAND2_X1 U6933 ( .A1(n5359), .A2(SI_23_), .ZN(n5360) );
  OR2_X1 U6934 ( .A1(n5362), .A2(n5361), .ZN(n5363) );
  NAND2_X1 U6935 ( .A1(n5367), .A2(n5363), .ZN(n7575) );
  NAND2_X1 U6936 ( .A1(n7575), .A2(n5434), .ZN(n5365) );
  OR2_X1 U6937 ( .A1(n5173), .A2(n8913), .ZN(n5364) );
  INV_X1 U6938 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7620) );
  MUX2_X1 U6939 ( .A(n7673), .B(n7620), .S(n4499), .Z(n5369) );
  INV_X1 U6940 ( .A(SI_24_), .ZN(n5368) );
  NAND2_X1 U6941 ( .A1(n5369), .A2(n5368), .ZN(n5376) );
  INV_X1 U6942 ( .A(n5369), .ZN(n5370) );
  NAND2_X1 U6943 ( .A1(n5370), .A2(SI_24_), .ZN(n5371) );
  XNOR2_X1 U6944 ( .A(n5375), .B(n5374), .ZN(n7619) );
  NAND2_X1 U6945 ( .A1(n7619), .A2(n5434), .ZN(n5373) );
  NAND2_X1 U6946 ( .A1(n5406), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5372) );
  INV_X1 U6947 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7746) );
  INV_X1 U6948 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7743) );
  MUX2_X1 U6949 ( .A(n7746), .B(n7743), .S(n4500), .Z(n5378) );
  INV_X1 U6950 ( .A(SI_25_), .ZN(n5377) );
  NAND2_X1 U6951 ( .A1(n5378), .A2(n5377), .ZN(n5385) );
  INV_X1 U6952 ( .A(n5378), .ZN(n5379) );
  NAND2_X1 U6953 ( .A1(n5379), .A2(SI_25_), .ZN(n5380) );
  XNOR2_X1 U6954 ( .A(n5384), .B(n5383), .ZN(n7742) );
  NAND2_X1 U6955 ( .A1(n7742), .A2(n5434), .ZN(n5382) );
  NAND2_X1 U6956 ( .A1(n5406), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5381) );
  NAND2_X1 U6957 ( .A1(n5384), .A2(n5383), .ZN(n5386) );
  NAND2_X1 U6958 ( .A1(n5386), .A2(n5385), .ZN(n5394) );
  INV_X1 U6959 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7777) );
  INV_X1 U6960 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7804) );
  NAND2_X1 U6961 ( .A1(n5388), .A2(n5387), .ZN(n5395) );
  INV_X1 U6962 ( .A(n5388), .ZN(n5389) );
  NAND2_X1 U6963 ( .A1(n5389), .A2(SI_26_), .ZN(n5390) );
  XNOR2_X1 U6964 ( .A(n5394), .B(n5393), .ZN(n7775) );
  NAND2_X1 U6965 ( .A1(n7775), .A2(n5434), .ZN(n5392) );
  NAND2_X1 U6966 ( .A1(n5406), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5391) );
  NAND2_X1 U6967 ( .A1(n5394), .A2(n5393), .ZN(n5396) );
  NAND2_X1 U6968 ( .A1(n5396), .A2(n5395), .ZN(n5404) );
  INV_X1 U6969 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9021) );
  INV_X1 U6970 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7803) );
  MUX2_X1 U6971 ( .A(n9021), .B(n7803), .S(n4500), .Z(n5398) );
  INV_X1 U6972 ( .A(SI_27_), .ZN(n5397) );
  NAND2_X1 U6973 ( .A1(n5398), .A2(n5397), .ZN(n5405) );
  INV_X1 U6974 ( .A(n5398), .ZN(n5399) );
  NAND2_X1 U6975 ( .A1(n5399), .A2(SI_27_), .ZN(n5400) );
  XNOR2_X1 U6976 ( .A(n5404), .B(n5403), .ZN(n7802) );
  NAND2_X1 U6977 ( .A1(n7802), .A2(n5434), .ZN(n5402) );
  NAND2_X1 U6978 ( .A1(n5406), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5401) );
  NAND2_X1 U6979 ( .A1(n9612), .A2(n9885), .ZN(n5765) );
  INV_X1 U6980 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7818) );
  XNOR2_X1 U6981 ( .A(n5412), .B(SI_28_), .ZN(n5409) );
  XNOR2_X1 U6982 ( .A(n5410), .B(n5409), .ZN(n7817) );
  NAND2_X1 U6983 ( .A1(n7817), .A2(n5434), .ZN(n5408) );
  NAND2_X1 U6984 ( .A1(n5406), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5407) );
  INV_X1 U6985 ( .A(SI_28_), .ZN(n5411) );
  NAND2_X1 U6986 ( .A1(n5412), .A2(n5411), .ZN(n5413) );
  INV_X1 U6987 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8552) );
  MUX2_X1 U6988 ( .A(n7801), .B(n8552), .S(n4835), .Z(n5416) );
  XNOR2_X1 U6989 ( .A(n5419), .B(SI_29_), .ZN(n7799) );
  NAND2_X1 U6990 ( .A1(n7799), .A2(n5434), .ZN(n5415) );
  OR2_X1 U6991 ( .A1(n5173), .A2(n7801), .ZN(n5414) );
  OR2_X1 U6992 ( .A1(n5417), .A2(n5416), .ZN(n5418) );
  INV_X1 U6993 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7882) );
  MUX2_X1 U6994 ( .A(n7882), .B(n7886), .S(n4835), .Z(n5421) );
  INV_X1 U6995 ( .A(SI_30_), .ZN(n5420) );
  NAND2_X1 U6996 ( .A1(n5421), .A2(n5420), .ZN(n5429) );
  INV_X1 U6997 ( .A(n5421), .ZN(n5422) );
  NAND2_X1 U6998 ( .A1(n5422), .A2(SI_30_), .ZN(n5423) );
  NAND2_X1 U6999 ( .A1(n5429), .A2(n5423), .ZN(n5424) );
  NAND2_X1 U7000 ( .A1(n5425), .A2(n5424), .ZN(n5426) );
  NAND2_X1 U7001 ( .A1(n5430), .A2(n5426), .ZN(n7885) );
  NAND2_X1 U7002 ( .A1(n7885), .A2(n5434), .ZN(n5428) );
  OR2_X1 U7003 ( .A1(n5173), .A2(n7882), .ZN(n5427) );
  NAND2_X1 U7004 ( .A1(n5430), .A2(n5429), .ZN(n5433) );
  INV_X1 U7005 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5435) );
  INV_X1 U7006 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n7892) );
  MUX2_X1 U7007 ( .A(n5435), .B(n7892), .S(n4835), .Z(n5431) );
  XNOR2_X1 U7008 ( .A(n5431), .B(SI_31_), .ZN(n5432) );
  XNOR2_X1 U7009 ( .A(n5433), .B(n5432), .ZN(n8546) );
  NAND2_X1 U7010 ( .A1(n8546), .A2(n5434), .ZN(n5437) );
  OR2_X1 U7011 ( .A1(n5173), .A2(n5435), .ZN(n5436) );
  INV_X1 U7012 ( .A(n5440), .ZN(n5441) );
  NAND2_X1 U7013 ( .A1(n5442), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5443) );
  NAND2_X1 U7014 ( .A1(n5447), .A2(n5446), .ZN(n5448) );
  NAND2_X1 U7015 ( .A1(n4494), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5453) );
  INV_X1 U7016 ( .A(n7884), .ZN(n5495) );
  NAND2_X1 U7017 ( .A1(n5079), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5452) );
  NAND2_X1 U7018 ( .A1(n7785), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5451) );
  AND3_X1 U7019 ( .A1(n5453), .A2(n5452), .A3(n5451), .ZN(n9452) );
  NAND2_X1 U7020 ( .A1(n5726), .A2(n9365), .ZN(n6538) );
  INV_X1 U7021 ( .A(n5456), .ZN(n9987) );
  NAND2_X1 U7022 ( .A1(n9987), .A2(P1_B_REG_SCAN_IN), .ZN(n5457) );
  NAND2_X1 U7023 ( .A1(n9184), .A2(n5457), .ZN(n7789) );
  NOR2_X1 U7024 ( .A1(n9452), .A2(n7789), .ZN(n9603) );
  NOR2_X1 U7025 ( .A1(n9602), .A2(n9603), .ZN(n6385) );
  NAND2_X1 U7026 ( .A1(n5460), .A2(n5459), .ZN(n5462) );
  OR2_X1 U7027 ( .A1(n5460), .A2(n5459), .ZN(n5461) );
  NAND2_X1 U7028 ( .A1(n7744), .A2(P1_B_REG_SCAN_IN), .ZN(n5465) );
  MUX2_X1 U7029 ( .A(n5465), .B(P1_B_REG_SCAN_IN), .S(n5467), .Z(n5466) );
  OAI22_X1 U7030 ( .A1(n5475), .A2(P1_D_REG_0__SCAN_IN), .B1(n5468), .B2(n5467), .ZN(n6537) );
  INV_X1 U7031 ( .A(n6537), .ZN(n5474) );
  NAND2_X1 U7032 ( .A1(n5470), .A2(n5469), .ZN(n5471) );
  NAND2_X1 U7033 ( .A1(n5471), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5473) );
  INV_X4 U7034 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  AND2_X1 U7035 ( .A1(n5474), .A2(n9475), .ZN(n6465) );
  INV_X1 U7036 ( .A(n5468), .ZN(n7806) );
  NAND2_X1 U7037 ( .A1(n7806), .A2(n7744), .ZN(n6851) );
  OAI21_X1 U7038 ( .B1(n5475), .B2(P1_D_REG_1__SCAN_IN), .A(n6851), .ZN(n6534)
         );
  NOR4_X1 U7039 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5484) );
  NOR4_X1 U7040 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n5483) );
  INV_X1 U7041 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10078) );
  INV_X1 U7042 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n10094) );
  INV_X1 U7043 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10077) );
  INV_X1 U7044 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10089) );
  NAND4_X1 U7045 ( .A1(n10078), .A2(n10094), .A3(n10077), .A4(n10089), .ZN(
        n5481) );
  NOR4_X1 U7046 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n5479) );
  NOR4_X1 U7047 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n5478) );
  NOR4_X1 U7048 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5477) );
  NOR4_X1 U7049 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n5476) );
  NAND4_X1 U7050 ( .A1(n5479), .A2(n5478), .A3(n5477), .A4(n5476), .ZN(n5480)
         );
  NOR4_X1 U7051 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n5481), .A4(n5480), .ZN(n5482) );
  NAND3_X1 U7052 ( .A1(n5484), .A2(n5483), .A3(n5482), .ZN(n5485) );
  NAND2_X1 U7053 ( .A1(n6849), .A2(n5485), .ZN(n6535) );
  INV_X1 U7054 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n5486) );
  NOR2_X1 U7055 ( .A1(n10192), .A2(n5486), .ZN(n5487) );
  NOR2_X1 U7056 ( .A1(n5488), .A2(n5487), .ZN(n5489) );
  OAI21_X1 U7057 ( .B1(n6385), .B2(n5490), .A(n5489), .ZN(P1_U3553) );
  NAND2_X1 U7058 ( .A1(n5079), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5499) );
  NAND2_X1 U7059 ( .A1(n5527), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5497) );
  NAND2_X1 U7060 ( .A1(n5503), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U7061 ( .A1(n4494), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6493) );
  NAND2_X1 U7062 ( .A1(n5503), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6492) );
  NAND2_X1 U7063 ( .A1(n5079), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6491) );
  NAND2_X1 U7064 ( .A1(n5518), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6490) );
  NAND4_X1 U7065 ( .A1(n6493), .A2(n6492), .A3(n6491), .A4(n6490), .ZN(n6533)
         );
  NAND2_X1 U7066 ( .A1(n6533), .A2(n7172), .ZN(n7280) );
  INV_X1 U7067 ( .A(n6633), .ZN(n5729) );
  NAND2_X1 U7068 ( .A1(n5729), .A2(n10104), .ZN(n5501) );
  NAND2_X1 U7069 ( .A1(n5079), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U7070 ( .A1(n5518), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5504) );
  NAND3_X1 U7071 ( .A1(n5506), .A2(n5505), .A3(n5504), .ZN(n9517) );
  NAND2_X1 U7072 ( .A1(n6930), .A2(n6763), .ZN(n5732) );
  NAND2_X1 U7073 ( .A1(n7266), .A2(n7262), .ZN(n5509) );
  NAND2_X1 U7074 ( .A1(n6930), .A2(n5507), .ZN(n5508) );
  NAND2_X1 U7075 ( .A1(n5509), .A2(n5508), .ZN(n10061) );
  NAND2_X1 U7076 ( .A1(n4494), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5514) );
  INV_X1 U7077 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U7078 ( .A1(n5518), .A2(n5510), .ZN(n5513) );
  NAND2_X1 U7079 ( .A1(n5079), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5512) );
  NAND2_X1 U7080 ( .A1(n5503), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5511) );
  NAND2_X1 U7081 ( .A1(n9516), .A2(n10118), .ZN(n9386) );
  NAND2_X1 U7082 ( .A1(n6919), .A2(n5515), .ZN(n9389) );
  NAND2_X1 U7083 ( .A1(n9386), .A2(n9389), .ZN(n10062) );
  NAND2_X1 U7084 ( .A1(n10061), .A2(n10062), .ZN(n5517) );
  NAND2_X1 U7085 ( .A1(n6919), .A2(n10118), .ZN(n5516) );
  NAND2_X1 U7086 ( .A1(n5517), .A2(n5516), .ZN(n7310) );
  NAND2_X1 U7087 ( .A1(n4494), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5523) );
  NAND2_X1 U7088 ( .A1(n5079), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5522) );
  AND2_X1 U7089 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5528) );
  NOR2_X1 U7090 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5519) );
  NOR2_X1 U7091 ( .A1(n5528), .A2(n5519), .ZN(n7313) );
  NAND2_X1 U7092 ( .A1(n5518), .A2(n7313), .ZN(n5521) );
  NAND2_X1 U7093 ( .A1(n5503), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U7094 ( .A1(n5524), .A2(n7314), .ZN(n9393) );
  INV_X1 U7095 ( .A(n5524), .ZN(n9515) );
  NAND2_X1 U7096 ( .A1(n7310), .A2(n9334), .ZN(n5526) );
  NAND2_X1 U7097 ( .A1(n5524), .A2(n10125), .ZN(n5525) );
  NAND2_X1 U7098 ( .A1(n5526), .A2(n5525), .ZN(n7288) );
  NAND2_X1 U7099 ( .A1(n4494), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5533) );
  NAND2_X1 U7100 ( .A1(n7785), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5532) );
  NAND2_X1 U7101 ( .A1(n5528), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5537) );
  OAI21_X1 U7102 ( .B1(n5528), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5537), .ZN(
        n5529) );
  INV_X1 U7103 ( .A(n5529), .ZN(n7297) );
  NAND2_X1 U7104 ( .A1(n5518), .A2(n7297), .ZN(n5531) );
  NAND2_X1 U7105 ( .A1(n5672), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5530) );
  NAND2_X1 U7106 ( .A1(n7326), .A2(n7298), .ZN(n9394) );
  INV_X1 U7107 ( .A(n7326), .ZN(n9514) );
  INV_X1 U7108 ( .A(n7298), .ZN(n10132) );
  NAND2_X1 U7109 ( .A1(n9514), .A2(n10132), .ZN(n9397) );
  NAND2_X1 U7110 ( .A1(n7288), .A2(n9335), .ZN(n5535) );
  NAND2_X1 U7111 ( .A1(n7326), .A2(n10132), .ZN(n5534) );
  NAND2_X1 U7112 ( .A1(n5535), .A2(n5534), .ZN(n7355) );
  NAND2_X1 U7113 ( .A1(n7785), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5542) );
  NAND2_X1 U7114 ( .A1(n4494), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5541) );
  INV_X1 U7115 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5536) );
  NOR2_X1 U7116 ( .A1(n5537), .A2(n5536), .ZN(n5545) );
  AND2_X1 U7117 ( .A1(n5537), .A2(n5536), .ZN(n5538) );
  NOR2_X1 U7118 ( .A1(n5545), .A2(n5538), .ZN(n7360) );
  NAND2_X1 U7119 ( .A1(n5518), .A2(n7360), .ZN(n5540) );
  NAND2_X1 U7120 ( .A1(n5672), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5539) );
  NAND2_X1 U7121 ( .A1(n7246), .A2(n7361), .ZN(n10034) );
  INV_X1 U7122 ( .A(n7246), .ZN(n9513) );
  NAND2_X1 U7123 ( .A1(n9513), .A2(n10138), .ZN(n9223) );
  NAND2_X1 U7124 ( .A1(n7355), .A2(n7356), .ZN(n5544) );
  NAND2_X1 U7125 ( .A1(n7246), .A2(n10138), .ZN(n5543) );
  NAND2_X1 U7126 ( .A1(n5544), .A2(n5543), .ZN(n10032) );
  NAND2_X1 U7127 ( .A1(n7785), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5550) );
  NAND2_X1 U7128 ( .A1(n4494), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5549) );
  NAND2_X1 U7129 ( .A1(n5545), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5552) );
  OR2_X1 U7130 ( .A1(n5545), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5546) );
  AND2_X1 U7131 ( .A1(n5552), .A2(n5546), .ZN(n10041) );
  NAND2_X1 U7132 ( .A1(n5518), .A2(n10041), .ZN(n5548) );
  NAND2_X1 U7133 ( .A1(n5672), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5547) );
  NAND2_X1 U7134 ( .A1(n7339), .A2(n10044), .ZN(n7337) );
  INV_X1 U7135 ( .A(n7339), .ZN(n9512) );
  NAND2_X1 U7136 ( .A1(n9512), .A2(n10145), .ZN(n5738) );
  NAND2_X1 U7137 ( .A1(n7337), .A2(n5738), .ZN(n10033) );
  NAND2_X1 U7138 ( .A1(n7339), .A2(n10145), .ZN(n5551) );
  NAND2_X1 U7139 ( .A1(n4494), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5557) );
  NAND2_X1 U7140 ( .A1(n5672), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5556) );
  NAND2_X1 U7141 ( .A1(n5552), .A2(n7521), .ZN(n5553) );
  AND2_X1 U7142 ( .A1(n5559), .A2(n5553), .ZN(n7524) );
  NAND2_X1 U7143 ( .A1(n5518), .A2(n7524), .ZN(n5555) );
  NAND2_X1 U7144 ( .A1(n7785), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5554) );
  NAND2_X1 U7145 ( .A1(n7516), .A2(n7510), .ZN(n9236) );
  INV_X1 U7146 ( .A(n7516), .ZN(n9511) );
  NAND2_X1 U7147 ( .A1(n9511), .A2(n5006), .ZN(n5739) );
  NAND2_X1 U7148 ( .A1(n4494), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U7149 ( .A1(n7785), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5563) );
  INV_X1 U7150 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5558) );
  NOR2_X1 U7151 ( .A1(n5559), .A2(n5558), .ZN(n5567) );
  AND2_X1 U7152 ( .A1(n5559), .A2(n5558), .ZN(n5560) );
  NOR2_X1 U7153 ( .A1(n5567), .A2(n5560), .ZN(n7600) );
  NAND2_X1 U7154 ( .A1(n5518), .A2(n7600), .ZN(n5562) );
  NAND2_X1 U7155 ( .A1(n5672), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U7156 ( .A1(n7597), .A2(n7605), .ZN(n9243) );
  INV_X1 U7157 ( .A(n7597), .ZN(n9510) );
  NAND2_X1 U7158 ( .A1(n9510), .A2(n10161), .ZN(n9246) );
  NAND2_X1 U7159 ( .A1(n9243), .A2(n9246), .ZN(n7404) );
  NAND2_X1 U7160 ( .A1(n7403), .A2(n7404), .ZN(n5566) );
  NAND2_X1 U7161 ( .A1(n7597), .A2(n10161), .ZN(n5565) );
  NAND2_X1 U7162 ( .A1(n5566), .A2(n5565), .ZN(n7396) );
  NAND2_X1 U7163 ( .A1(n7785), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U7164 ( .A1(n4494), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5572) );
  NOR2_X1 U7165 ( .A1(n5567), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5568) );
  OR2_X1 U7166 ( .A1(n5576), .A2(n5568), .ZN(n8706) );
  INV_X1 U7167 ( .A(n8706), .ZN(n5569) );
  NAND2_X1 U7168 ( .A1(n5518), .A2(n5569), .ZN(n5571) );
  NAND2_X1 U7169 ( .A1(n5672), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U7170 ( .A1(n7638), .A2(n8713), .ZN(n9402) );
  INV_X1 U7171 ( .A(n7638), .ZN(n9509) );
  NAND2_X1 U7172 ( .A1(n9509), .A2(n10169), .ZN(n9399) );
  NAND2_X1 U7173 ( .A1(n7396), .A2(n9342), .ZN(n5575) );
  NAND2_X1 U7174 ( .A1(n7638), .A2(n10169), .ZN(n5574) );
  NAND2_X1 U7175 ( .A1(n5575), .A2(n5574), .ZN(n7435) );
  NAND2_X1 U7176 ( .A1(n5576), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5585) );
  OR2_X1 U7177 ( .A1(n5576), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5577) );
  AND2_X1 U7178 ( .A1(n5585), .A2(n5577), .ZN(n7691) );
  NAND2_X1 U7179 ( .A1(n5518), .A2(n7691), .ZN(n5581) );
  NAND2_X1 U7180 ( .A1(n4494), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5580) );
  NAND2_X1 U7181 ( .A1(n5672), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5579) );
  NAND2_X1 U7182 ( .A1(n7785), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5578) );
  NAND4_X1 U7183 ( .A1(n5581), .A2(n5580), .A3(n5579), .A4(n5578), .ZN(n9508)
         );
  NOR2_X1 U7184 ( .A1(n7693), .A2(n9508), .ZN(n5583) );
  NAND2_X1 U7185 ( .A1(n7693), .A2(n9508), .ZN(n5582) );
  NAND2_X1 U7186 ( .A1(n4494), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5590) );
  NAND2_X1 U7187 ( .A1(n7785), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5589) );
  NAND2_X1 U7188 ( .A1(n5079), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U7189 ( .A1(n5585), .A2(n5584), .ZN(n5586) );
  NAND2_X1 U7190 ( .A1(n5594), .A2(n5586), .ZN(n9969) );
  INV_X1 U7191 ( .A(n9969), .ZN(n7504) );
  NAND2_X1 U7192 ( .A1(n5518), .A2(n7504), .ZN(n5587) );
  OR2_X1 U7193 ( .A1(n7653), .A2(n7655), .ZN(n9255) );
  NAND2_X1 U7194 ( .A1(n7653), .A2(n7655), .ZN(n9257) );
  NAND2_X1 U7195 ( .A1(n9255), .A2(n9257), .ZN(n7497) );
  NAND2_X1 U7196 ( .A1(n7495), .A2(n7497), .ZN(n5592) );
  INV_X1 U7197 ( .A(n7655), .ZN(n9507) );
  NAND2_X1 U7198 ( .A1(n7653), .A2(n9507), .ZN(n5591) );
  NAND2_X1 U7199 ( .A1(n5592), .A2(n5591), .ZN(n7586) );
  NAND2_X1 U7200 ( .A1(n5527), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U7201 ( .A1(n7785), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U7202 ( .A1(n5594), .A2(n5593), .ZN(n5595) );
  AND2_X1 U7203 ( .A1(n5601), .A2(n5595), .ZN(n7669) );
  NAND2_X1 U7204 ( .A1(n5518), .A2(n7669), .ZN(n5597) );
  NAND2_X1 U7205 ( .A1(n5672), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5596) );
  OR2_X1 U7206 ( .A1(n7625), .A2(n7708), .ZN(n9409) );
  NAND2_X1 U7207 ( .A1(n7625), .A2(n7708), .ZN(n9258) );
  INV_X1 U7208 ( .A(n7708), .ZN(n9506) );
  NAND2_X1 U7209 ( .A1(n7625), .A2(n9506), .ZN(n5600) );
  NAND2_X1 U7210 ( .A1(n7785), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U7211 ( .A1(n4494), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5605) );
  AND2_X1 U7212 ( .A1(n5601), .A2(n8683), .ZN(n5602) );
  NOR2_X1 U7213 ( .A1(n5609), .A2(n5602), .ZN(n8687) );
  NAND2_X1 U7214 ( .A1(n5518), .A2(n8687), .ZN(n5604) );
  NAND2_X1 U7215 ( .A1(n5672), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5603) );
  NAND4_X1 U7216 ( .A1(n5606), .A2(n5605), .A3(n5604), .A4(n5603), .ZN(n9505)
         );
  AND2_X1 U7217 ( .A1(n9263), .A2(n9505), .ZN(n5608) );
  OR2_X1 U7218 ( .A1(n9263), .A2(n9505), .ZN(n5607) );
  NAND2_X1 U7219 ( .A1(n5527), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5614) );
  NAND2_X1 U7220 ( .A1(n5672), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5613) );
  OR2_X1 U7221 ( .A1(n5609), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5610) );
  NAND2_X1 U7222 ( .A1(n5609), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5615) );
  AND2_X1 U7223 ( .A1(n5610), .A2(n5615), .ZN(n9210) );
  NAND2_X1 U7224 ( .A1(n5518), .A2(n9210), .ZN(n5612) );
  NAND2_X1 U7225 ( .A1(n7785), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5611) );
  NAND4_X1 U7226 ( .A1(n5614), .A2(n5613), .A3(n5612), .A4(n5611), .ZN(n9503)
         );
  NOR2_X1 U7227 ( .A1(n9218), .A2(n9503), .ZN(n7719) );
  NAND2_X1 U7228 ( .A1(n4494), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5620) );
  NAND2_X1 U7229 ( .A1(n7785), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5619) );
  NAND2_X1 U7230 ( .A1(n5615), .A2(n8773), .ZN(n5616) );
  AND2_X1 U7231 ( .A1(n5624), .A2(n5616), .ZN(n9797) );
  NAND2_X1 U7232 ( .A1(n5518), .A2(n9797), .ZN(n5618) );
  NAND2_X1 U7233 ( .A1(n5672), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5617) );
  OR2_X1 U7234 ( .A1(n9796), .A2(n9142), .ZN(n9416) );
  NAND2_X1 U7235 ( .A1(n9796), .A2(n9142), .ZN(n9418) );
  NAND2_X1 U7236 ( .A1(n9416), .A2(n9418), .ZN(n9788) );
  NAND2_X1 U7237 ( .A1(n9785), .A2(n9788), .ZN(n5622) );
  INV_X1 U7238 ( .A(n9142), .ZN(n9502) );
  NAND2_X1 U7239 ( .A1(n9796), .A2(n9502), .ZN(n5621) );
  NAND2_X1 U7240 ( .A1(n4494), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5629) );
  NAND2_X1 U7241 ( .A1(n7785), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5628) );
  INV_X1 U7242 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5623) );
  AND2_X1 U7243 ( .A1(n5624), .A2(n5623), .ZN(n5625) );
  NOR2_X1 U7244 ( .A1(n5631), .A2(n5625), .ZN(n9779) );
  NAND2_X1 U7245 ( .A1(n5518), .A2(n9779), .ZN(n5627) );
  NAND2_X1 U7246 ( .A1(n5672), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5626) );
  NAND4_X1 U7247 ( .A1(n5629), .A2(n5628), .A3(n5627), .A4(n5626), .ZN(n9501)
         );
  OR2_X1 U7248 ( .A1(n9333), .A2(n9501), .ZN(n5630) );
  NAND2_X1 U7249 ( .A1(n7785), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5636) );
  NAND2_X1 U7250 ( .A1(n4494), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5635) );
  NOR2_X1 U7251 ( .A1(n5631), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5632) );
  OR2_X1 U7252 ( .A1(n5637), .A2(n5632), .ZN(n9188) );
  INV_X1 U7253 ( .A(n9188), .ZN(n9766) );
  NAND2_X1 U7254 ( .A1(n5518), .A2(n9766), .ZN(n5634) );
  NAND2_X1 U7255 ( .A1(n5672), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5633) );
  NAND4_X1 U7256 ( .A1(n5636), .A2(n5635), .A3(n5634), .A4(n5633), .ZN(n9500)
         );
  NAND2_X1 U7257 ( .A1(n4494), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5642) );
  NAND2_X1 U7258 ( .A1(n7785), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5641) );
  NOR2_X1 U7259 ( .A1(n5637), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5638) );
  OR2_X1 U7260 ( .A1(n5644), .A2(n5638), .ZN(n8723) );
  INV_X1 U7261 ( .A(n8723), .ZN(n9749) );
  NAND2_X1 U7262 ( .A1(n5518), .A2(n9749), .ZN(n5640) );
  NAND2_X1 U7263 ( .A1(n5672), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5639) );
  NAND4_X1 U7264 ( .A1(n5642), .A2(n5641), .A3(n5640), .A4(n5639), .ZN(n9499)
         );
  OR2_X1 U7265 ( .A1(n9748), .A2(n9499), .ZN(n5643) );
  NAND2_X1 U7266 ( .A1(n4494), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5649) );
  NAND2_X1 U7267 ( .A1(n7785), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5648) );
  NOR2_X1 U7268 ( .A1(n5644), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5645) );
  NOR2_X1 U7269 ( .A1(n5652), .A2(n5645), .ZN(n9735) );
  NAND2_X1 U7270 ( .A1(n5518), .A2(n9735), .ZN(n5647) );
  NAND2_X1 U7271 ( .A1(n5672), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5646) );
  NAND4_X1 U7272 ( .A1(n5649), .A2(n5648), .A3(n5647), .A4(n5646), .ZN(n9498)
         );
  NAND2_X1 U7273 ( .A1(n9913), .A2(n9498), .ZN(n9288) );
  INV_X1 U7274 ( .A(n9498), .ZN(n8720) );
  NAND2_X1 U7275 ( .A1(n9734), .A2(n8720), .ZN(n9286) );
  NAND2_X1 U7276 ( .A1(n9913), .A2(n8720), .ZN(n5651) );
  NAND2_X1 U7277 ( .A1(n9726), .A2(n5651), .ZN(n9710) );
  NAND2_X1 U7278 ( .A1(n7785), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5657) );
  NAND2_X1 U7279 ( .A1(n4494), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5656) );
  OR2_X1 U7280 ( .A1(n5652), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5653) );
  NAND2_X1 U7281 ( .A1(n5652), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5662) );
  AND2_X1 U7282 ( .A1(n5653), .A2(n5662), .ZN(n9721) );
  NAND2_X1 U7283 ( .A1(n5518), .A2(n9721), .ZN(n5655) );
  NAND2_X1 U7284 ( .A1(n5672), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5654) );
  NAND4_X1 U7285 ( .A1(n5657), .A2(n5656), .A3(n5655), .A4(n5654), .ZN(n9497)
         );
  NAND2_X1 U7286 ( .A1(n9715), .A2(n9497), .ZN(n5658) );
  NAND2_X1 U7287 ( .A1(n9710), .A2(n5658), .ZN(n5660) );
  OR2_X1 U7288 ( .A1(n9715), .A2(n9497), .ZN(n5659) );
  NAND2_X1 U7289 ( .A1(n5660), .A2(n5659), .ZN(n9694) );
  NAND2_X1 U7290 ( .A1(n4494), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5668) );
  NAND2_X1 U7291 ( .A1(n7785), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5667) );
  INV_X1 U7292 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U7293 ( .A1(n5661), .A2(n5662), .ZN(n5664) );
  INV_X1 U7294 ( .A(n5662), .ZN(n5663) );
  NAND2_X1 U7295 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(n5663), .ZN(n5670) );
  AND2_X1 U7296 ( .A1(n5664), .A2(n5670), .ZN(n9704) );
  NAND2_X1 U7297 ( .A1(n5518), .A2(n9704), .ZN(n5666) );
  NAND2_X1 U7298 ( .A1(n5672), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5665) );
  NAND4_X1 U7299 ( .A1(n5668), .A2(n5667), .A3(n5666), .A4(n5665), .ZN(n9496)
         );
  NAND2_X1 U7300 ( .A1(n7785), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5676) );
  NAND2_X1 U7301 ( .A1(n5527), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5675) );
  INV_X1 U7302 ( .A(n5670), .ZN(n5669) );
  NAND2_X1 U7303 ( .A1(n5669), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5679) );
  INV_X1 U7304 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8700) );
  NAND2_X1 U7305 ( .A1(n5670), .A2(n8700), .ZN(n5671) );
  AND2_X1 U7306 ( .A1(n5679), .A2(n5671), .ZN(n9681) );
  NAND2_X1 U7307 ( .A1(n5518), .A2(n9681), .ZN(n5674) );
  NAND2_X1 U7308 ( .A1(n5672), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5673) );
  OR2_X1 U7309 ( .A1(n9690), .A2(n9171), .ZN(n9297) );
  INV_X1 U7310 ( .A(n9664), .ZN(n5685) );
  NAND2_X1 U7311 ( .A1(n7785), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5684) );
  NAND2_X1 U7312 ( .A1(n4494), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5683) );
  INV_X1 U7313 ( .A(n5679), .ZN(n5678) );
  NAND2_X1 U7314 ( .A1(n5678), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5688) );
  INV_X1 U7315 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9155) );
  NAND2_X1 U7316 ( .A1(n5679), .A2(n9155), .ZN(n5680) );
  AND2_X1 U7317 ( .A1(n5688), .A2(n5680), .ZN(n9672) );
  NAND2_X1 U7318 ( .A1(n5518), .A2(n9672), .ZN(n5682) );
  NAND2_X1 U7319 ( .A1(n5672), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5681) );
  NAND4_X1 U7320 ( .A1(n5684), .A2(n5683), .A3(n5682), .A4(n5681), .ZN(n9494)
         );
  NAND2_X1 U7321 ( .A1(n9671), .A2(n9494), .ZN(n5686) );
  NAND2_X1 U7322 ( .A1(n7785), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5693) );
  NAND2_X1 U7323 ( .A1(n4494), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5692) );
  INV_X1 U7324 ( .A(n5688), .ZN(n5687) );
  NAND2_X1 U7325 ( .A1(n5687), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5698) );
  INV_X1 U7326 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8766) );
  NAND2_X1 U7327 ( .A1(n5688), .A2(n8766), .ZN(n5689) );
  AND2_X1 U7328 ( .A1(n5698), .A2(n5689), .ZN(n9657) );
  NAND2_X1 U7329 ( .A1(n5518), .A2(n9657), .ZN(n5691) );
  NAND2_X1 U7330 ( .A1(n5079), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5690) );
  NAND4_X1 U7331 ( .A1(n5693), .A2(n5692), .A3(n5691), .A4(n5690), .ZN(n9493)
         );
  OR2_X1 U7332 ( .A1(n9656), .A2(n9493), .ZN(n5694) );
  NAND2_X1 U7333 ( .A1(n5527), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5703) );
  NAND2_X1 U7334 ( .A1(n7785), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5702) );
  INV_X1 U7335 ( .A(n5698), .ZN(n5696) );
  NAND2_X1 U7336 ( .A1(n5696), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5707) );
  INV_X1 U7337 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5697) );
  NAND2_X1 U7338 ( .A1(n5698), .A2(n5697), .ZN(n5699) );
  AND2_X1 U7339 ( .A1(n5707), .A2(n5699), .ZN(n9640) );
  NAND2_X1 U7340 ( .A1(n5518), .A2(n9640), .ZN(n5701) );
  NAND2_X1 U7341 ( .A1(n5079), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5700) );
  NAND4_X1 U7342 ( .A1(n5703), .A2(n5702), .A3(n5701), .A4(n5700), .ZN(n9492)
         );
  NOR2_X1 U7343 ( .A1(n9639), .A2(n9492), .ZN(n5704) );
  INV_X1 U7344 ( .A(n9492), .ZN(n8673) );
  NAND2_X1 U7345 ( .A1(n5527), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5712) );
  NAND2_X1 U7346 ( .A1(n7785), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5711) );
  INV_X1 U7347 ( .A(n5707), .ZN(n5705) );
  NAND2_X1 U7348 ( .A1(n5705), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5716) );
  INV_X1 U7349 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5706) );
  NAND2_X1 U7350 ( .A1(n5707), .A2(n5706), .ZN(n5708) );
  AND2_X1 U7351 ( .A1(n5716), .A2(n5708), .ZN(n8672) );
  NAND2_X1 U7352 ( .A1(n5518), .A2(n8672), .ZN(n5710) );
  NAND2_X1 U7353 ( .A1(n5079), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5709) );
  OR2_X1 U7354 ( .A1(n9628), .A2(n9196), .ZN(n9313) );
  NAND2_X1 U7355 ( .A1(n9628), .A2(n9196), .ZN(n9310) );
  OR2_X1 U7356 ( .A1(n9628), .A2(n9491), .ZN(n5713) );
  INV_X1 U7357 ( .A(n5724), .ZN(n5723) );
  NAND2_X1 U7358 ( .A1(n4494), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5721) );
  NAND2_X1 U7359 ( .A1(n7785), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5720) );
  INV_X1 U7360 ( .A(n5716), .ZN(n5714) );
  NAND2_X1 U7361 ( .A1(n5714), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n5757) );
  INV_X1 U7362 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5715) );
  NAND2_X1 U7363 ( .A1(n5716), .A2(n5715), .ZN(n5717) );
  NAND2_X1 U7364 ( .A1(n5518), .A2(n8740), .ZN(n5719) );
  NAND2_X1 U7365 ( .A1(n5079), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5718) );
  OR2_X1 U7366 ( .A1(n8745), .A2(n8736), .ZN(n9368) );
  NAND2_X1 U7367 ( .A1(n8745), .A2(n8736), .ZN(n9318) );
  NAND2_X1 U7368 ( .A1(n9368), .A2(n9318), .ZN(n9360) );
  INV_X1 U7369 ( .A(n9360), .ZN(n5722) );
  NAND2_X1 U7370 ( .A1(n5723), .A2(n9360), .ZN(n7778) );
  NAND2_X1 U7371 ( .A1(n5724), .A2(n5722), .ZN(n5725) );
  NAND2_X1 U7372 ( .A1(n9365), .A2(n9720), .ZN(n6528) );
  NAND2_X1 U7373 ( .A1(n5726), .A2(n7225), .ZN(n6527) );
  OR2_X1 U7374 ( .A1(n6528), .A2(n6527), .ZN(n9473) );
  INV_X1 U7375 ( .A(n6545), .ZN(n9469) );
  NAND2_X1 U7376 ( .A1(n6528), .A2(n9469), .ZN(n5727) );
  NAND3_X1 U7377 ( .A1(n9473), .A2(n7164), .A3(n5727), .ZN(n10031) );
  INV_X2 U7378 ( .A(n9321), .ZN(n9325) );
  OR2_X1 U7379 ( .A1(n9325), .A2(n9467), .ZN(n10143) );
  NOR2_X1 U7380 ( .A1(n6533), .A2(n7275), .ZN(n7271) );
  NAND2_X1 U7381 ( .A1(n9337), .A2(n7271), .ZN(n5731) );
  NAND2_X1 U7382 ( .A1(n5729), .A2(n7279), .ZN(n5730) );
  INV_X1 U7383 ( .A(n5732), .ZN(n7305) );
  INV_X1 U7384 ( .A(n9389), .ZN(n5733) );
  INV_X1 U7385 ( .A(n9386), .ZN(n5735) );
  INV_X1 U7386 ( .A(n9391), .ZN(n5734) );
  INV_X1 U7387 ( .A(n9232), .ZN(n5737) );
  NAND2_X1 U7388 ( .A1(n5737), .A2(n9393), .ZN(n7289) );
  INV_X1 U7389 ( .A(n9335), .ZN(n7291) );
  NAND2_X1 U7390 ( .A1(n7289), .A2(n7291), .ZN(n7290) );
  NAND2_X1 U7391 ( .A1(n7337), .A2(n9236), .ZN(n9233) );
  AND2_X1 U7392 ( .A1(n5739), .A2(n5738), .ZN(n9235) );
  NAND3_X1 U7393 ( .A1(n9235), .A2(n9223), .A3(n9246), .ZN(n9341) );
  NAND2_X1 U7394 ( .A1(n4552), .A2(n9341), .ZN(n9400) );
  INV_X1 U7395 ( .A(n9342), .ZN(n7387) );
  AND2_X1 U7396 ( .A1(n9400), .A2(n7387), .ZN(n5740) );
  INV_X1 U7397 ( .A(n9508), .ZN(n7644) );
  OR2_X1 U7398 ( .A1(n7644), .A2(n7693), .ZN(n9254) );
  NAND2_X1 U7399 ( .A1(n7644), .A2(n7693), .ZN(n9401) );
  NAND2_X1 U7400 ( .A1(n9254), .A2(n9401), .ZN(n7436) );
  INV_X1 U7401 ( .A(n9254), .ZN(n5742) );
  NOR2_X1 U7402 ( .A1(n7497), .A2(n5742), .ZN(n5743) );
  NAND2_X1 U7403 ( .A1(n7496), .A2(n5743), .ZN(n5744) );
  NAND2_X1 U7404 ( .A1(n5744), .A2(n9257), .ZN(n7587) );
  XNOR2_X1 U7405 ( .A(n9263), .B(n9505), .ZN(n9349) );
  INV_X1 U7406 ( .A(n9503), .ZN(n8579) );
  NAND2_X1 U7407 ( .A1(n9218), .A2(n8579), .ZN(n9265) );
  INV_X1 U7408 ( .A(n9505), .ZN(n9262) );
  NAND2_X1 U7409 ( .A1(n9263), .A2(n9262), .ZN(n7718) );
  AND2_X1 U7410 ( .A1(n9265), .A2(n7718), .ZN(n9414) );
  OR2_X1 U7411 ( .A1(n9218), .A2(n8579), .ZN(n9787) );
  NAND2_X1 U7412 ( .A1(n9789), .A2(n9787), .ZN(n5747) );
  INV_X1 U7413 ( .A(n9788), .ZN(n9786) );
  NAND2_X1 U7414 ( .A1(n5747), .A2(n9786), .ZN(n9791) );
  INV_X1 U7415 ( .A(n9501), .ZN(n9332) );
  NAND2_X1 U7416 ( .A1(n9333), .A2(n9332), .ZN(n9276) );
  INV_X1 U7417 ( .A(n9500), .ZN(n8721) );
  OR2_X1 U7418 ( .A1(n9765), .A2(n8721), .ZN(n9331) );
  OR2_X1 U7419 ( .A1(n9333), .A2(n9332), .ZN(n9756) );
  AND2_X1 U7420 ( .A1(n9331), .A2(n9756), .ZN(n9421) );
  NAND2_X1 U7421 ( .A1(n9765), .A2(n8721), .ZN(n9330) );
  INV_X1 U7422 ( .A(n9499), .ZN(n9282) );
  OR2_X1 U7423 ( .A1(n9748), .A2(n9282), .ZN(n9284) );
  NAND2_X1 U7424 ( .A1(n9748), .A2(n9282), .ZN(n9423) );
  NAND2_X1 U7425 ( .A1(n9742), .A2(n9743), .ZN(n5748) );
  NAND2_X1 U7426 ( .A1(n5748), .A2(n9423), .ZN(n9446) );
  NAND2_X1 U7427 ( .A1(n9446), .A2(n9728), .ZN(n5749) );
  NAND2_X1 U7428 ( .A1(n5749), .A2(n9286), .ZN(n9711) );
  XNOR2_X1 U7429 ( .A(n9715), .B(n9497), .ZN(n9712) );
  NAND2_X1 U7430 ( .A1(n9711), .A2(n9712), .ZN(n5750) );
  INV_X1 U7431 ( .A(n9497), .ZN(n9287) );
  NAND2_X1 U7432 ( .A1(n9715), .A2(n9287), .ZN(n9292) );
  NAND2_X1 U7433 ( .A1(n5750), .A2(n9292), .ZN(n9696) );
  INV_X1 U7434 ( .A(n9496), .ZN(n8626) );
  OR2_X1 U7435 ( .A1(n9703), .A2(n8626), .ZN(n9295) );
  NAND2_X1 U7436 ( .A1(n9703), .A2(n8626), .ZN(n9296) );
  INV_X1 U7437 ( .A(n9494), .ZN(n5751) );
  OR2_X1 U7438 ( .A1(n9671), .A2(n5751), .ZN(n9647) );
  NAND2_X1 U7439 ( .A1(n9671), .A2(n5751), .ZN(n9431) );
  NAND2_X1 U7440 ( .A1(n9647), .A2(n9431), .ZN(n9663) );
  NAND2_X1 U7441 ( .A1(n4522), .A2(n5752), .ZN(n9665) );
  INV_X1 U7442 ( .A(n9493), .ZN(n5753) );
  OR2_X1 U7443 ( .A1(n9656), .A2(n5753), .ZN(n9377) );
  NAND2_X1 U7444 ( .A1(n9656), .A2(n5753), .ZN(n9307) );
  NAND2_X1 U7445 ( .A1(n9377), .A2(n9307), .ZN(n9648) );
  INV_X1 U7446 ( .A(n9647), .ZN(n5754) );
  NOR2_X1 U7447 ( .A1(n9648), .A2(n5754), .ZN(n5755) );
  NAND2_X1 U7448 ( .A1(n9665), .A2(n5755), .ZN(n9650) );
  NAND2_X1 U7449 ( .A1(n9650), .A2(n9307), .ZN(n9634) );
  OR2_X1 U7450 ( .A1(n9639), .A2(n8673), .ZN(n9309) );
  NAND2_X1 U7451 ( .A1(n9639), .A2(n8673), .ZN(n9222) );
  NAND2_X1 U7452 ( .A1(n9634), .A2(n9633), .ZN(n9618) );
  NAND2_X1 U7453 ( .A1(n9365), .A2(n9598), .ZN(n5756) );
  NAND2_X1 U7454 ( .A1(n5726), .A2(n9467), .ZN(n9364) );
  NAND2_X1 U7455 ( .A1(n7785), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5761) );
  NAND2_X1 U7456 ( .A1(n4494), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5760) );
  INV_X1 U7457 ( .A(n5757), .ZN(n7794) );
  NAND2_X1 U7458 ( .A1(n5518), .A2(n7794), .ZN(n5759) );
  NAND2_X1 U7459 ( .A1(n5079), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5758) );
  NAND4_X1 U7460 ( .A1(n5761), .A2(n5760), .A3(n5759), .A4(n5758), .ZN(n9490)
         );
  NAND2_X1 U7461 ( .A1(n9490), .A2(n9184), .ZN(n5763) );
  INV_X1 U7462 ( .A(n5454), .ZN(n10005) );
  NAND2_X1 U7463 ( .A1(n9491), .A2(n9197), .ZN(n5762) );
  NAND2_X1 U7464 ( .A1(n5763), .A2(n5762), .ZN(n8741) );
  AOI21_X1 U7465 ( .B1(n5765), .B2(n8745), .A(n9794), .ZN(n5766) );
  NAND2_X1 U7466 ( .A1(n5766), .A2(n7793), .ZN(n7874) );
  NAND2_X1 U7467 ( .A1(n5958), .A2(n10192), .ZN(n5771) );
  INV_X1 U7468 ( .A(n8745), .ZN(n7876) );
  INV_X1 U7469 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n5767) );
  NOR2_X1 U7470 ( .A1(n10192), .A2(n5767), .ZN(n5768) );
  NAND2_X1 U7471 ( .A1(n5771), .A2(n5770), .ZN(P1_U3550) );
  NAND2_X1 U7472 ( .A1(n5922), .A2(n5842), .ZN(n5836) );
  INV_X1 U7473 ( .A(n5836), .ZN(n5774) );
  NAND4_X1 U7474 ( .A1(n5776), .A2(n5832), .A3(n5820), .A4(n5775), .ZN(n5781)
         );
  NAND4_X1 U7475 ( .A1(n5825), .A2(n5779), .A3(n5778), .A4(n5777), .ZN(n5780)
         );
  NOR2_X1 U7476 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5792) );
  NOR2_X1 U7477 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5791) );
  NOR2_X1 U7478 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n5790) );
  NOR2_X1 U7479 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5789) );
  NAND2_X1 U7480 ( .A1(n5794), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5793) );
  MUX2_X1 U7481 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5793), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5797) );
  NAND2_X1 U7482 ( .A1(n6293), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5806) );
  MUX2_X1 U7483 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5806), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n5807) );
  NAND2_X1 U7484 ( .A1(n6374), .A2(n8106), .ZN(n5808) );
  NAND2_X1 U7485 ( .A1(n5808), .A2(n5951), .ZN(n5949) );
  NAND2_X1 U7486 ( .A1(n5949), .A2(n6322), .ZN(n5812) );
  NAND2_X1 U7487 ( .A1(n5812), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NAND2_X1 U7488 ( .A1(n5813), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5814) );
  XNOR2_X1 U7489 ( .A(n5814), .B(P2_IR_REG_18__SCAN_IN), .ZN(n9950) );
  INV_X1 U7490 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9114) );
  AOI22_X1 U7491 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n4914), .B1(n9950), .B2(
        n9114), .ZN(n9949) );
  OR2_X1 U7492 ( .A1(n5815), .A2(n4674), .ZN(n5816) );
  XNOR2_X1 U7493 ( .A(n5816), .B(P2_IR_REG_17__SCAN_IN), .ZN(n10341) );
  NAND2_X1 U7494 ( .A1(n5817), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5818) );
  XNOR2_X1 U7495 ( .A(n5818), .B(P2_IR_REG_16__SCAN_IN), .ZN(n10322) );
  INV_X1 U7496 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n5880) );
  INV_X1 U7497 ( .A(n10322), .ZN(n6831) );
  AOI22_X1 U7498 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n6831), .B1(n10322), .B2(
        n5880), .ZN(n10325) );
  NOR2_X1 U7499 ( .A1(n5819), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5861) );
  AND2_X1 U7500 ( .A1(n5861), .A2(n5820), .ZN(n5831) );
  NOR2_X1 U7501 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5821) );
  NAND2_X1 U7502 ( .A1(n5831), .A2(n5821), .ZN(n5868) );
  OAI21_X1 U7503 ( .B1(n5870), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5829) );
  INV_X1 U7504 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5822) );
  NAND2_X1 U7505 ( .A1(n5829), .A2(n5822), .ZN(n5823) );
  NAND2_X1 U7506 ( .A1(n5823), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5826) );
  NAND2_X1 U7507 ( .A1(n5826), .A2(n5825), .ZN(n5828) );
  NAND2_X1 U7508 ( .A1(n5828), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5824) );
  XNOR2_X1 U7509 ( .A(n5824), .B(P2_IR_REG_15__SCAN_IN), .ZN(n10307) );
  OR2_X1 U7510 ( .A1(n5826), .A2(n5825), .ZN(n5827) );
  NAND2_X1 U7511 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n6522), .ZN(n5877) );
  INV_X1 U7512 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6135) );
  AOI22_X1 U7513 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n6522), .B1(n10290), .B2(
        n6135), .ZN(n10293) );
  XNOR2_X1 U7514 ( .A(n5829), .B(P2_IR_REG_13__SCAN_IN), .ZN(n10274) );
  NAND2_X1 U7515 ( .A1(n5870), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5830) );
  XNOR2_X1 U7516 ( .A(n5830), .B(P2_IR_REG_12__SCAN_IN), .ZN(n10257) );
  INV_X1 U7517 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n5874) );
  INV_X1 U7518 ( .A(n10257), .ZN(n6487) );
  AOI22_X1 U7519 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n6487), .B1(n10257), .B2(
        n5874), .ZN(n10260) );
  OR2_X1 U7520 ( .A1(n5831), .A2(n4674), .ZN(n5835) );
  NAND2_X1 U7521 ( .A1(n5835), .A2(n5832), .ZN(n5833) );
  NAND2_X1 U7522 ( .A1(n5833), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5834) );
  XNOR2_X1 U7523 ( .A(n5834), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10225) );
  INV_X1 U7524 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n5867) );
  INV_X1 U7525 ( .A(n10225), .ZN(n6462) );
  AOI22_X1 U7526 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n6462), .B1(n10225), .B2(
        n5867), .ZN(n10228) );
  XNOR2_X1 U7527 ( .A(n5835), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10209) );
  NAND2_X1 U7528 ( .A1(n4601), .A2(n5840), .ZN(n5853) );
  OAI21_X1 U7529 ( .B1(n5853), .B2(P2_IR_REG_5__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5837) );
  MUX2_X1 U7530 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5837), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5838) );
  AND2_X1 U7531 ( .A1(n5838), .A2(n5819), .ZN(n6869) );
  INV_X1 U7532 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7006) );
  NAND2_X1 U7533 ( .A1(n5839), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5841) );
  XNOR2_X1 U7534 ( .A(n5841), .B(n5840), .ZN(n6984) );
  INV_X1 U7535 ( .A(n7036), .ZN(n5893) );
  INV_X1 U7536 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10380) );
  INV_X1 U7537 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5844) );
  NAND2_X1 U7538 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5843) );
  XNOR2_X1 U7539 ( .A(n5844), .B(n5843), .ZN(n10193) );
  NAND2_X1 U7540 ( .A1(n4492), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5846) );
  INV_X1 U7541 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5988) );
  NOR3_X1 U7542 ( .A1(n4492), .A2(P2_IR_REG_0__SCAN_IN), .A3(n5988), .ZN(n5845) );
  AOI21_X1 U7543 ( .B1(n10193), .B2(n5846), .A(n5845), .ZN(n10195) );
  INV_X1 U7544 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10194) );
  INV_X1 U7545 ( .A(n4492), .ZN(n5847) );
  OAI22_X1 U7546 ( .A1(n10195), .A2(n10194), .B1(n5988), .B2(n5847), .ZN(n7028) );
  MUX2_X1 U7547 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10380), .S(n7036), .Z(n7029)
         );
  NAND2_X1 U7548 ( .A1(n7028), .A2(n7029), .ZN(n7027) );
  OAI21_X1 U7549 ( .B1(n5893), .B2(n10380), .A(n7027), .ZN(n5851) );
  XNOR2_X1 U7550 ( .A(n5849), .B(n5848), .ZN(n6999) );
  INV_X1 U7551 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10369) );
  MUX2_X1 U7552 ( .A(n10369), .B(P2_REG2_REG_4__SCAN_IN), .S(n6984), .Z(n6968)
         );
  NAND2_X1 U7553 ( .A1(n5853), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5855) );
  XNOR2_X1 U7554 ( .A(n5855), .B(n5854), .ZN(n6437) );
  INV_X1 U7555 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6747) );
  INV_X1 U7556 ( .A(n6437), .ZN(n6845) );
  OAI22_X1 U7557 ( .A1(n6840), .A2(n6747), .B1(n5856), .B2(n6845), .ZN(n6861)
         );
  MUX2_X1 U7558 ( .A(n7006), .B(P2_REG2_REG_6__SCAN_IN), .S(n6869), .Z(n6862)
         );
  NAND2_X1 U7559 ( .A1(n6861), .A2(n6862), .ZN(n6860) );
  NAND2_X1 U7560 ( .A1(n5819), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5857) );
  MUX2_X1 U7561 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5857), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n5859) );
  INV_X1 U7562 ( .A(n5861), .ZN(n5858) );
  NAND2_X1 U7563 ( .A1(n5859), .A2(n5858), .ZN(n7084) );
  INV_X1 U7564 ( .A(n7084), .ZN(n6060) );
  XNOR2_X1 U7565 ( .A(n5860), .B(n6060), .ZN(n7090) );
  INV_X1 U7566 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n5863) );
  OR2_X1 U7567 ( .A1(n5861), .A2(n4674), .ZN(n5862) );
  XNOR2_X1 U7568 ( .A(n5862), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6886) );
  MUX2_X1 U7569 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n5863), .S(n6886), .Z(n6874)
         );
  INV_X1 U7570 ( .A(n6872), .ZN(n5864) );
  NAND2_X1 U7571 ( .A1(n6456), .A2(n5865), .ZN(n5866) );
  NAND2_X1 U7572 ( .A1(n5868), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5869) );
  MUX2_X1 U7573 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5869), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n5871) );
  INV_X1 U7574 ( .A(n10241), .ZN(n6482) );
  NAND2_X1 U7575 ( .A1(n5872), .A2(n6482), .ZN(n5873) );
  XNOR2_X1 U7576 ( .A(n5872), .B(n10241), .ZN(n10243) );
  NAND2_X1 U7577 ( .A1(n6497), .A2(n5875), .ZN(n5876) );
  XNOR2_X1 U7578 ( .A(n5875), .B(n10274), .ZN(n10276) );
  NAND2_X1 U7579 ( .A1(n6601), .A2(n5878), .ZN(n5879) );
  NAND2_X1 U7580 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n10309), .ZN(n10308) );
  NAND2_X1 U7581 ( .A1(n5879), .A2(n10308), .ZN(n10324) );
  NAND2_X1 U7582 ( .A1(n10325), .A2(n10324), .ZN(n10323) );
  OAI21_X1 U7583 ( .B1(n10322), .B2(n5880), .A(n10323), .ZN(n5881) );
  NAND2_X1 U7584 ( .A1(n6834), .A2(n5881), .ZN(n5882) );
  NAND2_X1 U7585 ( .A1(n5882), .A2(n10342), .ZN(n9948) );
  INV_X1 U7586 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n5885) );
  NAND2_X1 U7587 ( .A1(n5883), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5884) );
  MUX2_X1 U7588 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n5885), .S(n8124), .Z(n5887)
         );
  NOR2_X1 U7589 ( .A1(n5886), .A2(P2_U3151), .ZN(n8556) );
  INV_X1 U7590 ( .A(n5946), .ZN(n6890) );
  INV_X1 U7591 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8483) );
  XNOR2_X1 U7592 ( .A(n8124), .B(n8483), .ZN(n5943) );
  MUX2_X1 U7593 ( .A(n5887), .B(n5943), .S(n5948), .Z(n5920) );
  MUX2_X1 U7594 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n5948), .Z(n5914) );
  INV_X1 U7595 ( .A(n5914), .ZN(n5915) );
  INV_X1 U7596 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7539) );
  INV_X1 U7597 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7532) );
  MUX2_X1 U7598 ( .A(n7539), .B(n7532), .S(n5948), .Z(n5913) );
  MUX2_X1 U7599 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n5948), .Z(n5911) );
  INV_X1 U7600 ( .A(n5911), .ZN(n5912) );
  MUX2_X1 U7601 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n5948), .Z(n5909) );
  INV_X1 U7602 ( .A(n5909), .ZN(n5910) );
  MUX2_X1 U7603 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n5948), .Z(n5907) );
  INV_X1 U7604 ( .A(n5907), .ZN(n5908) );
  INV_X1 U7605 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7186) );
  INV_X1 U7606 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6101) );
  MUX2_X1 U7607 ( .A(n7186), .B(n6101), .S(n5948), .Z(n5906) );
  MUX2_X1 U7608 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n5948), .Z(n5904) );
  INV_X1 U7609 ( .A(n5904), .ZN(n5905) );
  MUX2_X1 U7610 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n5948), .Z(n5888) );
  INV_X1 U7611 ( .A(n5888), .ZN(n5903) );
  XNOR2_X1 U7612 ( .A(n5888), .B(n6456), .ZN(n10218) );
  INV_X1 U7613 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6065) );
  MUX2_X1 U7614 ( .A(n5863), .B(n6065), .S(n5948), .Z(n5902) );
  MUX2_X1 U7615 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n5948), .Z(n5899) );
  NOR2_X1 U7616 ( .A1(n5899), .A2(n7084), .ZN(n5901) );
  INV_X1 U7617 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6023) );
  MUX2_X1 U7618 ( .A(n7006), .B(n6023), .S(n5948), .Z(n5898) );
  MUX2_X1 U7619 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n5948), .Z(n5895) );
  MUX2_X1 U7620 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n5889), .Z(n5890) );
  XOR2_X1 U7621 ( .A(n10193), .B(n5890), .Z(n10204) );
  INV_X1 U7622 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5987) );
  MUX2_X1 U7623 ( .A(n5988), .B(n5987), .S(n5948), .Z(n6891) );
  NAND2_X1 U7624 ( .A1(n6891), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n10203) );
  AOI22_X1 U7625 ( .A1(n10204), .A2(n10203), .B1(n5890), .B2(n10193), .ZN(
        n7030) );
  MUX2_X1 U7626 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n5948), .Z(n5891) );
  XNOR2_X1 U7627 ( .A(n5891), .B(n7036), .ZN(n7031) );
  INV_X1 U7628 ( .A(n5891), .ZN(n5892) );
  MUX2_X1 U7629 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n5948), .Z(n5894) );
  XNOR2_X1 U7630 ( .A(n5894), .B(n6999), .ZN(n6991) );
  NOR2_X1 U7631 ( .A1(n5894), .A2(n6999), .ZN(n6979) );
  XNOR2_X1 U7632 ( .A(n5895), .B(n6984), .ZN(n6978) );
  MUX2_X1 U7633 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n5948), .Z(n5896) );
  XNOR2_X1 U7634 ( .A(n5896), .B(n6437), .ZN(n6837) );
  INV_X1 U7635 ( .A(n5896), .ZN(n5897) );
  XNOR2_X1 U7636 ( .A(n5898), .B(n6869), .ZN(n6856) );
  AOI21_X1 U7637 ( .B1(n5899), .B2(n7084), .A(n5901), .ZN(n5900) );
  INV_X1 U7638 ( .A(n5900), .ZN(n7082) );
  NOR2_X1 U7639 ( .A1(n7083), .A2(n7082), .ZN(n7081) );
  XNOR2_X1 U7640 ( .A(n5902), .B(n6886), .ZN(n6877) );
  XNOR2_X1 U7641 ( .A(n5904), .B(n6462), .ZN(n10235) );
  XNOR2_X1 U7642 ( .A(n5906), .B(n10241), .ZN(n10250) );
  XNOR2_X1 U7643 ( .A(n5907), .B(n6487), .ZN(n10267) );
  XNOR2_X1 U7644 ( .A(n5909), .B(n6497), .ZN(n10283) );
  NOR2_X1 U7645 ( .A1(n10284), .A2(n10283), .ZN(n10282) );
  XNOR2_X1 U7646 ( .A(n5911), .B(n6522), .ZN(n10300) );
  XNOR2_X1 U7647 ( .A(n10307), .B(n5913), .ZN(n10315) );
  XNOR2_X1 U7648 ( .A(n5914), .B(n6831), .ZN(n10332) );
  NOR2_X1 U7649 ( .A1(n10333), .A2(n10332), .ZN(n10331) );
  AOI21_X1 U7650 ( .B1(n10322), .B2(n5915), .A(n10331), .ZN(n10353) );
  MUX2_X1 U7651 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n5948), .Z(n5916) );
  XNOR2_X1 U7652 ( .A(n5916), .B(n6834), .ZN(n10352) );
  INV_X1 U7653 ( .A(n5916), .ZN(n5917) );
  NAND2_X1 U7654 ( .A1(n5917), .A2(n10341), .ZN(n5918) );
  MUX2_X1 U7655 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n5948), .Z(n5919) );
  NOR2_X1 U7656 ( .A1(n5921), .A2(n10354), .ZN(n5956) );
  INV_X1 U7657 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n5942) );
  AOI22_X1 U7658 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n4914), .B1(n9950), .B2(
        n5942), .ZN(n9940) );
  INV_X1 U7659 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n7680) );
  AOI22_X1 U7660 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n6831), .B1(n10322), .B2(
        n7680), .ZN(n10328) );
  INV_X1 U7661 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9120) );
  AOI22_X1 U7662 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n6522), .B1(n10290), .B2(
        n9120), .ZN(n10296) );
  INV_X1 U7663 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9052) );
  AOI22_X1 U7664 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n6487), .B1(n10257), .B2(
        n9052), .ZN(n10263) );
  INV_X1 U7665 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10442) );
  AOI22_X1 U7666 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n6462), .B1(n10225), .B2(
        n10442), .ZN(n10231) );
  MUX2_X1 U7667 ( .A(n6065), .B(P2_REG1_REG_8__SCAN_IN), .S(n6886), .Z(n6879)
         );
  NAND2_X1 U7668 ( .A1(n4492), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5924) );
  NOR3_X1 U7669 ( .A1(n4492), .A2(P2_IR_REG_0__SCAN_IN), .A3(n5987), .ZN(n5923) );
  AOI21_X1 U7670 ( .B1(n10193), .B2(n5924), .A(n5923), .ZN(n10196) );
  INV_X1 U7671 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n5925) );
  OAI21_X1 U7672 ( .B1(n10196), .B2(n5925), .A(n5924), .ZN(n7021) );
  INV_X1 U7673 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6593) );
  XNOR2_X1 U7674 ( .A(n7036), .B(n6593), .ZN(n7022) );
  AOI22_X1 U7675 ( .A1(n7021), .A2(n7022), .B1(P2_REG1_REG_2__SCAN_IN), .B2(
        n7036), .ZN(n5926) );
  XNOR2_X1 U7676 ( .A(n5926), .B(n6999), .ZN(n6985) );
  INV_X1 U7677 ( .A(n5926), .ZN(n5927) );
  INV_X1 U7678 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9037) );
  MUX2_X1 U7679 ( .A(n9037), .B(P2_REG1_REG_4__SCAN_IN), .S(n6984), .Z(n6973)
         );
  INV_X1 U7680 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5929) );
  OAI22_X1 U7681 ( .A1(n6839), .A2(n5929), .B1(n6845), .B2(n5928), .ZN(n6858)
         );
  MUX2_X1 U7682 ( .A(n6023), .B(P2_REG1_REG_6__SCAN_IN), .S(n6869), .Z(n6859)
         );
  NAND2_X1 U7683 ( .A1(n6858), .A2(n6859), .ZN(n6857) );
  NAND2_X1 U7684 ( .A1(n7084), .A2(n5930), .ZN(n5931) );
  NAND2_X1 U7685 ( .A1(n6879), .A2(n6880), .ZN(n6878) );
  NAND2_X1 U7686 ( .A1(n6456), .A2(n5932), .ZN(n5933) );
  NAND2_X1 U7687 ( .A1(n10231), .A2(n10230), .ZN(n10229) );
  OAI21_X1 U7688 ( .B1(n10225), .B2(n10442), .A(n10229), .ZN(n5934) );
  NAND2_X1 U7689 ( .A1(n5934), .A2(n6482), .ZN(n5935) );
  XNOR2_X1 U7690 ( .A(n5934), .B(n10241), .ZN(n10245) );
  NAND2_X1 U7691 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n10245), .ZN(n10244) );
  NAND2_X1 U7692 ( .A1(n6497), .A2(n5936), .ZN(n5937) );
  NAND2_X1 U7693 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n10278), .ZN(n10277) );
  NAND2_X1 U7694 ( .A1(n6601), .A2(n5938), .ZN(n5939) );
  NAND2_X1 U7695 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n10311), .ZN(n10310) );
  NAND2_X1 U7696 ( .A1(n6834), .A2(n5940), .ZN(n5941) );
  NAND2_X1 U7697 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n10345), .ZN(n10344) );
  NAND2_X1 U7698 ( .A1(n5941), .A2(n10344), .ZN(n9939) );
  NAND2_X1 U7699 ( .A1(n9940), .A2(n9939), .ZN(n9938) );
  OAI21_X1 U7700 ( .B1(n9950), .B2(n5942), .A(n9938), .ZN(n5945) );
  INV_X1 U7701 ( .A(n5943), .ZN(n5944) );
  XNOR2_X1 U7702 ( .A(n5945), .B(n5944), .ZN(n5947) );
  NOR2_X1 U7703 ( .A1(n5948), .A2(P2_U3151), .ZN(n8559) );
  AND2_X1 U7704 ( .A1(n5949), .A2(n8559), .ZN(n5950) );
  NAND2_X1 U7705 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3151), .ZN(n5954) );
  INV_X1 U7706 ( .A(n5951), .ZN(n6695) );
  NOR2_X1 U7707 ( .A1(n6374), .A2(n6695), .ZN(n5952) );
  NAND2_X1 U7708 ( .A1(n10339), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5953) );
  OAI211_X1 U7709 ( .C1(n9945), .C2(n7138), .A(n5954), .B(n5953), .ZN(n5955)
         );
  AND2_X1 U7710 ( .A1(n10175), .A2(n5959), .ZN(n6387) );
  NOR2_X1 U7711 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6014) );
  INV_X1 U7712 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6706) );
  NAND2_X1 U7713 ( .A1(n6014), .A2(n6706), .ZN(n6037) );
  NOR2_X1 U7714 ( .A1(n6053), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6052) );
  INV_X1 U7715 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U7716 ( .A1(n6066), .A2(n7158), .ZN(n6093) );
  NAND2_X1 U7717 ( .A1(n6113), .A2(n8206), .ZN(n6133) );
  INV_X1 U7718 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5963) );
  INV_X1 U7719 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5964) );
  INV_X1 U7720 ( .A(n6190), .ZN(n6191) );
  NAND2_X1 U7721 ( .A1(n6181), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U7722 ( .A1(n6191), .A2(n5965), .ZN(n8416) );
  XNOR2_X2 U7723 ( .A(n5969), .B(n5968), .ZN(n5973) );
  NAND2_X4 U7724 ( .A1(n5975), .A2(n5974), .ZN(n6285) );
  NAND2_X1 U7725 ( .A1(n8416), .A2(n6266), .ZN(n5978) );
  AND2_X4 U7726 ( .A1(n5973), .A2(n8553), .ZN(n6314) );
  AOI22_X1 U7727 ( .A1(n6314), .A2(P2_REG0_REG_19__SCAN_IN), .B1(n6315), .B2(
        P2_REG1_REG_19__SCAN_IN), .ZN(n5977) );
  CLKBUF_X3 U7728 ( .A(n6013), .Z(n7902) );
  OR2_X1 U7729 ( .A1(n7902), .A2(n5885), .ZN(n5976) );
  NAND2_X1 U7730 ( .A1(n7136), .A2(n7891), .ZN(n5980) );
  AOI22_X1 U7731 ( .A1(n6176), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6175), .B2(
        n8124), .ZN(n5979) );
  NAND2_X1 U7732 ( .A1(n6314), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5986) );
  INV_X1 U7733 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n5981) );
  OR2_X1 U7734 ( .A1(n6285), .A2(n5981), .ZN(n5985) );
  OR2_X1 U7735 ( .A1(n6013), .A2(n10194), .ZN(n5984) );
  NAND2_X1 U7736 ( .A1(n5982), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5983) );
  NAND2_X1 U7737 ( .A1(n6314), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5993) );
  OR2_X1 U7738 ( .A1(n7900), .A2(n5987), .ZN(n5992) );
  OR2_X1 U7739 ( .A1(n6013), .A2(n5988), .ZN(n5991) );
  INV_X1 U7740 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n5989) );
  OR2_X1 U7741 ( .A1(n6285), .A2(n5989), .ZN(n5990) );
  NAND2_X1 U7742 ( .A1(n4835), .A2(SI_0_), .ZN(n5994) );
  XNOR2_X1 U7743 ( .A(n5994), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8564) );
  MUX2_X1 U7744 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8564), .S(n6322), .Z(n6673) );
  NAND2_X1 U7745 ( .A1(n5995), .A2(n10383), .ZN(n5996) );
  NAND2_X1 U7746 ( .A1(n5982), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6000) );
  OR2_X1 U7747 ( .A1(n6013), .A2(n10380), .ZN(n5998) );
  INV_X1 U7748 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10372) );
  OR2_X1 U7749 ( .A1(n6285), .A2(n10372), .ZN(n5997) );
  OR2_X1 U7750 ( .A1(n6080), .A2(n6430), .ZN(n6002) );
  OR2_X1 U7751 ( .A1(n6031), .A2(n4589), .ZN(n6001) );
  INV_X1 U7752 ( .A(n7971), .ZN(n6585) );
  NAND2_X1 U7753 ( .A1(n6942), .A2(n10371), .ZN(n7012) );
  NAND2_X1 U7754 ( .A1(n5982), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6008) );
  INV_X1 U7755 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6003) );
  OR2_X1 U7756 ( .A1(n6050), .A2(n6003), .ZN(n6007) );
  OR2_X1 U7757 ( .A1(n6285), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6006) );
  INV_X1 U7758 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6004) );
  OR2_X1 U7759 ( .A1(n6013), .A2(n6004), .ZN(n6005) );
  OR2_X1 U7760 ( .A1(n6080), .A2(n6431), .ZN(n6010) );
  OR2_X1 U7761 ( .A1(n6031), .A2(n6432), .ZN(n6009) );
  OAI211_X1 U7762 ( .C1(n6322), .C2(n6999), .A(n6010), .B(n6009), .ZN(n10390)
         );
  NAND2_X1 U7763 ( .A1(n6692), .A2(n7017), .ZN(n6011) );
  AND2_X1 U7764 ( .A1(n7012), .A2(n6011), .ZN(n6012) );
  NAND2_X1 U7765 ( .A1(n7013), .A2(n6012), .ZN(n6578) );
  NAND2_X1 U7766 ( .A1(n6314), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6019) );
  OR2_X1 U7767 ( .A1(n7900), .A2(n9037), .ZN(n6018) );
  OR2_X1 U7768 ( .A1(n6013), .A2(n10369), .ZN(n6017) );
  INV_X1 U7769 ( .A(n6014), .ZN(n6035) );
  NAND2_X1 U7770 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6015) );
  AND2_X1 U7771 ( .A1(n6035), .A2(n6015), .ZN(n10366) );
  OR2_X1 U7772 ( .A1(n6285), .A2(n10366), .ZN(n6016) );
  OR2_X1 U7773 ( .A1(n6031), .A2(n6434), .ZN(n6020) );
  INV_X1 U7774 ( .A(n6579), .ZN(n6021) );
  NOR2_X1 U7775 ( .A1(n7981), .A2(n6021), .ZN(n6022) );
  NAND2_X1 U7776 ( .A1(n6578), .A2(n6022), .ZN(n6737) );
  NAND2_X1 U7777 ( .A1(n6314), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6028) );
  OR2_X1 U7778 ( .A1(n7900), .A2(n6023), .ZN(n6027) );
  NAND2_X1 U7779 ( .A1(n6037), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6024) );
  AND2_X1 U7780 ( .A1(n6053), .A2(n6024), .ZN(n7007) );
  OR2_X1 U7781 ( .A1(n6285), .A2(n7007), .ZN(n6026) );
  OR2_X1 U7782 ( .A1(n7902), .A2(n7006), .ZN(n6025) );
  OR2_X1 U7783 ( .A1(n6443), .A2(n6080), .ZN(n6030) );
  AOI22_X1 U7784 ( .A1(n6176), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6175), .B2(
        n6869), .ZN(n6029) );
  NAND2_X1 U7785 ( .A1(n6030), .A2(n6029), .ZN(n10398) );
  NAND2_X1 U7786 ( .A1(n7063), .A2(n7008), .ZN(n6046) );
  INV_X1 U7787 ( .A(n8287), .ZN(n6754) );
  INV_X1 U7788 ( .A(n6694), .ZN(n10364) );
  NAND2_X1 U7789 ( .A1(n6754), .A2(n10364), .ZN(n6738) );
  OR2_X1 U7790 ( .A1(n6438), .A2(n6080), .ZN(n6034) );
  OR2_X1 U7791 ( .A1(n6322), .A2(n6437), .ZN(n6033) );
  OR2_X1 U7792 ( .A1(n7893), .A2(n6439), .ZN(n6032) );
  NAND2_X1 U7793 ( .A1(n5982), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6042) );
  OR2_X1 U7794 ( .A1(n7902), .A2(n6747), .ZN(n6041) );
  NAND2_X1 U7795 ( .A1(n6035), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6036) );
  AND2_X1 U7796 ( .A1(n6037), .A2(n6036), .ZN(n6748) );
  OR2_X1 U7797 ( .A1(n6285), .A2(n6748), .ZN(n6040) );
  INV_X1 U7798 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6038) );
  OR2_X1 U7799 ( .A1(n6050), .A2(n6038), .ZN(n6039) );
  NAND2_X1 U7800 ( .A1(n6736), .A2(n6043), .ZN(n6044) );
  AND2_X1 U7801 ( .A1(n6738), .A2(n6044), .ZN(n6739) );
  AND2_X1 U7802 ( .A1(n6046), .A2(n6739), .ZN(n6045) );
  NAND2_X1 U7803 ( .A1(n6737), .A2(n6045), .ZN(n6049) );
  INV_X1 U7804 ( .A(n6046), .ZN(n6047) );
  NAND2_X1 U7805 ( .A1(n10394), .A2(n8286), .ZN(n7000) );
  NAND2_X1 U7806 ( .A1(n6049), .A2(n6048), .ZN(n7099) );
  NAND2_X1 U7807 ( .A1(n6315), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6059) );
  INV_X1 U7808 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6051) );
  OR2_X1 U7809 ( .A1(n6050), .A2(n6051), .ZN(n6058) );
  INV_X1 U7810 ( .A(n6052), .ZN(n6067) );
  NAND2_X1 U7811 ( .A1(n6053), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6054) );
  AND2_X1 U7812 ( .A1(n6067), .A2(n6054), .ZN(n7104) );
  OR2_X1 U7813 ( .A1(n6285), .A2(n7104), .ZN(n6057) );
  INV_X1 U7814 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6055) );
  OR2_X1 U7815 ( .A1(n7902), .A2(n6055), .ZN(n6056) );
  OR2_X1 U7816 ( .A1(n6446), .A2(n6080), .ZN(n6062) );
  AOI22_X1 U7817 ( .A1(n6176), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6175), .B2(
        n6060), .ZN(n6061) );
  NAND2_X1 U7818 ( .A1(n6062), .A2(n6061), .ZN(n10406) );
  AND2_X1 U7819 ( .A1(n8284), .A2(n10406), .ZN(n6064) );
  OR2_X1 U7820 ( .A1(n8284), .A2(n10406), .ZN(n6063) );
  OAI21_X2 U7821 ( .B1(n7099), .B2(n6064), .A(n6063), .ZN(n6947) );
  NAND2_X1 U7822 ( .A1(n6314), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6072) );
  OR2_X1 U7823 ( .A1(n7900), .A2(n6065), .ZN(n6071) );
  INV_X1 U7824 ( .A(n6066), .ZN(n6082) );
  NAND2_X1 U7825 ( .A1(n6067), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6068) );
  AND2_X1 U7826 ( .A1(n6082), .A2(n6068), .ZN(n6953) );
  OR2_X1 U7827 ( .A1(n6285), .A2(n6953), .ZN(n6070) );
  OR2_X1 U7828 ( .A1(n7902), .A2(n5863), .ZN(n6069) );
  NAND4_X1 U7829 ( .A1(n6072), .A2(n6071), .A3(n6070), .A4(n6069), .ZN(n8282)
         );
  NAND2_X1 U7830 ( .A1(n6947), .A2(n7152), .ZN(n6075) );
  OR2_X1 U7831 ( .A1(n6449), .A2(n6080), .ZN(n6074) );
  AOI22_X1 U7832 ( .A1(n6176), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6175), .B2(
        n6886), .ZN(n6073) );
  INV_X1 U7833 ( .A(n7114), .ZN(n10407) );
  NAND2_X1 U7834 ( .A1(n6075), .A2(n10407), .ZN(n6078) );
  INV_X1 U7835 ( .A(n6947), .ZN(n6076) );
  NAND2_X1 U7836 ( .A1(n6076), .A2(n8282), .ZN(n6077) );
  AOI22_X1 U7837 ( .A1(n6176), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6175), .B2(
        n10209), .ZN(n6079) );
  NAND2_X1 U7838 ( .A1(n6314), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6087) );
  INV_X1 U7839 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6081) );
  OR2_X1 U7840 ( .A1(n7900), .A2(n6081), .ZN(n6086) );
  NAND2_X1 U7841 ( .A1(n6082), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6083) );
  AND2_X1 U7842 ( .A1(n6093), .A2(n6083), .ZN(n7201) );
  OR2_X1 U7843 ( .A1(n6285), .A2(n7201), .ZN(n6085) );
  INV_X1 U7844 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7202) );
  OR2_X1 U7845 ( .A1(n7902), .A2(n7202), .ZN(n6084) );
  INV_X1 U7846 ( .A(n7426), .ZN(n8281) );
  NAND2_X1 U7847 ( .A1(n6088), .A2(n7426), .ZN(n6089) );
  NAND2_X1 U7848 ( .A1(n6460), .A2(n7891), .ZN(n6091) );
  AOI22_X1 U7849 ( .A1(n6176), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6175), .B2(
        n10225), .ZN(n6090) );
  INV_X1 U7850 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n6092) );
  OR2_X1 U7851 ( .A1(n6050), .A2(n6092), .ZN(n6098) );
  OR2_X1 U7852 ( .A1(n7900), .A2(n10442), .ZN(n6097) );
  NAND2_X1 U7853 ( .A1(n6093), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6094) );
  AND2_X1 U7854 ( .A1(n6102), .A2(n6094), .ZN(n7430) );
  OR2_X1 U7855 ( .A1(n6285), .A2(n7430), .ZN(n6096) );
  OR2_X1 U7856 ( .A1(n7902), .A2(n5867), .ZN(n6095) );
  NAND4_X1 U7857 ( .A1(n6098), .A2(n6097), .A3(n6096), .A4(n6095), .ZN(n8280)
         );
  OR2_X1 U7858 ( .A1(n10419), .A2(n7457), .ZN(n7181) );
  NAND2_X1 U7859 ( .A1(n6480), .A2(n7891), .ZN(n6100) );
  AOI22_X1 U7860 ( .A1(n6176), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6175), .B2(
        n10241), .ZN(n6099) );
  NAND2_X1 U7861 ( .A1(n6100), .A2(n6099), .ZN(n10428) );
  NAND2_X1 U7862 ( .A1(n6314), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6107) );
  OR2_X1 U7863 ( .A1(n7900), .A2(n6101), .ZN(n6106) );
  NAND2_X1 U7864 ( .A1(n6102), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6103) );
  AND2_X1 U7865 ( .A1(n6114), .A2(n6103), .ZN(n7464) );
  OR2_X1 U7866 ( .A1(n6285), .A2(n7464), .ZN(n6105) );
  OR2_X1 U7867 ( .A1(n7902), .A2(n7186), .ZN(n6104) );
  INV_X1 U7868 ( .A(n7558), .ZN(n8279) );
  NAND2_X1 U7869 ( .A1(n10428), .A2(n8279), .ZN(n6108) );
  AND2_X1 U7870 ( .A1(n7181), .A2(n6108), .ZN(n6110) );
  INV_X1 U7871 ( .A(n6108), .ZN(n6109) );
  OR2_X1 U7872 ( .A1(n10428), .A2(n7558), .ZN(n8010) );
  NAND2_X1 U7873 ( .A1(n10428), .A2(n7558), .ZN(n8006) );
  NAND2_X1 U7874 ( .A1(n6486), .A2(n7891), .ZN(n6112) );
  AOI22_X1 U7875 ( .A1(n6176), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6175), .B2(
        n10257), .ZN(n6111) );
  NAND2_X1 U7876 ( .A1(n6112), .A2(n6111), .ZN(n7568) );
  NAND2_X1 U7877 ( .A1(n6314), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6119) );
  OR2_X1 U7878 ( .A1(n7900), .A2(n9052), .ZN(n6118) );
  OR2_X1 U7879 ( .A1(n7902), .A2(n5874), .ZN(n6117) );
  INV_X1 U7880 ( .A(n6113), .ZN(n6123) );
  NAND2_X1 U7881 ( .A1(n6114), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6115) );
  AND2_X1 U7882 ( .A1(n6123), .A2(n6115), .ZN(n7566) );
  OR2_X1 U7883 ( .A1(n6285), .A2(n7566), .ZN(n6116) );
  INV_X1 U7884 ( .A(n7749), .ZN(n8278) );
  AND2_X1 U7885 ( .A1(n7568), .A2(n8278), .ZN(n6120) );
  OAI22_X1 U7886 ( .A1(n7254), .A2(n6120), .B1(n8278), .B2(n7568), .ZN(n7414)
         );
  NAND2_X1 U7887 ( .A1(n6496), .A2(n7891), .ZN(n6122) );
  AOI22_X1 U7888 ( .A1(n6176), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6175), .B2(
        n10274), .ZN(n6121) );
  NAND2_X1 U7889 ( .A1(n6314), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6128) );
  INV_X1 U7890 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7421) );
  OR2_X1 U7891 ( .A1(n7900), .A2(n7421), .ZN(n6127) );
  NAND2_X1 U7892 ( .A1(n6123), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6124) );
  AND2_X1 U7893 ( .A1(n6133), .A2(n6124), .ZN(n8209) );
  OR2_X1 U7894 ( .A1(n6285), .A2(n8209), .ZN(n6126) );
  INV_X1 U7895 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7454) );
  OR2_X1 U7896 ( .A1(n7902), .A2(n7454), .ZN(n6125) );
  OR2_X1 U7897 ( .A1(n8217), .A2(n8277), .ZN(n8022) );
  INV_X1 U7898 ( .A(n8022), .ZN(n6129) );
  OR2_X1 U7899 ( .A1(n7414), .A2(n6129), .ZN(n6130) );
  NAND2_X1 U7900 ( .A1(n8217), .A2(n8277), .ZN(n8023) );
  NAND2_X1 U7901 ( .A1(n6516), .A2(n7891), .ZN(n6132) );
  AOI22_X1 U7902 ( .A1(n6176), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6175), .B2(
        n10290), .ZN(n6131) );
  NAND2_X1 U7903 ( .A1(n6314), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6139) );
  OR2_X1 U7904 ( .A1(n7900), .A2(n9120), .ZN(n6138) );
  NAND2_X1 U7905 ( .A1(n6133), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6134) );
  AND2_X1 U7906 ( .A1(n6144), .A2(n6134), .ZN(n7755) );
  OR2_X1 U7907 ( .A1(n6285), .A2(n7755), .ZN(n6137) );
  OR2_X1 U7908 ( .A1(n7902), .A2(n6135), .ZN(n6136) );
  INV_X1 U7909 ( .A(n8259), .ZN(n8276) );
  AND2_X1 U7910 ( .A1(n7751), .A2(n8276), .ZN(n6140) );
  NAND2_X1 U7911 ( .A1(n6599), .A2(n7891), .ZN(n6142) );
  AOI22_X1 U7912 ( .A1(n6176), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n10307), 
        .B2(n6175), .ZN(n6141) );
  NAND2_X1 U7913 ( .A1(n6314), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6149) );
  OR2_X1 U7914 ( .A1(n7900), .A2(n7532), .ZN(n6148) );
  INV_X1 U7915 ( .A(n6143), .ZN(n6155) );
  NAND2_X1 U7916 ( .A1(n6144), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6145) );
  AND2_X1 U7917 ( .A1(n6155), .A2(n6145), .ZN(n7540) );
  OR2_X1 U7918 ( .A1(n6285), .A2(n7540), .ZN(n6147) );
  OR2_X1 U7919 ( .A1(n7902), .A2(n7539), .ZN(n6146) );
  NAND2_X1 U7920 ( .A1(n8250), .A2(n8275), .ZN(n6150) );
  NAND2_X1 U7921 ( .A1(n6151), .A2(n6150), .ZN(n7675) );
  NAND2_X1 U7922 ( .A1(n6723), .A2(n7891), .ZN(n6153) );
  AOI22_X1 U7923 ( .A1(n6176), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6175), .B2(
        n10322), .ZN(n6152) );
  INV_X1 U7924 ( .A(n6154), .ZN(n6168) );
  NAND2_X1 U7925 ( .A1(n6155), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6156) );
  NAND2_X1 U7926 ( .A1(n6168), .A2(n6156), .ZN(n8175) );
  NAND2_X1 U7927 ( .A1(n6266), .A2(n8175), .ZN(n6160) );
  OR2_X1 U7928 ( .A1(n7900), .A2(n7680), .ZN(n6159) );
  OR2_X1 U7929 ( .A1(n7902), .A2(n5880), .ZN(n6158) );
  INV_X1 U7930 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n7677) );
  OR2_X1 U7931 ( .A1(n6050), .A2(n7677), .ZN(n6157) );
  NAND2_X1 U7932 ( .A1(n8181), .A2(n8187), .ZN(n8038) );
  INV_X1 U7933 ( .A(n8037), .ZN(n6161) );
  NAND2_X1 U7934 ( .A1(n7675), .A2(n6161), .ZN(n6163) );
  INV_X1 U7935 ( .A(n8187), .ZN(n8274) );
  NAND2_X1 U7936 ( .A1(n8181), .A2(n8274), .ZN(n6162) );
  NAND2_X1 U7937 ( .A1(n6163), .A2(n6162), .ZN(n7735) );
  NAND2_X1 U7938 ( .A1(n6779), .A2(n7891), .ZN(n6165) );
  AOI22_X1 U7939 ( .A1(n6176), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6175), .B2(
        n10341), .ZN(n6164) );
  INV_X1 U7940 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8964) );
  OR2_X1 U7941 ( .A1(n7900), .A2(n8964), .ZN(n6167) );
  INV_X1 U7942 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8788) );
  OR2_X1 U7943 ( .A1(n6050), .A2(n8788), .ZN(n6166) );
  AND2_X1 U7944 ( .A1(n6167), .A2(n6166), .ZN(n6172) );
  NAND2_X1 U7945 ( .A1(n6168), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6169) );
  NAND2_X1 U7946 ( .A1(n6179), .A2(n6169), .ZN(n8184) );
  NAND2_X1 U7947 ( .A1(n8184), .A2(n6266), .ZN(n6171) );
  INV_X1 U7948 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n7738) );
  OR2_X1 U7949 ( .A1(n7902), .A2(n7738), .ZN(n6170) );
  OR2_X1 U7950 ( .A1(n8491), .A2(n8235), .ZN(n8050) );
  NAND2_X1 U7951 ( .A1(n8491), .A2(n8235), .ZN(n8051) );
  NAND2_X1 U7952 ( .A1(n8050), .A2(n8051), .ZN(n8043) );
  NAND2_X1 U7953 ( .A1(n7735), .A2(n8043), .ZN(n6174) );
  NAND2_X1 U7954 ( .A1(n8491), .A2(n8428), .ZN(n6173) );
  NAND2_X1 U7955 ( .A1(n6174), .A2(n6173), .ZN(n8425) );
  NAND2_X1 U7956 ( .A1(n7051), .A2(n7891), .ZN(n6178) );
  AOI22_X1 U7957 ( .A1(n6176), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6175), .B2(
        n9950), .ZN(n6177) );
  NAND2_X1 U7958 ( .A1(n6179), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6180) );
  NAND2_X1 U7959 ( .A1(n6181), .A2(n6180), .ZN(n8431) );
  NAND2_X1 U7960 ( .A1(n8431), .A2(n6266), .ZN(n6184) );
  AOI22_X1 U7961 ( .A1(n6315), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n6316), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U7962 ( .A1(n6314), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6182) );
  AND2_X1 U7963 ( .A1(n8435), .A2(n8412), .ZN(n6185) );
  OR2_X1 U7964 ( .A1(n8435), .A2(n8412), .ZN(n6186) );
  NAND2_X1 U7965 ( .A1(n8476), .A2(n8202), .ZN(n8055) );
  NOR2_X1 U7966 ( .A1(n7893), .A2(n8894), .ZN(n6188) );
  AOI21_X1 U7967 ( .B1(n7223), .B2(n7891), .A(n6188), .ZN(n7837) );
  INV_X1 U7968 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n6189) );
  INV_X1 U7969 ( .A(n6202), .ZN(n6203) );
  NAND2_X1 U7970 ( .A1(n6191), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6192) );
  NAND2_X1 U7971 ( .A1(n6203), .A2(n6192), .ZN(n8403) );
  NAND2_X1 U7972 ( .A1(n8403), .A2(n6266), .ZN(n6197) );
  INV_X1 U7973 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8532) );
  NAND2_X1 U7974 ( .A1(n6316), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U7975 ( .A1(n6315), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6193) );
  OAI211_X1 U7976 ( .C1(n6050), .C2(n8532), .A(n6194), .B(n6193), .ZN(n6195)
         );
  INV_X1 U7977 ( .A(n6195), .ZN(n6196) );
  NAND2_X1 U7978 ( .A1(n6197), .A2(n6196), .ZN(n8413) );
  INV_X1 U7979 ( .A(n7837), .ZN(n8534) );
  NAND2_X1 U7980 ( .A1(n8534), .A2(n8390), .ZN(n8380) );
  NAND2_X1 U7981 ( .A1(n4567), .A2(n8380), .ZN(n8400) );
  NAND2_X1 U7982 ( .A1(n7367), .A2(n7891), .ZN(n6200) );
  OR2_X1 U7983 ( .A1(n7893), .A2(n7384), .ZN(n6199) );
  INV_X1 U7984 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6201) );
  NAND2_X1 U7985 ( .A1(n6203), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6204) );
  NAND2_X1 U7986 ( .A1(n6211), .A2(n6204), .ZN(n8392) );
  INV_X1 U7987 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8528) );
  NAND2_X1 U7988 ( .A1(n6316), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6206) );
  NAND2_X1 U7989 ( .A1(n6315), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6205) );
  OAI211_X1 U7990 ( .C1(n6050), .C2(n8528), .A(n6206), .B(n6205), .ZN(n6207)
         );
  NAND2_X1 U7991 ( .A1(n8469), .A2(n8222), .ZN(n8066) );
  NAND2_X1 U7992 ( .A1(n7492), .A2(n7891), .ZN(n6210) );
  OR2_X1 U7993 ( .A1(n7893), .A2(n9038), .ZN(n6209) );
  NAND2_X1 U7994 ( .A1(n6211), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U7995 ( .A1(n6221), .A2(n6212), .ZN(n8371) );
  NAND2_X1 U7996 ( .A1(n8371), .A2(n6266), .ZN(n6218) );
  INV_X1 U7997 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n6215) );
  NAND2_X1 U7998 ( .A1(n6316), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6214) );
  NAND2_X1 U7999 ( .A1(n6315), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6213) );
  OAI211_X1 U8000 ( .C1(n6050), .C2(n6215), .A(n6214), .B(n6213), .ZN(n6216)
         );
  INV_X1 U8001 ( .A(n6216), .ZN(n6217) );
  NAND2_X1 U8002 ( .A1(n7575), .A2(n7891), .ZN(n6220) );
  OR2_X1 U8003 ( .A1(n7893), .A2(n7573), .ZN(n6219) );
  NAND2_X1 U8004 ( .A1(n6221), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6222) );
  NAND2_X1 U8005 ( .A1(n6231), .A2(n6222), .ZN(n8362) );
  NAND2_X1 U8006 ( .A1(n8362), .A2(n6266), .ZN(n6227) );
  INV_X1 U8007 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8523) );
  NAND2_X1 U8008 ( .A1(n6315), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6224) );
  NAND2_X1 U8009 ( .A1(n6316), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6223) );
  OAI211_X1 U8010 ( .C1(n6050), .C2(n8523), .A(n6224), .B(n6223), .ZN(n6225)
         );
  INV_X1 U8011 ( .A(n6225), .ZN(n6226) );
  NOR2_X1 U8012 ( .A1(n8460), .A2(n8369), .ZN(n6228) );
  NAND2_X1 U8013 ( .A1(n7619), .A2(n7891), .ZN(n6230) );
  OR2_X1 U8014 ( .A1(n7893), .A2(n7673), .ZN(n6229) );
  INV_X1 U8015 ( .A(n6244), .ZN(n6245) );
  NAND2_X1 U8016 ( .A1(n6231), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U8017 ( .A1(n6245), .A2(n6232), .ZN(n8354) );
  NAND2_X1 U8018 ( .A1(n8354), .A2(n6266), .ZN(n6237) );
  INV_X1 U8019 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8928) );
  NAND2_X1 U8020 ( .A1(n6315), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6234) );
  NAND2_X1 U8021 ( .A1(n6316), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6233) );
  OAI211_X1 U8022 ( .C1(n6050), .C2(n8928), .A(n6234), .B(n6233), .ZN(n6235)
         );
  INV_X1 U8023 ( .A(n6235), .ZN(n6236) );
  INV_X1 U8024 ( .A(n8361), .ZN(n8338) );
  INV_X1 U8025 ( .A(n8518), .ZN(n8352) );
  NAND2_X1 U8026 ( .A1(n7742), .A2(n7891), .ZN(n6242) );
  OR2_X1 U8027 ( .A1(n7893), .A2(n7746), .ZN(n6241) );
  INV_X1 U8028 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6243) );
  INV_X1 U8029 ( .A(n6256), .ZN(n6247) );
  NAND2_X1 U8030 ( .A1(n6245), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6246) );
  NAND2_X1 U8031 ( .A1(n6247), .A2(n6246), .ZN(n8340) );
  NAND2_X1 U8032 ( .A1(n8340), .A2(n6266), .ZN(n6252) );
  INV_X1 U8033 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8916) );
  NAND2_X1 U8034 ( .A1(n6316), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6249) );
  INV_X1 U8035 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8886) );
  OR2_X1 U8036 ( .A1(n7900), .A2(n8886), .ZN(n6248) );
  OAI211_X1 U8037 ( .C1(n6050), .C2(n8916), .A(n6249), .B(n6248), .ZN(n6250)
         );
  INV_X1 U8038 ( .A(n6250), .ZN(n6251) );
  NAND2_X1 U8039 ( .A1(n8513), .A2(n8326), .ZN(n8091) );
  NAND2_X1 U8040 ( .A1(n7775), .A2(n7891), .ZN(n6254) );
  OR2_X1 U8041 ( .A1(n7893), .A2(n7777), .ZN(n6253) );
  INV_X1 U8042 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6255) );
  NOR2_X1 U8043 ( .A1(n6256), .A2(n6255), .ZN(n6257) );
  INV_X1 U8044 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8329) );
  NAND2_X1 U8045 ( .A1(n6315), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6259) );
  NAND2_X1 U8046 ( .A1(n6314), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6258) );
  OAI211_X1 U8047 ( .C1(n7902), .C2(n8329), .A(n6259), .B(n6258), .ZN(n6260)
         );
  INV_X1 U8048 ( .A(n8316), .ZN(n8337) );
  NOR2_X1 U8049 ( .A1(n8331), .A2(n8337), .ZN(n6261) );
  NAND2_X1 U8050 ( .A1(n7802), .A2(n7891), .ZN(n6263) );
  OR2_X1 U8051 ( .A1(n7893), .A2(n9021), .ZN(n6262) );
  OR2_X1 U8052 ( .A1(n6264), .A2(n9044), .ZN(n6265) );
  NAND2_X1 U8053 ( .A1(n9044), .A2(n6264), .ZN(n6277) );
  NAND2_X1 U8054 ( .A1(n6265), .A2(n6277), .ZN(n8317) );
  NAND2_X1 U8055 ( .A1(n8317), .A2(n6266), .ZN(n6271) );
  NAND2_X1 U8056 ( .A1(n6314), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6268) );
  NAND2_X1 U8057 ( .A1(n6315), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6267) );
  OAI211_X1 U8058 ( .C1(n7902), .C2(n9095), .A(n6268), .B(n6267), .ZN(n6269)
         );
  INV_X1 U8059 ( .A(n6269), .ZN(n6270) );
  NAND2_X1 U8060 ( .A1(n8448), .A2(n8327), .ZN(n8095) );
  NAND2_X1 U8061 ( .A1(n8094), .A2(n8095), .ZN(n8312) );
  NAND2_X1 U8062 ( .A1(n7817), .A2(n7891), .ZN(n6274) );
  OR2_X1 U8063 ( .A1(n7893), .A2(n6272), .ZN(n6273) );
  NAND2_X1 U8064 ( .A1(n6314), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6282) );
  INV_X1 U8065 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6366) );
  OR2_X1 U8066 ( .A1(n7900), .A2(n6366), .ZN(n6281) );
  INV_X1 U8067 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6276) );
  INV_X1 U8068 ( .A(n6277), .ZN(n6275) );
  NAND2_X1 U8069 ( .A1(n6276), .A2(n6275), .ZN(n7808) );
  NAND2_X1 U8070 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(n6277), .ZN(n6278) );
  OR2_X1 U8071 ( .A1(n6285), .A2(n8300), .ZN(n6280) );
  INV_X1 U8072 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8301) );
  OR2_X1 U8073 ( .A1(n7902), .A2(n8301), .ZN(n6279) );
  NAND4_X1 U8074 ( .A1(n6282), .A2(n6281), .A3(n6280), .A4(n6279), .ZN(n8271)
         );
  XNOR2_X1 U8075 ( .A(n8303), .B(n8271), .ZN(n7936) );
  INV_X1 U8076 ( .A(n8303), .ZN(n8114) );
  INV_X1 U8077 ( .A(n8271), .ZN(n8315) );
  NAND2_X1 U8078 ( .A1(n7799), .A2(n7891), .ZN(n6284) );
  OR2_X1 U8079 ( .A1(n7893), .A2(n8552), .ZN(n6283) );
  INV_X1 U8080 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8906) );
  OR2_X1 U8081 ( .A1(n7900), .A2(n8906), .ZN(n6289) );
  INV_X1 U8082 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n7810) );
  OR2_X1 U8083 ( .A1(n7902), .A2(n7810), .ZN(n6288) );
  INV_X1 U8084 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6286) );
  OR2_X1 U8085 ( .A1(n6050), .A2(n6286), .ZN(n6287) );
  NOR2_X1 U8086 ( .A1(n7815), .A2(n7861), .ZN(n7897) );
  INV_X1 U8087 ( .A(n7897), .ZN(n8111) );
  NAND2_X1 U8088 ( .A1(n7815), .A2(n7861), .ZN(n7890) );
  NAND2_X1 U8089 ( .A1(n8111), .A2(n7890), .ZN(n8100) );
  XNOR2_X1 U8090 ( .A(n6290), .B(n8100), .ZN(n6326) );
  NAND2_X1 U8091 ( .A1(n8128), .A2(n8124), .ZN(n6375) );
  NAND2_X1 U8092 ( .A1(n6291), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6292) );
  MUX2_X1 U8093 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6292), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n6294) );
  NAND2_X1 U8094 ( .A1(n7957), .A2(n8118), .ZN(n6295) );
  NAND2_X1 U8095 ( .A1(n6942), .A2(n6658), .ZN(n7975) );
  NAND2_X1 U8096 ( .A1(n6588), .A2(n7975), .ZN(n7016) );
  NAND2_X1 U8097 ( .A1(n6692), .A2(n10390), .ZN(n7983) );
  INV_X1 U8098 ( .A(n6692), .ZN(n8288) );
  NAND2_X1 U8099 ( .A1(n8288), .A2(n7017), .ZN(n7992) );
  NAND2_X1 U8100 ( .A1(n7016), .A2(n7911), .ZN(n6298) );
  NAND2_X1 U8101 ( .A1(n6298), .A2(n7983), .ZN(n6576) );
  NAND2_X1 U8102 ( .A1(n6754), .A2(n6694), .ZN(n7993) );
  NAND2_X1 U8103 ( .A1(n8286), .A2(n6736), .ZN(n7984) );
  NAND2_X1 U8104 ( .A1(n6043), .A2(n10394), .ZN(n7994) );
  NAND2_X1 U8105 ( .A1(n7063), .A2(n10398), .ZN(n7997) );
  AND2_X1 U8106 ( .A1(n7994), .A2(n7997), .ZN(n7987) );
  NAND2_X1 U8107 ( .A1(n7008), .A2(n8285), .ZN(n7988) );
  NAND2_X1 U8108 ( .A1(n6299), .A2(n7988), .ZN(n7096) );
  OR2_X1 U8109 ( .A1(n7058), .A2(n10406), .ZN(n7944) );
  NAND2_X1 U8110 ( .A1(n10406), .A2(n7058), .ZN(n7948) );
  NAND2_X1 U8111 ( .A1(n7096), .A2(n8001), .ZN(n7098) );
  OR2_X1 U8112 ( .A1(n10416), .A2(n7426), .ZN(n7946) );
  AND2_X1 U8113 ( .A1(n7114), .A2(n8282), .ZN(n7190) );
  INV_X1 U8114 ( .A(n7190), .ZN(n7945) );
  NAND2_X1 U8115 ( .A1(n7946), .A2(n7945), .ZN(n7953) );
  AND2_X1 U8116 ( .A1(n10419), .A2(n8280), .ZN(n7142) );
  OR2_X1 U8117 ( .A1(n7953), .A2(n7142), .ZN(n7176) );
  INV_X1 U8118 ( .A(n8010), .ZN(n8005) );
  NAND2_X1 U8119 ( .A1(n7432), .A2(n7457), .ZN(n7950) );
  AND2_X1 U8120 ( .A1(n8006), .A2(n7950), .ZN(n8008) );
  INV_X1 U8121 ( .A(n7946), .ZN(n6300) );
  NAND2_X1 U8122 ( .A1(n10416), .A2(n7426), .ZN(n7951) );
  NAND2_X1 U8123 ( .A1(n10407), .A2(n7152), .ZN(n7949) );
  OR2_X1 U8124 ( .A1(n7142), .A2(n7140), .ZN(n7177) );
  OR2_X1 U8125 ( .A1(n7568), .A2(n7749), .ZN(n8013) );
  NAND2_X1 U8126 ( .A1(n7568), .A2(n7749), .ZN(n8012) );
  NAND2_X1 U8127 ( .A1(n7252), .A2(n8013), .ZN(n7417) );
  NAND2_X1 U8128 ( .A1(n8217), .A2(n8020), .ZN(n6301) );
  OR2_X1 U8129 ( .A1(n8217), .A2(n8020), .ZN(n6302) );
  NOR2_X1 U8130 ( .A1(n7751), .A2(n8259), .ZN(n8030) );
  INV_X1 U8131 ( .A(n8030), .ZN(n6303) );
  NAND2_X1 U8132 ( .A1(n7751), .A2(n8259), .ZN(n8029) );
  AND2_X1 U8133 ( .A1(n8250), .A2(n8179), .ZN(n7527) );
  OR2_X1 U8134 ( .A1(n8250), .A2(n8179), .ZN(n8036) );
  NAND2_X1 U8135 ( .A1(n7674), .A2(n8038), .ZN(n6305) );
  NAND2_X1 U8136 ( .A1(n6305), .A2(n8041), .ZN(n7732) );
  NAND2_X1 U8137 ( .A1(n8435), .A2(n8154), .ZN(n7929) );
  NAND2_X1 U8138 ( .A1(n7928), .A2(n7929), .ZN(n8437) );
  AND2_X1 U8139 ( .A1(n8066), .A2(n8380), .ZN(n7939) );
  INV_X1 U8140 ( .A(n8273), .ZN(n8388) );
  OR2_X1 U8141 ( .A1(n8463), .A2(n8388), .ZN(n8071) );
  AND2_X1 U8142 ( .A1(n7845), .A2(n8369), .ZN(n7909) );
  NAND2_X1 U8143 ( .A1(n8460), .A2(n8221), .ZN(n8078) );
  NAND2_X1 U8144 ( .A1(n8334), .A2(n8091), .ZN(n6308) );
  NOR2_X1 U8145 ( .A1(n8331), .A2(n8316), .ZN(n7907) );
  INV_X1 U8146 ( .A(n8312), .ZN(n6309) );
  NAND2_X1 U8147 ( .A1(n8331), .A2(n8316), .ZN(n8307) );
  AND2_X1 U8148 ( .A1(n6309), .A2(n8307), .ZN(n6310) );
  OR2_X1 U8149 ( .A1(n8303), .A2(n8315), .ZN(n6311) );
  INV_X1 U8150 ( .A(n8100), .ZN(n6312) );
  INV_X1 U8151 ( .A(n8118), .ZN(n7261) );
  INV_X1 U8152 ( .A(n8128), .ZN(n7493) );
  AOI21_X1 U8153 ( .B1(n7493), .B2(n8118), .A(n8124), .ZN(n6313) );
  NAND3_X1 U8154 ( .A1(n6675), .A2(n6313), .A3(n10418), .ZN(n7200) );
  NOR2_X1 U8155 ( .A1(n7812), .A2(n7200), .ZN(n6325) );
  NAND2_X1 U8156 ( .A1(n6314), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6319) );
  NAND2_X1 U8157 ( .A1(n6315), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6318) );
  NAND2_X1 U8158 ( .A1(n6316), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6317) );
  AND4_X1 U8159 ( .A1(n7906), .A2(n6319), .A3(n6318), .A4(n6317), .ZN(n7889)
         );
  INV_X1 U8160 ( .A(n7889), .ZN(n8269) );
  OR2_X1 U8161 ( .A1(n5886), .A2(n5948), .ZN(n6320) );
  NAND2_X1 U8162 ( .A1(n6322), .A2(P2_B_REG_SCAN_IN), .ZN(n6323) );
  AND2_X1 U8163 ( .A1(n6321), .A2(n6323), .ZN(n8291) );
  AOI22_X1 U8164 ( .A1(n8269), .A2(n8291), .B1(n8427), .B2(n8271), .ZN(n6324)
         );
  INV_X1 U8165 ( .A(n7812), .ZN(n6329) );
  INV_X1 U8166 ( .A(n6714), .ZN(n6327) );
  NAND2_X1 U8167 ( .A1(n6331), .A2(n7776), .ZN(n6648) );
  NAND2_X1 U8168 ( .A1(n6332), .A2(n7776), .ZN(n6334) );
  NAND2_X1 U8169 ( .A1(n8118), .A2(n7138), .ZN(n6336) );
  NAND2_X1 U8170 ( .A1(n7963), .A2(n6336), .ZN(n6337) );
  NAND2_X1 U8171 ( .A1(n8128), .A2(n6337), .ZN(n6664) );
  NAND2_X1 U8172 ( .A1(n6667), .A2(n6664), .ZN(n6338) );
  AND2_X1 U8173 ( .A1(n6373), .A2(n6338), .ZN(n6355) );
  INV_X1 U8174 ( .A(n6452), .ZN(n6349) );
  NOR4_X1 U8175 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6347) );
  INV_X1 U8176 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n8930) );
  INV_X1 U8177 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n8961) );
  INV_X1 U8178 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n9050) );
  INV_X1 U8179 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n9094) );
  NAND4_X1 U8180 ( .A1(n8930), .A2(n8961), .A3(n9050), .A4(n9094), .ZN(n6344)
         );
  NOR4_X1 U8181 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6342) );
  NOR4_X1 U8182 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6341) );
  NOR4_X1 U8183 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6340) );
  NOR4_X1 U8184 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6339) );
  NAND4_X1 U8185 ( .A1(n6342), .A2(n6341), .A3(n6340), .A4(n6339), .ZN(n6343)
         );
  NOR4_X1 U8186 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        n6344), .A4(n6343), .ZN(n6346) );
  NOR4_X1 U8187 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6345) );
  NAND3_X1 U8188 ( .A1(n6347), .A2(n6346), .A3(n6345), .ZN(n6348) );
  OR2_X1 U8189 ( .A1(n8106), .A2(n6649), .ZN(n6350) );
  AND2_X1 U8190 ( .A1(n6374), .A2(n6350), .ZN(n6620) );
  NAND2_X1 U8191 ( .A1(n6620), .A2(n6627), .ZN(n6351) );
  NAND2_X1 U8192 ( .A1(n6328), .A2(n7963), .ZN(n6603) );
  INV_X1 U8193 ( .A(n6603), .ZN(n6352) );
  INV_X1 U8194 ( .A(n6664), .ZN(n6666) );
  NAND2_X1 U8195 ( .A1(n6665), .A2(n6666), .ZN(n6353) );
  INV_X1 U8196 ( .A(n7815), .ZN(n6390) );
  NAND2_X1 U8197 ( .A1(n10446), .A2(n10429), .ZN(n8451) );
  NAND2_X1 U8198 ( .A1(n10444), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6356) );
  NAND2_X1 U8199 ( .A1(n6359), .A2(n6358), .ZN(P2_U3488) );
  XNOR2_X1 U8200 ( .A(n6360), .B(n7936), .ZN(n6364) );
  MUX2_X1 U8201 ( .A(n6366), .B(n6381), .S(n10446), .Z(n6372) );
  OAI21_X1 U8202 ( .B1(n6368), .B2(n7936), .A(n6367), .ZN(n8306) );
  NAND2_X1 U8203 ( .A1(n6370), .A2(n6369), .ZN(n6371) );
  NAND2_X1 U8204 ( .A1(n6372), .A2(n6371), .ZN(P2_U3487) );
  INV_X1 U8205 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6382) );
  INV_X1 U8206 ( .A(n6623), .ZN(n6451) );
  NAND2_X1 U8207 ( .A1(n6615), .A2(n6451), .ZN(n6606) );
  NAND2_X1 U8208 ( .A1(n7963), .A2(n8118), .ZN(n6376) );
  OR2_X1 U8209 ( .A1(n6376), .A2(n6375), .ZN(n6607) );
  AND2_X1 U8210 ( .A1(n6607), .A2(n6675), .ZN(n6377) );
  OR2_X1 U8211 ( .A1(n6606), .A2(n6377), .ZN(n6380) );
  NAND2_X1 U8212 ( .A1(n6667), .A2(n6665), .ZN(n6670) );
  NAND3_X1 U8213 ( .A1(n6607), .A2(n8106), .A3(n10418), .ZN(n6605) );
  NAND2_X1 U8214 ( .A1(n6605), .A2(n10370), .ZN(n6616) );
  NAND2_X1 U8215 ( .A1(n6610), .A2(n6616), .ZN(n6379) );
  MUX2_X1 U8216 ( .A(n6382), .B(n6381), .S(n10430), .Z(n6384) );
  INV_X1 U8217 ( .A(n10408), .ZN(n10424) );
  NAND2_X1 U8218 ( .A1(n6370), .A2(n7418), .ZN(n6383) );
  NAND2_X1 U8219 ( .A1(n6384), .A2(n6383), .ZN(P2_U3455) );
  INV_X1 U8220 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6386) );
  MUX2_X1 U8221 ( .A(n6386), .B(n6385), .S(n10175), .Z(n6388) );
  NAND2_X1 U8222 ( .A1(n6388), .A2(n5082), .ZN(P1_U3521) );
  OR2_X1 U8223 ( .A1(n10430), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6389) );
  NAND2_X1 U8224 ( .A1(n6391), .A2(n5081), .ZN(P2_U3456) );
  NAND2_X1 U8225 ( .A1(n7576), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6392) );
  INV_X1 U8226 ( .A(n6435), .ZN(n6800) );
  INV_X1 U8227 ( .A(n6426), .ZN(n9525) );
  INV_X1 U8228 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6393) );
  MUX2_X1 U8229 ( .A(n6393), .B(P1_REG2_REG_1__SCAN_IN), .S(n6422), .Z(n6726)
         );
  NAND2_X1 U8230 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10002) );
  NOR2_X1 U8231 ( .A1(n6726), .A2(n10002), .ZN(n6725) );
  AOI21_X1 U8232 ( .B1(n6422), .B2(P1_REG2_REG_1__SCAN_IN), .A(n6725), .ZN(
        n9998) );
  NAND2_X1 U8233 ( .A1(n10001), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6394) );
  OAI21_X1 U8234 ( .B1(n10001), .B2(P1_REG2_REG_2__SCAN_IN), .A(n6394), .ZN(
        n9997) );
  XOR2_X1 U8235 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6426), .Z(n9519) );
  NAND2_X1 U8236 ( .A1(n10024), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6395) );
  OAI21_X1 U8237 ( .B1(n10024), .B2(P1_REG2_REG_4__SCAN_IN), .A(n6395), .ZN(
        n10020) );
  NOR2_X1 U8238 ( .A1(n10021), .A2(n10020), .ZN(n10019) );
  XOR2_X1 U8239 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n6435), .Z(n6795) );
  OR2_X1 U8240 ( .A1(n6825), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6397) );
  NAND2_X1 U8241 ( .A1(n6825), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6396) );
  NAND2_X1 U8242 ( .A1(n6397), .A2(n6396), .ZN(n6820) );
  AOI21_X1 U8243 ( .B1(n6825), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6819), .ZN(
        n6403) );
  MUX2_X1 U8244 ( .A(n4935), .B(P1_REG2_REG_7__SCAN_IN), .S(n6554), .Z(n6398)
         );
  INV_X1 U8245 ( .A(n6398), .ZN(n6402) );
  NOR2_X1 U8246 ( .A1(n6403), .A2(n6402), .ZN(n6555) );
  INV_X1 U8247 ( .A(n7576), .ZN(n6399) );
  OAI21_X1 U8248 ( .B1(n6530), .B2(n6399), .A(P1_STATE_REG_SCAN_IN), .ZN(n6414) );
  NAND2_X1 U8249 ( .A1(n9463), .A2(n7576), .ZN(n6400) );
  NAND2_X1 U8250 ( .A1(n5151), .A2(n6400), .ZN(n6413) );
  OR2_X1 U8251 ( .A1(n6414), .A2(n6413), .ZN(n9991) );
  INV_X1 U8252 ( .A(n9991), .ZN(n6401) );
  NAND2_X1 U8253 ( .A1(n6401), .A2(n9987), .ZN(n9595) );
  NOR2_X1 U8254 ( .A1(n9595), .A2(n5454), .ZN(n9593) );
  AOI211_X1 U8255 ( .C1(n6403), .C2(n6402), .A(n6555), .B(n10018), .ZN(n6421)
         );
  INV_X1 U8256 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10176) );
  XNOR2_X1 U8257 ( .A(n6422), .B(n10176), .ZN(n6729) );
  AND2_X1 U8258 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6728) );
  NAND2_X1 U8259 ( .A1(n6729), .A2(n6728), .ZN(n6727) );
  NAND2_X1 U8260 ( .A1(n6422), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6404) );
  AND2_X1 U8261 ( .A1(n6727), .A2(n6404), .ZN(n9995) );
  XNOR2_X1 U8262 ( .A(n6426), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9528) );
  NAND2_X1 U8263 ( .A1(n9527), .A2(n9528), .ZN(n9526) );
  INV_X1 U8264 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6405) );
  OR2_X1 U8265 ( .A1(n6426), .A2(n6405), .ZN(n6406) );
  NAND2_X1 U8266 ( .A1(n9526), .A2(n6406), .ZN(n10013) );
  OR2_X1 U8267 ( .A1(n10024), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6408) );
  NAND2_X1 U8268 ( .A1(n10024), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6407) );
  AND2_X1 U8269 ( .A1(n6408), .A2(n6407), .ZN(n10014) );
  XOR2_X1 U8270 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6435), .Z(n6798) );
  AOI21_X1 U8271 ( .B1(n6800), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6797), .ZN(
        n6824) );
  INV_X1 U8272 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6409) );
  MUX2_X1 U8273 ( .A(n6409), .B(P1_REG1_REG_6__SCAN_IN), .S(n6825), .Z(n6823)
         );
  NOR2_X1 U8274 ( .A1(n6824), .A2(n6823), .ZN(n6822) );
  AOI21_X1 U8275 ( .B1(n6825), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6822), .ZN(
        n6412) );
  INV_X1 U8276 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6410) );
  MUX2_X1 U8277 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n6410), .S(n6554), .Z(n6411)
         );
  NOR2_X1 U8278 ( .A1(n6412), .A2(n6411), .ZN(n6559) );
  AOI211_X1 U8279 ( .C1(n6412), .C2(n6411), .A(n6559), .B(n9993), .ZN(n6420)
         );
  NOR2_X2 U8280 ( .A1(n9991), .A2(n10005), .ZN(n10025) );
  INV_X1 U8281 ( .A(n10025), .ZN(n7132) );
  NOR2_X1 U8282 ( .A1(n7132), .A2(n6554), .ZN(n6419) );
  INV_X1 U8283 ( .A(n6413), .ZN(n6415) );
  INV_X1 U8284 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6417) );
  NAND2_X1 U8285 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n6416) );
  OAI21_X1 U8286 ( .B1(n9601), .B2(n6417), .A(n6416), .ZN(n6418) );
  OR4_X1 U8287 ( .A1(n6421), .A2(n6420), .A3(n6419), .A4(n6418), .ZN(P1_U3250)
         );
  INV_X1 U8288 ( .A(n6422), .ZN(n6732) );
  OAI222_X1 U8289 ( .A1(n7819), .A2(n6423), .B1(n4496), .B2(n6444), .C1(
        P1_U3086), .C2(n6732), .ZN(P1_U3354) );
  OAI222_X1 U8290 ( .A1(n7819), .A2(n6425), .B1(n4496), .B2(n6430), .C1(
        P1_U3086), .C2(n6424), .ZN(P1_U3353) );
  OAI222_X1 U8291 ( .A1(n7819), .A2(n6427), .B1(n4496), .B2(n6431), .C1(
        P1_U3086), .C2(n6426), .ZN(P1_U3352) );
  OAI222_X1 U8292 ( .A1(n7819), .A2(n6429), .B1(n4496), .B2(n6433), .C1(
        P1_U3086), .C2(n6428), .ZN(P1_U3351) );
  NOR2_X1 U8293 ( .A1(n4835), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8560) );
  INV_X2 U8294 ( .A(n8560), .ZN(n8551) );
  NAND2_X1 U8295 ( .A1(n4835), .A2(P2_U3151), .ZN(n8562) );
  OAI222_X1 U8296 ( .A1(n8551), .A2(n4589), .B1(n8562), .B2(n6430), .C1(
        P2_U3151), .C2(n7036), .ZN(P2_U3293) );
  OAI222_X1 U8297 ( .A1(n8551), .A2(n6432), .B1(n8562), .B2(n6431), .C1(
        P2_U3151), .C2(n6999), .ZN(P2_U3292) );
  OAI222_X1 U8298 ( .A1(n8551), .A2(n6434), .B1(n8562), .B2(n6433), .C1(
        P2_U3151), .C2(n6984), .ZN(P2_U3291) );
  OAI222_X1 U8299 ( .A1(n7819), .A2(n6436), .B1(n4496), .B2(n6438), .C1(
        P1_U3086), .C2(n6435), .ZN(P1_U3350) );
  OAI222_X1 U8300 ( .A1(n8551), .A2(n6439), .B1(n8562), .B2(n6438), .C1(
        P2_U3151), .C2(n6437), .ZN(P2_U3290) );
  OAI222_X1 U8301 ( .A1(n7819), .A2(n6441), .B1(n4496), .B2(n6443), .C1(
        P1_U3086), .C2(n6440), .ZN(P1_U3349) );
  INV_X1 U8302 ( .A(n8562), .ZN(n7571) );
  INV_X1 U8303 ( .A(n7571), .ZN(n8555) );
  AOI22_X1 U8304 ( .A1(n6869), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n8560), .ZN(n6442) );
  OAI21_X1 U8305 ( .B1(n6443), .B2(n8555), .A(n6442), .ZN(P2_U3289) );
  OAI222_X1 U8306 ( .A1(n8551), .A2(n4836), .B1(n8555), .B2(n6444), .C1(
        P2_U3151), .C2(n10193), .ZN(P2_U3294) );
  INV_X1 U8307 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6445) );
  OAI222_X1 U8308 ( .A1(n8551), .A2(n6445), .B1(n8562), .B2(n6446), .C1(
        P2_U3151), .C2(n7084), .ZN(P2_U3288) );
  OAI222_X1 U8309 ( .A1(n7819), .A2(n6447), .B1(n4496), .B2(n6446), .C1(
        P1_U3086), .C2(n6554), .ZN(P1_U3348) );
  OAI222_X1 U8310 ( .A1(n8551), .A2(n9062), .B1(n8562), .B2(n6449), .C1(
        P2_U3151), .C2(n4873), .ZN(P2_U3287) );
  OAI222_X1 U8311 ( .A1(n7819), .A2(n6450), .B1(n4496), .B2(n6449), .C1(
        P1_U3086), .C2(n6448), .ZN(P1_U3347) );
  INV_X1 U8312 ( .A(n6648), .ZN(n6453) );
  AOI22_X1 U8313 ( .A1(n6467), .A2(n4973), .B1(n6627), .B2(n6453), .ZN(
        P2_U3376) );
  INV_X1 U8314 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6455) );
  AND2_X1 U8315 ( .A1(n6627), .A2(n7776), .ZN(n6454) );
  AOI22_X1 U8316 ( .A1(n6467), .A2(n6455), .B1(n6454), .B2(n6332), .ZN(
        P2_U3377) );
  OAI222_X1 U8317 ( .A1(n8551), .A2(n6457), .B1(n8562), .B2(n6458), .C1(n6456), 
        .C2(P2_U3151), .ZN(P2_U3286) );
  OAI222_X1 U8318 ( .A1(n7819), .A2(n6459), .B1(n4496), .B2(n6458), .C1(n6567), 
        .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U8319 ( .A(n6460), .ZN(n6463) );
  INV_X1 U8320 ( .A(n7819), .ZN(n9934) );
  AOI22_X1 U8321 ( .A1(n7071), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9934), .ZN(n6461) );
  OAI21_X1 U8322 ( .B1(n6463), .B2(n4496), .A(n6461), .ZN(P1_U3345) );
  INV_X1 U8323 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6464) );
  OAI222_X1 U8324 ( .A1(n8551), .A2(n6464), .B1(n8555), .B2(n6463), .C1(n6462), 
        .C2(P2_U3151), .ZN(P2_U3285) );
  AOI21_X1 U8325 ( .B1(P1_D_REG_0__SCAN_IN), .B2(n6850), .A(n6465), .ZN(n6466)
         );
  INV_X1 U8326 ( .A(n6466), .ZN(P1_U3439) );
  INV_X1 U8327 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n6468) );
  NOR2_X1 U8328 ( .A1(n6501), .A2(n6468), .ZN(P2_U3258) );
  NOR2_X1 U8329 ( .A1(n6501), .A2(n8930), .ZN(P2_U3261) );
  INV_X1 U8330 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n6469) );
  NOR2_X1 U8331 ( .A1(n6501), .A2(n6469), .ZN(P2_U3262) );
  INV_X1 U8332 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n6470) );
  NOR2_X1 U8333 ( .A1(n6501), .A2(n6470), .ZN(P2_U3252) );
  INV_X1 U8334 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n6471) );
  NOR2_X1 U8335 ( .A1(n6501), .A2(n6471), .ZN(P2_U3253) );
  INV_X1 U8336 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n6472) );
  NOR2_X1 U8337 ( .A1(n6501), .A2(n6472), .ZN(P2_U3249) );
  INV_X1 U8338 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n6473) );
  NOR2_X1 U8339 ( .A1(n6501), .A2(n6473), .ZN(P2_U3259) );
  INV_X1 U8340 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n6474) );
  NOR2_X1 U8341 ( .A1(n6501), .A2(n6474), .ZN(P2_U3260) );
  INV_X1 U8342 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n6475) );
  NOR2_X1 U8343 ( .A1(n6501), .A2(n6475), .ZN(P2_U3246) );
  INV_X1 U8344 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n6476) );
  NOR2_X1 U8345 ( .A1(n6501), .A2(n6476), .ZN(P2_U3247) );
  INV_X1 U8346 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n6477) );
  NOR2_X1 U8347 ( .A1(n6501), .A2(n6477), .ZN(P2_U3250) );
  INV_X1 U8348 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n6478) );
  NOR2_X1 U8349 ( .A1(n6501), .A2(n6478), .ZN(P2_U3248) );
  INV_X1 U8350 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n6479) );
  NOR2_X1 U8351 ( .A1(n6501), .A2(n6479), .ZN(P2_U3251) );
  INV_X1 U8352 ( .A(n6480), .ZN(n6483) );
  AOI22_X1 U8353 ( .A1(n7123), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9934), .ZN(n6481) );
  OAI21_X1 U8354 ( .B1(n6483), .B2(n4496), .A(n6481), .ZN(P1_U3344) );
  OAI222_X1 U8355 ( .A1(n8551), .A2(n6484), .B1(n8555), .B2(n6483), .C1(
        P2_U3151), .C2(n6482), .ZN(P2_U3284) );
  INV_X1 U8356 ( .A(n9601), .ZN(n10026) );
  INV_X2 U8357 ( .A(n9504), .ZN(P1_U3973) );
  NOR2_X1 U8358 ( .A1(n10026), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8359 ( .A(n9452), .ZN(n9322) );
  NAND2_X1 U8360 ( .A1(n9322), .A2(P1_U3973), .ZN(n6485) );
  OAI21_X1 U8361 ( .B1(P1_U3973), .B2(n7892), .A(n6485), .ZN(P1_U3585) );
  INV_X1 U8362 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6488) );
  INV_X1 U8363 ( .A(n6486), .ZN(n6489) );
  OAI222_X1 U8364 ( .A1(n8551), .A2(n6488), .B1(n8555), .B2(n6489), .C1(n6487), 
        .C2(P2_U3151), .ZN(P2_U3283) );
  INV_X1 U8365 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9043) );
  INV_X1 U8366 ( .A(n7374), .ZN(n7131) );
  OAI222_X1 U8367 ( .A1(n7819), .A2(n9043), .B1(n4496), .B2(n6489), .C1(n7131), 
        .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U8368 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6495) );
  NAND2_X1 U8369 ( .A1(n6533), .A2(P1_U3973), .ZN(n6494) );
  OAI21_X1 U8370 ( .B1(P1_U3973), .B2(n6495), .A(n6494), .ZN(P1_U3554) );
  INV_X1 U8371 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6498) );
  INV_X1 U8372 ( .A(n6496), .ZN(n6500) );
  OAI222_X1 U8373 ( .A1(n8551), .A2(n6498), .B1(n8555), .B2(n6500), .C1(
        P2_U3151), .C2(n6497), .ZN(P2_U3282) );
  INV_X1 U8374 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9023) );
  INV_X1 U8375 ( .A(n7482), .ZN(n6499) );
  OAI222_X1 U8376 ( .A1(n7819), .A2(n9023), .B1(n4496), .B2(n6500), .C1(
        P1_U3086), .C2(n6499), .ZN(P1_U3342) );
  INV_X1 U8377 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n6502) );
  NOR2_X1 U8378 ( .A1(n6501), .A2(n6502), .ZN(P2_U3244) );
  INV_X1 U8379 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n6503) );
  NOR2_X1 U8380 ( .A1(n6501), .A2(n6503), .ZN(P2_U3238) );
  INV_X1 U8381 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n6504) );
  NOR2_X1 U8382 ( .A1(n6501), .A2(n6504), .ZN(P2_U3256) );
  INV_X1 U8383 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n6505) );
  NOR2_X1 U8384 ( .A1(n6501), .A2(n6505), .ZN(P2_U3245) );
  INV_X1 U8385 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n6506) );
  NOR2_X1 U8386 ( .A1(n6501), .A2(n6506), .ZN(P2_U3255) );
  INV_X1 U8387 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n6507) );
  NOR2_X1 U8388 ( .A1(n6501), .A2(n6507), .ZN(P2_U3237) );
  NOR2_X1 U8389 ( .A1(n6501), .A2(n8961), .ZN(P2_U3240) );
  INV_X1 U8390 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n6508) );
  NOR2_X1 U8391 ( .A1(n6501), .A2(n6508), .ZN(P2_U3243) );
  INV_X1 U8392 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n6509) );
  NOR2_X1 U8393 ( .A1(n6501), .A2(n6509), .ZN(P2_U3257) );
  INV_X1 U8394 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n6510) );
  NOR2_X1 U8395 ( .A1(n6501), .A2(n6510), .ZN(P2_U3241) );
  INV_X1 U8396 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n6511) );
  NOR2_X1 U8397 ( .A1(n6501), .A2(n6511), .ZN(P2_U3236) );
  INV_X1 U8398 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n6512) );
  NOR2_X1 U8399 ( .A1(n6501), .A2(n6512), .ZN(P2_U3263) );
  INV_X1 U8400 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n6513) );
  NOR2_X1 U8401 ( .A1(n6501), .A2(n6513), .ZN(P2_U3234) );
  NOR2_X1 U8402 ( .A1(n6501), .A2(n9050), .ZN(P2_U3239) );
  NOR2_X1 U8403 ( .A1(n6501), .A2(n9094), .ZN(P2_U3254) );
  INV_X1 U8404 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n6514) );
  NOR2_X1 U8405 ( .A1(n6501), .A2(n6514), .ZN(P2_U3242) );
  INV_X1 U8406 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n6515) );
  NOR2_X1 U8407 ( .A1(n6501), .A2(n6515), .ZN(P2_U3235) );
  INV_X1 U8408 ( .A(n6516), .ZN(n6523) );
  AOI22_X1 U8409 ( .A1(n7767), .A2(P1_STATE_REG_SCAN_IN), .B1(n9934), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n6517) );
  OAI21_X1 U8410 ( .B1(n6523), .B2(n4496), .A(n6517), .ZN(P1_U3341) );
  INV_X1 U8411 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6521) );
  AND2_X1 U8412 ( .A1(n6533), .A2(n7275), .ZN(n9382) );
  OR2_X1 U8413 ( .A1(n9382), .A2(n7271), .ZN(n9336) );
  OAI21_X1 U8414 ( .B1(n10054), .B2(n10172), .A(n9336), .ZN(n6519) );
  NOR2_X1 U8415 ( .A1(n5729), .A2(n9195), .ZN(n7166) );
  INV_X1 U8416 ( .A(n7166), .ZN(n6518) );
  OAI211_X1 U8417 ( .C1(n7164), .C2(n7275), .A(n6519), .B(n6518), .ZN(n9876)
         );
  NAND2_X1 U8418 ( .A1(n9876), .A2(n10175), .ZN(n6520) );
  OAI21_X1 U8419 ( .B1(n10175), .B2(n6521), .A(n6520), .ZN(P1_U3453) );
  OAI222_X1 U8420 ( .A1(n8551), .A2(n6524), .B1(n8555), .B2(n6523), .C1(
        P2_U3151), .C2(n6522), .ZN(P2_U3281) );
  INV_X1 U8421 ( .A(n6530), .ZN(n6532) );
  INV_X1 U8422 ( .A(n6527), .ZN(n6525) );
  NAND2_X1 U8423 ( .A1(n6545), .A2(n5455), .ZN(n6526) );
  OAI22_X1 U8424 ( .A1(n6642), .A2(n8627), .B1(n6531), .B2(n7275), .ZN(n6630)
         );
  XNOR2_X1 U8425 ( .A(n6632), .B(n4501), .ZN(n10003) );
  INV_X1 U8426 ( .A(n6534), .ZN(n6536) );
  NAND2_X1 U8427 ( .A1(n6536), .A2(n6535), .ZN(n7167) );
  OR2_X1 U8428 ( .A1(n7167), .A2(n6537), .ZN(n6543) );
  AND2_X1 U8429 ( .A1(n10168), .A2(n6538), .ZN(n6539) );
  NAND2_X1 U8430 ( .A1(n6543), .A2(n10168), .ZN(n6541) );
  NAND2_X1 U8431 ( .A1(n6541), .A2(n6540), .ZN(n6927) );
  INV_X1 U8432 ( .A(n6927), .ZN(n6544) );
  OR2_X1 U8433 ( .A1(n7164), .A2(n7225), .ZN(n7171) );
  NOR2_X1 U8434 ( .A1(n7171), .A2(P1_U3086), .ZN(n6542) );
  NAND2_X1 U8435 ( .A1(n6543), .A2(n6542), .ZN(n6928) );
  NAND3_X1 U8436 ( .A1(n6544), .A2(n9475), .A3(n6928), .ZN(n6776) );
  AOI22_X1 U8437 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n6776), .B1(n7166), .B2(
        n9960), .ZN(n6552) );
  INV_X1 U8438 ( .A(n6546), .ZN(n6547) );
  OR2_X1 U8439 ( .A1(n6547), .A2(n7171), .ZN(n6550) );
  NAND2_X1 U8440 ( .A1(n9217), .A2(n7172), .ZN(n6551) );
  OAI211_X1 U8441 ( .C1(n10003), .C2(n9220), .A(n6552), .B(n6551), .ZN(
        P1_U3232) );
  NOR2_X1 U8442 ( .A1(n6785), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6553) );
  AOI21_X1 U8443 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n6785), .A(n6553), .ZN(
        n6558) );
  INV_X1 U8444 ( .A(n6554), .ZN(n6560) );
  NAND2_X1 U8445 ( .A1(n6812), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6556) );
  OAI21_X1 U8446 ( .B1(n6812), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6556), .ZN(
        n6807) );
  OAI21_X1 U8447 ( .B1(n6558), .B2(n6557), .A(n6781), .ZN(n6569) );
  AND2_X1 U8448 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7603) );
  AOI21_X1 U8449 ( .B1(n10026), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n7603), .ZN(
        n6566) );
  INV_X1 U8450 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10189) );
  AOI22_X1 U8451 ( .A1(n6785), .A2(P1_REG1_REG_9__SCAN_IN), .B1(n10189), .B2(
        n6567), .ZN(n6563) );
  AOI21_X1 U8452 ( .B1(n6560), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6559), .ZN(
        n6811) );
  NAND2_X1 U8453 ( .A1(n6812), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6561) );
  OAI21_X1 U8454 ( .B1(n6812), .B2(P1_REG1_REG_8__SCAN_IN), .A(n6561), .ZN(
        n6810) );
  OAI21_X1 U8455 ( .B1(n6563), .B2(n6562), .A(n6784), .ZN(n6564) );
  NAND2_X1 U8456 ( .A1(n10017), .A2(n6564), .ZN(n6565) );
  OAI211_X1 U8457 ( .C1(n7132), .C2(n6567), .A(n6566), .B(n6565), .ZN(n6568)
         );
  AOI21_X1 U8458 ( .B1(n9593), .B2(n6569), .A(n6568), .ZN(n6570) );
  INV_X1 U8459 ( .A(n6570), .ZN(P1_U3252) );
  INV_X1 U8460 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9118) );
  INV_X1 U8461 ( .A(n6717), .ZN(n8290) );
  NAND2_X1 U8462 ( .A1(n8290), .A2(n6654), .ZN(n7960) );
  AND2_X1 U8463 ( .A1(n6712), .A2(n7960), .ZN(n7910) );
  NOR2_X1 U8464 ( .A1(n10408), .A2(n8430), .ZN(n6571) );
  OR2_X1 U8465 ( .A1(n7910), .A2(n6571), .ZN(n6574) );
  OR2_X1 U8466 ( .A1(n5995), .A2(n8389), .ZN(n6674) );
  OAI21_X1 U8467 ( .B1(n10418), .B2(n6654), .A(n6674), .ZN(n6572) );
  INV_X1 U8468 ( .A(n6572), .ZN(n6573) );
  NAND2_X1 U8469 ( .A1(n6574), .A2(n6573), .ZN(n8494) );
  NAND2_X1 U8470 ( .A1(n10430), .A2(n8494), .ZN(n6575) );
  OAI21_X1 U8471 ( .B1(n10430), .B2(n9118), .A(n6575), .ZN(P2_U3390) );
  OAI21_X1 U8472 ( .B1(n6576), .B2(n7981), .A(n6577), .ZN(n10361) );
  AND2_X1 U8473 ( .A1(n6579), .A2(n6578), .ZN(n6580) );
  XNOR2_X1 U8474 ( .A(n6580), .B(n7981), .ZN(n6581) );
  OAI222_X1 U8475 ( .A1(n8391), .A2(n6692), .B1(n8389), .B2(n6043), .C1(n6581), 
        .C2(n8387), .ZN(n10360) );
  AOI21_X1 U8476 ( .B1(n10408), .B2(n10361), .A(n10360), .ZN(n6598) );
  OAI22_X1 U8477 ( .A1(n8451), .A2(n10364), .B1(n10446), .B2(n9037), .ZN(n6582) );
  INV_X1 U8478 ( .A(n6582), .ZN(n6583) );
  OAI21_X1 U8479 ( .B1(n6598), .B2(n10444), .A(n6583), .ZN(P2_U3463) );
  OAI21_X1 U8480 ( .B1(n6585), .B2(n6584), .A(n7013), .ZN(n6587) );
  OAI22_X1 U8481 ( .A1(n5995), .A2(n8391), .B1(n6692), .B2(n8389), .ZN(n6586)
         );
  AOI21_X1 U8482 ( .B1(n6587), .B2(n8430), .A(n6586), .ZN(n6591) );
  OAI21_X1 U8483 ( .B1(n6589), .B2(n7971), .A(n6588), .ZN(n10377) );
  INV_X1 U8484 ( .A(n7200), .ZN(n6746) );
  NAND2_X1 U8485 ( .A1(n10377), .A2(n6746), .ZN(n6590) );
  AND2_X1 U8486 ( .A1(n6591), .A2(n6590), .ZN(n10374) );
  AOI22_X1 U8487 ( .A1(n10377), .A2(n6328), .B1(n10429), .B2(n6658), .ZN(n6592) );
  AND2_X1 U8488 ( .A1(n10374), .A2(n6592), .ZN(n10388) );
  MUX2_X1 U8489 ( .A(n6593), .B(n10388), .S(n10446), .Z(n6594) );
  INV_X1 U8490 ( .A(n6594), .ZN(P2_U3461) );
  INV_X1 U8491 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6595) );
  OAI22_X1 U8492 ( .A1(n10364), .A2(n8507), .B1(n10430), .B2(n6595), .ZN(n6596) );
  INV_X1 U8493 ( .A(n6596), .ZN(n6597) );
  OAI21_X1 U8494 ( .B1(n6598), .B2(n10432), .A(n6597), .ZN(P2_U3402) );
  INV_X1 U8495 ( .A(n6599), .ZN(n6602) );
  OAI222_X1 U8496 ( .A1(P1_U3086), .A2(n9542), .B1(n4496), .B2(n6602), .C1(
        n6600), .C2(n7819), .ZN(P1_U3340) );
  OAI222_X1 U8497 ( .A1(n8551), .A2(n9103), .B1(n8555), .B2(n6602), .C1(n6601), 
        .C2(P2_U3151), .ZN(P2_U3280) );
  OR2_X1 U8498 ( .A1(n6606), .A2(n10418), .ZN(n6604) );
  INV_X1 U8499 ( .A(n8237), .ZN(n8266) );
  OR2_X1 U8500 ( .A1(n6606), .A2(n6605), .ZN(n6609) );
  INV_X1 U8501 ( .A(n6607), .ZN(n6618) );
  NAND2_X1 U8502 ( .A1(n6610), .A2(n6618), .ZN(n6608) );
  INV_X1 U8503 ( .A(n7910), .ZN(n6614) );
  INV_X1 U8504 ( .A(n6610), .ZN(n6611) );
  NOR2_X1 U8505 ( .A1(n6611), .A2(n6675), .ZN(n6657) );
  INV_X1 U8506 ( .A(n6656), .ZN(n6612) );
  AOI22_X1 U8507 ( .A1(n8242), .A2(n6614), .B1(n8257), .B2(n6652), .ZN(n6629)
         );
  INV_X1 U8508 ( .A(n6615), .ZN(n6617) );
  NAND2_X1 U8509 ( .A1(n6617), .A2(n6616), .ZN(n6621) );
  NAND2_X1 U8510 ( .A1(n6624), .A2(n6618), .ZN(n6619) );
  NAND3_X1 U8511 ( .A1(n6621), .A2(n6620), .A3(n6619), .ZN(n6622) );
  NAND2_X1 U8512 ( .A1(n6622), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6626) );
  NOR2_X1 U8513 ( .A1(n6623), .A2(n6675), .ZN(n8126) );
  NAND2_X1 U8514 ( .A1(n6624), .A2(n8126), .ZN(n6625) );
  NAND2_X1 U8515 ( .A1(n6696), .A2(n6627), .ZN(n6944) );
  NAND2_X1 U8516 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(n6944), .ZN(n6628) );
  OAI211_X1 U8517 ( .C1(n8266), .C2(n6654), .A(n6629), .B(n6628), .ZN(P2_U3172) );
  OAI22_X1 U8518 ( .A1(n6632), .A2(n4501), .B1(n7517), .B2(n6630), .ZN(n6641)
         );
  NAND2_X1 U8519 ( .A1(n6633), .A2(n8733), .ZN(n6635) );
  NAND2_X1 U8520 ( .A1(n7279), .A2(n7040), .ZN(n6634) );
  NAND2_X1 U8521 ( .A1(n6633), .A2(n8653), .ZN(n6637) );
  NAND2_X1 U8522 ( .A1(n7279), .A2(n8733), .ZN(n6636) );
  AND2_X1 U8523 ( .A1(n6637), .A2(n6636), .ZN(n6638) );
  OAI21_X1 U8524 ( .B1(n6639), .B2(n6638), .A(n6761), .ZN(n6640) );
  AOI21_X1 U8525 ( .B1(n6641), .B2(n6640), .A(n6771), .ZN(n6645) );
  OAI22_X1 U8526 ( .A1(n6642), .A2(n9141), .B1(n6930), .B2(n9195), .ZN(n7272)
         );
  AOI22_X1 U8527 ( .A1(n7272), .A2(n9960), .B1(n6776), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n6644) );
  NAND2_X1 U8528 ( .A1(n9217), .A2(n7279), .ZN(n6643) );
  OAI211_X1 U8529 ( .C1(n6645), .C2(n9220), .A(n6644), .B(n6643), .ZN(P1_U3222) );
  NAND2_X1 U8530 ( .A1(n9504), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6646) );
  OAI21_X1 U8531 ( .B1(n8736), .B2(n9504), .A(n6646), .ZN(P1_U3582) );
  XNOR2_X1 U8532 ( .A(n7963), .B(n8118), .ZN(n6647) );
  XNOR2_X1 U8533 ( .A(n6653), .B(n10371), .ZN(n6682) );
  XNOR2_X1 U8534 ( .A(n6682), .B(n6942), .ZN(n6684) );
  AOI21_X1 U8535 ( .B1(n6681), .B2(n6654), .A(n6296), .ZN(n6939) );
  XOR2_X1 U8536 ( .A(n6684), .B(n6685), .Z(n6662) );
  AOI22_X1 U8537 ( .A1(n8244), .A2(n6652), .B1(n8237), .B2(n6658), .ZN(n6659)
         );
  OAI21_X1 U8538 ( .B1(n6692), .B2(n8246), .A(n6659), .ZN(n6660) );
  AOI21_X1 U8539 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n6944), .A(n6660), .ZN(
        n6661) );
  OAI21_X1 U8540 ( .B1(n8251), .B2(n6662), .A(n6661), .ZN(P2_U3177) );
  INV_X1 U8541 ( .A(n6663), .ZN(n6671) );
  OR2_X1 U8542 ( .A1(n6665), .A2(n6664), .ZN(n6669) );
  OR2_X1 U8543 ( .A1(n6667), .A2(n6666), .ZN(n6668) );
  NAND4_X1 U8544 ( .A1(n6671), .A2(n6670), .A3(n6669), .A4(n6668), .ZN(n6672)
         );
  AOI22_X1 U8545 ( .A1(n8434), .A2(n6673), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n8404), .ZN(n6680) );
  INV_X1 U8546 ( .A(n6674), .ZN(n6678) );
  INV_X1 U8547 ( .A(n6675), .ZN(n6676) );
  NOR3_X1 U8548 ( .A1(n7910), .A2(n10429), .A3(n6676), .ZN(n6677) );
  OAI21_X1 U8549 ( .B1(n6678), .B2(n6677), .A(n4495), .ZN(n6679) );
  OAI211_X1 U8550 ( .C1(n5988), .C2(n4495), .A(n6680), .B(n6679), .ZN(P2_U3233) );
  XNOR2_X1 U8551 ( .A(n6653), .B(n10364), .ZN(n6701) );
  XNOR2_X1 U8552 ( .A(n6701), .B(n8287), .ZN(n6691) );
  INV_X1 U8553 ( .A(n6682), .ZN(n6683) );
  XNOR2_X1 U8554 ( .A(n6653), .B(n7017), .ZN(n6686) );
  XNOR2_X1 U8555 ( .A(n6686), .B(n6692), .ZN(n6757) );
  NAND2_X1 U8556 ( .A1(n6758), .A2(n6757), .ZN(n6756) );
  NAND2_X1 U8557 ( .A1(n6686), .A2(n8288), .ZN(n6687) );
  NAND2_X1 U8558 ( .A1(n6756), .A2(n6687), .ZN(n6690) );
  AOI21_X1 U8559 ( .B1(n6691), .B2(n6690), .A(n6689), .ZN(n6700) );
  INV_X1 U8560 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n8892) );
  NOR2_X1 U8561 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8892), .ZN(n6969) );
  OAI22_X1 U8562 ( .A1(n6043), .A2(n8246), .B1(n8260), .B2(n6692), .ZN(n6693)
         );
  AOI211_X1 U8563 ( .C1(n6694), .C2(n8237), .A(n6969), .B(n6693), .ZN(n6699)
         );
  NAND2_X1 U8564 ( .A1(n6695), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8130) );
  INV_X1 U8565 ( .A(n10366), .ZN(n6697) );
  NAND2_X1 U8566 ( .A1(n8262), .A2(n6697), .ZN(n6698) );
  OAI211_X1 U8567 ( .C1(n6700), .C2(n8251), .A(n6699), .B(n6698), .ZN(P2_U3170) );
  INV_X1 U8568 ( .A(n6701), .ZN(n6702) );
  XNOR2_X1 U8569 ( .A(n6958), .B(n6957), .ZN(n6705) );
  NAND2_X1 U8570 ( .A1(n6705), .A2(n8242), .ZN(n6709) );
  NOR2_X1 U8571 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6706), .ZN(n6844) );
  OAI22_X1 U8572 ( .A1(n6754), .A2(n8260), .B1(n8246), .B2(n7063), .ZN(n6707)
         );
  AOI211_X1 U8573 ( .C1(n10394), .C2(n8237), .A(n6844), .B(n6707), .ZN(n6708)
         );
  OAI211_X1 U8574 ( .C1(n6748), .C2(n8210), .A(n6709), .B(n6708), .ZN(P2_U3167) );
  NAND2_X1 U8575 ( .A1(n6711), .A2(n6712), .ZN(n6713) );
  AND2_X1 U8576 ( .A1(n6714), .A2(n7957), .ZN(n10378) );
  NAND2_X1 U8577 ( .A1(n4495), .A2(n10378), .ZN(n7811) );
  OAI21_X1 U8578 ( .B1(n6716), .B2(n6711), .A(n6715), .ZN(n6720) );
  OAI22_X1 U8579 ( .A1(n6942), .A2(n8389), .B1(n6717), .B2(n8391), .ZN(n6719)
         );
  NOR2_X1 U8580 ( .A1(n10384), .A2(n7200), .ZN(n6718) );
  AOI211_X1 U8581 ( .C1(n8430), .C2(n6720), .A(n6719), .B(n6718), .ZN(n10382)
         );
  MUX2_X1 U8582 ( .A(n10194), .B(n10382), .S(n4495), .Z(n6722) );
  AOI22_X1 U8583 ( .A1(n8419), .A2(n6940), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8404), .ZN(n6721) );
  OAI211_X1 U8584 ( .C1(n10384), .C2(n7811), .A(n6722), .B(n6721), .ZN(
        P2_U3232) );
  INV_X1 U8585 ( .A(n6723), .ZN(n6832) );
  AOI22_X1 U8586 ( .A1(n9561), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9934), .ZN(n6724) );
  OAI21_X1 U8587 ( .B1(n6832), .B2(n4496), .A(n6724), .ZN(P1_U3339) );
  AOI211_X1 U8588 ( .C1(n10002), .C2(n6726), .A(n6725), .B(n10018), .ZN(n6734)
         );
  AOI22_X1 U8589 ( .A1(n10026), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n6731) );
  OAI211_X1 U8590 ( .C1(n6729), .C2(n6728), .A(n10017), .B(n6727), .ZN(n6730)
         );
  OAI211_X1 U8591 ( .C1(n7132), .C2(n6732), .A(n6731), .B(n6730), .ZN(n6733)
         );
  OR2_X1 U8592 ( .A1(n6734), .A2(n6733), .ZN(P1_U3244) );
  XNOR2_X1 U8593 ( .A(n8286), .B(n6736), .ZN(n7912) );
  INV_X1 U8594 ( .A(n7912), .ZN(n6743) );
  XNOR2_X1 U8595 ( .A(n6735), .B(n6743), .ZN(n10395) );
  INV_X1 U8596 ( .A(n10395), .ZN(n6752) );
  OAI22_X1 U8597 ( .A1(n6754), .A2(n8391), .B1(n7063), .B2(n8389), .ZN(n6745)
         );
  NAND2_X1 U8598 ( .A1(n6737), .A2(n6738), .ZN(n6742) );
  NAND2_X1 U8599 ( .A1(n6737), .A2(n6739), .ZN(n7001) );
  INV_X1 U8600 ( .A(n7000), .ZN(n6740) );
  NOR2_X1 U8601 ( .A1(n7001), .A2(n6740), .ZN(n6741) );
  AOI211_X1 U8602 ( .C1(n6743), .C2(n6742), .A(n8387), .B(n6741), .ZN(n6744)
         );
  AOI211_X1 U8603 ( .C1(n6746), .C2(n10395), .A(n6745), .B(n6744), .ZN(n10397)
         );
  MUX2_X1 U8604 ( .A(n6747), .B(n10397), .S(n4495), .Z(n6751) );
  INV_X1 U8605 ( .A(n6748), .ZN(n6749) );
  AOI22_X1 U8606 ( .A1(n8419), .A2(n10394), .B1(n8404), .B2(n6749), .ZN(n6750)
         );
  OAI211_X1 U8607 ( .C1(n6752), .C2(n7811), .A(n6751), .B(n6750), .ZN(P2_U3228) );
  INV_X1 U8608 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6753) );
  NOR2_X1 U8609 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6753), .ZN(n6986) );
  OAI22_X1 U8610 ( .A1(n6942), .A2(n8260), .B1(n8246), .B2(n6754), .ZN(n6755)
         );
  AOI211_X1 U8611 ( .C1(n10390), .C2(n8237), .A(n6986), .B(n6755), .ZN(n6760)
         );
  OAI211_X1 U8612 ( .C1(n6758), .C2(n6757), .A(n6756), .B(n8242), .ZN(n6759)
         );
  OAI211_X1 U8613 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8210), .A(n6760), .B(
        n6759), .ZN(P2_U3158) );
  INV_X1 U8614 ( .A(n6761), .ZN(n6773) );
  INV_X1 U8615 ( .A(n7040), .ZN(n8609) );
  XNOR2_X1 U8616 ( .A(n6762), .B(n8731), .ZN(n6766) );
  OR2_X1 U8617 ( .A1(n6930), .A2(n4503), .ZN(n6765) );
  NAND2_X1 U8618 ( .A1(n6763), .A2(n8733), .ZN(n6764) );
  AND2_X1 U8619 ( .A1(n6765), .A2(n6764), .ZN(n6767) );
  NAND2_X1 U8620 ( .A1(n6766), .A2(n6767), .ZN(n6922) );
  INV_X1 U8621 ( .A(n6766), .ZN(n6769) );
  INV_X1 U8622 ( .A(n6767), .ZN(n6768) );
  NAND2_X1 U8623 ( .A1(n6769), .A2(n6768), .ZN(n6770) );
  INV_X1 U8624 ( .A(n6923), .ZN(n6775) );
  NOR3_X1 U8625 ( .A1(n6771), .A2(n6773), .A3(n6772), .ZN(n6774) );
  OAI21_X1 U8626 ( .B1(n6775), .B2(n6774), .A(n9966), .ZN(n6778) );
  OAI22_X1 U8627 ( .A1(n5729), .A2(n9141), .B1(n6919), .B2(n9195), .ZN(n7263)
         );
  AOI22_X1 U8628 ( .A1(n7263), .A2(n9960), .B1(n6776), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n6777) );
  OAI211_X1 U8629 ( .C1(n5507), .C2(n9963), .A(n6778), .B(n6777), .ZN(P1_U3237) );
  INV_X1 U8630 ( .A(n6779), .ZN(n6835) );
  AOI22_X1 U8631 ( .A1(n9578), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9934), .ZN(n6780) );
  OAI21_X1 U8632 ( .B1(n6835), .B2(n4496), .A(n6780), .ZN(P1_U3338) );
  OAI21_X1 U8633 ( .B1(n6785), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6781), .ZN(
        n6783) );
  INV_X1 U8634 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7392) );
  MUX2_X1 U8635 ( .A(n7392), .B(P1_REG2_REG_10__SCAN_IN), .S(n7071), .Z(n6782)
         );
  NOR2_X1 U8636 ( .A1(n6782), .A2(n6783), .ZN(n7067) );
  AOI211_X1 U8637 ( .C1(n6783), .C2(n6782), .A(n7067), .B(n10018), .ZN(n6793)
         );
  INV_X1 U8638 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6786) );
  MUX2_X1 U8639 ( .A(n6786), .B(P1_REG1_REG_10__SCAN_IN), .S(n7071), .Z(n6787)
         );
  NOR2_X1 U8640 ( .A1(n6787), .A2(n6788), .ZN(n7070) );
  AOI211_X1 U8641 ( .C1(n6788), .C2(n6787), .A(n7070), .B(n9993), .ZN(n6792)
         );
  INV_X1 U8642 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9115) );
  NAND2_X1 U8643 ( .A1(n10025), .A2(n7071), .ZN(n6790) );
  NAND2_X1 U8644 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n6789) );
  OAI211_X1 U8645 ( .C1(n9115), .C2(n9601), .A(n6790), .B(n6789), .ZN(n6791)
         );
  OR3_X1 U8646 ( .A1(n6793), .A2(n6792), .A3(n6791), .ZN(P1_U3253) );
  AOI211_X1 U8647 ( .C1(n6796), .C2(n6795), .A(n6794), .B(n10018), .ZN(n6805)
         );
  AOI211_X1 U8648 ( .C1(n6799), .C2(n6798), .A(n6797), .B(n9993), .ZN(n6804)
         );
  INV_X1 U8649 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6802) );
  NAND2_X1 U8650 ( .A1(n10025), .A2(n6800), .ZN(n6801) );
  NAND2_X1 U8651 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n7219) );
  OAI211_X1 U8652 ( .C1(n6802), .C2(n9601), .A(n6801), .B(n7219), .ZN(n6803)
         );
  OR3_X1 U8653 ( .A1(n6805), .A2(n6804), .A3(n6803), .ZN(P1_U3248) );
  AOI211_X1 U8654 ( .C1(n6808), .C2(n6807), .A(n6806), .B(n10018), .ZN(n6818)
         );
  AOI211_X1 U8655 ( .C1(n6811), .C2(n6810), .A(n6809), .B(n9993), .ZN(n6817)
         );
  INV_X1 U8656 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6815) );
  NAND2_X1 U8657 ( .A1(n10025), .A2(n6812), .ZN(n6814) );
  NAND2_X1 U8658 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n6813) );
  OAI211_X1 U8659 ( .C1(n6815), .C2(n9601), .A(n6814), .B(n6813), .ZN(n6816)
         );
  OR3_X1 U8660 ( .A1(n6818), .A2(n6817), .A3(n6816), .ZN(P1_U3251) );
  AOI211_X1 U8661 ( .C1(n6821), .C2(n6820), .A(n10018), .B(n6819), .ZN(n6830)
         );
  AOI211_X1 U8662 ( .C1(n6824), .C2(n6823), .A(n6822), .B(n9993), .ZN(n6829)
         );
  INV_X1 U8663 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6827) );
  NAND2_X1 U8664 ( .A1(n10025), .A2(n6825), .ZN(n6826) );
  NAND2_X1 U8665 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7329) );
  OAI211_X1 U8666 ( .C1(n6827), .C2(n9601), .A(n6826), .B(n7329), .ZN(n6828)
         );
  OR3_X1 U8667 ( .A1(n6830), .A2(n6829), .A3(n6828), .ZN(P1_U3249) );
  OAI222_X1 U8668 ( .A1(n8551), .A2(n6833), .B1(n8555), .B2(n6832), .C1(
        P2_U3151), .C2(n6831), .ZN(P2_U3279) );
  OAI222_X1 U8669 ( .A1(n8551), .A2(n6836), .B1(n8555), .B2(n6835), .C1(n6834), 
        .C2(P2_U3151), .ZN(P2_U3278) );
  XNOR2_X1 U8670 ( .A(n6838), .B(n6837), .ZN(n6848) );
  INV_X1 U8671 ( .A(n10347), .ZN(n7025) );
  XNOR2_X1 U8672 ( .A(n6839), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n6842) );
  XNOR2_X1 U8673 ( .A(n6840), .B(P2_REG2_REG_5__SCAN_IN), .ZN(n6841) );
  OAI22_X1 U8674 ( .A1(n7025), .A2(n6842), .B1(n6841), .B2(n6993), .ZN(n6843)
         );
  AOI211_X1 U8675 ( .C1(n10339), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n6844), .B(
        n6843), .ZN(n6847) );
  NAND2_X1 U8676 ( .A1(n10340), .A2(n6845), .ZN(n6846) );
  OAI211_X1 U8677 ( .C1(n6848), .C2(n10354), .A(n6847), .B(n6846), .ZN(
        P2_U3187) );
  INV_X1 U8678 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6853) );
  OAI21_X1 U8679 ( .B1(n10102), .B2(P1_D_REG_1__SCAN_IN), .A(n6851), .ZN(n6852) );
  OAI21_X1 U8680 ( .B1(n9475), .B2(n6853), .A(n6852), .ZN(P1_U3440) );
  AOI21_X1 U8681 ( .B1(n6856), .B2(n6855), .A(n6854), .ZN(n6871) );
  INV_X1 U8682 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6867) );
  OAI21_X1 U8683 ( .B1(n6859), .B2(n6858), .A(n6857), .ZN(n6864) );
  OAI21_X1 U8684 ( .B1(n6862), .B2(n6861), .A(n6860), .ZN(n6863) );
  AOI22_X1 U8685 ( .A1(n10347), .A2(n6864), .B1(n10348), .B2(n6863), .ZN(n6866) );
  INV_X1 U8686 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9035) );
  NOR2_X1 U8687 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9035), .ZN(n6963) );
  INV_X1 U8688 ( .A(n6963), .ZN(n6865) );
  OAI211_X1 U8689 ( .C1(n10200), .C2(n6867), .A(n6866), .B(n6865), .ZN(n6868)
         );
  AOI21_X1 U8690 ( .B1(n6869), .B2(n10340), .A(n6868), .ZN(n6870) );
  OAI21_X1 U8691 ( .B1(n6871), .B2(n10354), .A(n6870), .ZN(P2_U3188) );
  AOI21_X1 U8692 ( .B1(n6874), .B2(n6873), .A(n6872), .ZN(n6889) );
  AOI21_X1 U8693 ( .B1(n6877), .B2(n6876), .A(n6875), .ZN(n6884) );
  OAI21_X1 U8694 ( .B1(n6880), .B2(n6879), .A(n6878), .ZN(n6881) );
  NAND2_X1 U8695 ( .A1(n10347), .A2(n6881), .ZN(n6883) );
  NOR2_X1 U8696 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5962), .ZN(n7111) );
  INV_X1 U8697 ( .A(n7111), .ZN(n6882) );
  OAI211_X1 U8698 ( .C1(n6884), .C2(n10354), .A(n6883), .B(n6882), .ZN(n6885)
         );
  AOI21_X1 U8699 ( .B1(n10339), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6885), .ZN(
        n6888) );
  NAND2_X1 U8700 ( .A1(n10340), .A2(n6886), .ZN(n6887) );
  OAI211_X1 U8701 ( .C1(n6889), .C2(n6993), .A(n6888), .B(n6887), .ZN(P2_U3190) );
  INV_X1 U8702 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6896) );
  NAND2_X1 U8703 ( .A1(n6890), .A2(n10354), .ZN(n6893) );
  OAI21_X1 U8704 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6891), .A(n10203), .ZN(
        n6892) );
  AOI22_X1 U8705 ( .A1(n6893), .A2(n6892), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        P2_U3151), .ZN(n6895) );
  NAND2_X1 U8706 ( .A1(n10340), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6894) );
  OAI211_X1 U8707 ( .C1(n10200), .C2(n6896), .A(n6895), .B(n6894), .ZN(
        P2_U3182) );
  INV_X1 U8708 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10453) );
  NOR2_X1 U8709 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n6897) );
  AOI21_X1 U8710 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n6897), .ZN(n10458) );
  NOR2_X1 U8711 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(P2_ADDR_REG_16__SCAN_IN), 
        .ZN(n6898) );
  AOI21_X1 U8712 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n6898), .ZN(n10461) );
  NOR2_X1 U8713 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n6899) );
  AOI21_X1 U8714 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n6899), .ZN(n10464) );
  NOR2_X1 U8715 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n6900) );
  AOI21_X1 U8716 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n6900), .ZN(n10467) );
  NOR2_X1 U8717 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n6901) );
  AOI21_X1 U8718 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n6901), .ZN(n10470) );
  NOR2_X1 U8719 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n6902) );
  AOI21_X1 U8720 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n6902), .ZN(n10473) );
  NOR2_X1 U8721 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n6903) );
  AOI21_X1 U8722 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n6903), .ZN(n10476) );
  NOR2_X1 U8723 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n6904) );
  AOI21_X1 U8724 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n6904), .ZN(n10479) );
  NOR2_X1 U8725 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(P2_ADDR_REG_9__SCAN_IN), 
        .ZN(n6905) );
  AOI21_X1 U8726 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n6905), .ZN(n10488) );
  NOR2_X1 U8727 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n6906) );
  AOI21_X1 U8728 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n6906), .ZN(n10494) );
  NOR2_X1 U8729 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n6907) );
  AOI21_X1 U8730 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n6907), .ZN(n10491) );
  NOR2_X1 U8731 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n6908) );
  AOI21_X1 U8732 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n6908), .ZN(n10482) );
  NOR2_X1 U8733 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n6909) );
  AOI21_X1 U8734 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n6909), .ZN(n10485) );
  AND2_X1 U8735 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n6910) );
  NOR2_X1 U8736 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n6910), .ZN(n10448) );
  INV_X1 U8737 ( .A(n10448), .ZN(n10449) );
  INV_X1 U8738 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10451) );
  NAND3_X1 U8739 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10450) );
  NAND2_X1 U8740 ( .A1(n10451), .A2(n10450), .ZN(n10447) );
  NAND2_X1 U8741 ( .A1(n10449), .A2(n10447), .ZN(n10497) );
  NAND2_X1 U8742 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n6911) );
  OAI21_X1 U8743 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n6911), .ZN(n10496) );
  NOR2_X1 U8744 ( .A1(n10497), .A2(n10496), .ZN(n10495) );
  AOI21_X1 U8745 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10495), .ZN(n10500) );
  NAND2_X1 U8746 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n6912) );
  OAI21_X1 U8747 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n6912), .ZN(n10499) );
  NOR2_X1 U8748 ( .A1(n10500), .A2(n10499), .ZN(n10498) );
  AOI21_X1 U8749 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10498), .ZN(n10503) );
  NOR2_X1 U8750 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n6913) );
  AOI21_X1 U8751 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n6913), .ZN(n10502) );
  NAND2_X1 U8752 ( .A1(n10503), .A2(n10502), .ZN(n10501) );
  OAI21_X1 U8753 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10501), .ZN(n10484) );
  NAND2_X1 U8754 ( .A1(n10485), .A2(n10484), .ZN(n10483) );
  OAI21_X1 U8755 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10483), .ZN(n10481) );
  NAND2_X1 U8756 ( .A1(n10482), .A2(n10481), .ZN(n10480) );
  OAI21_X1 U8757 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n10480), .ZN(n10490) );
  NAND2_X1 U8758 ( .A1(n10491), .A2(n10490), .ZN(n10489) );
  OAI21_X1 U8759 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10489), .ZN(n10493) );
  NAND2_X1 U8760 ( .A1(n10494), .A2(n10493), .ZN(n10492) );
  OAI21_X1 U8761 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10492), .ZN(n10487) );
  NAND2_X1 U8762 ( .A1(n10488), .A2(n10487), .ZN(n10486) );
  OAI21_X1 U8763 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n10486), .ZN(n10478) );
  NAND2_X1 U8764 ( .A1(n10479), .A2(n10478), .ZN(n10477) );
  OAI21_X1 U8765 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10477), .ZN(n10475) );
  NAND2_X1 U8766 ( .A1(n10476), .A2(n10475), .ZN(n10474) );
  OAI21_X1 U8767 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10474), .ZN(n10472) );
  NAND2_X1 U8768 ( .A1(n10473), .A2(n10472), .ZN(n10471) );
  OAI21_X1 U8769 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10471), .ZN(n10469) );
  NAND2_X1 U8770 ( .A1(n10470), .A2(n10469), .ZN(n10468) );
  OAI21_X1 U8771 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10468), .ZN(n10466) );
  NAND2_X1 U8772 ( .A1(n10467), .A2(n10466), .ZN(n10465) );
  OAI21_X1 U8773 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10465), .ZN(n10463) );
  NAND2_X1 U8774 ( .A1(n10464), .A2(n10463), .ZN(n10462) );
  OAI21_X1 U8775 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10462), .ZN(n10460) );
  NAND2_X1 U8776 ( .A1(n10461), .A2(n10460), .ZN(n10459) );
  OAI21_X1 U8777 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n10459), .ZN(n10457) );
  NAND2_X1 U8778 ( .A1(n10458), .A2(n10457), .ZN(n10456) );
  OAI21_X1 U8779 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10456), .ZN(n10454) );
  NOR2_X1 U8780 ( .A1(n10453), .A2(n10454), .ZN(n6914) );
  NAND2_X1 U8781 ( .A1(n10453), .A2(n10454), .ZN(n10452) );
  OAI21_X1 U8782 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n6914), .A(n10452), .ZN(
        n6917) );
  XNOR2_X1 U8783 ( .A(n6915), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n6916) );
  XNOR2_X1 U8784 ( .A(n6917), .B(n6916), .ZN(ADD_1068_U4) );
  AOI22_X1 U8785 ( .A1(n9516), .A2(n8733), .B1(n5515), .B2(n8727), .ZN(n6918)
         );
  XNOR2_X1 U8786 ( .A(n6918), .B(n7517), .ZN(n7039) );
  OR2_X1 U8787 ( .A1(n6919), .A2(n4503), .ZN(n6921) );
  NAND2_X1 U8788 ( .A1(n5515), .A2(n8733), .ZN(n6920) );
  NAND2_X1 U8789 ( .A1(n6921), .A2(n6920), .ZN(n7037) );
  XNOR2_X1 U8790 ( .A(n7039), .B(n7037), .ZN(n6925) );
  OAI21_X1 U8791 ( .B1(n6925), .B2(n6924), .A(n7044), .ZN(n6936) );
  OAI21_X1 U8792 ( .B1(n6927), .B2(n6926), .A(P1_STATE_REG_SCAN_IN), .ZN(n6929) );
  OR2_X1 U8793 ( .A1(n6930), .A2(n9141), .ZN(n6932) );
  OR2_X1 U8794 ( .A1(n5524), .A2(n9195), .ZN(n6931) );
  NAND2_X1 U8795 ( .A1(n6932), .A2(n6931), .ZN(n10053) );
  AOI22_X1 U8796 ( .A1(n10053), .A2(n9960), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        P1_U3086), .ZN(n6934) );
  NAND2_X1 U8797 ( .A1(n9217), .A2(n5515), .ZN(n6933) );
  OAI211_X1 U8798 ( .C1(n9970), .C2(P1_REG3_REG_3__SCAN_IN), .A(n6934), .B(
        n6933), .ZN(n6935) );
  AOI21_X1 U8799 ( .B1(n6936), .B2(n9966), .A(n6935), .ZN(n6937) );
  INV_X1 U8800 ( .A(n6937), .ZN(P1_U3218) );
  XOR2_X1 U8801 ( .A(n6939), .B(n6938), .Z(n6946) );
  AOI22_X1 U8802 ( .A1(n8244), .A2(n8290), .B1(n8237), .B2(n6940), .ZN(n6941)
         );
  OAI21_X1 U8803 ( .B1(n6942), .B2(n8246), .A(n6941), .ZN(n6943) );
  AOI21_X1 U8804 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n6944), .A(n6943), .ZN(
        n6945) );
  OAI21_X1 U8805 ( .B1(n8251), .B2(n6946), .A(n6945), .ZN(P2_U3162) );
  AND2_X1 U8806 ( .A1(n7945), .A2(n7949), .ZN(n7916) );
  INV_X1 U8807 ( .A(n7916), .ZN(n6951) );
  XNOR2_X1 U8808 ( .A(n6947), .B(n6951), .ZN(n6949) );
  OAI22_X1 U8809 ( .A1(n7058), .A2(n8391), .B1(n7426), .B2(n8389), .ZN(n6948)
         );
  AOI21_X1 U8810 ( .B1(n6949), .B2(n8430), .A(n6948), .ZN(n10411) );
  XNOR2_X1 U8811 ( .A(n6950), .B(n6951), .ZN(n10409) );
  INV_X1 U8812 ( .A(n10378), .ZN(n6952) );
  NAND2_X1 U8813 ( .A1(n7200), .A2(n6952), .ZN(n10362) );
  INV_X1 U8814 ( .A(n8419), .ZN(n10365) );
  INV_X1 U8815 ( .A(n6953), .ZN(n7116) );
  AOI22_X1 U8816 ( .A1(n10381), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n8404), .B2(
        n7116), .ZN(n6954) );
  OAI21_X1 U8817 ( .B1(n7114), .B2(n10365), .A(n6954), .ZN(n6955) );
  AOI21_X1 U8818 ( .B1(n10409), .B2(n8438), .A(n6955), .ZN(n6956) );
  OAI21_X1 U8819 ( .B1(n10411), .B2(n10381), .A(n6956), .ZN(P2_U3225) );
  XNOR2_X1 U8820 ( .A(n7856), .B(n7008), .ZN(n7055) );
  XNOR2_X1 U8821 ( .A(n7055), .B(n8285), .ZN(n6960) );
  AOI211_X1 U8822 ( .C1(n6960), .C2(n6959), .A(n8251), .B(n7057), .ZN(n6961)
         );
  INV_X1 U8823 ( .A(n6961), .ZN(n6965) );
  OAI22_X1 U8824 ( .A1(n6043), .A2(n8260), .B1(n8246), .B2(n7058), .ZN(n6962)
         );
  AOI211_X1 U8825 ( .C1(n10398), .C2(n8237), .A(n6963), .B(n6962), .ZN(n6964)
         );
  OAI211_X1 U8826 ( .C1(n7007), .C2(n8210), .A(n6965), .B(n6964), .ZN(P2_U3179) );
  AOI21_X1 U8827 ( .B1(n6968), .B2(n6967), .A(n6966), .ZN(n6971) );
  INV_X1 U8828 ( .A(n6969), .ZN(n6970) );
  OAI21_X1 U8829 ( .B1(n6993), .B2(n6971), .A(n6970), .ZN(n6976) );
  AOI21_X1 U8830 ( .B1(n6973), .B2(n6972), .A(n4585), .ZN(n6974) );
  NOR2_X1 U8831 ( .A1(n7025), .A2(n6974), .ZN(n6975) );
  AOI211_X1 U8832 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n10339), .A(n6976), .B(
        n6975), .ZN(n6983) );
  INV_X1 U8833 ( .A(n6977), .ZN(n6981) );
  INV_X1 U8834 ( .A(n10354), .ZN(n10206) );
  OAI21_X1 U8835 ( .B1(n6989), .B2(n6979), .A(n6978), .ZN(n6980) );
  NAND3_X1 U8836 ( .A1(n6981), .A2(n10206), .A3(n6980), .ZN(n6982) );
  OAI211_X1 U8837 ( .C1(n9945), .C2(n6984), .A(n6983), .B(n6982), .ZN(P2_U3186) );
  XOR2_X1 U8838 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6985), .Z(n6988) );
  INV_X1 U8839 ( .A(n6986), .ZN(n6987) );
  OAI21_X1 U8840 ( .B1(n7025), .B2(n6988), .A(n6987), .ZN(n6997) );
  AOI21_X1 U8841 ( .B1(n6991), .B2(n6990), .A(n6989), .ZN(n6995) );
  XOR2_X1 U8842 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6992), .Z(n6994) );
  OAI22_X1 U8843 ( .A1(n6995), .A2(n10354), .B1(n6994), .B2(n6993), .ZN(n6996)
         );
  AOI211_X1 U8844 ( .C1(n10339), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n6997), .B(
        n6996), .ZN(n6998) );
  OAI21_X1 U8845 ( .B1(n6999), .B2(n9945), .A(n6998), .ZN(P2_U3185) );
  NAND2_X1 U8846 ( .A1(n7001), .A2(n7000), .ZN(n7002) );
  XNOR2_X1 U8847 ( .A(n10398), .B(n8285), .ZN(n7915) );
  XNOR2_X1 U8848 ( .A(n7002), .B(n7915), .ZN(n7003) );
  AOI222_X1 U8849 ( .A1(n8430), .A2(n7003), .B1(n8284), .B2(n6321), .C1(n8286), 
        .C2(n8427), .ZN(n10401) );
  NAND2_X1 U8850 ( .A1(n7004), .A2(n7994), .ZN(n7005) );
  XNOR2_X1 U8851 ( .A(n7005), .B(n7915), .ZN(n10399) );
  NOR2_X1 U8852 ( .A1(n4495), .A2(n7006), .ZN(n7010) );
  OAI22_X1 U8853 ( .A1(n10365), .A2(n7008), .B1(n7007), .B2(n10373), .ZN(n7009) );
  AOI211_X1 U8854 ( .C1(n10399), .C2(n8438), .A(n7010), .B(n7009), .ZN(n7011)
         );
  OAI21_X1 U8855 ( .B1(n10401), .B2(n10381), .A(n7011), .ZN(P2_U3227) );
  NAND2_X1 U8856 ( .A1(n7013), .A2(n7012), .ZN(n7014) );
  XOR2_X1 U8857 ( .A(n7911), .B(n7014), .Z(n7015) );
  AOI222_X1 U8858 ( .A1(n8430), .A2(n7015), .B1(n8287), .B2(n6321), .C1(n8289), 
        .C2(n8427), .ZN(n10393) );
  XNOR2_X1 U8859 ( .A(n7016), .B(n7911), .ZN(n10391) );
  NOR2_X1 U8860 ( .A1(n4495), .A2(n6004), .ZN(n7019) );
  OAI22_X1 U8861 ( .A1(n10365), .A2(n7017), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n10373), .ZN(n7018) );
  AOI211_X1 U8862 ( .C1(n10391), .C2(n8438), .A(n7019), .B(n7018), .ZN(n7020)
         );
  OAI21_X1 U8863 ( .B1(n10381), .B2(n10393), .A(n7020), .ZN(P2_U3230) );
  XOR2_X1 U8864 ( .A(n7022), .B(n7021), .Z(n7024) );
  NAND2_X1 U8865 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(P2_U3151), .ZN(n7023) );
  OAI21_X1 U8866 ( .B1(n7025), .B2(n7024), .A(n7023), .ZN(n7026) );
  AOI21_X1 U8867 ( .B1(n10339), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n7026), .ZN(
        n7035) );
  OAI21_X1 U8868 ( .B1(n7029), .B2(n7028), .A(n7027), .ZN(n7033) );
  XOR2_X1 U8869 ( .A(n7031), .B(n7030), .Z(n7032) );
  AOI22_X1 U8870 ( .A1(n10348), .A2(n7033), .B1(n10206), .B2(n7032), .ZN(n7034) );
  OAI211_X1 U8871 ( .C1(n7036), .C2(n9945), .A(n7035), .B(n7034), .ZN(P2_U3184) );
  INV_X1 U8872 ( .A(n7313), .ZN(n7050) );
  INV_X1 U8873 ( .A(n7037), .ZN(n7038) );
  NAND2_X1 U8874 ( .A1(n7039), .A2(n7038), .ZN(n7042) );
  AND2_X1 U8875 ( .A1(n7044), .A2(n7042), .ZN(n7046) );
  OAI22_X1 U8876 ( .A1(n5524), .A2(n4503), .B1(n10125), .B2(n8728), .ZN(n7209)
         );
  OAI22_X1 U8877 ( .A1(n5524), .A2(n8728), .B1(n10125), .B2(n8609), .ZN(n7041)
         );
  XNOR2_X1 U8878 ( .A(n7041), .B(n7517), .ZN(n7208) );
  XOR2_X1 U8879 ( .A(n7209), .B(n7208), .Z(n7045) );
  AND2_X1 U8880 ( .A1(n7045), .A2(n7042), .ZN(n7043) );
  OAI211_X1 U8881 ( .C1(n7046), .C2(n7045), .A(n9966), .B(n7212), .ZN(n7049)
         );
  AOI22_X1 U8882 ( .A1(n9197), .A2(n9516), .B1(n9514), .B2(n9184), .ZN(n7308)
         );
  NAND2_X1 U8883 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n10029) );
  OAI21_X1 U8884 ( .B1(n7308), .B2(n9214), .A(n10029), .ZN(n7047) );
  AOI21_X1 U8885 ( .B1(n7314), .B2(n9217), .A(n7047), .ZN(n7048) );
  OAI211_X1 U8886 ( .C1(n9970), .C2(n7050), .A(n7049), .B(n7048), .ZN(P1_U3230) );
  INV_X1 U8887 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7052) );
  INV_X1 U8888 ( .A(n7051), .ZN(n7053) );
  OAI222_X1 U8889 ( .A1(n8551), .A2(n7052), .B1(n8555), .B2(n7053), .C1(n4914), 
        .C2(P2_U3151), .ZN(P2_U3277) );
  INV_X1 U8890 ( .A(n9587), .ZN(n7054) );
  INV_X1 U8891 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n9025) );
  OAI222_X1 U8892 ( .A1(P1_U3086), .A2(n7054), .B1(n4496), .B2(n7053), .C1(
        n9025), .C2(n7819), .ZN(P1_U3337) );
  AND2_X1 U8893 ( .A1(n7055), .A2(n8285), .ZN(n7056) );
  OAI21_X1 U8894 ( .B1(n7060), .B2(n7059), .A(n7110), .ZN(n7061) );
  NAND2_X1 U8895 ( .A1(n7061), .A2(n8242), .ZN(n7066) );
  INV_X1 U8896 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7062) );
  NOR2_X1 U8897 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7062), .ZN(n7086) );
  OAI22_X1 U8898 ( .A1(n7152), .A2(n8246), .B1(n8260), .B2(n7063), .ZN(n7064)
         );
  AOI211_X1 U8899 ( .C1(n10406), .C2(n8237), .A(n7086), .B(n7064), .ZN(n7065)
         );
  OAI211_X1 U8900 ( .C1(n7104), .C2(n8210), .A(n7066), .B(n7065), .ZN(P2_U3153) );
  XNOR2_X1 U8901 ( .A(n7123), .B(P1_REG2_REG_11__SCAN_IN), .ZN(n7068) );
  AOI211_X1 U8902 ( .C1(n7069), .C2(n7068), .A(n7119), .B(n10018), .ZN(n7080)
         );
  INV_X1 U8903 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7072) );
  MUX2_X1 U8904 ( .A(n7072), .B(P1_REG1_REG_11__SCAN_IN), .S(n7123), .Z(n7073)
         );
  AOI211_X1 U8905 ( .C1(n7074), .C2(n7073), .A(n7125), .B(n9993), .ZN(n7079)
         );
  INV_X1 U8906 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7077) );
  NAND2_X1 U8907 ( .A1(n10025), .A2(n7123), .ZN(n7076) );
  NAND2_X1 U8908 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n7075) );
  OAI211_X1 U8909 ( .C1(n7077), .C2(n9601), .A(n7076), .B(n7075), .ZN(n7078)
         );
  OR3_X1 U8910 ( .A1(n7080), .A2(n7079), .A3(n7078), .ZN(P1_U3254) );
  AOI21_X1 U8911 ( .B1(n7083), .B2(n7082), .A(n7081), .ZN(n7095) );
  NOR2_X1 U8912 ( .A1(n9945), .A2(n7084), .ZN(n7085) );
  AOI211_X1 U8913 ( .C1(n10339), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n7086), .B(
        n7085), .ZN(n7094) );
  OAI21_X1 U8914 ( .B1(P2_REG1_REG_7__SCAN_IN), .B2(n7088), .A(n7087), .ZN(
        n7092) );
  OAI21_X1 U8915 ( .B1(n7090), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7089), .ZN(
        n7091) );
  AOI22_X1 U8916 ( .A1(n7092), .A2(n10347), .B1(n10348), .B2(n7091), .ZN(n7093) );
  OAI211_X1 U8917 ( .C1(n7095), .C2(n10354), .A(n7094), .B(n7093), .ZN(
        P2_U3189) );
  OR2_X1 U8918 ( .A1(n7096), .A2(n8001), .ZN(n7097) );
  NAND2_X1 U8919 ( .A1(n7098), .A2(n7097), .ZN(n10403) );
  XNOR2_X1 U8920 ( .A(n7099), .B(n8001), .ZN(n7100) );
  NAND2_X1 U8921 ( .A1(n7100), .A2(n8430), .ZN(n7102) );
  AOI22_X1 U8922 ( .A1(n8285), .A2(n8427), .B1(n6321), .B2(n8282), .ZN(n7101)
         );
  OAI211_X1 U8923 ( .C1(n10403), .C2(n7200), .A(n7102), .B(n7101), .ZN(n10404)
         );
  MUX2_X1 U8924 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10404), .S(n4495), .Z(n7103)
         );
  INV_X1 U8925 ( .A(n7103), .ZN(n7107) );
  INV_X1 U8926 ( .A(n7104), .ZN(n7105) );
  AOI22_X1 U8927 ( .A1(n8434), .A2(n10406), .B1(n8404), .B2(n7105), .ZN(n7106)
         );
  OAI211_X1 U8928 ( .C1(n10403), .C2(n7811), .A(n7107), .B(n7106), .ZN(
        P2_U3226) );
  XNOR2_X1 U8929 ( .A(n7856), .B(n7114), .ZN(n7151) );
  XNOR2_X1 U8930 ( .A(n7151), .B(n7152), .ZN(n7154) );
  XOR2_X1 U8931 ( .A(n7155), .B(n7154), .Z(n7118) );
  AOI21_X1 U8932 ( .B1(n8244), .B2(n8284), .A(n7111), .ZN(n7113) );
  NAND2_X1 U8933 ( .A1(n8257), .A2(n8281), .ZN(n7112) );
  OAI211_X1 U8934 ( .C1(n7114), .C2(n8266), .A(n7113), .B(n7112), .ZN(n7115)
         );
  AOI21_X1 U8935 ( .B1(n7116), .B2(n8262), .A(n7115), .ZN(n7117) );
  OAI21_X1 U8936 ( .B1(n7118), .B2(n8251), .A(n7117), .ZN(P2_U3161) );
  NOR2_X1 U8937 ( .A1(n7374), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7120) );
  AOI21_X1 U8938 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7374), .A(n7120), .ZN(
        n7121) );
  OAI21_X1 U8939 ( .B1(n7122), .B2(n7121), .A(n7369), .ZN(n7134) );
  AND2_X1 U8940 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9959) );
  AOI21_X1 U8941 ( .B1(n10026), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n9959), .ZN(
        n7130) );
  AND2_X1 U8942 ( .A1(n7123), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7124) );
  INV_X1 U8943 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7581) );
  AOI22_X1 U8944 ( .A1(n7374), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n7581), .B2(
        n7131), .ZN(n7126) );
  OAI21_X1 U8945 ( .B1(n7127), .B2(n7126), .A(n7373), .ZN(n7128) );
  NAND2_X1 U8946 ( .A1(n10017), .A2(n7128), .ZN(n7129) );
  OAI211_X1 U8947 ( .C1(n7132), .C2(n7131), .A(n7130), .B(n7129), .ZN(n7133)
         );
  AOI21_X1 U8948 ( .B1(n9593), .B2(n7134), .A(n7133), .ZN(n7135) );
  INV_X1 U8949 ( .A(n7135), .ZN(P1_U3255) );
  INV_X1 U8950 ( .A(n7136), .ZN(n7139) );
  OAI222_X1 U8951 ( .A1(n7819), .A2(n7137), .B1(n4496), .B2(n7139), .C1(
        P1_U3086), .C2(n9720), .ZN(P1_U3336) );
  OAI222_X1 U8952 ( .A1(n8551), .A2(n8883), .B1(n8555), .B2(n7139), .C1(n7138), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  OR2_X1 U8953 ( .A1(n6950), .A2(n7953), .ZN(n7141) );
  AND2_X1 U8954 ( .A1(n7141), .A2(n7140), .ZN(n7143) );
  INV_X1 U8955 ( .A(n7142), .ZN(n8004) );
  XNOR2_X1 U8956 ( .A(n7143), .B(n7921), .ZN(n10421) );
  XOR2_X1 U8957 ( .A(n7144), .B(n7921), .Z(n7145) );
  NAND2_X1 U8958 ( .A1(n7145), .A2(n8430), .ZN(n7147) );
  AOI22_X1 U8959 ( .A1(n8427), .A2(n8281), .B1(n8279), .B2(n6321), .ZN(n7146)
         );
  OAI211_X1 U8960 ( .C1(n10421), .C2(n7200), .A(n7147), .B(n7146), .ZN(n10423)
         );
  NAND2_X1 U8961 ( .A1(n10423), .A2(n4495), .ZN(n7150) );
  OAI22_X1 U8962 ( .A1(n4495), .A2(n5867), .B1(n7430), .B2(n10373), .ZN(n7148)
         );
  AOI21_X1 U8963 ( .B1(n8419), .B2(n7432), .A(n7148), .ZN(n7149) );
  OAI211_X1 U8964 ( .C1(n10421), .C2(n7811), .A(n7150), .B(n7149), .ZN(
        P2_U3223) );
  INV_X1 U8965 ( .A(n7151), .ZN(n7153) );
  XNOR2_X1 U8966 ( .A(n10416), .B(n7856), .ZN(n7425) );
  XOR2_X1 U8967 ( .A(n7426), .B(n7425), .Z(n7156) );
  OAI211_X1 U8968 ( .C1(n7157), .C2(n7156), .A(n7424), .B(n8242), .ZN(n7163)
         );
  NOR2_X1 U8969 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7158), .ZN(n10216) );
  AOI21_X1 U8970 ( .B1(n8244), .B2(n8282), .A(n10216), .ZN(n7160) );
  NAND2_X1 U8971 ( .A1(n8257), .A2(n8280), .ZN(n7159) );
  OAI211_X1 U8972 ( .C1(n8210), .C2(n7201), .A(n7160), .B(n7159), .ZN(n7161)
         );
  AOI21_X1 U8973 ( .B1(n10416), .B2(n8237), .A(n7161), .ZN(n7162) );
  NAND2_X1 U8974 ( .A1(n7163), .A2(n7162), .ZN(P2_U3171) );
  INV_X2 U8975 ( .A(n10056), .ZN(n10042) );
  AND3_X1 U8976 ( .A1(n9336), .A2(n9473), .A3(n7164), .ZN(n7165) );
  AOI211_X1 U8977 ( .C1(n10042), .C2(P1_REG3_REG_0__SCAN_IN), .A(n7166), .B(
        n7165), .ZN(n7175) );
  INV_X1 U8978 ( .A(n7167), .ZN(n7169) );
  NAND3_X1 U8979 ( .A1(n7169), .A2(n9475), .A3(n7168), .ZN(n7170) );
  OAI21_X1 U8980 ( .B1(n9611), .B2(n9794), .A(n9800), .ZN(n7173) );
  AOI22_X1 U8981 ( .A1(n7173), .A2(n7172), .B1(n10043), .B2(
        P1_REG2_REG_0__SCAN_IN), .ZN(n7174) );
  OAI21_X1 U8982 ( .B1(n7175), .B2(n10043), .A(n7174), .ZN(P1_U3293) );
  OR2_X1 U8983 ( .A1(n6950), .A2(n7176), .ZN(n7178) );
  AND2_X1 U8984 ( .A1(n7178), .A2(n7177), .ZN(n7179) );
  NAND2_X1 U8985 ( .A1(n7179), .A2(n7950), .ZN(n7180) );
  XNOR2_X1 U8986 ( .A(n7180), .B(n7183), .ZN(n10425) );
  NAND2_X1 U8987 ( .A1(n7182), .A2(n7181), .ZN(n7184) );
  XNOR2_X1 U8988 ( .A(n7184), .B(n7183), .ZN(n7185) );
  OAI222_X1 U8989 ( .A1(n8391), .A2(n7457), .B1(n8389), .B2(n7749), .C1(n7185), 
        .C2(n8387), .ZN(n10426) );
  NAND2_X1 U8990 ( .A1(n10426), .A2(n4495), .ZN(n7189) );
  OAI22_X1 U8991 ( .A1(n4495), .A2(n7186), .B1(n7464), .B2(n10373), .ZN(n7187)
         );
  AOI21_X1 U8992 ( .B1(n8434), .B2(n10428), .A(n7187), .ZN(n7188) );
  OAI211_X1 U8993 ( .C1(n8407), .C2(n10425), .A(n7189), .B(n7188), .ZN(
        P2_U3222) );
  OR2_X1 U8994 ( .A1(n6950), .A2(n7190), .ZN(n7192) );
  AND2_X1 U8995 ( .A1(n7192), .A2(n7949), .ZN(n7195) );
  NAND2_X1 U8996 ( .A1(n7192), .A2(n7191), .ZN(n7193) );
  OAI21_X1 U8997 ( .B1(n7195), .B2(n7194), .A(n7193), .ZN(n10413) );
  XOR2_X1 U8998 ( .A(n7918), .B(n7196), .Z(n7197) );
  NAND2_X1 U8999 ( .A1(n7197), .A2(n8430), .ZN(n7199) );
  AOI22_X1 U9000 ( .A1(n8427), .A2(n8282), .B1(n8280), .B2(n6321), .ZN(n7198)
         );
  OAI211_X1 U9001 ( .C1(n7200), .C2(n10413), .A(n7199), .B(n7198), .ZN(n10414)
         );
  NAND2_X1 U9002 ( .A1(n10414), .A2(n4495), .ZN(n7205) );
  OAI22_X1 U9003 ( .A1(n4495), .A2(n7202), .B1(n7201), .B2(n10373), .ZN(n7203)
         );
  AOI21_X1 U9004 ( .B1(n8419), .B2(n10416), .A(n7203), .ZN(n7204) );
  OAI211_X1 U9005 ( .C1(n10413), .C2(n7811), .A(n7205), .B(n7204), .ZN(
        P2_U3224) );
  OR2_X1 U9006 ( .A1(n7326), .A2(n4503), .ZN(n7207) );
  NAND2_X1 U9007 ( .A1(n7298), .A2(n8733), .ZN(n7206) );
  NAND2_X1 U9008 ( .A1(n7207), .A2(n7206), .ZN(n7230) );
  INV_X1 U9009 ( .A(n7208), .ZN(n7211) );
  INV_X1 U9010 ( .A(n7209), .ZN(n7210) );
  OAI22_X1 U9011 ( .A1(n7326), .A2(n8728), .B1(n10132), .B2(n8609), .ZN(n7213)
         );
  XNOR2_X1 U9012 ( .A(n7213), .B(n7517), .ZN(n7231) );
  INV_X1 U9013 ( .A(n7231), .ZN(n7214) );
  NAND2_X1 U9014 ( .A1(n4580), .A2(n7214), .ZN(n7320) );
  OAI21_X1 U9015 ( .B1(n4580), .B2(n7214), .A(n7320), .ZN(n7215) );
  NOR2_X1 U9016 ( .A1(n7215), .A2(n7230), .ZN(n7323) );
  AOI21_X1 U9017 ( .B1(n7230), .B2(n7215), .A(n7323), .ZN(n7222) );
  OR2_X1 U9018 ( .A1(n5524), .A2(n9141), .ZN(n7217) );
  OR2_X1 U9019 ( .A1(n7246), .A2(n9195), .ZN(n7216) );
  NAND2_X1 U9020 ( .A1(n7217), .A2(n7216), .ZN(n7293) );
  NAND2_X1 U9021 ( .A1(n7293), .A2(n9960), .ZN(n7218) );
  OAI211_X1 U9022 ( .C1(n9963), .C2(n10132), .A(n7219), .B(n7218), .ZN(n7220)
         );
  AOI21_X1 U9023 ( .B1(n7297), .B2(n9211), .A(n7220), .ZN(n7221) );
  OAI21_X1 U9024 ( .B1(n7222), .B2(n9220), .A(n7221), .ZN(P1_U3227) );
  INV_X1 U9025 ( .A(n7223), .ZN(n7260) );
  OAI222_X1 U9026 ( .A1(P1_U3086), .A2(n7225), .B1(n4496), .B2(n7260), .C1(
        n7224), .C2(n7819), .ZN(P1_U3335) );
  OR2_X1 U9027 ( .A1(n7231), .A2(n7230), .ZN(n7226) );
  OAI22_X1 U9028 ( .A1(n7246), .A2(n8728), .B1(n10138), .B2(n8609), .ZN(n7227)
         );
  XNOR2_X1 U9029 ( .A(n7227), .B(n8731), .ZN(n7235) );
  OR2_X1 U9030 ( .A1(n7246), .A2(n4503), .ZN(n7229) );
  NAND2_X1 U9031 ( .A1(n7361), .A2(n8733), .ZN(n7228) );
  NAND2_X1 U9032 ( .A1(n7229), .A2(n7228), .ZN(n7236) );
  XNOR2_X1 U9033 ( .A(n7235), .B(n7236), .ZN(n7322) );
  NAND2_X1 U9034 ( .A1(n7231), .A2(n7230), .ZN(n7232) );
  INV_X1 U9035 ( .A(n7236), .ZN(n7237) );
  NAND2_X1 U9036 ( .A1(n7235), .A2(n7237), .ZN(n7238) );
  OAI22_X1 U9037 ( .A1(n7339), .A2(n8728), .B1(n10145), .B2(n8609), .ZN(n7239)
         );
  XNOR2_X1 U9038 ( .A(n7239), .B(n4493), .ZN(n7243) );
  OR2_X1 U9039 ( .A1(n7339), .A2(n4503), .ZN(n7241) );
  NAND2_X1 U9040 ( .A1(n10044), .A2(n8733), .ZN(n7240) );
  NAND2_X1 U9041 ( .A1(n7241), .A2(n7240), .ZN(n7242) );
  NOR2_X1 U9042 ( .A1(n7243), .A2(n7242), .ZN(n7514) );
  INV_X1 U9043 ( .A(n7514), .ZN(n7244) );
  NAND2_X1 U9044 ( .A1(n7243), .A2(n7242), .ZN(n7513) );
  NAND2_X1 U9045 ( .A1(n7244), .A2(n7513), .ZN(n7245) );
  XNOR2_X1 U9046 ( .A(n7515), .B(n7245), .ZN(n7250) );
  OAI22_X1 U9047 ( .A1(n7516), .A2(n9195), .B1(n7246), .B2(n9141), .ZN(n10040)
         );
  AOI22_X1 U9048 ( .A1(n10040), .A2(n9960), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3086), .ZN(n7247) );
  OAI21_X1 U9049 ( .B1(n10145), .B2(n9963), .A(n7247), .ZN(n7248) );
  AOI21_X1 U9050 ( .B1(n10041), .B2(n9211), .A(n7248), .ZN(n7249) );
  OAI21_X1 U9051 ( .B1(n7250), .B2(n9220), .A(n7249), .ZN(P1_U3213) );
  OR2_X1 U9052 ( .A1(n7251), .A2(n7923), .ZN(n7253) );
  INV_X1 U9053 ( .A(n7285), .ZN(n7259) );
  INV_X1 U9054 ( .A(n7923), .ZN(n8018) );
  XNOR2_X1 U9055 ( .A(n7254), .B(n8018), .ZN(n7255) );
  OAI222_X1 U9056 ( .A1(n8391), .A2(n7558), .B1(n8389), .B2(n8020), .C1(n7255), 
        .C2(n8387), .ZN(n7283) );
  NAND2_X1 U9057 ( .A1(n7283), .A2(n4495), .ZN(n7258) );
  OAI22_X1 U9058 ( .A1(n4495), .A2(n5874), .B1(n7566), .B2(n10373), .ZN(n7256)
         );
  AOI21_X1 U9059 ( .B1(n8434), .B2(n7568), .A(n7256), .ZN(n7257) );
  OAI211_X1 U9060 ( .C1(n7259), .C2(n8407), .A(n7258), .B(n7257), .ZN(P2_U3221) );
  OAI222_X1 U9061 ( .A1(n8551), .A2(n8894), .B1(P2_U3151), .B2(n7261), .C1(
        n8562), .C2(n7260), .ZN(P2_U3275) );
  XOR2_X1 U9062 ( .A(n7304), .B(n7262), .Z(n7264) );
  AOI21_X1 U9063 ( .B1(n7264), .B2(n10054), .A(n7263), .ZN(n10112) );
  AND2_X1 U9064 ( .A1(n10031), .A2(n10045), .ZN(n7265) );
  XNOR2_X1 U9065 ( .A(n7266), .B(n7262), .ZN(n10115) );
  NAND2_X1 U9066 ( .A1(n10110), .A2(n10066), .ZN(n7268) );
  AOI22_X1 U9067 ( .A1(n10070), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n10042), .ZN(n7267) );
  OAI211_X1 U9068 ( .C1(n5507), .C2(n9800), .A(n7268), .B(n7267), .ZN(n7269)
         );
  AOI21_X1 U9069 ( .B1(n10067), .B2(n10115), .A(n7269), .ZN(n7270) );
  OAI21_X1 U9070 ( .B1(n10043), .B2(n10112), .A(n7270), .ZN(P1_U3291) );
  XNOR2_X1 U9071 ( .A(n9337), .B(n7271), .ZN(n7273) );
  AOI21_X1 U9072 ( .B1(n7273), .B2(n10054), .A(n7272), .ZN(n10105) );
  OAI211_X1 U9073 ( .C1(n7275), .C2(n10104), .A(n10063), .B(n7274), .ZN(n10103) );
  NOR2_X1 U9074 ( .A1(n9611), .A2(n10103), .ZN(n7278) );
  INV_X1 U9075 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7276) );
  OAI22_X1 U9076 ( .A1(n10058), .A2(n6393), .B1(n7276), .B2(n10056), .ZN(n7277) );
  AOI211_X1 U9077 ( .C1(n10060), .C2(n7279), .A(n7278), .B(n7277), .ZN(n7282)
         );
  XNOR2_X1 U9078 ( .A(n7280), .B(n5728), .ZN(n10108) );
  NAND2_X1 U9079 ( .A1(n10108), .A2(n10067), .ZN(n7281) );
  OAI211_X1 U9080 ( .C1(n10070), .C2(n10105), .A(n7282), .B(n7281), .ZN(
        P1_U3292) );
  AOI21_X1 U9081 ( .B1(n10429), .B2(n7568), .A(n7283), .ZN(n7287) );
  INV_X1 U9082 ( .A(n8544), .ZN(n7418) );
  AOI22_X1 U9083 ( .A1(n7285), .A2(n7418), .B1(P2_REG0_REG_12__SCAN_IN), .B2(
        n10432), .ZN(n7284) );
  OAI21_X1 U9084 ( .B1(n7287), .B2(n10432), .A(n7284), .ZN(P2_U3426) );
  AOI22_X1 U9085 ( .A1(n7285), .A2(n6369), .B1(P2_REG1_REG_12__SCAN_IN), .B2(
        n10444), .ZN(n7286) );
  OAI21_X1 U9086 ( .B1(n7287), .B2(n10444), .A(n7286), .ZN(P2_U3471) );
  XNOR2_X1 U9087 ( .A(n7288), .B(n9335), .ZN(n10130) );
  INV_X1 U9088 ( .A(n10130), .ZN(n7303) );
  OAI21_X1 U9089 ( .B1(n7291), .B2(n7289), .A(n7290), .ZN(n7292) );
  NAND2_X1 U9090 ( .A1(n7292), .A2(n10054), .ZN(n7295) );
  INV_X1 U9091 ( .A(n7293), .ZN(n7294) );
  NAND2_X1 U9092 ( .A1(n7295), .A2(n7294), .ZN(n10135) );
  AOI21_X1 U9093 ( .B1(n7312), .B2(n7298), .A(n9794), .ZN(n7296) );
  NAND2_X1 U9094 ( .A1(n7296), .A2(n7357), .ZN(n10131) );
  AOI22_X1 U9095 ( .A1(n10070), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7297), .B2(
        n10042), .ZN(n7300) );
  NAND2_X1 U9096 ( .A1(n10060), .A2(n7298), .ZN(n7299) );
  OAI211_X1 U9097 ( .C1(n10131), .C2(n9611), .A(n7300), .B(n7299), .ZN(n7301)
         );
  AOI21_X1 U9098 ( .B1(n10135), .B2(n10058), .A(n7301), .ZN(n7302) );
  OAI21_X1 U9099 ( .B1(n7303), .B2(n9803), .A(n7302), .ZN(P1_U3288) );
  INV_X1 U9100 ( .A(n7304), .ZN(n7306) );
  NAND2_X1 U9101 ( .A1(n7306), .A2(n5732), .ZN(n9388) );
  NAND2_X1 U9102 ( .A1(n9388), .A2(n9385), .ZN(n10052) );
  OAI21_X1 U9103 ( .B1(n10052), .B2(n10062), .A(n9389), .ZN(n7307) );
  XNOR2_X1 U9104 ( .A(n9334), .B(n7307), .ZN(n7309) );
  OAI21_X1 U9105 ( .B1(n7309), .B2(n10036), .A(n7308), .ZN(n10126) );
  INV_X1 U9106 ( .A(n10126), .ZN(n7319) );
  XNOR2_X1 U9107 ( .A(n7310), .B(n9334), .ZN(n10128) );
  OAI211_X1 U9108 ( .C1(n5162), .C2(n10125), .A(n10063), .B(n7312), .ZN(n10124) );
  AOI22_X1 U9109 ( .A1(n10070), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7313), .B2(
        n10042), .ZN(n7316) );
  NAND2_X1 U9110 ( .A1(n10060), .A2(n7314), .ZN(n7315) );
  OAI211_X1 U9111 ( .C1(n10124), .C2(n9611), .A(n7316), .B(n7315), .ZN(n7317)
         );
  AOI21_X1 U9112 ( .B1(n10128), .B2(n10067), .A(n7317), .ZN(n7318) );
  OAI21_X1 U9113 ( .B1(n7319), .B2(n10070), .A(n7318), .ZN(P1_U3289) );
  INV_X1 U9114 ( .A(n7320), .ZN(n7321) );
  OR3_X1 U9115 ( .A1(n7323), .A2(n7322), .A3(n7321), .ZN(n7325) );
  AOI21_X1 U9116 ( .B1(n7325), .B2(n7324), .A(n9220), .ZN(n7335) );
  INV_X1 U9117 ( .A(n7360), .ZN(n7333) );
  OR2_X1 U9118 ( .A1(n7339), .A2(n9195), .ZN(n7328) );
  OR2_X1 U9119 ( .A1(n7326), .A2(n9141), .ZN(n7327) );
  NAND2_X1 U9120 ( .A1(n7328), .A2(n7327), .ZN(n7352) );
  INV_X1 U9121 ( .A(n7329), .ZN(n7330) );
  AOI21_X1 U9122 ( .B1(n7352), .B2(n9960), .A(n7330), .ZN(n7332) );
  NAND2_X1 U9123 ( .A1(n9217), .A2(n7361), .ZN(n7331) );
  OAI211_X1 U9124 ( .C1(n9970), .C2(n7333), .A(n7332), .B(n7331), .ZN(n7334)
         );
  OR2_X1 U9125 ( .A1(n7335), .A2(n7334), .ZN(P1_U3239) );
  NAND2_X1 U9126 ( .A1(n7351), .A2(n9223), .ZN(n10035) );
  NAND2_X1 U9127 ( .A1(n10035), .A2(n10034), .ZN(n7336) );
  NAND2_X1 U9128 ( .A1(n7336), .A2(n4783), .ZN(n10038) );
  AOI21_X1 U9129 ( .B1(n10038), .B2(n7337), .A(n7344), .ZN(n7400) );
  AND3_X1 U9130 ( .A1(n10038), .A2(n7337), .A3(n7344), .ZN(n7338) );
  OAI21_X1 U9131 ( .B1(n7400), .B2(n7338), .A(n10054), .ZN(n7342) );
  OR2_X1 U9132 ( .A1(n7339), .A2(n9141), .ZN(n7341) );
  OR2_X1 U9133 ( .A1(n7597), .A2(n9195), .ZN(n7340) );
  AND2_X1 U9134 ( .A1(n7341), .A2(n7340), .ZN(n7522) );
  NAND2_X1 U9135 ( .A1(n7342), .A2(n7522), .ZN(n10158) );
  INV_X1 U9136 ( .A(n10158), .ZN(n7350) );
  XNOR2_X1 U9137 ( .A(n7343), .B(n7344), .ZN(n10152) );
  AOI21_X1 U9138 ( .B1(n10046), .B2(n7510), .A(n9794), .ZN(n7345) );
  NAND2_X1 U9139 ( .A1(n7345), .A2(n5080), .ZN(n10151) );
  AOI22_X1 U9140 ( .A1(n10070), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7524), .B2(
        n10042), .ZN(n7347) );
  NAND2_X1 U9141 ( .A1(n10060), .A2(n7510), .ZN(n7346) );
  OAI211_X1 U9142 ( .C1(n10151), .C2(n9611), .A(n7347), .B(n7346), .ZN(n7348)
         );
  AOI21_X1 U9143 ( .B1(n10152), .B2(n10067), .A(n7348), .ZN(n7349) );
  OAI21_X1 U9144 ( .B1(n7350), .B2(n10070), .A(n7349), .ZN(P1_U3285) );
  XNOR2_X1 U9145 ( .A(n7351), .B(n7356), .ZN(n7354) );
  INV_X1 U9146 ( .A(n7352), .ZN(n7353) );
  OAI21_X1 U9147 ( .B1(n7354), .B2(n10036), .A(n7353), .ZN(n10139) );
  INV_X1 U9148 ( .A(n10139), .ZN(n7366) );
  XNOR2_X1 U9149 ( .A(n7355), .B(n7356), .ZN(n10141) );
  INV_X1 U9150 ( .A(n7357), .ZN(n7359) );
  INV_X1 U9151 ( .A(n10047), .ZN(n7358) );
  OAI211_X1 U9152 ( .C1(n10138), .C2(n7359), .A(n7358), .B(n10063), .ZN(n10137) );
  AOI22_X1 U9153 ( .A1(n10043), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7360), .B2(
        n10042), .ZN(n7363) );
  NAND2_X1 U9154 ( .A1(n10060), .A2(n7361), .ZN(n7362) );
  OAI211_X1 U9155 ( .C1(n10137), .C2(n9611), .A(n7363), .B(n7362), .ZN(n7364)
         );
  AOI21_X1 U9156 ( .B1(n10141), .B2(n10067), .A(n7364), .ZN(n7365) );
  OAI21_X1 U9157 ( .B1(n7366), .B2(n10070), .A(n7365), .ZN(P1_U3287) );
  INV_X1 U9158 ( .A(n7367), .ZN(n7383) );
  OAI222_X1 U9159 ( .A1(P1_U3086), .A2(n9381), .B1(n4496), .B2(n7383), .C1(
        n7368), .C2(n7819), .ZN(P1_U3334) );
  OAI21_X1 U9160 ( .B1(n7374), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7369), .ZN(
        n7372) );
  NAND2_X1 U9161 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7482), .ZN(n7370) );
  OAI21_X1 U9162 ( .B1(n7482), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7370), .ZN(
        n7371) );
  NOR2_X1 U9163 ( .A1(n7371), .A2(n7372), .ZN(n7477) );
  AOI211_X1 U9164 ( .C1(n7372), .C2(n7371), .A(n7477), .B(n10018), .ZN(n7382)
         );
  OAI21_X1 U9165 ( .B1(n7374), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7373), .ZN(
        n7377) );
  INV_X1 U9166 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7375) );
  MUX2_X1 U9167 ( .A(n7375), .B(P1_REG1_REG_13__SCAN_IN), .S(n7482), .Z(n7376)
         );
  NOR2_X1 U9168 ( .A1(n7376), .A2(n7377), .ZN(n7481) );
  AOI211_X1 U9169 ( .C1(n7377), .C2(n7376), .A(n7481), .B(n9993), .ZN(n7381)
         );
  INV_X1 U9170 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7379) );
  NAND2_X1 U9171 ( .A1(n10025), .A2(n7482), .ZN(n7378) );
  NAND2_X1 U9172 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n7666) );
  OAI211_X1 U9173 ( .C1(n7379), .C2(n9601), .A(n7378), .B(n7666), .ZN(n7380)
         );
  OR3_X1 U9174 ( .A1(n7382), .A2(n7381), .A3(n7380), .ZN(P1_U3256) );
  OAI222_X1 U9175 ( .A1(n8551), .A2(n7384), .B1(P2_U3151), .B2(n7963), .C1(
        n8562), .C2(n7383), .ZN(P2_U3274) );
  AND2_X1 U9176 ( .A1(n7385), .A2(n9400), .ZN(n7388) );
  OAI21_X1 U9177 ( .B1(n7388), .B2(n7387), .A(n7386), .ZN(n7391) );
  OR2_X1 U9178 ( .A1(n7597), .A2(n9141), .ZN(n7390) );
  NAND2_X1 U9179 ( .A1(n9508), .A2(n9184), .ZN(n7389) );
  NAND2_X1 U9180 ( .A1(n7390), .A2(n7389), .ZN(n8704) );
  AOI21_X1 U9181 ( .B1(n7391), .B2(n10054), .A(n8704), .ZN(n10167) );
  OAI22_X1 U9182 ( .A1(n10058), .A2(n7392), .B1(n8706), .B2(n10056), .ZN(n7395) );
  INV_X1 U9183 ( .A(n7442), .ZN(n7393) );
  OAI211_X1 U9184 ( .C1(n10169), .C2(n7406), .A(n7393), .B(n10063), .ZN(n10166) );
  NOR2_X1 U9185 ( .A1(n10166), .A2(n9611), .ZN(n7394) );
  AOI211_X1 U9186 ( .C1(n10060), .C2(n8713), .A(n7395), .B(n7394), .ZN(n7398)
         );
  XNOR2_X1 U9187 ( .A(n7396), .B(n9342), .ZN(n10171) );
  NAND2_X1 U9188 ( .A1(n10171), .A2(n10067), .ZN(n7397) );
  OAI211_X1 U9189 ( .C1(n10070), .C2(n10167), .A(n7398), .B(n7397), .ZN(
        P1_U3283) );
  INV_X1 U9190 ( .A(n9236), .ZN(n7399) );
  NOR2_X1 U9191 ( .A1(n7400), .A2(n7399), .ZN(n7401) );
  XOR2_X1 U9192 ( .A(n7404), .B(n7401), .Z(n7402) );
  OR2_X1 U9193 ( .A1(n7516), .A2(n9141), .ZN(n7601) );
  OAI21_X1 U9194 ( .B1(n7402), .B2(n10036), .A(n7601), .ZN(n10162) );
  INV_X1 U9195 ( .A(n10162), .ZN(n7413) );
  XNOR2_X1 U9196 ( .A(n7403), .B(n7404), .ZN(n10164) );
  NAND2_X1 U9197 ( .A1(n5080), .A2(n7605), .ZN(n7405) );
  NAND2_X1 U9198 ( .A1(n7405), .A2(n10063), .ZN(n7407) );
  OR2_X1 U9199 ( .A1(n7407), .A2(n7406), .ZN(n7408) );
  OR2_X1 U9200 ( .A1(n7638), .A2(n9195), .ZN(n7602) );
  AND2_X1 U9201 ( .A1(n7408), .A2(n7602), .ZN(n10160) );
  AOI22_X1 U9202 ( .A1(n10043), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7600), .B2(
        n10042), .ZN(n7410) );
  NAND2_X1 U9203 ( .A1(n10060), .A2(n7605), .ZN(n7409) );
  OAI211_X1 U9204 ( .C1(n10160), .C2(n9611), .A(n7410), .B(n7409), .ZN(n7411)
         );
  AOI21_X1 U9205 ( .B1(n10164), .B2(n10067), .A(n7411), .ZN(n7412) );
  OAI21_X1 U9206 ( .B1(n7413), .B2(n10043), .A(n7412), .ZN(P1_U3284) );
  INV_X1 U9207 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7416) );
  XNOR2_X1 U9208 ( .A(n7414), .B(n7925), .ZN(n7415) );
  AOI222_X1 U9209 ( .A1(n8430), .A2(n7415), .B1(n8276), .B2(n6321), .C1(n8278), 
        .C2(n8427), .ZN(n7448) );
  MUX2_X1 U9210 ( .A(n7416), .B(n7448), .S(n10430), .Z(n7420) );
  XNOR2_X1 U9211 ( .A(n7417), .B(n7925), .ZN(n7451) );
  AOI22_X1 U9212 ( .A1(n7451), .A2(n7418), .B1(n8533), .B2(n8217), .ZN(n7419)
         );
  NAND2_X1 U9213 ( .A1(n7420), .A2(n7419), .ZN(P2_U3429) );
  MUX2_X1 U9214 ( .A(n7421), .B(n7448), .S(n10446), .Z(n7423) );
  AOI22_X1 U9215 ( .A1(n7451), .A2(n6369), .B1(n8473), .B2(n8217), .ZN(n7422)
         );
  NAND2_X1 U9216 ( .A1(n7423), .A2(n7422), .ZN(P2_U3472) );
  XNOR2_X1 U9217 ( .A(n7455), .B(n7457), .ZN(n7459) );
  XNOR2_X1 U9218 ( .A(n7432), .B(n7856), .ZN(n7458) );
  XOR2_X1 U9219 ( .A(n7459), .B(n7458), .Z(n7434) );
  NAND2_X1 U9220 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n10238) );
  INV_X1 U9221 ( .A(n10238), .ZN(n7427) );
  AOI21_X1 U9222 ( .B1(n8244), .B2(n8281), .A(n7427), .ZN(n7429) );
  NAND2_X1 U9223 ( .A1(n8257), .A2(n8279), .ZN(n7428) );
  OAI211_X1 U9224 ( .C1(n8210), .C2(n7430), .A(n7429), .B(n7428), .ZN(n7431)
         );
  AOI21_X1 U9225 ( .B1(n7432), .B2(n8237), .A(n7431), .ZN(n7433) );
  OAI21_X1 U9226 ( .B1(n7434), .B2(n8251), .A(n7433), .ZN(P2_U3157) );
  XNOR2_X1 U9227 ( .A(n7435), .B(n5741), .ZN(n7470) );
  AOI21_X1 U9228 ( .B1(n7437), .B2(n7436), .A(n10036), .ZN(n7440) );
  OR2_X1 U9229 ( .A1(n7655), .A2(n9195), .ZN(n7439) );
  OR2_X1 U9230 ( .A1(n7638), .A2(n9141), .ZN(n7438) );
  NAND2_X1 U9231 ( .A1(n7439), .A2(n7438), .ZN(n7692) );
  AOI21_X1 U9232 ( .B1(n7440), .B2(n7496), .A(n7692), .ZN(n7469) );
  INV_X1 U9233 ( .A(n7469), .ZN(n7446) );
  OAI211_X1 U9234 ( .C1(n7442), .C2(n7645), .A(n10063), .B(n7441), .ZN(n7468)
         );
  AOI22_X1 U9235 ( .A1(n10070), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7691), .B2(
        n10042), .ZN(n7444) );
  NAND2_X1 U9236 ( .A1(n10060), .A2(n7693), .ZN(n7443) );
  OAI211_X1 U9237 ( .C1(n7468), .C2(n9611), .A(n7444), .B(n7443), .ZN(n7445)
         );
  AOI21_X1 U9238 ( .B1(n7446), .B2(n10058), .A(n7445), .ZN(n7447) );
  OAI21_X1 U9239 ( .B1(n7470), .B2(n9803), .A(n7447), .ZN(P1_U3282) );
  INV_X1 U9240 ( .A(n7448), .ZN(n7450) );
  INV_X1 U9241 ( .A(n8217), .ZN(n8019) );
  OAI22_X1 U9242 ( .A1(n8019), .A2(n10370), .B1(n8209), .B2(n10373), .ZN(n7449) );
  OAI21_X1 U9243 ( .B1(n7450), .B2(n7449), .A(n4495), .ZN(n7453) );
  NAND2_X1 U9244 ( .A1(n7451), .A2(n8438), .ZN(n7452) );
  OAI211_X1 U9245 ( .C1(n4495), .C2(n7454), .A(n7453), .B(n7452), .ZN(P2_U3220) );
  INV_X1 U9246 ( .A(n7455), .ZN(n7456) );
  XNOR2_X1 U9247 ( .A(n7922), .B(n7856), .ZN(n7559) );
  NAND2_X1 U9248 ( .A1(n7460), .A2(n7559), .ZN(n7561) );
  OAI211_X1 U9249 ( .C1(n7460), .C2(n7559), .A(n7561), .B(n8242), .ZN(n7467)
         );
  INV_X1 U9250 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7461) );
  NOR2_X1 U9251 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7461), .ZN(n10248) );
  AOI21_X1 U9252 ( .B1(n8244), .B2(n8280), .A(n10248), .ZN(n7463) );
  NAND2_X1 U9253 ( .A1(n8257), .A2(n8278), .ZN(n7462) );
  OAI211_X1 U9254 ( .C1(n8210), .C2(n7464), .A(n7463), .B(n7462), .ZN(n7465)
         );
  AOI21_X1 U9255 ( .B1(n10428), .B2(n8237), .A(n7465), .ZN(n7466) );
  NAND2_X1 U9256 ( .A1(n7467), .A2(n7466), .ZN(P2_U3176) );
  OAI211_X1 U9257 ( .C1(n7470), .C2(n9815), .A(n7469), .B(n7468), .ZN(n7475)
         );
  OAI22_X1 U9258 ( .A1(n9875), .A2(n7645), .B1(n10192), .B2(n7072), .ZN(n7471)
         );
  AOI21_X1 U9259 ( .B1(n7475), .B2(n10192), .A(n7471), .ZN(n7472) );
  INV_X1 U9260 ( .A(n7472), .ZN(P1_U3533) );
  INV_X1 U9261 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7473) );
  OAI22_X1 U9262 ( .A1(n9929), .A2(n7645), .B1(n10175), .B2(n7473), .ZN(n7474)
         );
  AOI21_X1 U9263 ( .B1(n7475), .B2(n10175), .A(n7474), .ZN(n7476) );
  INV_X1 U9264 ( .A(n7476), .ZN(P1_U3486) );
  INV_X1 U9265 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7478) );
  MUX2_X1 U9266 ( .A(n7478), .B(P1_REG2_REG_14__SCAN_IN), .S(n7767), .Z(n7479)
         );
  AOI211_X1 U9267 ( .C1(n7480), .C2(n7479), .A(n7763), .B(n10018), .ZN(n7491)
         );
  INV_X1 U9268 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7483) );
  MUX2_X1 U9269 ( .A(n7483), .B(P1_REG1_REG_14__SCAN_IN), .S(n7767), .Z(n7484)
         );
  AOI211_X1 U9270 ( .C1(n7485), .C2(n7484), .A(n7766), .B(n9993), .ZN(n7490)
         );
  INV_X1 U9271 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7488) );
  NAND2_X1 U9272 ( .A1(n10025), .A2(n7767), .ZN(n7487) );
  NAND2_X1 U9273 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n7486) );
  OAI211_X1 U9274 ( .C1(n7488), .C2(n9601), .A(n7487), .B(n7486), .ZN(n7489)
         );
  OR3_X1 U9275 ( .A1(n7491), .A2(n7490), .A3(n7489), .ZN(P1_U3257) );
  INV_X1 U9276 ( .A(n7492), .ZN(n7494) );
  OAI222_X1 U9277 ( .A1(n8551), .A2(n9038), .B1(n8555), .B2(n7494), .C1(
        P2_U3151), .C2(n7493), .ZN(P2_U3273) );
  OAI222_X1 U9278 ( .A1(n7819), .A2(n9041), .B1(n4496), .B2(n7494), .C1(
        P1_U3086), .C2(n5455), .ZN(P1_U3333) );
  INV_X1 U9279 ( .A(n7497), .ZN(n9345) );
  XNOR2_X1 U9280 ( .A(n7495), .B(n9345), .ZN(n7580) );
  INV_X1 U9281 ( .A(n7580), .ZN(n7509) );
  NAND2_X1 U9282 ( .A1(n7496), .A2(n9254), .ZN(n7498) );
  XNOR2_X1 U9283 ( .A(n7498), .B(n7497), .ZN(n7499) );
  NAND2_X1 U9284 ( .A1(n7499), .A2(n10054), .ZN(n7502) );
  OR2_X1 U9285 ( .A1(n7708), .A2(n9195), .ZN(n7501) );
  NAND2_X1 U9286 ( .A1(n9508), .A2(n9197), .ZN(n7500) );
  AND2_X1 U9287 ( .A1(n7501), .A2(n7500), .ZN(n9958) );
  NAND2_X1 U9288 ( .A1(n7502), .A2(n9958), .ZN(n7578) );
  INV_X1 U9289 ( .A(n7589), .ZN(n7503) );
  NAND2_X1 U9290 ( .A1(n7579), .A2(n10066), .ZN(n7506) );
  AOI22_X1 U9291 ( .A1(n10043), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7504), .B2(
        n10042), .ZN(n7505) );
  OAI211_X1 U9292 ( .C1(n9964), .C2(n9800), .A(n7506), .B(n7505), .ZN(n7507)
         );
  AOI21_X1 U9293 ( .B1(n10058), .B2(n7578), .A(n7507), .ZN(n7508) );
  OAI21_X1 U9294 ( .B1(n9803), .B2(n7509), .A(n7508), .ZN(P1_U3281) );
  OR2_X1 U9295 ( .A1(n7516), .A2(n4503), .ZN(n7512) );
  NAND2_X1 U9296 ( .A1(n7510), .A2(n8733), .ZN(n7511) );
  NAND2_X1 U9297 ( .A1(n7512), .A2(n7511), .ZN(n7630) );
  INV_X1 U9298 ( .A(n7630), .ZN(n7628) );
  OAI22_X1 U9299 ( .A1(n7516), .A2(n8728), .B1(n5006), .B2(n8609), .ZN(n7518)
         );
  INV_X1 U9300 ( .A(n7631), .ZN(n7627) );
  XNOR2_X1 U9301 ( .A(n7637), .B(n7627), .ZN(n7519) );
  NAND2_X1 U9302 ( .A1(n7519), .A2(n7628), .ZN(n7595) );
  OAI21_X1 U9303 ( .B1(n7628), .B2(n7519), .A(n7595), .ZN(n7520) );
  NAND2_X1 U9304 ( .A1(n7520), .A2(n9966), .ZN(n7526) );
  OAI22_X1 U9305 ( .A1(n7522), .A2(n9214), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7521), .ZN(n7523) );
  AOI21_X1 U9306 ( .B1(n7524), .B2(n9211), .A(n7523), .ZN(n7525) );
  OAI211_X1 U9307 ( .C1(n5006), .C2(n9963), .A(n7526), .B(n7525), .ZN(P1_U3221) );
  INV_X1 U9308 ( .A(n7527), .ZN(n8040) );
  XOR2_X1 U9309 ( .A(n7528), .B(n8034), .Z(n7543) );
  XNOR2_X1 U9310 ( .A(n7529), .B(n4635), .ZN(n7531) );
  OAI22_X1 U9311 ( .A1(n8259), .A2(n8391), .B1(n8187), .B2(n8389), .ZN(n7530)
         );
  AOI21_X1 U9312 ( .B1(n7531), .B2(n8430), .A(n7530), .ZN(n7538) );
  MUX2_X1 U9313 ( .A(n7532), .B(n7538), .S(n10446), .Z(n7534) );
  NAND2_X1 U9314 ( .A1(n8250), .A2(n8473), .ZN(n7533) );
  OAI211_X1 U9315 ( .C1(n8493), .C2(n7543), .A(n7534), .B(n7533), .ZN(P2_U3474) );
  INV_X1 U9316 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n7535) );
  MUX2_X1 U9317 ( .A(n7535), .B(n7538), .S(n10430), .Z(n7537) );
  NAND2_X1 U9318 ( .A1(n8250), .A2(n8533), .ZN(n7536) );
  OAI211_X1 U9319 ( .C1(n7543), .C2(n8544), .A(n7537), .B(n7536), .ZN(P2_U3435) );
  MUX2_X1 U9320 ( .A(n7539), .B(n7538), .S(n4495), .Z(n7542) );
  INV_X1 U9321 ( .A(n7540), .ZN(n8263) );
  AOI22_X1 U9322 ( .A1(n8250), .A2(n8434), .B1(n8404), .B2(n8263), .ZN(n7541)
         );
  OAI211_X1 U9323 ( .C1(n7543), .C2(n8407), .A(n7542), .B(n7541), .ZN(P2_U3218) );
  XNOR2_X1 U9324 ( .A(n7544), .B(n8025), .ZN(n7557) );
  INV_X1 U9325 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7547) );
  XNOR2_X1 U9326 ( .A(n7545), .B(n8025), .ZN(n7546) );
  AOI222_X1 U9327 ( .A1(n8430), .A2(n7546), .B1(n8275), .B2(n6321), .C1(n8277), 
        .C2(n8427), .ZN(n7552) );
  MUX2_X1 U9328 ( .A(n7547), .B(n7552), .S(n10430), .Z(n7549) );
  NAND2_X1 U9329 ( .A1(n7751), .A2(n8533), .ZN(n7548) );
  OAI211_X1 U9330 ( .C1(n7557), .C2(n8544), .A(n7549), .B(n7548), .ZN(P2_U3432) );
  MUX2_X1 U9331 ( .A(n9120), .B(n7552), .S(n10446), .Z(n7551) );
  NAND2_X1 U9332 ( .A1(n7751), .A2(n8473), .ZN(n7550) );
  OAI211_X1 U9333 ( .C1(n7557), .C2(n8493), .A(n7551), .B(n7550), .ZN(P2_U3473) );
  INV_X1 U9334 ( .A(n7552), .ZN(n7554) );
  INV_X1 U9335 ( .A(n7751), .ZN(n7762) );
  OAI22_X1 U9336 ( .A1(n7762), .A2(n10370), .B1(n7755), .B2(n10373), .ZN(n7553) );
  OAI21_X1 U9337 ( .B1(n7554), .B2(n7553), .A(n4495), .ZN(n7556) );
  NAND2_X1 U9338 ( .A1(n10381), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7555) );
  OAI211_X1 U9339 ( .C1(n7557), .C2(n8407), .A(n7556), .B(n7555), .ZN(P2_U3219) );
  OR2_X1 U9340 ( .A1(n7559), .A2(n7558), .ZN(n7560) );
  NAND2_X1 U9341 ( .A1(n7561), .A2(n7560), .ZN(n7563) );
  XNOR2_X1 U9342 ( .A(n7568), .B(n7856), .ZN(n7748) );
  XOR2_X1 U9343 ( .A(n7749), .B(n7748), .Z(n7562) );
  NAND2_X1 U9344 ( .A1(n7563), .A2(n7562), .ZN(n7747) );
  OAI211_X1 U9345 ( .C1(n7563), .C2(n7562), .A(n7747), .B(n8242), .ZN(n7570)
         );
  INV_X1 U9346 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8914) );
  NOR2_X1 U9347 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8914), .ZN(n10266) );
  AOI21_X1 U9348 ( .B1(n8244), .B2(n8279), .A(n10266), .ZN(n7565) );
  NAND2_X1 U9349 ( .A1(n8257), .A2(n8277), .ZN(n7564) );
  OAI211_X1 U9350 ( .C1(n8210), .C2(n7566), .A(n7565), .B(n7564), .ZN(n7567)
         );
  AOI21_X1 U9351 ( .B1(n7568), .B2(n8237), .A(n7567), .ZN(n7569) );
  NAND2_X1 U9352 ( .A1(n7570), .A2(n7569), .ZN(P2_U3164) );
  NAND2_X1 U9353 ( .A1(n7575), .A2(n7571), .ZN(n7572) );
  OAI211_X1 U9354 ( .C1(n7573), .C2(n8551), .A(n7572), .B(n8130), .ZN(P2_U3272) );
  NAND2_X1 U9355 ( .A1(n7575), .A2(n7574), .ZN(n7577) );
  OR2_X1 U9356 ( .A1(n7576), .A2(P1_U3086), .ZN(n9470) );
  OAI211_X1 U9357 ( .C1(n8913), .C2(n7819), .A(n7577), .B(n9470), .ZN(P1_U3332) );
  AOI211_X1 U9358 ( .C1(n7580), .C2(n10172), .A(n7579), .B(n7578), .ZN(n7583)
         );
  MUX2_X1 U9359 ( .A(n7581), .B(n7583), .S(n10192), .Z(n7582) );
  OAI21_X1 U9360 ( .B1(n9964), .B2(n9875), .A(n7582), .ZN(P1_U3534) );
  INV_X1 U9361 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7584) );
  MUX2_X1 U9362 ( .A(n7584), .B(n7583), .S(n10175), .Z(n7585) );
  OAI21_X1 U9363 ( .B1(n9964), .B2(n9929), .A(n7585), .ZN(P1_U3489) );
  XOR2_X1 U9364 ( .A(n7586), .B(n9347), .Z(n7614) );
  INV_X1 U9365 ( .A(n7614), .ZN(n7594) );
  XNOR2_X1 U9366 ( .A(n7587), .B(n9347), .ZN(n7588) );
  AOI22_X1 U9367 ( .A1(n9507), .A2(n9197), .B1(n9184), .B2(n9505), .ZN(n7667)
         );
  OAI21_X1 U9368 ( .B1(n7588), .B2(n10036), .A(n7667), .ZN(n7612) );
  AOI211_X1 U9369 ( .C1(n7625), .C2(n7589), .A(n9794), .B(n7712), .ZN(n7613)
         );
  NAND2_X1 U9370 ( .A1(n7613), .A2(n10066), .ZN(n7591) );
  AOI22_X1 U9371 ( .A1(n10043), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7669), .B2(
        n10042), .ZN(n7590) );
  OAI211_X1 U9372 ( .C1(n5031), .C2(n9800), .A(n7591), .B(n7590), .ZN(n7592)
         );
  AOI21_X1 U9373 ( .B1(n10058), .B2(n7612), .A(n7592), .ZN(n7593) );
  OAI21_X1 U9374 ( .B1(n7594), .B2(n9803), .A(n7593), .ZN(P1_U3280) );
  OAI21_X1 U9375 ( .B1(n7631), .B2(n7637), .A(n7595), .ZN(n7599) );
  OAI22_X1 U9376 ( .A1(n7597), .A2(n8728), .B1(n10161), .B2(n8609), .ZN(n7596)
         );
  XNOR2_X1 U9377 ( .A(n7596), .B(n8731), .ZN(n7634) );
  OAI22_X1 U9378 ( .A1(n7597), .A2(n4503), .B1(n10161), .B2(n8728), .ZN(n7629)
         );
  XNOR2_X1 U9379 ( .A(n7634), .B(n7629), .ZN(n7598) );
  XNOR2_X1 U9380 ( .A(n7599), .B(n7598), .ZN(n7610) );
  INV_X1 U9381 ( .A(n7600), .ZN(n7608) );
  NAND2_X1 U9382 ( .A1(n7602), .A2(n7601), .ZN(n7604) );
  AOI21_X1 U9383 ( .B1(n7604), .B2(n9960), .A(n7603), .ZN(n7607) );
  NAND2_X1 U9384 ( .A1(n9217), .A2(n7605), .ZN(n7606) );
  OAI211_X1 U9385 ( .C1(n9970), .C2(n7608), .A(n7607), .B(n7606), .ZN(n7609)
         );
  AOI21_X1 U9386 ( .B1(n7610), .B2(n9966), .A(n7609), .ZN(n7611) );
  INV_X1 U9387 ( .A(n7611), .ZN(P1_U3231) );
  AOI211_X1 U9388 ( .C1(n7614), .C2(n10172), .A(n7613), .B(n7612), .ZN(n7616)
         );
  MUX2_X1 U9389 ( .A(n7375), .B(n7616), .S(n10192), .Z(n7615) );
  OAI21_X1 U9390 ( .B1(n5031), .B2(n9875), .A(n7615), .ZN(P1_U3535) );
  INV_X1 U9391 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7617) );
  MUX2_X1 U9392 ( .A(n7617), .B(n7616), .S(n10175), .Z(n7618) );
  OAI21_X1 U9393 ( .B1(n5031), .B2(n9929), .A(n7618), .ZN(P1_U3492) );
  INV_X1 U9394 ( .A(n7619), .ZN(n7672) );
  OAI222_X1 U9395 ( .A1(P1_U3086), .A2(n7621), .B1(n4496), .B2(n7672), .C1(
        n7620), .C2(n7819), .ZN(P1_U3331) );
  NAND2_X1 U9396 ( .A1(n7625), .A2(n8727), .ZN(n7623) );
  OR2_X1 U9397 ( .A1(n7708), .A2(n8728), .ZN(n7622) );
  NAND2_X1 U9398 ( .A1(n7623), .A2(n7622), .ZN(n7624) );
  XNOR2_X1 U9399 ( .A(n7624), .B(n7517), .ZN(n8567) );
  AOI22_X1 U9400 ( .A1(n7625), .A2(n8733), .B1(n8653), .B2(n9506), .ZN(n8565)
         );
  XNOR2_X1 U9401 ( .A(n8567), .B(n8565), .ZN(n7664) );
  INV_X1 U9402 ( .A(n7629), .ZN(n7626) );
  OAI22_X1 U9403 ( .A1(n7628), .A2(n7627), .B1(n7634), .B2(n7626), .ZN(n7636)
         );
  OAI21_X1 U9404 ( .B1(n7631), .B2(n7630), .A(n7629), .ZN(n7633) );
  NOR3_X1 U9405 ( .A1(n7631), .A2(n7630), .A3(n7629), .ZN(n7632) );
  OR2_X1 U9406 ( .A1(n7638), .A2(n4503), .ZN(n7640) );
  NAND2_X1 U9407 ( .A1(n8713), .A2(n8733), .ZN(n7639) );
  NOR2_X1 U9408 ( .A1(n7685), .A2(n7684), .ZN(n7647) );
  NAND2_X1 U9409 ( .A1(n7693), .A2(n8727), .ZN(n7642) );
  NAND2_X1 U9410 ( .A1(n9508), .A2(n8733), .ZN(n7641) );
  NAND2_X1 U9411 ( .A1(n7642), .A2(n7641), .ZN(n7643) );
  XNOR2_X1 U9412 ( .A(n7643), .B(n7517), .ZN(n7688) );
  OAI22_X1 U9413 ( .A1(n7645), .A2(n8728), .B1(n7644), .B2(n4503), .ZN(n7687)
         );
  NAND2_X1 U9414 ( .A1(n7688), .A2(n7687), .ZN(n7686) );
  INV_X1 U9415 ( .A(n7687), .ZN(n7648) );
  AOI21_X1 U9416 ( .B1(n7685), .B2(n7684), .A(n7648), .ZN(n7650) );
  NAND3_X1 U9417 ( .A1(n7685), .A2(n7684), .A3(n7648), .ZN(n7649) );
  OAI21_X1 U9418 ( .B1(n7650), .B2(n7688), .A(n7649), .ZN(n7651) );
  INV_X1 U9419 ( .A(n7651), .ZN(n7652) );
  AOI22_X1 U9420 ( .A1(n7653), .A2(n8727), .B1(n9507), .B2(n8733), .ZN(n7654)
         );
  XOR2_X1 U9421 ( .A(n7517), .B(n7654), .Z(n7657) );
  OAI22_X1 U9422 ( .A1(n9964), .A2(n8728), .B1(n7655), .B2(n4503), .ZN(n7656)
         );
  NOR2_X1 U9423 ( .A1(n7657), .A2(n7656), .ZN(n7658) );
  AOI21_X1 U9424 ( .B1(n7657), .B2(n7656), .A(n7658), .ZN(n9957) );
  NAND2_X1 U9425 ( .A1(n7662), .A2(n9957), .ZN(n9956) );
  INV_X1 U9426 ( .A(n7658), .ZN(n7659) );
  NAND2_X1 U9427 ( .A1(n9956), .A2(n7659), .ZN(n7663) );
  AND2_X1 U9428 ( .A1(n9957), .A2(n7664), .ZN(n7661) );
  INV_X1 U9429 ( .A(n7664), .ZN(n7660) );
  OAI21_X1 U9430 ( .B1(n7664), .B2(n7663), .A(n8569), .ZN(n7665) );
  NAND2_X1 U9431 ( .A1(n7665), .A2(n9966), .ZN(n7671) );
  OAI21_X1 U9432 ( .B1(n7667), .B2(n9214), .A(n7666), .ZN(n7668) );
  AOI21_X1 U9433 ( .B1(n7669), .B2(n9211), .A(n7668), .ZN(n7670) );
  OAI211_X1 U9434 ( .C1(n5031), .C2(n9963), .A(n7671), .B(n7670), .ZN(P1_U3234) );
  OAI222_X1 U9435 ( .A1(n8551), .A2(n7673), .B1(P2_U3151), .B2(n6331), .C1(
        n8562), .C2(n7672), .ZN(P2_U3271) );
  XNOR2_X1 U9436 ( .A(n7674), .B(n8037), .ZN(n7703) );
  XNOR2_X1 U9437 ( .A(n7675), .B(n8037), .ZN(n7676) );
  AOI222_X1 U9438 ( .A1(n8430), .A2(n7676), .B1(n8275), .B2(n8427), .C1(n8428), 
        .C2(n6321), .ZN(n7700) );
  MUX2_X1 U9439 ( .A(n7677), .B(n7700), .S(n10430), .Z(n7679) );
  NAND2_X1 U9440 ( .A1(n8181), .A2(n8533), .ZN(n7678) );
  OAI211_X1 U9441 ( .C1(n7703), .C2(n8544), .A(n7679), .B(n7678), .ZN(P2_U3438) );
  MUX2_X1 U9442 ( .A(n7680), .B(n7700), .S(n10446), .Z(n7682) );
  NAND2_X1 U9443 ( .A1(n8181), .A2(n8473), .ZN(n7681) );
  OAI211_X1 U9444 ( .C1(n7703), .C2(n8493), .A(n7682), .B(n7681), .ZN(P2_U3475) );
  XNOR2_X1 U9445 ( .A(n7683), .B(n7685), .ZN(n8709) );
  INV_X1 U9446 ( .A(n7684), .ZN(n8708) );
  NOR2_X1 U9447 ( .A1(n8709), .A2(n8708), .ZN(n8707) );
  AOI21_X1 U9448 ( .B1(n7685), .B2(n7683), .A(n8707), .ZN(n7690) );
  OAI21_X1 U9449 ( .B1(n7688), .B2(n7687), .A(n7686), .ZN(n7689) );
  XNOR2_X1 U9450 ( .A(n7690), .B(n7689), .ZN(n7698) );
  INV_X1 U9451 ( .A(n7691), .ZN(n7696) );
  AOI22_X1 U9452 ( .A1(n7692), .A2(n9960), .B1(P1_REG3_REG_11__SCAN_IN), .B2(
        P1_U3086), .ZN(n7695) );
  NAND2_X1 U9453 ( .A1(n9217), .A2(n7693), .ZN(n7694) );
  OAI211_X1 U9454 ( .C1(n9970), .C2(n7696), .A(n7695), .B(n7694), .ZN(n7697)
         );
  AOI21_X1 U9455 ( .B1(n7698), .B2(n9966), .A(n7697), .ZN(n7699) );
  INV_X1 U9456 ( .A(n7699), .ZN(P1_U3236) );
  MUX2_X1 U9457 ( .A(n5880), .B(n7700), .S(n4495), .Z(n7702) );
  AOI22_X1 U9458 ( .A1(n8181), .A2(n8434), .B1(n8404), .B2(n8175), .ZN(n7701)
         );
  OAI211_X1 U9459 ( .C1(n7703), .C2(n8407), .A(n7702), .B(n7701), .ZN(P2_U3217) );
  XNOR2_X1 U9460 ( .A(n7704), .B(n9349), .ZN(n9873) );
  INV_X1 U9461 ( .A(n9873), .ZN(n7717) );
  OAI21_X1 U9462 ( .B1(n7706), .B2(n9349), .A(n7705), .ZN(n7707) );
  NAND2_X1 U9463 ( .A1(n7707), .A2(n10054), .ZN(n7711) );
  OR2_X1 U9464 ( .A1(n7708), .A2(n9141), .ZN(n7710) );
  NAND2_X1 U9465 ( .A1(n9503), .A2(n9184), .ZN(n7709) );
  AND2_X1 U9466 ( .A1(n7710), .A2(n7709), .ZN(n8684) );
  NAND2_X1 U9467 ( .A1(n7711), .A2(n8684), .ZN(n9871) );
  AOI211_X1 U9468 ( .C1(n9263), .C2(n5033), .A(n9794), .B(n7726), .ZN(n9872)
         );
  NAND2_X1 U9469 ( .A1(n9872), .A2(n10066), .ZN(n7714) );
  AOI22_X1 U9470 ( .A1(n10043), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8687), .B2(
        n10042), .ZN(n7713) );
  OAI211_X1 U9471 ( .C1(n9930), .C2(n9800), .A(n7714), .B(n7713), .ZN(n7715)
         );
  AOI21_X1 U9472 ( .B1(n10058), .B2(n9871), .A(n7715), .ZN(n7716) );
  OAI21_X1 U9473 ( .B1(n7717), .B2(n9803), .A(n7716), .ZN(P1_U3279) );
  NAND2_X1 U9474 ( .A1(n7705), .A2(n7718), .ZN(n7720) );
  OR2_X1 U9475 ( .A1(n7719), .A2(n4579), .ZN(n9350) );
  XNOR2_X1 U9476 ( .A(n7720), .B(n9350), .ZN(n7724) );
  OR2_X1 U9477 ( .A1(n9142), .A2(n9195), .ZN(n7722) );
  NAND2_X1 U9478 ( .A1(n9505), .A2(n9197), .ZN(n7721) );
  AND2_X1 U9479 ( .A1(n7722), .A2(n7721), .ZN(n9215) );
  INV_X1 U9480 ( .A(n9215), .ZN(n7723) );
  AOI21_X1 U9481 ( .B1(n7724), .B2(n10054), .A(n7723), .ZN(n9977) );
  XOR2_X1 U9482 ( .A(n7725), .B(n9350), .Z(n9980) );
  NAND2_X1 U9483 ( .A1(n9980), .A2(n10067), .ZN(n7731) );
  OAI211_X1 U9484 ( .C1(n7726), .C2(n9978), .A(n10063), .B(n9795), .ZN(n9976)
         );
  INV_X1 U9485 ( .A(n9976), .ZN(n7729) );
  AOI22_X1 U9486 ( .A1(n10070), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9210), .B2(
        n10042), .ZN(n7727) );
  OAI21_X1 U9487 ( .B1(n9978), .B2(n9800), .A(n7727), .ZN(n7728) );
  AOI21_X1 U9488 ( .B1(n7729), .B2(n10066), .A(n7728), .ZN(n7730) );
  OAI211_X1 U9489 ( .C1(n10043), .C2(n9977), .A(n7731), .B(n7730), .ZN(
        P1_U3278) );
  INV_X1 U9490 ( .A(n7733), .ZN(n7734) );
  AOI21_X1 U9491 ( .B1(n8043), .B2(n7732), .A(n7734), .ZN(n8545) );
  XNOR2_X1 U9492 ( .A(n7735), .B(n8043), .ZN(n7736) );
  OAI222_X1 U9493 ( .A1(n8391), .A2(n8187), .B1(n8389), .B2(n8154), .C1(n7736), 
        .C2(n8387), .ZN(n8490) );
  NAND2_X1 U9494 ( .A1(n8490), .A2(n4495), .ZN(n7741) );
  INV_X1 U9495 ( .A(n8184), .ZN(n7737) );
  OAI22_X1 U9496 ( .A1(n4495), .A2(n7738), .B1(n7737), .B2(n10373), .ZN(n7739)
         );
  AOI21_X1 U9497 ( .B1(n8491), .B2(n8434), .A(n7739), .ZN(n7740) );
  OAI211_X1 U9498 ( .C1(n8545), .C2(n8407), .A(n7741), .B(n7740), .ZN(P2_U3216) );
  INV_X1 U9499 ( .A(n7742), .ZN(n7745) );
  OAI222_X1 U9500 ( .A1(P1_U3086), .A2(n7744), .B1(n4496), .B2(n7745), .C1(
        n7743), .C2(n7819), .ZN(P1_U3330) );
  OAI222_X1 U9501 ( .A1(n8551), .A2(n7746), .B1(P2_U3151), .B2(n6332), .C1(
        n8562), .C2(n7745), .ZN(P2_U3270) );
  XNOR2_X1 U9502 ( .A(n8217), .B(n7856), .ZN(n8211) );
  INV_X1 U9503 ( .A(n8211), .ZN(n7750) );
  XNOR2_X1 U9504 ( .A(n7751), .B(n7856), .ZN(n7820) );
  XOR2_X1 U9505 ( .A(n8259), .B(n7820), .Z(n7752) );
  OAI21_X1 U9506 ( .B1(n7753), .B2(n7752), .A(n7822), .ZN(n7754) );
  NAND2_X1 U9507 ( .A1(n7754), .A2(n8242), .ZN(n7761) );
  INV_X1 U9508 ( .A(n7755), .ZN(n7759) );
  NAND2_X1 U9509 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n10304) );
  INV_X1 U9510 ( .A(n10304), .ZN(n7756) );
  AOI21_X1 U9511 ( .B1(n8257), .B2(n8275), .A(n7756), .ZN(n7757) );
  OAI21_X1 U9512 ( .B1(n8260), .B2(n8020), .A(n7757), .ZN(n7758) );
  AOI21_X1 U9513 ( .B1(n7759), .B2(n8262), .A(n7758), .ZN(n7760) );
  OAI211_X1 U9514 ( .C1(n7762), .C2(n8266), .A(n7761), .B(n7760), .ZN(P2_U3155) );
  INV_X1 U9515 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7764) );
  NOR2_X1 U9516 ( .A1(n7764), .A2(n7765), .ZN(n9544) );
  AOI211_X1 U9517 ( .C1(n7765), .C2(n7764), .A(n9544), .B(n10018), .ZN(n7774)
         );
  INV_X1 U9518 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9981) );
  NOR2_X1 U9519 ( .A1(n9981), .A2(n7768), .ZN(n9533) );
  AOI211_X1 U9520 ( .C1(n7768), .C2(n9981), .A(n9533), .B(n9993), .ZN(n7773)
         );
  INV_X1 U9521 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7771) );
  NAND2_X1 U9522 ( .A1(n10025), .A2(n7769), .ZN(n7770) );
  NAND2_X1 U9523 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9212) );
  OAI211_X1 U9524 ( .C1(n7771), .C2(n9601), .A(n7770), .B(n9212), .ZN(n7772)
         );
  OR3_X1 U9525 ( .A1(n7774), .A2(n7773), .A3(n7772), .ZN(P1_U3258) );
  INV_X1 U9526 ( .A(n7775), .ZN(n7805) );
  OAI222_X1 U9527 ( .A1(n8551), .A2(n7777), .B1(P2_U3151), .B2(n7776), .C1(
        n8555), .C2(n7805), .ZN(P2_U3269) );
  NAND2_X1 U9528 ( .A1(n7778), .A2(n5083), .ZN(n7780) );
  INV_X1 U9529 ( .A(n9490), .ZN(n7779) );
  OR2_X1 U9530 ( .A1(n9810), .A2(n7779), .ZN(n9369) );
  NAND2_X1 U9531 ( .A1(n9810), .A2(n7779), .ZN(n9367) );
  NAND2_X1 U9532 ( .A1(n9369), .A2(n9367), .ZN(n9359) );
  XNOR2_X1 U9533 ( .A(n7780), .B(n9359), .ZN(n9816) );
  INV_X1 U9534 ( .A(n9318), .ZN(n7781) );
  AOI21_X1 U9535 ( .B1(n7782), .B2(n5722), .A(n7781), .ZN(n7783) );
  XNOR2_X1 U9536 ( .A(n7783), .B(n9359), .ZN(n7784) );
  NAND2_X1 U9537 ( .A1(n4494), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n7788) );
  NAND2_X1 U9538 ( .A1(n5079), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7787) );
  NAND2_X1 U9539 ( .A1(n7785), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7786) );
  AND3_X1 U9540 ( .A1(n7788), .A2(n7787), .A3(n7786), .ZN(n9371) );
  AOI211_X1 U9541 ( .C1(n9810), .C2(n7793), .A(n9794), .B(n9607), .ZN(n9809)
         );
  NAND2_X1 U9542 ( .A1(n9809), .A2(n10066), .ZN(n7796) );
  AOI22_X1 U9543 ( .A1(n10070), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n7794), .B2(
        n10042), .ZN(n7795) );
  OAI211_X1 U9544 ( .C1(n5012), .C2(n9800), .A(n7796), .B(n7795), .ZN(n7797)
         );
  AOI21_X1 U9545 ( .B1(n9813), .B2(n10058), .A(n7797), .ZN(n7798) );
  OAI21_X1 U9546 ( .B1(n9816), .B2(n9803), .A(n7798), .ZN(P1_U3356) );
  INV_X1 U9547 ( .A(n7799), .ZN(n8554) );
  OAI222_X1 U9548 ( .A1(n7819), .A2(n7801), .B1(n4496), .B2(n8554), .C1(n7800), 
        .C2(P1_U3086), .ZN(P1_U3326) );
  INV_X1 U9549 ( .A(n7802), .ZN(n8563) );
  OAI222_X1 U9550 ( .A1(n7819), .A2(n7803), .B1(n4496), .B2(n8563), .C1(n5456), 
        .C2(P1_U3086), .ZN(P1_U3328) );
  OAI222_X1 U9551 ( .A1(P1_U3086), .A2(n7806), .B1(n4496), .B2(n7805), .C1(
        n7804), .C2(n7819), .ZN(P1_U3329) );
  INV_X1 U9552 ( .A(n7808), .ZN(n7809) );
  NAND2_X1 U9553 ( .A1(n8404), .A2(n7809), .ZN(n8294) );
  OAI21_X1 U9554 ( .B1(n4495), .B2(n7810), .A(n8294), .ZN(n7814) );
  NOR2_X1 U9555 ( .A1(n7812), .A2(n7811), .ZN(n7813) );
  AOI211_X1 U9556 ( .C1(n8419), .C2(n7815), .A(n7814), .B(n7813), .ZN(n7816)
         );
  OAI21_X1 U9557 ( .B1(n7807), .B2(n10381), .A(n7816), .ZN(P2_U3204) );
  INV_X1 U9558 ( .A(n7817), .ZN(n8558) );
  OAI222_X1 U9559 ( .A1(n7819), .A2(n7818), .B1(n4496), .B2(n8558), .C1(n5454), 
        .C2(P1_U3086), .ZN(P1_U3327) );
  INV_X1 U9560 ( .A(n7885), .ZN(n7883) );
  OAI222_X1 U9561 ( .A1(n8551), .A2(n7886), .B1(n8562), .B2(n7883), .C1(n5973), 
        .C2(P2_U3151), .ZN(P2_U3265) );
  NAND2_X1 U9562 ( .A1(n7820), .A2(n8259), .ZN(n7821) );
  XNOR2_X1 U9563 ( .A(n8250), .B(n7856), .ZN(n7823) );
  XNOR2_X1 U9564 ( .A(n7823), .B(n8179), .ZN(n8252) );
  INV_X1 U9565 ( .A(n7823), .ZN(n7824) );
  NAND2_X1 U9566 ( .A1(n7824), .A2(n8275), .ZN(n7825) );
  NAND2_X1 U9567 ( .A1(n8254), .A2(n7825), .ZN(n8174) );
  XNOR2_X1 U9568 ( .A(n8181), .B(n7856), .ZN(n8172) );
  NAND2_X1 U9569 ( .A1(n8172), .A2(n8187), .ZN(n7826) );
  XNOR2_X1 U9570 ( .A(n8491), .B(n7856), .ZN(n7831) );
  XOR2_X1 U9571 ( .A(n8235), .B(n7831), .Z(n8228) );
  XNOR2_X1 U9572 ( .A(n8435), .B(n7856), .ZN(n7827) );
  NAND2_X1 U9573 ( .A1(n7827), .A2(n8154), .ZN(n7832) );
  INV_X1 U9574 ( .A(n7832), .ZN(n7828) );
  XNOR2_X1 U9575 ( .A(n7827), .B(n8412), .ZN(n8232) );
  OR2_X1 U9576 ( .A1(n7828), .A2(n8232), .ZN(n7830) );
  AND2_X1 U9577 ( .A1(n8228), .A2(n7830), .ZN(n8147) );
  XNOR2_X1 U9578 ( .A(n8476), .B(n7856), .ZN(n7836) );
  XOR2_X1 U9579 ( .A(n8202), .B(n7836), .Z(n8151) );
  AND2_X1 U9580 ( .A1(n8147), .A2(n8151), .ZN(n7829) );
  INV_X1 U9581 ( .A(n8151), .ZN(n7835) );
  INV_X1 U9582 ( .A(n7830), .ZN(n7834) );
  NAND2_X1 U9583 ( .A1(n7831), .A2(n8235), .ZN(n8229) );
  AND2_X1 U9584 ( .A1(n8229), .A2(n7832), .ZN(n7833) );
  OR2_X1 U9585 ( .A1(n7834), .A2(n7833), .ZN(n8148) );
  XNOR2_X1 U9586 ( .A(n7837), .B(n7856), .ZN(n7838) );
  XNOR2_X1 U9587 ( .A(n7838), .B(n8390), .ZN(n8199) );
  INV_X1 U9588 ( .A(n7838), .ZN(n7839) );
  NAND2_X1 U9589 ( .A1(n7839), .A2(n8390), .ZN(n7840) );
  XNOR2_X1 U9590 ( .A(n8469), .B(n7856), .ZN(n7841) );
  XOR2_X1 U9591 ( .A(n8222), .B(n7841), .Z(n8159) );
  XOR2_X1 U9592 ( .A(n7856), .B(n8463), .Z(n7843) );
  INV_X1 U9593 ( .A(n7843), .ZN(n7842) );
  XNOR2_X1 U9594 ( .A(n7842), .B(n8273), .ZN(n8220) );
  NOR2_X1 U9595 ( .A1(n7843), .A2(n8273), .ZN(n7844) );
  AOI21_X1 U9596 ( .B1(n8219), .B2(n8220), .A(n7844), .ZN(n7848) );
  XNOR2_X1 U9597 ( .A(n7845), .B(n6681), .ZN(n7846) );
  XNOR2_X1 U9598 ( .A(n7848), .B(n7846), .ZN(n8140) );
  INV_X1 U9599 ( .A(n7846), .ZN(n7847) );
  OR2_X1 U9600 ( .A1(n7848), .A2(n7847), .ZN(n7849) );
  XNOR2_X1 U9601 ( .A(n8518), .B(n7856), .ZN(n7850) );
  XOR2_X1 U9602 ( .A(n8361), .B(n7850), .Z(n8192) );
  NAND2_X1 U9603 ( .A1(n7850), .A2(n8361), .ZN(n7851) );
  XNOR2_X1 U9604 ( .A(n8513), .B(n7856), .ZN(n7852) );
  XOR2_X1 U9605 ( .A(n8326), .B(n7852), .Z(n8166) );
  XNOR2_X1 U9606 ( .A(n8331), .B(n7856), .ZN(n7853) );
  XOR2_X1 U9607 ( .A(n8316), .B(n7853), .Z(n8241) );
  NAND2_X1 U9608 ( .A1(n8240), .A2(n8241), .ZN(n7855) );
  NAND2_X1 U9609 ( .A1(n7853), .A2(n8316), .ZN(n7854) );
  NAND2_X1 U9610 ( .A1(n7855), .A2(n7854), .ZN(n8132) );
  XNOR2_X1 U9611 ( .A(n8448), .B(n6681), .ZN(n7865) );
  NAND2_X1 U9612 ( .A1(n7865), .A2(n8272), .ZN(n7858) );
  OAI21_X1 U9613 ( .B1(n7865), .B2(n8272), .A(n7858), .ZN(n8131) );
  XNOR2_X1 U9614 ( .A(n7856), .B(n8315), .ZN(n7857) );
  XNOR2_X1 U9615 ( .A(n8303), .B(n7857), .ZN(n7864) );
  NAND2_X1 U9616 ( .A1(n7864), .A2(n8242), .ZN(n7872) );
  INV_X1 U9617 ( .A(n7858), .ZN(n7859) );
  NOR3_X1 U9618 ( .A1(n7859), .A2(n7864), .A3(n8251), .ZN(n7860) );
  NAND2_X1 U9619 ( .A1(n8133), .A2(n7860), .ZN(n7871) );
  AOI22_X1 U9620 ( .A1(n8272), .A2(n8244), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n7863) );
  INV_X1 U9621 ( .A(n7861), .ZN(n8270) );
  NAND2_X1 U9622 ( .A1(n8257), .A2(n8270), .ZN(n7862) );
  OAI211_X1 U9623 ( .C1(n8300), .C2(n8210), .A(n7863), .B(n7862), .ZN(n7869)
         );
  INV_X1 U9624 ( .A(n7864), .ZN(n7867) );
  INV_X1 U9625 ( .A(n7865), .ZN(n7866) );
  NOR4_X1 U9626 ( .A1(n7867), .A2(n7866), .A3(n8327), .A4(n8251), .ZN(n7868)
         );
  AOI211_X1 U9627 ( .C1(n8303), .C2(n8237), .A(n7869), .B(n7868), .ZN(n7870)
         );
  OAI211_X1 U9628 ( .C1(n8133), .C2(n7872), .A(n7871), .B(n7870), .ZN(P2_U3160) );
  INV_X1 U9629 ( .A(n7873), .ZN(n7879) );
  NOR2_X1 U9630 ( .A1(n7874), .A2(n9611), .ZN(n7878) );
  AOI22_X1 U9631 ( .A1(n10070), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n8740), .B2(
        n10042), .ZN(n7875) );
  OAI21_X1 U9632 ( .B1(n7876), .B2(n9800), .A(n7875), .ZN(n7877) );
  AOI211_X1 U9633 ( .C1(n7879), .C2(n10058), .A(n7878), .B(n7877), .ZN(n7880)
         );
  OAI21_X1 U9634 ( .B1(n7881), .B2(n9803), .A(n7880), .ZN(P1_U3265) );
  OAI222_X1 U9635 ( .A1(P1_U3086), .A2(n7884), .B1(n4496), .B2(n7883), .C1(
        n7882), .C2(n7819), .ZN(P1_U3325) );
  NAND2_X1 U9636 ( .A1(n7885), .A2(n7891), .ZN(n7888) );
  OR2_X1 U9637 ( .A1(n7893), .A2(n7886), .ZN(n7887) );
  NAND2_X1 U9638 ( .A1(n7888), .A2(n7887), .ZN(n8498) );
  NAND2_X1 U9639 ( .A1(n8498), .A2(n7889), .ZN(n8107) );
  NAND2_X1 U9640 ( .A1(n8546), .A2(n7891), .ZN(n7895) );
  OR2_X1 U9641 ( .A1(n7893), .A2(n7892), .ZN(n7894) );
  INV_X1 U9642 ( .A(n8443), .ZN(n8495) );
  INV_X1 U9643 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n7899) );
  OR2_X1 U9644 ( .A1(n6050), .A2(n7899), .ZN(n7905) );
  INV_X1 U9645 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9040) );
  OR2_X1 U9646 ( .A1(n7900), .A2(n9040), .ZN(n7904) );
  INV_X1 U9647 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n7901) );
  OR2_X1 U9648 ( .A1(n7902), .A2(n7901), .ZN(n7903) );
  INV_X1 U9649 ( .A(n8498), .ZN(n8298) );
  AND2_X1 U9650 ( .A1(n8298), .A2(n8269), .ZN(n8105) );
  INV_X1 U9651 ( .A(n7907), .ZN(n8092) );
  NAND2_X1 U9652 ( .A1(n8092), .A2(n8307), .ZN(n8089) );
  NAND2_X1 U9653 ( .A1(n8083), .A2(n4759), .ZN(n8349) );
  INV_X1 U9654 ( .A(n7909), .ZN(n8084) );
  NAND4_X1 U9655 ( .A1(n7911), .A2(n7910), .A3(n6297), .A4(n7971), .ZN(n7914)
         );
  INV_X1 U9656 ( .A(n7981), .ZN(n7913) );
  NOR3_X1 U9657 ( .A1(n7914), .A2(n7913), .A3(n7912), .ZN(n7917) );
  NAND4_X1 U9658 ( .A1(n7917), .A2(n7916), .A3(n8001), .A4(n7915), .ZN(n7919)
         );
  NOR2_X1 U9659 ( .A1(n7919), .A2(n7918), .ZN(n7920) );
  NAND4_X1 U9660 ( .A1(n7923), .A2(n7922), .A3(n7921), .A4(n7920), .ZN(n7924)
         );
  NOR2_X1 U9661 ( .A1(n7925), .A2(n7924), .ZN(n7926) );
  NAND4_X1 U9662 ( .A1(n8037), .A2(n8025), .A3(n8034), .A4(n7926), .ZN(n7927)
         );
  NOR2_X1 U9663 ( .A1(n8043), .A2(n7927), .ZN(n7930) );
  NAND4_X1 U9664 ( .A1(n8420), .A2(n7930), .A3(n7929), .A4(n7928), .ZN(n7931)
         );
  NOR2_X1 U9665 ( .A1(n8400), .A2(n7931), .ZN(n7932) );
  NAND4_X1 U9666 ( .A1(n8358), .A2(n8384), .A3(n7932), .A4(n8375), .ZN(n7933)
         );
  NOR2_X1 U9667 ( .A1(n8349), .A2(n7933), .ZN(n7934) );
  NAND2_X1 U9668 ( .A1(n8335), .A2(n7934), .ZN(n7935) );
  NOR2_X1 U9669 ( .A1(n8089), .A2(n7935), .ZN(n7937) );
  NAND4_X1 U9670 ( .A1(n8107), .A2(n6309), .A3(n7937), .A4(n7936), .ZN(n7938)
         );
  INV_X1 U9671 ( .A(n8293), .ZN(n8268) );
  NAND2_X1 U9672 ( .A1(n8495), .A2(n8293), .ZN(n8122) );
  INV_X1 U9673 ( .A(n7939), .ZN(n7940) );
  NAND2_X1 U9674 ( .A1(n7940), .A2(n8106), .ZN(n8062) );
  INV_X1 U9675 ( .A(n7941), .ZN(n7942) );
  OAI21_X1 U9676 ( .B1(n8400), .B2(n7942), .A(n8106), .ZN(n8060) );
  NAND2_X1 U9677 ( .A1(n7951), .A2(n7949), .ZN(n7943) );
  MUX2_X1 U9678 ( .A(n7953), .B(n7943), .S(n8106), .Z(n8000) );
  AND2_X1 U9679 ( .A1(n7945), .A2(n7944), .ZN(n7947) );
  OAI211_X1 U9680 ( .C1(n8000), .C2(n7947), .A(n7946), .B(n8004), .ZN(n7955)
         );
  AND2_X1 U9681 ( .A1(n7949), .A2(n7948), .ZN(n7952) );
  OAI211_X1 U9682 ( .C1(n7953), .C2(n7952), .A(n7951), .B(n7950), .ZN(n7954)
         );
  MUX2_X1 U9683 ( .A(n7955), .B(n7954), .S(n8112), .Z(n7956) );
  INV_X1 U9684 ( .A(n7956), .ZN(n8003) );
  NAND2_X1 U9685 ( .A1(n7960), .A2(n7957), .ZN(n7958) );
  NAND2_X1 U9686 ( .A1(n7958), .A2(n8106), .ZN(n7962) );
  NAND3_X1 U9687 ( .A1(n7960), .A2(n7959), .A3(n8128), .ZN(n7961) );
  NAND2_X1 U9688 ( .A1(n7962), .A2(n7961), .ZN(n7965) );
  NAND2_X1 U9689 ( .A1(n6296), .A2(n7963), .ZN(n7964) );
  NAND2_X1 U9690 ( .A1(n7965), .A2(n7964), .ZN(n7968) );
  INV_X1 U9691 ( .A(n7966), .ZN(n7967) );
  MUX2_X1 U9692 ( .A(n7968), .B(n8106), .S(n7967), .Z(n7973) );
  INV_X1 U9693 ( .A(n7959), .ZN(n7969) );
  NAND2_X1 U9694 ( .A1(n7969), .A2(n8106), .ZN(n7970) );
  AND2_X1 U9695 ( .A1(n7971), .A2(n7970), .ZN(n7972) );
  NAND2_X1 U9696 ( .A1(n7973), .A2(n7972), .ZN(n7980) );
  NAND2_X1 U9697 ( .A1(n8289), .A2(n10371), .ZN(n7974) );
  NAND2_X1 U9698 ( .A1(n7992), .A2(n7974), .ZN(n7977) );
  NAND2_X1 U9699 ( .A1(n7983), .A2(n7975), .ZN(n7976) );
  MUX2_X1 U9700 ( .A(n7977), .B(n7976), .S(n8106), .Z(n7978) );
  INV_X1 U9701 ( .A(n7978), .ZN(n7979) );
  NAND2_X1 U9702 ( .A1(n7980), .A2(n7979), .ZN(n7982) );
  INV_X1 U9703 ( .A(n7983), .ZN(n7986) );
  AND2_X1 U9704 ( .A1(n7988), .A2(n7984), .ZN(n7998) );
  NAND2_X1 U9705 ( .A1(n8287), .A2(n10364), .ZN(n7985) );
  OAI211_X1 U9706 ( .C1(n7996), .C2(n7986), .A(n7998), .B(n7985), .ZN(n7991)
         );
  INV_X1 U9707 ( .A(n7987), .ZN(n7989) );
  NAND2_X1 U9708 ( .A1(n7989), .A2(n7988), .ZN(n7990) );
  INV_X1 U9709 ( .A(n7992), .ZN(n7995) );
  OAI211_X1 U9710 ( .C1(n7996), .C2(n7995), .A(n7994), .B(n7993), .ZN(n7999)
         );
  INV_X1 U9711 ( .A(n8000), .ZN(n8002) );
  NAND2_X1 U9712 ( .A1(n8009), .A2(n8004), .ZN(n8007) );
  NAND2_X1 U9713 ( .A1(n8009), .A2(n8008), .ZN(n8011) );
  INV_X1 U9714 ( .A(n8012), .ZN(n8015) );
  INV_X1 U9715 ( .A(n8013), .ZN(n8014) );
  MUX2_X1 U9716 ( .A(n8015), .B(n8014), .S(n8112), .Z(n8016) );
  INV_X1 U9717 ( .A(n8016), .ZN(n8017) );
  MUX2_X1 U9718 ( .A(n8020), .B(n8019), .S(n8112), .Z(n8021) );
  OAI21_X1 U9719 ( .B1(n8024), .B2(n8022), .A(n8021), .ZN(n8028) );
  INV_X1 U9720 ( .A(n8025), .ZN(n8026) );
  AOI21_X1 U9721 ( .B1(n8028), .B2(n8027), .A(n8026), .ZN(n8033) );
  INV_X1 U9722 ( .A(n8029), .ZN(n8031) );
  MUX2_X1 U9723 ( .A(n8031), .B(n8030), .S(n8112), .Z(n8032) );
  OR2_X1 U9724 ( .A1(n8033), .A2(n8032), .ZN(n8035) );
  XNOR2_X1 U9725 ( .A(n8038), .B(n8112), .ZN(n8039) );
  AND2_X1 U9726 ( .A1(n8412), .A2(n8112), .ZN(n8048) );
  NAND2_X1 U9727 ( .A1(n8154), .A2(n8106), .ZN(n8047) );
  NAND2_X1 U9728 ( .A1(n8435), .A2(n8047), .ZN(n8042) );
  OAI21_X1 U9729 ( .B1(n8435), .B2(n8048), .A(n8042), .ZN(n8045) );
  INV_X1 U9730 ( .A(n8043), .ZN(n8044) );
  AND2_X1 U9731 ( .A1(n8045), .A2(n8044), .ZN(n8046) );
  INV_X1 U9732 ( .A(n8047), .ZN(n8049) );
  AOI22_X1 U9733 ( .A1(n8049), .A2(n8050), .B1(n8051), .B2(n8048), .ZN(n8054)
         );
  OAI211_X1 U9734 ( .C1(n8050), .C2(n8154), .A(n8106), .B(n8435), .ZN(n8053)
         );
  INV_X1 U9735 ( .A(n8435), .ZN(n8489) );
  OAI211_X1 U9736 ( .C1(n8412), .C2(n8051), .A(n8489), .B(n8112), .ZN(n8052)
         );
  NAND4_X1 U9737 ( .A1(n8420), .A2(n8054), .A3(n8053), .A4(n8052), .ZN(n8058)
         );
  NAND2_X1 U9738 ( .A1(n8380), .A2(n8055), .ZN(n8056) );
  NAND2_X1 U9739 ( .A1(n8056), .A2(n8112), .ZN(n8057) );
  NAND4_X1 U9740 ( .A1(n8060), .A2(n8059), .A3(n8058), .A4(n8057), .ZN(n8061)
         );
  NAND2_X1 U9741 ( .A1(n8062), .A2(n8061), .ZN(n8070) );
  NAND3_X1 U9742 ( .A1(n8375), .A2(n8070), .A3(n8067), .ZN(n8064) );
  NAND2_X1 U9743 ( .A1(n8463), .A2(n8388), .ZN(n8063) );
  NAND3_X1 U9744 ( .A1(n8064), .A2(n8063), .A3(n8078), .ZN(n8065) );
  NAND2_X1 U9745 ( .A1(n8065), .A2(n8106), .ZN(n8077) );
  AND2_X1 U9746 ( .A1(n8066), .A2(n8112), .ZN(n8069) );
  NAND2_X1 U9747 ( .A1(n8067), .A2(n4567), .ZN(n8068) );
  AOI22_X1 U9748 ( .A1(n8070), .A2(n8384), .B1(n8069), .B2(n8068), .ZN(n8074)
         );
  OAI21_X1 U9749 ( .B1(n8074), .B2(n4762), .A(n8073), .ZN(n8075) );
  NAND3_X1 U9750 ( .A1(n8085), .A2(n8078), .A3(n4759), .ZN(n8079) );
  NAND3_X1 U9751 ( .A1(n8079), .A2(n8112), .A3(n8083), .ZN(n8080) );
  NAND2_X1 U9752 ( .A1(n8080), .A2(n8335), .ZN(n8081) );
  OAI21_X1 U9753 ( .B1(n8082), .B2(n8106), .A(n8081), .ZN(n8088) );
  NAND3_X1 U9754 ( .A1(n8085), .A2(n8084), .A3(n8083), .ZN(n8086) );
  NAND3_X1 U9755 ( .A1(n8086), .A2(n8106), .A3(n4759), .ZN(n8087) );
  NAND2_X1 U9756 ( .A1(n8088), .A2(n8087), .ZN(n8090) );
  OAI211_X1 U9757 ( .C1(n8112), .C2(n8091), .A(n8090), .B(n8323), .ZN(n8098)
         );
  MUX2_X1 U9758 ( .A(n8307), .B(n8092), .S(n8106), .Z(n8093) );
  MUX2_X1 U9759 ( .A(n8095), .B(n8094), .S(n8112), .Z(n8096) );
  MUX2_X1 U9760 ( .A(n8315), .B(n8114), .S(n8106), .Z(n8102) );
  OR2_X1 U9761 ( .A1(n8100), .A2(n8102), .ZN(n8101) );
  NAND2_X1 U9762 ( .A1(n8103), .A2(n8101), .ZN(n8115) );
  NAND2_X1 U9763 ( .A1(n8115), .A2(n8315), .ZN(n8104) );
  NAND3_X1 U9764 ( .A1(n8104), .A2(n5092), .A3(n8113), .ZN(n8110) );
  NAND2_X1 U9765 ( .A1(n4982), .A2(n8106), .ZN(n8108) );
  NAND2_X1 U9766 ( .A1(n8108), .A2(n8107), .ZN(n8109) );
  NAND2_X1 U9767 ( .A1(n8110), .A2(n8109), .ZN(n8121) );
  NAND4_X1 U9768 ( .A1(n8113), .A2(n8112), .A3(n8111), .A4(n4982), .ZN(n8117)
         );
  AND2_X1 U9769 ( .A1(n8115), .A2(n8114), .ZN(n8116) );
  INV_X1 U9770 ( .A(n5886), .ZN(n8125) );
  NAND3_X1 U9771 ( .A1(n8126), .A2(n8125), .A3(n5948), .ZN(n8127) );
  OAI211_X1 U9772 ( .C1(n8128), .C2(n8130), .A(n8127), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8129) );
  AOI21_X1 U9773 ( .B1(n8132), .B2(n8131), .A(n8251), .ZN(n8134) );
  NAND2_X1 U9774 ( .A1(n8134), .A2(n8133), .ZN(n8139) );
  AOI22_X1 U9775 ( .A1(n8257), .A2(n8271), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8136) );
  NAND2_X1 U9776 ( .A1(n8262), .A2(n8317), .ZN(n8135) );
  OAI211_X1 U9777 ( .C1(n8316), .C2(n8260), .A(n8136), .B(n8135), .ZN(n8137)
         );
  AOI21_X1 U9778 ( .B1(n8448), .B2(n8237), .A(n8137), .ZN(n8138) );
  NAND2_X1 U9779 ( .A1(n8139), .A2(n8138), .ZN(P2_U3154) );
  XNOR2_X1 U9780 ( .A(n8140), .B(n8369), .ZN(n8145) );
  NAND2_X1 U9781 ( .A1(n8262), .A2(n8362), .ZN(n8142) );
  AOI22_X1 U9782 ( .A1(n8244), .A2(n8273), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8141) );
  OAI211_X1 U9783 ( .C1(n8361), .C2(n8246), .A(n8142), .B(n8141), .ZN(n8143)
         );
  AOI21_X1 U9784 ( .B1(n8460), .B2(n8237), .A(n8143), .ZN(n8144) );
  OAI21_X1 U9785 ( .B1(n8145), .B2(n8251), .A(n8144), .ZN(P2_U3156) );
  NAND2_X1 U9786 ( .A1(n8146), .A2(n8147), .ZN(n8149) );
  NAND2_X1 U9787 ( .A1(n8149), .A2(n8148), .ZN(n8150) );
  XOR2_X1 U9788 ( .A(n8151), .B(n8150), .Z(n8157) );
  NAND2_X1 U9789 ( .A1(n8262), .A2(n8416), .ZN(n8153) );
  AOI22_X1 U9790 ( .A1(n8257), .A2(n8413), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3151), .ZN(n8152) );
  OAI211_X1 U9791 ( .C1(n8154), .C2(n8260), .A(n8153), .B(n8152), .ZN(n8155)
         );
  AOI21_X1 U9792 ( .B1(n8476), .B2(n8237), .A(n8155), .ZN(n8156) );
  OAI21_X1 U9793 ( .B1(n8157), .B2(n8251), .A(n8156), .ZN(P2_U3159) );
  XOR2_X1 U9794 ( .A(n8158), .B(n8159), .Z(n8164) );
  NAND2_X1 U9795 ( .A1(n8262), .A2(n8392), .ZN(n8161) );
  AOI22_X1 U9796 ( .A1(n8257), .A2(n8273), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8160) );
  OAI211_X1 U9797 ( .C1(n8390), .C2(n8260), .A(n8161), .B(n8160), .ZN(n8162)
         );
  AOI21_X1 U9798 ( .B1(n8469), .B2(n8237), .A(n8162), .ZN(n8163) );
  OAI21_X1 U9799 ( .B1(n8164), .B2(n8251), .A(n8163), .ZN(P2_U3163) );
  XOR2_X1 U9800 ( .A(n8166), .B(n8165), .Z(n8171) );
  AOI22_X1 U9801 ( .A1(n8337), .A2(n8257), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8168) );
  NAND2_X1 U9802 ( .A1(n8262), .A2(n8340), .ZN(n8167) );
  OAI211_X1 U9803 ( .C1(n8361), .C2(n8260), .A(n8168), .B(n8167), .ZN(n8169)
         );
  AOI21_X1 U9804 ( .B1(n8513), .B2(n8237), .A(n8169), .ZN(n8170) );
  OAI21_X1 U9805 ( .B1(n8171), .B2(n8251), .A(n8170), .ZN(P2_U3165) );
  XNOR2_X1 U9806 ( .A(n8172), .B(n8274), .ZN(n8173) );
  XNOR2_X1 U9807 ( .A(n8174), .B(n8173), .ZN(n8183) );
  NAND2_X1 U9808 ( .A1(n8262), .A2(n8175), .ZN(n8178) );
  NAND2_X1 U9809 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n10336) );
  INV_X1 U9810 ( .A(n10336), .ZN(n8176) );
  AOI21_X1 U9811 ( .B1(n8257), .B2(n8428), .A(n8176), .ZN(n8177) );
  OAI211_X1 U9812 ( .C1(n8179), .C2(n8260), .A(n8178), .B(n8177), .ZN(n8180)
         );
  AOI21_X1 U9813 ( .B1(n8181), .B2(n8237), .A(n8180), .ZN(n8182) );
  OAI21_X1 U9814 ( .B1(n8183), .B2(n8251), .A(n8182), .ZN(P2_U3166) );
  XOR2_X1 U9815 ( .A(n8146), .B(n8228), .Z(n8190) );
  NAND2_X1 U9816 ( .A1(n8262), .A2(n8184), .ZN(n8186) );
  AOI22_X1 U9817 ( .A1(n8257), .A2(n8412), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3151), .ZN(n8185) );
  OAI211_X1 U9818 ( .C1(n8187), .C2(n8260), .A(n8186), .B(n8185), .ZN(n8188)
         );
  AOI21_X1 U9819 ( .B1(n8491), .B2(n8237), .A(n8188), .ZN(n8189) );
  OAI21_X1 U9820 ( .B1(n8190), .B2(n8251), .A(n8189), .ZN(P2_U3168) );
  XOR2_X1 U9821 ( .A(n8192), .B(n8191), .Z(n8197) );
  AOI22_X1 U9822 ( .A1(n8350), .A2(n8257), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8194) );
  NAND2_X1 U9823 ( .A1(n8262), .A2(n8354), .ZN(n8193) );
  OAI211_X1 U9824 ( .C1(n8221), .C2(n8260), .A(n8194), .B(n8193), .ZN(n8195)
         );
  AOI21_X1 U9825 ( .B1(n8518), .B2(n8237), .A(n8195), .ZN(n8196) );
  OAI21_X1 U9826 ( .B1(n8197), .B2(n8251), .A(n8196), .ZN(P2_U3169) );
  XOR2_X1 U9827 ( .A(n8198), .B(n8199), .Z(n8205) );
  NAND2_X1 U9828 ( .A1(n8262), .A2(n8403), .ZN(n8201) );
  AOI22_X1 U9829 ( .A1(n8257), .A2(n6208), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8200) );
  OAI211_X1 U9830 ( .C1(n8202), .C2(n8260), .A(n8201), .B(n8200), .ZN(n8203)
         );
  AOI21_X1 U9831 ( .B1(n8534), .B2(n8237), .A(n8203), .ZN(n8204) );
  OAI21_X1 U9832 ( .B1(n8205), .B2(n8251), .A(n8204), .ZN(P2_U3173) );
  NOR2_X1 U9833 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8206), .ZN(n10281) );
  AOI21_X1 U9834 ( .B1(n8257), .B2(n8276), .A(n10281), .ZN(n8208) );
  NAND2_X1 U9835 ( .A1(n8244), .A2(n8278), .ZN(n8207) );
  OAI211_X1 U9836 ( .C1(n8210), .C2(n8209), .A(n8208), .B(n8207), .ZN(n8216)
         );
  XNOR2_X1 U9837 ( .A(n8211), .B(n8277), .ZN(n8212) );
  XNOR2_X1 U9838 ( .A(n8213), .B(n8212), .ZN(n8214) );
  NOR2_X1 U9839 ( .A1(n8214), .A2(n8251), .ZN(n8215) );
  AOI211_X1 U9840 ( .C1(n8217), .C2(n8237), .A(n8216), .B(n8215), .ZN(n8218)
         );
  INV_X1 U9841 ( .A(n8218), .ZN(P2_U3174) );
  XOR2_X1 U9842 ( .A(n8220), .B(n8219), .Z(n8227) );
  NOR2_X1 U9843 ( .A1(n8246), .A2(n8221), .ZN(n8224) );
  INV_X1 U9844 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9080) );
  OAI22_X1 U9845 ( .A1(n8260), .A2(n8222), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9080), .ZN(n8223) );
  AOI211_X1 U9846 ( .C1(n8371), .C2(n8262), .A(n8224), .B(n8223), .ZN(n8226)
         );
  NAND2_X1 U9847 ( .A1(n8463), .A2(n8237), .ZN(n8225) );
  OAI211_X1 U9848 ( .C1(n8227), .C2(n8251), .A(n8226), .B(n8225), .ZN(P2_U3175) );
  NAND2_X1 U9849 ( .A1(n8146), .A2(n8228), .ZN(n8230) );
  NAND2_X1 U9850 ( .A1(n8230), .A2(n8229), .ZN(n8231) );
  XOR2_X1 U9851 ( .A(n8232), .B(n8231), .Z(n8239) );
  NAND2_X1 U9852 ( .A1(n8262), .A2(n8431), .ZN(n8234) );
  AOI22_X1 U9853 ( .A1(n8257), .A2(n8426), .B1(P2_REG3_REG_18__SCAN_IN), .B2(
        P2_U3151), .ZN(n8233) );
  OAI211_X1 U9854 ( .C1(n8235), .C2(n8260), .A(n8234), .B(n8233), .ZN(n8236)
         );
  AOI21_X1 U9855 ( .B1(n8435), .B2(n8237), .A(n8236), .ZN(n8238) );
  OAI21_X1 U9856 ( .B1(n8239), .B2(n8251), .A(n8238), .ZN(P2_U3178) );
  XNOR2_X1 U9857 ( .A(n8240), .B(n8241), .ZN(n8243) );
  NAND2_X1 U9858 ( .A1(n8243), .A2(n8242), .ZN(n8249) );
  AOI22_X1 U9859 ( .A1(n8350), .A2(n8244), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8245) );
  OAI21_X1 U9860 ( .B1(n8327), .B2(n8246), .A(n8245), .ZN(n8247) );
  AOI21_X1 U9861 ( .B1(n8330), .B2(n8262), .A(n8247), .ZN(n8248) );
  OAI211_X1 U9862 ( .C1(n8508), .C2(n8266), .A(n8249), .B(n8248), .ZN(P2_U3180) );
  INV_X1 U9863 ( .A(n8250), .ZN(n8267) );
  AOI21_X1 U9864 ( .B1(n8253), .B2(n8252), .A(n8251), .ZN(n8255) );
  NAND2_X1 U9865 ( .A1(n8255), .A2(n8254), .ZN(n8265) );
  INV_X1 U9866 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8256) );
  NOR2_X1 U9867 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8256), .ZN(n10314) );
  AOI21_X1 U9868 ( .B1(n8257), .B2(n8274), .A(n10314), .ZN(n8258) );
  OAI21_X1 U9869 ( .B1(n8260), .B2(n8259), .A(n8258), .ZN(n8261) );
  AOI21_X1 U9870 ( .B1(n8263), .B2(n8262), .A(n8261), .ZN(n8264) );
  OAI211_X1 U9871 ( .C1(n8267), .C2(n8266), .A(n8265), .B(n8264), .ZN(P2_U3181) );
  MUX2_X1 U9872 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8268), .S(n8283), .Z(
        P2_U3522) );
  MUX2_X1 U9873 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8269), .S(n8283), .Z(
        P2_U3521) );
  MUX2_X1 U9874 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8270), .S(n8283), .Z(
        P2_U3520) );
  MUX2_X1 U9875 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8271), .S(n8283), .Z(
        P2_U3519) );
  MUX2_X1 U9876 ( .A(n8272), .B(P2_DATAO_REG_27__SCAN_IN), .S(n9946), .Z(
        P2_U3518) );
  MUX2_X1 U9877 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8337), .S(n8283), .Z(
        P2_U3517) );
  MUX2_X1 U9878 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8350), .S(n8283), .Z(
        P2_U3516) );
  MUX2_X1 U9879 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8338), .S(n8283), .Z(
        P2_U3515) );
  MUX2_X1 U9880 ( .A(n8369), .B(P2_DATAO_REG_23__SCAN_IN), .S(n9946), .Z(
        P2_U3514) );
  MUX2_X1 U9881 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8273), .S(n8283), .Z(
        P2_U3513) );
  MUX2_X1 U9882 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n6208), .S(n8283), .Z(
        P2_U3512) );
  MUX2_X1 U9883 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8413), .S(n8283), .Z(
        P2_U3511) );
  MUX2_X1 U9884 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8426), .S(n8283), .Z(
        P2_U3510) );
  MUX2_X1 U9885 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8412), .S(n8283), .Z(
        P2_U3509) );
  MUX2_X1 U9886 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8428), .S(n8283), .Z(
        P2_U3508) );
  MUX2_X1 U9887 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8274), .S(n8283), .Z(
        P2_U3507) );
  MUX2_X1 U9888 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8275), .S(n8283), .Z(
        P2_U3506) );
  MUX2_X1 U9889 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8276), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U9890 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8277), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U9891 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8278), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U9892 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8279), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U9893 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8280), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U9894 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8281), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U9895 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8282), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U9896 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8284), .S(n8283), .Z(
        P2_U3498) );
  MUX2_X1 U9897 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8285), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U9898 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8286), .S(P2_U3893), .Z(
        P2_U3496) );
  MUX2_X1 U9899 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8287), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U9900 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8288), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U9901 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8289), .S(P2_U3893), .Z(
        P2_U3493) );
  MUX2_X1 U9902 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n6652), .S(P2_U3893), .Z(
        P2_U3492) );
  MUX2_X1 U9903 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8290), .S(P2_U3893), .Z(
        P2_U3491) );
  INV_X1 U9904 ( .A(n8291), .ZN(n8292) );
  AOI21_X1 U9905 ( .B1(n8294), .B2(n8441), .A(n10381), .ZN(n8296) );
  AOI21_X1 U9906 ( .B1(n10381), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8296), .ZN(
        n8295) );
  OAI21_X1 U9907 ( .B1(n8443), .B2(n10365), .A(n8295), .ZN(P2_U3202) );
  AOI21_X1 U9908 ( .B1(n10381), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8296), .ZN(
        n8297) );
  OAI21_X1 U9909 ( .B1(n8298), .B2(n10365), .A(n8297), .ZN(P2_U3203) );
  NAND2_X1 U9910 ( .A1(n8299), .A2(n4495), .ZN(n8305) );
  OAI22_X1 U9911 ( .A1(n4495), .A2(n8301), .B1(n8300), .B2(n10373), .ZN(n8302)
         );
  AOI21_X1 U9912 ( .B1(n8303), .B2(n8419), .A(n8302), .ZN(n8304) );
  OAI211_X1 U9913 ( .C1(n8306), .C2(n8407), .A(n8305), .B(n8304), .ZN(P2_U3205) );
  NAND2_X1 U9914 ( .A1(n8308), .A2(n8307), .ZN(n8309) );
  NAND2_X1 U9915 ( .A1(n8309), .A2(n8312), .ZN(n8310) );
  NAND2_X1 U9916 ( .A1(n8311), .A2(n8310), .ZN(n8505) );
  XNOR2_X1 U9917 ( .A(n8313), .B(n8312), .ZN(n8314) );
  OAI222_X1 U9918 ( .A1(n8391), .A2(n8316), .B1(n8389), .B2(n8315), .C1(n8314), 
        .C2(n8387), .ZN(n8447) );
  NAND2_X1 U9919 ( .A1(n8447), .A2(n4495), .ZN(n8321) );
  NAND2_X1 U9920 ( .A1(n8317), .A2(n8404), .ZN(n8318) );
  OAI21_X1 U9921 ( .B1(n4495), .B2(n9095), .A(n8318), .ZN(n8319) );
  AOI21_X1 U9922 ( .B1(n8448), .B2(n8434), .A(n8319), .ZN(n8320) );
  OAI211_X1 U9923 ( .C1(n8407), .C2(n8505), .A(n8321), .B(n8320), .ZN(P2_U3206) );
  XNOR2_X1 U9924 ( .A(n8322), .B(n8323), .ZN(n8509) );
  XNOR2_X1 U9925 ( .A(n8324), .B(n8323), .ZN(n8325) );
  OAI222_X1 U9926 ( .A1(n8389), .A2(n8327), .B1(n8391), .B2(n8326), .C1(n8387), 
        .C2(n8325), .ZN(n8506) );
  INV_X1 U9927 ( .A(n8506), .ZN(n8328) );
  MUX2_X1 U9928 ( .A(n8329), .B(n8328), .S(n4495), .Z(n8333) );
  AOI22_X1 U9929 ( .A1(n8331), .A2(n8434), .B1(n8404), .B2(n8330), .ZN(n8332)
         );
  OAI211_X1 U9930 ( .C1(n8509), .C2(n8407), .A(n8333), .B(n8332), .ZN(P2_U3207) );
  XNOR2_X1 U9931 ( .A(n8334), .B(n8335), .ZN(n8516) );
  XNOR2_X1 U9932 ( .A(n8336), .B(n8335), .ZN(n8339) );
  AOI222_X1 U9933 ( .A1(n8430), .A2(n8339), .B1(n8338), .B2(n8427), .C1(n8337), 
        .C2(n6321), .ZN(n8512) );
  INV_X1 U9934 ( .A(n8512), .ZN(n8344) );
  INV_X1 U9935 ( .A(n8513), .ZN(n8342) );
  INV_X1 U9936 ( .A(n8340), .ZN(n8341) );
  OAI22_X1 U9937 ( .A1(n8342), .A2(n10370), .B1(n8341), .B2(n10373), .ZN(n8343) );
  OAI21_X1 U9938 ( .B1(n8344), .B2(n8343), .A(n4495), .ZN(n8346) );
  NAND2_X1 U9939 ( .A1(n10381), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8345) );
  OAI211_X1 U9940 ( .C1(n8516), .C2(n8407), .A(n8346), .B(n8345), .ZN(P2_U3208) );
  XNOR2_X1 U9941 ( .A(n8347), .B(n8349), .ZN(n8521) );
  XOR2_X1 U9942 ( .A(n8349), .B(n8348), .Z(n8351) );
  AOI222_X1 U9943 ( .A1(n8430), .A2(n8351), .B1(n8369), .B2(n8427), .C1(n8350), 
        .C2(n6321), .ZN(n8517) );
  OAI21_X1 U9944 ( .B1(n8352), .B2(n10370), .A(n8517), .ZN(n8353) );
  NAND2_X1 U9945 ( .A1(n8353), .A2(n4495), .ZN(n8356) );
  AOI22_X1 U9946 ( .A1(n10381), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8404), .B2(
        n8354), .ZN(n8355) );
  OAI211_X1 U9947 ( .C1(n8521), .C2(n8407), .A(n8356), .B(n8355), .ZN(P2_U3209) );
  XNOR2_X1 U9948 ( .A(n8357), .B(n8358), .ZN(n8525) );
  XNOR2_X1 U9949 ( .A(n8359), .B(n8358), .ZN(n8360) );
  OAI222_X1 U9950 ( .A1(n8391), .A2(n8388), .B1(n8389), .B2(n8361), .C1(n8387), 
        .C2(n8360), .ZN(n8459) );
  NAND2_X1 U9951 ( .A1(n8459), .A2(n4495), .ZN(n8367) );
  INV_X1 U9952 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8364) );
  INV_X1 U9953 ( .A(n8362), .ZN(n8363) );
  OAI22_X1 U9954 ( .A1(n4495), .A2(n8364), .B1(n8363), .B2(n10373), .ZN(n8365)
         );
  AOI21_X1 U9955 ( .B1(n8460), .B2(n8434), .A(n8365), .ZN(n8366) );
  OAI211_X1 U9956 ( .C1(n8525), .C2(n8407), .A(n8367), .B(n8366), .ZN(P2_U3210) );
  XNOR2_X1 U9957 ( .A(n8368), .B(n8375), .ZN(n8370) );
  AOI222_X1 U9958 ( .A1(n8430), .A2(n8370), .B1(n8369), .B2(n6321), .C1(n6208), 
        .C2(n8427), .ZN(n8466) );
  INV_X1 U9959 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8373) );
  INV_X1 U9960 ( .A(n8371), .ZN(n8372) );
  OAI22_X1 U9961 ( .A1(n4495), .A2(n8373), .B1(n8372), .B2(n10373), .ZN(n8374)
         );
  AOI21_X1 U9962 ( .B1(n8463), .B2(n8419), .A(n8374), .ZN(n8379) );
  OR2_X1 U9963 ( .A1(n8376), .A2(n8375), .ZN(n8464) );
  NAND3_X1 U9964 ( .A1(n8464), .A2(n8438), .A3(n8377), .ZN(n8378) );
  OAI211_X1 U9965 ( .C1(n8466), .C2(n10381), .A(n8379), .B(n8378), .ZN(
        P2_U3211) );
  NAND2_X1 U9966 ( .A1(n8381), .A2(n8380), .ZN(n8383) );
  XNOR2_X1 U9967 ( .A(n8383), .B(n8382), .ZN(n8530) );
  XNOR2_X1 U9968 ( .A(n8385), .B(n8384), .ZN(n8386) );
  OAI222_X1 U9969 ( .A1(n8391), .A2(n8390), .B1(n8389), .B2(n8388), .C1(n8387), 
        .C2(n8386), .ZN(n8468) );
  NAND2_X1 U9970 ( .A1(n8468), .A2(n4495), .ZN(n8397) );
  INV_X1 U9971 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8394) );
  INV_X1 U9972 ( .A(n8392), .ZN(n8393) );
  OAI22_X1 U9973 ( .A1(n4495), .A2(n8394), .B1(n8393), .B2(n10373), .ZN(n8395)
         );
  AOI21_X1 U9974 ( .B1(n8469), .B2(n8434), .A(n8395), .ZN(n8396) );
  OAI211_X1 U9975 ( .C1(n8530), .C2(n8407), .A(n8397), .B(n8396), .ZN(P2_U3212) );
  XOR2_X1 U9976 ( .A(n8400), .B(n8398), .Z(n8537) );
  INV_X1 U9977 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8402) );
  OAI21_X1 U9978 ( .B1(n4518), .B2(n8400), .A(n8399), .ZN(n8401) );
  AOI222_X1 U9979 ( .A1(n8430), .A2(n8401), .B1(n8426), .B2(n8427), .C1(n6208), 
        .C2(n6321), .ZN(n8531) );
  MUX2_X1 U9980 ( .A(n8402), .B(n8531), .S(n4495), .Z(n8406) );
  AOI22_X1 U9981 ( .A1(n8534), .A2(n8419), .B1(n8404), .B2(n8403), .ZN(n8405)
         );
  OAI211_X1 U9982 ( .C1(n8537), .C2(n8407), .A(n8406), .B(n8405), .ZN(P2_U3213) );
  NAND2_X1 U9983 ( .A1(n8408), .A2(n8420), .ZN(n8409) );
  NAND2_X1 U9984 ( .A1(n8409), .A2(n8430), .ZN(n8410) );
  OR2_X1 U9985 ( .A1(n8411), .A2(n8410), .ZN(n8415) );
  AOI22_X1 U9986 ( .A1(n8413), .A2(n6321), .B1(n8427), .B2(n8412), .ZN(n8414)
         );
  NAND2_X1 U9987 ( .A1(n8415), .A2(n8414), .ZN(n8482) );
  INV_X1 U9988 ( .A(n8482), .ZN(n8424) );
  INV_X1 U9989 ( .A(n8416), .ZN(n8417) );
  OAI22_X1 U9990 ( .A1(n4495), .A2(n5885), .B1(n8417), .B2(n10373), .ZN(n8418)
         );
  AOI21_X1 U9991 ( .B1(n8476), .B2(n8419), .A(n8418), .ZN(n8423) );
  OR2_X1 U9992 ( .A1(n8421), .A2(n8420), .ZN(n8478) );
  NAND3_X1 U9993 ( .A1(n8478), .A2(n8438), .A3(n8477), .ZN(n8422) );
  OAI211_X1 U9994 ( .C1(n8424), .C2(n10381), .A(n8423), .B(n8422), .ZN(
        P2_U3214) );
  XOR2_X1 U9995 ( .A(n8425), .B(n8437), .Z(n8429) );
  AOI222_X1 U9996 ( .A1(n8430), .A2(n8429), .B1(n8428), .B2(n8427), .C1(n8426), 
        .C2(n6321), .ZN(n8488) );
  INV_X1 U9997 ( .A(n8431), .ZN(n8432) );
  OAI22_X1 U9998 ( .A1(n4495), .A2(n9114), .B1(n8432), .B2(n10373), .ZN(n8433)
         );
  AOI21_X1 U9999 ( .B1(n8435), .B2(n8434), .A(n8433), .ZN(n8440) );
  NAND2_X1 U10000 ( .A1(n8436), .A2(n8437), .ZN(n8485) );
  NAND3_X1 U10001 ( .A1(n8486), .A2(n8485), .A3(n8438), .ZN(n8439) );
  OAI211_X1 U10002 ( .C1(n8488), .C2(n10381), .A(n8440), .B(n8439), .ZN(
        P2_U3215) );
  NAND2_X1 U10003 ( .A1(n10446), .A2(n8496), .ZN(n8444) );
  NAND2_X1 U10004 ( .A1(n10444), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8442) );
  OAI211_X1 U10005 ( .C1(n8443), .C2(n8451), .A(n8444), .B(n8442), .ZN(
        P2_U3490) );
  INV_X1 U10006 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8446) );
  NAND2_X1 U10007 ( .A1(n8498), .A2(n8473), .ZN(n8445) );
  OAI211_X1 U10008 ( .C1(n10446), .C2(n8446), .A(n8445), .B(n8444), .ZN(
        P2_U3489) );
  INV_X1 U10009 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8449) );
  AOI21_X1 U10010 ( .B1(n10429), .B2(n8448), .A(n8447), .ZN(n8502) );
  OAI21_X1 U10011 ( .B1(n8493), .B2(n8505), .A(n8450), .ZN(P2_U3486) );
  MUX2_X1 U10012 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8506), .S(n10446), .Z(
        n8453) );
  OAI22_X1 U10013 ( .A1(n8509), .A2(n8493), .B1(n8508), .B2(n8451), .ZN(n8452)
         );
  OR2_X1 U10014 ( .A1(n8453), .A2(n8452), .ZN(P2_U3485) );
  MUX2_X1 U10015 ( .A(n8886), .B(n8512), .S(n10446), .Z(n8455) );
  NAND2_X1 U10016 ( .A1(n8513), .A2(n8473), .ZN(n8454) );
  OAI211_X1 U10017 ( .C1(n8516), .C2(n8493), .A(n8455), .B(n8454), .ZN(
        P2_U3484) );
  INV_X1 U10018 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8456) );
  MUX2_X1 U10019 ( .A(n8456), .B(n8517), .S(n10446), .Z(n8458) );
  NAND2_X1 U10020 ( .A1(n8518), .A2(n8473), .ZN(n8457) );
  OAI211_X1 U10021 ( .C1(n8493), .C2(n8521), .A(n8458), .B(n8457), .ZN(
        P2_U3483) );
  INV_X1 U10022 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8461) );
  AOI21_X1 U10023 ( .B1(n10429), .B2(n8460), .A(n8459), .ZN(n8522) );
  MUX2_X1 U10024 ( .A(n8461), .B(n8522), .S(n10446), .Z(n8462) );
  OAI21_X1 U10025 ( .B1(n8525), .B2(n8493), .A(n8462), .ZN(P2_U3482) );
  INV_X1 U10026 ( .A(n8463), .ZN(n8467) );
  NAND3_X1 U10027 ( .A1(n8464), .A2(n8377), .A3(n10408), .ZN(n8465) );
  OAI211_X1 U10028 ( .C1(n8467), .C2(n10418), .A(n8466), .B(n8465), .ZN(n8526)
         );
  MUX2_X1 U10029 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8526), .S(n10446), .Z(
        P2_U3481) );
  INV_X1 U10030 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8470) );
  AOI21_X1 U10031 ( .B1(n10429), .B2(n8469), .A(n8468), .ZN(n8527) );
  MUX2_X1 U10032 ( .A(n8470), .B(n8527), .S(n10446), .Z(n8471) );
  OAI21_X1 U10033 ( .B1(n8493), .B2(n8530), .A(n8471), .ZN(P2_U3480) );
  INV_X1 U10034 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8472) );
  MUX2_X1 U10035 ( .A(n8472), .B(n8531), .S(n10446), .Z(n8475) );
  NAND2_X1 U10036 ( .A1(n8534), .A2(n8473), .ZN(n8474) );
  OAI211_X1 U10037 ( .C1(n8537), .C2(n8493), .A(n8475), .B(n8474), .ZN(
        P2_U3479) );
  INV_X1 U10038 ( .A(n8476), .ZN(n8480) );
  NAND3_X1 U10039 ( .A1(n8478), .A2(n8477), .A3(n10408), .ZN(n8479) );
  OAI21_X1 U10040 ( .B1(n8480), .B2(n10418), .A(n8479), .ZN(n8481) );
  NOR2_X1 U10041 ( .A1(n8482), .A2(n8481), .ZN(n8538) );
  MUX2_X1 U10042 ( .A(n8483), .B(n8538), .S(n10446), .Z(n8484) );
  INV_X1 U10043 ( .A(n8484), .ZN(P2_U3478) );
  NAND3_X1 U10044 ( .A1(n8486), .A2(n10408), .A3(n8485), .ZN(n8487) );
  OAI211_X1 U10045 ( .C1(n8489), .C2(n10418), .A(n8488), .B(n8487), .ZN(n8541)
         );
  MUX2_X1 U10046 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8541), .S(n10446), .Z(
        P2_U3477) );
  AOI21_X1 U10047 ( .B1(n10429), .B2(n8491), .A(n8490), .ZN(n8542) );
  MUX2_X1 U10048 ( .A(n8964), .B(n8542), .S(n10446), .Z(n8492) );
  OAI21_X1 U10049 ( .B1(n8545), .B2(n8493), .A(n8492), .ZN(P2_U3476) );
  MUX2_X1 U10050 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n8494), .S(n10446), .Z(
        P2_U3459) );
  NAND2_X1 U10051 ( .A1(n8495), .A2(n8533), .ZN(n8497) );
  NAND2_X1 U10052 ( .A1(n10430), .A2(n8496), .ZN(n8499) );
  OAI211_X1 U10053 ( .C1(n7899), .C2(n10430), .A(n8497), .B(n8499), .ZN(
        P2_U3458) );
  INV_X1 U10054 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8501) );
  NAND2_X1 U10055 ( .A1(n8498), .A2(n8533), .ZN(n8500) );
  OAI211_X1 U10056 ( .C1(n8501), .C2(n10430), .A(n8500), .B(n8499), .ZN(
        P2_U3457) );
  INV_X1 U10057 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8503) );
  OAI21_X1 U10058 ( .B1(n8505), .B2(n8544), .A(n8504), .ZN(P2_U3454) );
  MUX2_X1 U10059 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8506), .S(n10430), .Z(
        n8511) );
  OAI22_X1 U10060 ( .A1(n8509), .A2(n8544), .B1(n8508), .B2(n8507), .ZN(n8510)
         );
  OR2_X1 U10061 ( .A1(n8511), .A2(n8510), .ZN(P2_U3453) );
  MUX2_X1 U10062 ( .A(n8916), .B(n8512), .S(n10430), .Z(n8515) );
  NAND2_X1 U10063 ( .A1(n8513), .A2(n8533), .ZN(n8514) );
  OAI211_X1 U10064 ( .C1(n8516), .C2(n8544), .A(n8515), .B(n8514), .ZN(
        P2_U3452) );
  MUX2_X1 U10065 ( .A(n8928), .B(n8517), .S(n10430), .Z(n8520) );
  NAND2_X1 U10066 ( .A1(n8518), .A2(n8533), .ZN(n8519) );
  OAI211_X1 U10067 ( .C1(n8521), .C2(n8544), .A(n8520), .B(n8519), .ZN(
        P2_U3451) );
  MUX2_X1 U10068 ( .A(n8523), .B(n8522), .S(n10430), .Z(n8524) );
  OAI21_X1 U10069 ( .B1(n8525), .B2(n8544), .A(n8524), .ZN(P2_U3450) );
  MUX2_X1 U10070 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8526), .S(n10430), .Z(
        P2_U3449) );
  MUX2_X1 U10071 ( .A(n8528), .B(n8527), .S(n10430), .Z(n8529) );
  OAI21_X1 U10072 ( .B1(n8530), .B2(n8544), .A(n8529), .ZN(P2_U3448) );
  MUX2_X1 U10073 ( .A(n8532), .B(n8531), .S(n10430), .Z(n8536) );
  NAND2_X1 U10074 ( .A1(n8534), .A2(n8533), .ZN(n8535) );
  OAI211_X1 U10075 ( .C1(n8537), .C2(n8544), .A(n8536), .B(n8535), .ZN(
        P2_U3447) );
  INV_X1 U10076 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8539) );
  MUX2_X1 U10077 ( .A(n8539), .B(n8538), .S(n10430), .Z(n8540) );
  INV_X1 U10078 ( .A(n8540), .ZN(P2_U3446) );
  MUX2_X1 U10079 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8541), .S(n10430), .Z(
        P2_U3444) );
  MUX2_X1 U10080 ( .A(n8788), .B(n8542), .S(n10430), .Z(n8543) );
  OAI21_X1 U10081 ( .B1(n8545), .B2(n8544), .A(n8543), .ZN(P2_U3441) );
  INV_X1 U10082 ( .A(n8546), .ZN(n9936) );
  INV_X1 U10083 ( .A(n8547), .ZN(n8548) );
  NOR4_X1 U10084 ( .A1(n8548), .A2(P2_IR_REG_30__SCAN_IN), .A3(n4674), .A4(
        P2_U3151), .ZN(n8549) );
  AOI21_X1 U10085 ( .B1(n8560), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8549), .ZN(
        n8550) );
  OAI21_X1 U10086 ( .B1(n9936), .B2(n8562), .A(n8550), .ZN(P2_U3264) );
  AOI21_X1 U10087 ( .B1(n8560), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n8556), .ZN(
        n8557) );
  OAI21_X1 U10088 ( .B1(n8558), .B2(n8562), .A(n8557), .ZN(P2_U3267) );
  AOI21_X1 U10089 ( .B1(n8560), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n8559), .ZN(
        n8561) );
  OAI21_X1 U10090 ( .B1(n8563), .B2(n8562), .A(n8561), .ZN(P2_U3268) );
  MUX2_X1 U10091 ( .A(n8564), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10092 ( .A(n8565), .ZN(n8566) );
  NAND2_X1 U10093 ( .A1(n8569), .A2(n8568), .ZN(n8572) );
  AOI22_X1 U10094 ( .A1(n9263), .A2(n8727), .B1(n8733), .B2(n9505), .ZN(n8570)
         );
  XNOR2_X1 U10095 ( .A(n8570), .B(n7517), .ZN(n8571) );
  NOR2_X2 U10096 ( .A1(n8572), .A2(n8571), .ZN(n8680) );
  OAI22_X1 U10097 ( .A1(n9930), .A2(n8728), .B1(n9262), .B2(n4503), .ZN(n8681)
         );
  NAND2_X1 U10098 ( .A1(n8572), .A2(n8571), .ZN(n8678) );
  INV_X1 U10099 ( .A(n8577), .ZN(n8575) );
  AOI22_X1 U10100 ( .A1(n9218), .A2(n8727), .B1(n8655), .B2(n9503), .ZN(n8573)
         );
  XNOR2_X1 U10101 ( .A(n8573), .B(n7517), .ZN(n8576) );
  INV_X1 U10102 ( .A(n8576), .ZN(n8574) );
  NAND2_X1 U10103 ( .A1(n8575), .A2(n8574), .ZN(n8578) );
  OAI22_X1 U10104 ( .A1(n9978), .A2(n8728), .B1(n8579), .B2(n4503), .ZN(n9209)
         );
  INV_X1 U10105 ( .A(n9209), .ZN(n8580) );
  AOI22_X1 U10106 ( .A1(n9796), .A2(n8727), .B1(n8733), .B2(n9502), .ZN(n8582)
         );
  XOR2_X1 U10107 ( .A(n7517), .B(n8582), .Z(n8584) );
  OAI22_X1 U10108 ( .A1(n9925), .A2(n8728), .B1(n9142), .B2(n4503), .ZN(n8583)
         );
  NOR2_X1 U10109 ( .A1(n8584), .A2(n8583), .ZN(n8589) );
  AOI21_X1 U10110 ( .B1(n8584), .B2(n8583), .A(n8589), .ZN(n8771) );
  NAND2_X1 U10111 ( .A1(n9333), .A2(n8727), .ZN(n8586) );
  NAND2_X1 U10112 ( .A1(n9501), .A2(n8733), .ZN(n8585) );
  NAND2_X1 U10113 ( .A1(n8586), .A2(n8585), .ZN(n8588) );
  XNOR2_X1 U10114 ( .A(n8588), .B(n7517), .ZN(n8594) );
  AOI22_X1 U10115 ( .A1(n9333), .A2(n8655), .B1(n8653), .B2(n9501), .ZN(n8592)
         );
  XNOR2_X1 U10116 ( .A(n8594), .B(n8592), .ZN(n9139) );
  AND2_X1 U10117 ( .A1(n8771), .A2(n9139), .ZN(n8591) );
  INV_X1 U10118 ( .A(n9139), .ZN(n8590) );
  INV_X1 U10119 ( .A(n8589), .ZN(n9135) );
  INV_X1 U10120 ( .A(n8592), .ZN(n8593) );
  NAND2_X1 U10121 ( .A1(n9765), .A2(n8727), .ZN(n8597) );
  NAND2_X1 U10122 ( .A1(n9500), .A2(n8655), .ZN(n8596) );
  NAND2_X1 U10123 ( .A1(n8597), .A2(n8596), .ZN(n8598) );
  XNOR2_X1 U10124 ( .A(n8598), .B(n7517), .ZN(n8602) );
  NAND2_X1 U10125 ( .A1(n9765), .A2(n8655), .ZN(n8600) );
  NAND2_X1 U10126 ( .A1(n9500), .A2(n8653), .ZN(n8599) );
  NAND2_X1 U10127 ( .A1(n8600), .A2(n8599), .ZN(n8601) );
  NOR2_X1 U10128 ( .A1(n8602), .A2(n8601), .ZN(n9179) );
  NAND2_X1 U10129 ( .A1(n8602), .A2(n8601), .ZN(n9180) );
  NAND2_X1 U10130 ( .A1(n9748), .A2(n8727), .ZN(n8604) );
  NAND2_X1 U10131 ( .A1(n9499), .A2(n8733), .ZN(n8603) );
  NAND2_X1 U10132 ( .A1(n8604), .A2(n8603), .ZN(n8605) );
  XNOR2_X1 U10133 ( .A(n8605), .B(n8731), .ZN(n8608) );
  AND2_X1 U10134 ( .A1(n9499), .A2(n8653), .ZN(n8606) );
  AOI21_X1 U10135 ( .B1(n9748), .B2(n8655), .A(n8606), .ZN(n8607) );
  NOR2_X1 U10136 ( .A1(n8608), .A2(n8607), .ZN(n8717) );
  NAND2_X1 U10137 ( .A1(n8608), .A2(n8607), .ZN(n8715) );
  OAI22_X1 U10138 ( .A1(n9913), .A2(n8609), .B1(n8720), .B2(n8728), .ZN(n8610)
         );
  XNOR2_X1 U10139 ( .A(n8610), .B(n7517), .ZN(n8612) );
  OAI22_X1 U10140 ( .A1(n9913), .A2(n8728), .B1(n8720), .B2(n4503), .ZN(n8611)
         );
  NOR2_X1 U10141 ( .A1(n8612), .A2(n8611), .ZN(n8613) );
  AOI21_X1 U10142 ( .B1(n8612), .B2(n8611), .A(n8613), .ZN(n9161) );
  NAND2_X1 U10143 ( .A1(n9160), .A2(n9161), .ZN(n9159) );
  INV_X1 U10144 ( .A(n8613), .ZN(n8614) );
  NAND2_X1 U10145 ( .A1(n9159), .A2(n8614), .ZN(n8753) );
  NAND2_X1 U10146 ( .A1(n9715), .A2(n8727), .ZN(n8616) );
  NAND2_X1 U10147 ( .A1(n9497), .A2(n8655), .ZN(n8615) );
  NAND2_X1 U10148 ( .A1(n8616), .A2(n8615), .ZN(n8617) );
  XNOR2_X1 U10149 ( .A(n8617), .B(n4493), .ZN(n8620) );
  AOI22_X1 U10150 ( .A1(n9715), .A2(n8733), .B1(n8653), .B2(n9497), .ZN(n8618)
         );
  XNOR2_X1 U10151 ( .A(n8620), .B(n8618), .ZN(n8754) );
  NAND2_X1 U10152 ( .A1(n8753), .A2(n8754), .ZN(n8752) );
  INV_X1 U10153 ( .A(n8618), .ZN(n8619) );
  AOI22_X1 U10154 ( .A1(n9703), .A2(n8727), .B1(n8655), .B2(n9496), .ZN(n8622)
         );
  XNOR2_X1 U10155 ( .A(n8622), .B(n4493), .ZN(n8623) );
  NAND2_X2 U10156 ( .A1(n8624), .A2(n8623), .ZN(n8693) );
  OAI22_X1 U10157 ( .A1(n9905), .A2(n8728), .B1(n8626), .B2(n4503), .ZN(n9170)
         );
  NAND2_X1 U10158 ( .A1(n9690), .A2(n8727), .ZN(n8629) );
  OR2_X1 U10159 ( .A1(n9171), .A2(n8728), .ZN(n8628) );
  NAND2_X1 U10160 ( .A1(n8629), .A2(n8628), .ZN(n8630) );
  XNOR2_X1 U10161 ( .A(n8630), .B(n8731), .ZN(n8634) );
  NOR2_X1 U10162 ( .A1(n9171), .A2(n4503), .ZN(n8631) );
  AOI21_X1 U10163 ( .B1(n9690), .B2(n8655), .A(n8631), .ZN(n8633) );
  OR2_X1 U10164 ( .A1(n8634), .A2(n8633), .ZN(n8691) );
  INV_X1 U10165 ( .A(n8691), .ZN(n8636) );
  OR2_X1 U10166 ( .A1(n9170), .A2(n8636), .ZN(n8632) );
  NAND2_X1 U10167 ( .A1(n8634), .A2(n8633), .ZN(n9148) );
  NAND2_X1 U10168 ( .A1(n9671), .A2(n8727), .ZN(n8638) );
  NAND2_X1 U10169 ( .A1(n9494), .A2(n8655), .ZN(n8637) );
  NAND2_X1 U10170 ( .A1(n8638), .A2(n8637), .ZN(n8639) );
  XNOR2_X1 U10171 ( .A(n8639), .B(n8731), .ZN(n8641) );
  AND2_X1 U10172 ( .A1(n9494), .A2(n8653), .ZN(n8640) );
  AOI21_X1 U10173 ( .B1(n9671), .B2(n8655), .A(n8640), .ZN(n8642) );
  NAND2_X1 U10174 ( .A1(n8641), .A2(n8642), .ZN(n8646) );
  INV_X1 U10175 ( .A(n8641), .ZN(n8644) );
  INV_X1 U10176 ( .A(n8642), .ZN(n8643) );
  NAND2_X1 U10177 ( .A1(n8644), .A2(n8643), .ZN(n8645) );
  AND2_X1 U10178 ( .A1(n8646), .A2(n8645), .ZN(n9149) );
  NAND2_X1 U10179 ( .A1(n9656), .A2(n8727), .ZN(n8648) );
  NAND2_X1 U10180 ( .A1(n9493), .A2(n8655), .ZN(n8647) );
  NAND2_X1 U10181 ( .A1(n8648), .A2(n8647), .ZN(n8649) );
  XNOR2_X1 U10182 ( .A(n8649), .B(n4493), .ZN(n8656) );
  AOI22_X1 U10183 ( .A1(n9656), .A2(n8733), .B1(n8653), .B2(n9493), .ZN(n8657)
         );
  XNOR2_X1 U10184 ( .A(n8656), .B(n8657), .ZN(n8762) );
  NAND2_X1 U10185 ( .A1(n8761), .A2(n8762), .ZN(n8760) );
  NAND2_X1 U10186 ( .A1(n9639), .A2(n8727), .ZN(n8651) );
  NAND2_X1 U10187 ( .A1(n9492), .A2(n8733), .ZN(n8650) );
  NAND2_X1 U10188 ( .A1(n8651), .A2(n8650), .ZN(n8652) );
  XNOR2_X1 U10189 ( .A(n8652), .B(n4493), .ZN(n8662) );
  AND2_X1 U10190 ( .A1(n9492), .A2(n8653), .ZN(n8654) );
  AOI21_X1 U10191 ( .B1(n9639), .B2(n8655), .A(n8654), .ZN(n8660) );
  XNOR2_X1 U10192 ( .A(n8662), .B(n8660), .ZN(n9193) );
  INV_X1 U10193 ( .A(n8656), .ZN(n8658) );
  NAND2_X1 U10194 ( .A1(n8658), .A2(n8657), .ZN(n9194) );
  NAND2_X1 U10195 ( .A1(n8760), .A2(n8659), .ZN(n9192) );
  INV_X1 U10196 ( .A(n8660), .ZN(n8661) );
  NAND2_X1 U10197 ( .A1(n8662), .A2(n8661), .ZN(n8667) );
  AOI22_X1 U10198 ( .A1(n9628), .A2(n8727), .B1(n8655), .B2(n9491), .ZN(n8663)
         );
  XOR2_X1 U10199 ( .A(n4493), .B(n8663), .Z(n8665) );
  OAI22_X1 U10200 ( .A1(n9885), .A2(n8728), .B1(n9196), .B2(n4503), .ZN(n8664)
         );
  NOR2_X1 U10201 ( .A1(n8665), .A2(n8664), .ZN(n8747) );
  AOI21_X1 U10202 ( .B1(n8665), .B2(n8664), .A(n8747), .ZN(n8666) );
  AOI21_X1 U10203 ( .B1(n9192), .B2(n8667), .A(n8666), .ZN(n8671) );
  INV_X1 U10204 ( .A(n8666), .ZN(n8669) );
  INV_X1 U10205 ( .A(n8667), .ZN(n8668) );
  NOR2_X1 U10206 ( .A1(n8669), .A2(n8668), .ZN(n8670) );
  OAI21_X1 U10207 ( .B1(n8671), .B2(n8739), .A(n9966), .ZN(n8677) );
  INV_X1 U10208 ( .A(n8672), .ZN(n9625) );
  OAI22_X1 U10209 ( .A1(n8673), .A2(n9141), .B1(n8736), .B2(n9195), .ZN(n9620)
         );
  AOI22_X1 U10210 ( .A1(n9620), .A2(n9960), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n8674) );
  OAI21_X1 U10211 ( .B1(n9970), .B2(n9625), .A(n8674), .ZN(n8675) );
  AOI21_X1 U10212 ( .B1(n9628), .B2(n9217), .A(n8675), .ZN(n8676) );
  NAND2_X1 U10213 ( .A1(n8677), .A2(n8676), .ZN(P1_U3214) );
  INV_X1 U10214 ( .A(n8678), .ZN(n8679) );
  NOR2_X1 U10215 ( .A1(n8680), .A2(n8679), .ZN(n8682) );
  XNOR2_X1 U10216 ( .A(n8682), .B(n8681), .ZN(n8689) );
  OAI22_X1 U10217 ( .A1(n9214), .A2(n8684), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8683), .ZN(n8686) );
  NOR2_X1 U10218 ( .A1(n9930), .A2(n9963), .ZN(n8685) );
  AOI211_X1 U10219 ( .C1(n8687), .C2(n9211), .A(n8686), .B(n8685), .ZN(n8688)
         );
  OAI21_X1 U10220 ( .B1(n8689), .B2(n9220), .A(n8688), .ZN(P1_U3215) );
  OR2_X1 U10221 ( .A1(n8690), .A2(n9170), .ZN(n8694) );
  INV_X1 U10222 ( .A(n8694), .ZN(n9169) );
  INV_X1 U10223 ( .A(n8693), .ZN(n8692) );
  AND2_X1 U10224 ( .A1(n9148), .A2(n8691), .ZN(n8695) );
  NOR3_X1 U10225 ( .A1(n9169), .A2(n8692), .A3(n8695), .ZN(n8697) );
  NAND2_X1 U10226 ( .A1(n8694), .A2(n8693), .ZN(n8696) );
  OAI21_X1 U10227 ( .B1(n8697), .B2(n9151), .A(n9966), .ZN(n8703) );
  NAND2_X1 U10228 ( .A1(n9496), .A2(n9197), .ZN(n8699) );
  NAND2_X1 U10229 ( .A1(n9494), .A2(n9184), .ZN(n8698) );
  AND2_X1 U10230 ( .A1(n8699), .A2(n8698), .ZN(n9684) );
  OAI22_X1 U10231 ( .A1(n9214), .A2(n9684), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8700), .ZN(n8701) );
  AOI21_X1 U10232 ( .B1(n9681), .B2(n9211), .A(n8701), .ZN(n8702) );
  OAI211_X1 U10233 ( .C1(n9901), .C2(n9963), .A(n8703), .B(n8702), .ZN(
        P1_U3216) );
  AOI22_X1 U10234 ( .A1(n9960), .A2(n8704), .B1(P1_REG3_REG_10__SCAN_IN), .B2(
        P1_U3086), .ZN(n8705) );
  OAI21_X1 U10235 ( .B1(n9970), .B2(n8706), .A(n8705), .ZN(n8712) );
  AOI21_X1 U10236 ( .B1(n8709), .B2(n8708), .A(n8707), .ZN(n8710) );
  NOR2_X1 U10237 ( .A1(n8710), .A2(n9220), .ZN(n8711) );
  AOI211_X1 U10238 ( .C1(n8713), .C2(n9217), .A(n8712), .B(n8711), .ZN(n8714)
         );
  INV_X1 U10239 ( .A(n8714), .ZN(P1_U3217) );
  INV_X1 U10240 ( .A(n8715), .ZN(n8716) );
  NOR2_X1 U10241 ( .A1(n8717), .A2(n8716), .ZN(n8718) );
  XNOR2_X1 U10242 ( .A(n8719), .B(n8718), .ZN(n8726) );
  OAI22_X1 U10243 ( .A1(n8721), .A2(n9141), .B1(n8720), .B2(n9195), .ZN(n9744)
         );
  AOI22_X1 U10244 ( .A1(n9744), .A2(n9960), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        P1_U3086), .ZN(n8722) );
  OAI21_X1 U10245 ( .B1(n9970), .B2(n8723), .A(n8722), .ZN(n8724) );
  AOI21_X1 U10246 ( .B1(n9748), .B2(n9217), .A(n8724), .ZN(n8725) );
  OAI21_X1 U10247 ( .B1(n8726), .B2(n9220), .A(n8725), .ZN(P1_U3219) );
  NAND2_X1 U10248 ( .A1(n8745), .A2(n8727), .ZN(n8730) );
  OR2_X1 U10249 ( .A1(n8736), .A2(n8728), .ZN(n8729) );
  NAND2_X1 U10250 ( .A1(n8730), .A2(n8729), .ZN(n8732) );
  XNOR2_X1 U10251 ( .A(n8732), .B(n8731), .ZN(n8738) );
  NAND2_X1 U10252 ( .A1(n8745), .A2(n8655), .ZN(n8734) );
  OAI21_X1 U10253 ( .B1(n8736), .B2(n4503), .A(n8734), .ZN(n8737) );
  XNOR2_X1 U10254 ( .A(n8738), .B(n8737), .ZN(n8746) );
  NAND3_X1 U10255 ( .A1(n8739), .A2(n9966), .A3(n8746), .ZN(n8750) );
  INV_X1 U10256 ( .A(n8740), .ZN(n8743) );
  AOI22_X1 U10257 ( .A1(n9960), .A2(n8741), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n8742) );
  OAI21_X1 U10258 ( .B1(n9970), .B2(n8743), .A(n8742), .ZN(n8744) );
  AOI21_X1 U10259 ( .B1(n8745), .B2(n9217), .A(n8744), .ZN(n8749) );
  NAND3_X1 U10260 ( .A1(n8747), .A2(n9966), .A3(n8746), .ZN(n8748) );
  NAND4_X1 U10261 ( .A1(n8751), .A2(n8750), .A3(n8749), .A4(n8748), .ZN(
        P1_U3220) );
  OAI21_X1 U10262 ( .B1(n8754), .B2(n8753), .A(n8752), .ZN(n8755) );
  NAND2_X1 U10263 ( .A1(n8755), .A2(n9966), .ZN(n8759) );
  AOI22_X1 U10264 ( .A1(n9197), .A2(n9498), .B1(n9496), .B2(n9184), .ZN(n9713)
         );
  INV_X1 U10265 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8756) );
  OAI22_X1 U10266 ( .A1(n9214), .A2(n9713), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8756), .ZN(n8757) );
  AOI21_X1 U10267 ( .B1(n9721), .B2(n9211), .A(n8757), .ZN(n8758) );
  OAI211_X1 U10268 ( .C1(n9909), .C2(n9963), .A(n8759), .B(n8758), .ZN(
        P1_U3223) );
  OAI21_X1 U10269 ( .B1(n8762), .B2(n8761), .A(n8760), .ZN(n8763) );
  NAND2_X1 U10270 ( .A1(n8763), .A2(n9966), .ZN(n8769) );
  NAND2_X1 U10271 ( .A1(n9494), .A2(n9197), .ZN(n8765) );
  NAND2_X1 U10272 ( .A1(n9492), .A2(n9184), .ZN(n8764) );
  AND2_X1 U10273 ( .A1(n8765), .A2(n8764), .ZN(n9653) );
  OAI22_X1 U10274 ( .A1(n9214), .A2(n9653), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8766), .ZN(n8767) );
  AOI21_X1 U10275 ( .B1(n9657), .B2(n9211), .A(n8767), .ZN(n8768) );
  OAI211_X1 U10276 ( .C1(n9893), .C2(n9963), .A(n8769), .B(n8768), .ZN(
        P1_U3225) );
  NAND2_X1 U10277 ( .A1(n8770), .A2(n8771), .ZN(n9136) );
  OAI21_X1 U10278 ( .B1(n8771), .B2(n8770), .A(n9136), .ZN(n8772) );
  NAND2_X1 U10279 ( .A1(n8772), .A2(n9966), .ZN(n8776) );
  AOI22_X1 U10280 ( .A1(n9197), .A2(n9503), .B1(n9501), .B2(n9184), .ZN(n9792)
         );
  OAI22_X1 U10281 ( .A1(n9214), .A2(n9792), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8773), .ZN(n8774) );
  AOI21_X1 U10282 ( .B1(n9797), .B2(n9211), .A(n8774), .ZN(n8775) );
  OAI211_X1 U10283 ( .C1(n9925), .C2(n9963), .A(n8776), .B(n8775), .ZN(n9134)
         );
  OAI22_X1 U10284 ( .A1(SI_9_), .A2(keyinput253), .B1(keyinput144), .B2(
        P1_REG0_REG_21__SCAN_IN), .ZN(n8777) );
  AOI221_X1 U10285 ( .B1(SI_9_), .B2(keyinput253), .C1(P1_REG0_REG_21__SCAN_IN), .C2(keyinput144), .A(n8777), .ZN(n8784) );
  OAI22_X1 U10286 ( .A1(n5929), .A2(keyinput243), .B1(keyinput215), .B2(
        P1_REG1_REG_26__SCAN_IN), .ZN(n8778) );
  AOI221_X1 U10287 ( .B1(n5929), .B2(keyinput243), .C1(P1_REG1_REG_26__SCAN_IN), .C2(keyinput215), .A(n8778), .ZN(n8783) );
  OAI22_X1 U10288 ( .A1(n10089), .A2(keyinput244), .B1(n5786), .B2(keyinput188), .ZN(n8779) );
  AOI221_X1 U10289 ( .B1(n10089), .B2(keyinput244), .C1(keyinput188), .C2(
        n5786), .A(n8779), .ZN(n8782) );
  INV_X1 U10290 ( .A(SI_5_), .ZN(n9067) );
  OAI22_X1 U10291 ( .A1(n9067), .A2(keyinput234), .B1(n8301), .B2(keyinput146), 
        .ZN(n8780) );
  AOI221_X1 U10292 ( .B1(n9067), .B2(keyinput234), .C1(keyinput146), .C2(n8301), .A(n8780), .ZN(n8781) );
  NAND4_X1 U10293 ( .A1(n8784), .A2(n8783), .A3(n8782), .A4(n8781), .ZN(n8808)
         );
  INV_X1 U10294 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n8786) );
  AOI22_X1 U10295 ( .A1(n8786), .A2(keyinput183), .B1(n9043), .B2(keyinput143), 
        .ZN(n8785) );
  OAI221_X1 U10296 ( .B1(n8786), .B2(keyinput183), .C1(n9043), .C2(keyinput143), .A(n8785), .ZN(n8807) );
  OAI22_X1 U10297 ( .A1(n8788), .A2(keyinput148), .B1(n9037), .B2(keyinput168), 
        .ZN(n8787) );
  AOI221_X1 U10298 ( .B1(n8788), .B2(keyinput148), .C1(keyinput168), .C2(n9037), .A(n8787), .ZN(n8795) );
  INV_X1 U10299 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n9028) );
  XNOR2_X1 U10300 ( .A(n9028), .B(keyinput209), .ZN(n8793) );
  XOR2_X1 U10301 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput242), .Z(n8792) );
  XOR2_X1 U10302 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput224), .Z(n8791) );
  XNOR2_X1 U10303 ( .A(n8789), .B(keyinput192), .ZN(n8790) );
  NOR4_X1 U10304 ( .A1(n8793), .A2(n8792), .A3(n8791), .A4(n8790), .ZN(n8794)
         );
  NAND2_X1 U10305 ( .A1(n8795), .A2(n8794), .ZN(n8806) );
  OAI22_X1 U10306 ( .A1(n5108), .A2(keyinput158), .B1(n9118), .B2(keyinput136), 
        .ZN(n8796) );
  AOI221_X1 U10307 ( .B1(n5108), .B2(keyinput158), .C1(keyinput136), .C2(n9118), .A(n8796), .ZN(n8804) );
  OAI22_X1 U10308 ( .A1(n10094), .A2(keyinput159), .B1(n5310), .B2(keyinput174), .ZN(n8797) );
  AOI221_X1 U10309 ( .B1(n10094), .B2(keyinput159), .C1(keyinput174), .C2(
        n5310), .A(n8797), .ZN(n8803) );
  INV_X1 U10310 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n8965) );
  OAI22_X1 U10311 ( .A1(n7478), .A2(keyinput231), .B1(n8965), .B2(keyinput140), 
        .ZN(n8798) );
  AOI221_X1 U10312 ( .B1(n7478), .B2(keyinput231), .C1(keyinput140), .C2(n8965), .A(n8798), .ZN(n8802) );
  XOR2_X1 U10313 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput171), .Z(n8800) );
  XNOR2_X1 U10314 ( .A(n10176), .B(keyinput245), .ZN(n8799) );
  NOR2_X1 U10315 ( .A1(n8800), .A2(n8799), .ZN(n8801) );
  NAND4_X1 U10316 ( .A1(n8804), .A2(n8803), .A3(n8802), .A4(n8801), .ZN(n8805)
         );
  NOR4_X1 U10317 ( .A1(n8808), .A2(n8807), .A3(n8806), .A4(n8805), .ZN(n8943)
         );
  OAI22_X1 U10318 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(keyinput186), .B1(
        keyinput236), .B2(P1_REG3_REG_9__SCAN_IN), .ZN(n8809) );
  AOI221_X1 U10319 ( .B1(P1_IR_REG_12__SCAN_IN), .B2(keyinput186), .C1(
        P1_REG3_REG_9__SCAN_IN), .C2(keyinput236), .A(n8809), .ZN(n8816) );
  OAI22_X1 U10320 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(keyinput254), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(keyinput179), .ZN(n8810) );
  AOI221_X1 U10321 ( .B1(P1_IR_REG_9__SCAN_IN), .B2(keyinput254), .C1(
        keyinput179), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n8810), .ZN(n8815) );
  OAI22_X1 U10322 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(keyinput226), .B1(
        keyinput205), .B2(P2_ADDR_REG_11__SCAN_IN), .ZN(n8811) );
  AOI221_X1 U10323 ( .B1(P2_IR_REG_4__SCAN_IN), .B2(keyinput226), .C1(
        P2_ADDR_REG_11__SCAN_IN), .C2(keyinput205), .A(n8811), .ZN(n8814) );
  OAI22_X1 U10324 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(keyinput131), .B1(
        keyinput167), .B2(P2_ADDR_REG_8__SCAN_IN), .ZN(n8812) );
  AOI221_X1 U10325 ( .B1(P2_DATAO_REG_0__SCAN_IN), .B2(keyinput131), .C1(
        P2_ADDR_REG_8__SCAN_IN), .C2(keyinput167), .A(n8812), .ZN(n8813) );
  NAND4_X1 U10326 ( .A1(n8816), .A2(n8815), .A3(n8814), .A4(n8813), .ZN(n8844)
         );
  OAI22_X1 U10327 ( .A1(P1_D_REG_4__SCAN_IN), .A2(keyinput137), .B1(
        keyinput151), .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8817) );
  AOI221_X1 U10328 ( .B1(P1_D_REG_4__SCAN_IN), .B2(keyinput137), .C1(
        P1_DATAO_REG_27__SCAN_IN), .C2(keyinput151), .A(n8817), .ZN(n8824) );
  OAI22_X1 U10329 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(keyinput189), .B1(
        keyinput197), .B2(P2_REG3_REG_6__SCAN_IN), .ZN(n8818) );
  AOI221_X1 U10330 ( .B1(P1_IR_REG_4__SCAN_IN), .B2(keyinput189), .C1(
        P2_REG3_REG_6__SCAN_IN), .C2(keyinput197), .A(n8818), .ZN(n8823) );
  OAI22_X1 U10331 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(keyinput162), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput184), .ZN(n8819) );
  AOI221_X1 U10332 ( .B1(P1_DATAO_REG_8__SCAN_IN), .B2(keyinput162), .C1(
        keyinput184), .C2(P2_REG3_REG_18__SCAN_IN), .A(n8819), .ZN(n8822) );
  OAI22_X1 U10333 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(keyinput139), .B1(
        P2_IR_REG_15__SCAN_IN), .B2(keyinput228), .ZN(n8820) );
  AOI221_X1 U10334 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(keyinput139), .C1(
        keyinput228), .C2(P2_IR_REG_15__SCAN_IN), .A(n8820), .ZN(n8821) );
  NAND4_X1 U10335 ( .A1(n8824), .A2(n8823), .A3(n8822), .A4(n8821), .ZN(n8843)
         );
  OAI22_X1 U10336 ( .A1(SI_12_), .A2(keyinput200), .B1(P1_REG2_REG_30__SCAN_IN), .B2(keyinput217), .ZN(n8825) );
  AOI221_X1 U10337 ( .B1(SI_12_), .B2(keyinput200), .C1(keyinput217), .C2(
        P1_REG2_REG_30__SCAN_IN), .A(n8825), .ZN(n8832) );
  OAI22_X1 U10338 ( .A1(P1_REG2_REG_19__SCAN_IN), .A2(keyinput190), .B1(
        P2_IR_REG_31__SCAN_IN), .B2(keyinput246), .ZN(n8826) );
  AOI221_X1 U10339 ( .B1(P1_REG2_REG_19__SCAN_IN), .B2(keyinput190), .C1(
        keyinput246), .C2(P2_IR_REG_31__SCAN_IN), .A(n8826), .ZN(n8831) );
  OAI22_X1 U10340 ( .A1(SI_2_), .A2(keyinput227), .B1(P2_REG0_REG_10__SCAN_IN), 
        .B2(keyinput157), .ZN(n8827) );
  AOI221_X1 U10341 ( .B1(SI_2_), .B2(keyinput227), .C1(keyinput157), .C2(
        P2_REG0_REG_10__SCAN_IN), .A(n8827), .ZN(n8830) );
  OAI22_X1 U10342 ( .A1(P1_REG0_REG_19__SCAN_IN), .A2(keyinput154), .B1(
        keyinput166), .B2(P2_REG0_REG_31__SCAN_IN), .ZN(n8828) );
  AOI221_X1 U10343 ( .B1(P1_REG0_REG_19__SCAN_IN), .B2(keyinput154), .C1(
        P2_REG0_REG_31__SCAN_IN), .C2(keyinput166), .A(n8828), .ZN(n8829) );
  NAND4_X1 U10344 ( .A1(n8832), .A2(n8831), .A3(n8830), .A4(n8829), .ZN(n8842)
         );
  OAI22_X1 U10345 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(keyinput181), .B1(
        keyinput241), .B2(P1_ADDR_REG_16__SCAN_IN), .ZN(n8833) );
  AOI221_X1 U10346 ( .B1(P2_DATAO_REG_16__SCAN_IN), .B2(keyinput181), .C1(
        P1_ADDR_REG_16__SCAN_IN), .C2(keyinput241), .A(n8833), .ZN(n8840) );
  OAI22_X1 U10347 ( .A1(SI_11_), .A2(keyinput145), .B1(P2_DATAO_REG_6__SCAN_IN), .B2(keyinput129), .ZN(n8834) );
  AOI221_X1 U10348 ( .B1(SI_11_), .B2(keyinput145), .C1(keyinput129), .C2(
        P2_DATAO_REG_6__SCAN_IN), .A(n8834), .ZN(n8839) );
  OAI22_X1 U10349 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(keyinput161), .B1(
        keyinput191), .B2(P2_REG0_REG_7__SCAN_IN), .ZN(n8835) );
  AOI221_X1 U10350 ( .B1(P2_IR_REG_3__SCAN_IN), .B2(keyinput161), .C1(
        P2_REG0_REG_7__SCAN_IN), .C2(keyinput191), .A(n8835), .ZN(n8838) );
  OAI22_X1 U10351 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(keyinput210), .B1(
        keyinput176), .B2(P2_REG2_REG_31__SCAN_IN), .ZN(n8836) );
  AOI221_X1 U10352 ( .B1(P1_REG3_REG_19__SCAN_IN), .B2(keyinput210), .C1(
        P2_REG2_REG_31__SCAN_IN), .C2(keyinput176), .A(n8836), .ZN(n8837) );
  NAND4_X1 U10353 ( .A1(n8840), .A2(n8839), .A3(n8838), .A4(n8837), .ZN(n8841)
         );
  NOR4_X1 U10354 ( .A1(n8844), .A2(n8843), .A3(n8842), .A4(n8841), .ZN(n8942)
         );
  OAI22_X1 U10355 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(keyinput160), .B1(
        P2_IR_REG_2__SCAN_IN), .B2(keyinput165), .ZN(n8845) );
  AOI221_X1 U10356 ( .B1(P1_DATAO_REG_26__SCAN_IN), .B2(keyinput160), .C1(
        keyinput165), .C2(P2_IR_REG_2__SCAN_IN), .A(n8845), .ZN(n8852) );
  OAI22_X1 U10357 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(keyinput180), .B1(
        P1_REG2_REG_29__SCAN_IN), .B2(keyinput169), .ZN(n8846) );
  AOI221_X1 U10358 ( .B1(P1_IR_REG_15__SCAN_IN), .B2(keyinput180), .C1(
        keyinput169), .C2(P1_REG2_REG_29__SCAN_IN), .A(n8846), .ZN(n8851) );
  OAI22_X1 U10359 ( .A1(P1_REG1_REG_28__SCAN_IN), .A2(keyinput202), .B1(
        P1_REG0_REG_10__SCAN_IN), .B2(keyinput142), .ZN(n8847) );
  AOI221_X1 U10360 ( .B1(P1_REG1_REG_28__SCAN_IN), .B2(keyinput202), .C1(
        keyinput142), .C2(P1_REG0_REG_10__SCAN_IN), .A(n8847), .ZN(n8850) );
  OAI22_X1 U10361 ( .A1(P1_REG0_REG_20__SCAN_IN), .A2(keyinput196), .B1(
        keyinput135), .B2(P2_REG3_REG_28__SCAN_IN), .ZN(n8848) );
  AOI221_X1 U10362 ( .B1(P1_REG0_REG_20__SCAN_IN), .B2(keyinput196), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput135), .A(n8848), .ZN(n8849) );
  NAND4_X1 U10363 ( .A1(n8852), .A2(n8851), .A3(n8850), .A4(n8849), .ZN(n8880)
         );
  OAI22_X1 U10364 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(keyinput207), .B1(
        P2_D_REG_25__SCAN_IN), .B2(keyinput223), .ZN(n8853) );
  AOI221_X1 U10365 ( .B1(P1_REG3_REG_14__SCAN_IN), .B2(keyinput207), .C1(
        keyinput223), .C2(P2_D_REG_25__SCAN_IN), .A(n8853), .ZN(n8860) );
  OAI22_X1 U10366 ( .A1(SI_6_), .A2(keyinput177), .B1(keyinput249), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8854) );
  AOI221_X1 U10367 ( .B1(SI_6_), .B2(keyinput177), .C1(P2_REG2_REG_27__SCAN_IN), .C2(keyinput249), .A(n8854), .ZN(n8859) );
  OAI22_X1 U10368 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(keyinput163), .B1(
        keyinput133), .B2(P2_D_REG_11__SCAN_IN), .ZN(n8855) );
  AOI221_X1 U10369 ( .B1(P1_DATAO_REG_10__SCAN_IN), .B2(keyinput163), .C1(
        P2_D_REG_11__SCAN_IN), .C2(keyinput133), .A(n8855), .ZN(n8858) );
  OAI22_X1 U10370 ( .A1(P1_REG1_REG_17__SCAN_IN), .A2(keyinput255), .B1(
        keyinput240), .B2(P2_REG1_REG_17__SCAN_IN), .ZN(n8856) );
  AOI221_X1 U10371 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(keyinput255), .C1(
        P2_REG1_REG_17__SCAN_IN), .C2(keyinput240), .A(n8856), .ZN(n8857) );
  NAND4_X1 U10372 ( .A1(n8860), .A2(n8859), .A3(n8858), .A4(n8857), .ZN(n8879)
         );
  OAI22_X1 U10373 ( .A1(SI_16_), .A2(keyinput170), .B1(keyinput201), .B2(
        P1_REG1_REG_19__SCAN_IN), .ZN(n8861) );
  AOI221_X1 U10374 ( .B1(SI_16_), .B2(keyinput170), .C1(
        P1_REG1_REG_19__SCAN_IN), .C2(keyinput201), .A(n8861), .ZN(n8868) );
  OAI22_X1 U10375 ( .A1(P2_REG2_REG_26__SCAN_IN), .A2(keyinput251), .B1(
        P1_ADDR_REG_6__SCAN_IN), .B2(keyinput213), .ZN(n8862) );
  AOI221_X1 U10376 ( .B1(P2_REG2_REG_26__SCAN_IN), .B2(keyinput251), .C1(
        keyinput213), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n8862), .ZN(n8867) );
  OAI22_X1 U10377 ( .A1(P1_REG0_REG_11__SCAN_IN), .A2(keyinput203), .B1(
        keyinput248), .B2(P2_REG1_REG_31__SCAN_IN), .ZN(n8863) );
  AOI221_X1 U10378 ( .B1(P1_REG0_REG_11__SCAN_IN), .B2(keyinput203), .C1(
        P2_REG1_REG_31__SCAN_IN), .C2(keyinput248), .A(n8863), .ZN(n8866) );
  OAI22_X1 U10379 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(keyinput214), .B1(SI_7_), .B2(keyinput182), .ZN(n8864) );
  AOI221_X1 U10380 ( .B1(P2_DATAO_REG_22__SCAN_IN), .B2(keyinput214), .C1(
        keyinput182), .C2(SI_7_), .A(n8864), .ZN(n8865) );
  NAND4_X1 U10381 ( .A1(n8868), .A2(n8867), .A3(n8866), .A4(n8865), .ZN(n8878)
         );
  OAI22_X1 U10382 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(keyinput204), .B1(
        P2_ADDR_REG_15__SCAN_IN), .B2(keyinput233), .ZN(n8869) );
  AOI221_X1 U10383 ( .B1(P2_IR_REG_9__SCAN_IN), .B2(keyinput204), .C1(
        keyinput233), .C2(P2_ADDR_REG_15__SCAN_IN), .A(n8869), .ZN(n8876) );
  OAI22_X1 U10384 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(keyinput211), .B1(
        P2_REG1_REG_14__SCAN_IN), .B2(keyinput141), .ZN(n8870) );
  AOI221_X1 U10385 ( .B1(P1_DATAO_REG_15__SCAN_IN), .B2(keyinput211), .C1(
        keyinput141), .C2(P2_REG1_REG_14__SCAN_IN), .A(n8870), .ZN(n8875) );
  OAI22_X1 U10386 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(keyinput134), .B1(SI_10_), 
        .B2(keyinput194), .ZN(n8871) );
  AOI221_X1 U10387 ( .B1(P1_IR_REG_18__SCAN_IN), .B2(keyinput134), .C1(
        keyinput194), .C2(SI_10_), .A(n8871), .ZN(n8874) );
  OAI22_X1 U10388 ( .A1(P1_D_REG_25__SCAN_IN), .A2(keyinput220), .B1(
        P1_REG2_REG_1__SCAN_IN), .B2(keyinput238), .ZN(n8872) );
  AOI221_X1 U10389 ( .B1(P1_D_REG_25__SCAN_IN), .B2(keyinput220), .C1(
        keyinput238), .C2(P1_REG2_REG_1__SCAN_IN), .A(n8872), .ZN(n8873) );
  NAND4_X1 U10390 ( .A1(n8876), .A2(n8875), .A3(n8874), .A4(n8873), .ZN(n8877)
         );
  NOR4_X1 U10391 ( .A1(n8880), .A2(n8879), .A3(n8878), .A4(n8877), .ZN(n8940)
         );
  INV_X1 U10392 ( .A(P1_B_REG_SCAN_IN), .ZN(n9471) );
  AOI22_X1 U10393 ( .A1(n9471), .A2(keyinput252), .B1(keyinput138), .B2(n6409), 
        .ZN(n8881) );
  OAI221_X1 U10394 ( .B1(n9471), .B2(keyinput252), .C1(n6409), .C2(keyinput138), .A(n8881), .ZN(n8890) );
  AOI22_X1 U10395 ( .A1(n9025), .A2(keyinput232), .B1(n8883), .B2(keyinput187), 
        .ZN(n8882) );
  OAI221_X1 U10396 ( .B1(n9025), .B2(keyinput232), .C1(n8883), .C2(keyinput187), .A(n8882), .ZN(n8889) );
  AOI22_X1 U10397 ( .A1(n5311), .A2(keyinput132), .B1(keyinput195), .B2(n5459), 
        .ZN(n8884) );
  OAI221_X1 U10398 ( .B1(n5311), .B2(keyinput132), .C1(n5459), .C2(keyinput195), .A(n8884), .ZN(n8888) );
  AOI22_X1 U10399 ( .A1(n8886), .A2(keyinput152), .B1(n5962), .B2(keyinput212), 
        .ZN(n8885) );
  OAI221_X1 U10400 ( .B1(n8886), .B2(keyinput152), .C1(n5962), .C2(keyinput212), .A(n8885), .ZN(n8887) );
  NOR4_X1 U10401 ( .A1(n8890), .A2(n8889), .A3(n8888), .A4(n8887), .ZN(n8939)
         );
  AOI22_X1 U10402 ( .A1(n8892), .A2(keyinput193), .B1(n7392), .B2(keyinput230), 
        .ZN(n8891) );
  OAI221_X1 U10403 ( .B1(n8892), .B2(keyinput193), .C1(n7392), .C2(keyinput230), .A(n8891), .ZN(n8900) );
  INV_X1 U10404 ( .A(P2_WR_REG_SCAN_IN), .ZN(n8967) );
  AOI22_X1 U10405 ( .A1(n8894), .A2(keyinput178), .B1(keyinput175), .B2(n8967), 
        .ZN(n8893) );
  OAI221_X1 U10406 ( .B1(n8894), .B2(keyinput178), .C1(n8967), .C2(keyinput175), .A(n8893), .ZN(n8899) );
  AOI22_X1 U10407 ( .A1(n9023), .A2(keyinput222), .B1(keyinput128), .B2(
        P2_U3151), .ZN(n8895) );
  OAI221_X1 U10408 ( .B1(n9023), .B2(keyinput222), .C1(P2_U3151), .C2(
        keyinput128), .A(n8895), .ZN(n8898) );
  INV_X1 U10409 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10438) );
  AOI22_X1 U10410 ( .A1(n10438), .A2(keyinput239), .B1(keyinput237), .B2(n9107), .ZN(n8896) );
  OAI221_X1 U10411 ( .B1(n10438), .B2(keyinput239), .C1(n9107), .C2(
        keyinput237), .A(n8896), .ZN(n8897) );
  NOR4_X1 U10412 ( .A1(n8900), .A2(n8899), .A3(n8898), .A4(n8897), .ZN(n8938)
         );
  AOI22_X1 U10413 ( .A1(n5267), .A2(keyinput216), .B1(keyinput199), .B2(n9044), 
        .ZN(n8901) );
  OAI221_X1 U10414 ( .B1(n5267), .B2(keyinput216), .C1(n9044), .C2(keyinput199), .A(n8901), .ZN(n8910) );
  INV_X1 U10415 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9883) );
  AOI22_X1 U10416 ( .A1(n9114), .A2(keyinput221), .B1(n9883), .B2(keyinput185), 
        .ZN(n8902) );
  OAI221_X1 U10417 ( .B1(n9114), .B2(keyinput221), .C1(n9883), .C2(keyinput185), .A(n8902), .ZN(n8909) );
  INV_X1 U10418 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n8904) );
  AOI22_X1 U10419 ( .A1(n8904), .A2(keyinput218), .B1(keyinput164), .B2(n9052), 
        .ZN(n8903) );
  OAI221_X1 U10420 ( .B1(n8904), .B2(keyinput218), .C1(n9052), .C2(keyinput164), .A(n8903), .ZN(n8908) );
  AOI22_X1 U10421 ( .A1(n8906), .A2(keyinput229), .B1(n9092), .B2(keyinput172), 
        .ZN(n8905) );
  OAI221_X1 U10422 ( .B1(n8906), .B2(keyinput229), .C1(n9092), .C2(keyinput172), .A(n8905), .ZN(n8907) );
  NOR4_X1 U10423 ( .A1(n8910), .A2(n8909), .A3(n8908), .A4(n8907), .ZN(n8936)
         );
  INV_X1 U10424 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10165) );
  AOI22_X1 U10425 ( .A1(n10078), .A2(keyinput156), .B1(keyinput206), .B2(
        n10165), .ZN(n8911) );
  OAI221_X1 U10426 ( .B1(n10078), .B2(keyinput156), .C1(n10165), .C2(
        keyinput206), .A(n8911), .ZN(n8919) );
  AOI22_X1 U10427 ( .A1(n8914), .A2(keyinput149), .B1(n8913), .B2(keyinput155), 
        .ZN(n8912) );
  OAI221_X1 U10428 ( .B1(n8914), .B2(keyinput149), .C1(n8913), .C2(keyinput155), .A(n8912), .ZN(n8918) );
  AOI22_X1 U10429 ( .A1(n8916), .A2(keyinput219), .B1(n9038), .B2(keyinput150), 
        .ZN(n8915) );
  OAI221_X1 U10430 ( .B1(n8916), .B2(keyinput219), .C1(n9038), .C2(keyinput150), .A(n8915), .ZN(n8917) );
  NOR3_X1 U10431 ( .A1(n8919), .A2(n8918), .A3(n8917), .ZN(n8935) );
  INV_X1 U10432 ( .A(SI_13_), .ZN(n9053) );
  AOI22_X1 U10433 ( .A1(n5469), .A2(keyinput225), .B1(keyinput130), .B2(n9053), 
        .ZN(n8920) );
  OAI221_X1 U10434 ( .B1(n5469), .B2(keyinput225), .C1(n9053), .C2(keyinput130), .A(n8920), .ZN(n8926) );
  XNOR2_X1 U10435 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(keyinput247), .ZN(n8924)
         );
  XNOR2_X1 U10436 ( .A(P2_REG1_REG_2__SCAN_IN), .B(keyinput235), .ZN(n8923) );
  XNOR2_X1 U10437 ( .A(keyinput153), .B(P2_IR_REG_24__SCAN_IN), .ZN(n8922) );
  XNOR2_X1 U10438 ( .A(keyinput250), .B(P1_ADDR_REG_9__SCAN_IN), .ZN(n8921) );
  NAND4_X1 U10439 ( .A1(n8924), .A2(n8923), .A3(n8922), .A4(n8921), .ZN(n8925)
         );
  NOR2_X1 U10440 ( .A1(n8926), .A2(n8925), .ZN(n8934) );
  AOI22_X1 U10441 ( .A1(n8928), .A2(keyinput173), .B1(n9050), .B2(keyinput208), 
        .ZN(n8927) );
  OAI221_X1 U10442 ( .B1(n8928), .B2(keyinput173), .C1(n9050), .C2(keyinput208), .A(n8927), .ZN(n8932) );
  AOI22_X1 U10443 ( .A1(n10451), .A2(keyinput198), .B1(n8930), .B2(keyinput147), .ZN(n8929) );
  OAI221_X1 U10444 ( .B1(n10451), .B2(keyinput198), .C1(n8930), .C2(
        keyinput147), .A(n8929), .ZN(n8931) );
  NOR2_X1 U10445 ( .A1(n8932), .A2(n8931), .ZN(n8933) );
  AND4_X1 U10446 ( .A1(n8936), .A2(n8935), .A3(n8934), .A4(n8933), .ZN(n8937)
         );
  AND4_X1 U10447 ( .A1(n8940), .A2(n8939), .A3(n8938), .A4(n8937), .ZN(n8941)
         );
  NAND3_X1 U10448 ( .A1(n8943), .A2(n8942), .A3(n8941), .ZN(n9132) );
  OAI22_X1 U10449 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(keyinput32), .B1(
        keyinput91), .B2(P2_REG0_REG_25__SCAN_IN), .ZN(n8944) );
  AOI221_X1 U10450 ( .B1(P1_DATAO_REG_26__SCAN_IN), .B2(keyinput32), .C1(
        P2_REG0_REG_25__SCAN_IN), .C2(keyinput91), .A(n8944), .ZN(n8951) );
  OAI22_X1 U10451 ( .A1(P1_REG2_REG_29__SCAN_IN), .A2(keyinput41), .B1(
        keyinput39), .B2(P2_ADDR_REG_8__SCAN_IN), .ZN(n8945) );
  AOI221_X1 U10452 ( .B1(P1_REG2_REG_29__SCAN_IN), .B2(keyinput41), .C1(
        P2_ADDR_REG_8__SCAN_IN), .C2(keyinput39), .A(n8945), .ZN(n8950) );
  OAI22_X1 U10453 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(keyinput33), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput56), .ZN(n8946) );
  AOI221_X1 U10454 ( .B1(P2_IR_REG_3__SCAN_IN), .B2(keyinput33), .C1(
        keyinput56), .C2(P2_REG3_REG_18__SCAN_IN), .A(n8946), .ZN(n8949) );
  OAI22_X1 U10455 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(keyinput4), .B1(
        P2_REG1_REG_25__SCAN_IN), .B2(keyinput24), .ZN(n8947) );
  AOI221_X1 U10456 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(keyinput4), .C1(
        keyinput24), .C2(P2_REG1_REG_25__SCAN_IN), .A(n8947), .ZN(n8948) );
  NAND4_X1 U10457 ( .A1(n8951), .A2(n8950), .A3(n8949), .A4(n8948), .ZN(n8983)
         );
  OAI22_X1 U10458 ( .A1(P1_REG0_REG_27__SCAN_IN), .A2(keyinput57), .B1(
        P1_REG0_REG_20__SCAN_IN), .B2(keyinput68), .ZN(n8952) );
  AOI221_X1 U10459 ( .B1(P1_REG0_REG_27__SCAN_IN), .B2(keyinput57), .C1(
        keyinput68), .C2(P1_REG0_REG_20__SCAN_IN), .A(n8952), .ZN(n8959) );
  OAI22_X1 U10460 ( .A1(P1_D_REG_4__SCAN_IN), .A2(keyinput9), .B1(keyinput74), 
        .B2(P1_REG1_REG_28__SCAN_IN), .ZN(n8953) );
  AOI221_X1 U10461 ( .B1(P1_D_REG_4__SCAN_IN), .B2(keyinput9), .C1(
        P1_REG1_REG_28__SCAN_IN), .C2(keyinput74), .A(n8953), .ZN(n8958) );
  OAI22_X1 U10462 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(keyinput52), .B1(
        keyinput53), .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8954) );
  AOI221_X1 U10463 ( .B1(P1_IR_REG_15__SCAN_IN), .B2(keyinput52), .C1(
        P2_DATAO_REG_16__SCAN_IN), .C2(keyinput53), .A(n8954), .ZN(n8957) );
  OAI22_X1 U10464 ( .A1(P1_REG1_REG_26__SCAN_IN), .A2(keyinput87), .B1(
        keyinput115), .B2(P2_REG1_REG_5__SCAN_IN), .ZN(n8955) );
  AOI221_X1 U10465 ( .B1(P1_REG1_REG_26__SCAN_IN), .B2(keyinput87), .C1(
        P2_REG1_REG_5__SCAN_IN), .C2(keyinput115), .A(n8955), .ZN(n8956) );
  NAND4_X1 U10466 ( .A1(n8959), .A2(n8958), .A3(n8957), .A4(n8956), .ZN(n8982)
         );
  OAI22_X1 U10467 ( .A1(n8961), .A2(keyinput95), .B1(keyinput123), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8960) );
  AOI221_X1 U10468 ( .B1(n8961), .B2(keyinput95), .C1(P2_REG2_REG_26__SCAN_IN), 
        .C2(keyinput123), .A(n8960), .ZN(n8971) );
  OAI22_X1 U10469 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(keyinput79), .B1(
        keyinput38), .B2(P2_REG0_REG_31__SCAN_IN), .ZN(n8962) );
  AOI221_X1 U10470 ( .B1(P1_REG3_REG_14__SCAN_IN), .B2(keyinput79), .C1(
        P2_REG0_REG_31__SCAN_IN), .C2(keyinput38), .A(n8962), .ZN(n8970) );
  OAI22_X1 U10471 ( .A1(n8965), .A2(keyinput12), .B1(n8964), .B2(keyinput112), 
        .ZN(n8963) );
  AOI221_X1 U10472 ( .B1(n8965), .B2(keyinput12), .C1(keyinput112), .C2(n8964), 
        .A(n8963), .ZN(n8969) );
  OAI22_X1 U10473 ( .A1(n6092), .A2(keyinput29), .B1(n8967), .B2(keyinput47), 
        .ZN(n8966) );
  AOI221_X1 U10474 ( .B1(n6092), .B2(keyinput29), .C1(keyinput47), .C2(n8967), 
        .A(n8966), .ZN(n8968) );
  NAND4_X1 U10475 ( .A1(n8971), .A2(n8970), .A3(n8969), .A4(n8968), .ZN(n8981)
         );
  OAI22_X1 U10476 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(keyinput35), .B1(
        keyinput98), .B2(P2_IR_REG_4__SCAN_IN), .ZN(n8972) );
  AOI221_X1 U10477 ( .B1(P1_DATAO_REG_10__SCAN_IN), .B2(keyinput35), .C1(
        P2_IR_REG_4__SCAN_IN), .C2(keyinput98), .A(n8972), .ZN(n8979) );
  OAI22_X1 U10478 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(keyinput108), .B1(
        P2_REG3_REG_4__SCAN_IN), .B2(keyinput65), .ZN(n8973) );
  AOI221_X1 U10479 ( .B1(P1_REG3_REG_9__SCAN_IN), .B2(keyinput108), .C1(
        keyinput65), .C2(P2_REG3_REG_4__SCAN_IN), .A(n8973), .ZN(n8978) );
  OAI22_X1 U10480 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput0), .B1(keyinput20), 
        .B2(P2_REG0_REG_17__SCAN_IN), .ZN(n8974) );
  AOI221_X1 U10481 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput0), .C1(
        P2_REG0_REG_17__SCAN_IN), .C2(keyinput20), .A(n8974), .ZN(n8977) );
  OAI22_X1 U10482 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(keyinput90), .B1(
        P1_REG0_REG_19__SCAN_IN), .B2(keyinput26), .ZN(n8975) );
  AOI221_X1 U10483 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(keyinput90), .C1(
        keyinput26), .C2(P1_REG0_REG_19__SCAN_IN), .A(n8975), .ZN(n8976) );
  NAND4_X1 U10484 ( .A1(n8979), .A2(n8978), .A3(n8977), .A4(n8976), .ZN(n8980)
         );
  NOR4_X1 U10485 ( .A1(n8983), .A2(n8982), .A3(n8981), .A4(n8980), .ZN(n9131)
         );
  OAI22_X1 U10486 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(keyinput55), .B1(
        P2_IR_REG_9__SCAN_IN), .B2(keyinput76), .ZN(n8984) );
  AOI221_X1 U10487 ( .B1(P1_REG1_REG_0__SCAN_IN), .B2(keyinput55), .C1(
        keyinput76), .C2(P2_IR_REG_9__SCAN_IN), .A(n8984), .ZN(n8991) );
  OAI22_X1 U10488 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(keyinput59), .B1(
        keyinput45), .B2(P2_REG0_REG_24__SCAN_IN), .ZN(n8985) );
  AOI221_X1 U10489 ( .B1(P1_DATAO_REG_19__SCAN_IN), .B2(keyinput59), .C1(
        P2_REG0_REG_24__SCAN_IN), .C2(keyinput45), .A(n8985), .ZN(n8990) );
  OAI22_X1 U10490 ( .A1(SI_6_), .A2(keyinput49), .B1(SI_2_), .B2(keyinput99), 
        .ZN(n8986) );
  AOI221_X1 U10491 ( .B1(SI_6_), .B2(keyinput49), .C1(keyinput99), .C2(SI_2_), 
        .A(n8986), .ZN(n8989) );
  OAI22_X1 U10492 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(keyinput43), .B1(
        P2_REG1_REG_7__SCAN_IN), .B2(keyinput111), .ZN(n8987) );
  AOI221_X1 U10493 ( .B1(P2_IR_REG_18__SCAN_IN), .B2(keyinput43), .C1(
        keyinput111), .C2(P2_REG1_REG_7__SCAN_IN), .A(n8987), .ZN(n8988) );
  NAND4_X1 U10494 ( .A1(n8991), .A2(n8990), .A3(n8989), .A4(n8988), .ZN(n9019)
         );
  OAI22_X1 U10495 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(keyinput64), .B1(
        P1_B_REG_SCAN_IN), .B2(keyinput124), .ZN(n8992) );
  AOI221_X1 U10496 ( .B1(P1_IR_REG_8__SCAN_IN), .B2(keyinput64), .C1(
        keyinput124), .C2(P1_B_REG_SCAN_IN), .A(n8992), .ZN(n8999) );
  OAI22_X1 U10497 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(keyinput27), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(keyinput113), .ZN(n8993) );
  AOI221_X1 U10498 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(keyinput27), .C1(
        keyinput113), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n8993), .ZN(n8998) );
  OAI22_X1 U10499 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(keyinput1), .B1(
        keyinput75), .B2(P1_REG0_REG_11__SCAN_IN), .ZN(n8994) );
  AOI221_X1 U10500 ( .B1(P2_DATAO_REG_6__SCAN_IN), .B2(keyinput1), .C1(
        P1_REG0_REG_11__SCAN_IN), .C2(keyinput75), .A(n8994), .ZN(n8997) );
  OAI22_X1 U10501 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(keyinput58), .B1(
        keyinput54), .B2(SI_7_), .ZN(n8995) );
  AOI221_X1 U10502 ( .B1(P1_IR_REG_12__SCAN_IN), .B2(keyinput58), .C1(SI_7_), 
        .C2(keyinput54), .A(n8995), .ZN(n8996) );
  NAND4_X1 U10503 ( .A1(n8999), .A2(n8998), .A3(n8997), .A4(n8996), .ZN(n9018)
         );
  OAI22_X1 U10504 ( .A1(P1_D_REG_14__SCAN_IN), .A2(keyinput116), .B1(
        keyinput14), .B2(P1_REG0_REG_10__SCAN_IN), .ZN(n9000) );
  AOI221_X1 U10505 ( .B1(P1_D_REG_14__SCAN_IN), .B2(keyinput116), .C1(
        P1_REG0_REG_10__SCAN_IN), .C2(keyinput14), .A(n9000), .ZN(n9007) );
  OAI22_X1 U10506 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(keyinput118), .B1(
        keyinput85), .B2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9001) );
  AOI221_X1 U10507 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(keyinput118), .C1(
        P1_ADDR_REG_6__SCAN_IN), .C2(keyinput85), .A(n9001), .ZN(n9006) );
  OAI22_X1 U10508 ( .A1(SI_10_), .A2(keyinput66), .B1(keyinput82), .B2(
        P1_REG3_REG_19__SCAN_IN), .ZN(n9002) );
  AOI221_X1 U10509 ( .B1(SI_10_), .B2(keyinput66), .C1(P1_REG3_REG_19__SCAN_IN), .C2(keyinput82), .A(n9002), .ZN(n9005) );
  OAI22_X1 U10510 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(keyinput50), .B1(
        keyinput19), .B2(P2_D_REG_4__SCAN_IN), .ZN(n9003) );
  AOI221_X1 U10511 ( .B1(P1_DATAO_REG_20__SCAN_IN), .B2(keyinput50), .C1(
        P2_D_REG_4__SCAN_IN), .C2(keyinput19), .A(n9003), .ZN(n9004) );
  NAND4_X1 U10512 ( .A1(n9007), .A2(n9006), .A3(n9005), .A4(n9004), .ZN(n9017)
         );
  OAI22_X1 U10513 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(keyinput67), .B1(
        keyinput77), .B2(P2_ADDR_REG_11__SCAN_IN), .ZN(n9008) );
  AOI221_X1 U10514 ( .B1(P1_IR_REG_25__SCAN_IN), .B2(keyinput67), .C1(
        P2_ADDR_REG_11__SCAN_IN), .C2(keyinput77), .A(n9008), .ZN(n9015) );
  OAI22_X1 U10515 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput21), .B1(
        keyinput18), .B2(P2_REG2_REG_28__SCAN_IN), .ZN(n9009) );
  AOI221_X1 U10516 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput21), .C1(
        P2_REG2_REG_28__SCAN_IN), .C2(keyinput18), .A(n9009), .ZN(n9014) );
  OAI22_X1 U10517 ( .A1(SI_9_), .A2(keyinput125), .B1(P2_REG1_REG_29__SCAN_IN), 
        .B2(keyinput101), .ZN(n9010) );
  AOI221_X1 U10518 ( .B1(SI_9_), .B2(keyinput125), .C1(keyinput101), .C2(
        P2_REG1_REG_29__SCAN_IN), .A(n9010), .ZN(n9013) );
  OAI22_X1 U10519 ( .A1(P1_D_REG_9__SCAN_IN), .A2(keyinput31), .B1(
        P1_REG2_REG_9__SCAN_IN), .B2(keyinput11), .ZN(n9011) );
  AOI221_X1 U10520 ( .B1(P1_D_REG_9__SCAN_IN), .B2(keyinput31), .C1(keyinput11), .C2(P1_REG2_REG_9__SCAN_IN), .A(n9011), .ZN(n9012) );
  NAND4_X1 U10521 ( .A1(n9015), .A2(n9014), .A3(n9013), .A4(n9012), .ZN(n9016)
         );
  NOR4_X1 U10522 ( .A1(n9019), .A2(n9018), .A3(n9017), .A4(n9016), .ZN(n9130)
         );
  AOI22_X1 U10523 ( .A1(n9021), .A2(keyinput23), .B1(n5469), .B2(keyinput97), 
        .ZN(n9020) );
  OAI221_X1 U10524 ( .B1(n9021), .B2(keyinput23), .C1(n5469), .C2(keyinput97), 
        .A(n9020), .ZN(n9033) );
  AOI22_X1 U10525 ( .A1(n7392), .A2(keyinput102), .B1(n9023), .B2(keyinput94), 
        .ZN(n9022) );
  OAI221_X1 U10526 ( .B1(n7392), .B2(keyinput102), .C1(n9023), .C2(keyinput94), 
        .A(n9022), .ZN(n9032) );
  AOI22_X1 U10527 ( .A1(n9026), .A2(keyinput72), .B1(n9025), .B2(keyinput104), 
        .ZN(n9024) );
  OAI221_X1 U10528 ( .B1(n9026), .B2(keyinput72), .C1(n9025), .C2(keyinput104), 
        .A(n9024), .ZN(n9031) );
  INV_X1 U10529 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n9029) );
  AOI22_X1 U10530 ( .A1(n9029), .A2(keyinput105), .B1(keyinput81), .B2(n9028), 
        .ZN(n9027) );
  OAI221_X1 U10531 ( .B1(n9029), .B2(keyinput105), .C1(n9028), .C2(keyinput81), 
        .A(n9027), .ZN(n9030) );
  NOR4_X1 U10532 ( .A1(n9033), .A2(n9032), .A3(n9031), .A4(n9030), .ZN(n9089)
         );
  AOI22_X1 U10533 ( .A1(n6276), .A2(keyinput7), .B1(keyinput69), .B2(n9035), 
        .ZN(n9034) );
  OAI221_X1 U10534 ( .B1(n6276), .B2(keyinput7), .C1(n9035), .C2(keyinput69), 
        .A(n9034), .ZN(n9048) );
  AOI22_X1 U10535 ( .A1(n9038), .A2(keyinput22), .B1(keyinput40), .B2(n9037), 
        .ZN(n9036) );
  OAI221_X1 U10536 ( .B1(n9038), .B2(keyinput22), .C1(n9037), .C2(keyinput40), 
        .A(n9036), .ZN(n9047) );
  AOI22_X1 U10537 ( .A1(n9041), .A2(keyinput86), .B1(keyinput120), .B2(n9040), 
        .ZN(n9039) );
  OAI221_X1 U10538 ( .B1(n9041), .B2(keyinput86), .C1(n9040), .C2(keyinput120), 
        .A(n9039), .ZN(n9046) );
  AOI22_X1 U10539 ( .A1(n9044), .A2(keyinput71), .B1(n9043), .B2(keyinput15), 
        .ZN(n9042) );
  OAI221_X1 U10540 ( .B1(n9044), .B2(keyinput71), .C1(n9043), .C2(keyinput15), 
        .A(n9042), .ZN(n9045) );
  NOR4_X1 U10541 ( .A1(n9048), .A2(n9047), .A3(n9046), .A4(n9045), .ZN(n9088)
         );
  AOI22_X1 U10542 ( .A1(n5842), .A2(keyinput37), .B1(keyinput80), .B2(n9050), 
        .ZN(n9049) );
  OAI221_X1 U10543 ( .B1(n5842), .B2(keyinput37), .C1(n9050), .C2(keyinput80), 
        .A(n9049), .ZN(n9060) );
  AOI22_X1 U10544 ( .A1(n9053), .A2(keyinput2), .B1(keyinput36), .B2(n9052), 
        .ZN(n9051) );
  OAI221_X1 U10545 ( .B1(n9053), .B2(keyinput2), .C1(n9052), .C2(keyinput36), 
        .A(n9051), .ZN(n9059) );
  XNOR2_X1 U10546 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput61), .ZN(n9057) );
  XNOR2_X1 U10547 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput126), .ZN(n9056) );
  XNOR2_X1 U10548 ( .A(P2_REG1_REG_2__SCAN_IN), .B(keyinput107), .ZN(n9055) );
  XNOR2_X1 U10549 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput114), .ZN(n9054) );
  NAND4_X1 U10550 ( .A1(n9057), .A2(n9056), .A3(n9055), .A4(n9054), .ZN(n9058)
         );
  NOR3_X1 U10551 ( .A1(n9060), .A2(n9059), .A3(n9058), .ZN(n9086) );
  AOI22_X1 U10552 ( .A1(n9062), .A2(keyinput34), .B1(keyinput25), .B2(n5798), 
        .ZN(n9061) );
  OAI221_X1 U10553 ( .B1(n9062), .B2(keyinput34), .C1(n5798), .C2(keyinput25), 
        .A(n9061), .ZN(n9070) );
  INV_X1 U10554 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9907) );
  AOI22_X1 U10555 ( .A1(n9064), .A2(keyinput42), .B1(keyinput16), .B2(n9907), 
        .ZN(n9063) );
  OAI221_X1 U10556 ( .B1(n9064), .B2(keyinput42), .C1(n9907), .C2(keyinput16), 
        .A(n9063), .ZN(n9069) );
  AOI22_X1 U10557 ( .A1(n9067), .A2(keyinput106), .B1(n9066), .B2(keyinput17), 
        .ZN(n9065) );
  OAI221_X1 U10558 ( .B1(n9067), .B2(keyinput106), .C1(n9066), .C2(keyinput17), 
        .A(n9065), .ZN(n9068) );
  NOR3_X1 U10559 ( .A1(n9070), .A2(n9069), .A3(n9068), .ZN(n9085) );
  AOI22_X1 U10560 ( .A1(n6393), .A2(keyinput110), .B1(n10176), .B2(keyinput117), .ZN(n9071) );
  OAI221_X1 U10561 ( .B1(n6393), .B2(keyinput110), .C1(n10176), .C2(
        keyinput117), .A(n9071), .ZN(n9077) );
  XNOR2_X1 U10562 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(keyinput119), .ZN(n9075)
         );
  XNOR2_X1 U10563 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(keyinput3), .ZN(n9074) );
  XNOR2_X1 U10564 ( .A(keyinput103), .B(P1_REG2_REG_14__SCAN_IN), .ZN(n9073)
         );
  XNOR2_X1 U10565 ( .A(keyinput6), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9072) );
  NAND4_X1 U10566 ( .A1(n9075), .A2(n9074), .A3(n9073), .A4(n9072), .ZN(n9076)
         );
  NOR2_X1 U10567 ( .A1(n9077), .A2(n9076), .ZN(n9084) );
  AOI22_X1 U10568 ( .A1(n5962), .A2(keyinput84), .B1(keyinput48), .B2(n7901), 
        .ZN(n9078) );
  OAI221_X1 U10569 ( .B1(n5962), .B2(keyinput84), .C1(n7901), .C2(keyinput48), 
        .A(n9078), .ZN(n9082) );
  AOI22_X1 U10570 ( .A1(n10165), .A2(keyinput78), .B1(keyinput96), .B2(n9080), 
        .ZN(n9079) );
  OAI221_X1 U10571 ( .B1(n10165), .B2(keyinput78), .C1(n9080), .C2(keyinput96), 
        .A(n9079), .ZN(n9081) );
  NOR2_X1 U10572 ( .A1(n9082), .A2(n9081), .ZN(n9083) );
  AND4_X1 U10573 ( .A1(n9086), .A2(n9085), .A3(n9084), .A4(n9083), .ZN(n9087)
         );
  AND3_X1 U10574 ( .A1(n9089), .A2(n9088), .A3(n9087), .ZN(n9128) );
  INV_X1 U10575 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9975) );
  AOI22_X1 U10576 ( .A1(n9975), .A2(keyinput127), .B1(keyinput63), .B2(n6051), 
        .ZN(n9090) );
  OAI221_X1 U10577 ( .B1(n9975), .B2(keyinput127), .C1(n6051), .C2(keyinput63), 
        .A(n9090), .ZN(n9100) );
  INV_X1 U10578 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9859) );
  AOI22_X1 U10579 ( .A1(n9859), .A2(keyinput73), .B1(n9092), .B2(keyinput44), 
        .ZN(n9091) );
  OAI221_X1 U10580 ( .B1(n9859), .B2(keyinput73), .C1(n9092), .C2(keyinput44), 
        .A(n9091), .ZN(n9099) );
  INV_X1 U10581 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n9095) );
  AOI22_X1 U10582 ( .A1(n9095), .A2(keyinput121), .B1(n9094), .B2(keyinput5), 
        .ZN(n9093) );
  OAI221_X1 U10583 ( .B1(n9095), .B2(keyinput121), .C1(n9094), .C2(keyinput5), 
        .A(n9093), .ZN(n9098) );
  AOI22_X1 U10584 ( .A1(n5310), .A2(keyinput46), .B1(keyinput70), .B2(n10451), 
        .ZN(n9096) );
  OAI221_X1 U10585 ( .B1(n5310), .B2(keyinput46), .C1(n10451), .C2(keyinput70), 
        .A(n9096), .ZN(n9097) );
  NOR4_X1 U10586 ( .A1(n9100), .A2(n9099), .A3(n9098), .A4(n9097), .ZN(n9127)
         );
  AOI22_X1 U10587 ( .A1(n5786), .A2(keyinput60), .B1(n6409), .B2(keyinput10), 
        .ZN(n9101) );
  OAI221_X1 U10588 ( .B1(n5786), .B2(keyinput60), .C1(n6409), .C2(keyinput10), 
        .A(n9101), .ZN(n9111) );
  AOI22_X1 U10589 ( .A1(n5267), .A2(keyinput88), .B1(keyinput83), .B2(n9103), 
        .ZN(n9102) );
  OAI221_X1 U10590 ( .B1(n5267), .B2(keyinput88), .C1(n9103), .C2(keyinput83), 
        .A(n9102), .ZN(n9110) );
  INV_X1 U10591 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9591) );
  INV_X1 U10592 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9105) );
  AOI22_X1 U10593 ( .A1(n9591), .A2(keyinput62), .B1(keyinput89), .B2(n9105), 
        .ZN(n9104) );
  OAI221_X1 U10594 ( .B1(n9591), .B2(keyinput62), .C1(n9105), .C2(keyinput89), 
        .A(n9104), .ZN(n9109) );
  AOI22_X1 U10595 ( .A1(n9107), .A2(keyinput109), .B1(n5779), .B2(keyinput100), 
        .ZN(n9106) );
  OAI221_X1 U10596 ( .B1(n9107), .B2(keyinput109), .C1(n5779), .C2(keyinput100), .A(n9106), .ZN(n9108) );
  NOR4_X1 U10597 ( .A1(n9111), .A2(n9110), .A3(n9109), .A4(n9108), .ZN(n9126)
         );
  AOI22_X1 U10598 ( .A1(n10078), .A2(keyinput28), .B1(keyinput92), .B2(n10077), 
        .ZN(n9112) );
  OAI221_X1 U10599 ( .B1(n10078), .B2(keyinput28), .C1(n10077), .C2(keyinput92), .A(n9112), .ZN(n9124) );
  AOI22_X1 U10600 ( .A1(n9115), .A2(keyinput51), .B1(n9114), .B2(keyinput93), 
        .ZN(n9113) );
  OAI221_X1 U10601 ( .B1(n9115), .B2(keyinput51), .C1(n9114), .C2(keyinput93), 
        .A(n9113), .ZN(n9123) );
  INV_X1 U10602 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9117) );
  AOI22_X1 U10603 ( .A1(n9118), .A2(keyinput8), .B1(keyinput122), .B2(n9117), 
        .ZN(n9116) );
  OAI221_X1 U10604 ( .B1(n9118), .B2(keyinput8), .C1(n9117), .C2(keyinput122), 
        .A(n9116), .ZN(n9122) );
  AOI22_X1 U10605 ( .A1(n9120), .A2(keyinput13), .B1(n5108), .B2(keyinput30), 
        .ZN(n9119) );
  OAI221_X1 U10606 ( .B1(n9120), .B2(keyinput13), .C1(n5108), .C2(keyinput30), 
        .A(n9119), .ZN(n9121) );
  NOR4_X1 U10607 ( .A1(n9124), .A2(n9123), .A3(n9122), .A4(n9121), .ZN(n9125)
         );
  AND4_X1 U10608 ( .A1(n9128), .A2(n9127), .A3(n9126), .A4(n9125), .ZN(n9129)
         );
  NAND4_X1 U10609 ( .A1(n9132), .A2(n9131), .A3(n9130), .A4(n9129), .ZN(n9133)
         );
  XNOR2_X1 U10610 ( .A(n9134), .B(n9133), .ZN(P1_U3226) );
  NAND2_X1 U10611 ( .A1(n9136), .A2(n9135), .ZN(n9138) );
  OAI21_X1 U10612 ( .B1(n9139), .B2(n9138), .A(n9137), .ZN(n9140) );
  NAND2_X1 U10613 ( .A1(n9140), .A2(n9966), .ZN(n9147) );
  OR2_X1 U10614 ( .A1(n9142), .A2(n9141), .ZN(n9144) );
  NAND2_X1 U10615 ( .A1(n9500), .A2(n9184), .ZN(n9143) );
  AND2_X1 U10616 ( .A1(n9144), .A2(n9143), .ZN(n9773) );
  NAND2_X1 U10617 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9564) );
  OAI21_X1 U10618 ( .B1(n9214), .B2(n9773), .A(n9564), .ZN(n9145) );
  AOI21_X1 U10619 ( .B1(n9779), .B2(n9211), .A(n9145), .ZN(n9146) );
  OAI211_X1 U10620 ( .C1(n5011), .C2(n9963), .A(n9147), .B(n9146), .ZN(
        P1_U3228) );
  INV_X1 U10621 ( .A(n9148), .ZN(n9150) );
  NOR3_X1 U10622 ( .A1(n9151), .A2(n9150), .A3(n9149), .ZN(n9154) );
  INV_X1 U10623 ( .A(n9152), .ZN(n9153) );
  OAI21_X1 U10624 ( .B1(n9154), .B2(n9153), .A(n9966), .ZN(n9158) );
  INV_X1 U10625 ( .A(n9171), .ZN(n9495) );
  AOI22_X1 U10626 ( .A1(n9495), .A2(n9197), .B1(n9184), .B2(n9493), .ZN(n9666)
         );
  OAI22_X1 U10627 ( .A1(n9666), .A2(n9214), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9155), .ZN(n9156) );
  AOI21_X1 U10628 ( .B1(n9672), .B2(n9211), .A(n9156), .ZN(n9157) );
  OAI211_X1 U10629 ( .C1(n9897), .C2(n9963), .A(n9158), .B(n9157), .ZN(
        P1_U3229) );
  OAI21_X1 U10630 ( .B1(n9161), .B2(n9160), .A(n9159), .ZN(n9162) );
  NAND2_X1 U10631 ( .A1(n9162), .A2(n9966), .ZN(n9168) );
  NAND2_X1 U10632 ( .A1(n9499), .A2(n9197), .ZN(n9164) );
  NAND2_X1 U10633 ( .A1(n9497), .A2(n9184), .ZN(n9163) );
  AND2_X1 U10634 ( .A1(n9164), .A2(n9163), .ZN(n9730) );
  INV_X1 U10635 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9165) );
  OAI22_X1 U10636 ( .A1(n9214), .A2(n9730), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9165), .ZN(n9166) );
  AOI21_X1 U10637 ( .B1(n9735), .B2(n9211), .A(n9166), .ZN(n9167) );
  OAI211_X1 U10638 ( .C1(n9913), .C2(n9963), .A(n9168), .B(n9167), .ZN(
        P1_U3233) );
  AOI21_X1 U10639 ( .B1(n9170), .B2(n8690), .A(n9169), .ZN(n9178) );
  INV_X1 U10640 ( .A(n9704), .ZN(n9175) );
  OR2_X1 U10641 ( .A1(n9171), .A2(n9195), .ZN(n9173) );
  NAND2_X1 U10642 ( .A1(n9497), .A2(n9197), .ZN(n9172) );
  NAND2_X1 U10643 ( .A1(n9173), .A2(n9172), .ZN(n9699) );
  AOI22_X1 U10644 ( .A1(n9960), .A2(n9699), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9174) );
  OAI21_X1 U10645 ( .B1(n9970), .B2(n9175), .A(n9174), .ZN(n9176) );
  AOI21_X1 U10646 ( .B1(n9703), .B2(n9217), .A(n9176), .ZN(n9177) );
  OAI21_X1 U10647 ( .B1(n9178), .B2(n9220), .A(n9177), .ZN(P1_U3235) );
  INV_X1 U10648 ( .A(n9179), .ZN(n9181) );
  NAND2_X1 U10649 ( .A1(n9181), .A2(n9180), .ZN(n9182) );
  XNOR2_X1 U10650 ( .A(n9183), .B(n9182), .ZN(n9191) );
  NAND2_X1 U10651 ( .A1(n9499), .A2(n9184), .ZN(n9186) );
  NAND2_X1 U10652 ( .A1(n9501), .A2(n9197), .ZN(n9185) );
  NAND2_X1 U10653 ( .A1(n9186), .A2(n9185), .ZN(n9761) );
  AOI22_X1 U10654 ( .A1(n9960), .A2(n9761), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3086), .ZN(n9187) );
  OAI21_X1 U10655 ( .B1(n9970), .B2(n9188), .A(n9187), .ZN(n9189) );
  AOI21_X1 U10656 ( .B1(n9765), .B2(n9217), .A(n9189), .ZN(n9190) );
  OAI21_X1 U10657 ( .B1(n9191), .B2(n9220), .A(n9190), .ZN(P1_U3238) );
  NAND2_X1 U10658 ( .A1(n9192), .A2(n9966), .ZN(n9205) );
  AOI21_X1 U10659 ( .B1(n8760), .B2(n9194), .A(n9193), .ZN(n9204) );
  INV_X1 U10660 ( .A(n9640), .ZN(n9201) );
  OR2_X1 U10661 ( .A1(n9196), .A2(n9195), .ZN(n9199) );
  NAND2_X1 U10662 ( .A1(n9493), .A2(n9197), .ZN(n9198) );
  NAND2_X1 U10663 ( .A1(n9199), .A2(n9198), .ZN(n9636) );
  AOI22_X1 U10664 ( .A1(n9960), .A2(n9636), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9200) );
  OAI21_X1 U10665 ( .B1(n9970), .B2(n9201), .A(n9200), .ZN(n9202) );
  AOI21_X1 U10666 ( .B1(n9639), .B2(n9217), .A(n9202), .ZN(n9203) );
  OAI21_X1 U10667 ( .B1(n9205), .B2(n9204), .A(n9203), .ZN(P1_U3240) );
  INV_X1 U10668 ( .A(n9206), .ZN(n9207) );
  AOI21_X1 U10669 ( .B1(n9209), .B2(n9208), .A(n9207), .ZN(n9221) );
  NAND2_X1 U10670 ( .A1(n9211), .A2(n9210), .ZN(n9213) );
  OAI211_X1 U10671 ( .C1(n9215), .C2(n9214), .A(n9213), .B(n9212), .ZN(n9216)
         );
  AOI21_X1 U10672 ( .B1(n9218), .B2(n9217), .A(n9216), .ZN(n9219) );
  OAI21_X1 U10673 ( .B1(n9221), .B2(n9220), .A(n9219), .ZN(P1_U3241) );
  INV_X1 U10674 ( .A(n9222), .ZN(n9616) );
  NAND2_X1 U10675 ( .A1(n9318), .A2(n9310), .ZN(n9439) );
  NAND4_X1 U10676 ( .A1(n10034), .A2(n9394), .A3(n9393), .A4(n9325), .ZN(n9231) );
  NAND2_X1 U10677 ( .A1(n9223), .A2(n9397), .ZN(n9225) );
  INV_X1 U10678 ( .A(n9225), .ZN(n9224) );
  NAND3_X1 U10679 ( .A1(n7289), .A2(n9321), .A3(n9224), .ZN(n9230) );
  NOR3_X1 U10680 ( .A1(n9225), .A2(n9394), .A3(n9325), .ZN(n9228) );
  NAND3_X1 U10681 ( .A1(n9225), .A2(n10034), .A3(n9325), .ZN(n9226) );
  OAI21_X1 U10682 ( .B1(n9325), .B2(n10034), .A(n9226), .ZN(n9227) );
  NOR3_X1 U10683 ( .A1(n9228), .A2(n9227), .A3(n10033), .ZN(n9229) );
  OAI211_X1 U10684 ( .C1(n9232), .C2(n9231), .A(n9230), .B(n9229), .ZN(n9242)
         );
  INV_X1 U10685 ( .A(n9233), .ZN(n9234) );
  MUX2_X1 U10686 ( .A(n9235), .B(n9234), .S(n9325), .Z(n9241) );
  NAND2_X1 U10687 ( .A1(n9236), .A2(n9243), .ZN(n9239) );
  INV_X1 U10688 ( .A(n9237), .ZN(n9238) );
  MUX2_X1 U10689 ( .A(n9239), .B(n9238), .S(n9325), .Z(n9240) );
  INV_X1 U10690 ( .A(n9243), .ZN(n9244) );
  OAI21_X1 U10691 ( .B1(n9248), .B2(n9244), .A(n9399), .ZN(n9245) );
  NAND4_X1 U10692 ( .A1(n9245), .A2(n9402), .A3(n9325), .A4(n9401), .ZN(n9251)
         );
  INV_X1 U10693 ( .A(n9246), .ZN(n9247) );
  OAI21_X1 U10694 ( .B1(n9248), .B2(n9247), .A(n9402), .ZN(n9249) );
  NAND4_X1 U10695 ( .A1(n9249), .A2(n9321), .A3(n9399), .A4(n9254), .ZN(n9250)
         );
  NAND2_X1 U10696 ( .A1(n9251), .A2(n9250), .ZN(n9256) );
  NAND2_X1 U10697 ( .A1(n9257), .A2(n9401), .ZN(n9252) );
  OAI211_X1 U10698 ( .C1(n9256), .C2(n9252), .A(n9409), .B(n9255), .ZN(n9253)
         );
  NAND2_X1 U10699 ( .A1(n9255), .A2(n9254), .ZN(n9405) );
  NOR2_X1 U10700 ( .A1(n9256), .A2(n9405), .ZN(n9259) );
  NAND2_X1 U10701 ( .A1(n9258), .A2(n9257), .ZN(n9406) );
  NAND2_X1 U10702 ( .A1(n9261), .A2(n9349), .ZN(n9269) );
  OR2_X1 U10703 ( .A1(n9263), .A2(n9262), .ZN(n9264) );
  AND2_X1 U10704 ( .A1(n9787), .A2(n9264), .ZN(n9410) );
  MUX2_X1 U10705 ( .A(n9414), .B(n9410), .S(n9325), .Z(n9268) );
  INV_X1 U10706 ( .A(n9787), .ZN(n9415) );
  INV_X1 U10707 ( .A(n9265), .ZN(n9266) );
  MUX2_X1 U10708 ( .A(n9415), .B(n9266), .S(n9325), .Z(n9267) );
  AOI211_X1 U10709 ( .C1(n9269), .C2(n9268), .A(n9267), .B(n9788), .ZN(n9273)
         );
  NAND2_X1 U10710 ( .A1(n9276), .A2(n9418), .ZN(n9271) );
  INV_X1 U10711 ( .A(n9416), .ZN(n9270) );
  MUX2_X1 U10712 ( .A(n9271), .B(n9270), .S(n9325), .Z(n9272) );
  INV_X1 U10713 ( .A(n9421), .ZN(n9274) );
  INV_X1 U10714 ( .A(n9275), .ZN(n9280) );
  NAND2_X1 U10715 ( .A1(n9330), .A2(n9276), .ZN(n9420) );
  AOI21_X1 U10716 ( .B1(n9277), .B2(n9756), .A(n9420), .ZN(n9278) );
  NAND2_X1 U10717 ( .A1(n9284), .A2(n9331), .ZN(n9424) );
  NOR2_X1 U10718 ( .A1(n9278), .A2(n9424), .ZN(n9279) );
  MUX2_X1 U10719 ( .A(n9280), .B(n9279), .S(n9325), .Z(n9291) );
  INV_X1 U10720 ( .A(n9288), .ZN(n9281) );
  OAI22_X1 U10721 ( .A1(n5650), .A2(n9748), .B1(n9281), .B2(n9325), .ZN(n9285)
         );
  NOR2_X1 U10722 ( .A1(n9282), .A2(n9321), .ZN(n9283) );
  AOI22_X1 U10723 ( .A1(n9285), .A2(n9284), .B1(n9283), .B2(n9286), .ZN(n9290)
         );
  AND2_X1 U10724 ( .A1(n9292), .A2(n9286), .ZN(n9432) );
  OR2_X1 U10725 ( .A1(n9715), .A2(n9287), .ZN(n9428) );
  AND2_X1 U10726 ( .A1(n9428), .A2(n9288), .ZN(n9378) );
  MUX2_X1 U10727 ( .A(n9432), .B(n9378), .S(n9325), .Z(n9289) );
  OAI21_X1 U10728 ( .B1(n9291), .B2(n9290), .A(n9289), .ZN(n9294) );
  MUX2_X1 U10729 ( .A(n9428), .B(n9292), .S(n9325), .Z(n9293) );
  AOI21_X1 U10730 ( .B1(n9294), .B2(n9293), .A(n4723), .ZN(n9300) );
  NAND2_X1 U10731 ( .A1(n9297), .A2(n9295), .ZN(n9373) );
  NAND2_X1 U10732 ( .A1(n9372), .A2(n9296), .ZN(n9429) );
  MUX2_X1 U10733 ( .A(n9373), .B(n9429), .S(n9325), .Z(n9299) );
  MUX2_X1 U10734 ( .A(n9372), .B(n9297), .S(n9325), .Z(n9298) );
  OAI211_X1 U10735 ( .C1(n9300), .C2(n9299), .A(n5752), .B(n9298), .ZN(n9302)
         );
  MUX2_X1 U10736 ( .A(n9647), .B(n9431), .S(n9325), .Z(n9301) );
  NAND2_X1 U10737 ( .A1(n9302), .A2(n9301), .ZN(n9308) );
  INV_X1 U10738 ( .A(n9377), .ZN(n9303) );
  INV_X1 U10739 ( .A(n9368), .ZN(n9305) );
  NOR2_X1 U10740 ( .A1(n9306), .A2(n9305), .ZN(n9316) );
  INV_X1 U10741 ( .A(n9307), .ZN(n9434) );
  AOI211_X1 U10742 ( .C1(n9308), .C2(n9377), .A(n9616), .B(n9434), .ZN(n9312)
         );
  INV_X1 U10743 ( .A(n9309), .ZN(n9311) );
  OAI21_X1 U10744 ( .B1(n9312), .B2(n9311), .A(n9310), .ZN(n9314) );
  NAND3_X1 U10745 ( .A1(n9314), .A2(n9368), .A3(n9313), .ZN(n9315) );
  MUX2_X1 U10746 ( .A(n9316), .B(n9315), .S(n9325), .Z(n9317) );
  OAI21_X1 U10747 ( .B1(n9321), .B2(n9318), .A(n9317), .ZN(n9320) );
  MUX2_X1 U10748 ( .A(n9367), .B(n9369), .S(n9325), .Z(n9319) );
  OAI21_X1 U10749 ( .B1(n9320), .B2(n9359), .A(n9319), .ZN(n9324) );
  OR2_X1 U10750 ( .A1(n9327), .A2(n9452), .ZN(n9460) );
  INV_X1 U10751 ( .A(n9371), .ZN(n9489) );
  NAND2_X1 U10752 ( .A1(n9489), .A2(n9322), .ZN(n9459) );
  NAND3_X1 U10753 ( .A1(n9323), .A2(n9460), .A3(n9459), .ZN(n9329) );
  NAND3_X1 U10754 ( .A1(n9326), .A2(n9489), .A3(n9327), .ZN(n9328) );
  NAND2_X1 U10755 ( .A1(n9327), .A2(n9452), .ZN(n9462) );
  NAND3_X1 U10756 ( .A1(n9329), .A2(n9328), .A3(n9462), .ZN(n9363) );
  AOI21_X1 U10757 ( .B1(n9363), .B2(n9365), .A(n9381), .ZN(n9488) );
  XNOR2_X1 U10758 ( .A(n9458), .B(n9371), .ZN(n9361) );
  INV_X1 U10759 ( .A(n9648), .ZN(n9357) );
  NAND2_X1 U10760 ( .A1(n9331), .A2(n9330), .ZN(n9758) );
  XNOR2_X1 U10761 ( .A(n9333), .B(n9332), .ZN(n9777) );
  NOR2_X1 U10762 ( .A1(n9334), .A2(n7262), .ZN(n9340) );
  NOR2_X1 U10763 ( .A1(n9335), .A2(n10062), .ZN(n9339) );
  NOR2_X1 U10764 ( .A1(n9336), .A2(n5726), .ZN(n9338) );
  NAND4_X1 U10765 ( .A1(n9340), .A2(n9339), .A3(n9338), .A4(n9337), .ZN(n9343)
         );
  NOR3_X1 U10766 ( .A1(n9343), .A2(n9342), .A3(n9341), .ZN(n9346) );
  INV_X1 U10767 ( .A(n9396), .ZN(n9344) );
  NAND4_X1 U10768 ( .A1(n9346), .A2(n9345), .A3(n9344), .A4(n5741), .ZN(n9348)
         );
  NOR2_X1 U10769 ( .A1(n9348), .A2(n9347), .ZN(n9351) );
  NAND4_X1 U10770 ( .A1(n9786), .A2(n9351), .A3(n9350), .A4(n9349), .ZN(n9352)
         );
  NOR3_X1 U10771 ( .A1(n9758), .A2(n9777), .A3(n9352), .ZN(n9353) );
  AND3_X1 U10772 ( .A1(n9728), .A2(n9743), .A3(n9353), .ZN(n9354) );
  NAND4_X1 U10773 ( .A1(n9687), .A2(n9697), .A3(n9354), .A4(n9712), .ZN(n9355)
         );
  NOR2_X1 U10774 ( .A1(n9663), .A2(n9355), .ZN(n9356) );
  NAND4_X1 U10775 ( .A1(n9624), .A2(n9357), .A3(n9633), .A4(n9356), .ZN(n9358)
         );
  NOR4_X1 U10776 ( .A1(n9361), .A2(n9360), .A3(n9359), .A4(n9358), .ZN(n9362)
         );
  NAND3_X1 U10777 ( .A1(n9460), .A2(n9362), .A3(n9462), .ZN(n9465) );
  INV_X1 U10778 ( .A(n9470), .ZN(n9472) );
  NAND4_X1 U10779 ( .A1(n9465), .A2(n9467), .A3(n9598), .A4(n9472), .ZN(n9487)
         );
  NAND2_X1 U10780 ( .A1(n9363), .A2(n5091), .ZN(n9485) );
  NOR2_X1 U10781 ( .A1(n9460), .A2(n9720), .ZN(n9366) );
  NOR4_X1 U10782 ( .A1(n9366), .A2(n9365), .A3(n9364), .A4(n9470), .ZN(n9484)
         );
  NAND2_X1 U10783 ( .A1(n9369), .A2(n9368), .ZN(n9455) );
  INV_X1 U10784 ( .A(n9455), .ZN(n9370) );
  OR2_X1 U10785 ( .A1(n9441), .A2(n9370), .ZN(n9444) );
  OR2_X1 U10786 ( .A1(n9458), .A2(n9371), .ZN(n9443) );
  NAND2_X1 U10787 ( .A1(n9373), .A2(n9372), .ZN(n9374) );
  NAND2_X1 U10788 ( .A1(n9647), .A2(n9374), .ZN(n9375) );
  NAND2_X1 U10789 ( .A1(n9375), .A2(n9431), .ZN(n9376) );
  AND2_X1 U10790 ( .A1(n9377), .A2(n9376), .ZN(n9436) );
  INV_X1 U10791 ( .A(n9436), .ZN(n9380) );
  INV_X1 U10792 ( .A(n9378), .ZN(n9379) );
  NOR2_X1 U10793 ( .A1(n9380), .A2(n9379), .ZN(n9447) );
  AOI21_X1 U10794 ( .B1(n6633), .B2(n10104), .A(n9381), .ZN(n9384) );
  INV_X1 U10795 ( .A(n9382), .ZN(n9383) );
  AND2_X1 U10796 ( .A1(n9384), .A2(n9383), .ZN(n9387) );
  OAI211_X1 U10797 ( .C1(n9388), .C2(n9387), .A(n9386), .B(n9385), .ZN(n9390)
         );
  NAND2_X1 U10798 ( .A1(n9390), .A2(n9389), .ZN(n9392) );
  NAND2_X1 U10799 ( .A1(n9392), .A2(n9391), .ZN(n9395) );
  NAND3_X1 U10800 ( .A1(n9395), .A2(n9394), .A3(n9393), .ZN(n9398) );
  AOI21_X1 U10801 ( .B1(n9398), .B2(n9397), .A(n9396), .ZN(n9404) );
  NAND2_X1 U10802 ( .A1(n9400), .A2(n9399), .ZN(n9403) );
  OAI211_X1 U10803 ( .C1(n9404), .C2(n9403), .A(n9402), .B(n9401), .ZN(n9408)
         );
  INV_X1 U10804 ( .A(n9405), .ZN(n9407) );
  AOI21_X1 U10805 ( .B1(n9408), .B2(n9407), .A(n9406), .ZN(n9412) );
  INV_X1 U10806 ( .A(n9410), .ZN(n9411) );
  OR3_X1 U10807 ( .A1(n9412), .A2(n5745), .A3(n9411), .ZN(n9413) );
  OAI21_X1 U10808 ( .B1(n9415), .B2(n9414), .A(n9413), .ZN(n9417) );
  NAND2_X1 U10809 ( .A1(n9417), .A2(n9416), .ZN(n9419) );
  NAND2_X1 U10810 ( .A1(n9419), .A2(n9418), .ZN(n9422) );
  AOI21_X1 U10811 ( .B1(n9422), .B2(n9421), .A(n9420), .ZN(n9425) );
  OAI21_X1 U10812 ( .B1(n9425), .B2(n9424), .A(n9423), .ZN(n9426) );
  AOI21_X1 U10813 ( .B1(n9447), .B2(n9426), .A(n9616), .ZN(n9427) );
  NOR2_X1 U10814 ( .A1(n9427), .A2(n9448), .ZN(n9440) );
  INV_X1 U10815 ( .A(n9428), .ZN(n9433) );
  INV_X1 U10816 ( .A(n9429), .ZN(n9430) );
  OAI211_X1 U10817 ( .C1(n9433), .C2(n9432), .A(n9431), .B(n9430), .ZN(n9435)
         );
  AOI21_X1 U10818 ( .B1(n9436), .B2(n9435), .A(n9434), .ZN(n9437) );
  NOR2_X1 U10819 ( .A1(n9448), .A2(n9437), .ZN(n9438) );
  OR2_X1 U10820 ( .A1(n9439), .A2(n9438), .ZN(n9451) );
  OR3_X1 U10821 ( .A1(n9441), .A2(n9440), .A3(n9451), .ZN(n9442) );
  NAND4_X1 U10822 ( .A1(n9462), .A2(n9444), .A3(n9443), .A4(n9442), .ZN(n9445)
         );
  NAND2_X1 U10823 ( .A1(n9445), .A2(n9460), .ZN(n9482) );
  OR3_X1 U10824 ( .A1(n9470), .A2(n9467), .A3(n9720), .ZN(n9481) );
  AOI21_X1 U10825 ( .B1(n9447), .B2(n9446), .A(n9616), .ZN(n9449) );
  NOR2_X1 U10826 ( .A1(n9449), .A2(n9448), .ZN(n9450) );
  NOR2_X1 U10827 ( .A1(n9451), .A2(n9450), .ZN(n9456) );
  NAND2_X1 U10828 ( .A1(n9458), .A2(n9452), .ZN(n9453) );
  OAI211_X1 U10829 ( .C1(n9456), .C2(n9455), .A(n9454), .B(n9453), .ZN(n9457)
         );
  OAI21_X1 U10830 ( .B1(n9459), .B2(n9458), .A(n9457), .ZN(n9461) );
  NAND2_X1 U10831 ( .A1(n9461), .A2(n9460), .ZN(n9464) );
  NAND3_X1 U10832 ( .A1(n9464), .A2(n9463), .A3(n9462), .ZN(n9466) );
  NAND2_X1 U10833 ( .A1(n9466), .A2(n9465), .ZN(n9468) );
  NAND4_X1 U10834 ( .A1(n9468), .A2(n9467), .A3(n9472), .A4(n9720), .ZN(n9480)
         );
  NOR2_X1 U10835 ( .A1(n9470), .A2(n9469), .ZN(n9478) );
  AOI21_X1 U10836 ( .B1(n9472), .B2(n5455), .A(n9471), .ZN(n9477) );
  INV_X1 U10837 ( .A(n9473), .ZN(n9474) );
  NAND4_X1 U10838 ( .A1(n9475), .A2(n10005), .A3(n9987), .A4(n9474), .ZN(n9476) );
  AOI22_X1 U10839 ( .A1(n9482), .A2(n9478), .B1(n9477), .B2(n9476), .ZN(n9479)
         );
  OAI211_X1 U10840 ( .C1(n9482), .C2(n9481), .A(n9480), .B(n9479), .ZN(n9483)
         );
  AOI21_X1 U10841 ( .B1(n9485), .B2(n9484), .A(n9483), .ZN(n9486) );
  OAI21_X1 U10842 ( .B1(n9488), .B2(n9487), .A(n9486), .ZN(P1_U3242) );
  MUX2_X1 U10843 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9489), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10844 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9490), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10845 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9491), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10846 ( .A(n9492), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9504), .Z(
        P1_U3580) );
  MUX2_X1 U10847 ( .A(n9493), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9504), .Z(
        P1_U3579) );
  MUX2_X1 U10848 ( .A(n9494), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9504), .Z(
        P1_U3578) );
  MUX2_X1 U10849 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9495), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10850 ( .A(n9496), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9504), .Z(
        P1_U3576) );
  MUX2_X1 U10851 ( .A(n9497), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9504), .Z(
        P1_U3575) );
  MUX2_X1 U10852 ( .A(n9498), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9504), .Z(
        P1_U3574) );
  MUX2_X1 U10853 ( .A(n9499), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9504), .Z(
        P1_U3573) );
  MUX2_X1 U10854 ( .A(n9500), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9504), .Z(
        P1_U3572) );
  MUX2_X1 U10855 ( .A(n9501), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9504), .Z(
        P1_U3571) );
  MUX2_X1 U10856 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9502), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10857 ( .A(n9503), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9504), .Z(
        P1_U3569) );
  MUX2_X1 U10858 ( .A(n9505), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9504), .Z(
        P1_U3568) );
  MUX2_X1 U10859 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9506), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10860 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9507), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10861 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9508), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10862 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9509), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10863 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9510), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10864 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9511), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10865 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9512), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10866 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9513), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10867 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9514), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10868 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9515), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10869 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9516), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10870 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9517), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10871 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6633), .S(P1_U3973), .Z(
        P1_U3555) );
  AOI211_X1 U10872 ( .C1(n9520), .C2(n9519), .A(n9518), .B(n10018), .ZN(n9521)
         );
  INV_X1 U10873 ( .A(n9521), .ZN(n9531) );
  INV_X1 U10874 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9523) );
  NAND2_X1 U10875 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9522) );
  OAI21_X1 U10876 ( .B1(n9601), .B2(n9523), .A(n9522), .ZN(n9524) );
  AOI21_X1 U10877 ( .B1(n9525), .B2(n10025), .A(n9524), .ZN(n9530) );
  OAI211_X1 U10878 ( .C1(n9528), .C2(n9527), .A(n10017), .B(n9526), .ZN(n9529)
         );
  NAND3_X1 U10879 ( .A1(n9531), .A2(n9530), .A3(n9529), .ZN(P1_U3246) );
  NOR2_X1 U10880 ( .A1(n9532), .A2(n9542), .ZN(n9534) );
  NAND2_X1 U10881 ( .A1(n9561), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9535) );
  OAI21_X1 U10882 ( .B1(n9561), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9535), .ZN(
        n9536) );
  INV_X1 U10883 ( .A(n9536), .ZN(n9537) );
  OAI21_X1 U10884 ( .B1(n9538), .B2(n9537), .A(n9560), .ZN(n9551) );
  INV_X1 U10885 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9541) );
  NAND2_X1 U10886 ( .A1(n10025), .A2(n9561), .ZN(n9540) );
  NAND2_X1 U10887 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n9539) );
  OAI211_X1 U10888 ( .C1(n9541), .C2(n9601), .A(n9540), .B(n9539), .ZN(n9550)
         );
  NOR2_X1 U10889 ( .A1(n9543), .A2(n9542), .ZN(n9545) );
  XNOR2_X1 U10890 ( .A(n9561), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n9547) );
  INV_X1 U10891 ( .A(n9555), .ZN(n9546) );
  AOI211_X1 U10892 ( .C1(n9548), .C2(n9547), .A(n10018), .B(n9546), .ZN(n9549)
         );
  AOI211_X1 U10893 ( .C1(n10017), .C2(n9551), .A(n9550), .B(n9549), .ZN(n9552)
         );
  INV_X1 U10894 ( .A(n9552), .ZN(P1_U3259) );
  INV_X1 U10895 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9553) );
  XNOR2_X1 U10896 ( .A(n9578), .B(n9553), .ZN(n9557) );
  NAND2_X1 U10897 ( .A1(n9561), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9554) );
  OAI21_X1 U10898 ( .B1(n9557), .B2(n9556), .A(n9580), .ZN(n9558) );
  NAND2_X1 U10899 ( .A1(n9558), .A2(n9593), .ZN(n9570) );
  NOR2_X1 U10900 ( .A1(n9578), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9559) );
  AOI21_X1 U10901 ( .B1(n9578), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9559), .ZN(
        n9563) );
  OAI21_X1 U10902 ( .B1(n9563), .B2(n9562), .A(n9573), .ZN(n9568) );
  INV_X1 U10903 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9566) );
  NAND2_X1 U10904 ( .A1(n10025), .A2(n9578), .ZN(n9565) );
  OAI211_X1 U10905 ( .C1(n9566), .C2(n9601), .A(n9565), .B(n9564), .ZN(n9567)
         );
  AOI21_X1 U10906 ( .B1(n9568), .B2(n10017), .A(n9567), .ZN(n9569) );
  NAND2_X1 U10907 ( .A1(n9570), .A2(n9569), .ZN(P1_U3260) );
  NAND2_X1 U10908 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n9571) );
  OAI21_X1 U10909 ( .B1(n9601), .B2(n10453), .A(n9571), .ZN(n9577) );
  INV_X1 U10910 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9864) );
  NOR2_X1 U10911 ( .A1(n9587), .A2(n9864), .ZN(n9572) );
  AOI21_X1 U10912 ( .B1(n9864), .B2(n9587), .A(n9572), .ZN(n9575) );
  OAI21_X1 U10913 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n9578), .A(n9573), .ZN(
        n9574) );
  NOR2_X1 U10914 ( .A1(n9574), .A2(n9575), .ZN(n9586) );
  AOI211_X1 U10915 ( .C1(n9575), .C2(n9574), .A(n9993), .B(n9586), .ZN(n9576)
         );
  AOI211_X1 U10916 ( .C1(n10025), .C2(n9587), .A(n9577), .B(n9576), .ZN(n9585)
         );
  OR2_X1 U10917 ( .A1(n9578), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9579) );
  AND2_X1 U10918 ( .A1(n9580), .A2(n9579), .ZN(n9583) );
  NAND2_X1 U10919 ( .A1(n9587), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9589) );
  OR2_X1 U10920 ( .A1(n9587), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9581) );
  AND2_X1 U10921 ( .A1(n9589), .A2(n9581), .ZN(n9582) );
  NAND2_X1 U10922 ( .A1(n9583), .A2(n9582), .ZN(n9590) );
  OAI211_X1 U10923 ( .C1(n9583), .C2(n9582), .A(n9590), .B(n9593), .ZN(n9584)
         );
  NAND2_X1 U10924 ( .A1(n9585), .A2(n9584), .ZN(P1_U3261) );
  AOI21_X1 U10925 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n9587), .A(n9586), .ZN(
        n9588) );
  XNOR2_X1 U10926 ( .A(n9588), .B(n9859), .ZN(n9597) );
  INV_X1 U10927 ( .A(n9597), .ZN(n9594) );
  NAND2_X1 U10928 ( .A1(n9590), .A2(n9589), .ZN(n9592) );
  XNOR2_X1 U10929 ( .A(n9592), .B(n9591), .ZN(n9596) );
  AOI22_X1 U10930 ( .A1(n9594), .A2(n10017), .B1(n9593), .B2(n9596), .ZN(n9599) );
  NAND2_X1 U10931 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9600) );
  NAND2_X1 U10932 ( .A1(n9602), .A2(n10066), .ZN(n9605) );
  INV_X1 U10933 ( .A(n9603), .ZN(n9805) );
  NOR2_X1 U10934 ( .A1(n9805), .A2(n10070), .ZN(n9609) );
  AOI21_X1 U10935 ( .B1(n10043), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9609), .ZN(
        n9604) );
  OAI211_X1 U10936 ( .C1(n5018), .C2(n9800), .A(n9605), .B(n9604), .ZN(
        P1_U3263) );
  OAI211_X1 U10937 ( .C1(n9607), .C2(n9880), .A(n10063), .B(n9606), .ZN(n9806)
         );
  NOR2_X1 U10938 ( .A1(n9880), .A2(n9800), .ZN(n9608) );
  AOI211_X1 U10939 ( .C1(n10043), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9609), .B(
        n9608), .ZN(n9610) );
  OAI21_X1 U10940 ( .B1(n9611), .B2(n9806), .A(n9610), .ZN(P1_U3264) );
  INV_X1 U10941 ( .A(n9612), .ZN(n9614) );
  INV_X1 U10942 ( .A(n5765), .ZN(n9613) );
  AOI211_X1 U10943 ( .C1(n9628), .C2(n9614), .A(n9794), .B(n9613), .ZN(n9818)
         );
  INV_X1 U10944 ( .A(n9615), .ZN(n9619) );
  OAI21_X1 U10945 ( .B1(n9624), .B2(n9616), .A(n9615), .ZN(n9617) );
  OAI211_X1 U10946 ( .C1(n9619), .C2(n9618), .A(n10054), .B(n9617), .ZN(n9622)
         );
  INV_X1 U10947 ( .A(n9620), .ZN(n9621) );
  NAND2_X1 U10948 ( .A1(n9622), .A2(n9621), .ZN(n9817) );
  AOI21_X1 U10949 ( .B1(n9818), .B2(n9720), .A(n9817), .ZN(n9631) );
  XNOR2_X1 U10950 ( .A(n9623), .B(n9624), .ZN(n9819) );
  NAND2_X1 U10951 ( .A1(n9819), .A2(n10067), .ZN(n9630) );
  INV_X1 U10952 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9626) );
  OAI22_X1 U10953 ( .A1(n10058), .A2(n9626), .B1(n9625), .B2(n10056), .ZN(
        n9627) );
  AOI21_X1 U10954 ( .B1(n9628), .B2(n10060), .A(n9627), .ZN(n9629) );
  OAI211_X1 U10955 ( .C1(n10043), .C2(n9631), .A(n9630), .B(n9629), .ZN(
        P1_U3266) );
  XOR2_X1 U10956 ( .A(n9633), .B(n9632), .Z(n9824) );
  INV_X1 U10957 ( .A(n9824), .ZN(n9645) );
  XNOR2_X1 U10958 ( .A(n9634), .B(n9633), .ZN(n9635) );
  NAND2_X1 U10959 ( .A1(n9635), .A2(n10054), .ZN(n9638) );
  INV_X1 U10960 ( .A(n9636), .ZN(n9637) );
  NAND2_X1 U10961 ( .A1(n9638), .A2(n9637), .ZN(n9822) );
  AOI211_X1 U10962 ( .C1(n9639), .C2(n5027), .A(n9794), .B(n9612), .ZN(n9823)
         );
  NAND2_X1 U10963 ( .A1(n9823), .A2(n10066), .ZN(n9642) );
  AOI22_X1 U10964 ( .A1(n10043), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9640), 
        .B2(n10042), .ZN(n9641) );
  OAI211_X1 U10965 ( .C1(n9889), .C2(n9800), .A(n9642), .B(n9641), .ZN(n9643)
         );
  AOI21_X1 U10966 ( .B1(n9822), .B2(n10058), .A(n9643), .ZN(n9644) );
  OAI21_X1 U10967 ( .B1(n9645), .B2(n9803), .A(n9644), .ZN(P1_U3267) );
  XOR2_X1 U10968 ( .A(n9646), .B(n9648), .Z(n9829) );
  INV_X1 U10969 ( .A(n9829), .ZN(n9662) );
  NAND2_X1 U10970 ( .A1(n9665), .A2(n9647), .ZN(n9649) );
  NAND2_X1 U10971 ( .A1(n9649), .A2(n9648), .ZN(n9651) );
  NAND2_X1 U10972 ( .A1(n9651), .A2(n9650), .ZN(n9652) );
  NAND2_X1 U10973 ( .A1(n9652), .A2(n10054), .ZN(n9654) );
  NAND2_X1 U10974 ( .A1(n9654), .A2(n9653), .ZN(n9827) );
  AOI211_X1 U10975 ( .C1(n9656), .C2(n9669), .A(n9794), .B(n9655), .ZN(n9828)
         );
  NAND2_X1 U10976 ( .A1(n9828), .A2(n10066), .ZN(n9659) );
  AOI22_X1 U10977 ( .A1(n10043), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9657), 
        .B2(n10042), .ZN(n9658) );
  OAI211_X1 U10978 ( .C1(n9893), .C2(n9800), .A(n9659), .B(n9658), .ZN(n9660)
         );
  AOI21_X1 U10979 ( .B1(n10058), .B2(n9827), .A(n9660), .ZN(n9661) );
  OAI21_X1 U10980 ( .B1(n9662), .B2(n9803), .A(n9661), .ZN(P1_U3268) );
  XNOR2_X1 U10981 ( .A(n9664), .B(n9663), .ZN(n9834) );
  INV_X1 U10982 ( .A(n9834), .ZN(n9677) );
  OAI211_X1 U10983 ( .C1(n4522), .C2(n5752), .A(n10054), .B(n9665), .ZN(n9667)
         );
  NAND2_X1 U10984 ( .A1(n9667), .A2(n9666), .ZN(n9832) );
  INV_X1 U10985 ( .A(n9669), .ZN(n9670) );
  AOI211_X1 U10986 ( .C1(n9671), .C2(n9668), .A(n9794), .B(n9670), .ZN(n9833)
         );
  NAND2_X1 U10987 ( .A1(n9833), .A2(n10066), .ZN(n9674) );
  AOI22_X1 U10988 ( .A1(n10043), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9672), 
        .B2(n10042), .ZN(n9673) );
  OAI211_X1 U10989 ( .C1(n9897), .C2(n9800), .A(n9674), .B(n9673), .ZN(n9675)
         );
  AOI21_X1 U10990 ( .B1(n10058), .B2(n9832), .A(n9675), .ZN(n9676) );
  OAI21_X1 U10991 ( .B1(n9677), .B2(n9803), .A(n9676), .ZN(P1_U3269) );
  INV_X1 U10992 ( .A(n9678), .ZN(n9680) );
  INV_X1 U10993 ( .A(n9668), .ZN(n9679) );
  AOI211_X1 U10994 ( .C1(n9690), .C2(n9680), .A(n9794), .B(n9679), .ZN(n9838)
         );
  INV_X1 U10995 ( .A(n9681), .ZN(n9682) );
  NOR2_X1 U10996 ( .A1(n10056), .A2(n9682), .ZN(n9686) );
  XOR2_X1 U10997 ( .A(n9687), .B(n9683), .Z(n9685) );
  OAI21_X1 U10998 ( .B1(n9685), .B2(n10036), .A(n9684), .ZN(n9837) );
  AOI211_X1 U10999 ( .C1(n9838), .C2(n9720), .A(n9686), .B(n9837), .ZN(n9693)
         );
  OAI21_X1 U11000 ( .B1(n9689), .B2(n5677), .A(n9688), .ZN(n9839) );
  NAND2_X1 U11001 ( .A1(n9839), .A2(n10067), .ZN(n9692) );
  AOI22_X1 U11002 ( .A1(n9690), .A2(n10060), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n10043), .ZN(n9691) );
  OAI211_X1 U11003 ( .C1(n9693), .C2(n10070), .A(n9692), .B(n9691), .ZN(
        P1_U3270) );
  XNOR2_X1 U11004 ( .A(n9694), .B(n4723), .ZN(n9844) );
  INV_X1 U11005 ( .A(n9844), .ZN(n9709) );
  OAI21_X1 U11006 ( .B1(n9697), .B2(n9696), .A(n9695), .ZN(n9698) );
  NAND2_X1 U11007 ( .A1(n9698), .A2(n10054), .ZN(n9701) );
  INV_X1 U11008 ( .A(n9699), .ZN(n9700) );
  NAND2_X1 U11009 ( .A1(n9701), .A2(n9700), .ZN(n9842) );
  INV_X1 U11010 ( .A(n9702), .ZN(n9716) );
  AOI211_X1 U11011 ( .C1(n9703), .C2(n9716), .A(n9794), .B(n9678), .ZN(n9843)
         );
  NAND2_X1 U11012 ( .A1(n9843), .A2(n10066), .ZN(n9706) );
  AOI22_X1 U11013 ( .A1(n10043), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9704), 
        .B2(n10042), .ZN(n9705) );
  OAI211_X1 U11014 ( .C1(n9905), .C2(n9800), .A(n9706), .B(n9705), .ZN(n9707)
         );
  AOI21_X1 U11015 ( .B1(n10058), .B2(n9842), .A(n9707), .ZN(n9708) );
  OAI21_X1 U11016 ( .B1(n9709), .B2(n9803), .A(n9708), .ZN(P1_U3271) );
  XOR2_X1 U11017 ( .A(n9710), .B(n9712), .Z(n9848) );
  XOR2_X1 U11018 ( .A(n9712), .B(n9711), .Z(n9714) );
  OAI21_X1 U11019 ( .B1(n9714), .B2(n10036), .A(n9713), .ZN(n9719) );
  AOI21_X1 U11020 ( .B1(n4519), .B2(n9715), .A(n9794), .ZN(n9717) );
  AOI21_X1 U11021 ( .B1(n9717), .B2(n9716), .A(n9719), .ZN(n9718) );
  INV_X1 U11022 ( .A(n9718), .ZN(n9847) );
  OAI211_X1 U11023 ( .C1(n9720), .C2(n9719), .A(n9847), .B(n10058), .ZN(n9723)
         );
  AOI22_X1 U11024 ( .A1(n10070), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9721), 
        .B2(n10042), .ZN(n9722) );
  OAI211_X1 U11025 ( .C1(n9909), .C2(n9800), .A(n9723), .B(n9722), .ZN(n9724)
         );
  AOI21_X1 U11026 ( .B1(n10067), .B2(n9848), .A(n9724), .ZN(n9725) );
  INV_X1 U11027 ( .A(n9725), .ZN(P1_U3272) );
  OAI21_X1 U11028 ( .B1(n9727), .B2(n5650), .A(n9726), .ZN(n9853) );
  INV_X1 U11029 ( .A(n9853), .ZN(n9740) );
  XNOR2_X1 U11030 ( .A(n9446), .B(n9728), .ZN(n9729) );
  NAND2_X1 U11031 ( .A1(n9729), .A2(n10054), .ZN(n9731) );
  NAND2_X1 U11032 ( .A1(n9731), .A2(n9730), .ZN(n9851) );
  INV_X1 U11033 ( .A(n4519), .ZN(n9733) );
  AOI211_X1 U11034 ( .C1(n9734), .C2(n9732), .A(n9794), .B(n9733), .ZN(n9852)
         );
  NAND2_X1 U11035 ( .A1(n9852), .A2(n10066), .ZN(n9737) );
  AOI22_X1 U11036 ( .A1(n10043), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9735), 
        .B2(n10042), .ZN(n9736) );
  OAI211_X1 U11037 ( .C1(n9913), .C2(n9800), .A(n9737), .B(n9736), .ZN(n9738)
         );
  AOI21_X1 U11038 ( .B1(n10058), .B2(n9851), .A(n9738), .ZN(n9739) );
  OAI21_X1 U11039 ( .B1(n9740), .B2(n9803), .A(n9739), .ZN(P1_U3273) );
  XNOR2_X1 U11040 ( .A(n9741), .B(n9743), .ZN(n9858) );
  INV_X1 U11041 ( .A(n9858), .ZN(n9754) );
  XOR2_X1 U11042 ( .A(n9742), .B(n9743), .Z(n9746) );
  INV_X1 U11043 ( .A(n9744), .ZN(n9745) );
  OAI21_X1 U11044 ( .B1(n9746), .B2(n10036), .A(n9745), .ZN(n9856) );
  INV_X1 U11045 ( .A(n9732), .ZN(n9747) );
  AOI211_X1 U11046 ( .C1(n9748), .C2(n5010), .A(n9794), .B(n9747), .ZN(n9857)
         );
  NAND2_X1 U11047 ( .A1(n9857), .A2(n10066), .ZN(n9751) );
  AOI22_X1 U11048 ( .A1(n10043), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9749), 
        .B2(n10042), .ZN(n9750) );
  OAI211_X1 U11049 ( .C1(n9917), .C2(n9800), .A(n9751), .B(n9750), .ZN(n9752)
         );
  AOI21_X1 U11050 ( .B1(n10058), .B2(n9856), .A(n9752), .ZN(n9753) );
  OAI21_X1 U11051 ( .B1(n9754), .B2(n9803), .A(n9753), .ZN(P1_U3274) );
  XNOR2_X1 U11052 ( .A(n9755), .B(n9758), .ZN(n9863) );
  INV_X1 U11053 ( .A(n9863), .ZN(n9771) );
  NAND2_X1 U11054 ( .A1(n9757), .A2(n9756), .ZN(n9759) );
  XNOR2_X1 U11055 ( .A(n9759), .B(n9758), .ZN(n9760) );
  NAND2_X1 U11056 ( .A1(n9760), .A2(n10054), .ZN(n9763) );
  INV_X1 U11057 ( .A(n9761), .ZN(n9762) );
  NAND2_X1 U11058 ( .A1(n9763), .A2(n9762), .ZN(n9861) );
  INV_X1 U11059 ( .A(n9765), .ZN(n9921) );
  AOI211_X1 U11060 ( .C1(n9765), .C2(n9778), .A(n9794), .B(n9764), .ZN(n9862)
         );
  NAND2_X1 U11061 ( .A1(n9862), .A2(n10066), .ZN(n9768) );
  AOI22_X1 U11062 ( .A1(n10043), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9766), 
        .B2(n10042), .ZN(n9767) );
  OAI211_X1 U11063 ( .C1(n9921), .C2(n9800), .A(n9768), .B(n9767), .ZN(n9769)
         );
  AOI21_X1 U11064 ( .B1(n10058), .B2(n9861), .A(n9769), .ZN(n9770) );
  OAI21_X1 U11065 ( .B1(n9771), .B2(n9803), .A(n9770), .ZN(P1_U3275) );
  XNOR2_X1 U11066 ( .A(n9772), .B(n9777), .ZN(n9775) );
  INV_X1 U11067 ( .A(n9773), .ZN(n9774) );
  AOI21_X1 U11068 ( .B1(n9775), .B2(n10054), .A(n9774), .ZN(n9972) );
  XOR2_X1 U11069 ( .A(n9777), .B(n9776), .Z(n9974) );
  NAND2_X1 U11070 ( .A1(n9974), .A2(n10067), .ZN(n9784) );
  OAI211_X1 U11071 ( .C1(n5295), .C2(n5011), .A(n10063), .B(n9778), .ZN(n9971)
         );
  INV_X1 U11072 ( .A(n9971), .ZN(n9782) );
  AOI22_X1 U11073 ( .A1(n10070), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9779), 
        .B2(n10042), .ZN(n9780) );
  OAI21_X1 U11074 ( .B1(n5011), .B2(n9800), .A(n9780), .ZN(n9781) );
  AOI21_X1 U11075 ( .B1(n9782), .B2(n10066), .A(n9781), .ZN(n9783) );
  OAI211_X1 U11076 ( .C1(n10070), .C2(n9972), .A(n9784), .B(n9783), .ZN(
        P1_U3276) );
  XNOR2_X1 U11077 ( .A(n9785), .B(n9786), .ZN(n9868) );
  INV_X1 U11078 ( .A(n9868), .ZN(n9804) );
  NAND3_X1 U11079 ( .A1(n9789), .A2(n9788), .A3(n9787), .ZN(n9790) );
  NAND3_X1 U11080 ( .A1(n9791), .A2(n10054), .A3(n9790), .ZN(n9793) );
  NAND2_X1 U11081 ( .A1(n9793), .A2(n9792), .ZN(n9866) );
  AOI211_X1 U11082 ( .C1(n9796), .C2(n9795), .A(n9794), .B(n5295), .ZN(n9867)
         );
  NAND2_X1 U11083 ( .A1(n9867), .A2(n10066), .ZN(n9799) );
  AOI22_X1 U11084 ( .A1(n10043), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9797), 
        .B2(n10042), .ZN(n9798) );
  OAI211_X1 U11085 ( .C1(n9925), .C2(n9800), .A(n9799), .B(n9798), .ZN(n9801)
         );
  AOI21_X1 U11086 ( .B1(n10058), .B2(n9866), .A(n9801), .ZN(n9802) );
  OAI21_X1 U11087 ( .B1(n9804), .B2(n9803), .A(n9802), .ZN(P1_U3277) );
  INV_X1 U11088 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9807) );
  AND2_X1 U11089 ( .A1(n9806), .A2(n9805), .ZN(n9877) );
  MUX2_X1 U11090 ( .A(n9807), .B(n9877), .S(n10192), .Z(n9808) );
  OAI21_X1 U11091 ( .B1(n9880), .B2(n9875), .A(n9808), .ZN(P1_U3552) );
  INV_X1 U11092 ( .A(n9809), .ZN(n9811) );
  OAI21_X1 U11093 ( .B1(n9816), .B2(n9815), .A(n9814), .ZN(n9881) );
  MUX2_X1 U11094 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9881), .S(n10192), .Z(
        P1_U3551) );
  INV_X1 U11095 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9820) );
  AOI211_X1 U11096 ( .C1(n9819), .C2(n10172), .A(n9818), .B(n9817), .ZN(n9882)
         );
  MUX2_X1 U11097 ( .A(n9820), .B(n9882), .S(n10192), .Z(n9821) );
  OAI21_X1 U11098 ( .B1(n9885), .B2(n9875), .A(n9821), .ZN(P1_U3549) );
  INV_X1 U11099 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9825) );
  AOI211_X1 U11100 ( .C1(n9824), .C2(n10172), .A(n9823), .B(n9822), .ZN(n9886)
         );
  MUX2_X1 U11101 ( .A(n9825), .B(n9886), .S(n10192), .Z(n9826) );
  OAI21_X1 U11102 ( .B1(n9889), .B2(n9875), .A(n9826), .ZN(P1_U3548) );
  INV_X1 U11103 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9830) );
  AOI211_X1 U11104 ( .C1(n9829), .C2(n10172), .A(n9828), .B(n9827), .ZN(n9890)
         );
  MUX2_X1 U11105 ( .A(n9830), .B(n9890), .S(n10192), .Z(n9831) );
  OAI21_X1 U11106 ( .B1(n9893), .B2(n9875), .A(n9831), .ZN(P1_U3547) );
  INV_X1 U11107 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9835) );
  AOI211_X1 U11108 ( .C1(n9834), .C2(n10172), .A(n9833), .B(n9832), .ZN(n9894)
         );
  MUX2_X1 U11109 ( .A(n9835), .B(n9894), .S(n10192), .Z(n9836) );
  OAI21_X1 U11110 ( .B1(n9897), .B2(n9875), .A(n9836), .ZN(P1_U3546) );
  INV_X1 U11111 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9840) );
  AOI211_X1 U11112 ( .C1(n9839), .C2(n10172), .A(n9838), .B(n9837), .ZN(n9898)
         );
  MUX2_X1 U11113 ( .A(n9840), .B(n9898), .S(n10192), .Z(n9841) );
  OAI21_X1 U11114 ( .B1(n9901), .B2(n9875), .A(n9841), .ZN(P1_U3545) );
  INV_X1 U11115 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9845) );
  AOI211_X1 U11116 ( .C1(n9844), .C2(n10172), .A(n9843), .B(n9842), .ZN(n9902)
         );
  MUX2_X1 U11117 ( .A(n9845), .B(n9902), .S(n10192), .Z(n9846) );
  OAI21_X1 U11118 ( .B1(n9905), .B2(n9875), .A(n9846), .ZN(P1_U3544) );
  INV_X1 U11119 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9849) );
  AOI21_X1 U11120 ( .B1(n9848), .B2(n10172), .A(n9847), .ZN(n9906) );
  MUX2_X1 U11121 ( .A(n9849), .B(n9906), .S(n10192), .Z(n9850) );
  OAI21_X1 U11122 ( .B1(n9909), .B2(n9875), .A(n9850), .ZN(P1_U3543) );
  INV_X1 U11123 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9854) );
  AOI211_X1 U11124 ( .C1(n9853), .C2(n10172), .A(n9852), .B(n9851), .ZN(n9910)
         );
  MUX2_X1 U11125 ( .A(n9854), .B(n9910), .S(n10192), .Z(n9855) );
  OAI21_X1 U11126 ( .B1(n9913), .B2(n9875), .A(n9855), .ZN(P1_U3542) );
  AOI211_X1 U11127 ( .C1(n9858), .C2(n10172), .A(n9857), .B(n9856), .ZN(n9914)
         );
  MUX2_X1 U11128 ( .A(n9859), .B(n9914), .S(n10192), .Z(n9860) );
  OAI21_X1 U11129 ( .B1(n9917), .B2(n9875), .A(n9860), .ZN(P1_U3541) );
  AOI211_X1 U11130 ( .C1(n9863), .C2(n10172), .A(n9862), .B(n9861), .ZN(n9918)
         );
  MUX2_X1 U11131 ( .A(n9864), .B(n9918), .S(n10192), .Z(n9865) );
  OAI21_X1 U11132 ( .B1(n9921), .B2(n9875), .A(n9865), .ZN(P1_U3540) );
  INV_X1 U11133 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9869) );
  AOI211_X1 U11134 ( .C1(n9868), .C2(n10172), .A(n9867), .B(n9866), .ZN(n9922)
         );
  MUX2_X1 U11135 ( .A(n9869), .B(n9922), .S(n10192), .Z(n9870) );
  OAI21_X1 U11136 ( .B1(n9925), .B2(n9875), .A(n9870), .ZN(P1_U3538) );
  AOI211_X1 U11137 ( .C1(n9873), .C2(n10172), .A(n9872), .B(n9871), .ZN(n9926)
         );
  MUX2_X1 U11138 ( .A(n7483), .B(n9926), .S(n10192), .Z(n9874) );
  OAI21_X1 U11139 ( .B1(n9930), .B2(n9875), .A(n9874), .ZN(P1_U3536) );
  MUX2_X1 U11140 ( .A(n9876), .B(P1_REG1_REG_0__SCAN_IN), .S(n5490), .Z(
        P1_U3522) );
  INV_X1 U11141 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9878) );
  MUX2_X1 U11142 ( .A(n9878), .B(n9877), .S(n10175), .Z(n9879) );
  OAI21_X1 U11143 ( .B1(n9880), .B2(n9929), .A(n9879), .ZN(P1_U3520) );
  MUX2_X1 U11144 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9881), .S(n10175), .Z(
        P1_U3519) );
  MUX2_X1 U11145 ( .A(n9883), .B(n9882), .S(n10175), .Z(n9884) );
  OAI21_X1 U11146 ( .B1(n9885), .B2(n9929), .A(n9884), .ZN(P1_U3517) );
  INV_X1 U11147 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9887) );
  MUX2_X1 U11148 ( .A(n9887), .B(n9886), .S(n10175), .Z(n9888) );
  OAI21_X1 U11149 ( .B1(n9889), .B2(n9929), .A(n9888), .ZN(P1_U3516) );
  INV_X1 U11150 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9891) );
  MUX2_X1 U11151 ( .A(n9891), .B(n9890), .S(n10175), .Z(n9892) );
  OAI21_X1 U11152 ( .B1(n9893), .B2(n9929), .A(n9892), .ZN(P1_U3515) );
  INV_X1 U11153 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9895) );
  MUX2_X1 U11154 ( .A(n9895), .B(n9894), .S(n10175), .Z(n9896) );
  OAI21_X1 U11155 ( .B1(n9897), .B2(n9929), .A(n9896), .ZN(P1_U3514) );
  INV_X1 U11156 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9899) );
  MUX2_X1 U11157 ( .A(n9899), .B(n9898), .S(n10175), .Z(n9900) );
  OAI21_X1 U11158 ( .B1(n9901), .B2(n9929), .A(n9900), .ZN(P1_U3513) );
  INV_X1 U11159 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9903) );
  MUX2_X1 U11160 ( .A(n9903), .B(n9902), .S(n10175), .Z(n9904) );
  OAI21_X1 U11161 ( .B1(n9905), .B2(n9929), .A(n9904), .ZN(P1_U3512) );
  MUX2_X1 U11162 ( .A(n9907), .B(n9906), .S(n10175), .Z(n9908) );
  OAI21_X1 U11163 ( .B1(n9909), .B2(n9929), .A(n9908), .ZN(P1_U3511) );
  INV_X1 U11164 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9911) );
  MUX2_X1 U11165 ( .A(n9911), .B(n9910), .S(n10175), .Z(n9912) );
  OAI21_X1 U11166 ( .B1(n9913), .B2(n9929), .A(n9912), .ZN(P1_U3510) );
  INV_X1 U11167 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9915) );
  MUX2_X1 U11168 ( .A(n9915), .B(n9914), .S(n10175), .Z(n9916) );
  OAI21_X1 U11169 ( .B1(n9917), .B2(n9929), .A(n9916), .ZN(P1_U3509) );
  INV_X1 U11170 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9919) );
  MUX2_X1 U11171 ( .A(n9919), .B(n9918), .S(n10175), .Z(n9920) );
  OAI21_X1 U11172 ( .B1(n9921), .B2(n9929), .A(n9920), .ZN(P1_U3507) );
  INV_X1 U11173 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9923) );
  MUX2_X1 U11174 ( .A(n9923), .B(n9922), .S(n10175), .Z(n9924) );
  OAI21_X1 U11175 ( .B1(n9925), .B2(n9929), .A(n9924), .ZN(P1_U3501) );
  INV_X1 U11176 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9927) );
  MUX2_X1 U11177 ( .A(n9927), .B(n9926), .S(n10175), .Z(n9928) );
  OAI21_X1 U11178 ( .B1(n9930), .B2(n9929), .A(n9928), .ZN(P1_U3495) );
  NOR4_X1 U11179 ( .A1(n9932), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9931), .A4(
        P1_U3086), .ZN(n9933) );
  AOI21_X1 U11180 ( .B1(n9934), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9933), .ZN(
        n9935) );
  OAI21_X1 U11181 ( .B1(n9936), .B2(n4496), .A(n9935), .ZN(P1_U3324) );
  MUX2_X1 U11182 ( .A(n9937), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  OAI21_X1 U11183 ( .B1(n9940), .B2(n9939), .A(n9938), .ZN(n9941) );
  AOI22_X1 U11184 ( .A1(n9941), .A2(n10347), .B1(n10339), .B2(
        P2_ADDR_REG_18__SCAN_IN), .ZN(n9955) );
  INV_X1 U11185 ( .A(n9942), .ZN(n9944) );
  NAND2_X1 U11186 ( .A1(n9944), .A2(n9943), .ZN(n9952) );
  OAI21_X1 U11187 ( .B1(n9952), .B2(n9946), .A(n9945), .ZN(n9951) );
  NAND2_X1 U11188 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3151), .ZN(n9954) );
  NAND3_X1 U11189 ( .A1(n9952), .A2(n10206), .A3(n4914), .ZN(n9953) );
  OAI21_X1 U11190 ( .B1(n9957), .B2(n7662), .A(n9956), .ZN(n9967) );
  INV_X1 U11191 ( .A(n9958), .ZN(n9961) );
  AOI21_X1 U11192 ( .B1(n9961), .B2(n9960), .A(n9959), .ZN(n9962) );
  OAI21_X1 U11193 ( .B1(n9964), .B2(n9963), .A(n9962), .ZN(n9965) );
  AOI21_X1 U11194 ( .B1(n9967), .B2(n9966), .A(n9965), .ZN(n9968) );
  OAI21_X1 U11195 ( .B1(n9970), .B2(n9969), .A(n9968), .ZN(P1_U3224) );
  OAI211_X1 U11196 ( .C1(n5011), .C2(n10168), .A(n9972), .B(n9971), .ZN(n9973)
         );
  AOI21_X1 U11197 ( .B1(n9974), .B2(n10172), .A(n9973), .ZN(n9983) );
  AOI22_X1 U11198 ( .A1(n10192), .A2(n9983), .B1(n9975), .B2(n5490), .ZN(
        P1_U3539) );
  OAI211_X1 U11199 ( .C1(n9978), .C2(n10168), .A(n9977), .B(n9976), .ZN(n9979)
         );
  AOI21_X1 U11200 ( .B1(n9980), .B2(n10172), .A(n9979), .ZN(n9985) );
  AOI22_X1 U11201 ( .A1(n10192), .A2(n9985), .B1(n9981), .B2(n5490), .ZN(
        P1_U3537) );
  INV_X1 U11202 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9982) );
  AOI22_X1 U11203 ( .A1(n10175), .A2(n9983), .B1(n9982), .B2(n10173), .ZN(
        P1_U3504) );
  INV_X1 U11204 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9984) );
  AOI22_X1 U11205 ( .A1(n10175), .A2(n9985), .B1(n9984), .B2(n10173), .ZN(
        P1_U3498) );
  XNOR2_X1 U11206 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11207 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11208 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9986) );
  AOI21_X1 U11209 ( .B1(n9987), .B2(n9986), .A(n5454), .ZN(n10009) );
  OAI21_X1 U11210 ( .B1(n9987), .B2(P1_REG1_REG_0__SCAN_IN), .A(n10009), .ZN(
        n9988) );
  XOR2_X1 U11211 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9988), .Z(n9992) );
  AOI22_X1 U11212 ( .A1(n10026), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9990) );
  OAI21_X1 U11213 ( .B1(n9992), .B2(n9991), .A(n9990), .ZN(P1_U3243) );
  AOI22_X1 U11214 ( .A1(n10026), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n10011) );
  AOI211_X1 U11215 ( .C1(n9995), .C2(n9994), .A(n4587), .B(n9993), .ZN(n10000)
         );
  AOI211_X1 U11216 ( .C1(n9998), .C2(n9997), .A(n9996), .B(n10018), .ZN(n9999)
         );
  AOI211_X1 U11217 ( .C1(n10025), .C2(n10001), .A(n10000), .B(n9999), .ZN(
        n10010) );
  INV_X1 U11218 ( .A(n10002), .ZN(n10004) );
  MUX2_X1 U11219 ( .A(n10004), .B(n10003), .S(n5456), .Z(n10006) );
  NAND2_X1 U11220 ( .A1(n10006), .A2(n10005), .ZN(n10008) );
  OAI211_X1 U11221 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n10009), .A(n10008), .B(
        P1_U3973), .ZN(n10028) );
  NAND3_X1 U11222 ( .A1(n10011), .A2(n10010), .A3(n10028), .ZN(P1_U3245) );
  OAI21_X1 U11223 ( .B1(n10014), .B2(n10013), .A(n10012), .ZN(n10015) );
  INV_X1 U11224 ( .A(n10015), .ZN(n10016) );
  AND2_X1 U11225 ( .A1(n10017), .A2(n10016), .ZN(n10023) );
  AOI211_X1 U11226 ( .C1(n10021), .C2(n10020), .A(n10019), .B(n10018), .ZN(
        n10022) );
  AOI211_X1 U11227 ( .C1(n10025), .C2(n10024), .A(n10023), .B(n10022), .ZN(
        n10030) );
  NAND2_X1 U11228 ( .A1(n10026), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n10027) );
  NAND4_X1 U11229 ( .A1(n10030), .A2(n10029), .A3(n10028), .A4(n10027), .ZN(
        P1_U3247) );
  INV_X1 U11230 ( .A(n10031), .ZN(n10154) );
  XNOR2_X1 U11231 ( .A(n10032), .B(n10033), .ZN(n10149) );
  NAND3_X1 U11232 ( .A1(n10035), .A2(n10034), .A3(n10033), .ZN(n10037) );
  AOI21_X1 U11233 ( .B1(n10038), .B2(n10037), .A(n10036), .ZN(n10039) );
  AOI211_X1 U11234 ( .C1(n10154), .C2(n10149), .A(n10040), .B(n10039), .ZN(
        n10146) );
  AOI222_X1 U11235 ( .A1(n10044), .A2(n10060), .B1(P1_REG2_REG_7__SCAN_IN), 
        .B2(n10043), .C1(n10042), .C2(n10041), .ZN(n10051) );
  NOR2_X1 U11236 ( .A1(n10070), .A2(n10045), .ZN(n10049) );
  OAI211_X1 U11237 ( .C1(n10047), .C2(n10145), .A(n10046), .B(n10063), .ZN(
        n10144) );
  INV_X1 U11238 ( .A(n10144), .ZN(n10048) );
  AOI22_X1 U11239 ( .A1(n10149), .A2(n10049), .B1(n10066), .B2(n10048), .ZN(
        n10050) );
  OAI211_X1 U11240 ( .C1(n10070), .C2(n10146), .A(n10051), .B(n10050), .ZN(
        P1_U3286) );
  XNOR2_X1 U11241 ( .A(n10052), .B(n10062), .ZN(n10055) );
  AOI21_X1 U11242 ( .B1(n10055), .B2(n10054), .A(n10053), .ZN(n10119) );
  INV_X1 U11243 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10057) );
  OAI22_X1 U11244 ( .A1(n10058), .A2(n10057), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n10056), .ZN(n10059) );
  AOI21_X1 U11245 ( .B1(n10060), .B2(n5515), .A(n10059), .ZN(n10069) );
  XNOR2_X1 U11246 ( .A(n10062), .B(n10061), .ZN(n10122) );
  OAI211_X1 U11247 ( .C1(n10064), .C2(n10118), .A(n7311), .B(n10063), .ZN(
        n10117) );
  INV_X1 U11248 ( .A(n10117), .ZN(n10065) );
  AOI22_X1 U11249 ( .A1(n10122), .A2(n10067), .B1(n10066), .B2(n10065), .ZN(
        n10068) );
  OAI211_X1 U11250 ( .C1(n10070), .C2(n10119), .A(n10069), .B(n10068), .ZN(
        P1_U3290) );
  INV_X1 U11251 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10071) );
  NOR2_X1 U11252 ( .A1(n10102), .A2(n10071), .ZN(P1_U3294) );
  INV_X1 U11253 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10072) );
  NOR2_X1 U11254 ( .A1(n10102), .A2(n10072), .ZN(P1_U3295) );
  INV_X1 U11255 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10073) );
  NOR2_X1 U11256 ( .A1(n10102), .A2(n10073), .ZN(P1_U3296) );
  INV_X1 U11257 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10074) );
  NOR2_X1 U11258 ( .A1(n10084), .A2(n10074), .ZN(P1_U3297) );
  INV_X1 U11259 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10075) );
  NOR2_X1 U11260 ( .A1(n10084), .A2(n10075), .ZN(P1_U3298) );
  INV_X1 U11261 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10076) );
  NOR2_X1 U11262 ( .A1(n10084), .A2(n10076), .ZN(P1_U3299) );
  NOR2_X1 U11263 ( .A1(n10084), .A2(n10077), .ZN(P1_U3300) );
  NOR2_X1 U11264 ( .A1(n10084), .A2(n10078), .ZN(P1_U3301) );
  INV_X1 U11265 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10079) );
  NOR2_X1 U11266 ( .A1(n10084), .A2(n10079), .ZN(P1_U3302) );
  INV_X1 U11267 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10080) );
  NOR2_X1 U11268 ( .A1(n10084), .A2(n10080), .ZN(P1_U3303) );
  INV_X1 U11269 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10081) );
  NOR2_X1 U11270 ( .A1(n10084), .A2(n10081), .ZN(P1_U3304) );
  INV_X1 U11271 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10082) );
  NOR2_X1 U11272 ( .A1(n10084), .A2(n10082), .ZN(P1_U3305) );
  INV_X1 U11273 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10083) );
  NOR2_X1 U11274 ( .A1(n10084), .A2(n10083), .ZN(P1_U3306) );
  INV_X1 U11275 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10085) );
  NOR2_X1 U11276 ( .A1(n10102), .A2(n10085), .ZN(P1_U3307) );
  INV_X1 U11277 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10086) );
  NOR2_X1 U11278 ( .A1(n10102), .A2(n10086), .ZN(P1_U3308) );
  INV_X1 U11279 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10087) );
  NOR2_X1 U11280 ( .A1(n10102), .A2(n10087), .ZN(P1_U3309) );
  INV_X1 U11281 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10088) );
  NOR2_X1 U11282 ( .A1(n10102), .A2(n10088), .ZN(P1_U3310) );
  NOR2_X1 U11283 ( .A1(n10102), .A2(n10089), .ZN(P1_U3311) );
  INV_X1 U11284 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10090) );
  NOR2_X1 U11285 ( .A1(n10102), .A2(n10090), .ZN(P1_U3312) );
  INV_X1 U11286 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10091) );
  NOR2_X1 U11287 ( .A1(n10102), .A2(n10091), .ZN(P1_U3313) );
  INV_X1 U11288 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10092) );
  NOR2_X1 U11289 ( .A1(n10102), .A2(n10092), .ZN(P1_U3314) );
  INV_X1 U11290 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10093) );
  NOR2_X1 U11291 ( .A1(n10102), .A2(n10093), .ZN(P1_U3315) );
  NOR2_X1 U11292 ( .A1(n10102), .A2(n10094), .ZN(P1_U3316) );
  INV_X1 U11293 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10095) );
  NOR2_X1 U11294 ( .A1(n10102), .A2(n10095), .ZN(P1_U3317) );
  INV_X1 U11295 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10096) );
  NOR2_X1 U11296 ( .A1(n10102), .A2(n10096), .ZN(P1_U3318) );
  INV_X1 U11297 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10097) );
  NOR2_X1 U11298 ( .A1(n10102), .A2(n10097), .ZN(P1_U3319) );
  INV_X1 U11299 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10098) );
  NOR2_X1 U11300 ( .A1(n10102), .A2(n10098), .ZN(P1_U3320) );
  INV_X1 U11301 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10099) );
  NOR2_X1 U11302 ( .A1(n10102), .A2(n10099), .ZN(P1_U3321) );
  INV_X1 U11303 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10100) );
  NOR2_X1 U11304 ( .A1(n10102), .A2(n10100), .ZN(P1_U3322) );
  INV_X1 U11305 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10101) );
  NOR2_X1 U11306 ( .A1(n10102), .A2(n10101), .ZN(P1_U3323) );
  OAI21_X1 U11307 ( .B1(n10104), .B2(n10168), .A(n10103), .ZN(n10107) );
  INV_X1 U11308 ( .A(n10105), .ZN(n10106) );
  AOI211_X1 U11309 ( .C1(n10108), .C2(n10172), .A(n10107), .B(n10106), .ZN(
        n10177) );
  INV_X1 U11310 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10109) );
  AOI22_X1 U11311 ( .A1(n10175), .A2(n10177), .B1(n10109), .B2(n10173), .ZN(
        P1_U3456) );
  INV_X1 U11312 ( .A(n10110), .ZN(n10111) );
  OAI21_X1 U11313 ( .B1(n5507), .B2(n10168), .A(n10111), .ZN(n10114) );
  INV_X1 U11314 ( .A(n10112), .ZN(n10113) );
  AOI211_X1 U11315 ( .C1(n10172), .C2(n10115), .A(n10114), .B(n10113), .ZN(
        n10179) );
  INV_X1 U11316 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10116) );
  AOI22_X1 U11317 ( .A1(n10175), .A2(n10179), .B1(n10116), .B2(n10173), .ZN(
        P1_U3459) );
  OAI21_X1 U11318 ( .B1(n10118), .B2(n10168), .A(n10117), .ZN(n10121) );
  INV_X1 U11319 ( .A(n10119), .ZN(n10120) );
  AOI211_X1 U11320 ( .C1(n10172), .C2(n10122), .A(n10121), .B(n10120), .ZN(
        n10180) );
  INV_X1 U11321 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10123) );
  AOI22_X1 U11322 ( .A1(n10175), .A2(n10180), .B1(n10123), .B2(n10173), .ZN(
        P1_U3462) );
  OAI21_X1 U11323 ( .B1(n10125), .B2(n10168), .A(n10124), .ZN(n10127) );
  AOI211_X1 U11324 ( .C1(n10172), .C2(n10128), .A(n10127), .B(n10126), .ZN(
        n10182) );
  INV_X1 U11325 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10129) );
  AOI22_X1 U11326 ( .A1(n10175), .A2(n10182), .B1(n10129), .B2(n10173), .ZN(
        P1_U3465) );
  AND2_X1 U11327 ( .A1(n10130), .A2(n10172), .ZN(n10134) );
  OAI21_X1 U11328 ( .B1(n10132), .B2(n10168), .A(n10131), .ZN(n10133) );
  NOR3_X1 U11329 ( .A1(n10135), .A2(n10134), .A3(n10133), .ZN(n10184) );
  INV_X1 U11330 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10136) );
  AOI22_X1 U11331 ( .A1(n10175), .A2(n10184), .B1(n10136), .B2(n10173), .ZN(
        P1_U3468) );
  OAI21_X1 U11332 ( .B1(n10138), .B2(n10168), .A(n10137), .ZN(n10140) );
  AOI211_X1 U11333 ( .C1(n10172), .C2(n10141), .A(n10140), .B(n10139), .ZN(
        n10185) );
  INV_X1 U11334 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10142) );
  AOI22_X1 U11335 ( .A1(n10175), .A2(n10185), .B1(n10142), .B2(n10173), .ZN(
        P1_U3471) );
  INV_X1 U11336 ( .A(n10143), .ZN(n10153) );
  OAI21_X1 U11337 ( .B1(n10145), .B2(n10168), .A(n10144), .ZN(n10148) );
  INV_X1 U11338 ( .A(n10146), .ZN(n10147) );
  AOI211_X1 U11339 ( .C1(n10153), .C2(n10149), .A(n10148), .B(n10147), .ZN(
        n10186) );
  INV_X1 U11340 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10150) );
  AOI22_X1 U11341 ( .A1(n10175), .A2(n10186), .B1(n10150), .B2(n10173), .ZN(
        P1_U3474) );
  OAI21_X1 U11342 ( .B1(n5006), .B2(n10168), .A(n10151), .ZN(n10157) );
  OAI21_X1 U11343 ( .B1(n10154), .B2(n10153), .A(n10152), .ZN(n10155) );
  INV_X1 U11344 ( .A(n10155), .ZN(n10156) );
  NOR3_X1 U11345 ( .A1(n10158), .A2(n10157), .A3(n10156), .ZN(n10188) );
  INV_X1 U11346 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10159) );
  AOI22_X1 U11347 ( .A1(n10175), .A2(n10188), .B1(n10159), .B2(n10173), .ZN(
        P1_U3477) );
  OAI21_X1 U11348 ( .B1(n10161), .B2(n10168), .A(n10160), .ZN(n10163) );
  AOI211_X1 U11349 ( .C1(n10172), .C2(n10164), .A(n10163), .B(n10162), .ZN(
        n10190) );
  AOI22_X1 U11350 ( .A1(n10175), .A2(n10190), .B1(n10165), .B2(n10173), .ZN(
        P1_U3480) );
  OAI211_X1 U11351 ( .C1(n10169), .C2(n10168), .A(n10167), .B(n10166), .ZN(
        n10170) );
  AOI21_X1 U11352 ( .B1(n10172), .B2(n10171), .A(n10170), .ZN(n10191) );
  INV_X1 U11353 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10174) );
  AOI22_X1 U11354 ( .A1(n10175), .A2(n10191), .B1(n10174), .B2(n10173), .ZN(
        P1_U3483) );
  AOI22_X1 U11355 ( .A1(n10192), .A2(n10177), .B1(n10176), .B2(n5490), .ZN(
        P1_U3523) );
  INV_X1 U11356 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10178) );
  AOI22_X1 U11357 ( .A1(n10192), .A2(n10179), .B1(n10178), .B2(n5490), .ZN(
        P1_U3524) );
  AOI22_X1 U11358 ( .A1(n10192), .A2(n10180), .B1(n6405), .B2(n5490), .ZN(
        P1_U3525) );
  INV_X1 U11359 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10181) );
  AOI22_X1 U11360 ( .A1(n10192), .A2(n10182), .B1(n10181), .B2(n5490), .ZN(
        P1_U3526) );
  INV_X1 U11361 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10183) );
  AOI22_X1 U11362 ( .A1(n10192), .A2(n10184), .B1(n10183), .B2(n5490), .ZN(
        P1_U3527) );
  AOI22_X1 U11363 ( .A1(n10192), .A2(n10185), .B1(n6409), .B2(n5490), .ZN(
        P1_U3528) );
  AOI22_X1 U11364 ( .A1(n10192), .A2(n10186), .B1(n6410), .B2(n5490), .ZN(
        P1_U3529) );
  INV_X1 U11365 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10187) );
  AOI22_X1 U11366 ( .A1(n10192), .A2(n10188), .B1(n10187), .B2(n5490), .ZN(
        P1_U3530) );
  AOI22_X1 U11367 ( .A1(n10192), .A2(n10190), .B1(n10189), .B2(n5490), .ZN(
        P1_U3531) );
  AOI22_X1 U11368 ( .A1(n10192), .A2(n10191), .B1(n6786), .B2(n5490), .ZN(
        P1_U3532) );
  INV_X1 U11369 ( .A(n10193), .ZN(n10202) );
  XNOR2_X1 U11370 ( .A(n10195), .B(n10194), .ZN(n10198) );
  XOR2_X1 U11371 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n10196), .Z(n10197) );
  AOI22_X1 U11372 ( .A1(n10348), .A2(n10198), .B1(n10347), .B2(n10197), .ZN(
        n10199) );
  OAI21_X1 U11373 ( .B1(n10451), .B2(n10200), .A(n10199), .ZN(n10201) );
  AOI21_X1 U11374 ( .B1(n10202), .B2(n10340), .A(n10201), .ZN(n10208) );
  XOR2_X1 U11375 ( .A(n10204), .B(n10203), .Z(n10205) );
  NAND2_X1 U11376 ( .A1(n10206), .A2(n10205), .ZN(n10207) );
  OAI211_X1 U11377 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n5981), .A(n10208), .B(
        n10207), .ZN(P2_U3183) );
  AOI22_X1 U11378 ( .A1(n10209), .A2(n10340), .B1(n10339), .B2(
        P2_ADDR_REG_9__SCAN_IN), .ZN(n10224) );
  OAI21_X1 U11379 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n10211), .A(n10210), .ZN(
        n10215) );
  OAI21_X1 U11380 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n10213), .A(n10212), .ZN(
        n10214) );
  AOI22_X1 U11381 ( .A1(n10215), .A2(n10348), .B1(n10214), .B2(n10347), .ZN(
        n10223) );
  INV_X1 U11382 ( .A(n10216), .ZN(n10222) );
  AOI21_X1 U11383 ( .B1(n10219), .B2(n10218), .A(n10217), .ZN(n10220) );
  OR2_X1 U11384 ( .A1(n10354), .A2(n10220), .ZN(n10221) );
  NAND4_X1 U11385 ( .A1(n10224), .A2(n10223), .A3(n10222), .A4(n10221), .ZN(
        P2_U3191) );
  AOI22_X1 U11386 ( .A1(n10225), .A2(n10340), .B1(n10339), .B2(
        P2_ADDR_REG_10__SCAN_IN), .ZN(n10240) );
  OAI21_X1 U11387 ( .B1(n10228), .B2(n10227), .A(n10226), .ZN(n10233) );
  OAI21_X1 U11388 ( .B1(n10231), .B2(n10230), .A(n10229), .ZN(n10232) );
  AOI22_X1 U11389 ( .A1(n10233), .A2(n10348), .B1(n10232), .B2(n10347), .ZN(
        n10239) );
  AOI21_X1 U11390 ( .B1(n4530), .B2(n10235), .A(n10234), .ZN(n10236) );
  OR2_X1 U11391 ( .A1(n10236), .A2(n10354), .ZN(n10237) );
  NAND4_X1 U11392 ( .A1(n10240), .A2(n10239), .A3(n10238), .A4(n10237), .ZN(
        P2_U3192) );
  AOI22_X1 U11393 ( .A1(n10339), .A2(P2_ADDR_REG_11__SCAN_IN), .B1(n10340), 
        .B2(n10241), .ZN(n10256) );
  OAI21_X1 U11394 ( .B1(n10243), .B2(P2_REG2_REG_11__SCAN_IN), .A(n10242), 
        .ZN(n10247) );
  OAI21_X1 U11395 ( .B1(n10245), .B2(P2_REG1_REG_11__SCAN_IN), .A(n10244), 
        .ZN(n10246) );
  AOI22_X1 U11396 ( .A1(n10247), .A2(n10348), .B1(n10246), .B2(n10347), .ZN(
        n10255) );
  INV_X1 U11397 ( .A(n10248), .ZN(n10254) );
  AOI21_X1 U11398 ( .B1(n10251), .B2(n10250), .A(n10249), .ZN(n10252) );
  OR2_X1 U11399 ( .A1(n10252), .A2(n10354), .ZN(n10253) );
  NAND4_X1 U11400 ( .A1(n10256), .A2(n10255), .A3(n10254), .A4(n10253), .ZN(
        P2_U3193) );
  AOI22_X1 U11401 ( .A1(n10257), .A2(n10340), .B1(n10339), .B2(
        P2_ADDR_REG_12__SCAN_IN), .ZN(n10273) );
  OAI21_X1 U11402 ( .B1(n10260), .B2(n10259), .A(n10258), .ZN(n10265) );
  OAI21_X1 U11403 ( .B1(n10263), .B2(n10262), .A(n10261), .ZN(n10264) );
  AOI22_X1 U11404 ( .A1(n10265), .A2(n10348), .B1(n10264), .B2(n10347), .ZN(
        n10272) );
  INV_X1 U11405 ( .A(n10266), .ZN(n10271) );
  AOI21_X1 U11406 ( .B1(n10268), .B2(n10267), .A(n4884), .ZN(n10269) );
  OR2_X1 U11407 ( .A1(n10269), .A2(n10354), .ZN(n10270) );
  NAND4_X1 U11408 ( .A1(n10273), .A2(n10272), .A3(n10271), .A4(n10270), .ZN(
        P2_U3194) );
  AOI22_X1 U11409 ( .A1(n10274), .A2(n10340), .B1(n10339), .B2(
        P2_ADDR_REG_13__SCAN_IN), .ZN(n10289) );
  OAI21_X1 U11410 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n10276), .A(n10275), 
        .ZN(n10280) );
  OAI21_X1 U11411 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n10278), .A(n10277), 
        .ZN(n10279) );
  AOI22_X1 U11412 ( .A1(n10280), .A2(n10348), .B1(n10347), .B2(n10279), .ZN(
        n10288) );
  INV_X1 U11413 ( .A(n10281), .ZN(n10287) );
  AOI21_X1 U11414 ( .B1(n10284), .B2(n10283), .A(n10282), .ZN(n10285) );
  OR2_X1 U11415 ( .A1(n10285), .A2(n10354), .ZN(n10286) );
  NAND4_X1 U11416 ( .A1(n10289), .A2(n10288), .A3(n10287), .A4(n10286), .ZN(
        P2_U3195) );
  AOI22_X1 U11417 ( .A1(n10290), .A2(n10340), .B1(P2_ADDR_REG_14__SCAN_IN), 
        .B2(n10339), .ZN(n10306) );
  OAI21_X1 U11418 ( .B1(n10293), .B2(n10292), .A(n10291), .ZN(n10298) );
  OAI21_X1 U11419 ( .B1(n10296), .B2(n10295), .A(n10294), .ZN(n10297) );
  AOI22_X1 U11420 ( .A1(n10298), .A2(n10348), .B1(n10347), .B2(n10297), .ZN(
        n10305) );
  AOI21_X1 U11421 ( .B1(n10301), .B2(n10300), .A(n10299), .ZN(n10302) );
  OR2_X1 U11422 ( .A1(n10302), .A2(n10354), .ZN(n10303) );
  NAND4_X1 U11423 ( .A1(n10306), .A2(n10305), .A3(n10304), .A4(n10303), .ZN(
        P2_U3196) );
  AOI22_X1 U11424 ( .A1(n10307), .A2(n10340), .B1(P2_ADDR_REG_15__SCAN_IN), 
        .B2(n10339), .ZN(n10321) );
  OAI21_X1 U11425 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n10309), .A(n10308), 
        .ZN(n10313) );
  OAI21_X1 U11426 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n10311), .A(n10310), 
        .ZN(n10312) );
  AOI22_X1 U11427 ( .A1(n10313), .A2(n10348), .B1(n10347), .B2(n10312), .ZN(
        n10320) );
  INV_X1 U11428 ( .A(n10314), .ZN(n10319) );
  AOI21_X1 U11429 ( .B1(n10316), .B2(n10315), .A(n4576), .ZN(n10317) );
  OR2_X1 U11430 ( .A1(n10317), .A2(n10354), .ZN(n10318) );
  NAND4_X1 U11431 ( .A1(n10321), .A2(n10320), .A3(n10319), .A4(n10318), .ZN(
        P2_U3197) );
  AOI22_X1 U11432 ( .A1(n10322), .A2(n10340), .B1(n10339), .B2(
        P2_ADDR_REG_16__SCAN_IN), .ZN(n10338) );
  OAI21_X1 U11433 ( .B1(n10325), .B2(n10324), .A(n10323), .ZN(n10330) );
  OAI21_X1 U11434 ( .B1(n10328), .B2(n10327), .A(n10326), .ZN(n10329) );
  AOI22_X1 U11435 ( .A1(n10330), .A2(n10348), .B1(n10347), .B2(n10329), .ZN(
        n10337) );
  AOI21_X1 U11436 ( .B1(n10333), .B2(n10332), .A(n10331), .ZN(n10334) );
  OR2_X1 U11437 ( .A1(n10334), .A2(n10354), .ZN(n10335) );
  NAND4_X1 U11438 ( .A1(n10338), .A2(n10337), .A3(n10336), .A4(n10335), .ZN(
        P2_U3198) );
  AOI22_X1 U11439 ( .A1(n10341), .A2(n10340), .B1(n10339), .B2(
        P2_ADDR_REG_17__SCAN_IN), .ZN(n10359) );
  OAI21_X1 U11440 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n10343), .A(n10342), 
        .ZN(n10349) );
  OAI21_X1 U11441 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n10345), .A(n10344), 
        .ZN(n10346) );
  AOI22_X1 U11442 ( .A1(n10349), .A2(n10348), .B1(n10347), .B2(n10346), .ZN(
        n10358) );
  NAND2_X1 U11443 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3151), .ZN(n10357)
         );
  AOI21_X1 U11444 ( .B1(n10353), .B2(n10352), .A(n10351), .ZN(n10355) );
  OR2_X1 U11445 ( .A1(n10355), .A2(n10354), .ZN(n10356) );
  NAND4_X1 U11446 ( .A1(n10359), .A2(n10358), .A3(n10357), .A4(n10356), .ZN(
        P2_U3199) );
  AOI21_X1 U11447 ( .B1(n10362), .B2(n10361), .A(n10360), .ZN(n10363) );
  OAI222_X1 U11448 ( .A1(n10373), .A2(n10366), .B1(n10365), .B2(n10364), .C1(
        n10381), .C2(n10363), .ZN(n10367) );
  INV_X1 U11449 ( .A(n10367), .ZN(n10368) );
  OAI21_X1 U11450 ( .B1(n4495), .B2(n10369), .A(n10368), .ZN(P2_U3229) );
  OAI22_X1 U11451 ( .A1(n10373), .A2(n10372), .B1(n10371), .B2(n10370), .ZN(
        n10376) );
  INV_X1 U11452 ( .A(n10374), .ZN(n10375) );
  AOI211_X1 U11453 ( .C1(n10378), .C2(n10377), .A(n10376), .B(n10375), .ZN(
        n10379) );
  AOI22_X1 U11454 ( .A1(n10381), .A2(n10380), .B1(n10379), .B2(n4495), .ZN(
        P2_U3231) );
  INV_X1 U11455 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10387) );
  INV_X1 U11456 ( .A(n10382), .ZN(n10386) );
  OAI22_X1 U11457 ( .A1(n10384), .A2(n10420), .B1(n10383), .B2(n10418), .ZN(
        n10385) );
  NOR2_X1 U11458 ( .A1(n10386), .A2(n10385), .ZN(n10433) );
  AOI22_X1 U11459 ( .A1(n10432), .A2(n10387), .B1(n10433), .B2(n10430), .ZN(
        P2_U3393) );
  INV_X1 U11460 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10389) );
  AOI22_X1 U11461 ( .A1(n10432), .A2(n10389), .B1(n10388), .B2(n10430), .ZN(
        P2_U3396) );
  AOI22_X1 U11462 ( .A1(n10391), .A2(n10408), .B1(n10429), .B2(n10390), .ZN(
        n10392) );
  AND2_X1 U11463 ( .A1(n10393), .A2(n10392), .ZN(n10435) );
  AOI22_X1 U11464 ( .A1(n10432), .A2(n6003), .B1(n10435), .B2(n10430), .ZN(
        P2_U3399) );
  AOI22_X1 U11465 ( .A1(n10395), .A2(n6328), .B1(n10429), .B2(n10394), .ZN(
        n10396) );
  AND2_X1 U11466 ( .A1(n10397), .A2(n10396), .ZN(n10436) );
  AOI22_X1 U11467 ( .A1(n10432), .A2(n6038), .B1(n10436), .B2(n10430), .ZN(
        P2_U3405) );
  INV_X1 U11468 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10402) );
  AOI22_X1 U11469 ( .A1(n10399), .A2(n10408), .B1(n10429), .B2(n10398), .ZN(
        n10400) );
  AND2_X1 U11470 ( .A1(n10401), .A2(n10400), .ZN(n10437) );
  AOI22_X1 U11471 ( .A1(n10432), .A2(n10402), .B1(n10437), .B2(n10430), .ZN(
        P2_U3408) );
  NOR2_X1 U11472 ( .A1(n10403), .A2(n10420), .ZN(n10405) );
  AOI211_X1 U11473 ( .C1(n10429), .C2(n10406), .A(n10405), .B(n10404), .ZN(
        n10439) );
  AOI22_X1 U11474 ( .A1(n10432), .A2(n6051), .B1(n10439), .B2(n10430), .ZN(
        P2_U3411) );
  INV_X1 U11475 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10412) );
  AOI22_X1 U11476 ( .A1(n10409), .A2(n10408), .B1(n10429), .B2(n10407), .ZN(
        n10410) );
  AND2_X1 U11477 ( .A1(n10411), .A2(n10410), .ZN(n10440) );
  AOI22_X1 U11478 ( .A1(n10432), .A2(n10412), .B1(n10440), .B2(n10430), .ZN(
        P2_U3414) );
  INV_X1 U11479 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10417) );
  NOR2_X1 U11480 ( .A1(n10413), .A2(n10420), .ZN(n10415) );
  AOI211_X1 U11481 ( .C1(n10429), .C2(n10416), .A(n10415), .B(n10414), .ZN(
        n10441) );
  AOI22_X1 U11482 ( .A1(n10432), .A2(n10417), .B1(n10441), .B2(n10430), .ZN(
        P2_U3417) );
  OAI22_X1 U11483 ( .A1(n10421), .A2(n10420), .B1(n10419), .B2(n10418), .ZN(
        n10422) );
  NOR2_X1 U11484 ( .A1(n10423), .A2(n10422), .ZN(n10443) );
  AOI22_X1 U11485 ( .A1(n10432), .A2(n6092), .B1(n10443), .B2(n10430), .ZN(
        P2_U3420) );
  INV_X1 U11486 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10431) );
  NOR2_X1 U11487 ( .A1(n10425), .A2(n10424), .ZN(n10427) );
  AOI211_X1 U11488 ( .C1(n10429), .C2(n10428), .A(n10427), .B(n10426), .ZN(
        n10445) );
  AOI22_X1 U11489 ( .A1(n10432), .A2(n10431), .B1(n10445), .B2(n10430), .ZN(
        P2_U3423) );
  AOI22_X1 U11490 ( .A1(n10446), .A2(n10433), .B1(n5925), .B2(n10444), .ZN(
        P2_U3460) );
  INV_X1 U11491 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10434) );
  AOI22_X1 U11492 ( .A1(n10446), .A2(n10435), .B1(n10434), .B2(n10444), .ZN(
        P2_U3462) );
  AOI22_X1 U11493 ( .A1(n10446), .A2(n10436), .B1(n5929), .B2(n10444), .ZN(
        P2_U3464) );
  AOI22_X1 U11494 ( .A1(n10446), .A2(n10437), .B1(n6023), .B2(n10444), .ZN(
        P2_U3465) );
  AOI22_X1 U11495 ( .A1(n10446), .A2(n10439), .B1(n10438), .B2(n10444), .ZN(
        P2_U3466) );
  AOI22_X1 U11496 ( .A1(n10446), .A2(n10440), .B1(n6065), .B2(n10444), .ZN(
        P2_U3467) );
  AOI22_X1 U11497 ( .A1(n10446), .A2(n10441), .B1(n6081), .B2(n10444), .ZN(
        P2_U3468) );
  AOI22_X1 U11498 ( .A1(n10446), .A2(n10443), .B1(n10442), .B2(n10444), .ZN(
        P2_U3469) );
  AOI22_X1 U11499 ( .A1(n10446), .A2(n10445), .B1(n6101), .B2(n10444), .ZN(
        P2_U3470) );
  OAI222_X1 U11500 ( .A1(n10451), .A2(n10450), .B1(n10451), .B2(n10449), .C1(
        n10448), .C2(n10447), .ZN(ADD_1068_U5) );
  XOR2_X1 U11501 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI21_X1 U11502 ( .B1(n10454), .B2(n10453), .A(n10452), .ZN(n10455) );
  XNOR2_X1 U11503 ( .A(n10455), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1068_U55)
         );
  OAI21_X1 U11504 ( .B1(n10458), .B2(n10457), .A(n10456), .ZN(ADD_1068_U56) );
  OAI21_X1 U11505 ( .B1(n10461), .B2(n10460), .A(n10459), .ZN(ADD_1068_U57) );
  OAI21_X1 U11506 ( .B1(n10464), .B2(n10463), .A(n10462), .ZN(ADD_1068_U58) );
  OAI21_X1 U11507 ( .B1(n10467), .B2(n10466), .A(n10465), .ZN(ADD_1068_U59) );
  OAI21_X1 U11508 ( .B1(n10470), .B2(n10469), .A(n10468), .ZN(ADD_1068_U60) );
  OAI21_X1 U11509 ( .B1(n10473), .B2(n10472), .A(n10471), .ZN(ADD_1068_U61) );
  OAI21_X1 U11510 ( .B1(n10476), .B2(n10475), .A(n10474), .ZN(ADD_1068_U62) );
  OAI21_X1 U11511 ( .B1(n10479), .B2(n10478), .A(n10477), .ZN(ADD_1068_U63) );
  OAI21_X1 U11512 ( .B1(n10482), .B2(n10481), .A(n10480), .ZN(ADD_1068_U50) );
  OAI21_X1 U11513 ( .B1(n10485), .B2(n10484), .A(n10483), .ZN(ADD_1068_U51) );
  OAI21_X1 U11514 ( .B1(n10488), .B2(n10487), .A(n10486), .ZN(ADD_1068_U47) );
  OAI21_X1 U11515 ( .B1(n10491), .B2(n10490), .A(n10489), .ZN(ADD_1068_U49) );
  OAI21_X1 U11516 ( .B1(n10494), .B2(n10493), .A(n10492), .ZN(ADD_1068_U48) );
  AOI21_X1 U11517 ( .B1(n10497), .B2(n10496), .A(n10495), .ZN(ADD_1068_U54) );
  AOI21_X1 U11518 ( .B1(n10500), .B2(n10499), .A(n10498), .ZN(ADD_1068_U53) );
  OAI21_X1 U11519 ( .B1(n10503), .B2(n10502), .A(n10501), .ZN(ADD_1068_U52) );
  NAND2_X2 U6090 ( .A1(n5127), .A2(n4835), .ZN(n5173) );
  CLKBUF_X2 U5020 ( .A(n7040), .Z(n8727) );
  CLKBUF_X1 U5033 ( .A(n5982), .Z(n6315) );
  CLKBUF_X2 U5052 ( .A(n5922), .Z(n4492) );
  CLKBUF_X2 U5057 ( .A(n5503), .Z(n7785) );
  CLKBUF_X1 U5118 ( .A(n5079), .Z(n5672) );
  CLKBUF_X1 U5134 ( .A(n6631), .Z(n4501) );
  CLKBUF_X1 U5175 ( .A(n5124), .Z(n4835) );
endmodule

